
module mult ( a, b, c );
  input [63:0] a;
  input [63:0] b;
  output [127:0] c;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
         n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
         n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
         n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873,
         n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
         n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889,
         n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
         n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905,
         n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
         n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
         n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
         n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937,
         n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
         n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
         n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
         n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
         n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985,
         n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
         n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
         n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009,
         n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017,
         n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025,
         n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
         n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041,
         n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049,
         n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057,
         n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065,
         n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
         n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081,
         n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089,
         n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
         n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105,
         n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113,
         n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121,
         n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129,
         n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137,
         n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145,
         n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153,
         n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161,
         n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169,
         n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177,
         n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185,
         n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193,
         n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201,
         n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209,
         n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217,
         n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225,
         n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233,
         n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241,
         n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249,
         n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257,
         n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265,
         n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273,
         n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281,
         n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289,
         n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297,
         n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305,
         n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313,
         n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321,
         n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329,
         n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337,
         n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345,
         n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353,
         n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361,
         n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369,
         n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377,
         n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385,
         n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393,
         n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401,
         n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409,
         n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417,
         n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425,
         n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433,
         n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441,
         n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449,
         n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457,
         n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465,
         n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473,
         n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481,
         n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489,
         n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497,
         n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505,
         n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513,
         n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521,
         n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529,
         n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537,
         n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545,
         n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553,
         n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561,
         n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569,
         n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577,
         n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585,
         n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593,
         n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601,
         n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609,
         n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617,
         n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625,
         n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633,
         n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641,
         n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649,
         n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657,
         n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665,
         n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673,
         n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681,
         n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689,
         n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697,
         n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705,
         n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713,
         n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721,
         n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729,
         n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737,
         n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745,
         n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753,
         n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761,
         n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769,
         n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777,
         n21778, n21779, n21780, n21781, n21782, n21783, n21784, n21785,
         n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793,
         n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801,
         n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809,
         n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817,
         n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825,
         n21826, n21827, n21828, n21829, n21830, n21831, n21832, n21833,
         n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841,
         n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849,
         n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857,
         n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865,
         n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873,
         n21874, n21875, n21876, n21877, n21878, n21879, n21880, n21881,
         n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889,
         n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897,
         n21898, n21899, n21900, n21901, n21902, n21903, n21904, n21905,
         n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913,
         n21914, n21915, n21916, n21917, n21918, n21919, n21920, n21921,
         n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929,
         n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937,
         n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945,
         n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953,
         n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961,
         n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969,
         n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977,
         n21978, n21979, n21980, n21981, n21982, n21983, n21984, n21985,
         n21986, n21987, n21988, n21989, n21990, n21991, n21992, n21993,
         n21994, n21995, n21996, n21997, n21998, n21999, n22000, n22001,
         n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009,
         n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017,
         n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025,
         n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033,
         n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041,
         n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049,
         n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057,
         n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065,
         n22066, n22067, n22068, n22069, n22070, n22071, n22072, n22073,
         n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081,
         n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089,
         n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097,
         n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105,
         n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113,
         n22114, n22115, n22116, n22117, n22118, n22119, n22120, n22121,
         n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129,
         n22130, n22131, n22132, n22133, n22134, n22135, n22136, n22137,
         n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145,
         n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153,
         n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161,
         n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169,
         n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177,
         n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185,
         n22186, n22187, n22188, n22189, n22190, n22191, n22192, n22193,
         n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201,
         n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209,
         n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217,
         n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225,
         n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233,
         n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241,
         n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249,
         n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257,
         n22258, n22259, n22260, n22261, n22262, n22263, n22264, n22265,
         n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273,
         n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281,
         n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289,
         n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297,
         n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305,
         n22306, n22307, n22308, n22309, n22310, n22311, n22312, n22313,
         n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321,
         n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329,
         n22330, n22331, n22332, n22333, n22334, n22335, n22336, n22337,
         n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345,
         n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353,
         n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361,
         n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369,
         n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377,
         n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385,
         n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393,
         n22394, n22395, n22396, n22397, n22398, n22399, n22400, n22401,
         n22402, n22403, n22404, n22405, n22406, n22407, n22408, n22409,
         n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417,
         n22418, n22419, n22420, n22421, n22422, n22423, n22424, n22425,
         n22426, n22427, n22428, n22429, n22430, n22431, n22432, n22433,
         n22434, n22435, n22436, n22437, n22438, n22439, n22440, n22441,
         n22442, n22443, n22444, n22445, n22446, n22447, n22448, n22449,
         n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457,
         n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465,
         n22466, n22467, n22468, n22469, n22470, n22471, n22472, n22473,
         n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22481,
         n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489,
         n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497,
         n22498, n22499, n22500, n22501, n22502, n22503, n22504, n22505,
         n22506, n22507, n22508, n22509, n22510, n22511, n22512, n22513,
         n22514, n22515, n22516, n22517, n22518, n22519, n22520, n22521,
         n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529,
         n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537,
         n22538, n22539, n22540, n22541, n22542, n22543, n22544, n22545,
         n22546, n22547, n22548, n22549, n22550, n22551, n22552, n22553,
         n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561,
         n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569,
         n22570, n22571, n22572, n22573, n22574, n22575, n22576, n22577,
         n22578, n22579, n22580, n22581, n22582, n22583, n22584, n22585,
         n22586, n22587, n22588, n22589, n22590, n22591, n22592, n22593,
         n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22601,
         n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609,
         n22610, n22611, n22612, n22613, n22614, n22615, n22616, n22617,
         n22618, n22619, n22620, n22621, n22622, n22623, n22624, n22625,
         n22626, n22627, n22628, n22629, n22630, n22631, n22632, n22633,
         n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641,
         n22642, n22643, n22644, n22645, n22646, n22647, n22648, n22649,
         n22650, n22651, n22652, n22653, n22654, n22655, n22656, n22657,
         n22658, n22659, n22660, n22661, n22662, n22663, n22664, n22665,
         n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673,
         n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681,
         n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689,
         n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697,
         n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705,
         n22706, n22707, n22708, n22709, n22710, n22711, n22712, n22713,
         n22714, n22715, n22716, n22717, n22718, n22719, n22720, n22721,
         n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729,
         n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737,
         n22738, n22739, n22740, n22741, n22742, n22743, n22744, n22745,
         n22746, n22747, n22748, n22749, n22750, n22751, n22752, n22753,
         n22754, n22755, n22756, n22757, n22758, n22759, n22760, n22761,
         n22762, n22763, n22764, n22765, n22766, n22767, n22768, n22769,
         n22770, n22771, n22772, n22773, n22774, n22775, n22776, n22777,
         n22778, n22779, n22780, n22781, n22782, n22783, n22784, n22785,
         n22786, n22787, n22788, n22789, n22790, n22791, n22792, n22793,
         n22794, n22795, n22796, n22797, n22798, n22799, n22800, n22801,
         n22802, n22803, n22804, n22805, n22806, n22807, n22808, n22809,
         n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22817,
         n22818, n22819, n22820, n22821, n22822, n22823, n22824, n22825,
         n22826, n22827, n22828, n22829, n22830, n22831, n22832, n22833,
         n22834, n22835, n22836, n22837, n22838, n22839, n22840, n22841,
         n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849,
         n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857,
         n22858, n22859, n22860, n22861, n22862, n22863, n22864, n22865,
         n22866, n22867, n22868, n22869, n22870, n22871, n22872, n22873,
         n22874, n22875, n22876, n22877, n22878, n22879, n22880, n22881,
         n22882, n22883, n22884, n22885, n22886, n22887, n22888, n22889,
         n22890, n22891, n22892, n22893, n22894, n22895, n22896, n22897,
         n22898, n22899, n22900, n22901, n22902, n22903, n22904, n22905,
         n22906, n22907, n22908, n22909, n22910, n22911, n22912, n22913,
         n22914, n22915, n22916, n22917, n22918, n22919, n22920, n22921,
         n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929,
         n22930, n22931, n22932, n22933, n22934, n22935, n22936, n22937,
         n22938, n22939, n22940, n22941, n22942, n22943, n22944, n22945,
         n22946, n22947, n22948, n22949, n22950, n22951, n22952, n22953,
         n22954, n22955, n22956, n22957, n22958, n22959, n22960, n22961,
         n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969,
         n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977,
         n22978, n22979, n22980, n22981, n22982, n22983, n22984, n22985,
         n22986, n22987, n22988, n22989, n22990, n22991, n22992, n22993,
         n22994, n22995, n22996, n22997, n22998, n22999, n23000, n23001,
         n23002, n23003, n23004, n23005, n23006, n23007, n23008, n23009,
         n23010, n23011, n23012, n23013, n23014, n23015, n23016, n23017,
         n23018, n23019, n23020, n23021, n23022, n23023, n23024, n23025,
         n23026, n23027, n23028, n23029, n23030, n23031, n23032, n23033,
         n23034, n23035, n23036, n23037, n23038, n23039, n23040, n23041,
         n23042, n23043, n23044, n23045, n23046, n23047, n23048, n23049,
         n23050, n23051, n23052, n23053, n23054, n23055, n23056, n23057,
         n23058, n23059, n23060, n23061, n23062, n23063, n23064, n23065,
         n23066, n23067, n23068, n23069, n23070, n23071, n23072, n23073,
         n23074, n23075, n23076, n23077, n23078, n23079, n23080, n23081,
         n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089,
         n23090, n23091, n23092, n23093, n23094, n23095, n23096, n23097,
         n23098, n23099, n23100, n23101, n23102, n23103, n23104, n23105,
         n23106, n23107, n23108, n23109, n23110, n23111, n23112, n23113,
         n23114, n23115, n23116, n23117, n23118, n23119, n23120, n23121,
         n23122, n23123, n23124, n23125, n23126, n23127, n23128, n23129,
         n23130, n23131, n23132, n23133, n23134, n23135, n23136, n23137,
         n23138, n23139, n23140, n23141, n23142, n23143, n23144, n23145,
         n23146, n23147, n23148, n23149, n23150, n23151, n23152, n23153,
         n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161,
         n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169,
         n23170, n23171, n23172, n23173, n23174, n23175, n23176, n23177,
         n23178, n23179, n23180, n23181, n23182, n23183, n23184, n23185,
         n23186, n23187, n23188, n23189, n23190, n23191, n23192, n23193,
         n23194, n23195, n23196, n23197, n23198, n23199, n23200, n23201,
         n23202, n23203, n23204, n23205, n23206, n23207, n23208, n23209,
         n23210, n23211, n23212, n23213, n23214, n23215, n23216, n23217,
         n23218, n23219, n23220, n23221, n23222, n23223, n23224, n23225,
         n23226, n23227, n23228, n23229, n23230, n23231, n23232, n23233,
         n23234, n23235, n23236, n23237, n23238, n23239, n23240, n23241,
         n23242, n23243, n23244, n23245, n23246, n23247, n23248, n23249,
         n23250, n23251, n23252, n23253, n23254, n23255, n23256, n23257,
         n23258, n23259, n23260, n23261, n23262, n23263, n23264, n23265,
         n23266, n23267, n23268, n23269, n23270, n23271, n23272, n23273,
         n23274, n23275, n23276, n23277, n23278, n23279, n23280, n23281,
         n23282, n23283, n23284, n23285, n23286, n23287, n23288, n23289,
         n23290, n23291, n23292, n23293, n23294, n23295, n23296, n23297,
         n23298, n23299, n23300, n23301, n23302, n23303, n23304, n23305,
         n23306, n23307, n23308, n23309, n23310, n23311, n23312, n23313,
         n23314, n23315, n23316, n23317, n23318, n23319, n23320, n23321,
         n23322, n23323, n23324, n23325, n23326, n23327, n23328, n23329,
         n23330, n23331, n23332, n23333, n23334, n23335, n23336, n23337,
         n23338, n23339, n23340, n23341, n23342, n23343, n23344, n23345,
         n23346, n23347, n23348, n23349, n23350, n23351, n23352, n23353,
         n23354, n23355, n23356, n23357, n23358, n23359, n23360, n23361,
         n23362, n23363, n23364, n23365, n23366, n23367, n23368, n23369,
         n23370, n23371, n23372, n23373, n23374, n23375, n23376, n23377,
         n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385,
         n23386, n23387, n23388, n23389, n23390, n23391, n23392, n23393,
         n23394, n23395, n23396, n23397, n23398, n23399, n23400, n23401,
         n23402, n23403, n23404, n23405, n23406, n23407, n23408, n23409,
         n23410, n23411, n23412, n23413, n23414, n23415, n23416, n23417,
         n23418, n23419, n23420, n23421, n23422, n23423, n23424, n23425,
         n23426, n23427, n23428, n23429, n23430, n23431, n23432, n23433,
         n23434, n23435, n23436, n23437, n23438, n23439, n23440, n23441,
         n23442, n23443, n23444, n23445, n23446, n23447, n23448, n23449,
         n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457,
         n23458, n23459, n23460, n23461, n23462, n23463, n23464, n23465,
         n23466, n23467, n23468, n23469, n23470, n23471, n23472, n23473,
         n23474, n23475, n23476, n23477, n23478, n23479, n23480, n23481,
         n23482, n23483, n23484, n23485, n23486, n23487, n23488, n23489,
         n23490, n23491, n23492, n23493, n23494, n23495, n23496, n23497,
         n23498, n23499, n23500, n23501, n23502, n23503, n23504, n23505,
         n23506, n23507, n23508, n23509, n23510, n23511, n23512, n23513,
         n23514, n23515, n23516, n23517, n23518, n23519, n23520, n23521,
         n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23529,
         n23530, n23531, n23532, n23533, n23534, n23535, n23536, n23537,
         n23538, n23539, n23540, n23541, n23542, n23543, n23544, n23545,
         n23546, n23547, n23548, n23549, n23550, n23551, n23552, n23553,
         n23554, n23555, n23556, n23557, n23558, n23559, n23560, n23561,
         n23562, n23563, n23564, n23565, n23566, n23567, n23568, n23569,
         n23570, n23571, n23572, n23573, n23574, n23575, n23576, n23577,
         n23578, n23579, n23580, n23581, n23582, n23583, n23584, n23585,
         n23586, n23587, n23588, n23589, n23590, n23591, n23592, n23593,
         n23594, n23595, n23596, n23597, n23598, n23599, n23600, n23601,
         n23602, n23603, n23604, n23605, n23606, n23607, n23608, n23609,
         n23610, n23611, n23612, n23613, n23614, n23615, n23616, n23617,
         n23618, n23619, n23620, n23621, n23622, n23623, n23624, n23625,
         n23626, n23627, n23628, n23629, n23630, n23631, n23632, n23633,
         n23634, n23635, n23636, n23637, n23638, n23639, n23640, n23641,
         n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649,
         n23650, n23651, n23652, n23653, n23654, n23655, n23656, n23657,
         n23658, n23659, n23660, n23661, n23662, n23663, n23664, n23665,
         n23666, n23667, n23668, n23669, n23670, n23671, n23672, n23673,
         n23674, n23675, n23676, n23677, n23678, n23679, n23680, n23681,
         n23682, n23683, n23684, n23685, n23686, n23687, n23688, n23689,
         n23690, n23691, n23692, n23693, n23694, n23695, n23696, n23697,
         n23698, n23699, n23700, n23701, n23702, n23703, n23704, n23705,
         n23706, n23707, n23708, n23709, n23710, n23711, n23712, n23713,
         n23714, n23715, n23716, n23717, n23718, n23719, n23720, n23721,
         n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729,
         n23730, n23731, n23732, n23733, n23734, n23735, n23736, n23737,
         n23738, n23739, n23740, n23741, n23742, n23743, n23744, n23745,
         n23746, n23747, n23748, n23749, n23750, n23751, n23752, n23753,
         n23754, n23755, n23756, n23757, n23758, n23759, n23760, n23761,
         n23762, n23763, n23764, n23765, n23766, n23767, n23768, n23769,
         n23770, n23771, n23772, n23773, n23774, n23775, n23776, n23777,
         n23778, n23779, n23780, n23781, n23782, n23783, n23784, n23785,
         n23786, n23787, n23788, n23789, n23790, n23791, n23792, n23793,
         n23794, n23795, n23796, n23797, n23798, n23799, n23800, n23801,
         n23802, n23803, n23804, n23805, n23806, n23807, n23808, n23809,
         n23810, n23811, n23812, n23813, n23814, n23815, n23816, n23817,
         n23818, n23819, n23820, n23821, n23822, n23823, n23824, n23825,
         n23826, n23827, n23828, n23829, n23830, n23831, n23832, n23833,
         n23834, n23835, n23836, n23837, n23838, n23839, n23840, n23841,
         n23842, n23843, n23844, n23845, n23846, n23847, n23848, n23849,
         n23850, n23851, n23852, n23853, n23854, n23855, n23856, n23857,
         n23858, n23859, n23860, n23861, n23862, n23863, n23864, n23865,
         n23866, n23867, n23868, n23869, n23870, n23871, n23872, n23873,
         n23874, n23875, n23876, n23877, n23878, n23879, n23880, n23881,
         n23882, n23883, n23884, n23885, n23886, n23887, n23888, n23889,
         n23890, n23891, n23892, n23893, n23894, n23895, n23896, n23897,
         n23898, n23899, n23900, n23901, n23902, n23903, n23904, n23905,
         n23906, n23907, n23908, n23909, n23910, n23911, n23912, n23913,
         n23914, n23915, n23916, n23917, n23918, n23919, n23920, n23921,
         n23922, n23923, n23924, n23925, n23926, n23927, n23928, n23929,
         n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937,
         n23938, n23939, n23940, n23941, n23942, n23943, n23944, n23945,
         n23946, n23947, n23948, n23949, n23950, n23951, n23952, n23953,
         n23954, n23955, n23956, n23957, n23958, n23959, n23960, n23961,
         n23962, n23963, n23964, n23965, n23966, n23967, n23968, n23969,
         n23970, n23971, n23972, n23973, n23974, n23975, n23976, n23977,
         n23978, n23979, n23980, n23981, n23982, n23983, n23984, n23985,
         n23986, n23987, n23988, n23989, n23990, n23991, n23992, n23993,
         n23994, n23995, n23996, n23997, n23998, n23999, n24000, n24001,
         n24002, n24003, n24004, n24005, n24006, n24007, n24008, n24009,
         n24010, n24011, n24012, n24013, n24014, n24015, n24016, n24017,
         n24018, n24019, n24020, n24021, n24022, n24023, n24024, n24025,
         n24026, n24027, n24028, n24029, n24030, n24031, n24032, n24033,
         n24034, n24035, n24036, n24037, n24038, n24039, n24040, n24041,
         n24042, n24043, n24044, n24045, n24046, n24047, n24048, n24049,
         n24050, n24051, n24052, n24053, n24054, n24055, n24056, n24057,
         n24058, n24059, n24060, n24061, n24062, n24063, n24064, n24065,
         n24066, n24067, n24068, n24069, n24070, n24071, n24072, n24073,
         n24074, n24075, n24076, n24077, n24078, n24079, n24080, n24081,
         n24082, n24083, n24084, n24085, n24086, n24087, n24088, n24089,
         n24090, n24091, n24092, n24093, n24094, n24095, n24096, n24097,
         n24098, n24099, n24100, n24101, n24102, n24103, n24104, n24105,
         n24106, n24107, n24108, n24109, n24110, n24111, n24112, n24113,
         n24114, n24115, n24116, n24117, n24118, n24119, n24120, n24121,
         n24122, n24123, n24124, n24125, n24126, n24127, n24128, n24129,
         n24130, n24131, n24132, n24133, n24134, n24135, n24136, n24137,
         n24138, n24139, n24140, n24141, n24142, n24143, n24144, n24145,
         n24146, n24147, n24148, n24149, n24150, n24151, n24152, n24153,
         n24154, n24155, n24156, n24157, n24158, n24159, n24160, n24161,
         n24162, n24163, n24164, n24165, n24166, n24167, n24168, n24169,
         n24170, n24171, n24172, n24173, n24174, n24175, n24176, n24177,
         n24178, n24179, n24180, n24181, n24182, n24183, n24184, n24185,
         n24186, n24187, n24188, n24189, n24190, n24191, n24192, n24193,
         n24194, n24195, n24196, n24197, n24198, n24199, n24200, n24201,
         n24202, n24203, n24204, n24205, n24206, n24207, n24208, n24209,
         n24210, n24211, n24212, n24213, n24214, n24215, n24216, n24217,
         n24218, n24219, n24220, n24221, n24222, n24223, n24224, n24225,
         n24226, n24227, n24228, n24229, n24230, n24231, n24232, n24233,
         n24234, n24235, n24236, n24237, n24238, n24239, n24240, n24241,
         n24242, n24243, n24244, n24245, n24246, n24247, n24248, n24249,
         n24250, n24251, n24252, n24253, n24254, n24255, n24256, n24257,
         n24258, n24259, n24260, n24261, n24262, n24263, n24264, n24265,
         n24266, n24267, n24268, n24269, n24270, n24271, n24272, n24273,
         n24274, n24275, n24276, n24277, n24278, n24279, n24280, n24281,
         n24282, n24283, n24284, n24285, n24286, n24287, n24288, n24289,
         n24290, n24291, n24292, n24293, n24294, n24295, n24296, n24297,
         n24298, n24299, n24300, n24301, n24302, n24303, n24304, n24305,
         n24306, n24307, n24308, n24309, n24310, n24311, n24312, n24313,
         n24314, n24315, n24316, n24317, n24318, n24319, n24320, n24321,
         n24322, n24323, n24324, n24325, n24326, n24327, n24328, n24329,
         n24330, n24331, n24332, n24333, n24334, n24335, n24336, n24337,
         n24338, n24339, n24340, n24341, n24342, n24343, n24344, n24345,
         n24346, n24347, n24348, n24349, n24350, n24351, n24352, n24353,
         n24354, n24355, n24356, n24357, n24358, n24359, n24360, n24361,
         n24362, n24363, n24364, n24365, n24366, n24367, n24368, n24369,
         n24370, n24371, n24372, n24373, n24374, n24375, n24376, n24377,
         n24378, n24379, n24380, n24381, n24382, n24383, n24384, n24385,
         n24386, n24387, n24388, n24389, n24390, n24391, n24392, n24393,
         n24394, n24395, n24396, n24397, n24398, n24399, n24400, n24401,
         n24402, n24403, n24404, n24405, n24406, n24407, n24408, n24409,
         n24410, n24411, n24412, n24413, n24414, n24415, n24416, n24417,
         n24418, n24419, n24420, n24421, n24422, n24423, n24424, n24425,
         n24426, n24427, n24428, n24429, n24430, n24431, n24432, n24433,
         n24434, n24435, n24436, n24437, n24438, n24439, n24440, n24441,
         n24442, n24443, n24444, n24445, n24446, n24447, n24448, n24449,
         n24450, n24451, n24452, n24453, n24454, n24455, n24456, n24457,
         n24458, n24459, n24460, n24461, n24462, n24463, n24464, n24465,
         n24466, n24467, n24468, n24469, n24470, n24471, n24472, n24473,
         n24474, n24475, n24476, n24477, n24478, n24479, n24480, n24481,
         n24482, n24483, n24484, n24485, n24486, n24487, n24488, n24489,
         n24490, n24491, n24492, n24493, n24494, n24495, n24496, n24497,
         n24498, n24499, n24500, n24501, n24502, n24503, n24504, n24505,
         n24506, n24507, n24508, n24509, n24510, n24511, n24512, n24513,
         n24514, n24515, n24516, n24517, n24518, n24519, n24520, n24521,
         n24522, n24523, n24524, n24525, n24526, n24527, n24528, n24529,
         n24530, n24531, n24532, n24533, n24534, n24535, n24536, n24537,
         n24538, n24539, n24540, n24541, n24542, n24543, n24544, n24545,
         n24546, n24547, n24548, n24549, n24550, n24551, n24552, n24553,
         n24554, n24555, n24556, n24557, n24558, n24559, n24560, n24561,
         n24562, n24563, n24564, n24565, n24566, n24567, n24568, n24569,
         n24570, n24571, n24572, n24573, n24574, n24575, n24576, n24577,
         n24578, n24579, n24580, n24581, n24582, n24583, n24584, n24585,
         n24586, n24587, n24588, n24589, n24590, n24591, n24592, n24593,
         n24594, n24595, n24596, n24597, n24598, n24599, n24600, n24601,
         n24602, n24603, n24604, n24605, n24606, n24607, n24608, n24609,
         n24610, n24611, n24612, n24613, n24614, n24615, n24616, n24617,
         n24618, n24619, n24620, n24621, n24622, n24623, n24624, n24625,
         n24626, n24627, n24628, n24629, n24630, n24631, n24632, n24633,
         n24634, n24635, n24636, n24637, n24638, n24639, n24640, n24641,
         n24642, n24643, n24644, n24645, n24646, n24647, n24648, n24649,
         n24650, n24651, n24652, n24653, n24654, n24655, n24656, n24657,
         n24658, n24659, n24660, n24661, n24662, n24663, n24664, n24665,
         n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673,
         n24674, n24675, n24676, n24677, n24678, n24679, n24680, n24681,
         n24682, n24683, n24684, n24685, n24686, n24687, n24688, n24689,
         n24690, n24691, n24692, n24693, n24694, n24695, n24696, n24697,
         n24698, n24699, n24700, n24701, n24702, n24703, n24704, n24705,
         n24706, n24707, n24708, n24709, n24710, n24711, n24712, n24713,
         n24714, n24715, n24716, n24717, n24718, n24719, n24720, n24721,
         n24722, n24723, n24724, n24725, n24726, n24727, n24728, n24729,
         n24730, n24731, n24732, n24733, n24734, n24735, n24736, n24737,
         n24738, n24739, n24740, n24741, n24742, n24743, n24744, n24745,
         n24746, n24747, n24748, n24749, n24750, n24751, n24752, n24753,
         n24754, n24755, n24756, n24757, n24758, n24759, n24760, n24761,
         n24762, n24763, n24764, n24765, n24766, n24767, n24768, n24769,
         n24770, n24771, n24772, n24773, n24774, n24775, n24776, n24777,
         n24778, n24779, n24780, n24781, n24782, n24783, n24784, n24785,
         n24786, n24787, n24788, n24789, n24790, n24791, n24792, n24793,
         n24794, n24795, n24796, n24797, n24798, n24799, n24800, n24801,
         n24802, n24803, n24804, n24805, n24806, n24807, n24808, n24809,
         n24810, n24811, n24812, n24813, n24814, n24815, n24816, n24817,
         n24818, n24819, n24820, n24821, n24822, n24823, n24824, n24825,
         n24826, n24827, n24828, n24829, n24830, n24831, n24832, n24833,
         n24834, n24835, n24836, n24837, n24838, n24839, n24840, n24841,
         n24842, n24843, n24844, n24845, n24846, n24847, n24848, n24849,
         n24850, n24851, n24852, n24853, n24854, n24855, n24856, n24857,
         n24858, n24859, n24860, n24861, n24862, n24863, n24864, n24865,
         n24866, n24867, n24868, n24869, n24870, n24871, n24872, n24873,
         n24874, n24875, n24876, n24877, n24878, n24879, n24880, n24881,
         n24882, n24883, n24884, n24885, n24886, n24887, n24888, n24889,
         n24890, n24891, n24892, n24893, n24894, n24895, n24896, n24897,
         n24898, n24899, n24900, n24901, n24902, n24903, n24904, n24905,
         n24906, n24907, n24908, n24909, n24910, n24911, n24912, n24913,
         n24914, n24915, n24916, n24917, n24918, n24919, n24920, n24921,
         n24922, n24923, n24924, n24925, n24926, n24927, n24928, n24929,
         n24930, n24931, n24932, n24933, n24934, n24935, n24936, n24937,
         n24938, n24939, n24940, n24941, n24942, n24943, n24944, n24945,
         n24946, n24947, n24948, n24949, n24950, n24951, n24952, n24953,
         n24954, n24955, n24956, n24957, n24958, n24959, n24960, n24961,
         n24962, n24963, n24964, n24965, n24966, n24967, n24968, n24969,
         n24970, n24971, n24972, n24973, n24974, n24975, n24976, n24977,
         n24978, n24979, n24980, n24981, n24982, n24983, n24984, n24985,
         n24986, n24987, n24988, n24989, n24990, n24991, n24992, n24993,
         n24994, n24995, n24996, n24997, n24998, n24999, n25000, n25001,
         n25002, n25003, n25004, n25005, n25006, n25007, n25008, n25009,
         n25010, n25011, n25012, n25013, n25014, n25015, n25016, n25017,
         n25018, n25019, n25020, n25021, n25022, n25023, n25024, n25025,
         n25026, n25027, n25028, n25029, n25030, n25031, n25032, n25033,
         n25034, n25035, n25036, n25037, n25038, n25039, n25040, n25041,
         n25042, n25043, n25044, n25045, n25046, n25047, n25048, n25049,
         n25050, n25051, n25052, n25053, n25054, n25055, n25056, n25057,
         n25058, n25059, n25060, n25061, n25062, n25063, n25064, n25065,
         n25066, n25067, n25068, n25069, n25070, n25071, n25072, n25073,
         n25074, n25075, n25076, n25077, n25078, n25079, n25080, n25081,
         n25082, n25083, n25084, n25085, n25086, n25087, n25088, n25089,
         n25090, n25091, n25092, n25093, n25094, n25095, n25096, n25097,
         n25098, n25099, n25100, n25101, n25102, n25103, n25104, n25105,
         n25106, n25107, n25108, n25109, n25110, n25111, n25112, n25113,
         n25114, n25115, n25116, n25117, n25118, n25119, n25120, n25121,
         n25122, n25123, n25124, n25125, n25126, n25127, n25128, n25129,
         n25130, n25131, n25132, n25133, n25134, n25135, n25136, n25137,
         n25138, n25139, n25140, n25141, n25142, n25143, n25144, n25145,
         n25146, n25147, n25148, n25149, n25150, n25151, n25152, n25153,
         n25154, n25155, n25156, n25157, n25158, n25159, n25160, n25161,
         n25162, n25163, n25164, n25165, n25166, n25167, n25168, n25169,
         n25170, n25171, n25172, n25173, n25174, n25175, n25176, n25177,
         n25178, n25179, n25180, n25181, n25182, n25183, n25184, n25185,
         n25186, n25187, n25188, n25189, n25190, n25191, n25192, n25193,
         n25194, n25195, n25196, n25197, n25198, n25199, n25200, n25201,
         n25202, n25203, n25204, n25205, n25206, n25207, n25208, n25209,
         n25210, n25211, n25212, n25213, n25214, n25215, n25216, n25217,
         n25218, n25219, n25220, n25221, n25222, n25223, n25224, n25225,
         n25226, n25227, n25228, n25229, n25230, n25231, n25232, n25233,
         n25234, n25235, n25236, n25237, n25238, n25239, n25240, n25241,
         n25242, n25243, n25244, n25245, n25246, n25247, n25248, n25249,
         n25250, n25251, n25252, n25253, n25254, n25255, n25256, n25257,
         n25258, n25259, n25260, n25261, n25262, n25263, n25264, n25265,
         n25266, n25267, n25268, n25269, n25270, n25271, n25272, n25273,
         n25274, n25275, n25276, n25277, n25278, n25279, n25280, n25281,
         n25282, n25283, n25284, n25285, n25286, n25287, n25288, n25289,
         n25290, n25291, n25292, n25293, n25294, n25295, n25296, n25297,
         n25298, n25299, n25300, n25301, n25302, n25303, n25304, n25305,
         n25306, n25307, n25308, n25309, n25310, n25311, n25312, n25313,
         n25314, n25315, n25316, n25317, n25318, n25319, n25320, n25321,
         n25322, n25323, n25324, n25325, n25326, n25327, n25328, n25329,
         n25330, n25331, n25332, n25333, n25334, n25335, n25336, n25337,
         n25338, n25339, n25340, n25341, n25342, n25343, n25344, n25345,
         n25346, n25347, n25348, n25349, n25350, n25351, n25352, n25353,
         n25354, n25355, n25356, n25357, n25358, n25359, n25360, n25361,
         n25362, n25363, n25364, n25365, n25366, n25367, n25368, n25369,
         n25370, n25371, n25372, n25373, n25374, n25375, n25376, n25377,
         n25378, n25379, n25380, n25381, n25382, n25383, n25384, n25385,
         n25386, n25387, n25388, n25389, n25390, n25391, n25392, n25393,
         n25394, n25395, n25396, n25397, n25398, n25399, n25400, n25401,
         n25402, n25403, n25404, n25405, n25406, n25407, n25408, n25409,
         n25410, n25411, n25412, n25413, n25414, n25415, n25416, n25417,
         n25418, n25419, n25420, n25421, n25422, n25423, n25424, n25425,
         n25426, n25427, n25428, n25429, n25430, n25431, n25432, n25433,
         n25434, n25435, n25436, n25437, n25438, n25439, n25440, n25441,
         n25442, n25443, n25444, n25445, n25446, n25447, n25448, n25449,
         n25450, n25451, n25452, n25453, n25454, n25455, n25456, n25457,
         n25458, n25459, n25460, n25461, n25462, n25463, n25464, n25465,
         n25466, n25467, n25468, n25469, n25470, n25471, n25472, n25473,
         n25474, n25475, n25476, n25477, n25478, n25479, n25480, n25481,
         n25482, n25483, n25484, n25485, n25486, n25487, n25488, n25489,
         n25490, n25491, n25492, n25493, n25494, n25495, n25496, n25497,
         n25498, n25499, n25500, n25501, n25502, n25503, n25504, n25505,
         n25506, n25507, n25508, n25509, n25510, n25511, n25512, n25513,
         n25514, n25515, n25516, n25517, n25518, n25519, n25520, n25521,
         n25522, n25523, n25524, n25525, n25526, n25527, n25528, n25529,
         n25530, n25531, n25532, n25533, n25534, n25535, n25536, n25537,
         n25538, n25539, n25540, n25541, n25542, n25543, n25544, n25545,
         n25546, n25547, n25548, n25549, n25550, n25551, n25552, n25553,
         n25554, n25555, n25556, n25557, n25558, n25559, n25560, n25561,
         n25562, n25563, n25564, n25565, n25566, n25567, n25568, n25569,
         n25570, n25571, n25572, n25573, n25574, n25575, n25576, n25577,
         n25578, n25579, n25580, n25581, n25582, n25583, n25584, n25585,
         n25586, n25587, n25588, n25589, n25590, n25591, n25592, n25593,
         n25594, n25595, n25596, n25597, n25598, n25599, n25600, n25601,
         n25602, n25603, n25604, n25605, n25606, n25607, n25608, n25609,
         n25610, n25611, n25612, n25613, n25614, n25615, n25616, n25617,
         n25618, n25619, n25620, n25621, n25622, n25623, n25624, n25625,
         n25626, n25627, n25628, n25629, n25630, n25631, n25632, n25633,
         n25634, n25635, n25636, n25637, n25638, n25639, n25640, n25641,
         n25642, n25643, n25644, n25645, n25646, n25647, n25648, n25649,
         n25650, n25651, n25652, n25653, n25654, n25655, n25656, n25657,
         n25658, n25659, n25660, n25661, n25662, n25663, n25664, n25665,
         n25666, n25667, n25668, n25669, n25670, n25671, n25672, n25673,
         n25674, n25675, n25676, n25677, n25678, n25679, n25680, n25681,
         n25682, n25683, n25684, n25685, n25686, n25687, n25688, n25689,
         n25690, n25691, n25692, n25693, n25694, n25695, n25696, n25697,
         n25698, n25699, n25700, n25701, n25702, n25703, n25704, n25705,
         n25706, n25707, n25708, n25709, n25710, n25711, n25712, n25713,
         n25714, n25715, n25716, n25717, n25718, n25719, n25720, n25721,
         n25722, n25723, n25724, n25725, n25726, n25727, n25728, n25729,
         n25730, n25731, n25732, n25733, n25734, n25735, n25736, n25737,
         n25738, n25739, n25740, n25741, n25742, n25743, n25744, n25745,
         n25746, n25747, n25748, n25749, n25750, n25751, n25752, n25753,
         n25754, n25755, n25756, n25757, n25758, n25759, n25760, n25761,
         n25762, n25763, n25764, n25765, n25766, n25767, n25768, n25769,
         n25770, n25771, n25772, n25773, n25774, n25775, n25776, n25777,
         n25778, n25779, n25780, n25781, n25782, n25783, n25784, n25785,
         n25786, n25787, n25788, n25789, n25790, n25791, n25792, n25793,
         n25794, n25795, n25796, n25797, n25798, n25799, n25800, n25801,
         n25802, n25803, n25804, n25805, n25806, n25807, n25808, n25809,
         n25810, n25811, n25812, n25813, n25814, n25815, n25816, n25817,
         n25818, n25819, n25820, n25821, n25822, n25823, n25824, n25825,
         n25826, n25827, n25828, n25829, n25830, n25831, n25832, n25833,
         n25834, n25835, n25836, n25837, n25838, n25839, n25840, n25841,
         n25842, n25843, n25844, n25845, n25846, n25847, n25848, n25849,
         n25850, n25851, n25852, n25853, n25854, n25855, n25856, n25857,
         n25858, n25859, n25860, n25861, n25862, n25863, n25864, n25865,
         n25866, n25867, n25868, n25869, n25870, n25871, n25872, n25873,
         n25874, n25875, n25876, n25877, n25878, n25879, n25880, n25881,
         n25882, n25883, n25884, n25885, n25886, n25887, n25888, n25889,
         n25890, n25891, n25892, n25893, n25894, n25895, n25896, n25897,
         n25898, n25899, n25900, n25901, n25902, n25903, n25904, n25905,
         n25906, n25907, n25908, n25909, n25910, n25911, n25912, n25913,
         n25914, n25915, n25916, n25917, n25918, n25919, n25920, n25921,
         n25922, n25923, n25924, n25925, n25926, n25927, n25928, n25929,
         n25930, n25931, n25932, n25933, n25934, n25935, n25936, n25937,
         n25938, n25939, n25940, n25941, n25942, n25943, n25944, n25945,
         n25946, n25947, n25948, n25949, n25950, n25951, n25952, n25953,
         n25954, n25955, n25956, n25957, n25958, n25959, n25960, n25961,
         n25962, n25963, n25964, n25965, n25966, n25967, n25968, n25969,
         n25970, n25971, n25972, n25973, n25974, n25975, n25976, n25977,
         n25978, n25979, n25980, n25981, n25982, n25983, n25984, n25985,
         n25986, n25987, n25988, n25989, n25990, n25991, n25992, n25993,
         n25994, n25995, n25996, n25997, n25998, n25999, n26000, n26001,
         n26002, n26003, n26004, n26005, n26006, n26007, n26008, n26009,
         n26010, n26011, n26012, n26013, n26014, n26015, n26016, n26017,
         n26018, n26019, n26020, n26021, n26022, n26023, n26024, n26025,
         n26026, n26027, n26028, n26029, n26030, n26031, n26032, n26033,
         n26034, n26035, n26036, n26037, n26038, n26039, n26040, n26041,
         n26042, n26043, n26044, n26045, n26046, n26047, n26048, n26049,
         n26050, n26051, n26052, n26053, n26054, n26055, n26056, n26057,
         n26058, n26059, n26060, n26061, n26062, n26063, n26064, n26065,
         n26066, n26067, n26068, n26069, n26070, n26071, n26072, n26073,
         n26074, n26075, n26076, n26077, n26078, n26079, n26080, n26081,
         n26082, n26083, n26084, n26085, n26086, n26087, n26088, n26089,
         n26090, n26091, n26092, n26093, n26094, n26095, n26096, n26097,
         n26098, n26099, n26100, n26101, n26102, n26103, n26104, n26105,
         n26106, n26107, n26108, n26109, n26110, n26111, n26112, n26113,
         n26114, n26115, n26116, n26117, n26118, n26119, n26120, n26121,
         n26122, n26123, n26124, n26125, n26126, n26127, n26128, n26129,
         n26130, n26131, n26132, n26133, n26134, n26135, n26136, n26137,
         n26138, n26139, n26140, n26141, n26142, n26143, n26144, n26145,
         n26146, n26147, n26148, n26149, n26150, n26151, n26152, n26153,
         n26154, n26155, n26156, n26157, n26158, n26159, n26160, n26161,
         n26162, n26163, n26164, n26165, n26166, n26167, n26168, n26169,
         n26170, n26171, n26172, n26173, n26174, n26175, n26176, n26177,
         n26178, n26179, n26180, n26181, n26182, n26183, n26184, n26185,
         n26186, n26187, n26188, n26189, n26190, n26191, n26192, n26193,
         n26194, n26195, n26196, n26197, n26198, n26199, n26200, n26201,
         n26202, n26203, n26204, n26205, n26206, n26207, n26208, n26209,
         n26210, n26211, n26212, n26213, n26214, n26215, n26216, n26217,
         n26218, n26219, n26220, n26221, n26222, n26223, n26224, n26225,
         n26226, n26227, n26228, n26229, n26230, n26231, n26232, n26233,
         n26234, n26235, n26236, n26237, n26238, n26239, n26240, n26241,
         n26242, n26243, n26244, n26245, n26246, n26247, n26248, n26249,
         n26250, n26251, n26252, n26253, n26254, n26255, n26256, n26257,
         n26258, n26259, n26260, n26261, n26262, n26263, n26264, n26265,
         n26266, n26267, n26268, n26269, n26270, n26271, n26272, n26273,
         n26274, n26275, n26276, n26277, n26278, n26279, n26280, n26281,
         n26282, n26283, n26284, n26285, n26286, n26287, n26288, n26289,
         n26290, n26291, n26292, n26293, n26294, n26295, n26296, n26297,
         n26298, n26299, n26300, n26301, n26302, n26303, n26304, n26305,
         n26306, n26307, n26308, n26309, n26310, n26311, n26312, n26313,
         n26314, n26315, n26316, n26317, n26318, n26319, n26320, n26321,
         n26322, n26323, n26324, n26325, n26326, n26327, n26328, n26329,
         n26330, n26331, n26332, n26333, n26334, n26335, n26336, n26337,
         n26338, n26339, n26340, n26341, n26342, n26343, n26344, n26345,
         n26346, n26347, n26348, n26349, n26350, n26351, n26352, n26353,
         n26354, n26355, n26356, n26357, n26358, n26359, n26360, n26361,
         n26362, n26363, n26364, n26365, n26366, n26367, n26368, n26369,
         n26370, n26371, n26372, n26373, n26374, n26375, n26376, n26377,
         n26378, n26379, n26380, n26381, n26382, n26383, n26384, n26385,
         n26386, n26387, n26388, n26389, n26390, n26391, n26392, n26393,
         n26394, n26395, n26396, n26397, n26398, n26399, n26400, n26401,
         n26402, n26403, n26404, n26405, n26406, n26407, n26408, n26409,
         n26410, n26411, n26412, n26413, n26414, n26415, n26416, n26417,
         n26418, n26419, n26420, n26421, n26422, n26423, n26424, n26425,
         n26426, n26427, n26428, n26429, n26430, n26431, n26432, n26433,
         n26434, n26435, n26436, n26437, n26438, n26439, n26440, n26441,
         n26442, n26443, n26444, n26445, n26446, n26447, n26448, n26449,
         n26450, n26451, n26452, n26453, n26454, n26455, n26456, n26457,
         n26458, n26459, n26460, n26461, n26462, n26463, n26464, n26465,
         n26466, n26467, n26468, n26469, n26470, n26471, n26472, n26473,
         n26474, n26475, n26476, n26477, n26478, n26479, n26480, n26481,
         n26482, n26483, n26484, n26485, n26486, n26487, n26488, n26489,
         n26490, n26491, n26492, n26493, n26494, n26495, n26496, n26497,
         n26498, n26499, n26500, n26501, n26502, n26503, n26504, n26505,
         n26506, n26507, n26508, n26509, n26510, n26511, n26512, n26513,
         n26514, n26515, n26516, n26517, n26518, n26519, n26520, n26521,
         n26522, n26523, n26524, n26525, n26526, n26527, n26528, n26529,
         n26530, n26531, n26532, n26533, n26534, n26535, n26536, n26537,
         n26538, n26539, n26540, n26541, n26542, n26543, n26544, n26545,
         n26546, n26547, n26548, n26549, n26550, n26551, n26552, n26553,
         n26554, n26555, n26556, n26557, n26558, n26559, n26560, n26561,
         n26562, n26563, n26564, n26565, n26566, n26567, n26568, n26569,
         n26570, n26571, n26572, n26573, n26574, n26575, n26576, n26577,
         n26578, n26579, n26580, n26581, n26582, n26583, n26584, n26585,
         n26586, n26587, n26588, n26589, n26590, n26591, n26592, n26593,
         n26594, n26595, n26596, n26597, n26598, n26599, n26600, n26601,
         n26602, n26603, n26604, n26605, n26606, n26607, n26608, n26609,
         n26610, n26611, n26612, n26613, n26614, n26615, n26616, n26617,
         n26618, n26619, n26620, n26621, n26622, n26623, n26624, n26625,
         n26626, n26627, n26628, n26629, n26630, n26631, n26632, n26633,
         n26634, n26635, n26636, n26637, n26638, n26639, n26640, n26641,
         n26642, n26643, n26644, n26645, n26646, n26647, n26648, n26649,
         n26650, n26651, n26652, n26653, n26654, n26655, n26656, n26657,
         n26658, n26659, n26660, n26661, n26662, n26663, n26664, n26665,
         n26666, n26667, n26668, n26669, n26670, n26671, n26672, n26673,
         n26674, n26675, n26676, n26677, n26678, n26679, n26680, n26681,
         n26682, n26683, n26684, n26685, n26686, n26687, n26688, n26689,
         n26690, n26691, n26692, n26693, n26694, n26695, n26696, n26697,
         n26698, n26699, n26700, n26701, n26702, n26703, n26704, n26705,
         n26706, n26707, n26708, n26709, n26710, n26711, n26712, n26713,
         n26714, n26715, n26716, n26717, n26718, n26719, n26720, n26721,
         n26722, n26723, n26724, n26725, n26726, n26727, n26728, n26729,
         n26730, n26731, n26732, n26733, n26734, n26735, n26736, n26737,
         n26738, n26739, n26740, n26741, n26742, n26743, n26744, n26745,
         n26746, n26747, n26748, n26749, n26750, n26751, n26752, n26753,
         n26754, n26755, n26756, n26757, n26758, n26759, n26760, n26761,
         n26762, n26763, n26764, n26765, n26766, n26767, n26768, n26769,
         n26770, n26771, n26772, n26773, n26774, n26775, n26776, n26777,
         n26778, n26779, n26780, n26781, n26782, n26783, n26784, n26785,
         n26786, n26787, n26788, n26789, n26790, n26791, n26792, n26793,
         n26794, n26795, n26796, n26797, n26798, n26799, n26800, n26801,
         n26802, n26803, n26804, n26805, n26806, n26807, n26808, n26809,
         n26810, n26811, n26812, n26813, n26814, n26815, n26816, n26817,
         n26818, n26819, n26820, n26821, n26822, n26823, n26824, n26825,
         n26826, n26827, n26828, n26829, n26830, n26831, n26832, n26833,
         n26834, n26835, n26836, n26837, n26838, n26839, n26840, n26841,
         n26842, n26843, n26844, n26845, n26846, n26847, n26848, n26849,
         n26850, n26851, n26852, n26853, n26854, n26855, n26856, n26857,
         n26858, n26859, n26860, n26861, n26862, n26863, n26864, n26865,
         n26866, n26867, n26868, n26869, n26870, n26871, n26872, n26873,
         n26874, n26875, n26876, n26877, n26878, n26879, n26880, n26881,
         n26882, n26883, n26884, n26885, n26886, n26887, n26888, n26889,
         n26890, n26891, n26892, n26893, n26894, n26895, n26896, n26897,
         n26898, n26899, n26900, n26901, n26902, n26903, n26904, n26905,
         n26906, n26907, n26908, n26909, n26910, n26911, n26912, n26913,
         n26914, n26915, n26916, n26917, n26918, n26919, n26920, n26921,
         n26922, n26923, n26924, n26925, n26926, n26927, n26928, n26929,
         n26930, n26931, n26932, n26933, n26934, n26935, n26936, n26937,
         n26938, n26939, n26940, n26941, n26942, n26943, n26944, n26945,
         n26946, n26947, n26948, n26949, n26950, n26951, n26952, n26953,
         n26954, n26955, n26956, n26957, n26958, n26959, n26960, n26961,
         n26962, n26963, n26964, n26965, n26966, n26967, n26968, n26969,
         n26970, n26971, n26972, n26973, n26974, n26975, n26976, n26977,
         n26978, n26979, n26980, n26981, n26982, n26983, n26984, n26985,
         n26986, n26987, n26988, n26989, n26990, n26991, n26992, n26993,
         n26994, n26995, n26996, n26997, n26998, n26999, n27000, n27001,
         n27002, n27003, n27004, n27005, n27006, n27007, n27008, n27009,
         n27010, n27011, n27012, n27013, n27014, n27015, n27016, n27017,
         n27018, n27019, n27020, n27021, n27022, n27023, n27024, n27025,
         n27026, n27027, n27028, n27029, n27030, n27031, n27032, n27033,
         n27034, n27035, n27036, n27037, n27038, n27039, n27040, n27041,
         n27042, n27043, n27044, n27045, n27046, n27047, n27048, n27049,
         n27050, n27051, n27052, n27053, n27054, n27055, n27056, n27057,
         n27058, n27059, n27060, n27061, n27062, n27063, n27064, n27065,
         n27066, n27067, n27068, n27069, n27070, n27071, n27072, n27073,
         n27074, n27075, n27076, n27077, n27078, n27079, n27080, n27081,
         n27082, n27083, n27084, n27085, n27086, n27087, n27088, n27089,
         n27090, n27091, n27092, n27093, n27094, n27095, n27096, n27097,
         n27098, n27099, n27100, n27101, n27102, n27103, n27104, n27105,
         n27106, n27107, n27108, n27109, n27110, n27111, n27112, n27113,
         n27114, n27115, n27116, n27117, n27118, n27119, n27120, n27121,
         n27122, n27123, n27124, n27125, n27126, n27127, n27128, n27129,
         n27130, n27131, n27132, n27133, n27134, n27135, n27136, n27137,
         n27138, n27139, n27140, n27141, n27142, n27143, n27144, n27145,
         n27146, n27147, n27148, n27149, n27150, n27151, n27152, n27153,
         n27154, n27155, n27156, n27157, n27158, n27159, n27160, n27161,
         n27162, n27163, n27164, n27165, n27166, n27167, n27168, n27169,
         n27170, n27171, n27172, n27173, n27174, n27175, n27176, n27177,
         n27178, n27179, n27180, n27181, n27182, n27183, n27184, n27185,
         n27186, n27187, n27188, n27189, n27190, n27191, n27192, n27193,
         n27194, n27195, n27196, n27197, n27198, n27199, n27200, n27201,
         n27202, n27203, n27204, n27205, n27206, n27207, n27208, n27209,
         n27210, n27211, n27212, n27213, n27214, n27215, n27216, n27217,
         n27218, n27219, n27220, n27221, n27222, n27223, n27224, n27225,
         n27226, n27227, n27228, n27229, n27230, n27231, n27232, n27233,
         n27234, n27235, n27236, n27237, n27238, n27239, n27240, n27241,
         n27242, n27243, n27244, n27245, n27246, n27247, n27248, n27249,
         n27250, n27251, n27252, n27253, n27254, n27255, n27256, n27257,
         n27258, n27259, n27260, n27261, n27262, n27263, n27264, n27265,
         n27266, n27267, n27268, n27269, n27270, n27271, n27272, n27273,
         n27274, n27275, n27276, n27277, n27278, n27279, n27280, n27281,
         n27282, n27283, n27284, n27285, n27286, n27287, n27288, n27289,
         n27290, n27291, n27292, n27293, n27294, n27295, n27296, n27297,
         n27298, n27299, n27300, n27301, n27302, n27303, n27304, n27305,
         n27306, n27307, n27308, n27309, n27310, n27311, n27312, n27313,
         n27314, n27315, n27316, n27317, n27318, n27319, n27320, n27321,
         n27322, n27323, n27324, n27325, n27326, n27327, n27328, n27329,
         n27330, n27331, n27332, n27333, n27334, n27335, n27336, n27337,
         n27338, n27339, n27340, n27341, n27342, n27343, n27344, n27345,
         n27346, n27347, n27348, n27349, n27350, n27351, n27352, n27353,
         n27354, n27355, n27356, n27357, n27358, n27359, n27360, n27361,
         n27362, n27363, n27364, n27365, n27366, n27367, n27368, n27369,
         n27370, n27371, n27372, n27373, n27374, n27375, n27376, n27377,
         n27378, n27379, n27380, n27381, n27382, n27383, n27384, n27385,
         n27386, n27387, n27388, n27389, n27390, n27391, n27392, n27393,
         n27394, n27395, n27396, n27397, n27398, n27399, n27400, n27401,
         n27402, n27403, n27404, n27405, n27406, n27407, n27408, n27409,
         n27410, n27411, n27412, n27413, n27414, n27415, n27416, n27417,
         n27418, n27419, n27420, n27421, n27422, n27423, n27424, n27425,
         n27426, n27427, n27428, n27429, n27430, n27431, n27432, n27433,
         n27434, n27435, n27436, n27437, n27438, n27439, n27440, n27441,
         n27442, n27443, n27444, n27445, n27446, n27447, n27448, n27449,
         n27450, n27451, n27452, n27453, n27454, n27455, n27456, n27457,
         n27458, n27459, n27460, n27461, n27462, n27463, n27464, n27465,
         n27466, n27467, n27468, n27469, n27470, n27471, n27472, n27473,
         n27474, n27475, n27476, n27477, n27478, n27479, n27480, n27481,
         n27482, n27483, n27484, n27485, n27486, n27487, n27488, n27489,
         n27490, n27491, n27492, n27493, n27494, n27495, n27496, n27497,
         n27498, n27499, n27500, n27501, n27502, n27503, n27504, n27505,
         n27506, n27507, n27508, n27509, n27510, n27511, n27512, n27513,
         n27514, n27515, n27516, n27517, n27518, n27519, n27520, n27521,
         n27522, n27523, n27524, n27525, n27526, n27527, n27528, n27529,
         n27530, n27531, n27532, n27533, n27534, n27535, n27536, n27537,
         n27538, n27539, n27540, n27541, n27542, n27543, n27544, n27545,
         n27546, n27547, n27548, n27549, n27550, n27551, n27552, n27553,
         n27554, n27555, n27556, n27557, n27558, n27559, n27560, n27561,
         n27562, n27563, n27564, n27565, n27566, n27567, n27568, n27569,
         n27570, n27571, n27572, n27573, n27574, n27575, n27576, n27577,
         n27578, n27579, n27580, n27581, n27582, n27583, n27584, n27585,
         n27586, n27587, n27588, n27589, n27590, n27591, n27592, n27593,
         n27594, n27595, n27596, n27597, n27598, n27599, n27600, n27601,
         n27602, n27603, n27604, n27605, n27606, n27607, n27608, n27609,
         n27610, n27611, n27612, n27613, n27614, n27615, n27616, n27617,
         n27618, n27619, n27620, n27621, n27622, n27623, n27624, n27625,
         n27626, n27627, n27628, n27629, n27630, n27631, n27632, n27633,
         n27634, n27635, n27636, n27637, n27638, n27639, n27640, n27641,
         n27642, n27643, n27644, n27645, n27646, n27647, n27648, n27649,
         n27650, n27651, n27652, n27653, n27654, n27655, n27656, n27657,
         n27658, n27659, n27660, n27661, n27662, n27663, n27664, n27665,
         n27666, n27667, n27668, n27669, n27670, n27671, n27672, n27673,
         n27674, n27675, n27676, n27677, n27678, n27679, n27680, n27681,
         n27682, n27683, n27684, n27685, n27686, n27687, n27688, n27689,
         n27690, n27691, n27692, n27693, n27694, n27695, n27696, n27697,
         n27698, n27699, n27700, n27701, n27702, n27703, n27704, n27705,
         n27706, n27707, n27708, n27709, n27710, n27711, n27712, n27713,
         n27714, n27715, n27716, n27717, n27718, n27719, n27720, n27721,
         n27722, n27723, n27724, n27725, n27726, n27727, n27728, n27729,
         n27730, n27731, n27732, n27733, n27734, n27735, n27736, n27737,
         n27738, n27739, n27740, n27741, n27742, n27743, n27744, n27745,
         n27746, n27747, n27748, n27749, n27750, n27751, n27752, n27753,
         n27754, n27755, n27756, n27757, n27758, n27759, n27760, n27761,
         n27762, n27763, n27764, n27765, n27766, n27767, n27768, n27769,
         n27770, n27771, n27772, n27773, n27774, n27775, n27776, n27777,
         n27778, n27779, n27780, n27781, n27782, n27783, n27784, n27785,
         n27786, n27787, n27788, n27789, n27790, n27791, n27792, n27793,
         n27794, n27795, n27796, n27797, n27798, n27799, n27800, n27801,
         n27802, n27803, n27804, n27805, n27806, n27807, n27808, n27809,
         n27810, n27811, n27812, n27813, n27814, n27815, n27816, n27817,
         n27818, n27819, n27820, n27821, n27822, n27823, n27824, n27825,
         n27826, n27827, n27828, n27829, n27830, n27831, n27832, n27833,
         n27834, n27835, n27836, n27837, n27838, n27839, n27840, n27841,
         n27842, n27843, n27844, n27845, n27846, n27847, n27848, n27849,
         n27850, n27851, n27852, n27853, n27854, n27855, n27856, n27857,
         n27858, n27859, n27860, n27861, n27862, n27863, n27864, n27865,
         n27866, n27867, n27868, n27869, n27870, n27871, n27872, n27873,
         n27874, n27875, n27876, n27877, n27878, n27879, n27880, n27881,
         n27882, n27883, n27884, n27885, n27886, n27887, n27888, n27889,
         n27890, n27891, n27892, n27893, n27894, n27895, n27896, n27897,
         n27898, n27899, n27900, n27901, n27902, n27903, n27904, n27905,
         n27906, n27907, n27908, n27909, n27910, n27911, n27912, n27913,
         n27914, n27915, n27916, n27917, n27918, n27919, n27920, n27921,
         n27922, n27923, n27924, n27925, n27926, n27927, n27928, n27929,
         n27930, n27931, n27932, n27933, n27934, n27935, n27936, n27937,
         n27938, n27939, n27940, n27941, n27942, n27943, n27944, n27945,
         n27946, n27947, n27948, n27949, n27950, n27951, n27952, n27953,
         n27954, n27955, n27956, n27957, n27958, n27959, n27960, n27961,
         n27962, n27963, n27964, n27965, n27966, n27967, n27968, n27969,
         n27970, n27971, n27972, n27973, n27974, n27975, n27976, n27977,
         n27978, n27979, n27980, n27981, n27982, n27983, n27984, n27985,
         n27986, n27987, n27988, n27989, n27990, n27991, n27992, n27993,
         n27994, n27995, n27996, n27997, n27998, n27999, n28000, n28001,
         n28002, n28003, n28004, n28005, n28006, n28007, n28008, n28009,
         n28010, n28011, n28012, n28013, n28014, n28015, n28016, n28017,
         n28018, n28019, n28020, n28021, n28022, n28023, n28024, n28025,
         n28026, n28027, n28028, n28029, n28030, n28031, n28032, n28033,
         n28034, n28035, n28036, n28037, n28038, n28039, n28040, n28041,
         n28042, n28043, n28044, n28045, n28046, n28047, n28048, n28049,
         n28050, n28051, n28052, n28053, n28054, n28055, n28056, n28057,
         n28058, n28059, n28060, n28061, n28062, n28063, n28064, n28065,
         n28066, n28067, n28068, n28069, n28070, n28071, n28072, n28073,
         n28074, n28075, n28076, n28077, n28078, n28079, n28080, n28081,
         n28082, n28083, n28084, n28085, n28086, n28087, n28088, n28089,
         n28090, n28091, n28092, n28093, n28094, n28095, n28096, n28097,
         n28098, n28099, n28100, n28101, n28102, n28103, n28104, n28105,
         n28106, n28107, n28108, n28109, n28110, n28111, n28112, n28113,
         n28114, n28115, n28116, n28117, n28118, n28119, n28120, n28121,
         n28122, n28123, n28124, n28125, n28126, n28127, n28128, n28129,
         n28130, n28131, n28132, n28133, n28134, n28135, n28136, n28137,
         n28138, n28139, n28140, n28141, n28142, n28143, n28144, n28145,
         n28146, n28147, n28148, n28149, n28150, n28151, n28152, n28153,
         n28154, n28155, n28156, n28157, n28158, n28159, n28160, n28161,
         n28162, n28163, n28164, n28165, n28166, n28167, n28168, n28169,
         n28170, n28171, n28172, n28173, n28174, n28175, n28176, n28177,
         n28178, n28179, n28180, n28181, n28182, n28183, n28184, n28185,
         n28186, n28187, n28188, n28189, n28190, n28191, n28192, n28193,
         n28194, n28195, n28196, n28197, n28198, n28199, n28200, n28201,
         n28202, n28203, n28204, n28205, n28206, n28207, n28208, n28209,
         n28210, n28211, n28212, n28213, n28214, n28215, n28216, n28217,
         n28218, n28219, n28220, n28221, n28222, n28223, n28224, n28225,
         n28226, n28227, n28228, n28229, n28230, n28231, n28232, n28233,
         n28234, n28235, n28236, n28237, n28238, n28239, n28240, n28241,
         n28242, n28243, n28244, n28245, n28246, n28247, n28248, n28249,
         n28250, n28251, n28252, n28253, n28254, n28255, n28256, n28257,
         n28258, n28259, n28260, n28261, n28262, n28263, n28264, n28265,
         n28266, n28267, n28268, n28269, n28270, n28271, n28272, n28273,
         n28274, n28275, n28276, n28277, n28278, n28279, n28280, n28281,
         n28282, n28283, n28284, n28285, n28286, n28287, n28288, n28289,
         n28290, n28291, n28292, n28293, n28294, n28295, n28296, n28297,
         n28298, n28299, n28300, n28301, n28302, n28303, n28304, n28305,
         n28306, n28307, n28308, n28309, n28310, n28311, n28312, n28313,
         n28314, n28315, n28316, n28317, n28318, n28319, n28320, n28321,
         n28322, n28323, n28324, n28325, n28326, n28327, n28328, n28329,
         n28330, n28331, n28332, n28333, n28334, n28335, n28336, n28337,
         n28338, n28339, n28340, n28341, n28342, n28343, n28344, n28345,
         n28346, n28347, n28348, n28349, n28350, n28351, n28352, n28353,
         n28354, n28355, n28356, n28357, n28358, n28359, n28360, n28361,
         n28362, n28363, n28364, n28365, n28366, n28367, n28368, n28369,
         n28370, n28371, n28372, n28373, n28374, n28375, n28376, n28377,
         n28378, n28379, n28380, n28381, n28382, n28383, n28384, n28385,
         n28386, n28387, n28388, n28389, n28390, n28391, n28392, n28393,
         n28394, n28395, n28396, n28397, n28398, n28399, n28400, n28401,
         n28402, n28403, n28404, n28405, n28406, n28407, n28408, n28409,
         n28410, n28411, n28412, n28413, n28414, n28415, n28416, n28417,
         n28418, n28419, n28420, n28421, n28422, n28423, n28424, n28425,
         n28426, n28427, n28428, n28429, n28430, n28431, n28432, n28433,
         n28434, n28435, n28436, n28437, n28438, n28439, n28440, n28441,
         n28442, n28443, n28444, n28445, n28446, n28447, n28448, n28449,
         n28450, n28451, n28452, n28453, n28454, n28455, n28456, n28457,
         n28458, n28459, n28460, n28461, n28462, n28463, n28464, n28465,
         n28466, n28467, n28468, n28469, n28470, n28471, n28472, n28473,
         n28474, n28475, n28476, n28477, n28478, n28479, n28480, n28481,
         n28482, n28483, n28484, n28485, n28486, n28487, n28488, n28489,
         n28490, n28491, n28492, n28493, n28494, n28495, n28496, n28497,
         n28498, n28499, n28500, n28501, n28502, n28503, n28504, n28505,
         n28506, n28507, n28508, n28509, n28510, n28511, n28512, n28513,
         n28514, n28515, n28516, n28517, n28518, n28519, n28520, n28521,
         n28522, n28523, n28524, n28525, n28526, n28527, n28528, n28529,
         n28530, n28531, n28532, n28533, n28534, n28535, n28536, n28537,
         n28538, n28539, n28540, n28541, n28542, n28543, n28544, n28545,
         n28546, n28547, n28548, n28549, n28550, n28551, n28552, n28553,
         n28554, n28555, n28556, n28557, n28558, n28559, n28560, n28561,
         n28562, n28563, n28564, n28565, n28566, n28567, n28568, n28569,
         n28570, n28571, n28572, n28573, n28574, n28575, n28576, n28577,
         n28578, n28579, n28580, n28581, n28582, n28583, n28584, n28585,
         n28586, n28587, n28588, n28589, n28590, n28591, n28592, n28593,
         n28594, n28595, n28596, n28597, n28598, n28599, n28600, n28601,
         n28602, n28603, n28604, n28605, n28606, n28607, n28608, n28609,
         n28610, n28611, n28612, n28613, n28614, n28615, n28616, n28617,
         n28618, n28619, n28620, n28621, n28622, n28623, n28624, n28625,
         n28626, n28627, n28628, n28629, n28630, n28631, n28632, n28633,
         n28634, n28635, n28636, n28637, n28638, n28639, n28640, n28641,
         n28642, n28643, n28644, n28645, n28646, n28647, n28648, n28649,
         n28650, n28651, n28652, n28653, n28654, n28655, n28656, n28657,
         n28658, n28659, n28660, n28661, n28662, n28663, n28664, n28665,
         n28666, n28667, n28668, n28669, n28670, n28671, n28672, n28673,
         n28674, n28675, n28676, n28677, n28678, n28679, n28680, n28681,
         n28682, n28683, n28684, n28685, n28686, n28687, n28688, n28689,
         n28690, n28691, n28692, n28693, n28694, n28695, n28696, n28697,
         n28698, n28699, n28700, n28701, n28702, n28703, n28704, n28705,
         n28706, n28707, n28708, n28709, n28710, n28711, n28712, n28713,
         n28714, n28715, n28716, n28717, n28718, n28719, n28720, n28721,
         n28722, n28723, n28724, n28725, n28726, n28727, n28728, n28729,
         n28730, n28731, n28732, n28733, n28734, n28735, n28736, n28737,
         n28738, n28739, n28740, n28741, n28742, n28743, n28744, n28745,
         n28746, n28747, n28748, n28749, n28750, n28751, n28752, n28753,
         n28754, n28755, n28756, n28757, n28758, n28759, n28760, n28761,
         n28762, n28763, n28764, n28765, n28766, n28767, n28768, n28769,
         n28770, n28771, n28772, n28773, n28774, n28775, n28776, n28777,
         n28778, n28779, n28780, n28781, n28782, n28783, n28784, n28785,
         n28786, n28787, n28788, n28789, n28790, n28791, n28792, n28793,
         n28794, n28795, n28796, n28797, n28798, n28799, n28800, n28801,
         n28802, n28803, n28804, n28805, n28806, n28807, n28808, n28809,
         n28810, n28811, n28812, n28813, n28814, n28815, n28816, n28817,
         n28818, n28819, n28820, n28821, n28822, n28823, n28824, n28825,
         n28826, n28827, n28828, n28829, n28830, n28831, n28832, n28833,
         n28834, n28835, n28836, n28837, n28838, n28839, n28840, n28841,
         n28842, n28843, n28844, n28845, n28846, n28847, n28848, n28849,
         n28850, n28851, n28852, n28853, n28854, n28855, n28856, n28857,
         n28858, n28859, n28860, n28861, n28862, n28863, n28864, n28865,
         n28866, n28867, n28868, n28869, n28870, n28871, n28872, n28873,
         n28874, n28875, n28876, n28877, n28878, n28879, n28880, n28881,
         n28882, n28883, n28884, n28885, n28886, n28887, n28888, n28889,
         n28890, n28891, n28892, n28893, n28894, n28895, n28896, n28897,
         n28898, n28899, n28900, n28901, n28902, n28903, n28904, n28905,
         n28906, n28907, n28908, n28909, n28910, n28911, n28912, n28913,
         n28914, n28915, n28916, n28917, n28918, n28919, n28920, n28921,
         n28922, n28923, n28924, n28925, n28926, n28927, n28928, n28929,
         n28930, n28931, n28932, n28933, n28934, n28935, n28936, n28937,
         n28938, n28939, n28940, n28941, n28942, n28943, n28944, n28945,
         n28946, n28947, n28948, n28949, n28950, n28951, n28952, n28953,
         n28954, n28955, n28956, n28957, n28958, n28959, n28960, n28961,
         n28962, n28963, n28964, n28965, n28966, n28967, n28968, n28969,
         n28970, n28971, n28972, n28973, n28974, n28975, n28976, n28977,
         n28978, n28979, n28980, n28981, n28982, n28983, n28984, n28985,
         n28986, n28987, n28988, n28989, n28990, n28991, n28992, n28993,
         n28994, n28995, n28996, n28997, n28998, n28999, n29000, n29001,
         n29002, n29003, n29004, n29005, n29006, n29007, n29008, n29009,
         n29010, n29011, n29012, n29013, n29014, n29015, n29016, n29017,
         n29018, n29019, n29020, n29021, n29022, n29023, n29024, n29025,
         n29026, n29027, n29028, n29029, n29030, n29031, n29032, n29033,
         n29034, n29035, n29036, n29037, n29038, n29039, n29040, n29041,
         n29042, n29043, n29044, n29045, n29046, n29047, n29048, n29049,
         n29050, n29051, n29052, n29053, n29054, n29055, n29056, n29057,
         n29058, n29059, n29060, n29061, n29062, n29063, n29064, n29065,
         n29066, n29067, n29068, n29069, n29070, n29071, n29072, n29073,
         n29074, n29075, n29076, n29077, n29078, n29079, n29080, n29081,
         n29082, n29083, n29084, n29085, n29086, n29087, n29088, n29089,
         n29090, n29091, n29092, n29093, n29094, n29095, n29096, n29097,
         n29098, n29099, n29100, n29101, n29102, n29103, n29104, n29105,
         n29106, n29107, n29108, n29109, n29110, n29111, n29112, n29113,
         n29114, n29115, n29116, n29117, n29118, n29119, n29120, n29121,
         n29122, n29123, n29124, n29125, n29126, n29127, n29128, n29129,
         n29130, n29131, n29132, n29133, n29134, n29135, n29136, n29137,
         n29138, n29139, n29140, n29141, n29142, n29143, n29144, n29145,
         n29146, n29147, n29148, n29149, n29150, n29151, n29152, n29153,
         n29154, n29155, n29156, n29157, n29158, n29159, n29160, n29161,
         n29162, n29163, n29164, n29165, n29166, n29167, n29168, n29169,
         n29170, n29171, n29172, n29173, n29174, n29175, n29176, n29177,
         n29178, n29179, n29180, n29181, n29182, n29183, n29184, n29185,
         n29186, n29187, n29188, n29189, n29190, n29191, n29192, n29193,
         n29194, n29195, n29196, n29197, n29198, n29199, n29200, n29201,
         n29202, n29203, n29204, n29205, n29206, n29207, n29208, n29209,
         n29210, n29211, n29212, n29213, n29214, n29215, n29216, n29217,
         n29218, n29219, n29220, n29221, n29222, n29223, n29224, n29225,
         n29226, n29227, n29228, n29229, n29230, n29231, n29232, n29233,
         n29234, n29235, n29236, n29237, n29238, n29239, n29240, n29241,
         n29242, n29243, n29244, n29245, n29246, n29247, n29248, n29249,
         n29250, n29251, n29252, n29253, n29254, n29255, n29256, n29257,
         n29258, n29259, n29260, n29261, n29262, n29263, n29264, n29265,
         n29266, n29267, n29268, n29269, n29270, n29271, n29272, n29273,
         n29274, n29275, n29276, n29277, n29278, n29279, n29280, n29281,
         n29282, n29283, n29284, n29285, n29286, n29287, n29288, n29289,
         n29290, n29291, n29292, n29293, n29294, n29295, n29296, n29297,
         n29298, n29299, n29300, n29301, n29302, n29303, n29304, n29305,
         n29306, n29307, n29308, n29309, n29310, n29311, n29312, n29313,
         n29314, n29315, n29316, n29317, n29318, n29319, n29320, n29321,
         n29322, n29323, n29324, n29325, n29326, n29327, n29328, n29329,
         n29330, n29331, n29332, n29333, n29334, n29335, n29336, n29337,
         n29338, n29339, n29340, n29341, n29342, n29343, n29344, n29345,
         n29346, n29347, n29348, n29349, n29350, n29351, n29352, n29353,
         n29354, n29355, n29356, n29357, n29358, n29359, n29360, n29361,
         n29362, n29363, n29364, n29365, n29366, n29367, n29368, n29369,
         n29370, n29371, n29372, n29373, n29374, n29375, n29376, n29377,
         n29378, n29379, n29380, n29381, n29382, n29383, n29384, n29385,
         n29386, n29387, n29388, n29389, n29390, n29391, n29392, n29393,
         n29394, n29395, n29396, n29397, n29398, n29399, n29400, n29401,
         n29402, n29403, n29404, n29405, n29406, n29407, n29408, n29409,
         n29410, n29411, n29412, n29413, n29414, n29415, n29416, n29417,
         n29418, n29419, n29420, n29421, n29422, n29423, n29424, n29425,
         n29426, n29427, n29428, n29429, n29430, n29431, n29432, n29433,
         n29434, n29435, n29436, n29437, n29438, n29439, n29440, n29441,
         n29442, n29443, n29444, n29445, n29446, n29447, n29448, n29449,
         n29450, n29451, n29452, n29453, n29454, n29455, n29456, n29457,
         n29458, n29459, n29460, n29461, n29462, n29463, n29464, n29465,
         n29466, n29467, n29468, n29469, n29470, n29471, n29472, n29473,
         n29474, n29475, n29476, n29477, n29478, n29479, n29480, n29481,
         n29482, n29483, n29484, n29485, n29486, n29487, n29488, n29489,
         n29490, n29491, n29492, n29493, n29494, n29495, n29496, n29497,
         n29498, n29499, n29500, n29501, n29502, n29503, n29504, n29505,
         n29506, n29507, n29508, n29509, n29510, n29511, n29512, n29513,
         n29514, n29515, n29516, n29517, n29518, n29519, n29520, n29521,
         n29522, n29523, n29524, n29525, n29526, n29527, n29528, n29529,
         n29530, n29531, n29532, n29533, n29534, n29535, n29536, n29537,
         n29538, n29539, n29540, n29541, n29542, n29543, n29544, n29545,
         n29546, n29547, n29548, n29549, n29550, n29551, n29552, n29553,
         n29554, n29555, n29556, n29557, n29558, n29559, n29560, n29561,
         n29562, n29563, n29564, n29565, n29566, n29567, n29568, n29569,
         n29570, n29571, n29572, n29573, n29574, n29575, n29576, n29577,
         n29578, n29579, n29580, n29581, n29582, n29583, n29584, n29585,
         n29586, n29587, n29588, n29589, n29590, n29591, n29592, n29593,
         n29594, n29595, n29596, n29597, n29598, n29599, n29600, n29601,
         n29602, n29603, n29604, n29605, n29606, n29607, n29608, n29609,
         n29610, n29611, n29612, n29613, n29614, n29615, n29616, n29617,
         n29618, n29619, n29620, n29621, n29622, n29623, n29624, n29625,
         n29626, n29627, n29628, n29629, n29630, n29631, n29632, n29633,
         n29634, n29635, n29636, n29637, n29638, n29639, n29640, n29641,
         n29642, n29643, n29644, n29645, n29646, n29647, n29648, n29649,
         n29650, n29651, n29652, n29653, n29654, n29655, n29656, n29657,
         n29658, n29659, n29660, n29661, n29662, n29663, n29664, n29665,
         n29666, n29667, n29668, n29669, n29670, n29671, n29672, n29673,
         n29674, n29675, n29676, n29677, n29678, n29679, n29680, n29681,
         n29682, n29683, n29684, n29685, n29686, n29687, n29688, n29689,
         n29690, n29691, n29692, n29693, n29694, n29695, n29696, n29697,
         n29698, n29699, n29700, n29701, n29702, n29703, n29704, n29705,
         n29706, n29707, n29708, n29709, n29710, n29711, n29712, n29713,
         n29714, n29715, n29716, n29717, n29718, n29719, n29720, n29721,
         n29722, n29723, n29724, n29725, n29726, n29727, n29728, n29729,
         n29730, n29731, n29732, n29733, n29734, n29735, n29736, n29737,
         n29738, n29739, n29740, n29741, n29742, n29743, n29744, n29745,
         n29746, n29747, n29748, n29749, n29750, n29751, n29752, n29753,
         n29754, n29755, n29756, n29757, n29758, n29759, n29760, n29761,
         n29762, n29763, n29764, n29765, n29766, n29767, n29768, n29769,
         n29770, n29771, n29772, n29773, n29774, n29775, n29776, n29777,
         n29778, n29779, n29780, n29781, n29782, n29783, n29784, n29785,
         n29786, n29787, n29788, n29789, n29790, n29791, n29792, n29793,
         n29794, n29795, n29796, n29797, n29798, n29799, n29800, n29801,
         n29802, n29803, n29804, n29805, n29806, n29807, n29808, n29809,
         n29810, n29811, n29812, n29813, n29814, n29815, n29816, n29817,
         n29818, n29819, n29820, n29821, n29822, n29823, n29824, n29825,
         n29826, n29827, n29828, n29829, n29830, n29831, n29832, n29833,
         n29834, n29835, n29836, n29837, n29838, n29839, n29840, n29841,
         n29842, n29843, n29844, n29845, n29846, n29847, n29848, n29849,
         n29850, n29851, n29852, n29853, n29854, n29855, n29856, n29857,
         n29858, n29859, n29860, n29861, n29862, n29863, n29864, n29865,
         n29866, n29867, n29868, n29869, n29870, n29871, n29872, n29873,
         n29874, n29875, n29876, n29877, n29878, n29879, n29880, n29881,
         n29882, n29883, n29884, n29885, n29886, n29887, n29888, n29889,
         n29890, n29891, n29892, n29893, n29894, n29895, n29896, n29897,
         n29898, n29899, n29900, n29901, n29902, n29903, n29904, n29905,
         n29906, n29907, n29908, n29909, n29910, n29911, n29912, n29913,
         n29914, n29915, n29916, n29917, n29918, n29919, n29920, n29921,
         n29922, n29923, n29924, n29925, n29926, n29927, n29928, n29929,
         n29930, n29931, n29932, n29933, n29934, n29935, n29936, n29937,
         n29938, n29939, n29940, n29941, n29942, n29943, n29944, n29945,
         n29946, n29947, n29948, n29949, n29950, n29951, n29952, n29953,
         n29954, n29955, n29956, n29957, n29958, n29959, n29960, n29961,
         n29962, n29963, n29964, n29965, n29966, n29967, n29968, n29969,
         n29970, n29971, n29972, n29973, n29974, n29975, n29976, n29977,
         n29978, n29979, n29980, n29981, n29982, n29983, n29984, n29985,
         n29986, n29987, n29988, n29989, n29990, n29991, n29992, n29993,
         n29994, n29995, n29996, n29997, n29998, n29999, n30000, n30001,
         n30002, n30003, n30004, n30005, n30006, n30007, n30008, n30009,
         n30010, n30011, n30012, n30013, n30014, n30015, n30016, n30017,
         n30018, n30019, n30020, n30021, n30022, n30023, n30024, n30025,
         n30026, n30027, n30028, n30029, n30030, n30031, n30032, n30033,
         n30034, n30035, n30036, n30037, n30038, n30039, n30040, n30041,
         n30042, n30043, n30044, n30045, n30046, n30047, n30048, n30049,
         n30050, n30051, n30052, n30053, n30054, n30055, n30056, n30057,
         n30058, n30059, n30060, n30061, n30062, n30063, n30064, n30065,
         n30066, n30067, n30068, n30069, n30070, n30071, n30072, n30073,
         n30074, n30075, n30076, n30077, n30078, n30079, n30080, n30081,
         n30082, n30083, n30084, n30085, n30086, n30087, n30088, n30089,
         n30090, n30091, n30092, n30093, n30094, n30095, n30096, n30097,
         n30098, n30099, n30100, n30101, n30102, n30103, n30104, n30105,
         n30106, n30107, n30108, n30109, n30110, n30111, n30112, n30113,
         n30114, n30115, n30116, n30117, n30118, n30119, n30120, n30121,
         n30122, n30123, n30124, n30125, n30126, n30127, n30128, n30129,
         n30130, n30131, n30132, n30133, n30134, n30135, n30136, n30137,
         n30138, n30139, n30140, n30141, n30142, n30143, n30144, n30145,
         n30146, n30147, n30148, n30149, n30150, n30151, n30152, n30153,
         n30154, n30155, n30156, n30157, n30158, n30159, n30160, n30161,
         n30162, n30163, n30164, n30165, n30166, n30167, n30168, n30169,
         n30170, n30171, n30172, n30173, n30174, n30175, n30176, n30177,
         n30178, n30179, n30180, n30181, n30182, n30183, n30184, n30185,
         n30186, n30187, n30188, n30189, n30190, n30191, n30192, n30193,
         n30194, n30195, n30196, n30197, n30198, n30199, n30200, n30201,
         n30202, n30203, n30204, n30205, n30206, n30207, n30208, n30209,
         n30210, n30211, n30212, n30213, n30214, n30215, n30216, n30217,
         n30218, n30219, n30220, n30221, n30222, n30223, n30224, n30225,
         n30226, n30227, n30228, n30229, n30230, n30231, n30232, n30233,
         n30234, n30235, n30236, n30237, n30238, n30239, n30240, n30241,
         n30242, n30243, n30244, n30245, n30246, n30247, n30248, n30249,
         n30250, n30251, n30252, n30253, n30254, n30255, n30256, n30257,
         n30258, n30259, n30260, n30261, n30262, n30263, n30264, n30265,
         n30266, n30267, n30268, n30269, n30270, n30271, n30272, n30273,
         n30274, n30275, n30276, n30277, n30278, n30279, n30280, n30281,
         n30282, n30283, n30284, n30285, n30286, n30287, n30288, n30289,
         n30290, n30291, n30292, n30293, n30294, n30295, n30296, n30297,
         n30298, n30299, n30300, n30301, n30302, n30303, n30304, n30305,
         n30306, n30307, n30308, n30309, n30310, n30311, n30312, n30313,
         n30314, n30315, n30316, n30317, n30318, n30319, n30320, n30321,
         n30322, n30323, n30324, n30325, n30326, n30327, n30328, n30329,
         n30330, n30331, n30332, n30333, n30334, n30335, n30336, n30337,
         n30338, n30339, n30340, n30341, n30342, n30343, n30344, n30345,
         n30346, n30347, n30348, n30349, n30350, n30351, n30352, n30353,
         n30354, n30355, n30356, n30357, n30358, n30359, n30360, n30361,
         n30362, n30363, n30364, n30365, n30366, n30367, n30368, n30369,
         n30370, n30371, n30372, n30373, n30374, n30375, n30376, n30377,
         n30378, n30379, n30380, n30381, n30382, n30383, n30384, n30385,
         n30386, n30387, n30388, n30389, n30390, n30391, n30392, n30393,
         n30394, n30395, n30396, n30397, n30398, n30399, n30400, n30401,
         n30402, n30403, n30404, n30405, n30406, n30407, n30408, n30409,
         n30410, n30411, n30412, n30413, n30414, n30415, n30416, n30417,
         n30418, n30419, n30420, n30421, n30422, n30423, n30424, n30425,
         n30426, n30427, n30428, n30429, n30430, n30431, n30432, n30433,
         n30434, n30435, n30436, n30437, n30438, n30439, n30440, n30441,
         n30442, n30443, n30444, n30445, n30446, n30447, n30448, n30449,
         n30450, n30451, n30452, n30453, n30454, n30455, n30456, n30457,
         n30458, n30459, n30460, n30461, n30462, n30463, n30464, n30465,
         n30466, n30467, n30468, n30469, n30470, n30471, n30472, n30473,
         n30474, n30475, n30476, n30477, n30478, n30479, n30480, n30481,
         n30482, n30483, n30484, n30485, n30486, n30487, n30488, n30489,
         n30490, n30491, n30492, n30493, n30494, n30495, n30496, n30497,
         n30498, n30499, n30500, n30501, n30502, n30503, n30504, n30505,
         n30506, n30507, n30508, n30509, n30510, n30511, n30512, n30513,
         n30514, n30515, n30516, n30517, n30518, n30519, n30520, n30521,
         n30522, n30523, n30524, n30525, n30526, n30527, n30528, n30529,
         n30530, n30531, n30532, n30533, n30534, n30535, n30536, n30537,
         n30538, n30539, n30540, n30541, n30542, n30543, n30544, n30545,
         n30546, n30547, n30548, n30549, n30550, n30551, n30552, n30553,
         n30554, n30555, n30556, n30557, n30558, n30559, n30560, n30561,
         n30562, n30563, n30564, n30565, n30566, n30567, n30568, n30569,
         n30570, n30571, n30572, n30573, n30574, n30575, n30576, n30577,
         n30578, n30579, n30580, n30581, n30582, n30583, n30584, n30585,
         n30586, n30587, n30588, n30589, n30590, n30591, n30592, n30593,
         n30594, n30595, n30596, n30597, n30598, n30599, n30600, n30601,
         n30602, n30603, n30604, n30605, n30606, n30607, n30608, n30609,
         n30610, n30611, n30612, n30613, n30614, n30615, n30616, n30617,
         n30618, n30619, n30620, n30621, n30622, n30623, n30624, n30625,
         n30626, n30627, n30628, n30629, n30630, n30631, n30632, n30633,
         n30634, n30635, n30636, n30637, n30638, n30639, n30640, n30641,
         n30642, n30643, n30644, n30645, n30646, n30647, n30648, n30649,
         n30650, n30651, n30652, n30653, n30654, n30655, n30656, n30657,
         n30658, n30659, n30660, n30661, n30662, n30663, n30664, n30665,
         n30666, n30667, n30668, n30669, n30670, n30671, n30672, n30673,
         n30674, n30675, n30676, n30677, n30678, n30679, n30680, n30681,
         n30682, n30683, n30684, n30685, n30686, n30687, n30688, n30689,
         n30690, n30691, n30692, n30693, n30694, n30695, n30696, n30697,
         n30698, n30699, n30700, n30701, n30702, n30703, n30704, n30705,
         n30706, n30707, n30708, n30709, n30710, n30711, n30712, n30713,
         n30714, n30715, n30716, n30717, n30718, n30719, n30720, n30721,
         n30722, n30723, n30724, n30725, n30726, n30727, n30728, n30729,
         n30730, n30731, n30732, n30733, n30734, n30735, n30736, n30737,
         n30738, n30739, n30740, n30741, n30742, n30743, n30744, n30745,
         n30746, n30747, n30748, n30749, n30750, n30751, n30752, n30753,
         n30754, n30755, n30756, n30757, n30758, n30759, n30760, n30761,
         n30762, n30763, n30764, n30765, n30766, n30767, n30768, n30769,
         n30770, n30771, n30772, n30773, n30774, n30775, n30776, n30777,
         n30778, n30779, n30780, n30781, n30782, n30783, n30784, n30785,
         n30786, n30787, n30788, n30789, n30790, n30791, n30792, n30793,
         n30794, n30795, n30796, n30797, n30798, n30799, n30800, n30801,
         n30802, n30803, n30804, n30805, n30806, n30807, n30808, n30809,
         n30810, n30811, n30812, n30813, n30814, n30815, n30816, n30817,
         n30818, n30819, n30820, n30821, n30822, n30823, n30824, n30825,
         n30826, n30827, n30828, n30829, n30830, n30831, n30832, n30833,
         n30834, n30835, n30836, n30837, n30838, n30839, n30840, n30841,
         n30842, n30843, n30844, n30845, n30846, n30847, n30848, n30849,
         n30850, n30851, n30852, n30853, n30854, n30855, n30856, n30857,
         n30858, n30859, n30860, n30861, n30862, n30863, n30864, n30865,
         n30866, n30867, n30868, n30869, n30870, n30871, n30872, n30873,
         n30874, n30875, n30876, n30877, n30878, n30879, n30880, n30881,
         n30882, n30883, n30884, n30885, n30886, n30887, n30888, n30889,
         n30890, n30891, n30892, n30893, n30894, n30895, n30896, n30897,
         n30898, n30899, n30900, n30901, n30902, n30903, n30904, n30905,
         n30906, n30907, n30908, n30909, n30910, n30911, n30912, n30913,
         n30914, n30915, n30916, n30917, n30918, n30919, n30920, n30921,
         n30922, n30923, n30924, n30925, n30926, n30927, n30928, n30929,
         n30930, n30931, n30932, n30933, n30934, n30935, n30936, n30937,
         n30938, n30939, n30940, n30941, n30942, n30943, n30944, n30945,
         n30946, n30947, n30948, n30949, n30950, n30951, n30952, n30953,
         n30954, n30955, n30956, n30957, n30958, n30959, n30960, n30961,
         n30962, n30963, n30964, n30965, n30966, n30967, n30968, n30969,
         n30970, n30971, n30972, n30973, n30974, n30975, n30976, n30977,
         n30978, n30979, n30980, n30981, n30982, n30983, n30984, n30985,
         n30986, n30987, n30988, n30989, n30990, n30991, n30992, n30993,
         n30994, n30995, n30996, n30997, n30998, n30999, n31000, n31001,
         n31002, n31003, n31004, n31005, n31006, n31007, n31008, n31009,
         n31010, n31011, n31012, n31013, n31014, n31015, n31016, n31017,
         n31018, n31019, n31020, n31021, n31022, n31023, n31024, n31025,
         n31026, n31027, n31028, n31029, n31030, n31031, n31032, n31033,
         n31034, n31035, n31036, n31037, n31038, n31039, n31040, n31041,
         n31042, n31043, n31044, n31045, n31046, n31047, n31048, n31049,
         n31050, n31051, n31052, n31053, n31054, n31055, n31056, n31057,
         n31058, n31059, n31060, n31061, n31062, n31063, n31064, n31065,
         n31066, n31067, n31068, n31069, n31070, n31071, n31072, n31073,
         n31074, n31075, n31076, n31077, n31078, n31079, n31080, n31081,
         n31082, n31083, n31084, n31085, n31086, n31087, n31088, n31089,
         n31090, n31091, n31092, n31093, n31094, n31095, n31096, n31097,
         n31098, n31099, n31100, n31101, n31102, n31103, n31104, n31105,
         n31106, n31107, n31108, n31109, n31110, n31111, n31112, n31113,
         n31114, n31115, n31116, n31117, n31118, n31119, n31120, n31121,
         n31122, n31123, n31124, n31125, n31126, n31127, n31128, n31129,
         n31130, n31131, n31132, n31133, n31134, n31135, n31136, n31137,
         n31138, n31139, n31140, n31141, n31142, n31143, n31144, n31145,
         n31146, n31147, n31148, n31149, n31150, n31151, n31152, n31153,
         n31154, n31155, n31156, n31157, n31158, n31159, n31160, n31161,
         n31162, n31163, n31164, n31165, n31166, n31167, n31168, n31169,
         n31170, n31171, n31172, n31173, n31174, n31175, n31176, n31177,
         n31178, n31179, n31180, n31181, n31182, n31183, n31184, n31185,
         n31186, n31187, n31188, n31189, n31190, n31191, n31192, n31193,
         n31194, n31195, n31196, n31197, n31198, n31199, n31200, n31201,
         n31202, n31203, n31204, n31205, n31206, n31207, n31208, n31209,
         n31210, n31211, n31212, n31213, n31214, n31215, n31216, n31217,
         n31218, n31219, n31220, n31221, n31222, n31223, n31224, n31225,
         n31226, n31227, n31228, n31229, n31230, n31231, n31232, n31233,
         n31234, n31235, n31236, n31237, n31238, n31239, n31240, n31241,
         n31242, n31243, n31244, n31245, n31246, n31247, n31248, n31249,
         n31250, n31251, n31252, n31253, n31254, n31255, n31256, n31257,
         n31258, n31259, n31260, n31261, n31262, n31263, n31264, n31265,
         n31266, n31267, n31268, n31269, n31270, n31271, n31272, n31273,
         n31274, n31275, n31276, n31277, n31278, n31279, n31280, n31281,
         n31282, n31283, n31284, n31285, n31286, n31287, n31288, n31289,
         n31290, n31291, n31292, n31293, n31294, n31295, n31296, n31297,
         n31298, n31299, n31300, n31301, n31302, n31303, n31304, n31305,
         n31306, n31307, n31308, n31309, n31310, n31311, n31312, n31313,
         n31314, n31315, n31316, n31317, n31318, n31319, n31320, n31321,
         n31322, n31323, n31324, n31325, n31326, n31327, n31328, n31329,
         n31330, n31331, n31332, n31333, n31334, n31335, n31336, n31337,
         n31338, n31339, n31340, n31341, n31342, n31343, n31344, n31345,
         n31346, n31347, n31348, n31349, n31350, n31351, n31352, n31353,
         n31354, n31355, n31356, n31357, n31358, n31359, n31360, n31361,
         n31362, n31363, n31364, n31365, n31366, n31367, n31368, n31369,
         n31370, n31371, n31372, n31373, n31374, n31375, n31376, n31377,
         n31378, n31379, n31380, n31381, n31382, n31383, n31384, n31385,
         n31386, n31387, n31388, n31389, n31390, n31391, n31392, n31393,
         n31394, n31395, n31396, n31397, n31398, n31399, n31400, n31401,
         n31402, n31403, n31404, n31405, n31406, n31407, n31408, n31409,
         n31410, n31411, n31412, n31413, n31414, n31415, n31416, n31417,
         n31418, n31419, n31420, n31421, n31422, n31423, n31424, n31425,
         n31426, n31427, n31428, n31429, n31430, n31431, n31432, n31433,
         n31434, n31435, n31436, n31437, n31438, n31439, n31440, n31441,
         n31442, n31443, n31444, n31445, n31446, n31447, n31448, n31449,
         n31450, n31451, n31452, n31453, n31454, n31455, n31456, n31457,
         n31458, n31459, n31460, n31461, n31462, n31463, n31464, n31465,
         n31466, n31467, n31468, n31469, n31470, n31471, n31472, n31473,
         n31474, n31475, n31476, n31477, n31478, n31479, n31480, n31481,
         n31482, n31483, n31484, n31485, n31486, n31487, n31488, n31489,
         n31490, n31491, n31492, n31493, n31494, n31495, n31496, n31497,
         n31498, n31499, n31500, n31501, n31502, n31503, n31504, n31505,
         n31506, n31507, n31508, n31509, n31510, n31511, n31512, n31513,
         n31514, n31515, n31516, n31517, n31518, n31519, n31520, n31521,
         n31522, n31523, n31524, n31525, n31526, n31527, n31528, n31529,
         n31530, n31531, n31532, n31533, n31534, n31535, n31536, n31537,
         n31538, n31539, n31540, n31541, n31542, n31543, n31544, n31545,
         n31546, n31547, n31548, n31549, n31550, n31551, n31552, n31553,
         n31554, n31555, n31556, n31557, n31558, n31559, n31560, n31561,
         n31562, n31563, n31564, n31565, n31566, n31567, n31568, n31569,
         n31570, n31571, n31572, n31573, n31574, n31575, n31576, n31577,
         n31578, n31579, n31580, n31581, n31582, n31583, n31584, n31585,
         n31586, n31587, n31588, n31589, n31590, n31591, n31592, n31593,
         n31594, n31595, n31596, n31597, n31598, n31599, n31600, n31601,
         n31602, n31603, n31604, n31605, n31606, n31607, n31608, n31609,
         n31610, n31611, n31612, n31613, n31614, n31615, n31616, n31617,
         n31618, n31619, n31620, n31621, n31622, n31623, n31624, n31625,
         n31626, n31627, n31628, n31629, n31630, n31631, n31632, n31633,
         n31634, n31635, n31636, n31637, n31638, n31639, n31640, n31641,
         n31642, n31643, n31644, n31645, n31646, n31647, n31648, n31649,
         n31650, n31651, n31652, n31653, n31654, n31655, n31656, n31657,
         n31658, n31659, n31660, n31661, n31662, n31663, n31664, n31665,
         n31666, n31667, n31668, n31669, n31670, n31671, n31672, n31673,
         n31674, n31675, n31676, n31677, n31678, n31679, n31680, n31681,
         n31682, n31683, n31684, n31685, n31686, n31687, n31688, n31689,
         n31690, n31691, n31692, n31693, n31694, n31695, n31696, n31697,
         n31698, n31699, n31700, n31701, n31702, n31703, n31704, n31705,
         n31706, n31707, n31708, n31709, n31710, n31711, n31712, n31713,
         n31714, n31715, n31716, n31717, n31718, n31719, n31720, n31721,
         n31722, n31723, n31724, n31725, n31726, n31727, n31728, n31729,
         n31730, n31731, n31732, n31733, n31734, n31735, n31736, n31737,
         n31738, n31739, n31740, n31741, n31742, n31743, n31744, n31745,
         n31746, n31747, n31748, n31749, n31750, n31751, n31752, n31753,
         n31754, n31755, n31756, n31757, n31758, n31759, n31760, n31761,
         n31762, n31763, n31764, n31765, n31766, n31767, n31768, n31769,
         n31770, n31771, n31772, n31773, n31774, n31775, n31776, n31777,
         n31778, n31779, n31780, n31781, n31782, n31783, n31784, n31785,
         n31786, n31787, n31788, n31789, n31790, n31791, n31792, n31793,
         n31794, n31795, n31796, n31797, n31798, n31799, n31800, n31801,
         n31802, n31803, n31804, n31805, n31806, n31807, n31808, n31809,
         n31810, n31811, n31812, n31813, n31814, n31815, n31816, n31817,
         n31818, n31819, n31820, n31821, n31822, n31823, n31824, n31825,
         n31826, n31827, n31828, n31829, n31830, n31831;

  IV U2 ( .A(n27489), .Z(n2) );
  IV U3 ( .A(n27488), .Z(n3) );
  IV U4 ( .A(n27491), .Z(n4) );
  NOR U5 ( .A(n4), .B(n2), .Z(n5) );
  XOR U6 ( .A(n27491), .B(n2), .Z(n6) );
  NOR U7 ( .A(n6), .B(n3), .Z(n7) );
  NOR U8 ( .A(n5), .B(n7), .Z(n8) );
  IV U9 ( .A(n8), .Z(n28005) );
  IV U10 ( .A(n7916), .Z(n9) );
  NOR U11 ( .A(n7916), .B(n7915), .Z(n10) );
  NOR U12 ( .A(n7528), .B(n9), .Z(n11) );
  NOR U13 ( .A(n7918), .B(n11), .Z(n12) );
  NOR U14 ( .A(n10), .B(n12), .Z(n7634) );
  IV U15 ( .A(n16282), .Z(n13) );
  NOR U16 ( .A(n16282), .B(n16283), .Z(n14) );
  NOR U17 ( .A(n15435), .B(n13), .Z(n15) );
  NOR U18 ( .A(n16285), .B(n15), .Z(n16) );
  NOR U19 ( .A(n14), .B(n16), .Z(n15785) );
  IV U20 ( .A(n18956), .Z(n17) );
  IV U21 ( .A(n18958), .Z(n18) );
  IV U22 ( .A(n18955), .Z(n19) );
  NOR U23 ( .A(n19), .B(n17), .Z(n20) );
  XOR U24 ( .A(n18955), .B(n17), .Z(n21) );
  NOR U25 ( .A(n21), .B(n18), .Z(n22) );
  NOR U26 ( .A(n20), .B(n22), .Z(n23) );
  IV U27 ( .A(n23), .Z(n18851) );
  IV U28 ( .A(n23992), .Z(n24) );
  IV U29 ( .A(n23990), .Z(n25) );
  NOR U30 ( .A(n25), .B(n24), .Z(n26) );
  NOR U31 ( .A(n23990), .B(n23992), .Z(n27) );
  NOR U32 ( .A(n23989), .B(n27), .Z(n28) );
  NOR U33 ( .A(n26), .B(n28), .Z(n23875) );
  NOR U34 ( .A(n31469), .B(n31465), .Z(n29) );
  IV U35 ( .A(n29), .Z(n30) );
  IV U36 ( .A(n31468), .Z(n31) );
  NOR U37 ( .A(n31469), .B(n31), .Z(n32) );
  NOR U38 ( .A(n31477), .B(n32), .Z(n33) );
  IV U39 ( .A(n33), .Z(n34) );
  NOR U40 ( .A(n31463), .B(n31464), .Z(n35) );
  NOR U41 ( .A(n30), .B(n35), .Z(n36) );
  NOR U42 ( .A(n36), .B(n34), .Z(n37) );
  NOR U43 ( .A(n31472), .B(n28502), .Z(n38) );
  NOR U44 ( .A(n37), .B(n38), .Z(n39) );
  NOR U45 ( .A(n31476), .B(n39), .Z(n40) );
  NOR U46 ( .A(n40), .B(n31481), .Z(n41) );
  IV U47 ( .A(n41), .Z(n31486) );
  IV U48 ( .A(b[37]), .Z(n42) );
  IV U49 ( .A(b[38]), .Z(n43) );
  IV U50 ( .A(b[36]), .Z(n44) );
  IV U51 ( .A(b[35]), .Z(n45) );
  IV U52 ( .A(b[34]), .Z(n46) );
  IV U53 ( .A(b[33]), .Z(n47) );
  IV U54 ( .A(b[32]), .Z(n48) );
  IV U55 ( .A(b[31]), .Z(n49) );
  IV U56 ( .A(b[30]), .Z(n50) );
  IV U57 ( .A(b[29]), .Z(n51) );
  IV U58 ( .A(b[28]), .Z(n52) );
  IV U59 ( .A(b[27]), .Z(n53) );
  IV U60 ( .A(b[26]), .Z(n54) );
  IV U61 ( .A(b[25]), .Z(n55) );
  IV U62 ( .A(b[24]), .Z(n56) );
  IV U63 ( .A(b[23]), .Z(n57) );
  IV U64 ( .A(b[22]), .Z(n58) );
  IV U65 ( .A(b[21]), .Z(n59) );
  IV U66 ( .A(b[20]), .Z(n60) );
  IV U67 ( .A(b[19]), .Z(n61) );
  IV U68 ( .A(b[18]), .Z(n62) );
  IV U69 ( .A(b[17]), .Z(n63) );
  IV U70 ( .A(b[16]), .Z(n64) );
  IV U71 ( .A(b[15]), .Z(n65) );
  IV U72 ( .A(b[14]), .Z(n66) );
  IV U73 ( .A(b[13]), .Z(n67) );
  IV U74 ( .A(b[12]), .Z(n68) );
  IV U75 ( .A(b[11]), .Z(n69) );
  IV U76 ( .A(b[10]), .Z(n70) );
  IV U77 ( .A(b[9]), .Z(n71) );
  IV U78 ( .A(b[8]), .Z(n72) );
  IV U79 ( .A(b[7]), .Z(n73) );
  IV U80 ( .A(b[6]), .Z(n74) );
  IV U81 ( .A(b[5]), .Z(n75) );
  IV U82 ( .A(b[4]), .Z(n76) );
  IV U83 ( .A(b[3]), .Z(n77) );
  IV U84 ( .A(b[2]), .Z(n78) );
  IV U85 ( .A(a[38]), .Z(n79) );
  IV U86 ( .A(a[36]), .Z(n80) );
  IV U87 ( .A(a[34]), .Z(n81) );
  IV U88 ( .A(a[32]), .Z(n82) );
  IV U89 ( .A(a[30]), .Z(n83) );
  IV U90 ( .A(a[28]), .Z(n84) );
  IV U91 ( .A(a[26]), .Z(n85) );
  IV U92 ( .A(a[24]), .Z(n86) );
  IV U93 ( .A(a[20]), .Z(n87) );
  IV U94 ( .A(a[18]), .Z(n88) );
  IV U95 ( .A(a[14]), .Z(n89) );
  IV U96 ( .A(a[12]), .Z(n90) );
  IV U97 ( .A(a[6]), .Z(n91) );
  IV U98 ( .A(b[1]), .Z(n92) );
  IV U99 ( .A(a[0]), .Z(n93) );
  IV U100 ( .A(a[2]), .Z(n94) );
  IV U101 ( .A(a[3]), .Z(n95) );
  IV U102 ( .A(a[4]), .Z(n96) );
  IV U103 ( .A(a[5]), .Z(n97) );
  IV U104 ( .A(a[7]), .Z(n98) );
  IV U105 ( .A(a[8]), .Z(n99) );
  IV U106 ( .A(a[9]), .Z(n100) );
  IV U107 ( .A(a[10]), .Z(n101) );
  IV U108 ( .A(a[11]), .Z(n102) );
  IV U109 ( .A(a[13]), .Z(n103) );
  IV U110 ( .A(a[15]), .Z(n104) );
  IV U111 ( .A(a[16]), .Z(n105) );
  IV U112 ( .A(a[17]), .Z(n106) );
  IV U113 ( .A(a[19]), .Z(n107) );
  IV U114 ( .A(a[21]), .Z(n108) );
  IV U115 ( .A(a[22]), .Z(n109) );
  IV U116 ( .A(a[23]), .Z(n110) );
  IV U117 ( .A(a[25]), .Z(n111) );
  IV U118 ( .A(a[27]), .Z(n112) );
  IV U119 ( .A(a[29]), .Z(n113) );
  IV U120 ( .A(a[31]), .Z(n114) );
  IV U121 ( .A(a[33]), .Z(n115) );
  IV U122 ( .A(a[35]), .Z(n116) );
  IV U123 ( .A(a[37]), .Z(n117) );
  IV U124 ( .A(b[39]), .Z(n118) );
  IV U125 ( .A(a[39]), .Z(n119) );
  IV U126 ( .A(a[40]), .Z(n120) );
  IV U127 ( .A(b[40]), .Z(n121) );
  IV U128 ( .A(b[41]), .Z(n122) );
  IV U129 ( .A(a[41]), .Z(n123) );
  IV U130 ( .A(b[42]), .Z(n124) );
  IV U131 ( .A(a[42]), .Z(n125) );
  IV U132 ( .A(a[43]), .Z(n126) );
  IV U133 ( .A(b[43]), .Z(n127) );
  IV U134 ( .A(a[44]), .Z(n128) );
  IV U135 ( .A(b[44]), .Z(n129) );
  IV U136 ( .A(b[45]), .Z(n130) );
  IV U137 ( .A(a[45]), .Z(n131) );
  IV U138 ( .A(b[46]), .Z(n132) );
  IV U139 ( .A(a[46]), .Z(n133) );
  IV U140 ( .A(b[47]), .Z(n134) );
  IV U141 ( .A(a[47]), .Z(n135) );
  IV U142 ( .A(b[48]), .Z(n136) );
  IV U143 ( .A(a[48]), .Z(n137) );
  IV U144 ( .A(b[49]), .Z(n138) );
  IV U145 ( .A(a[49]), .Z(n139) );
  IV U146 ( .A(b[50]), .Z(n140) );
  IV U147 ( .A(a[50]), .Z(n141) );
  IV U148 ( .A(b[51]), .Z(n142) );
  IV U149 ( .A(a[51]), .Z(n143) );
  IV U150 ( .A(b[52]), .Z(n144) );
  IV U151 ( .A(a[52]), .Z(n145) );
  IV U152 ( .A(b[53]), .Z(n146) );
  IV U153 ( .A(a[53]), .Z(n147) );
  IV U154 ( .A(a[54]), .Z(n148) );
  IV U155 ( .A(b[54]), .Z(n149) );
  IV U156 ( .A(a[55]), .Z(n150) );
  IV U157 ( .A(b[55]), .Z(n151) );
  IV U158 ( .A(b[56]), .Z(n152) );
  IV U159 ( .A(a[56]), .Z(n153) );
  IV U160 ( .A(b[57]), .Z(n154) );
  IV U161 ( .A(a[57]), .Z(n155) );
  IV U162 ( .A(a[58]), .Z(n156) );
  IV U163 ( .A(b[58]), .Z(n157) );
  IV U164 ( .A(a[59]), .Z(n158) );
  IV U165 ( .A(b[59]), .Z(n159) );
  IV U166 ( .A(b[60]), .Z(n160) );
  IV U167 ( .A(a[60]), .Z(n161) );
  IV U168 ( .A(b[61]), .Z(n162) );
  IV U169 ( .A(a[61]), .Z(n163) );
  IV U170 ( .A(b[62]), .Z(n164) );
  IV U171 ( .A(a[62]), .Z(n165) );
  IV U172 ( .A(b[63]), .Z(n166) );
  IV U173 ( .A(a[63]), .Z(n167) );
  IV U174 ( .A(a[1]), .Z(n168) );
  IV U175 ( .A(b[0]), .Z(n169) );
  NOR U176 ( .A(n139), .B(n118), .Z(n6708) );
  NOR U177 ( .A(n131), .B(n122), .Z(n5649) );
  NOR U178 ( .A(n123), .B(n127), .Z(n4706) );
  NOR U179 ( .A(n79), .B(n130), .Z(n3981) );
  NOR U180 ( .A(n81), .B(n134), .Z(n3200) );
  NOR U181 ( .A(n104), .B(n146), .Z(n869) );
  NOR U182 ( .A(n91), .B(n157), .Z(n342) );
  NOR U183 ( .A(n97), .B(n159), .Z(n314) );
  NOR U184 ( .A(n96), .B(n160), .Z(n335) );
  NOR U185 ( .A(n95), .B(n162), .Z(n321) );
  NOR U186 ( .A(n166), .B(n168), .Z(n170) );
  IV U187 ( .A(n170), .Z(n330) );
  NOR U188 ( .A(n164), .B(n93), .Z(n328) );
  NOR U189 ( .A(n330), .B(n328), .Z(n171) );
  NOR U190 ( .A(n164), .B(n94), .Z(n329) );
  IV U191 ( .A(n329), .Z(n453) );
  XOR U192 ( .A(n171), .B(n453), .Z(n323) );
  XOR U193 ( .A(n321), .B(n323), .Z(n324) );
  NOR U194 ( .A(n93), .B(n166), .Z(n174) );
  NOR U195 ( .A(n164), .B(n168), .Z(n172) );
  IV U196 ( .A(n172), .Z(n177) );
  NOR U197 ( .A(n93), .B(n162), .Z(n211) );
  NOR U198 ( .A(n177), .B(n211), .Z(n173) );
  XOR U199 ( .A(n174), .B(n173), .Z(n197) );
  IV U200 ( .A(n197), .Z(n176) );
  NOR U201 ( .A(n94), .B(n162), .Z(n175) );
  IV U202 ( .A(n175), .Z(n198) );
  NOR U203 ( .A(n176), .B(n198), .Z(n181) );
  IV U204 ( .A(n211), .Z(n178) );
  NOR U205 ( .A(n178), .B(n177), .Z(n186) );
  IV U206 ( .A(n186), .Z(n179) );
  NOR U207 ( .A(b[63]), .B(n179), .Z(n180) );
  NOR U208 ( .A(n181), .B(n180), .Z(n325) );
  XOR U209 ( .A(n324), .B(n325), .Z(n182) );
  IV U210 ( .A(n182), .Z(n337) );
  XOR U211 ( .A(n335), .B(n337), .Z(n338) );
  NOR U212 ( .A(n93), .B(n160), .Z(n243) );
  IV U213 ( .A(n243), .Z(n184) );
  NOR U214 ( .A(n162), .B(n168), .Z(n187) );
  IV U215 ( .A(n187), .Z(n183) );
  NOR U216 ( .A(n184), .B(n183), .Z(n209) );
  IV U217 ( .A(n209), .Z(n185) );
  NOR U218 ( .A(n186), .B(n185), .Z(n193) );
  XOR U219 ( .A(n187), .B(n328), .Z(n188) );
  NOR U220 ( .A(n209), .B(n188), .Z(n189) );
  NOR U221 ( .A(n193), .B(n189), .Z(n190) );
  IV U222 ( .A(n190), .Z(n222) );
  NOR U223 ( .A(n94), .B(n160), .Z(n221) );
  IV U224 ( .A(n221), .Z(n191) );
  NOR U225 ( .A(n222), .B(n191), .Z(n192) );
  NOR U226 ( .A(n193), .B(n192), .Z(n195) );
  NOR U227 ( .A(n95), .B(n160), .Z(n196) );
  IV U228 ( .A(n196), .Z(n194) );
  NOR U229 ( .A(n195), .B(n194), .Z(n200) );
  XOR U230 ( .A(n196), .B(n195), .Z(n202) );
  XOR U231 ( .A(n198), .B(n197), .Z(n203) );
  NOR U232 ( .A(n202), .B(n203), .Z(n199) );
  NOR U233 ( .A(n200), .B(n199), .Z(n339) );
  XOR U234 ( .A(n338), .B(n339), .Z(n201) );
  IV U235 ( .A(n201), .Z(n316) );
  XOR U236 ( .A(n314), .B(n316), .Z(n317) );
  NOR U237 ( .A(n96), .B(n159), .Z(n226) );
  IV U238 ( .A(n226), .Z(n205) );
  XOR U239 ( .A(n203), .B(n202), .Z(n204) );
  IV U240 ( .A(n204), .Z(n225) );
  NOR U241 ( .A(n205), .B(n225), .Z(n228) );
  NOR U242 ( .A(n93), .B(n159), .Z(n284) );
  IV U243 ( .A(n284), .Z(n207) );
  NOR U244 ( .A(n160), .B(n168), .Z(n210) );
  IV U245 ( .A(n210), .Z(n206) );
  NOR U246 ( .A(n207), .B(n206), .Z(n241) );
  IV U247 ( .A(n241), .Z(n208) );
  NOR U248 ( .A(n209), .B(n208), .Z(n217) );
  XOR U249 ( .A(n211), .B(n210), .Z(n212) );
  NOR U250 ( .A(n241), .B(n212), .Z(n213) );
  NOR U251 ( .A(n217), .B(n213), .Z(n214) );
  IV U252 ( .A(n214), .Z(n254) );
  NOR U253 ( .A(n94), .B(n159), .Z(n253) );
  IV U254 ( .A(n253), .Z(n215) );
  NOR U255 ( .A(n254), .B(n215), .Z(n216) );
  NOR U256 ( .A(n217), .B(n216), .Z(n219) );
  NOR U257 ( .A(n95), .B(n159), .Z(n220) );
  IV U258 ( .A(n220), .Z(n218) );
  NOR U259 ( .A(n219), .B(n218), .Z(n224) );
  XOR U260 ( .A(n220), .B(n219), .Z(n234) );
  XOR U261 ( .A(n222), .B(n221), .Z(n235) );
  NOR U262 ( .A(n234), .B(n235), .Z(n223) );
  NOR U263 ( .A(n224), .B(n223), .Z(n230) );
  XOR U264 ( .A(n226), .B(n225), .Z(n231) );
  NOR U265 ( .A(n230), .B(n231), .Z(n227) );
  NOR U266 ( .A(n228), .B(n227), .Z(n318) );
  XOR U267 ( .A(n317), .B(n318), .Z(n229) );
  IV U268 ( .A(n229), .Z(n344) );
  XOR U269 ( .A(n342), .B(n344), .Z(n345) );
  XOR U270 ( .A(n231), .B(n230), .Z(n232) );
  IV U271 ( .A(n232), .Z(n261) );
  NOR U272 ( .A(n97), .B(n157), .Z(n262) );
  IV U273 ( .A(n262), .Z(n233) );
  NOR U274 ( .A(n261), .B(n233), .Z(n264) );
  NOR U275 ( .A(n96), .B(n157), .Z(n258) );
  IV U276 ( .A(n258), .Z(n237) );
  XOR U277 ( .A(n235), .B(n234), .Z(n236) );
  IV U278 ( .A(n236), .Z(n257) );
  NOR U279 ( .A(n237), .B(n257), .Z(n260) );
  NOR U280 ( .A(n93), .B(n157), .Z(n376) );
  IV U281 ( .A(n376), .Z(n239) );
  NOR U282 ( .A(n159), .B(n168), .Z(n242) );
  IV U283 ( .A(n242), .Z(n238) );
  NOR U284 ( .A(n239), .B(n238), .Z(n282) );
  IV U285 ( .A(n282), .Z(n240) );
  NOR U286 ( .A(n241), .B(n240), .Z(n249) );
  XOR U287 ( .A(n243), .B(n242), .Z(n244) );
  NOR U288 ( .A(n282), .B(n244), .Z(n245) );
  NOR U289 ( .A(n249), .B(n245), .Z(n246) );
  IV U290 ( .A(n246), .Z(n295) );
  NOR U291 ( .A(n94), .B(n157), .Z(n294) );
  IV U292 ( .A(n294), .Z(n247) );
  NOR U293 ( .A(n295), .B(n247), .Z(n248) );
  NOR U294 ( .A(n249), .B(n248), .Z(n251) );
  NOR U295 ( .A(n95), .B(n157), .Z(n252) );
  IV U296 ( .A(n252), .Z(n250) );
  NOR U297 ( .A(n251), .B(n250), .Z(n256) );
  XOR U298 ( .A(n252), .B(n251), .Z(n275) );
  XOR U299 ( .A(n254), .B(n253), .Z(n276) );
  NOR U300 ( .A(n275), .B(n276), .Z(n255) );
  NOR U301 ( .A(n256), .B(n255), .Z(n271) );
  XOR U302 ( .A(n258), .B(n257), .Z(n272) );
  NOR U303 ( .A(n271), .B(n272), .Z(n259) );
  NOR U304 ( .A(n260), .B(n259), .Z(n267) );
  XOR U305 ( .A(n262), .B(n261), .Z(n268) );
  NOR U306 ( .A(n267), .B(n268), .Z(n263) );
  NOR U307 ( .A(n264), .B(n263), .Z(n346) );
  XOR U308 ( .A(n345), .B(n346), .Z(n265) );
  IV U309 ( .A(n265), .Z(n310) );
  NOR U310 ( .A(n98), .B(n154), .Z(n311) );
  IV U311 ( .A(n311), .Z(n266) );
  NOR U312 ( .A(n310), .B(n266), .Z(n313) );
  XOR U313 ( .A(n268), .B(n267), .Z(n269) );
  IV U314 ( .A(n269), .Z(n306) );
  NOR U315 ( .A(n91), .B(n154), .Z(n307) );
  IV U316 ( .A(n307), .Z(n270) );
  NOR U317 ( .A(n306), .B(n270), .Z(n309) );
  XOR U318 ( .A(n272), .B(n271), .Z(n273) );
  IV U319 ( .A(n273), .Z(n302) );
  NOR U320 ( .A(n97), .B(n154), .Z(n303) );
  IV U321 ( .A(n303), .Z(n274) );
  NOR U322 ( .A(n302), .B(n274), .Z(n305) );
  NOR U323 ( .A(n96), .B(n154), .Z(n299) );
  IV U324 ( .A(n299), .Z(n278) );
  XOR U325 ( .A(n276), .B(n275), .Z(n277) );
  IV U326 ( .A(n277), .Z(n298) );
  NOR U327 ( .A(n278), .B(n298), .Z(n301) );
  NOR U328 ( .A(n93), .B(n154), .Z(n499) );
  IV U329 ( .A(n499), .Z(n280) );
  NOR U330 ( .A(n157), .B(n168), .Z(n283) );
  IV U331 ( .A(n283), .Z(n279) );
  NOR U332 ( .A(n280), .B(n279), .Z(n374) );
  IV U333 ( .A(n374), .Z(n281) );
  NOR U334 ( .A(n282), .B(n281), .Z(n290) );
  XOR U335 ( .A(n284), .B(n283), .Z(n285) );
  NOR U336 ( .A(n374), .B(n285), .Z(n286) );
  NOR U337 ( .A(n290), .B(n286), .Z(n287) );
  IV U338 ( .A(n287), .Z(n387) );
  NOR U339 ( .A(n94), .B(n154), .Z(n386) );
  IV U340 ( .A(n386), .Z(n288) );
  NOR U341 ( .A(n387), .B(n288), .Z(n289) );
  NOR U342 ( .A(n290), .B(n289), .Z(n292) );
  NOR U343 ( .A(n95), .B(n154), .Z(n293) );
  IV U344 ( .A(n293), .Z(n291) );
  NOR U345 ( .A(n292), .B(n291), .Z(n297) );
  XOR U346 ( .A(n293), .B(n292), .Z(n367) );
  XOR U347 ( .A(n295), .B(n294), .Z(n368) );
  NOR U348 ( .A(n367), .B(n368), .Z(n296) );
  NOR U349 ( .A(n297), .B(n296), .Z(n363) );
  XOR U350 ( .A(n299), .B(n298), .Z(n364) );
  NOR U351 ( .A(n363), .B(n364), .Z(n300) );
  NOR U352 ( .A(n301), .B(n300), .Z(n359) );
  XOR U353 ( .A(n303), .B(n302), .Z(n360) );
  NOR U354 ( .A(n359), .B(n360), .Z(n304) );
  NOR U355 ( .A(n305), .B(n304), .Z(n355) );
  XOR U356 ( .A(n307), .B(n306), .Z(n356) );
  NOR U357 ( .A(n355), .B(n356), .Z(n308) );
  NOR U358 ( .A(n309), .B(n308), .Z(n351) );
  XOR U359 ( .A(n311), .B(n310), .Z(n352) );
  NOR U360 ( .A(n351), .B(n352), .Z(n312) );
  NOR U361 ( .A(n313), .B(n312), .Z(n418) );
  IV U362 ( .A(n418), .Z(n349) );
  NOR U363 ( .A(n99), .B(n154), .Z(n414) );
  IV U364 ( .A(n314), .Z(n315) );
  NOR U365 ( .A(n316), .B(n315), .Z(n320) );
  NOR U366 ( .A(n318), .B(n317), .Z(n319) );
  NOR U367 ( .A(n320), .B(n319), .Z(n433) );
  NOR U368 ( .A(n91), .B(n159), .Z(n429) );
  IV U369 ( .A(n321), .Z(n322) );
  NOR U370 ( .A(n323), .B(n322), .Z(n327) );
  NOR U371 ( .A(n325), .B(n324), .Z(n326) );
  NOR U372 ( .A(n327), .B(n326), .Z(n448) );
  NOR U373 ( .A(n96), .B(n162), .Z(n444) );
  NOR U374 ( .A(n329), .B(n328), .Z(n331) );
  NOR U375 ( .A(n331), .B(n330), .Z(n332) );
  IV U376 ( .A(n332), .Z(n456) );
  NOR U377 ( .A(n95), .B(n164), .Z(n334) );
  NOR U378 ( .A(n94), .B(n166), .Z(n333) );
  XOR U379 ( .A(n334), .B(n333), .Z(n454) );
  XOR U380 ( .A(n456), .B(n454), .Z(n446) );
  XOR U381 ( .A(n444), .B(n446), .Z(n447) );
  XOR U382 ( .A(n448), .B(n447), .Z(n439) );
  IV U383 ( .A(n335), .Z(n336) );
  NOR U384 ( .A(n337), .B(n336), .Z(n341) );
  NOR U385 ( .A(n339), .B(n338), .Z(n340) );
  NOR U386 ( .A(n341), .B(n340), .Z(n438) );
  NOR U387 ( .A(n97), .B(n160), .Z(n436) );
  XOR U388 ( .A(n438), .B(n436), .Z(n441) );
  XOR U389 ( .A(n439), .B(n441), .Z(n431) );
  XOR U390 ( .A(n429), .B(n431), .Z(n432) );
  XOR U391 ( .A(n433), .B(n432), .Z(n424) );
  IV U392 ( .A(n342), .Z(n343) );
  NOR U393 ( .A(n344), .B(n343), .Z(n348) );
  NOR U394 ( .A(n346), .B(n345), .Z(n347) );
  NOR U395 ( .A(n348), .B(n347), .Z(n423) );
  NOR U396 ( .A(n98), .B(n157), .Z(n421) );
  XOR U397 ( .A(n423), .B(n421), .Z(n425) );
  XOR U398 ( .A(n424), .B(n425), .Z(n416) );
  XOR U399 ( .A(n414), .B(n416), .Z(n417) );
  XOR U400 ( .A(n349), .B(n417), .Z(n410) );
  NOR U401 ( .A(n100), .B(n152), .Z(n411) );
  IV U402 ( .A(n411), .Z(n350) );
  NOR U403 ( .A(n410), .B(n350), .Z(n413) );
  XOR U404 ( .A(n352), .B(n351), .Z(n353) );
  IV U405 ( .A(n353), .Z(n406) );
  NOR U406 ( .A(n99), .B(n152), .Z(n407) );
  IV U407 ( .A(n407), .Z(n354) );
  NOR U408 ( .A(n406), .B(n354), .Z(n409) );
  XOR U409 ( .A(n356), .B(n355), .Z(n357) );
  IV U410 ( .A(n357), .Z(n402) );
  NOR U411 ( .A(n98), .B(n152), .Z(n403) );
  IV U412 ( .A(n403), .Z(n358) );
  NOR U413 ( .A(n402), .B(n358), .Z(n405) );
  XOR U414 ( .A(n360), .B(n359), .Z(n361) );
  IV U415 ( .A(n361), .Z(n398) );
  NOR U416 ( .A(n91), .B(n152), .Z(n399) );
  IV U417 ( .A(n399), .Z(n362) );
  NOR U418 ( .A(n398), .B(n362), .Z(n401) );
  XOR U419 ( .A(n364), .B(n363), .Z(n365) );
  IV U420 ( .A(n365), .Z(n394) );
  NOR U421 ( .A(n97), .B(n152), .Z(n395) );
  IV U422 ( .A(n395), .Z(n366) );
  NOR U423 ( .A(n394), .B(n366), .Z(n397) );
  NOR U424 ( .A(n96), .B(n152), .Z(n391) );
  IV U425 ( .A(n391), .Z(n370) );
  XOR U426 ( .A(n368), .B(n367), .Z(n369) );
  IV U427 ( .A(n369), .Z(n390) );
  NOR U428 ( .A(n370), .B(n390), .Z(n393) );
  NOR U429 ( .A(n93), .B(n152), .Z(n641) );
  IV U430 ( .A(n641), .Z(n372) );
  NOR U431 ( .A(n154), .B(n168), .Z(n375) );
  IV U432 ( .A(n375), .Z(n371) );
  NOR U433 ( .A(n372), .B(n371), .Z(n497) );
  IV U434 ( .A(n497), .Z(n373) );
  NOR U435 ( .A(n374), .B(n373), .Z(n382) );
  XOR U436 ( .A(n376), .B(n375), .Z(n377) );
  NOR U437 ( .A(n497), .B(n377), .Z(n378) );
  NOR U438 ( .A(n382), .B(n378), .Z(n379) );
  IV U439 ( .A(n379), .Z(n510) );
  NOR U440 ( .A(n94), .B(n152), .Z(n509) );
  IV U441 ( .A(n509), .Z(n380) );
  NOR U442 ( .A(n510), .B(n380), .Z(n381) );
  NOR U443 ( .A(n382), .B(n381), .Z(n384) );
  NOR U444 ( .A(n95), .B(n152), .Z(n385) );
  IV U445 ( .A(n385), .Z(n383) );
  NOR U446 ( .A(n384), .B(n383), .Z(n389) );
  XOR U447 ( .A(n385), .B(n384), .Z(n490) );
  XOR U448 ( .A(n387), .B(n386), .Z(n491) );
  NOR U449 ( .A(n490), .B(n491), .Z(n388) );
  NOR U450 ( .A(n389), .B(n388), .Z(n486) );
  XOR U451 ( .A(n391), .B(n390), .Z(n487) );
  NOR U452 ( .A(n486), .B(n487), .Z(n392) );
  NOR U453 ( .A(n393), .B(n392), .Z(n482) );
  XOR U454 ( .A(n395), .B(n394), .Z(n483) );
  NOR U455 ( .A(n482), .B(n483), .Z(n396) );
  NOR U456 ( .A(n397), .B(n396), .Z(n478) );
  XOR U457 ( .A(n399), .B(n398), .Z(n479) );
  NOR U458 ( .A(n478), .B(n479), .Z(n400) );
  NOR U459 ( .A(n401), .B(n400), .Z(n474) );
  XOR U460 ( .A(n403), .B(n402), .Z(n475) );
  NOR U461 ( .A(n474), .B(n475), .Z(n404) );
  NOR U462 ( .A(n405), .B(n404), .Z(n470) );
  XOR U463 ( .A(n407), .B(n406), .Z(n471) );
  NOR U464 ( .A(n470), .B(n471), .Z(n408) );
  NOR U465 ( .A(n409), .B(n408), .Z(n466) );
  XOR U466 ( .A(n411), .B(n410), .Z(n467) );
  NOR U467 ( .A(n466), .B(n467), .Z(n412) );
  NOR U468 ( .A(n413), .B(n412), .Z(n549) );
  IV U469 ( .A(n549), .Z(n464) );
  NOR U470 ( .A(n101), .B(n152), .Z(n545) );
  IV U471 ( .A(n414), .Z(n415) );
  NOR U472 ( .A(n416), .B(n415), .Z(n420) );
  NOR U473 ( .A(n418), .B(n417), .Z(n419) );
  NOR U474 ( .A(n420), .B(n419), .Z(n556) );
  IV U475 ( .A(n556), .Z(n463) );
  NOR U476 ( .A(n100), .B(n154), .Z(n552) );
  IV U477 ( .A(n421), .Z(n422) );
  NOR U478 ( .A(n423), .B(n422), .Z(n428) );
  IV U479 ( .A(n424), .Z(n426) );
  NOR U480 ( .A(n426), .B(n425), .Z(n427) );
  NOR U481 ( .A(n428), .B(n427), .Z(n563) );
  IV U482 ( .A(n563), .Z(n462) );
  NOR U483 ( .A(n99), .B(n157), .Z(n559) );
  IV U484 ( .A(n429), .Z(n430) );
  NOR U485 ( .A(n431), .B(n430), .Z(n435) );
  NOR U486 ( .A(n433), .B(n432), .Z(n434) );
  NOR U487 ( .A(n435), .B(n434), .Z(n570) );
  IV U488 ( .A(n570), .Z(n461) );
  NOR U489 ( .A(n98), .B(n159), .Z(n566) );
  IV U490 ( .A(n436), .Z(n437) );
  NOR U491 ( .A(n438), .B(n437), .Z(n443) );
  IV U492 ( .A(n439), .Z(n440) );
  NOR U493 ( .A(n441), .B(n440), .Z(n442) );
  NOR U494 ( .A(n443), .B(n442), .Z(n577) );
  IV U495 ( .A(n577), .Z(n460) );
  IV U496 ( .A(n444), .Z(n445) );
  NOR U497 ( .A(n446), .B(n445), .Z(n450) );
  NOR U498 ( .A(n448), .B(n447), .Z(n449) );
  NOR U499 ( .A(n450), .B(n449), .Z(n451) );
  IV U500 ( .A(n451), .Z(n583) );
  NOR U501 ( .A(n97), .B(n162), .Z(n581) );
  NOR U502 ( .A(n166), .B(n95), .Z(n452) );
  IV U503 ( .A(n452), .Z(n590) );
  NOR U504 ( .A(n453), .B(n590), .Z(n458) );
  IV U505 ( .A(n454), .Z(n455) );
  NOR U506 ( .A(n456), .B(n455), .Z(n457) );
  NOR U507 ( .A(n458), .B(n457), .Z(n588) );
  NOR U508 ( .A(n164), .B(n96), .Z(n586) );
  XOR U509 ( .A(n588), .B(n586), .Z(n589) );
  XOR U510 ( .A(n590), .B(n589), .Z(n580) );
  XOR U511 ( .A(n581), .B(n580), .Z(n459) );
  IV U512 ( .A(n459), .Z(n582) );
  XOR U513 ( .A(n583), .B(n582), .Z(n575) );
  NOR U514 ( .A(n91), .B(n160), .Z(n573) );
  XOR U515 ( .A(n575), .B(n573), .Z(n576) );
  XOR U516 ( .A(n460), .B(n576), .Z(n568) );
  XOR U517 ( .A(n566), .B(n568), .Z(n569) );
  XOR U518 ( .A(n461), .B(n569), .Z(n561) );
  XOR U519 ( .A(n559), .B(n561), .Z(n562) );
  XOR U520 ( .A(n462), .B(n562), .Z(n554) );
  XOR U521 ( .A(n552), .B(n554), .Z(n555) );
  XOR U522 ( .A(n463), .B(n555), .Z(n547) );
  XOR U523 ( .A(n545), .B(n547), .Z(n548) );
  XOR U524 ( .A(n464), .B(n548), .Z(n541) );
  NOR U525 ( .A(n102), .B(n151), .Z(n542) );
  IV U526 ( .A(n542), .Z(n465) );
  NOR U527 ( .A(n541), .B(n465), .Z(n544) );
  IV U528 ( .A(n466), .Z(n468) );
  XOR U529 ( .A(n468), .B(n467), .Z(n537) );
  NOR U530 ( .A(n101), .B(n151), .Z(n538) );
  IV U531 ( .A(n538), .Z(n469) );
  NOR U532 ( .A(n537), .B(n469), .Z(n540) );
  XOR U533 ( .A(n471), .B(n470), .Z(n472) );
  IV U534 ( .A(n472), .Z(n533) );
  NOR U535 ( .A(n100), .B(n151), .Z(n534) );
  IV U536 ( .A(n534), .Z(n473) );
  NOR U537 ( .A(n533), .B(n473), .Z(n536) );
  XOR U538 ( .A(n475), .B(n474), .Z(n476) );
  IV U539 ( .A(n476), .Z(n529) );
  NOR U540 ( .A(n99), .B(n151), .Z(n530) );
  IV U541 ( .A(n530), .Z(n477) );
  NOR U542 ( .A(n529), .B(n477), .Z(n532) );
  XOR U543 ( .A(n479), .B(n478), .Z(n480) );
  IV U544 ( .A(n480), .Z(n525) );
  NOR U545 ( .A(n98), .B(n151), .Z(n526) );
  IV U546 ( .A(n526), .Z(n481) );
  NOR U547 ( .A(n525), .B(n481), .Z(n528) );
  XOR U548 ( .A(n483), .B(n482), .Z(n484) );
  IV U549 ( .A(n484), .Z(n521) );
  NOR U550 ( .A(n91), .B(n151), .Z(n522) );
  IV U551 ( .A(n522), .Z(n485) );
  NOR U552 ( .A(n521), .B(n485), .Z(n524) );
  XOR U553 ( .A(n487), .B(n486), .Z(n488) );
  IV U554 ( .A(n488), .Z(n517) );
  NOR U555 ( .A(n97), .B(n151), .Z(n518) );
  IV U556 ( .A(n518), .Z(n489) );
  NOR U557 ( .A(n517), .B(n489), .Z(n520) );
  NOR U558 ( .A(n96), .B(n151), .Z(n514) );
  IV U559 ( .A(n514), .Z(n493) );
  XOR U560 ( .A(n491), .B(n490), .Z(n492) );
  IV U561 ( .A(n492), .Z(n513) );
  NOR U562 ( .A(n493), .B(n513), .Z(n516) );
  NOR U563 ( .A(n93), .B(n151), .Z(n809) );
  IV U564 ( .A(n809), .Z(n495) );
  NOR U565 ( .A(n152), .B(n168), .Z(n498) );
  IV U566 ( .A(n498), .Z(n494) );
  NOR U567 ( .A(n495), .B(n494), .Z(n639) );
  IV U568 ( .A(n639), .Z(n496) );
  NOR U569 ( .A(n497), .B(n496), .Z(n505) );
  XOR U570 ( .A(n499), .B(n498), .Z(n500) );
  NOR U571 ( .A(n639), .B(n500), .Z(n501) );
  NOR U572 ( .A(n505), .B(n501), .Z(n502) );
  IV U573 ( .A(n502), .Z(n652) );
  NOR U574 ( .A(n94), .B(n151), .Z(n651) );
  IV U575 ( .A(n651), .Z(n503) );
  NOR U576 ( .A(n652), .B(n503), .Z(n504) );
  NOR U577 ( .A(n505), .B(n504), .Z(n507) );
  NOR U578 ( .A(n95), .B(n151), .Z(n508) );
  IV U579 ( .A(n508), .Z(n506) );
  NOR U580 ( .A(n507), .B(n506), .Z(n512) );
  XOR U581 ( .A(n508), .B(n507), .Z(n632) );
  XOR U582 ( .A(n510), .B(n509), .Z(n633) );
  NOR U583 ( .A(n632), .B(n633), .Z(n511) );
  NOR U584 ( .A(n512), .B(n511), .Z(n628) );
  XOR U585 ( .A(n514), .B(n513), .Z(n629) );
  NOR U586 ( .A(n628), .B(n629), .Z(n515) );
  NOR U587 ( .A(n516), .B(n515), .Z(n624) );
  XOR U588 ( .A(n518), .B(n517), .Z(n625) );
  NOR U589 ( .A(n624), .B(n625), .Z(n519) );
  NOR U590 ( .A(n520), .B(n519), .Z(n620) );
  XOR U591 ( .A(n522), .B(n521), .Z(n621) );
  NOR U592 ( .A(n620), .B(n621), .Z(n523) );
  NOR U593 ( .A(n524), .B(n523), .Z(n616) );
  XOR U594 ( .A(n526), .B(n525), .Z(n617) );
  NOR U595 ( .A(n616), .B(n617), .Z(n527) );
  NOR U596 ( .A(n528), .B(n527), .Z(n612) );
  XOR U597 ( .A(n530), .B(n529), .Z(n613) );
  NOR U598 ( .A(n612), .B(n613), .Z(n531) );
  NOR U599 ( .A(n532), .B(n531), .Z(n608) );
  XOR U600 ( .A(n534), .B(n533), .Z(n609) );
  NOR U601 ( .A(n608), .B(n609), .Z(n535) );
  NOR U602 ( .A(n536), .B(n535), .Z(n604) );
  XOR U603 ( .A(n538), .B(n537), .Z(n605) );
  NOR U604 ( .A(n604), .B(n605), .Z(n539) );
  NOR U605 ( .A(n540), .B(n539), .Z(n600) );
  XOR U606 ( .A(n542), .B(n541), .Z(n601) );
  NOR U607 ( .A(n600), .B(n601), .Z(n543) );
  NOR U608 ( .A(n544), .B(n543), .Z(n699) );
  IV U609 ( .A(n699), .Z(n598) );
  NOR U610 ( .A(n90), .B(n151), .Z(n695) );
  IV U611 ( .A(n545), .Z(n546) );
  NOR U612 ( .A(n547), .B(n546), .Z(n551) );
  NOR U613 ( .A(n549), .B(n548), .Z(n550) );
  NOR U614 ( .A(n551), .B(n550), .Z(n706) );
  IV U615 ( .A(n706), .Z(n597) );
  NOR U616 ( .A(n102), .B(n152), .Z(n702) );
  IV U617 ( .A(n552), .Z(n553) );
  NOR U618 ( .A(n554), .B(n553), .Z(n558) );
  NOR U619 ( .A(n556), .B(n555), .Z(n557) );
  NOR U620 ( .A(n558), .B(n557), .Z(n713) );
  IV U621 ( .A(n713), .Z(n596) );
  NOR U622 ( .A(n101), .B(n154), .Z(n709) );
  IV U623 ( .A(n559), .Z(n560) );
  NOR U624 ( .A(n561), .B(n560), .Z(n565) );
  NOR U625 ( .A(n563), .B(n562), .Z(n564) );
  NOR U626 ( .A(n565), .B(n564), .Z(n720) );
  IV U627 ( .A(n720), .Z(n595) );
  NOR U628 ( .A(n100), .B(n157), .Z(n716) );
  IV U629 ( .A(n566), .Z(n567) );
  NOR U630 ( .A(n568), .B(n567), .Z(n572) );
  NOR U631 ( .A(n570), .B(n569), .Z(n571) );
  NOR U632 ( .A(n572), .B(n571), .Z(n727) );
  IV U633 ( .A(n727), .Z(n594) );
  NOR U634 ( .A(n99), .B(n159), .Z(n723) );
  IV U635 ( .A(n573), .Z(n574) );
  NOR U636 ( .A(n575), .B(n574), .Z(n579) );
  NOR U637 ( .A(n577), .B(n576), .Z(n578) );
  NOR U638 ( .A(n579), .B(n578), .Z(n734) );
  IV U639 ( .A(n734), .Z(n593) );
  NOR U640 ( .A(n98), .B(n160), .Z(n730) );
  NOR U641 ( .A(n581), .B(n580), .Z(n585) );
  NOR U642 ( .A(n583), .B(n582), .Z(n584) );
  NOR U643 ( .A(n585), .B(n584), .Z(n740) );
  NOR U644 ( .A(n91), .B(n162), .Z(n737) );
  NOR U645 ( .A(n166), .B(n96), .Z(n748) );
  IV U646 ( .A(n586), .Z(n587) );
  NOR U647 ( .A(n588), .B(n587), .Z(n592) );
  NOR U648 ( .A(n590), .B(n589), .Z(n591) );
  NOR U649 ( .A(n592), .B(n591), .Z(n747) );
  NOR U650 ( .A(n164), .B(n97), .Z(n745) );
  XOR U651 ( .A(n747), .B(n745), .Z(n750) );
  XOR U652 ( .A(n748), .B(n750), .Z(n739) );
  XOR U653 ( .A(n737), .B(n739), .Z(n742) );
  XOR U654 ( .A(n740), .B(n742), .Z(n732) );
  XOR U655 ( .A(n730), .B(n732), .Z(n733) );
  XOR U656 ( .A(n593), .B(n733), .Z(n725) );
  XOR U657 ( .A(n723), .B(n725), .Z(n726) );
  XOR U658 ( .A(n594), .B(n726), .Z(n718) );
  XOR U659 ( .A(n716), .B(n718), .Z(n719) );
  XOR U660 ( .A(n595), .B(n719), .Z(n711) );
  XOR U661 ( .A(n709), .B(n711), .Z(n712) );
  XOR U662 ( .A(n596), .B(n712), .Z(n704) );
  XOR U663 ( .A(n702), .B(n704), .Z(n705) );
  XOR U664 ( .A(n597), .B(n705), .Z(n697) );
  XOR U665 ( .A(n695), .B(n697), .Z(n698) );
  XOR U666 ( .A(n598), .B(n698), .Z(n691) );
  NOR U667 ( .A(n103), .B(n149), .Z(n692) );
  IV U668 ( .A(n692), .Z(n599) );
  NOR U669 ( .A(n691), .B(n599), .Z(n694) );
  IV U670 ( .A(n600), .Z(n602) );
  XOR U671 ( .A(n602), .B(n601), .Z(n687) );
  NOR U672 ( .A(n90), .B(n149), .Z(n688) );
  IV U673 ( .A(n688), .Z(n603) );
  NOR U674 ( .A(n687), .B(n603), .Z(n690) );
  IV U675 ( .A(n604), .Z(n606) );
  XOR U676 ( .A(n606), .B(n605), .Z(n683) );
  NOR U677 ( .A(n102), .B(n149), .Z(n684) );
  IV U678 ( .A(n684), .Z(n607) );
  NOR U679 ( .A(n683), .B(n607), .Z(n686) );
  XOR U680 ( .A(n609), .B(n608), .Z(n610) );
  IV U681 ( .A(n610), .Z(n679) );
  NOR U682 ( .A(n101), .B(n149), .Z(n680) );
  IV U683 ( .A(n680), .Z(n611) );
  NOR U684 ( .A(n679), .B(n611), .Z(n682) );
  XOR U685 ( .A(n613), .B(n612), .Z(n614) );
  IV U686 ( .A(n614), .Z(n675) );
  NOR U687 ( .A(n100), .B(n149), .Z(n676) );
  IV U688 ( .A(n676), .Z(n615) );
  NOR U689 ( .A(n675), .B(n615), .Z(n678) );
  XOR U690 ( .A(n617), .B(n616), .Z(n618) );
  IV U691 ( .A(n618), .Z(n671) );
  NOR U692 ( .A(n99), .B(n149), .Z(n672) );
  IV U693 ( .A(n672), .Z(n619) );
  NOR U694 ( .A(n671), .B(n619), .Z(n674) );
  XOR U695 ( .A(n621), .B(n620), .Z(n622) );
  IV U696 ( .A(n622), .Z(n667) );
  NOR U697 ( .A(n98), .B(n149), .Z(n668) );
  IV U698 ( .A(n668), .Z(n623) );
  NOR U699 ( .A(n667), .B(n623), .Z(n670) );
  XOR U700 ( .A(n625), .B(n624), .Z(n626) );
  IV U701 ( .A(n626), .Z(n663) );
  NOR U702 ( .A(n91), .B(n149), .Z(n664) );
  IV U703 ( .A(n664), .Z(n627) );
  NOR U704 ( .A(n663), .B(n627), .Z(n666) );
  XOR U705 ( .A(n629), .B(n628), .Z(n630) );
  IV U706 ( .A(n630), .Z(n659) );
  NOR U707 ( .A(n97), .B(n149), .Z(n660) );
  IV U708 ( .A(n660), .Z(n631) );
  NOR U709 ( .A(n659), .B(n631), .Z(n662) );
  NOR U710 ( .A(n96), .B(n149), .Z(n656) );
  IV U711 ( .A(n656), .Z(n635) );
  XOR U712 ( .A(n633), .B(n632), .Z(n634) );
  IV U713 ( .A(n634), .Z(n655) );
  NOR U714 ( .A(n635), .B(n655), .Z(n658) );
  NOR U715 ( .A(n93), .B(n149), .Z(n1003) );
  IV U716 ( .A(n1003), .Z(n637) );
  NOR U717 ( .A(n151), .B(n168), .Z(n640) );
  IV U718 ( .A(n640), .Z(n636) );
  NOR U719 ( .A(n637), .B(n636), .Z(n807) );
  IV U720 ( .A(n807), .Z(n638) );
  NOR U721 ( .A(n639), .B(n638), .Z(n647) );
  XOR U722 ( .A(n641), .B(n640), .Z(n642) );
  NOR U723 ( .A(n807), .B(n642), .Z(n643) );
  NOR U724 ( .A(n647), .B(n643), .Z(n644) );
  IV U725 ( .A(n644), .Z(n820) );
  NOR U726 ( .A(n94), .B(n149), .Z(n819) );
  IV U727 ( .A(n819), .Z(n645) );
  NOR U728 ( .A(n820), .B(n645), .Z(n646) );
  NOR U729 ( .A(n647), .B(n646), .Z(n649) );
  NOR U730 ( .A(n95), .B(n149), .Z(n650) );
  IV U731 ( .A(n650), .Z(n648) );
  NOR U732 ( .A(n649), .B(n648), .Z(n654) );
  XOR U733 ( .A(n650), .B(n649), .Z(n800) );
  XOR U734 ( .A(n652), .B(n651), .Z(n801) );
  NOR U735 ( .A(n800), .B(n801), .Z(n653) );
  NOR U736 ( .A(n654), .B(n653), .Z(n796) );
  XOR U737 ( .A(n656), .B(n655), .Z(n797) );
  NOR U738 ( .A(n796), .B(n797), .Z(n657) );
  NOR U739 ( .A(n658), .B(n657), .Z(n792) );
  XOR U740 ( .A(n660), .B(n659), .Z(n793) );
  NOR U741 ( .A(n792), .B(n793), .Z(n661) );
  NOR U742 ( .A(n662), .B(n661), .Z(n788) );
  XOR U743 ( .A(n664), .B(n663), .Z(n789) );
  NOR U744 ( .A(n788), .B(n789), .Z(n665) );
  NOR U745 ( .A(n666), .B(n665), .Z(n784) );
  XOR U746 ( .A(n668), .B(n667), .Z(n785) );
  NOR U747 ( .A(n784), .B(n785), .Z(n669) );
  NOR U748 ( .A(n670), .B(n669), .Z(n780) );
  XOR U749 ( .A(n672), .B(n671), .Z(n781) );
  NOR U750 ( .A(n780), .B(n781), .Z(n673) );
  NOR U751 ( .A(n674), .B(n673), .Z(n776) );
  XOR U752 ( .A(n676), .B(n675), .Z(n777) );
  NOR U753 ( .A(n776), .B(n777), .Z(n677) );
  NOR U754 ( .A(n678), .B(n677), .Z(n772) );
  XOR U755 ( .A(n680), .B(n679), .Z(n773) );
  NOR U756 ( .A(n772), .B(n773), .Z(n681) );
  NOR U757 ( .A(n682), .B(n681), .Z(n768) );
  XOR U758 ( .A(n684), .B(n683), .Z(n769) );
  NOR U759 ( .A(n768), .B(n769), .Z(n685) );
  NOR U760 ( .A(n686), .B(n685), .Z(n764) );
  XOR U761 ( .A(n688), .B(n687), .Z(n765) );
  NOR U762 ( .A(n764), .B(n765), .Z(n689) );
  NOR U763 ( .A(n690), .B(n689), .Z(n760) );
  XOR U764 ( .A(n692), .B(n691), .Z(n761) );
  NOR U765 ( .A(n760), .B(n761), .Z(n693) );
  NOR U766 ( .A(n694), .B(n693), .Z(n877) );
  NOR U767 ( .A(n89), .B(n149), .Z(n873) );
  IV U768 ( .A(n695), .Z(n696) );
  NOR U769 ( .A(n697), .B(n696), .Z(n701) );
  NOR U770 ( .A(n699), .B(n698), .Z(n700) );
  NOR U771 ( .A(n701), .B(n700), .Z(n884) );
  IV U772 ( .A(n884), .Z(n759) );
  NOR U773 ( .A(n103), .B(n151), .Z(n880) );
  IV U774 ( .A(n702), .Z(n703) );
  NOR U775 ( .A(n704), .B(n703), .Z(n708) );
  NOR U776 ( .A(n706), .B(n705), .Z(n707) );
  NOR U777 ( .A(n708), .B(n707), .Z(n891) );
  IV U778 ( .A(n891), .Z(n758) );
  NOR U779 ( .A(n90), .B(n152), .Z(n887) );
  IV U780 ( .A(n709), .Z(n710) );
  NOR U781 ( .A(n711), .B(n710), .Z(n715) );
  NOR U782 ( .A(n713), .B(n712), .Z(n714) );
  NOR U783 ( .A(n715), .B(n714), .Z(n898) );
  IV U784 ( .A(n898), .Z(n757) );
  NOR U785 ( .A(n102), .B(n154), .Z(n894) );
  IV U786 ( .A(n716), .Z(n717) );
  NOR U787 ( .A(n718), .B(n717), .Z(n722) );
  NOR U788 ( .A(n720), .B(n719), .Z(n721) );
  NOR U789 ( .A(n722), .B(n721), .Z(n938) );
  IV U790 ( .A(n938), .Z(n756) );
  NOR U791 ( .A(n101), .B(n157), .Z(n934) );
  IV U792 ( .A(n723), .Z(n724) );
  NOR U793 ( .A(n725), .B(n724), .Z(n729) );
  NOR U794 ( .A(n727), .B(n726), .Z(n728) );
  NOR U795 ( .A(n729), .B(n728), .Z(n905) );
  IV U796 ( .A(n905), .Z(n755) );
  NOR U797 ( .A(n99), .B(n160), .Z(n927) );
  IV U798 ( .A(n730), .Z(n731) );
  NOR U799 ( .A(n732), .B(n731), .Z(n736) );
  NOR U800 ( .A(n734), .B(n733), .Z(n735) );
  NOR U801 ( .A(n736), .B(n735), .Z(n925) );
  XOR U802 ( .A(n927), .B(n925), .Z(n929) );
  IV U803 ( .A(n737), .Z(n738) );
  NOR U804 ( .A(n739), .B(n738), .Z(n744) );
  IV U805 ( .A(n740), .Z(n741) );
  NOR U806 ( .A(n742), .B(n741), .Z(n743) );
  NOR U807 ( .A(n744), .B(n743), .Z(n911) );
  NOR U808 ( .A(n98), .B(n162), .Z(n910) );
  IV U809 ( .A(n910), .Z(n754) );
  IV U810 ( .A(n745), .Z(n746) );
  NOR U811 ( .A(n747), .B(n746), .Z(n752) );
  IV U812 ( .A(n748), .Z(n749) );
  NOR U813 ( .A(n750), .B(n749), .Z(n751) );
  NOR U814 ( .A(n752), .B(n751), .Z(n918) );
  NOR U815 ( .A(n164), .B(n91), .Z(n916) );
  XOR U816 ( .A(n918), .B(n916), .Z(n920) );
  NOR U817 ( .A(n166), .B(n97), .Z(n753) );
  IV U818 ( .A(n753), .Z(n919) );
  XOR U819 ( .A(n920), .B(n919), .Z(n909) );
  XOR U820 ( .A(n754), .B(n909), .Z(n912) );
  XOR U821 ( .A(n911), .B(n912), .Z(n928) );
  XOR U822 ( .A(n929), .B(n928), .Z(n903) );
  NOR U823 ( .A(n100), .B(n159), .Z(n901) );
  XOR U824 ( .A(n903), .B(n901), .Z(n904) );
  XOR U825 ( .A(n755), .B(n904), .Z(n936) );
  XOR U826 ( .A(n934), .B(n936), .Z(n937) );
  XOR U827 ( .A(n756), .B(n937), .Z(n896) );
  XOR U828 ( .A(n894), .B(n896), .Z(n897) );
  XOR U829 ( .A(n757), .B(n897), .Z(n889) );
  XOR U830 ( .A(n887), .B(n889), .Z(n890) );
  XOR U831 ( .A(n758), .B(n890), .Z(n882) );
  XOR U832 ( .A(n880), .B(n882), .Z(n883) );
  XOR U833 ( .A(n759), .B(n883), .Z(n875) );
  XOR U834 ( .A(n873), .B(n875), .Z(n876) );
  XOR U835 ( .A(n877), .B(n876), .Z(n868) );
  NOR U836 ( .A(n869), .B(n868), .Z(n872) );
  IV U837 ( .A(n760), .Z(n762) );
  XOR U838 ( .A(n762), .B(n761), .Z(n863) );
  NOR U839 ( .A(n89), .B(n146), .Z(n864) );
  IV U840 ( .A(n864), .Z(n763) );
  NOR U841 ( .A(n863), .B(n763), .Z(n866) );
  IV U842 ( .A(n764), .Z(n766) );
  XOR U843 ( .A(n766), .B(n765), .Z(n859) );
  NOR U844 ( .A(n103), .B(n146), .Z(n860) );
  IV U845 ( .A(n860), .Z(n767) );
  NOR U846 ( .A(n859), .B(n767), .Z(n862) );
  IV U847 ( .A(n768), .Z(n770) );
  XOR U848 ( .A(n770), .B(n769), .Z(n855) );
  NOR U849 ( .A(n90), .B(n146), .Z(n856) );
  IV U850 ( .A(n856), .Z(n771) );
  NOR U851 ( .A(n855), .B(n771), .Z(n858) );
  XOR U852 ( .A(n773), .B(n772), .Z(n774) );
  IV U853 ( .A(n774), .Z(n851) );
  NOR U854 ( .A(n102), .B(n146), .Z(n852) );
  IV U855 ( .A(n852), .Z(n775) );
  NOR U856 ( .A(n851), .B(n775), .Z(n854) );
  NOR U857 ( .A(n101), .B(n146), .Z(n848) );
  IV U858 ( .A(n848), .Z(n779) );
  XOR U859 ( .A(n777), .B(n776), .Z(n778) );
  IV U860 ( .A(n778), .Z(n847) );
  NOR U861 ( .A(n779), .B(n847), .Z(n850) );
  XOR U862 ( .A(n781), .B(n780), .Z(n782) );
  IV U863 ( .A(n782), .Z(n843) );
  NOR U864 ( .A(n100), .B(n146), .Z(n844) );
  IV U865 ( .A(n844), .Z(n783) );
  NOR U866 ( .A(n843), .B(n783), .Z(n846) );
  XOR U867 ( .A(n785), .B(n784), .Z(n786) );
  IV U868 ( .A(n786), .Z(n839) );
  NOR U869 ( .A(n99), .B(n146), .Z(n840) );
  IV U870 ( .A(n840), .Z(n787) );
  NOR U871 ( .A(n839), .B(n787), .Z(n842) );
  XOR U872 ( .A(n789), .B(n788), .Z(n790) );
  IV U873 ( .A(n790), .Z(n835) );
  NOR U874 ( .A(n98), .B(n146), .Z(n836) );
  IV U875 ( .A(n836), .Z(n791) );
  NOR U876 ( .A(n835), .B(n791), .Z(n838) );
  XOR U877 ( .A(n793), .B(n792), .Z(n794) );
  IV U878 ( .A(n794), .Z(n831) );
  NOR U879 ( .A(n91), .B(n146), .Z(n832) );
  IV U880 ( .A(n832), .Z(n795) );
  NOR U881 ( .A(n831), .B(n795), .Z(n834) );
  XOR U882 ( .A(n797), .B(n796), .Z(n798) );
  IV U883 ( .A(n798), .Z(n827) );
  NOR U884 ( .A(n97), .B(n146), .Z(n828) );
  IV U885 ( .A(n828), .Z(n799) );
  NOR U886 ( .A(n827), .B(n799), .Z(n830) );
  NOR U887 ( .A(n96), .B(n146), .Z(n824) );
  IV U888 ( .A(n824), .Z(n803) );
  XOR U889 ( .A(n801), .B(n800), .Z(n802) );
  IV U890 ( .A(n802), .Z(n823) );
  NOR U891 ( .A(n803), .B(n823), .Z(n826) );
  NOR U892 ( .A(n93), .B(n146), .Z(n1212) );
  IV U893 ( .A(n1212), .Z(n805) );
  NOR U894 ( .A(n149), .B(n168), .Z(n808) );
  IV U895 ( .A(n808), .Z(n804) );
  NOR U896 ( .A(n805), .B(n804), .Z(n1001) );
  IV U897 ( .A(n1001), .Z(n806) );
  NOR U898 ( .A(n807), .B(n806), .Z(n815) );
  XOR U899 ( .A(n809), .B(n808), .Z(n810) );
  NOR U900 ( .A(n1001), .B(n810), .Z(n811) );
  NOR U901 ( .A(n815), .B(n811), .Z(n812) );
  IV U902 ( .A(n812), .Z(n1014) );
  NOR U903 ( .A(n94), .B(n146), .Z(n1013) );
  IV U904 ( .A(n1013), .Z(n813) );
  NOR U905 ( .A(n1014), .B(n813), .Z(n814) );
  NOR U906 ( .A(n815), .B(n814), .Z(n817) );
  NOR U907 ( .A(n95), .B(n146), .Z(n818) );
  IV U908 ( .A(n818), .Z(n816) );
  NOR U909 ( .A(n817), .B(n816), .Z(n822) );
  XOR U910 ( .A(n818), .B(n817), .Z(n994) );
  XOR U911 ( .A(n820), .B(n819), .Z(n995) );
  NOR U912 ( .A(n994), .B(n995), .Z(n821) );
  NOR U913 ( .A(n822), .B(n821), .Z(n990) );
  XOR U914 ( .A(n824), .B(n823), .Z(n991) );
  NOR U915 ( .A(n990), .B(n991), .Z(n825) );
  NOR U916 ( .A(n826), .B(n825), .Z(n986) );
  XOR U917 ( .A(n828), .B(n827), .Z(n987) );
  NOR U918 ( .A(n986), .B(n987), .Z(n829) );
  NOR U919 ( .A(n830), .B(n829), .Z(n982) );
  XOR U920 ( .A(n832), .B(n831), .Z(n983) );
  NOR U921 ( .A(n982), .B(n983), .Z(n833) );
  NOR U922 ( .A(n834), .B(n833), .Z(n978) );
  XOR U923 ( .A(n836), .B(n835), .Z(n979) );
  NOR U924 ( .A(n978), .B(n979), .Z(n837) );
  NOR U925 ( .A(n838), .B(n837), .Z(n974) );
  XOR U926 ( .A(n840), .B(n839), .Z(n975) );
  NOR U927 ( .A(n974), .B(n975), .Z(n841) );
  NOR U928 ( .A(n842), .B(n841), .Z(n970) );
  XOR U929 ( .A(n844), .B(n843), .Z(n971) );
  NOR U930 ( .A(n970), .B(n971), .Z(n845) );
  NOR U931 ( .A(n846), .B(n845), .Z(n966) );
  XOR U932 ( .A(n848), .B(n847), .Z(n967) );
  NOR U933 ( .A(n966), .B(n967), .Z(n849) );
  NOR U934 ( .A(n850), .B(n849), .Z(n962) );
  XOR U935 ( .A(n852), .B(n851), .Z(n963) );
  NOR U936 ( .A(n962), .B(n963), .Z(n853) );
  NOR U937 ( .A(n854), .B(n853), .Z(n958) );
  XOR U938 ( .A(n856), .B(n855), .Z(n959) );
  NOR U939 ( .A(n958), .B(n959), .Z(n857) );
  NOR U940 ( .A(n858), .B(n857), .Z(n954) );
  XOR U941 ( .A(n860), .B(n859), .Z(n955) );
  NOR U942 ( .A(n954), .B(n955), .Z(n861) );
  NOR U943 ( .A(n862), .B(n861), .Z(n950) );
  XOR U944 ( .A(n864), .B(n863), .Z(n951) );
  NOR U945 ( .A(n950), .B(n951), .Z(n865) );
  NOR U946 ( .A(n866), .B(n865), .Z(n867) );
  IV U947 ( .A(n867), .Z(n948) );
  XOR U948 ( .A(n869), .B(n868), .Z(n870) );
  IV U949 ( .A(n870), .Z(n947) );
  NOR U950 ( .A(n948), .B(n947), .Z(n871) );
  NOR U951 ( .A(n872), .B(n871), .Z(n1076) );
  NOR U952 ( .A(n105), .B(n146), .Z(n1073) );
  IV U953 ( .A(n873), .Z(n874) );
  NOR U954 ( .A(n875), .B(n874), .Z(n879) );
  NOR U955 ( .A(n877), .B(n876), .Z(n878) );
  NOR U956 ( .A(n879), .B(n878), .Z(n1085) );
  IV U957 ( .A(n1085), .Z(n945) );
  NOR U958 ( .A(n104), .B(n149), .Z(n1081) );
  IV U959 ( .A(n880), .Z(n881) );
  NOR U960 ( .A(n882), .B(n881), .Z(n886) );
  NOR U961 ( .A(n884), .B(n883), .Z(n885) );
  NOR U962 ( .A(n886), .B(n885), .Z(n1092) );
  IV U963 ( .A(n1092), .Z(n944) );
  NOR U964 ( .A(n89), .B(n151), .Z(n1088) );
  IV U965 ( .A(n887), .Z(n888) );
  NOR U966 ( .A(n889), .B(n888), .Z(n893) );
  NOR U967 ( .A(n891), .B(n890), .Z(n892) );
  NOR U968 ( .A(n893), .B(n892), .Z(n1099) );
  IV U969 ( .A(n1099), .Z(n943) );
  NOR U970 ( .A(n103), .B(n152), .Z(n1095) );
  IV U971 ( .A(n894), .Z(n895) );
  NOR U972 ( .A(n896), .B(n895), .Z(n900) );
  NOR U973 ( .A(n898), .B(n897), .Z(n899) );
  NOR U974 ( .A(n900), .B(n899), .Z(n1106) );
  IV U975 ( .A(n1106), .Z(n942) );
  NOR U976 ( .A(n90), .B(n154), .Z(n1102) );
  IV U977 ( .A(n901), .Z(n902) );
  NOR U978 ( .A(n903), .B(n902), .Z(n907) );
  NOR U979 ( .A(n905), .B(n904), .Z(n906) );
  NOR U980 ( .A(n907), .B(n906), .Z(n908) );
  IV U981 ( .A(n908), .Z(n1112) );
  NOR U982 ( .A(n101), .B(n159), .Z(n1110) );
  NOR U983 ( .A(n910), .B(n909), .Z(n915) );
  IV U984 ( .A(n911), .Z(n913) );
  NOR U985 ( .A(n913), .B(n912), .Z(n914) );
  NOR U986 ( .A(n915), .B(n914), .Z(n1125) );
  NOR U987 ( .A(n99), .B(n162), .Z(n1123) );
  IV U988 ( .A(n1123), .Z(n924) );
  IV U989 ( .A(n916), .Z(n917) );
  NOR U990 ( .A(n918), .B(n917), .Z(n922) );
  NOR U991 ( .A(n920), .B(n919), .Z(n921) );
  NOR U992 ( .A(n922), .B(n921), .Z(n1130) );
  NOR U993 ( .A(n164), .B(n98), .Z(n1128) );
  XOR U994 ( .A(n1130), .B(n1128), .Z(n1132) );
  NOR U995 ( .A(n166), .B(n91), .Z(n923) );
  IV U996 ( .A(n923), .Z(n1131) );
  XOR U997 ( .A(n1132), .B(n1131), .Z(n1122) );
  XOR U998 ( .A(n924), .B(n1122), .Z(n1124) );
  XOR U999 ( .A(n1125), .B(n1124), .Z(n1117) );
  IV U1000 ( .A(n925), .Z(n926) );
  NOR U1001 ( .A(n927), .B(n926), .Z(n931) );
  NOR U1002 ( .A(n929), .B(n928), .Z(n930) );
  NOR U1003 ( .A(n931), .B(n930), .Z(n1115) );
  XOR U1004 ( .A(n1117), .B(n1115), .Z(n1119) );
  NOR U1005 ( .A(n100), .B(n160), .Z(n932) );
  IV U1006 ( .A(n932), .Z(n1118) );
  XOR U1007 ( .A(n1119), .B(n1118), .Z(n1109) );
  XOR U1008 ( .A(n1110), .B(n1109), .Z(n933) );
  IV U1009 ( .A(n933), .Z(n1111) );
  XOR U1010 ( .A(n1112), .B(n1111), .Z(n1142) );
  IV U1011 ( .A(n934), .Z(n935) );
  NOR U1012 ( .A(n936), .B(n935), .Z(n940) );
  NOR U1013 ( .A(n938), .B(n937), .Z(n939) );
  NOR U1014 ( .A(n940), .B(n939), .Z(n1140) );
  NOR U1015 ( .A(n102), .B(n157), .Z(n1138) );
  XOR U1016 ( .A(n1140), .B(n1138), .Z(n1141) );
  XOR U1017 ( .A(n1142), .B(n1141), .Z(n941) );
  IV U1018 ( .A(n941), .Z(n1104) );
  XOR U1019 ( .A(n1102), .B(n1104), .Z(n1105) );
  XOR U1020 ( .A(n942), .B(n1105), .Z(n1097) );
  XOR U1021 ( .A(n1095), .B(n1097), .Z(n1098) );
  XOR U1022 ( .A(n943), .B(n1098), .Z(n1090) );
  XOR U1023 ( .A(n1088), .B(n1090), .Z(n1091) );
  XOR U1024 ( .A(n944), .B(n1091), .Z(n1083) );
  XOR U1025 ( .A(n1081), .B(n1083), .Z(n1084) );
  XOR U1026 ( .A(n945), .B(n1084), .Z(n1075) );
  XOR U1027 ( .A(n1073), .B(n1075), .Z(n1078) );
  XOR U1028 ( .A(n1076), .B(n1078), .Z(n1069) );
  NOR U1029 ( .A(n106), .B(n144), .Z(n1070) );
  IV U1030 ( .A(n1070), .Z(n946) );
  NOR U1031 ( .A(n1069), .B(n946), .Z(n1072) );
  XOR U1032 ( .A(n948), .B(n947), .Z(n1066) );
  NOR U1033 ( .A(n105), .B(n144), .Z(n1065) );
  IV U1034 ( .A(n1065), .Z(n949) );
  NOR U1035 ( .A(n1066), .B(n949), .Z(n1068) );
  IV U1036 ( .A(n950), .Z(n952) );
  XOR U1037 ( .A(n952), .B(n951), .Z(n1061) );
  NOR U1038 ( .A(n104), .B(n144), .Z(n1062) );
  IV U1039 ( .A(n1062), .Z(n953) );
  NOR U1040 ( .A(n1061), .B(n953), .Z(n1064) );
  IV U1041 ( .A(n954), .Z(n956) );
  XOR U1042 ( .A(n956), .B(n955), .Z(n1057) );
  NOR U1043 ( .A(n89), .B(n144), .Z(n1058) );
  IV U1044 ( .A(n1058), .Z(n957) );
  NOR U1045 ( .A(n1057), .B(n957), .Z(n1060) );
  IV U1046 ( .A(n958), .Z(n960) );
  XOR U1047 ( .A(n960), .B(n959), .Z(n1053) );
  NOR U1048 ( .A(n103), .B(n144), .Z(n1054) );
  IV U1049 ( .A(n1054), .Z(n961) );
  NOR U1050 ( .A(n1053), .B(n961), .Z(n1056) );
  XOR U1051 ( .A(n963), .B(n962), .Z(n964) );
  IV U1052 ( .A(n964), .Z(n1049) );
  NOR U1053 ( .A(n90), .B(n144), .Z(n1050) );
  IV U1054 ( .A(n1050), .Z(n965) );
  NOR U1055 ( .A(n1049), .B(n965), .Z(n1052) );
  XOR U1056 ( .A(n967), .B(n966), .Z(n968) );
  IV U1057 ( .A(n968), .Z(n1045) );
  NOR U1058 ( .A(n102), .B(n144), .Z(n1046) );
  IV U1059 ( .A(n1046), .Z(n969) );
  NOR U1060 ( .A(n1045), .B(n969), .Z(n1048) );
  XOR U1061 ( .A(n971), .B(n970), .Z(n972) );
  IV U1062 ( .A(n972), .Z(n1041) );
  NOR U1063 ( .A(n101), .B(n144), .Z(n1042) );
  IV U1064 ( .A(n1042), .Z(n973) );
  NOR U1065 ( .A(n1041), .B(n973), .Z(n1044) );
  IV U1066 ( .A(n974), .Z(n976) );
  XOR U1067 ( .A(n976), .B(n975), .Z(n1037) );
  NOR U1068 ( .A(n100), .B(n144), .Z(n1038) );
  IV U1069 ( .A(n1038), .Z(n977) );
  NOR U1070 ( .A(n1037), .B(n977), .Z(n1040) );
  XOR U1071 ( .A(n979), .B(n978), .Z(n980) );
  IV U1072 ( .A(n980), .Z(n1033) );
  NOR U1073 ( .A(n99), .B(n144), .Z(n1034) );
  IV U1074 ( .A(n1034), .Z(n981) );
  NOR U1075 ( .A(n1033), .B(n981), .Z(n1036) );
  XOR U1076 ( .A(n983), .B(n982), .Z(n984) );
  IV U1077 ( .A(n984), .Z(n1029) );
  NOR U1078 ( .A(n98), .B(n144), .Z(n1030) );
  IV U1079 ( .A(n1030), .Z(n985) );
  NOR U1080 ( .A(n1029), .B(n985), .Z(n1032) );
  XOR U1081 ( .A(n987), .B(n986), .Z(n988) );
  IV U1082 ( .A(n988), .Z(n1025) );
  NOR U1083 ( .A(n91), .B(n144), .Z(n1026) );
  IV U1084 ( .A(n1026), .Z(n989) );
  NOR U1085 ( .A(n1025), .B(n989), .Z(n1028) );
  XOR U1086 ( .A(n991), .B(n990), .Z(n992) );
  IV U1087 ( .A(n992), .Z(n1021) );
  NOR U1088 ( .A(n97), .B(n144), .Z(n1022) );
  IV U1089 ( .A(n1022), .Z(n993) );
  NOR U1090 ( .A(n1021), .B(n993), .Z(n1024) );
  NOR U1091 ( .A(n96), .B(n144), .Z(n1018) );
  IV U1092 ( .A(n1018), .Z(n997) );
  XOR U1093 ( .A(n995), .B(n994), .Z(n996) );
  IV U1094 ( .A(n996), .Z(n1017) );
  NOR U1095 ( .A(n997), .B(n1017), .Z(n1020) );
  NOR U1096 ( .A(n93), .B(n144), .Z(n1448) );
  IV U1097 ( .A(n1448), .Z(n999) );
  NOR U1098 ( .A(n146), .B(n168), .Z(n1002) );
  IV U1099 ( .A(n1002), .Z(n998) );
  NOR U1100 ( .A(n999), .B(n998), .Z(n1210) );
  IV U1101 ( .A(n1210), .Z(n1000) );
  NOR U1102 ( .A(n1001), .B(n1000), .Z(n1009) );
  XOR U1103 ( .A(n1003), .B(n1002), .Z(n1004) );
  NOR U1104 ( .A(n1210), .B(n1004), .Z(n1005) );
  NOR U1105 ( .A(n1009), .B(n1005), .Z(n1006) );
  IV U1106 ( .A(n1006), .Z(n1223) );
  NOR U1107 ( .A(n94), .B(n144), .Z(n1222) );
  IV U1108 ( .A(n1222), .Z(n1007) );
  NOR U1109 ( .A(n1223), .B(n1007), .Z(n1008) );
  NOR U1110 ( .A(n1009), .B(n1008), .Z(n1011) );
  NOR U1111 ( .A(n95), .B(n144), .Z(n1012) );
  IV U1112 ( .A(n1012), .Z(n1010) );
  NOR U1113 ( .A(n1011), .B(n1010), .Z(n1016) );
  XOR U1114 ( .A(n1012), .B(n1011), .Z(n1203) );
  XOR U1115 ( .A(n1014), .B(n1013), .Z(n1204) );
  NOR U1116 ( .A(n1203), .B(n1204), .Z(n1015) );
  NOR U1117 ( .A(n1016), .B(n1015), .Z(n1199) );
  XOR U1118 ( .A(n1018), .B(n1017), .Z(n1200) );
  NOR U1119 ( .A(n1199), .B(n1200), .Z(n1019) );
  NOR U1120 ( .A(n1020), .B(n1019), .Z(n1195) );
  XOR U1121 ( .A(n1022), .B(n1021), .Z(n1196) );
  NOR U1122 ( .A(n1195), .B(n1196), .Z(n1023) );
  NOR U1123 ( .A(n1024), .B(n1023), .Z(n1191) );
  XOR U1124 ( .A(n1026), .B(n1025), .Z(n1192) );
  NOR U1125 ( .A(n1191), .B(n1192), .Z(n1027) );
  NOR U1126 ( .A(n1028), .B(n1027), .Z(n1187) );
  XOR U1127 ( .A(n1030), .B(n1029), .Z(n1188) );
  NOR U1128 ( .A(n1187), .B(n1188), .Z(n1031) );
  NOR U1129 ( .A(n1032), .B(n1031), .Z(n1183) );
  XOR U1130 ( .A(n1034), .B(n1033), .Z(n1184) );
  NOR U1131 ( .A(n1183), .B(n1184), .Z(n1035) );
  NOR U1132 ( .A(n1036), .B(n1035), .Z(n1179) );
  XOR U1133 ( .A(n1038), .B(n1037), .Z(n1180) );
  NOR U1134 ( .A(n1179), .B(n1180), .Z(n1039) );
  NOR U1135 ( .A(n1040), .B(n1039), .Z(n1175) );
  XOR U1136 ( .A(n1042), .B(n1041), .Z(n1176) );
  NOR U1137 ( .A(n1175), .B(n1176), .Z(n1043) );
  NOR U1138 ( .A(n1044), .B(n1043), .Z(n1171) );
  XOR U1139 ( .A(n1046), .B(n1045), .Z(n1172) );
  NOR U1140 ( .A(n1171), .B(n1172), .Z(n1047) );
  NOR U1141 ( .A(n1048), .B(n1047), .Z(n1167) );
  XOR U1142 ( .A(n1050), .B(n1049), .Z(n1168) );
  NOR U1143 ( .A(n1167), .B(n1168), .Z(n1051) );
  NOR U1144 ( .A(n1052), .B(n1051), .Z(n1163) );
  XOR U1145 ( .A(n1054), .B(n1053), .Z(n1164) );
  NOR U1146 ( .A(n1163), .B(n1164), .Z(n1055) );
  NOR U1147 ( .A(n1056), .B(n1055), .Z(n1159) );
  XOR U1148 ( .A(n1058), .B(n1057), .Z(n1160) );
  NOR U1149 ( .A(n1159), .B(n1160), .Z(n1059) );
  NOR U1150 ( .A(n1060), .B(n1059), .Z(n1155) );
  XOR U1151 ( .A(n1062), .B(n1061), .Z(n1156) );
  NOR U1152 ( .A(n1155), .B(n1156), .Z(n1063) );
  NOR U1153 ( .A(n1064), .B(n1063), .Z(n1154) );
  XOR U1154 ( .A(n1066), .B(n1065), .Z(n1153) );
  NOR U1155 ( .A(n1154), .B(n1153), .Z(n1067) );
  NOR U1156 ( .A(n1068), .B(n1067), .Z(n1152) );
  XOR U1157 ( .A(n1070), .B(n1069), .Z(n1151) );
  NOR U1158 ( .A(n1152), .B(n1151), .Z(n1071) );
  NOR U1159 ( .A(n1072), .B(n1071), .Z(n1296) );
  IV U1160 ( .A(n1296), .Z(n1147) );
  NOR U1161 ( .A(n88), .B(n144), .Z(n1292) );
  IV U1162 ( .A(n1073), .Z(n1074) );
  NOR U1163 ( .A(n1075), .B(n1074), .Z(n1080) );
  IV U1164 ( .A(n1076), .Z(n1077) );
  NOR U1165 ( .A(n1078), .B(n1077), .Z(n1079) );
  NOR U1166 ( .A(n1080), .B(n1079), .Z(n1303) );
  IV U1167 ( .A(n1303), .Z(n1146) );
  NOR U1168 ( .A(n106), .B(n146), .Z(n1299) );
  NOR U1169 ( .A(n105), .B(n149), .Z(n1309) );
  IV U1170 ( .A(n1081), .Z(n1082) );
  NOR U1171 ( .A(n1083), .B(n1082), .Z(n1087) );
  NOR U1172 ( .A(n1085), .B(n1084), .Z(n1086) );
  NOR U1173 ( .A(n1087), .B(n1086), .Z(n1308) );
  IV U1174 ( .A(n1088), .Z(n1089) );
  NOR U1175 ( .A(n1090), .B(n1089), .Z(n1094) );
  NOR U1176 ( .A(n1092), .B(n1091), .Z(n1093) );
  NOR U1177 ( .A(n1094), .B(n1093), .Z(n1318) );
  NOR U1178 ( .A(n104), .B(n151), .Z(n1314) );
  NOR U1179 ( .A(n89), .B(n152), .Z(n1324) );
  IV U1180 ( .A(n1095), .Z(n1096) );
  NOR U1181 ( .A(n1097), .B(n1096), .Z(n1101) );
  NOR U1182 ( .A(n1099), .B(n1098), .Z(n1100) );
  NOR U1183 ( .A(n1101), .B(n1100), .Z(n1323) );
  IV U1184 ( .A(n1102), .Z(n1103) );
  NOR U1185 ( .A(n1104), .B(n1103), .Z(n1108) );
  NOR U1186 ( .A(n1106), .B(n1105), .Z(n1107) );
  NOR U1187 ( .A(n1108), .B(n1107), .Z(n1333) );
  NOR U1188 ( .A(n103), .B(n154), .Z(n1329) );
  NOR U1189 ( .A(n1110), .B(n1109), .Z(n1114) );
  NOR U1190 ( .A(n1112), .B(n1111), .Z(n1113) );
  NOR U1191 ( .A(n1114), .B(n1113), .Z(n1347) );
  NOR U1192 ( .A(n102), .B(n159), .Z(n1345) );
  IV U1193 ( .A(n1345), .Z(n1137) );
  IV U1194 ( .A(n1115), .Z(n1116) );
  NOR U1195 ( .A(n1117), .B(n1116), .Z(n1121) );
  NOR U1196 ( .A(n1119), .B(n1118), .Z(n1120) );
  NOR U1197 ( .A(n1121), .B(n1120), .Z(n1352) );
  NOR U1198 ( .A(n101), .B(n160), .Z(n1351) );
  NOR U1199 ( .A(n1123), .B(n1122), .Z(n1127) );
  NOR U1200 ( .A(n1125), .B(n1124), .Z(n1126) );
  NOR U1201 ( .A(n1127), .B(n1126), .Z(n1362) );
  NOR U1202 ( .A(n100), .B(n162), .Z(n1359) );
  IV U1203 ( .A(n1128), .Z(n1129) );
  NOR U1204 ( .A(n1130), .B(n1129), .Z(n1134) );
  NOR U1205 ( .A(n1132), .B(n1131), .Z(n1133) );
  NOR U1206 ( .A(n1134), .B(n1133), .Z(n1367) );
  NOR U1207 ( .A(n164), .B(n99), .Z(n1365) );
  XOR U1208 ( .A(n1367), .B(n1365), .Z(n1369) );
  NOR U1209 ( .A(n166), .B(n98), .Z(n1135) );
  IV U1210 ( .A(n1135), .Z(n1368) );
  XOR U1211 ( .A(n1369), .B(n1368), .Z(n1358) );
  XOR U1212 ( .A(n1359), .B(n1358), .Z(n1360) );
  XOR U1213 ( .A(n1362), .B(n1360), .Z(n1350) );
  XOR U1214 ( .A(n1351), .B(n1350), .Z(n1136) );
  IV U1215 ( .A(n1136), .Z(n1353) );
  XOR U1216 ( .A(n1352), .B(n1353), .Z(n1344) );
  XOR U1217 ( .A(n1137), .B(n1344), .Z(n1346) );
  XOR U1218 ( .A(n1347), .B(n1346), .Z(n1341) );
  IV U1219 ( .A(n1341), .Z(n1145) );
  IV U1220 ( .A(n1138), .Z(n1139) );
  NOR U1221 ( .A(n1140), .B(n1139), .Z(n1144) );
  NOR U1222 ( .A(n1142), .B(n1141), .Z(n1143) );
  NOR U1223 ( .A(n1144), .B(n1143), .Z(n1339) );
  NOR U1224 ( .A(n90), .B(n157), .Z(n1337) );
  XOR U1225 ( .A(n1339), .B(n1337), .Z(n1340) );
  XOR U1226 ( .A(n1145), .B(n1340), .Z(n1331) );
  XOR U1227 ( .A(n1329), .B(n1331), .Z(n1332) );
  XOR U1228 ( .A(n1333), .B(n1332), .Z(n1321) );
  XOR U1229 ( .A(n1323), .B(n1321), .Z(n1326) );
  XOR U1230 ( .A(n1324), .B(n1326), .Z(n1316) );
  XOR U1231 ( .A(n1314), .B(n1316), .Z(n1317) );
  XOR U1232 ( .A(n1318), .B(n1317), .Z(n1306) );
  XOR U1233 ( .A(n1308), .B(n1306), .Z(n1311) );
  XOR U1234 ( .A(n1309), .B(n1311), .Z(n1301) );
  XOR U1235 ( .A(n1299), .B(n1301), .Z(n1302) );
  XOR U1236 ( .A(n1146), .B(n1302), .Z(n1294) );
  XOR U1237 ( .A(n1292), .B(n1294), .Z(n1295) );
  XOR U1238 ( .A(n1147), .B(n1295), .Z(n1149) );
  NOR U1239 ( .A(n107), .B(n142), .Z(n1150) );
  IV U1240 ( .A(n1150), .Z(n1148) );
  NOR U1241 ( .A(n1149), .B(n1148), .Z(n1291) );
  XOR U1242 ( .A(n1150), .B(n1149), .Z(n1526) );
  NOR U1243 ( .A(n88), .B(n142), .Z(n1285) );
  XOR U1244 ( .A(n1152), .B(n1151), .Z(n1284) );
  NOR U1245 ( .A(n1285), .B(n1284), .Z(n1288) );
  NOR U1246 ( .A(n106), .B(n142), .Z(n1280) );
  XOR U1247 ( .A(n1154), .B(n1153), .Z(n1279) );
  NOR U1248 ( .A(n1280), .B(n1279), .Z(n1283) );
  IV U1249 ( .A(n1155), .Z(n1157) );
  XOR U1250 ( .A(n1157), .B(n1156), .Z(n1274) );
  NOR U1251 ( .A(n105), .B(n142), .Z(n1275) );
  IV U1252 ( .A(n1275), .Z(n1158) );
  NOR U1253 ( .A(n1274), .B(n1158), .Z(n1277) );
  IV U1254 ( .A(n1159), .Z(n1161) );
  XOR U1255 ( .A(n1161), .B(n1160), .Z(n1270) );
  NOR U1256 ( .A(n104), .B(n142), .Z(n1271) );
  IV U1257 ( .A(n1271), .Z(n1162) );
  NOR U1258 ( .A(n1270), .B(n1162), .Z(n1273) );
  IV U1259 ( .A(n1163), .Z(n1165) );
  XOR U1260 ( .A(n1165), .B(n1164), .Z(n1266) );
  NOR U1261 ( .A(n89), .B(n142), .Z(n1267) );
  IV U1262 ( .A(n1267), .Z(n1166) );
  NOR U1263 ( .A(n1266), .B(n1166), .Z(n1269) );
  XOR U1264 ( .A(n1168), .B(n1167), .Z(n1169) );
  IV U1265 ( .A(n1169), .Z(n1262) );
  NOR U1266 ( .A(n103), .B(n142), .Z(n1263) );
  IV U1267 ( .A(n1263), .Z(n1170) );
  NOR U1268 ( .A(n1262), .B(n1170), .Z(n1265) );
  XOR U1269 ( .A(n1172), .B(n1171), .Z(n1173) );
  IV U1270 ( .A(n1173), .Z(n1258) );
  NOR U1271 ( .A(n90), .B(n142), .Z(n1259) );
  IV U1272 ( .A(n1259), .Z(n1174) );
  NOR U1273 ( .A(n1258), .B(n1174), .Z(n1261) );
  XOR U1274 ( .A(n1176), .B(n1175), .Z(n1177) );
  IV U1275 ( .A(n1177), .Z(n1254) );
  NOR U1276 ( .A(n102), .B(n142), .Z(n1255) );
  IV U1277 ( .A(n1255), .Z(n1178) );
  NOR U1278 ( .A(n1254), .B(n1178), .Z(n1257) );
  XOR U1279 ( .A(n1180), .B(n1179), .Z(n1181) );
  IV U1280 ( .A(n1181), .Z(n1250) );
  NOR U1281 ( .A(n101), .B(n142), .Z(n1251) );
  IV U1282 ( .A(n1251), .Z(n1182) );
  NOR U1283 ( .A(n1250), .B(n1182), .Z(n1253) );
  XOR U1284 ( .A(n1184), .B(n1183), .Z(n1185) );
  IV U1285 ( .A(n1185), .Z(n1246) );
  NOR U1286 ( .A(n100), .B(n142), .Z(n1247) );
  IV U1287 ( .A(n1247), .Z(n1186) );
  NOR U1288 ( .A(n1246), .B(n1186), .Z(n1249) );
  XOR U1289 ( .A(n1188), .B(n1187), .Z(n1189) );
  IV U1290 ( .A(n1189), .Z(n1242) );
  NOR U1291 ( .A(n99), .B(n142), .Z(n1243) );
  IV U1292 ( .A(n1243), .Z(n1190) );
  NOR U1293 ( .A(n1242), .B(n1190), .Z(n1245) );
  XOR U1294 ( .A(n1192), .B(n1191), .Z(n1193) );
  IV U1295 ( .A(n1193), .Z(n1238) );
  NOR U1296 ( .A(n98), .B(n142), .Z(n1239) );
  IV U1297 ( .A(n1239), .Z(n1194) );
  NOR U1298 ( .A(n1238), .B(n1194), .Z(n1241) );
  XOR U1299 ( .A(n1196), .B(n1195), .Z(n1197) );
  IV U1300 ( .A(n1197), .Z(n1234) );
  NOR U1301 ( .A(n91), .B(n142), .Z(n1235) );
  IV U1302 ( .A(n1235), .Z(n1198) );
  NOR U1303 ( .A(n1234), .B(n1198), .Z(n1237) );
  XOR U1304 ( .A(n1200), .B(n1199), .Z(n1201) );
  IV U1305 ( .A(n1201), .Z(n1230) );
  NOR U1306 ( .A(n97), .B(n142), .Z(n1231) );
  IV U1307 ( .A(n1231), .Z(n1202) );
  NOR U1308 ( .A(n1230), .B(n1202), .Z(n1233) );
  NOR U1309 ( .A(n96), .B(n142), .Z(n1227) );
  IV U1310 ( .A(n1227), .Z(n1206) );
  XOR U1311 ( .A(n1204), .B(n1203), .Z(n1205) );
  IV U1312 ( .A(n1205), .Z(n1226) );
  NOR U1313 ( .A(n1206), .B(n1226), .Z(n1229) );
  NOR U1314 ( .A(n93), .B(n142), .Z(n1707) );
  IV U1315 ( .A(n1707), .Z(n1208) );
  NOR U1316 ( .A(n144), .B(n168), .Z(n1211) );
  IV U1317 ( .A(n1211), .Z(n1207) );
  NOR U1318 ( .A(n1208), .B(n1207), .Z(n1446) );
  IV U1319 ( .A(n1446), .Z(n1209) );
  NOR U1320 ( .A(n1210), .B(n1209), .Z(n1218) );
  XOR U1321 ( .A(n1212), .B(n1211), .Z(n1213) );
  NOR U1322 ( .A(n1446), .B(n1213), .Z(n1214) );
  NOR U1323 ( .A(n1218), .B(n1214), .Z(n1215) );
  IV U1324 ( .A(n1215), .Z(n1459) );
  NOR U1325 ( .A(n94), .B(n142), .Z(n1458) );
  IV U1326 ( .A(n1458), .Z(n1216) );
  NOR U1327 ( .A(n1459), .B(n1216), .Z(n1217) );
  NOR U1328 ( .A(n1218), .B(n1217), .Z(n1220) );
  NOR U1329 ( .A(n95), .B(n142), .Z(n1221) );
  IV U1330 ( .A(n1221), .Z(n1219) );
  NOR U1331 ( .A(n1220), .B(n1219), .Z(n1225) );
  XOR U1332 ( .A(n1221), .B(n1220), .Z(n1439) );
  XOR U1333 ( .A(n1223), .B(n1222), .Z(n1440) );
  NOR U1334 ( .A(n1439), .B(n1440), .Z(n1224) );
  NOR U1335 ( .A(n1225), .B(n1224), .Z(n1435) );
  XOR U1336 ( .A(n1227), .B(n1226), .Z(n1436) );
  NOR U1337 ( .A(n1435), .B(n1436), .Z(n1228) );
  NOR U1338 ( .A(n1229), .B(n1228), .Z(n1431) );
  XOR U1339 ( .A(n1231), .B(n1230), .Z(n1432) );
  NOR U1340 ( .A(n1431), .B(n1432), .Z(n1232) );
  NOR U1341 ( .A(n1233), .B(n1232), .Z(n1427) );
  XOR U1342 ( .A(n1235), .B(n1234), .Z(n1428) );
  NOR U1343 ( .A(n1427), .B(n1428), .Z(n1236) );
  NOR U1344 ( .A(n1237), .B(n1236), .Z(n1423) );
  XOR U1345 ( .A(n1239), .B(n1238), .Z(n1424) );
  NOR U1346 ( .A(n1423), .B(n1424), .Z(n1240) );
  NOR U1347 ( .A(n1241), .B(n1240), .Z(n1419) );
  XOR U1348 ( .A(n1243), .B(n1242), .Z(n1420) );
  NOR U1349 ( .A(n1419), .B(n1420), .Z(n1244) );
  NOR U1350 ( .A(n1245), .B(n1244), .Z(n1415) );
  XOR U1351 ( .A(n1247), .B(n1246), .Z(n1416) );
  NOR U1352 ( .A(n1415), .B(n1416), .Z(n1248) );
  NOR U1353 ( .A(n1249), .B(n1248), .Z(n1411) );
  XOR U1354 ( .A(n1251), .B(n1250), .Z(n1412) );
  NOR U1355 ( .A(n1411), .B(n1412), .Z(n1252) );
  NOR U1356 ( .A(n1253), .B(n1252), .Z(n1407) );
  XOR U1357 ( .A(n1255), .B(n1254), .Z(n1408) );
  NOR U1358 ( .A(n1407), .B(n1408), .Z(n1256) );
  NOR U1359 ( .A(n1257), .B(n1256), .Z(n1403) );
  XOR U1360 ( .A(n1259), .B(n1258), .Z(n1404) );
  NOR U1361 ( .A(n1403), .B(n1404), .Z(n1260) );
  NOR U1362 ( .A(n1261), .B(n1260), .Z(n1399) );
  XOR U1363 ( .A(n1263), .B(n1262), .Z(n1400) );
  NOR U1364 ( .A(n1399), .B(n1400), .Z(n1264) );
  NOR U1365 ( .A(n1265), .B(n1264), .Z(n1395) );
  XOR U1366 ( .A(n1267), .B(n1266), .Z(n1396) );
  NOR U1367 ( .A(n1395), .B(n1396), .Z(n1268) );
  NOR U1368 ( .A(n1269), .B(n1268), .Z(n1391) );
  XOR U1369 ( .A(n1271), .B(n1270), .Z(n1392) );
  NOR U1370 ( .A(n1391), .B(n1392), .Z(n1272) );
  NOR U1371 ( .A(n1273), .B(n1272), .Z(n1387) );
  XOR U1372 ( .A(n1275), .B(n1274), .Z(n1388) );
  NOR U1373 ( .A(n1387), .B(n1388), .Z(n1276) );
  NOR U1374 ( .A(n1277), .B(n1276), .Z(n1278) );
  IV U1375 ( .A(n1278), .Z(n1385) );
  XOR U1376 ( .A(n1280), .B(n1279), .Z(n1281) );
  IV U1377 ( .A(n1281), .Z(n1384) );
  NOR U1378 ( .A(n1385), .B(n1384), .Z(n1282) );
  NOR U1379 ( .A(n1283), .B(n1282), .Z(n1382) );
  XOR U1380 ( .A(n1285), .B(n1284), .Z(n1286) );
  IV U1381 ( .A(n1286), .Z(n1381) );
  NOR U1382 ( .A(n1382), .B(n1381), .Z(n1287) );
  NOR U1383 ( .A(n1288), .B(n1287), .Z(n1527) );
  IV U1384 ( .A(n1527), .Z(n1289) );
  NOR U1385 ( .A(n1526), .B(n1289), .Z(n1290) );
  NOR U1386 ( .A(n1291), .B(n1290), .Z(n1544) );
  NOR U1387 ( .A(n87), .B(n142), .Z(n1540) );
  IV U1388 ( .A(n1292), .Z(n1293) );
  NOR U1389 ( .A(n1294), .B(n1293), .Z(n1298) );
  NOR U1390 ( .A(n1296), .B(n1295), .Z(n1297) );
  NOR U1391 ( .A(n1298), .B(n1297), .Z(n1551) );
  IV U1392 ( .A(n1551), .Z(n1380) );
  NOR U1393 ( .A(n107), .B(n144), .Z(n1547) );
  IV U1394 ( .A(n1299), .Z(n1300) );
  NOR U1395 ( .A(n1301), .B(n1300), .Z(n1305) );
  NOR U1396 ( .A(n1303), .B(n1302), .Z(n1304) );
  NOR U1397 ( .A(n1305), .B(n1304), .Z(n1558) );
  IV U1398 ( .A(n1558), .Z(n1379) );
  NOR U1399 ( .A(n88), .B(n146), .Z(n1554) );
  IV U1400 ( .A(n1306), .Z(n1307) );
  NOR U1401 ( .A(n1308), .B(n1307), .Z(n1313) );
  IV U1402 ( .A(n1309), .Z(n1310) );
  NOR U1403 ( .A(n1311), .B(n1310), .Z(n1312) );
  NOR U1404 ( .A(n1313), .B(n1312), .Z(n1565) );
  IV U1405 ( .A(n1565), .Z(n1378) );
  NOR U1406 ( .A(n106), .B(n149), .Z(n1561) );
  IV U1407 ( .A(n1314), .Z(n1315) );
  NOR U1408 ( .A(n1316), .B(n1315), .Z(n1320) );
  NOR U1409 ( .A(n1318), .B(n1317), .Z(n1319) );
  NOR U1410 ( .A(n1320), .B(n1319), .Z(n1572) );
  IV U1411 ( .A(n1572), .Z(n1377) );
  NOR U1412 ( .A(n105), .B(n151), .Z(n1568) );
  IV U1413 ( .A(n1321), .Z(n1322) );
  NOR U1414 ( .A(n1323), .B(n1322), .Z(n1328) );
  IV U1415 ( .A(n1324), .Z(n1325) );
  NOR U1416 ( .A(n1326), .B(n1325), .Z(n1327) );
  NOR U1417 ( .A(n1328), .B(n1327), .Z(n1579) );
  IV U1418 ( .A(n1579), .Z(n1376) );
  IV U1419 ( .A(n1329), .Z(n1330) );
  NOR U1420 ( .A(n1331), .B(n1330), .Z(n1335) );
  NOR U1421 ( .A(n1333), .B(n1332), .Z(n1334) );
  NOR U1422 ( .A(n1335), .B(n1334), .Z(n1336) );
  IV U1423 ( .A(n1336), .Z(n1585) );
  NOR U1424 ( .A(n89), .B(n154), .Z(n1583) );
  IV U1425 ( .A(n1337), .Z(n1338) );
  NOR U1426 ( .A(n1339), .B(n1338), .Z(n1343) );
  NOR U1427 ( .A(n1341), .B(n1340), .Z(n1342) );
  NOR U1428 ( .A(n1343), .B(n1342), .Z(n1592) );
  NOR U1429 ( .A(n1345), .B(n1344), .Z(n1349) );
  NOR U1430 ( .A(n1347), .B(n1346), .Z(n1348) );
  NOR U1431 ( .A(n1349), .B(n1348), .Z(n1598) );
  NOR U1432 ( .A(n90), .B(n159), .Z(n1596) );
  IV U1433 ( .A(n1596), .Z(n1374) );
  NOR U1434 ( .A(n1351), .B(n1350), .Z(n1356) );
  IV U1435 ( .A(n1352), .Z(n1354) );
  NOR U1436 ( .A(n1354), .B(n1353), .Z(n1355) );
  NOR U1437 ( .A(n1356), .B(n1355), .Z(n1357) );
  IV U1438 ( .A(n1357), .Z(n1603) );
  NOR U1439 ( .A(n102), .B(n160), .Z(n1601) );
  XOR U1440 ( .A(n1603), .B(n1601), .Z(n1604) );
  NOR U1441 ( .A(n1359), .B(n1358), .Z(n1364) );
  IV U1442 ( .A(n1360), .Z(n1361) );
  NOR U1443 ( .A(n1362), .B(n1361), .Z(n1363) );
  NOR U1444 ( .A(n1364), .B(n1363), .Z(n1611) );
  NOR U1445 ( .A(n101), .B(n162), .Z(n1609) );
  IV U1446 ( .A(n1609), .Z(n1373) );
  IV U1447 ( .A(n1365), .Z(n1366) );
  NOR U1448 ( .A(n1367), .B(n1366), .Z(n1371) );
  NOR U1449 ( .A(n1369), .B(n1368), .Z(n1370) );
  NOR U1450 ( .A(n1371), .B(n1370), .Z(n1616) );
  NOR U1451 ( .A(n164), .B(n100), .Z(n1614) );
  XOR U1452 ( .A(n1616), .B(n1614), .Z(n1618) );
  NOR U1453 ( .A(n166), .B(n99), .Z(n1372) );
  IV U1454 ( .A(n1372), .Z(n1617) );
  XOR U1455 ( .A(n1618), .B(n1617), .Z(n1608) );
  XOR U1456 ( .A(n1373), .B(n1608), .Z(n1610) );
  XOR U1457 ( .A(n1611), .B(n1610), .Z(n1605) );
  XOR U1458 ( .A(n1604), .B(n1605), .Z(n1595) );
  XOR U1459 ( .A(n1374), .B(n1595), .Z(n1597) );
  XOR U1460 ( .A(n1598), .B(n1597), .Z(n1590) );
  NOR U1461 ( .A(n103), .B(n157), .Z(n1588) );
  XOR U1462 ( .A(n1590), .B(n1588), .Z(n1591) );
  XOR U1463 ( .A(n1592), .B(n1591), .Z(n1582) );
  XOR U1464 ( .A(n1583), .B(n1582), .Z(n1375) );
  IV U1465 ( .A(n1375), .Z(n1584) );
  XOR U1466 ( .A(n1585), .B(n1584), .Z(n1577) );
  NOR U1467 ( .A(n104), .B(n152), .Z(n1575) );
  XOR U1468 ( .A(n1577), .B(n1575), .Z(n1578) );
  XOR U1469 ( .A(n1376), .B(n1578), .Z(n1570) );
  XOR U1470 ( .A(n1568), .B(n1570), .Z(n1571) );
  XOR U1471 ( .A(n1377), .B(n1571), .Z(n1563) );
  XOR U1472 ( .A(n1561), .B(n1563), .Z(n1564) );
  XOR U1473 ( .A(n1378), .B(n1564), .Z(n1556) );
  XOR U1474 ( .A(n1554), .B(n1556), .Z(n1557) );
  XOR U1475 ( .A(n1379), .B(n1557), .Z(n1549) );
  XOR U1476 ( .A(n1547), .B(n1549), .Z(n1550) );
  XOR U1477 ( .A(n1380), .B(n1550), .Z(n1542) );
  XOR U1478 ( .A(n1540), .B(n1542), .Z(n1543) );
  XOR U1479 ( .A(n1544), .B(n1543), .Z(n1536) );
  XOR U1480 ( .A(n1382), .B(n1381), .Z(n1523) );
  NOR U1481 ( .A(n107), .B(n140), .Z(n1522) );
  IV U1482 ( .A(n1522), .Z(n1383) );
  NOR U1483 ( .A(n1523), .B(n1383), .Z(n1525) );
  XOR U1484 ( .A(n1385), .B(n1384), .Z(n1519) );
  NOR U1485 ( .A(n88), .B(n140), .Z(n1518) );
  IV U1486 ( .A(n1518), .Z(n1386) );
  NOR U1487 ( .A(n1519), .B(n1386), .Z(n1521) );
  IV U1488 ( .A(n1387), .Z(n1389) );
  XOR U1489 ( .A(n1389), .B(n1388), .Z(n1514) );
  NOR U1490 ( .A(n106), .B(n140), .Z(n1515) );
  IV U1491 ( .A(n1515), .Z(n1390) );
  NOR U1492 ( .A(n1514), .B(n1390), .Z(n1517) );
  IV U1493 ( .A(n1391), .Z(n1393) );
  XOR U1494 ( .A(n1393), .B(n1392), .Z(n1510) );
  NOR U1495 ( .A(n105), .B(n140), .Z(n1511) );
  IV U1496 ( .A(n1511), .Z(n1394) );
  NOR U1497 ( .A(n1510), .B(n1394), .Z(n1513) );
  IV U1498 ( .A(n1395), .Z(n1397) );
  XOR U1499 ( .A(n1397), .B(n1396), .Z(n1506) );
  NOR U1500 ( .A(n104), .B(n140), .Z(n1507) );
  IV U1501 ( .A(n1507), .Z(n1398) );
  NOR U1502 ( .A(n1506), .B(n1398), .Z(n1509) );
  XOR U1503 ( .A(n1400), .B(n1399), .Z(n1401) );
  IV U1504 ( .A(n1401), .Z(n1502) );
  NOR U1505 ( .A(n89), .B(n140), .Z(n1503) );
  IV U1506 ( .A(n1503), .Z(n1402) );
  NOR U1507 ( .A(n1502), .B(n1402), .Z(n1505) );
  XOR U1508 ( .A(n1404), .B(n1403), .Z(n1405) );
  IV U1509 ( .A(n1405), .Z(n1498) );
  NOR U1510 ( .A(n103), .B(n140), .Z(n1499) );
  IV U1511 ( .A(n1499), .Z(n1406) );
  NOR U1512 ( .A(n1498), .B(n1406), .Z(n1501) );
  XOR U1513 ( .A(n1408), .B(n1407), .Z(n1409) );
  IV U1514 ( .A(n1409), .Z(n1494) );
  NOR U1515 ( .A(n90), .B(n140), .Z(n1495) );
  IV U1516 ( .A(n1495), .Z(n1410) );
  NOR U1517 ( .A(n1494), .B(n1410), .Z(n1497) );
  XOR U1518 ( .A(n1412), .B(n1411), .Z(n1413) );
  IV U1519 ( .A(n1413), .Z(n1490) );
  NOR U1520 ( .A(n102), .B(n140), .Z(n1491) );
  IV U1521 ( .A(n1491), .Z(n1414) );
  NOR U1522 ( .A(n1490), .B(n1414), .Z(n1493) );
  XOR U1523 ( .A(n1416), .B(n1415), .Z(n1417) );
  IV U1524 ( .A(n1417), .Z(n1486) );
  NOR U1525 ( .A(n101), .B(n140), .Z(n1487) );
  IV U1526 ( .A(n1487), .Z(n1418) );
  NOR U1527 ( .A(n1486), .B(n1418), .Z(n1489) );
  XOR U1528 ( .A(n1420), .B(n1419), .Z(n1421) );
  IV U1529 ( .A(n1421), .Z(n1482) );
  NOR U1530 ( .A(n100), .B(n140), .Z(n1483) );
  IV U1531 ( .A(n1483), .Z(n1422) );
  NOR U1532 ( .A(n1482), .B(n1422), .Z(n1485) );
  NOR U1533 ( .A(n99), .B(n140), .Z(n1479) );
  IV U1534 ( .A(n1479), .Z(n1426) );
  XOR U1535 ( .A(n1424), .B(n1423), .Z(n1425) );
  IV U1536 ( .A(n1425), .Z(n1478) );
  NOR U1537 ( .A(n1426), .B(n1478), .Z(n1481) );
  XOR U1538 ( .A(n1428), .B(n1427), .Z(n1429) );
  IV U1539 ( .A(n1429), .Z(n1474) );
  NOR U1540 ( .A(n98), .B(n140), .Z(n1475) );
  IV U1541 ( .A(n1475), .Z(n1430) );
  NOR U1542 ( .A(n1474), .B(n1430), .Z(n1477) );
  XOR U1543 ( .A(n1432), .B(n1431), .Z(n1433) );
  IV U1544 ( .A(n1433), .Z(n1470) );
  NOR U1545 ( .A(n91), .B(n140), .Z(n1471) );
  IV U1546 ( .A(n1471), .Z(n1434) );
  NOR U1547 ( .A(n1470), .B(n1434), .Z(n1473) );
  XOR U1548 ( .A(n1436), .B(n1435), .Z(n1437) );
  IV U1549 ( .A(n1437), .Z(n1466) );
  NOR U1550 ( .A(n97), .B(n140), .Z(n1467) );
  IV U1551 ( .A(n1467), .Z(n1438) );
  NOR U1552 ( .A(n1466), .B(n1438), .Z(n1469) );
  NOR U1553 ( .A(n96), .B(n140), .Z(n1463) );
  IV U1554 ( .A(n1463), .Z(n1442) );
  XOR U1555 ( .A(n1440), .B(n1439), .Z(n1441) );
  IV U1556 ( .A(n1441), .Z(n1462) );
  NOR U1557 ( .A(n1442), .B(n1462), .Z(n1465) );
  NOR U1558 ( .A(n93), .B(n140), .Z(n1983) );
  IV U1559 ( .A(n1983), .Z(n1444) );
  NOR U1560 ( .A(n142), .B(n168), .Z(n1447) );
  IV U1561 ( .A(n1447), .Z(n1443) );
  NOR U1562 ( .A(n1444), .B(n1443), .Z(n1705) );
  IV U1563 ( .A(n1705), .Z(n1445) );
  NOR U1564 ( .A(n1446), .B(n1445), .Z(n1454) );
  XOR U1565 ( .A(n1448), .B(n1447), .Z(n1449) );
  NOR U1566 ( .A(n1705), .B(n1449), .Z(n1450) );
  NOR U1567 ( .A(n1454), .B(n1450), .Z(n1451) );
  IV U1568 ( .A(n1451), .Z(n1718) );
  NOR U1569 ( .A(n94), .B(n140), .Z(n1717) );
  IV U1570 ( .A(n1717), .Z(n1452) );
  NOR U1571 ( .A(n1718), .B(n1452), .Z(n1453) );
  NOR U1572 ( .A(n1454), .B(n1453), .Z(n1456) );
  NOR U1573 ( .A(n95), .B(n140), .Z(n1457) );
  IV U1574 ( .A(n1457), .Z(n1455) );
  NOR U1575 ( .A(n1456), .B(n1455), .Z(n1461) );
  XOR U1576 ( .A(n1457), .B(n1456), .Z(n1698) );
  XOR U1577 ( .A(n1459), .B(n1458), .Z(n1699) );
  NOR U1578 ( .A(n1698), .B(n1699), .Z(n1460) );
  NOR U1579 ( .A(n1461), .B(n1460), .Z(n1694) );
  XOR U1580 ( .A(n1463), .B(n1462), .Z(n1695) );
  NOR U1581 ( .A(n1694), .B(n1695), .Z(n1464) );
  NOR U1582 ( .A(n1465), .B(n1464), .Z(n1690) );
  XOR U1583 ( .A(n1467), .B(n1466), .Z(n1691) );
  NOR U1584 ( .A(n1690), .B(n1691), .Z(n1468) );
  NOR U1585 ( .A(n1469), .B(n1468), .Z(n1686) );
  XOR U1586 ( .A(n1471), .B(n1470), .Z(n1687) );
  NOR U1587 ( .A(n1686), .B(n1687), .Z(n1472) );
  NOR U1588 ( .A(n1473), .B(n1472), .Z(n1682) );
  XOR U1589 ( .A(n1475), .B(n1474), .Z(n1683) );
  NOR U1590 ( .A(n1682), .B(n1683), .Z(n1476) );
  NOR U1591 ( .A(n1477), .B(n1476), .Z(n1678) );
  XOR U1592 ( .A(n1479), .B(n1478), .Z(n1679) );
  NOR U1593 ( .A(n1678), .B(n1679), .Z(n1480) );
  NOR U1594 ( .A(n1481), .B(n1480), .Z(n1674) );
  XOR U1595 ( .A(n1483), .B(n1482), .Z(n1675) );
  NOR U1596 ( .A(n1674), .B(n1675), .Z(n1484) );
  NOR U1597 ( .A(n1485), .B(n1484), .Z(n1670) );
  XOR U1598 ( .A(n1487), .B(n1486), .Z(n1671) );
  NOR U1599 ( .A(n1670), .B(n1671), .Z(n1488) );
  NOR U1600 ( .A(n1489), .B(n1488), .Z(n1666) );
  XOR U1601 ( .A(n1491), .B(n1490), .Z(n1667) );
  NOR U1602 ( .A(n1666), .B(n1667), .Z(n1492) );
  NOR U1603 ( .A(n1493), .B(n1492), .Z(n1662) );
  XOR U1604 ( .A(n1495), .B(n1494), .Z(n1663) );
  NOR U1605 ( .A(n1662), .B(n1663), .Z(n1496) );
  NOR U1606 ( .A(n1497), .B(n1496), .Z(n1658) );
  XOR U1607 ( .A(n1499), .B(n1498), .Z(n1659) );
  NOR U1608 ( .A(n1658), .B(n1659), .Z(n1500) );
  NOR U1609 ( .A(n1501), .B(n1500), .Z(n1654) );
  XOR U1610 ( .A(n1503), .B(n1502), .Z(n1655) );
  NOR U1611 ( .A(n1654), .B(n1655), .Z(n1504) );
  NOR U1612 ( .A(n1505), .B(n1504), .Z(n1650) );
  XOR U1613 ( .A(n1507), .B(n1506), .Z(n1651) );
  NOR U1614 ( .A(n1650), .B(n1651), .Z(n1508) );
  NOR U1615 ( .A(n1509), .B(n1508), .Z(n1646) );
  XOR U1616 ( .A(n1511), .B(n1510), .Z(n1647) );
  NOR U1617 ( .A(n1646), .B(n1647), .Z(n1512) );
  NOR U1618 ( .A(n1513), .B(n1512), .Z(n1642) );
  XOR U1619 ( .A(n1515), .B(n1514), .Z(n1643) );
  NOR U1620 ( .A(n1642), .B(n1643), .Z(n1516) );
  NOR U1621 ( .A(n1517), .B(n1516), .Z(n1641) );
  XOR U1622 ( .A(n1519), .B(n1518), .Z(n1640) );
  NOR U1623 ( .A(n1641), .B(n1640), .Z(n1520) );
  NOR U1624 ( .A(n1521), .B(n1520), .Z(n1639) );
  XOR U1625 ( .A(n1523), .B(n1522), .Z(n1638) );
  NOR U1626 ( .A(n1639), .B(n1638), .Z(n1524) );
  NOR U1627 ( .A(n1525), .B(n1524), .Z(n1528) );
  XOR U1628 ( .A(n1527), .B(n1526), .Z(n1529) );
  NOR U1629 ( .A(n1528), .B(n1529), .Z(n1533) );
  IV U1630 ( .A(n1528), .Z(n1530) );
  XOR U1631 ( .A(n1530), .B(n1529), .Z(n1637) );
  NOR U1632 ( .A(n87), .B(n140), .Z(n1531) );
  IV U1633 ( .A(n1531), .Z(n1636) );
  NOR U1634 ( .A(n1637), .B(n1636), .Z(n1532) );
  NOR U1635 ( .A(n1533), .B(n1532), .Z(n1535) );
  IV U1636 ( .A(n1535), .Z(n1534) );
  NOR U1637 ( .A(n1536), .B(n1534), .Z(n1538) );
  NOR U1638 ( .A(n108), .B(n140), .Z(n1632) );
  XOR U1639 ( .A(n1536), .B(n1535), .Z(n1631) );
  NOR U1640 ( .A(n1632), .B(n1631), .Z(n1537) );
  NOR U1641 ( .A(n1538), .B(n1537), .Z(n1539) );
  IV U1642 ( .A(n1539), .Z(n1895) );
  NOR U1643 ( .A(n109), .B(n140), .Z(n1893) );
  XOR U1644 ( .A(n1895), .B(n1893), .Z(n1898) );
  IV U1645 ( .A(n1540), .Z(n1541) );
  NOR U1646 ( .A(n1542), .B(n1541), .Z(n1546) );
  NOR U1647 ( .A(n1544), .B(n1543), .Z(n1545) );
  NOR U1648 ( .A(n1546), .B(n1545), .Z(n1808) );
  NOR U1649 ( .A(n108), .B(n142), .Z(n1804) );
  IV U1650 ( .A(n1547), .Z(n1548) );
  NOR U1651 ( .A(n1549), .B(n1548), .Z(n1553) );
  NOR U1652 ( .A(n1551), .B(n1550), .Z(n1552) );
  NOR U1653 ( .A(n1553), .B(n1552), .Z(n1815) );
  IV U1654 ( .A(n1815), .Z(n1629) );
  NOR U1655 ( .A(n87), .B(n144), .Z(n1811) );
  IV U1656 ( .A(n1554), .Z(n1555) );
  NOR U1657 ( .A(n1556), .B(n1555), .Z(n1560) );
  NOR U1658 ( .A(n1558), .B(n1557), .Z(n1559) );
  NOR U1659 ( .A(n1560), .B(n1559), .Z(n1822) );
  IV U1660 ( .A(n1822), .Z(n1628) );
  NOR U1661 ( .A(n88), .B(n149), .Z(n1827) );
  IV U1662 ( .A(n1561), .Z(n1562) );
  NOR U1663 ( .A(n1563), .B(n1562), .Z(n1567) );
  NOR U1664 ( .A(n1565), .B(n1564), .Z(n1566) );
  NOR U1665 ( .A(n1567), .B(n1566), .Z(n1825) );
  XOR U1666 ( .A(n1827), .B(n1825), .Z(n1829) );
  IV U1667 ( .A(n1568), .Z(n1569) );
  NOR U1668 ( .A(n1570), .B(n1569), .Z(n1574) );
  NOR U1669 ( .A(n1572), .B(n1571), .Z(n1573) );
  NOR U1670 ( .A(n1574), .B(n1573), .Z(n1835) );
  NOR U1671 ( .A(n106), .B(n151), .Z(n1834) );
  IV U1672 ( .A(n1834), .Z(n1627) );
  IV U1673 ( .A(n1575), .Z(n1576) );
  NOR U1674 ( .A(n1577), .B(n1576), .Z(n1581) );
  NOR U1675 ( .A(n1579), .B(n1578), .Z(n1580) );
  NOR U1676 ( .A(n1581), .B(n1580), .Z(n1885) );
  IV U1677 ( .A(n1885), .Z(n1625) );
  NOR U1678 ( .A(n1583), .B(n1582), .Z(n1587) );
  NOR U1679 ( .A(n1585), .B(n1584), .Z(n1586) );
  NOR U1680 ( .A(n1587), .B(n1586), .Z(n1843) );
  NOR U1681 ( .A(n104), .B(n154), .Z(n1841) );
  IV U1682 ( .A(n1841), .Z(n1624) );
  IV U1683 ( .A(n1588), .Z(n1589) );
  NOR U1684 ( .A(n1590), .B(n1589), .Z(n1594) );
  NOR U1685 ( .A(n1592), .B(n1591), .Z(n1593) );
  NOR U1686 ( .A(n1594), .B(n1593), .Z(n1846) );
  IV U1687 ( .A(n1846), .Z(n1622) );
  NOR U1688 ( .A(n1596), .B(n1595), .Z(n1600) );
  NOR U1689 ( .A(n1598), .B(n1597), .Z(n1599) );
  NOR U1690 ( .A(n1600), .B(n1599), .Z(n1856) );
  NOR U1691 ( .A(n103), .B(n159), .Z(n1854) );
  NOR U1692 ( .A(n90), .B(n160), .Z(n1863) );
  IV U1693 ( .A(n1601), .Z(n1602) );
  NOR U1694 ( .A(n1603), .B(n1602), .Z(n1607) );
  NOR U1695 ( .A(n1605), .B(n1604), .Z(n1606) );
  NOR U1696 ( .A(n1607), .B(n1606), .Z(n1859) );
  NOR U1697 ( .A(n1609), .B(n1608), .Z(n1613) );
  NOR U1698 ( .A(n1611), .B(n1610), .Z(n1612) );
  NOR U1699 ( .A(n1613), .B(n1612), .Z(n1871) );
  NOR U1700 ( .A(n102), .B(n162), .Z(n1868) );
  IV U1701 ( .A(n1614), .Z(n1615) );
  NOR U1702 ( .A(n1616), .B(n1615), .Z(n1620) );
  NOR U1703 ( .A(n1618), .B(n1617), .Z(n1619) );
  NOR U1704 ( .A(n1620), .B(n1619), .Z(n1876) );
  NOR U1705 ( .A(n164), .B(n101), .Z(n1874) );
  XOR U1706 ( .A(n1876), .B(n1874), .Z(n1878) );
  NOR U1707 ( .A(n166), .B(n100), .Z(n1621) );
  IV U1708 ( .A(n1621), .Z(n1877) );
  XOR U1709 ( .A(n1878), .B(n1877), .Z(n1867) );
  XOR U1710 ( .A(n1868), .B(n1867), .Z(n1869) );
  XOR U1711 ( .A(n1871), .B(n1869), .Z(n1860) );
  XOR U1712 ( .A(n1859), .B(n1860), .Z(n1862) );
  XOR U1713 ( .A(n1863), .B(n1862), .Z(n1852) );
  XOR U1714 ( .A(n1854), .B(n1852), .Z(n1855) );
  XOR U1715 ( .A(n1856), .B(n1855), .Z(n1847) );
  XOR U1716 ( .A(n1622), .B(n1847), .Z(n1849) );
  NOR U1717 ( .A(n89), .B(n157), .Z(n1623) );
  IV U1718 ( .A(n1623), .Z(n1848) );
  XOR U1719 ( .A(n1849), .B(n1848), .Z(n1840) );
  XOR U1720 ( .A(n1624), .B(n1840), .Z(n1842) );
  XOR U1721 ( .A(n1843), .B(n1842), .Z(n1886) );
  XOR U1722 ( .A(n1625), .B(n1886), .Z(n1888) );
  NOR U1723 ( .A(n105), .B(n152), .Z(n1626) );
  IV U1724 ( .A(n1626), .Z(n1887) );
  XOR U1725 ( .A(n1888), .B(n1887), .Z(n1833) );
  XOR U1726 ( .A(n1627), .B(n1833), .Z(n1836) );
  XOR U1727 ( .A(n1835), .B(n1836), .Z(n1828) );
  XOR U1728 ( .A(n1829), .B(n1828), .Z(n1820) );
  NOR U1729 ( .A(n107), .B(n146), .Z(n1818) );
  XOR U1730 ( .A(n1820), .B(n1818), .Z(n1821) );
  XOR U1731 ( .A(n1628), .B(n1821), .Z(n1813) );
  XOR U1732 ( .A(n1811), .B(n1813), .Z(n1814) );
  XOR U1733 ( .A(n1629), .B(n1814), .Z(n1806) );
  XOR U1734 ( .A(n1804), .B(n1806), .Z(n1807) );
  XOR U1735 ( .A(n1808), .B(n1807), .Z(n1896) );
  XOR U1736 ( .A(n1898), .B(n1896), .Z(n1800) );
  NOR U1737 ( .A(n110), .B(n138), .Z(n1801) );
  IV U1738 ( .A(n1801), .Z(n1630) );
  NOR U1739 ( .A(n1800), .B(n1630), .Z(n1803) );
  XOR U1740 ( .A(n1632), .B(n1631), .Z(n1635) );
  NOR U1741 ( .A(n109), .B(n138), .Z(n1634) );
  IV U1742 ( .A(n1634), .Z(n1633) );
  NOR U1743 ( .A(n1635), .B(n1633), .Z(n1799) );
  XOR U1744 ( .A(n1635), .B(n1634), .Z(n2073) );
  NOR U1745 ( .A(n108), .B(n138), .Z(n1792) );
  XOR U1746 ( .A(n1637), .B(n1636), .Z(n1793) );
  NOR U1747 ( .A(n1792), .B(n1793), .Z(n1796) );
  NOR U1748 ( .A(n87), .B(n138), .Z(n1788) );
  XOR U1749 ( .A(n1639), .B(n1638), .Z(n1787) );
  NOR U1750 ( .A(n1788), .B(n1787), .Z(n1791) );
  NOR U1751 ( .A(n107), .B(n138), .Z(n1783) );
  XOR U1752 ( .A(n1641), .B(n1640), .Z(n1782) );
  NOR U1753 ( .A(n1783), .B(n1782), .Z(n1786) );
  IV U1754 ( .A(n1642), .Z(n1644) );
  XOR U1755 ( .A(n1644), .B(n1643), .Z(n1777) );
  NOR U1756 ( .A(n88), .B(n138), .Z(n1778) );
  IV U1757 ( .A(n1778), .Z(n1645) );
  NOR U1758 ( .A(n1777), .B(n1645), .Z(n1780) );
  IV U1759 ( .A(n1646), .Z(n1648) );
  XOR U1760 ( .A(n1648), .B(n1647), .Z(n1773) );
  NOR U1761 ( .A(n106), .B(n138), .Z(n1774) );
  IV U1762 ( .A(n1774), .Z(n1649) );
  NOR U1763 ( .A(n1773), .B(n1649), .Z(n1776) );
  IV U1764 ( .A(n1650), .Z(n1652) );
  XOR U1765 ( .A(n1652), .B(n1651), .Z(n1769) );
  NOR U1766 ( .A(n105), .B(n138), .Z(n1770) );
  IV U1767 ( .A(n1770), .Z(n1653) );
  NOR U1768 ( .A(n1769), .B(n1653), .Z(n1772) );
  XOR U1769 ( .A(n1655), .B(n1654), .Z(n1656) );
  IV U1770 ( .A(n1656), .Z(n1765) );
  NOR U1771 ( .A(n104), .B(n138), .Z(n1766) );
  IV U1772 ( .A(n1766), .Z(n1657) );
  NOR U1773 ( .A(n1765), .B(n1657), .Z(n1768) );
  XOR U1774 ( .A(n1659), .B(n1658), .Z(n1660) );
  IV U1775 ( .A(n1660), .Z(n1761) );
  NOR U1776 ( .A(n89), .B(n138), .Z(n1762) );
  IV U1777 ( .A(n1762), .Z(n1661) );
  NOR U1778 ( .A(n1761), .B(n1661), .Z(n1764) );
  XOR U1779 ( .A(n1663), .B(n1662), .Z(n1664) );
  IV U1780 ( .A(n1664), .Z(n1757) );
  NOR U1781 ( .A(n103), .B(n138), .Z(n1758) );
  IV U1782 ( .A(n1758), .Z(n1665) );
  NOR U1783 ( .A(n1757), .B(n1665), .Z(n1760) );
  XOR U1784 ( .A(n1667), .B(n1666), .Z(n1668) );
  IV U1785 ( .A(n1668), .Z(n1753) );
  NOR U1786 ( .A(n90), .B(n138), .Z(n1754) );
  IV U1787 ( .A(n1754), .Z(n1669) );
  NOR U1788 ( .A(n1753), .B(n1669), .Z(n1756) );
  IV U1789 ( .A(n1670), .Z(n1672) );
  XOR U1790 ( .A(n1672), .B(n1671), .Z(n1749) );
  NOR U1791 ( .A(n102), .B(n138), .Z(n1750) );
  IV U1792 ( .A(n1750), .Z(n1673) );
  NOR U1793 ( .A(n1749), .B(n1673), .Z(n1752) );
  XOR U1794 ( .A(n1675), .B(n1674), .Z(n1676) );
  IV U1795 ( .A(n1676), .Z(n1745) );
  NOR U1796 ( .A(n101), .B(n138), .Z(n1746) );
  IV U1797 ( .A(n1746), .Z(n1677) );
  NOR U1798 ( .A(n1745), .B(n1677), .Z(n1748) );
  XOR U1799 ( .A(n1679), .B(n1678), .Z(n1680) );
  IV U1800 ( .A(n1680), .Z(n1741) );
  NOR U1801 ( .A(n100), .B(n138), .Z(n1742) );
  IV U1802 ( .A(n1742), .Z(n1681) );
  NOR U1803 ( .A(n1741), .B(n1681), .Z(n1744) );
  XOR U1804 ( .A(n1683), .B(n1682), .Z(n1684) );
  IV U1805 ( .A(n1684), .Z(n1737) );
  NOR U1806 ( .A(n99), .B(n138), .Z(n1738) );
  IV U1807 ( .A(n1738), .Z(n1685) );
  NOR U1808 ( .A(n1737), .B(n1685), .Z(n1740) );
  XOR U1809 ( .A(n1687), .B(n1686), .Z(n1688) );
  IV U1810 ( .A(n1688), .Z(n1733) );
  NOR U1811 ( .A(n98), .B(n138), .Z(n1734) );
  IV U1812 ( .A(n1734), .Z(n1689) );
  NOR U1813 ( .A(n1733), .B(n1689), .Z(n1736) );
  XOR U1814 ( .A(n1691), .B(n1690), .Z(n1692) );
  IV U1815 ( .A(n1692), .Z(n1729) );
  NOR U1816 ( .A(n91), .B(n138), .Z(n1730) );
  IV U1817 ( .A(n1730), .Z(n1693) );
  NOR U1818 ( .A(n1729), .B(n1693), .Z(n1732) );
  XOR U1819 ( .A(n1695), .B(n1694), .Z(n1696) );
  IV U1820 ( .A(n1696), .Z(n1725) );
  NOR U1821 ( .A(n97), .B(n138), .Z(n1726) );
  IV U1822 ( .A(n1726), .Z(n1697) );
  NOR U1823 ( .A(n1725), .B(n1697), .Z(n1728) );
  XOR U1824 ( .A(n1699), .B(n1698), .Z(n1700) );
  IV U1825 ( .A(n1700), .Z(n1721) );
  NOR U1826 ( .A(n96), .B(n138), .Z(n1722) );
  IV U1827 ( .A(n1722), .Z(n1701) );
  NOR U1828 ( .A(n1721), .B(n1701), .Z(n1724) );
  NOR U1829 ( .A(n93), .B(n138), .Z(n3056) );
  IV U1830 ( .A(n3056), .Z(n1703) );
  NOR U1831 ( .A(n140), .B(n168), .Z(n1706) );
  IV U1832 ( .A(n1706), .Z(n1702) );
  NOR U1833 ( .A(n1703), .B(n1702), .Z(n1981) );
  IV U1834 ( .A(n1981), .Z(n1704) );
  NOR U1835 ( .A(n1705), .B(n1704), .Z(n1713) );
  XOR U1836 ( .A(n1707), .B(n1706), .Z(n1708) );
  NOR U1837 ( .A(n1981), .B(n1708), .Z(n1709) );
  NOR U1838 ( .A(n1713), .B(n1709), .Z(n1710) );
  IV U1839 ( .A(n1710), .Z(n1994) );
  NOR U1840 ( .A(n94), .B(n138), .Z(n1993) );
  IV U1841 ( .A(n1993), .Z(n1711) );
  NOR U1842 ( .A(n1994), .B(n1711), .Z(n1712) );
  NOR U1843 ( .A(n1713), .B(n1712), .Z(n1715) );
  NOR U1844 ( .A(n95), .B(n138), .Z(n1716) );
  IV U1845 ( .A(n1716), .Z(n1714) );
  NOR U1846 ( .A(n1715), .B(n1714), .Z(n1720) );
  XOR U1847 ( .A(n1716), .B(n1715), .Z(n1974) );
  XOR U1848 ( .A(n1718), .B(n1717), .Z(n1975) );
  NOR U1849 ( .A(n1974), .B(n1975), .Z(n1719) );
  NOR U1850 ( .A(n1720), .B(n1719), .Z(n1970) );
  XOR U1851 ( .A(n1722), .B(n1721), .Z(n1971) );
  NOR U1852 ( .A(n1970), .B(n1971), .Z(n1723) );
  NOR U1853 ( .A(n1724), .B(n1723), .Z(n1966) );
  XOR U1854 ( .A(n1726), .B(n1725), .Z(n1967) );
  NOR U1855 ( .A(n1966), .B(n1967), .Z(n1727) );
  NOR U1856 ( .A(n1728), .B(n1727), .Z(n1962) );
  XOR U1857 ( .A(n1730), .B(n1729), .Z(n1963) );
  NOR U1858 ( .A(n1962), .B(n1963), .Z(n1731) );
  NOR U1859 ( .A(n1732), .B(n1731), .Z(n1958) );
  XOR U1860 ( .A(n1734), .B(n1733), .Z(n1959) );
  NOR U1861 ( .A(n1958), .B(n1959), .Z(n1735) );
  NOR U1862 ( .A(n1736), .B(n1735), .Z(n1954) );
  XOR U1863 ( .A(n1738), .B(n1737), .Z(n1955) );
  NOR U1864 ( .A(n1954), .B(n1955), .Z(n1739) );
  NOR U1865 ( .A(n1740), .B(n1739), .Z(n1950) );
  XOR U1866 ( .A(n1742), .B(n1741), .Z(n1951) );
  NOR U1867 ( .A(n1950), .B(n1951), .Z(n1743) );
  NOR U1868 ( .A(n1744), .B(n1743), .Z(n1946) );
  XOR U1869 ( .A(n1746), .B(n1745), .Z(n1947) );
  NOR U1870 ( .A(n1946), .B(n1947), .Z(n1747) );
  NOR U1871 ( .A(n1748), .B(n1747), .Z(n1942) );
  XOR U1872 ( .A(n1750), .B(n1749), .Z(n1943) );
  NOR U1873 ( .A(n1942), .B(n1943), .Z(n1751) );
  NOR U1874 ( .A(n1752), .B(n1751), .Z(n1938) );
  XOR U1875 ( .A(n1754), .B(n1753), .Z(n1939) );
  NOR U1876 ( .A(n1938), .B(n1939), .Z(n1755) );
  NOR U1877 ( .A(n1756), .B(n1755), .Z(n1934) );
  XOR U1878 ( .A(n1758), .B(n1757), .Z(n1935) );
  NOR U1879 ( .A(n1934), .B(n1935), .Z(n1759) );
  NOR U1880 ( .A(n1760), .B(n1759), .Z(n1930) );
  XOR U1881 ( .A(n1762), .B(n1761), .Z(n1931) );
  NOR U1882 ( .A(n1930), .B(n1931), .Z(n1763) );
  NOR U1883 ( .A(n1764), .B(n1763), .Z(n1926) );
  XOR U1884 ( .A(n1766), .B(n1765), .Z(n1927) );
  NOR U1885 ( .A(n1926), .B(n1927), .Z(n1767) );
  NOR U1886 ( .A(n1768), .B(n1767), .Z(n1922) );
  XOR U1887 ( .A(n1770), .B(n1769), .Z(n1923) );
  NOR U1888 ( .A(n1922), .B(n1923), .Z(n1771) );
  NOR U1889 ( .A(n1772), .B(n1771), .Z(n1918) );
  XOR U1890 ( .A(n1774), .B(n1773), .Z(n1919) );
  NOR U1891 ( .A(n1918), .B(n1919), .Z(n1775) );
  NOR U1892 ( .A(n1776), .B(n1775), .Z(n1914) );
  XOR U1893 ( .A(n1778), .B(n1777), .Z(n1915) );
  NOR U1894 ( .A(n1914), .B(n1915), .Z(n1779) );
  NOR U1895 ( .A(n1780), .B(n1779), .Z(n1781) );
  IV U1896 ( .A(n1781), .Z(n1912) );
  XOR U1897 ( .A(n1783), .B(n1782), .Z(n1784) );
  IV U1898 ( .A(n1784), .Z(n1911) );
  NOR U1899 ( .A(n1912), .B(n1911), .Z(n1785) );
  NOR U1900 ( .A(n1786), .B(n1785), .Z(n1909) );
  XOR U1901 ( .A(n1788), .B(n1787), .Z(n1789) );
  IV U1902 ( .A(n1789), .Z(n1908) );
  NOR U1903 ( .A(n1909), .B(n1908), .Z(n1790) );
  NOR U1904 ( .A(n1791), .B(n1790), .Z(n1906) );
  IV U1905 ( .A(n1792), .Z(n1794) );
  XOR U1906 ( .A(n1794), .B(n1793), .Z(n1905) );
  NOR U1907 ( .A(n1906), .B(n1905), .Z(n1795) );
  NOR U1908 ( .A(n1796), .B(n1795), .Z(n2074) );
  IV U1909 ( .A(n2074), .Z(n1797) );
  NOR U1910 ( .A(n2073), .B(n1797), .Z(n1798) );
  NOR U1911 ( .A(n1799), .B(n1798), .Z(n1904) );
  XOR U1912 ( .A(n1801), .B(n1800), .Z(n1903) );
  NOR U1913 ( .A(n1904), .B(n1903), .Z(n1802) );
  NOR U1914 ( .A(n1803), .B(n1802), .Z(n2095) );
  IV U1915 ( .A(n2095), .Z(n1901) );
  NOR U1916 ( .A(n86), .B(n138), .Z(n2091) );
  IV U1917 ( .A(n1804), .Z(n1805) );
  NOR U1918 ( .A(n1806), .B(n1805), .Z(n1810) );
  NOR U1919 ( .A(n1808), .B(n1807), .Z(n1809) );
  NOR U1920 ( .A(n1810), .B(n1809), .Z(n2110) );
  NOR U1921 ( .A(n108), .B(n144), .Z(n2190) );
  IV U1922 ( .A(n1811), .Z(n1812) );
  NOR U1923 ( .A(n1813), .B(n1812), .Z(n1817) );
  NOR U1924 ( .A(n1815), .B(n1814), .Z(n1816) );
  NOR U1925 ( .A(n1817), .B(n1816), .Z(n2186) );
  IV U1926 ( .A(n1818), .Z(n1819) );
  NOR U1927 ( .A(n1820), .B(n1819), .Z(n1824) );
  NOR U1928 ( .A(n1822), .B(n1821), .Z(n1823) );
  NOR U1929 ( .A(n1824), .B(n1823), .Z(n2116) );
  NOR U1930 ( .A(n87), .B(n146), .Z(n2115) );
  IV U1931 ( .A(n2115), .Z(n1892) );
  IV U1932 ( .A(n1825), .Z(n1826) );
  NOR U1933 ( .A(n1827), .B(n1826), .Z(n1831) );
  NOR U1934 ( .A(n1829), .B(n1828), .Z(n1830) );
  NOR U1935 ( .A(n1831), .B(n1830), .Z(n1832) );
  IV U1936 ( .A(n1832), .Z(n2182) );
  NOR U1937 ( .A(n1834), .B(n1833), .Z(n1839) );
  IV U1938 ( .A(n1835), .Z(n1837) );
  NOR U1939 ( .A(n1837), .B(n1836), .Z(n1838) );
  NOR U1940 ( .A(n1839), .B(n1838), .Z(n2124) );
  NOR U1941 ( .A(n88), .B(n151), .Z(n2122) );
  NOR U1942 ( .A(n1841), .B(n1840), .Z(n1845) );
  NOR U1943 ( .A(n1843), .B(n1842), .Z(n1844) );
  NOR U1944 ( .A(n1845), .B(n1844), .Z(n2137) );
  NOR U1945 ( .A(n105), .B(n154), .Z(n2135) );
  NOR U1946 ( .A(n1847), .B(n1846), .Z(n1851) );
  NOR U1947 ( .A(n1849), .B(n1848), .Z(n1850) );
  NOR U1948 ( .A(n1851), .B(n1850), .Z(n2173) );
  IV U1949 ( .A(n1852), .Z(n1853) );
  NOR U1950 ( .A(n1854), .B(n1853), .Z(n1858) );
  NOR U1951 ( .A(n1856), .B(n1855), .Z(n1857) );
  NOR U1952 ( .A(n1858), .B(n1857), .Z(n2143) );
  NOR U1953 ( .A(n89), .B(n159), .Z(n2141) );
  IV U1954 ( .A(n2141), .Z(n1883) );
  IV U1955 ( .A(n1859), .Z(n1861) );
  NOR U1956 ( .A(n1861), .B(n1860), .Z(n1865) );
  NOR U1957 ( .A(n1863), .B(n1862), .Z(n1864) );
  NOR U1958 ( .A(n1865), .B(n1864), .Z(n1866) );
  IV U1959 ( .A(n1866), .Z(n2148) );
  NOR U1960 ( .A(n103), .B(n160), .Z(n2146) );
  XOR U1961 ( .A(n2148), .B(n2146), .Z(n2149) );
  NOR U1962 ( .A(n1868), .B(n1867), .Z(n1873) );
  IV U1963 ( .A(n1869), .Z(n1870) );
  NOR U1964 ( .A(n1871), .B(n1870), .Z(n1872) );
  NOR U1965 ( .A(n1873), .B(n1872), .Z(n2156) );
  NOR U1966 ( .A(n90), .B(n162), .Z(n2154) );
  IV U1967 ( .A(n2154), .Z(n1882) );
  IV U1968 ( .A(n1874), .Z(n1875) );
  NOR U1969 ( .A(n1876), .B(n1875), .Z(n1880) );
  NOR U1970 ( .A(n1878), .B(n1877), .Z(n1879) );
  NOR U1971 ( .A(n1880), .B(n1879), .Z(n2161) );
  NOR U1972 ( .A(n164), .B(n102), .Z(n2159) );
  XOR U1973 ( .A(n2161), .B(n2159), .Z(n2163) );
  NOR U1974 ( .A(n166), .B(n101), .Z(n1881) );
  IV U1975 ( .A(n1881), .Z(n2162) );
  XOR U1976 ( .A(n2163), .B(n2162), .Z(n2153) );
  XOR U1977 ( .A(n1882), .B(n2153), .Z(n2155) );
  XOR U1978 ( .A(n2156), .B(n2155), .Z(n2150) );
  XOR U1979 ( .A(n2149), .B(n2150), .Z(n2140) );
  XOR U1980 ( .A(n1883), .B(n2140), .Z(n2142) );
  XOR U1981 ( .A(n2143), .B(n2142), .Z(n2171) );
  NOR U1982 ( .A(n104), .B(n157), .Z(n2169) );
  XOR U1983 ( .A(n2171), .B(n2169), .Z(n2172) );
  XOR U1984 ( .A(n2173), .B(n2172), .Z(n2134) );
  XOR U1985 ( .A(n2135), .B(n2134), .Z(n1884) );
  IV U1986 ( .A(n1884), .Z(n2136) );
  XOR U1987 ( .A(n2137), .B(n2136), .Z(n2131) );
  NOR U1988 ( .A(n1886), .B(n1885), .Z(n1890) );
  NOR U1989 ( .A(n1888), .B(n1887), .Z(n1889) );
  NOR U1990 ( .A(n1890), .B(n1889), .Z(n2129) );
  NOR U1991 ( .A(n106), .B(n152), .Z(n2127) );
  XOR U1992 ( .A(n2129), .B(n2127), .Z(n2130) );
  XOR U1993 ( .A(n2131), .B(n2130), .Z(n2121) );
  XOR U1994 ( .A(n2122), .B(n2121), .Z(n1891) );
  IV U1995 ( .A(n1891), .Z(n2123) );
  XOR U1996 ( .A(n2124), .B(n2123), .Z(n2180) );
  NOR U1997 ( .A(n107), .B(n149), .Z(n2178) );
  XOR U1998 ( .A(n2180), .B(n2178), .Z(n2181) );
  XOR U1999 ( .A(n2182), .B(n2181), .Z(n2114) );
  XOR U2000 ( .A(n1892), .B(n2114), .Z(n2117) );
  XOR U2001 ( .A(n2116), .B(n2117), .Z(n2187) );
  XOR U2002 ( .A(n2186), .B(n2187), .Z(n2189) );
  XOR U2003 ( .A(n2190), .B(n2189), .Z(n2108) );
  NOR U2004 ( .A(n109), .B(n142), .Z(n2106) );
  XOR U2005 ( .A(n2108), .B(n2106), .Z(n2109) );
  XOR U2006 ( .A(n2110), .B(n2109), .Z(n2101) );
  IV U2007 ( .A(n1893), .Z(n1894) );
  NOR U2008 ( .A(n1895), .B(n1894), .Z(n1900) );
  IV U2009 ( .A(n1896), .Z(n1897) );
  NOR U2010 ( .A(n1898), .B(n1897), .Z(n1899) );
  NOR U2011 ( .A(n1900), .B(n1899), .Z(n2100) );
  NOR U2012 ( .A(n110), .B(n140), .Z(n2098) );
  XOR U2013 ( .A(n2100), .B(n2098), .Z(n2103) );
  XOR U2014 ( .A(n2101), .B(n2103), .Z(n2093) );
  XOR U2015 ( .A(n2091), .B(n2093), .Z(n2094) );
  XOR U2016 ( .A(n1901), .B(n2094), .Z(n2086) );
  NOR U2017 ( .A(n111), .B(n136), .Z(n2087) );
  IV U2018 ( .A(n2087), .Z(n1902) );
  NOR U2019 ( .A(n2086), .B(n1902), .Z(n2090) );
  XOR U2020 ( .A(n1904), .B(n1903), .Z(n2083) );
  XOR U2021 ( .A(n1906), .B(n1905), .Z(n2070) );
  NOR U2022 ( .A(n109), .B(n136), .Z(n2069) );
  IV U2023 ( .A(n2069), .Z(n1907) );
  NOR U2024 ( .A(n2070), .B(n1907), .Z(n2072) );
  XOR U2025 ( .A(n1909), .B(n1908), .Z(n2066) );
  NOR U2026 ( .A(n108), .B(n136), .Z(n2065) );
  IV U2027 ( .A(n2065), .Z(n1910) );
  NOR U2028 ( .A(n2066), .B(n1910), .Z(n2068) );
  XOR U2029 ( .A(n1912), .B(n1911), .Z(n2062) );
  NOR U2030 ( .A(n87), .B(n136), .Z(n2061) );
  IV U2031 ( .A(n2061), .Z(n1913) );
  NOR U2032 ( .A(n2062), .B(n1913), .Z(n2064) );
  IV U2033 ( .A(n1914), .Z(n1916) );
  XOR U2034 ( .A(n1916), .B(n1915), .Z(n2057) );
  NOR U2035 ( .A(n107), .B(n136), .Z(n2058) );
  IV U2036 ( .A(n2058), .Z(n1917) );
  NOR U2037 ( .A(n2057), .B(n1917), .Z(n2060) );
  IV U2038 ( .A(n1918), .Z(n1920) );
  XOR U2039 ( .A(n1920), .B(n1919), .Z(n2053) );
  NOR U2040 ( .A(n88), .B(n136), .Z(n2054) );
  IV U2041 ( .A(n2054), .Z(n1921) );
  NOR U2042 ( .A(n2053), .B(n1921), .Z(n2056) );
  IV U2043 ( .A(n1922), .Z(n1924) );
  XOR U2044 ( .A(n1924), .B(n1923), .Z(n2049) );
  NOR U2045 ( .A(n106), .B(n136), .Z(n2050) );
  IV U2046 ( .A(n2050), .Z(n1925) );
  NOR U2047 ( .A(n2049), .B(n1925), .Z(n2052) );
  XOR U2048 ( .A(n1927), .B(n1926), .Z(n1928) );
  IV U2049 ( .A(n1928), .Z(n2045) );
  NOR U2050 ( .A(n105), .B(n136), .Z(n2046) );
  IV U2051 ( .A(n2046), .Z(n1929) );
  NOR U2052 ( .A(n2045), .B(n1929), .Z(n2048) );
  XOR U2053 ( .A(n1931), .B(n1930), .Z(n1932) );
  IV U2054 ( .A(n1932), .Z(n2041) );
  NOR U2055 ( .A(n104), .B(n136), .Z(n2042) );
  IV U2056 ( .A(n2042), .Z(n1933) );
  NOR U2057 ( .A(n2041), .B(n1933), .Z(n2044) );
  XOR U2058 ( .A(n1935), .B(n1934), .Z(n1936) );
  IV U2059 ( .A(n1936), .Z(n2037) );
  NOR U2060 ( .A(n89), .B(n136), .Z(n2038) );
  IV U2061 ( .A(n2038), .Z(n1937) );
  NOR U2062 ( .A(n2037), .B(n1937), .Z(n2040) );
  XOR U2063 ( .A(n1939), .B(n1938), .Z(n1940) );
  IV U2064 ( .A(n1940), .Z(n2033) );
  NOR U2065 ( .A(n103), .B(n136), .Z(n2034) );
  IV U2066 ( .A(n2034), .Z(n1941) );
  NOR U2067 ( .A(n2033), .B(n1941), .Z(n2036) );
  XOR U2068 ( .A(n1943), .B(n1942), .Z(n1944) );
  IV U2069 ( .A(n1944), .Z(n2029) );
  NOR U2070 ( .A(n90), .B(n136), .Z(n2030) );
  IV U2071 ( .A(n2030), .Z(n1945) );
  NOR U2072 ( .A(n2029), .B(n1945), .Z(n2032) );
  XOR U2073 ( .A(n1947), .B(n1946), .Z(n1948) );
  IV U2074 ( .A(n1948), .Z(n2025) );
  NOR U2075 ( .A(n102), .B(n136), .Z(n2026) );
  IV U2076 ( .A(n2026), .Z(n1949) );
  NOR U2077 ( .A(n2025), .B(n1949), .Z(n2028) );
  XOR U2078 ( .A(n1951), .B(n1950), .Z(n1952) );
  IV U2079 ( .A(n1952), .Z(n2021) );
  NOR U2080 ( .A(n101), .B(n136), .Z(n2022) );
  IV U2081 ( .A(n2022), .Z(n1953) );
  NOR U2082 ( .A(n2021), .B(n1953), .Z(n2024) );
  XOR U2083 ( .A(n1955), .B(n1954), .Z(n1956) );
  IV U2084 ( .A(n1956), .Z(n2017) );
  NOR U2085 ( .A(n100), .B(n136), .Z(n2018) );
  IV U2086 ( .A(n2018), .Z(n1957) );
  NOR U2087 ( .A(n2017), .B(n1957), .Z(n2020) );
  XOR U2088 ( .A(n1959), .B(n1958), .Z(n1960) );
  IV U2089 ( .A(n1960), .Z(n2013) );
  NOR U2090 ( .A(n99), .B(n136), .Z(n2014) );
  IV U2091 ( .A(n2014), .Z(n1961) );
  NOR U2092 ( .A(n2013), .B(n1961), .Z(n2016) );
  XOR U2093 ( .A(n1963), .B(n1962), .Z(n1964) );
  IV U2094 ( .A(n1964), .Z(n2009) );
  NOR U2095 ( .A(n98), .B(n136), .Z(n2010) );
  IV U2096 ( .A(n2010), .Z(n1965) );
  NOR U2097 ( .A(n2009), .B(n1965), .Z(n2012) );
  XOR U2098 ( .A(n1967), .B(n1966), .Z(n1968) );
  IV U2099 ( .A(n1968), .Z(n2005) );
  NOR U2100 ( .A(n91), .B(n136), .Z(n2006) );
  IV U2101 ( .A(n2006), .Z(n1969) );
  NOR U2102 ( .A(n2005), .B(n1969), .Z(n2008) );
  XOR U2103 ( .A(n1971), .B(n1970), .Z(n1972) );
  IV U2104 ( .A(n1972), .Z(n2001) );
  NOR U2105 ( .A(n97), .B(n136), .Z(n2002) );
  IV U2106 ( .A(n2002), .Z(n1973) );
  NOR U2107 ( .A(n2001), .B(n1973), .Z(n2004) );
  XOR U2108 ( .A(n1975), .B(n1974), .Z(n1976) );
  IV U2109 ( .A(n1976), .Z(n1997) );
  NOR U2110 ( .A(n96), .B(n136), .Z(n1998) );
  IV U2111 ( .A(n1998), .Z(n1977) );
  NOR U2112 ( .A(n1997), .B(n1977), .Z(n2000) );
  NOR U2113 ( .A(n93), .B(n136), .Z(n3407) );
  IV U2114 ( .A(n3407), .Z(n1979) );
  NOR U2115 ( .A(n138), .B(n168), .Z(n1982) );
  IV U2116 ( .A(n1982), .Z(n1978) );
  NOR U2117 ( .A(n1979), .B(n1978), .Z(n3054) );
  IV U2118 ( .A(n3054), .Z(n1980) );
  NOR U2119 ( .A(n1981), .B(n1980), .Z(n1989) );
  XOR U2120 ( .A(n1983), .B(n1982), .Z(n1984) );
  NOR U2121 ( .A(n3054), .B(n1984), .Z(n1985) );
  NOR U2122 ( .A(n1989), .B(n1985), .Z(n1986) );
  IV U2123 ( .A(n1986), .Z(n3067) );
  NOR U2124 ( .A(n94), .B(n136), .Z(n3066) );
  IV U2125 ( .A(n3066), .Z(n1987) );
  NOR U2126 ( .A(n3067), .B(n1987), .Z(n1988) );
  NOR U2127 ( .A(n1989), .B(n1988), .Z(n1991) );
  NOR U2128 ( .A(n95), .B(n136), .Z(n1992) );
  IV U2129 ( .A(n1992), .Z(n1990) );
  NOR U2130 ( .A(n1991), .B(n1990), .Z(n1996) );
  XOR U2131 ( .A(n1992), .B(n1991), .Z(n3047) );
  XOR U2132 ( .A(n1994), .B(n1993), .Z(n3048) );
  NOR U2133 ( .A(n3047), .B(n3048), .Z(n1995) );
  NOR U2134 ( .A(n1996), .B(n1995), .Z(n3043) );
  XOR U2135 ( .A(n1998), .B(n1997), .Z(n3044) );
  NOR U2136 ( .A(n3043), .B(n3044), .Z(n1999) );
  NOR U2137 ( .A(n2000), .B(n1999), .Z(n3039) );
  XOR U2138 ( .A(n2002), .B(n2001), .Z(n3040) );
  NOR U2139 ( .A(n3039), .B(n3040), .Z(n2003) );
  NOR U2140 ( .A(n2004), .B(n2003), .Z(n3035) );
  XOR U2141 ( .A(n2006), .B(n2005), .Z(n3036) );
  NOR U2142 ( .A(n3035), .B(n3036), .Z(n2007) );
  NOR U2143 ( .A(n2008), .B(n2007), .Z(n3031) );
  XOR U2144 ( .A(n2010), .B(n2009), .Z(n3032) );
  NOR U2145 ( .A(n3031), .B(n3032), .Z(n2011) );
  NOR U2146 ( .A(n2012), .B(n2011), .Z(n3027) );
  XOR U2147 ( .A(n2014), .B(n2013), .Z(n3028) );
  NOR U2148 ( .A(n3027), .B(n3028), .Z(n2015) );
  NOR U2149 ( .A(n2016), .B(n2015), .Z(n3023) );
  XOR U2150 ( .A(n2018), .B(n2017), .Z(n3024) );
  NOR U2151 ( .A(n3023), .B(n3024), .Z(n2019) );
  NOR U2152 ( .A(n2020), .B(n2019), .Z(n3019) );
  XOR U2153 ( .A(n2022), .B(n2021), .Z(n3020) );
  NOR U2154 ( .A(n3019), .B(n3020), .Z(n2023) );
  NOR U2155 ( .A(n2024), .B(n2023), .Z(n3015) );
  XOR U2156 ( .A(n2026), .B(n2025), .Z(n3016) );
  NOR U2157 ( .A(n3015), .B(n3016), .Z(n2027) );
  NOR U2158 ( .A(n2028), .B(n2027), .Z(n3011) );
  XOR U2159 ( .A(n2030), .B(n2029), .Z(n3012) );
  NOR U2160 ( .A(n3011), .B(n3012), .Z(n2031) );
  NOR U2161 ( .A(n2032), .B(n2031), .Z(n3007) );
  XOR U2162 ( .A(n2034), .B(n2033), .Z(n3008) );
  NOR U2163 ( .A(n3007), .B(n3008), .Z(n2035) );
  NOR U2164 ( .A(n2036), .B(n2035), .Z(n3003) );
  XOR U2165 ( .A(n2038), .B(n2037), .Z(n3004) );
  NOR U2166 ( .A(n3003), .B(n3004), .Z(n2039) );
  NOR U2167 ( .A(n2040), .B(n2039), .Z(n2999) );
  XOR U2168 ( .A(n2042), .B(n2041), .Z(n3000) );
  NOR U2169 ( .A(n2999), .B(n3000), .Z(n2043) );
  NOR U2170 ( .A(n2044), .B(n2043), .Z(n2995) );
  XOR U2171 ( .A(n2046), .B(n2045), .Z(n2996) );
  NOR U2172 ( .A(n2995), .B(n2996), .Z(n2047) );
  NOR U2173 ( .A(n2048), .B(n2047), .Z(n2991) );
  XOR U2174 ( .A(n2050), .B(n2049), .Z(n2992) );
  NOR U2175 ( .A(n2991), .B(n2992), .Z(n2051) );
  NOR U2176 ( .A(n2052), .B(n2051), .Z(n2988) );
  XOR U2177 ( .A(n2054), .B(n2053), .Z(n2987) );
  NOR U2178 ( .A(n2988), .B(n2987), .Z(n2055) );
  NOR U2179 ( .A(n2056), .B(n2055), .Z(n2983) );
  XOR U2180 ( .A(n2058), .B(n2057), .Z(n2984) );
  NOR U2181 ( .A(n2983), .B(n2984), .Z(n2059) );
  NOR U2182 ( .A(n2060), .B(n2059), .Z(n2982) );
  XOR U2183 ( .A(n2062), .B(n2061), .Z(n2981) );
  NOR U2184 ( .A(n2982), .B(n2981), .Z(n2063) );
  NOR U2185 ( .A(n2064), .B(n2063), .Z(n2980) );
  XOR U2186 ( .A(n2066), .B(n2065), .Z(n2979) );
  NOR U2187 ( .A(n2980), .B(n2979), .Z(n2067) );
  NOR U2188 ( .A(n2068), .B(n2067), .Z(n2978) );
  XOR U2189 ( .A(n2070), .B(n2069), .Z(n2977) );
  NOR U2190 ( .A(n2978), .B(n2977), .Z(n2071) );
  NOR U2191 ( .A(n2072), .B(n2071), .Z(n2075) );
  XOR U2192 ( .A(n2074), .B(n2073), .Z(n2076) );
  NOR U2193 ( .A(n2075), .B(n2076), .Z(n2080) );
  IV U2194 ( .A(n2075), .Z(n2077) );
  XOR U2195 ( .A(n2077), .B(n2076), .Z(n2976) );
  NOR U2196 ( .A(n110), .B(n136), .Z(n2078) );
  IV U2197 ( .A(n2078), .Z(n2975) );
  NOR U2198 ( .A(n2976), .B(n2975), .Z(n2079) );
  NOR U2199 ( .A(n2080), .B(n2079), .Z(n2082) );
  IV U2200 ( .A(n2082), .Z(n2081) );
  NOR U2201 ( .A(n2083), .B(n2081), .Z(n2085) );
  NOR U2202 ( .A(n86), .B(n136), .Z(n2971) );
  XOR U2203 ( .A(n2083), .B(n2082), .Z(n2970) );
  NOR U2204 ( .A(n2971), .B(n2970), .Z(n2084) );
  NOR U2205 ( .A(n2085), .B(n2084), .Z(n2968) );
  IV U2206 ( .A(n2968), .Z(n2088) );
  XOR U2207 ( .A(n2087), .B(n2086), .Z(n2967) );
  NOR U2208 ( .A(n2088), .B(n2967), .Z(n2089) );
  NOR U2209 ( .A(n2090), .B(n2089), .Z(n2198) );
  IV U2210 ( .A(n2091), .Z(n2092) );
  NOR U2211 ( .A(n2093), .B(n2092), .Z(n2097) );
  NOR U2212 ( .A(n2095), .B(n2094), .Z(n2096) );
  NOR U2213 ( .A(n2097), .B(n2096), .Z(n2206) );
  NOR U2214 ( .A(n111), .B(n138), .Z(n2202) );
  NOR U2215 ( .A(n86), .B(n140), .Z(n2301) );
  IV U2216 ( .A(n2098), .Z(n2099) );
  NOR U2217 ( .A(n2100), .B(n2099), .Z(n2105) );
  IV U2218 ( .A(n2101), .Z(n2102) );
  NOR U2219 ( .A(n2103), .B(n2102), .Z(n2104) );
  NOR U2220 ( .A(n2105), .B(n2104), .Z(n2299) );
  IV U2221 ( .A(n2299), .Z(n2195) );
  IV U2222 ( .A(n2106), .Z(n2107) );
  NOR U2223 ( .A(n2108), .B(n2107), .Z(n2112) );
  NOR U2224 ( .A(n2110), .B(n2109), .Z(n2111) );
  NOR U2225 ( .A(n2112), .B(n2111), .Z(n2113) );
  IV U2226 ( .A(n2113), .Z(n2213) );
  NOR U2227 ( .A(n110), .B(n142), .Z(n2211) );
  NOR U2228 ( .A(n2115), .B(n2114), .Z(n2120) );
  IV U2229 ( .A(n2116), .Z(n2118) );
  NOR U2230 ( .A(n2118), .B(n2117), .Z(n2119) );
  NOR U2231 ( .A(n2120), .B(n2119), .Z(n2219) );
  NOR U2232 ( .A(n108), .B(n146), .Z(n2217) );
  NOR U2233 ( .A(n2122), .B(n2121), .Z(n2126) );
  NOR U2234 ( .A(n2124), .B(n2123), .Z(n2125) );
  NOR U2235 ( .A(n2126), .B(n2125), .Z(n2232) );
  NOR U2236 ( .A(n107), .B(n151), .Z(n2230) );
  IV U2237 ( .A(n2127), .Z(n2128) );
  NOR U2238 ( .A(n2129), .B(n2128), .Z(n2133) );
  NOR U2239 ( .A(n2131), .B(n2130), .Z(n2132) );
  NOR U2240 ( .A(n2133), .B(n2132), .Z(n2284) );
  NOR U2241 ( .A(n2135), .B(n2134), .Z(n2139) );
  NOR U2242 ( .A(n2137), .B(n2136), .Z(n2138) );
  NOR U2243 ( .A(n2139), .B(n2138), .Z(n2238) );
  NOR U2244 ( .A(n106), .B(n154), .Z(n2236) );
  NOR U2245 ( .A(n2141), .B(n2140), .Z(n2145) );
  NOR U2246 ( .A(n2143), .B(n2142), .Z(n2144) );
  NOR U2247 ( .A(n2145), .B(n2144), .Z(n2251) );
  NOR U2248 ( .A(n104), .B(n159), .Z(n2249) );
  IV U2249 ( .A(n2146), .Z(n2147) );
  NOR U2250 ( .A(n2148), .B(n2147), .Z(n2152) );
  NOR U2251 ( .A(n2150), .B(n2149), .Z(n2151) );
  NOR U2252 ( .A(n2152), .B(n2151), .Z(n2273) );
  NOR U2253 ( .A(n2154), .B(n2153), .Z(n2158) );
  NOR U2254 ( .A(n2156), .B(n2155), .Z(n2157) );
  NOR U2255 ( .A(n2158), .B(n2157), .Z(n2257) );
  NOR U2256 ( .A(n103), .B(n162), .Z(n2255) );
  IV U2257 ( .A(n2255), .Z(n2167) );
  IV U2258 ( .A(n2159), .Z(n2160) );
  NOR U2259 ( .A(n2161), .B(n2160), .Z(n2165) );
  NOR U2260 ( .A(n2163), .B(n2162), .Z(n2164) );
  NOR U2261 ( .A(n2165), .B(n2164), .Z(n2262) );
  NOR U2262 ( .A(n164), .B(n90), .Z(n2260) );
  XOR U2263 ( .A(n2262), .B(n2260), .Z(n2264) );
  NOR U2264 ( .A(n166), .B(n102), .Z(n2166) );
  IV U2265 ( .A(n2166), .Z(n2263) );
  XOR U2266 ( .A(n2264), .B(n2263), .Z(n2254) );
  XOR U2267 ( .A(n2167), .B(n2254), .Z(n2256) );
  XOR U2268 ( .A(n2257), .B(n2256), .Z(n2271) );
  NOR U2269 ( .A(n89), .B(n160), .Z(n2269) );
  XOR U2270 ( .A(n2271), .B(n2269), .Z(n2272) );
  XOR U2271 ( .A(n2273), .B(n2272), .Z(n2248) );
  XOR U2272 ( .A(n2249), .B(n2248), .Z(n2168) );
  IV U2273 ( .A(n2168), .Z(n2250) );
  XOR U2274 ( .A(n2251), .B(n2250), .Z(n2245) );
  IV U2275 ( .A(n2169), .Z(n2170) );
  NOR U2276 ( .A(n2171), .B(n2170), .Z(n2175) );
  NOR U2277 ( .A(n2173), .B(n2172), .Z(n2174) );
  NOR U2278 ( .A(n2175), .B(n2174), .Z(n2243) );
  NOR U2279 ( .A(n105), .B(n157), .Z(n2241) );
  XOR U2280 ( .A(n2243), .B(n2241), .Z(n2244) );
  XOR U2281 ( .A(n2245), .B(n2244), .Z(n2235) );
  XOR U2282 ( .A(n2236), .B(n2235), .Z(n2176) );
  IV U2283 ( .A(n2176), .Z(n2237) );
  XOR U2284 ( .A(n2238), .B(n2237), .Z(n2282) );
  NOR U2285 ( .A(n88), .B(n152), .Z(n2280) );
  XOR U2286 ( .A(n2282), .B(n2280), .Z(n2283) );
  XOR U2287 ( .A(n2284), .B(n2283), .Z(n2229) );
  XOR U2288 ( .A(n2230), .B(n2229), .Z(n2177) );
  IV U2289 ( .A(n2177), .Z(n2231) );
  XOR U2290 ( .A(n2232), .B(n2231), .Z(n2226) );
  IV U2291 ( .A(n2178), .Z(n2179) );
  NOR U2292 ( .A(n2180), .B(n2179), .Z(n2184) );
  NOR U2293 ( .A(n2182), .B(n2181), .Z(n2183) );
  NOR U2294 ( .A(n2184), .B(n2183), .Z(n2224) );
  NOR U2295 ( .A(n87), .B(n149), .Z(n2222) );
  XOR U2296 ( .A(n2224), .B(n2222), .Z(n2225) );
  XOR U2297 ( .A(n2226), .B(n2225), .Z(n2216) );
  XOR U2298 ( .A(n2217), .B(n2216), .Z(n2185) );
  IV U2299 ( .A(n2185), .Z(n2218) );
  XOR U2300 ( .A(n2219), .B(n2218), .Z(n2293) );
  NOR U2301 ( .A(n109), .B(n144), .Z(n2291) );
  XOR U2302 ( .A(n2293), .B(n2291), .Z(n2295) );
  IV U2303 ( .A(n2186), .Z(n2188) );
  NOR U2304 ( .A(n2188), .B(n2187), .Z(n2192) );
  NOR U2305 ( .A(n2190), .B(n2189), .Z(n2191) );
  NOR U2306 ( .A(n2192), .B(n2191), .Z(n2193) );
  IV U2307 ( .A(n2193), .Z(n2294) );
  XOR U2308 ( .A(n2295), .B(n2294), .Z(n2210) );
  XOR U2309 ( .A(n2211), .B(n2210), .Z(n2194) );
  IV U2310 ( .A(n2194), .Z(n2212) );
  XOR U2311 ( .A(n2213), .B(n2212), .Z(n2300) );
  XOR U2312 ( .A(n2195), .B(n2300), .Z(n2303) );
  XOR U2313 ( .A(n2301), .B(n2303), .Z(n2204) );
  XOR U2314 ( .A(n2202), .B(n2204), .Z(n2205) );
  XOR U2315 ( .A(n2206), .B(n2205), .Z(n2197) );
  IV U2316 ( .A(n2197), .Z(n2196) );
  NOR U2317 ( .A(n2198), .B(n2196), .Z(n2201) );
  XOR U2318 ( .A(n2198), .B(n2197), .Z(n2964) );
  NOR U2319 ( .A(n85), .B(n136), .Z(n2965) );
  IV U2320 ( .A(n2965), .Z(n2199) );
  NOR U2321 ( .A(n2964), .B(n2199), .Z(n2200) );
  NOR U2322 ( .A(n2201), .B(n2200), .Z(n2308) );
  IV U2323 ( .A(n2308), .Z(n2306) );
  IV U2324 ( .A(n2202), .Z(n2203) );
  NOR U2325 ( .A(n2204), .B(n2203), .Z(n2208) );
  NOR U2326 ( .A(n2206), .B(n2205), .Z(n2207) );
  NOR U2327 ( .A(n2208), .B(n2207), .Z(n2209) );
  IV U2328 ( .A(n2209), .Z(n2317) );
  NOR U2329 ( .A(n85), .B(n138), .Z(n2314) );
  NOR U2330 ( .A(n2211), .B(n2210), .Z(n2215) );
  NOR U2331 ( .A(n2213), .B(n2212), .Z(n2214) );
  NOR U2332 ( .A(n2215), .B(n2214), .Z(n2330) );
  NOR U2333 ( .A(n86), .B(n142), .Z(n2328) );
  NOR U2334 ( .A(n2217), .B(n2216), .Z(n2221) );
  NOR U2335 ( .A(n2219), .B(n2218), .Z(n2220) );
  NOR U2336 ( .A(n2221), .B(n2220), .Z(n2343) );
  NOR U2337 ( .A(n109), .B(n146), .Z(n2341) );
  IV U2338 ( .A(n2341), .Z(n2290) );
  IV U2339 ( .A(n2222), .Z(n2223) );
  NOR U2340 ( .A(n2224), .B(n2223), .Z(n2228) );
  NOR U2341 ( .A(n2226), .B(n2225), .Z(n2227) );
  NOR U2342 ( .A(n2228), .B(n2227), .Z(n2346) );
  IV U2343 ( .A(n2346), .Z(n2288) );
  NOR U2344 ( .A(n2230), .B(n2229), .Z(n2234) );
  NOR U2345 ( .A(n2232), .B(n2231), .Z(n2233) );
  NOR U2346 ( .A(n2234), .B(n2233), .Z(n2355) );
  NOR U2347 ( .A(n87), .B(n151), .Z(n2353) );
  IV U2348 ( .A(n2353), .Z(n2287) );
  NOR U2349 ( .A(n2236), .B(n2235), .Z(n2240) );
  NOR U2350 ( .A(n2238), .B(n2237), .Z(n2239) );
  NOR U2351 ( .A(n2240), .B(n2239), .Z(n2368) );
  NOR U2352 ( .A(n88), .B(n154), .Z(n2366) );
  IV U2353 ( .A(n2366), .Z(n2279) );
  IV U2354 ( .A(n2241), .Z(n2242) );
  NOR U2355 ( .A(n2243), .B(n2242), .Z(n2247) );
  NOR U2356 ( .A(n2245), .B(n2244), .Z(n2246) );
  NOR U2357 ( .A(n2247), .B(n2246), .Z(n2371) );
  IV U2358 ( .A(n2371), .Z(n2277) );
  NOR U2359 ( .A(n2249), .B(n2248), .Z(n2253) );
  NOR U2360 ( .A(n2251), .B(n2250), .Z(n2252) );
  NOR U2361 ( .A(n2253), .B(n2252), .Z(n2380) );
  NOR U2362 ( .A(n105), .B(n159), .Z(n2378) );
  IV U2363 ( .A(n2378), .Z(n2276) );
  NOR U2364 ( .A(n2255), .B(n2254), .Z(n2259) );
  NOR U2365 ( .A(n2257), .B(n2256), .Z(n2258) );
  NOR U2366 ( .A(n2259), .B(n2258), .Z(n2393) );
  NOR U2367 ( .A(n89), .B(n162), .Z(n2391) );
  IV U2368 ( .A(n2391), .Z(n2268) );
  IV U2369 ( .A(n2260), .Z(n2261) );
  NOR U2370 ( .A(n2262), .B(n2261), .Z(n2266) );
  NOR U2371 ( .A(n2264), .B(n2263), .Z(n2265) );
  NOR U2372 ( .A(n2266), .B(n2265), .Z(n2398) );
  NOR U2373 ( .A(n164), .B(n103), .Z(n2396) );
  XOR U2374 ( .A(n2398), .B(n2396), .Z(n2400) );
  NOR U2375 ( .A(n166), .B(n90), .Z(n2267) );
  IV U2376 ( .A(n2267), .Z(n2399) );
  XOR U2377 ( .A(n2400), .B(n2399), .Z(n2390) );
  XOR U2378 ( .A(n2268), .B(n2390), .Z(n2392) );
  XOR U2379 ( .A(n2393), .B(n2392), .Z(n2387) );
  IV U2380 ( .A(n2269), .Z(n2270) );
  NOR U2381 ( .A(n2271), .B(n2270), .Z(n2275) );
  NOR U2382 ( .A(n2273), .B(n2272), .Z(n2274) );
  NOR U2383 ( .A(n2275), .B(n2274), .Z(n2385) );
  NOR U2384 ( .A(n104), .B(n160), .Z(n2383) );
  XOR U2385 ( .A(n2385), .B(n2383), .Z(n2386) );
  XOR U2386 ( .A(n2387), .B(n2386), .Z(n2377) );
  XOR U2387 ( .A(n2276), .B(n2377), .Z(n2379) );
  XOR U2388 ( .A(n2380), .B(n2379), .Z(n2372) );
  XOR U2389 ( .A(n2277), .B(n2372), .Z(n2374) );
  NOR U2390 ( .A(n106), .B(n157), .Z(n2278) );
  IV U2391 ( .A(n2278), .Z(n2373) );
  XOR U2392 ( .A(n2374), .B(n2373), .Z(n2365) );
  XOR U2393 ( .A(n2279), .B(n2365), .Z(n2367) );
  XOR U2394 ( .A(n2368), .B(n2367), .Z(n2362) );
  IV U2395 ( .A(n2280), .Z(n2281) );
  NOR U2396 ( .A(n2282), .B(n2281), .Z(n2286) );
  NOR U2397 ( .A(n2284), .B(n2283), .Z(n2285) );
  NOR U2398 ( .A(n2286), .B(n2285), .Z(n2360) );
  NOR U2399 ( .A(n107), .B(n152), .Z(n2358) );
  XOR U2400 ( .A(n2360), .B(n2358), .Z(n2361) );
  XOR U2401 ( .A(n2362), .B(n2361), .Z(n2352) );
  XOR U2402 ( .A(n2287), .B(n2352), .Z(n2354) );
  XOR U2403 ( .A(n2355), .B(n2354), .Z(n2347) );
  XOR U2404 ( .A(n2288), .B(n2347), .Z(n2349) );
  NOR U2405 ( .A(n108), .B(n149), .Z(n2289) );
  IV U2406 ( .A(n2289), .Z(n2348) );
  XOR U2407 ( .A(n2349), .B(n2348), .Z(n2340) );
  XOR U2408 ( .A(n2290), .B(n2340), .Z(n2342) );
  XOR U2409 ( .A(n2343), .B(n2342), .Z(n2337) );
  IV U2410 ( .A(n2291), .Z(n2292) );
  NOR U2411 ( .A(n2293), .B(n2292), .Z(n2297) );
  NOR U2412 ( .A(n2295), .B(n2294), .Z(n2296) );
  NOR U2413 ( .A(n2297), .B(n2296), .Z(n2335) );
  NOR U2414 ( .A(n110), .B(n144), .Z(n2333) );
  XOR U2415 ( .A(n2335), .B(n2333), .Z(n2336) );
  XOR U2416 ( .A(n2337), .B(n2336), .Z(n2327) );
  XOR U2417 ( .A(n2328), .B(n2327), .Z(n2298) );
  IV U2418 ( .A(n2298), .Z(n2329) );
  XOR U2419 ( .A(n2330), .B(n2329), .Z(n2324) );
  NOR U2420 ( .A(n2300), .B(n2299), .Z(n2305) );
  IV U2421 ( .A(n2301), .Z(n2302) );
  NOR U2422 ( .A(n2303), .B(n2302), .Z(n2304) );
  NOR U2423 ( .A(n2305), .B(n2304), .Z(n2322) );
  NOR U2424 ( .A(n111), .B(n140), .Z(n2320) );
  XOR U2425 ( .A(n2322), .B(n2320), .Z(n2323) );
  XOR U2426 ( .A(n2324), .B(n2323), .Z(n2313) );
  XOR U2427 ( .A(n2314), .B(n2313), .Z(n2315) );
  XOR U2428 ( .A(n2317), .B(n2315), .Z(n2307) );
  NOR U2429 ( .A(n2306), .B(n2307), .Z(n2310) );
  NOR U2430 ( .A(n112), .B(n136), .Z(n2962) );
  XOR U2431 ( .A(n2308), .B(n2307), .Z(n2961) );
  NOR U2432 ( .A(n2962), .B(n2961), .Z(n2309) );
  NOR U2433 ( .A(n2310), .B(n2309), .Z(n2311) );
  IV U2434 ( .A(n2311), .Z(n2414) );
  NOR U2435 ( .A(n84), .B(n136), .Z(n2413) );
  IV U2436 ( .A(n2413), .Z(n2312) );
  NOR U2437 ( .A(n2414), .B(n2312), .Z(n2416) );
  NOR U2438 ( .A(n2314), .B(n2313), .Z(n2319) );
  IV U2439 ( .A(n2315), .Z(n2316) );
  NOR U2440 ( .A(n2317), .B(n2316), .Z(n2318) );
  NOR U2441 ( .A(n2319), .B(n2318), .Z(n2421) );
  NOR U2442 ( .A(n112), .B(n138), .Z(n2419) );
  IV U2443 ( .A(n2419), .Z(n2412) );
  IV U2444 ( .A(n2320), .Z(n2321) );
  NOR U2445 ( .A(n2322), .B(n2321), .Z(n2326) );
  NOR U2446 ( .A(n2324), .B(n2323), .Z(n2325) );
  NOR U2447 ( .A(n2326), .B(n2325), .Z(n2516) );
  IV U2448 ( .A(n2516), .Z(n2410) );
  NOR U2449 ( .A(n2328), .B(n2327), .Z(n2332) );
  NOR U2450 ( .A(n2330), .B(n2329), .Z(n2331) );
  NOR U2451 ( .A(n2332), .B(n2331), .Z(n2427) );
  NOR U2452 ( .A(n111), .B(n142), .Z(n2424) );
  NOR U2453 ( .A(n86), .B(n144), .Z(n2435) );
  IV U2454 ( .A(n2333), .Z(n2334) );
  NOR U2455 ( .A(n2335), .B(n2334), .Z(n2339) );
  NOR U2456 ( .A(n2337), .B(n2336), .Z(n2338) );
  NOR U2457 ( .A(n2339), .B(n2338), .Z(n2434) );
  IV U2458 ( .A(n2434), .Z(n2409) );
  NOR U2459 ( .A(n2341), .B(n2340), .Z(n2345) );
  NOR U2460 ( .A(n2343), .B(n2342), .Z(n2344) );
  NOR U2461 ( .A(n2345), .B(n2344), .Z(n2444) );
  NOR U2462 ( .A(n110), .B(n146), .Z(n2441) );
  NOR U2463 ( .A(n109), .B(n149), .Z(n2452) );
  NOR U2464 ( .A(n2347), .B(n2346), .Z(n2351) );
  NOR U2465 ( .A(n2349), .B(n2348), .Z(n2350) );
  NOR U2466 ( .A(n2351), .B(n2350), .Z(n2450) );
  IV U2467 ( .A(n2450), .Z(n2408) );
  NOR U2468 ( .A(n2353), .B(n2352), .Z(n2357) );
  NOR U2469 ( .A(n2355), .B(n2354), .Z(n2356) );
  NOR U2470 ( .A(n2357), .B(n2356), .Z(n2460) );
  NOR U2471 ( .A(n108), .B(n151), .Z(n2458) );
  IV U2472 ( .A(n2458), .Z(n2407) );
  IV U2473 ( .A(n2358), .Z(n2359) );
  NOR U2474 ( .A(n2360), .B(n2359), .Z(n2364) );
  NOR U2475 ( .A(n2362), .B(n2361), .Z(n2363) );
  NOR U2476 ( .A(n2364), .B(n2363), .Z(n2510) );
  NOR U2477 ( .A(n2366), .B(n2365), .Z(n2370) );
  NOR U2478 ( .A(n2368), .B(n2367), .Z(n2369) );
  NOR U2479 ( .A(n2370), .B(n2369), .Z(n2466) );
  NOR U2480 ( .A(n107), .B(n154), .Z(n2464) );
  NOR U2481 ( .A(n2372), .B(n2371), .Z(n2376) );
  NOR U2482 ( .A(n2374), .B(n2373), .Z(n2375) );
  NOR U2483 ( .A(n2376), .B(n2375), .Z(n2473) );
  NOR U2484 ( .A(n2378), .B(n2377), .Z(n2382) );
  NOR U2485 ( .A(n2380), .B(n2379), .Z(n2381) );
  NOR U2486 ( .A(n2382), .B(n2381), .Z(n2479) );
  NOR U2487 ( .A(n106), .B(n159), .Z(n2477) );
  IV U2488 ( .A(n2383), .Z(n2384) );
  NOR U2489 ( .A(n2385), .B(n2384), .Z(n2389) );
  NOR U2490 ( .A(n2387), .B(n2386), .Z(n2388) );
  NOR U2491 ( .A(n2389), .B(n2388), .Z(n2501) );
  NOR U2492 ( .A(n2391), .B(n2390), .Z(n2395) );
  NOR U2493 ( .A(n2393), .B(n2392), .Z(n2394) );
  NOR U2494 ( .A(n2395), .B(n2394), .Z(n2485) );
  NOR U2495 ( .A(n104), .B(n162), .Z(n2483) );
  IV U2496 ( .A(n2483), .Z(n2404) );
  IV U2497 ( .A(n2396), .Z(n2397) );
  NOR U2498 ( .A(n2398), .B(n2397), .Z(n2402) );
  NOR U2499 ( .A(n2400), .B(n2399), .Z(n2401) );
  NOR U2500 ( .A(n2402), .B(n2401), .Z(n2490) );
  NOR U2501 ( .A(n164), .B(n89), .Z(n2488) );
  XOR U2502 ( .A(n2490), .B(n2488), .Z(n2492) );
  NOR U2503 ( .A(n166), .B(n103), .Z(n2403) );
  IV U2504 ( .A(n2403), .Z(n2491) );
  XOR U2505 ( .A(n2492), .B(n2491), .Z(n2482) );
  XOR U2506 ( .A(n2404), .B(n2482), .Z(n2484) );
  XOR U2507 ( .A(n2485), .B(n2484), .Z(n2499) );
  NOR U2508 ( .A(n105), .B(n160), .Z(n2497) );
  XOR U2509 ( .A(n2499), .B(n2497), .Z(n2500) );
  XOR U2510 ( .A(n2501), .B(n2500), .Z(n2476) );
  XOR U2511 ( .A(n2477), .B(n2476), .Z(n2405) );
  IV U2512 ( .A(n2405), .Z(n2478) );
  XOR U2513 ( .A(n2479), .B(n2478), .Z(n2471) );
  NOR U2514 ( .A(n88), .B(n157), .Z(n2469) );
  XOR U2515 ( .A(n2471), .B(n2469), .Z(n2472) );
  XOR U2516 ( .A(n2473), .B(n2472), .Z(n2463) );
  XOR U2517 ( .A(n2464), .B(n2463), .Z(n2406) );
  IV U2518 ( .A(n2406), .Z(n2465) );
  XOR U2519 ( .A(n2466), .B(n2465), .Z(n2508) );
  NOR U2520 ( .A(n87), .B(n152), .Z(n2506) );
  XOR U2521 ( .A(n2508), .B(n2506), .Z(n2509) );
  XOR U2522 ( .A(n2510), .B(n2509), .Z(n2457) );
  XOR U2523 ( .A(n2407), .B(n2457), .Z(n2459) );
  XOR U2524 ( .A(n2460), .B(n2459), .Z(n2451) );
  XOR U2525 ( .A(n2408), .B(n2451), .Z(n2454) );
  XOR U2526 ( .A(n2452), .B(n2454), .Z(n2443) );
  XOR U2527 ( .A(n2441), .B(n2443), .Z(n2446) );
  XOR U2528 ( .A(n2444), .B(n2446), .Z(n2433) );
  XOR U2529 ( .A(n2409), .B(n2433), .Z(n2437) );
  XOR U2530 ( .A(n2435), .B(n2437), .Z(n2426) );
  XOR U2531 ( .A(n2424), .B(n2426), .Z(n2429) );
  XOR U2532 ( .A(n2427), .B(n2429), .Z(n2515) );
  XOR U2533 ( .A(n2410), .B(n2515), .Z(n2518) );
  NOR U2534 ( .A(n85), .B(n140), .Z(n2411) );
  IV U2535 ( .A(n2411), .Z(n2517) );
  XOR U2536 ( .A(n2518), .B(n2517), .Z(n2418) );
  XOR U2537 ( .A(n2412), .B(n2418), .Z(n2420) );
  XOR U2538 ( .A(n2421), .B(n2420), .Z(n2959) );
  XOR U2539 ( .A(n2414), .B(n2413), .Z(n2960) );
  NOR U2540 ( .A(n2959), .B(n2960), .Z(n2415) );
  NOR U2541 ( .A(n2416), .B(n2415), .Z(n2523) );
  NOR U2542 ( .A(n113), .B(n136), .Z(n2522) );
  IV U2543 ( .A(n2522), .Z(n2417) );
  NOR U2544 ( .A(n2523), .B(n2417), .Z(n2525) );
  NOR U2545 ( .A(n2419), .B(n2418), .Z(n2423) );
  NOR U2546 ( .A(n2421), .B(n2420), .Z(n2422) );
  NOR U2547 ( .A(n2423), .B(n2422), .Z(n2530) );
  NOR U2548 ( .A(n84), .B(n138), .Z(n2528) );
  IV U2549 ( .A(n2424), .Z(n2425) );
  NOR U2550 ( .A(n2426), .B(n2425), .Z(n2431) );
  IV U2551 ( .A(n2427), .Z(n2428) );
  NOR U2552 ( .A(n2429), .B(n2428), .Z(n2430) );
  NOR U2553 ( .A(n2431), .B(n2430), .Z(n2432) );
  IV U2554 ( .A(n2432), .Z(n2536) );
  NOR U2555 ( .A(n85), .B(n142), .Z(n2534) );
  NOR U2556 ( .A(n2434), .B(n2433), .Z(n2439) );
  IV U2557 ( .A(n2435), .Z(n2436) );
  NOR U2558 ( .A(n2437), .B(n2436), .Z(n2438) );
  NOR U2559 ( .A(n2439), .B(n2438), .Z(n2440) );
  IV U2560 ( .A(n2440), .Z(n2542) );
  NOR U2561 ( .A(n111), .B(n144), .Z(n2540) );
  IV U2562 ( .A(n2441), .Z(n2442) );
  NOR U2563 ( .A(n2443), .B(n2442), .Z(n2448) );
  IV U2564 ( .A(n2444), .Z(n2445) );
  NOR U2565 ( .A(n2446), .B(n2445), .Z(n2447) );
  NOR U2566 ( .A(n2448), .B(n2447), .Z(n2449) );
  IV U2567 ( .A(n2449), .Z(n2551) );
  NOR U2568 ( .A(n86), .B(n146), .Z(n2548) );
  NOR U2569 ( .A(n2451), .B(n2450), .Z(n2456) );
  IV U2570 ( .A(n2452), .Z(n2453) );
  NOR U2571 ( .A(n2454), .B(n2453), .Z(n2455) );
  NOR U2572 ( .A(n2456), .B(n2455), .Z(n2617) );
  NOR U2573 ( .A(n2458), .B(n2457), .Z(n2462) );
  NOR U2574 ( .A(n2460), .B(n2459), .Z(n2461) );
  NOR U2575 ( .A(n2462), .B(n2461), .Z(n2557) );
  NOR U2576 ( .A(n109), .B(n151), .Z(n2555) );
  NOR U2577 ( .A(n2464), .B(n2463), .Z(n2468) );
  NOR U2578 ( .A(n2466), .B(n2465), .Z(n2467) );
  NOR U2579 ( .A(n2468), .B(n2467), .Z(n2563) );
  NOR U2580 ( .A(n87), .B(n154), .Z(n2561) );
  IV U2581 ( .A(n2561), .Z(n2505) );
  IV U2582 ( .A(n2469), .Z(n2470) );
  NOR U2583 ( .A(n2471), .B(n2470), .Z(n2475) );
  NOR U2584 ( .A(n2473), .B(n2472), .Z(n2474) );
  NOR U2585 ( .A(n2475), .B(n2474), .Z(n2568) );
  NOR U2586 ( .A(n107), .B(n157), .Z(n2567) );
  NOR U2587 ( .A(n2477), .B(n2476), .Z(n2481) );
  NOR U2588 ( .A(n2479), .B(n2478), .Z(n2480) );
  NOR U2589 ( .A(n2481), .B(n2480), .Z(n2578) );
  NOR U2590 ( .A(n88), .B(n159), .Z(n2575) );
  NOR U2591 ( .A(n2483), .B(n2482), .Z(n2487) );
  NOR U2592 ( .A(n2485), .B(n2484), .Z(n2486) );
  NOR U2593 ( .A(n2487), .B(n2486), .Z(n2584) );
  NOR U2594 ( .A(n105), .B(n162), .Z(n2582) );
  IV U2595 ( .A(n2582), .Z(n2496) );
  IV U2596 ( .A(n2488), .Z(n2489) );
  NOR U2597 ( .A(n2490), .B(n2489), .Z(n2494) );
  NOR U2598 ( .A(n2492), .B(n2491), .Z(n2493) );
  NOR U2599 ( .A(n2494), .B(n2493), .Z(n2589) );
  NOR U2600 ( .A(n164), .B(n104), .Z(n2587) );
  XOR U2601 ( .A(n2589), .B(n2587), .Z(n2591) );
  NOR U2602 ( .A(n166), .B(n89), .Z(n2495) );
  IV U2603 ( .A(n2495), .Z(n2590) );
  XOR U2604 ( .A(n2591), .B(n2590), .Z(n2581) );
  XOR U2605 ( .A(n2496), .B(n2581), .Z(n2583) );
  XOR U2606 ( .A(n2584), .B(n2583), .Z(n2600) );
  IV U2607 ( .A(n2497), .Z(n2498) );
  NOR U2608 ( .A(n2499), .B(n2498), .Z(n2503) );
  NOR U2609 ( .A(n2501), .B(n2500), .Z(n2502) );
  NOR U2610 ( .A(n2503), .B(n2502), .Z(n2598) );
  NOR U2611 ( .A(n106), .B(n160), .Z(n2596) );
  XOR U2612 ( .A(n2598), .B(n2596), .Z(n2599) );
  XOR U2613 ( .A(n2600), .B(n2599), .Z(n2574) );
  XOR U2614 ( .A(n2575), .B(n2574), .Z(n2576) );
  XOR U2615 ( .A(n2578), .B(n2576), .Z(n2566) );
  XOR U2616 ( .A(n2567), .B(n2566), .Z(n2504) );
  IV U2617 ( .A(n2504), .Z(n2569) );
  XOR U2618 ( .A(n2568), .B(n2569), .Z(n2560) );
  XOR U2619 ( .A(n2505), .B(n2560), .Z(n2562) );
  XOR U2620 ( .A(n2563), .B(n2562), .Z(n2609) );
  IV U2621 ( .A(n2506), .Z(n2507) );
  NOR U2622 ( .A(n2508), .B(n2507), .Z(n2512) );
  NOR U2623 ( .A(n2510), .B(n2509), .Z(n2511) );
  NOR U2624 ( .A(n2512), .B(n2511), .Z(n2607) );
  NOR U2625 ( .A(n108), .B(n152), .Z(n2605) );
  XOR U2626 ( .A(n2607), .B(n2605), .Z(n2608) );
  XOR U2627 ( .A(n2609), .B(n2608), .Z(n2554) );
  XOR U2628 ( .A(n2555), .B(n2554), .Z(n2513) );
  IV U2629 ( .A(n2513), .Z(n2556) );
  XOR U2630 ( .A(n2557), .B(n2556), .Z(n2615) );
  NOR U2631 ( .A(n110), .B(n149), .Z(n2613) );
  XOR U2632 ( .A(n2615), .B(n2613), .Z(n2616) );
  XOR U2633 ( .A(n2617), .B(n2616), .Z(n2547) );
  XOR U2634 ( .A(n2548), .B(n2547), .Z(n2549) );
  XOR U2635 ( .A(n2551), .B(n2549), .Z(n2539) );
  XOR U2636 ( .A(n2540), .B(n2539), .Z(n2541) );
  XOR U2637 ( .A(n2542), .B(n2541), .Z(n2533) );
  XOR U2638 ( .A(n2534), .B(n2533), .Z(n2514) );
  IV U2639 ( .A(n2514), .Z(n2535) );
  XOR U2640 ( .A(n2536), .B(n2535), .Z(n2626) );
  NOR U2641 ( .A(n2516), .B(n2515), .Z(n2520) );
  NOR U2642 ( .A(n2518), .B(n2517), .Z(n2519) );
  NOR U2643 ( .A(n2520), .B(n2519), .Z(n2624) );
  NOR U2644 ( .A(n112), .B(n140), .Z(n2622) );
  XOR U2645 ( .A(n2624), .B(n2622), .Z(n2625) );
  XOR U2646 ( .A(n2626), .B(n2625), .Z(n2527) );
  XOR U2647 ( .A(n2528), .B(n2527), .Z(n2521) );
  IV U2648 ( .A(n2521), .Z(n2529) );
  XOR U2649 ( .A(n2530), .B(n2529), .Z(n2958) );
  XOR U2650 ( .A(n2523), .B(n2522), .Z(n2957) );
  NOR U2651 ( .A(n2958), .B(n2957), .Z(n2524) );
  NOR U2652 ( .A(n2525), .B(n2524), .Z(n2631) );
  NOR U2653 ( .A(n83), .B(n136), .Z(n2630) );
  IV U2654 ( .A(n2630), .Z(n2526) );
  NOR U2655 ( .A(n2631), .B(n2526), .Z(n2633) );
  NOR U2656 ( .A(n2528), .B(n2527), .Z(n2532) );
  NOR U2657 ( .A(n2530), .B(n2529), .Z(n2531) );
  NOR U2658 ( .A(n2532), .B(n2531), .Z(n2638) );
  NOR U2659 ( .A(n113), .B(n138), .Z(n2636) );
  NOR U2660 ( .A(n2534), .B(n2533), .Z(n2538) );
  NOR U2661 ( .A(n2536), .B(n2535), .Z(n2537) );
  NOR U2662 ( .A(n2538), .B(n2537), .Z(n2651) );
  NOR U2663 ( .A(n112), .B(n142), .Z(n2649) );
  IV U2664 ( .A(n2649), .Z(n2621) );
  NOR U2665 ( .A(n2540), .B(n2539), .Z(n2545) );
  IV U2666 ( .A(n2541), .Z(n2543) );
  NOR U2667 ( .A(n2543), .B(n2542), .Z(n2544) );
  NOR U2668 ( .A(n2545), .B(n2544), .Z(n2546) );
  IV U2669 ( .A(n2546), .Z(n2658) );
  NOR U2670 ( .A(n2548), .B(n2547), .Z(n2553) );
  IV U2671 ( .A(n2549), .Z(n2550) );
  NOR U2672 ( .A(n2551), .B(n2550), .Z(n2552) );
  NOR U2673 ( .A(n2553), .B(n2552), .Z(n2664) );
  NOR U2674 ( .A(n111), .B(n146), .Z(n2662) );
  NOR U2675 ( .A(n2555), .B(n2554), .Z(n2559) );
  NOR U2676 ( .A(n2557), .B(n2556), .Z(n2558) );
  NOR U2677 ( .A(n2559), .B(n2558), .Z(n2670) );
  NOR U2678 ( .A(n110), .B(n151), .Z(n2668) );
  NOR U2679 ( .A(n2561), .B(n2560), .Z(n2565) );
  NOR U2680 ( .A(n2563), .B(n2562), .Z(n2564) );
  NOR U2681 ( .A(n2565), .B(n2564), .Z(n2683) );
  NOR U2682 ( .A(n108), .B(n154), .Z(n2681) );
  IV U2683 ( .A(n2681), .Z(n2604) );
  NOR U2684 ( .A(n2567), .B(n2566), .Z(n2572) );
  IV U2685 ( .A(n2568), .Z(n2570) );
  NOR U2686 ( .A(n2570), .B(n2569), .Z(n2571) );
  NOR U2687 ( .A(n2572), .B(n2571), .Z(n2573) );
  IV U2688 ( .A(n2573), .Z(n2688) );
  NOR U2689 ( .A(n87), .B(n157), .Z(n2686) );
  XOR U2690 ( .A(n2688), .B(n2686), .Z(n2689) );
  NOR U2691 ( .A(n2575), .B(n2574), .Z(n2580) );
  IV U2692 ( .A(n2576), .Z(n2577) );
  NOR U2693 ( .A(n2578), .B(n2577), .Z(n2579) );
  NOR U2694 ( .A(n2580), .B(n2579), .Z(n2696) );
  NOR U2695 ( .A(n107), .B(n159), .Z(n2694) );
  IV U2696 ( .A(n2694), .Z(n2603) );
  NOR U2697 ( .A(n2582), .B(n2581), .Z(n2586) );
  NOR U2698 ( .A(n2584), .B(n2583), .Z(n2585) );
  NOR U2699 ( .A(n2586), .B(n2585), .Z(n2709) );
  NOR U2700 ( .A(n106), .B(n162), .Z(n2707) );
  IV U2701 ( .A(n2707), .Z(n2595) );
  IV U2702 ( .A(n2587), .Z(n2588) );
  NOR U2703 ( .A(n2589), .B(n2588), .Z(n2593) );
  NOR U2704 ( .A(n2591), .B(n2590), .Z(n2592) );
  NOR U2705 ( .A(n2593), .B(n2592), .Z(n2714) );
  NOR U2706 ( .A(n164), .B(n105), .Z(n2712) );
  XOR U2707 ( .A(n2714), .B(n2712), .Z(n2716) );
  NOR U2708 ( .A(n166), .B(n104), .Z(n2594) );
  IV U2709 ( .A(n2594), .Z(n2715) );
  XOR U2710 ( .A(n2716), .B(n2715), .Z(n2706) );
  XOR U2711 ( .A(n2595), .B(n2706), .Z(n2708) );
  XOR U2712 ( .A(n2709), .B(n2708), .Z(n2703) );
  IV U2713 ( .A(n2596), .Z(n2597) );
  NOR U2714 ( .A(n2598), .B(n2597), .Z(n2602) );
  NOR U2715 ( .A(n2600), .B(n2599), .Z(n2601) );
  NOR U2716 ( .A(n2602), .B(n2601), .Z(n2701) );
  NOR U2717 ( .A(n88), .B(n160), .Z(n2699) );
  XOR U2718 ( .A(n2701), .B(n2699), .Z(n2702) );
  XOR U2719 ( .A(n2703), .B(n2702), .Z(n2693) );
  XOR U2720 ( .A(n2603), .B(n2693), .Z(n2695) );
  XOR U2721 ( .A(n2696), .B(n2695), .Z(n2690) );
  XOR U2722 ( .A(n2689), .B(n2690), .Z(n2680) );
  XOR U2723 ( .A(n2604), .B(n2680), .Z(n2682) );
  XOR U2724 ( .A(n2683), .B(n2682), .Z(n2677) );
  IV U2725 ( .A(n2605), .Z(n2606) );
  NOR U2726 ( .A(n2607), .B(n2606), .Z(n2611) );
  NOR U2727 ( .A(n2609), .B(n2608), .Z(n2610) );
  NOR U2728 ( .A(n2611), .B(n2610), .Z(n2675) );
  NOR U2729 ( .A(n109), .B(n152), .Z(n2673) );
  XOR U2730 ( .A(n2675), .B(n2673), .Z(n2676) );
  XOR U2731 ( .A(n2677), .B(n2676), .Z(n2667) );
  XOR U2732 ( .A(n2668), .B(n2667), .Z(n2612) );
  IV U2733 ( .A(n2612), .Z(n2669) );
  XOR U2734 ( .A(n2670), .B(n2669), .Z(n2732) );
  IV U2735 ( .A(n2613), .Z(n2614) );
  NOR U2736 ( .A(n2615), .B(n2614), .Z(n2619) );
  NOR U2737 ( .A(n2617), .B(n2616), .Z(n2618) );
  NOR U2738 ( .A(n2619), .B(n2618), .Z(n2730) );
  NOR U2739 ( .A(n86), .B(n149), .Z(n2728) );
  XOR U2740 ( .A(n2730), .B(n2728), .Z(n2731) );
  XOR U2741 ( .A(n2732), .B(n2731), .Z(n2661) );
  XOR U2742 ( .A(n2662), .B(n2661), .Z(n2620) );
  IV U2743 ( .A(n2620), .Z(n2663) );
  XOR U2744 ( .A(n2664), .B(n2663), .Z(n2656) );
  NOR U2745 ( .A(n85), .B(n144), .Z(n2654) );
  XOR U2746 ( .A(n2656), .B(n2654), .Z(n2657) );
  XOR U2747 ( .A(n2658), .B(n2657), .Z(n2648) );
  XOR U2748 ( .A(n2621), .B(n2648), .Z(n2650) );
  XOR U2749 ( .A(n2651), .B(n2650), .Z(n2645) );
  IV U2750 ( .A(n2622), .Z(n2623) );
  NOR U2751 ( .A(n2624), .B(n2623), .Z(n2628) );
  NOR U2752 ( .A(n2626), .B(n2625), .Z(n2627) );
  NOR U2753 ( .A(n2628), .B(n2627), .Z(n2643) );
  NOR U2754 ( .A(n84), .B(n140), .Z(n2641) );
  XOR U2755 ( .A(n2643), .B(n2641), .Z(n2644) );
  XOR U2756 ( .A(n2645), .B(n2644), .Z(n2635) );
  XOR U2757 ( .A(n2636), .B(n2635), .Z(n2629) );
  IV U2758 ( .A(n2629), .Z(n2637) );
  XOR U2759 ( .A(n2638), .B(n2637), .Z(n2956) );
  XOR U2760 ( .A(n2631), .B(n2630), .Z(n2955) );
  NOR U2761 ( .A(n2956), .B(n2955), .Z(n2632) );
  NOR U2762 ( .A(n2633), .B(n2632), .Z(n2739) );
  NOR U2763 ( .A(n114), .B(n136), .Z(n2738) );
  IV U2764 ( .A(n2738), .Z(n2634) );
  NOR U2765 ( .A(n2739), .B(n2634), .Z(n2741) );
  NOR U2766 ( .A(n2636), .B(n2635), .Z(n2640) );
  NOR U2767 ( .A(n2638), .B(n2637), .Z(n2639) );
  NOR U2768 ( .A(n2640), .B(n2639), .Z(n2746) );
  NOR U2769 ( .A(n83), .B(n138), .Z(n2744) );
  IV U2770 ( .A(n2641), .Z(n2642) );
  NOR U2771 ( .A(n2643), .B(n2642), .Z(n2647) );
  NOR U2772 ( .A(n2645), .B(n2644), .Z(n2646) );
  NOR U2773 ( .A(n2647), .B(n2646), .Z(n2834) );
  NOR U2774 ( .A(n2649), .B(n2648), .Z(n2653) );
  NOR U2775 ( .A(n2651), .B(n2650), .Z(n2652) );
  NOR U2776 ( .A(n2653), .B(n2652), .Z(n2752) );
  NOR U2777 ( .A(n84), .B(n142), .Z(n2750) );
  IV U2778 ( .A(n2654), .Z(n2655) );
  NOR U2779 ( .A(n2656), .B(n2655), .Z(n2660) );
  NOR U2780 ( .A(n2658), .B(n2657), .Z(n2659) );
  NOR U2781 ( .A(n2660), .B(n2659), .Z(n2826) );
  NOR U2782 ( .A(n2662), .B(n2661), .Z(n2666) );
  NOR U2783 ( .A(n2664), .B(n2663), .Z(n2665) );
  NOR U2784 ( .A(n2666), .B(n2665), .Z(n2758) );
  NOR U2785 ( .A(n85), .B(n146), .Z(n2756) );
  NOR U2786 ( .A(n2668), .B(n2667), .Z(n2672) );
  NOR U2787 ( .A(n2670), .B(n2669), .Z(n2671) );
  NOR U2788 ( .A(n2672), .B(n2671), .Z(n2764) );
  NOR U2789 ( .A(n86), .B(n151), .Z(n2762) );
  IV U2790 ( .A(n2673), .Z(n2674) );
  NOR U2791 ( .A(n2675), .B(n2674), .Z(n2679) );
  NOR U2792 ( .A(n2677), .B(n2676), .Z(n2678) );
  NOR U2793 ( .A(n2679), .B(n2678), .Z(n2771) );
  NOR U2794 ( .A(n2681), .B(n2680), .Z(n2685) );
  NOR U2795 ( .A(n2683), .B(n2682), .Z(n2684) );
  NOR U2796 ( .A(n2685), .B(n2684), .Z(n2777) );
  NOR U2797 ( .A(n109), .B(n154), .Z(n2775) );
  IV U2798 ( .A(n2775), .Z(n2726) );
  IV U2799 ( .A(n2686), .Z(n2687) );
  NOR U2800 ( .A(n2688), .B(n2687), .Z(n2692) );
  NOR U2801 ( .A(n2690), .B(n2689), .Z(n2691) );
  NOR U2802 ( .A(n2692), .B(n2691), .Z(n2780) );
  IV U2803 ( .A(n2780), .Z(n2724) );
  NOR U2804 ( .A(n2694), .B(n2693), .Z(n2698) );
  NOR U2805 ( .A(n2696), .B(n2695), .Z(n2697) );
  NOR U2806 ( .A(n2698), .B(n2697), .Z(n2789) );
  NOR U2807 ( .A(n87), .B(n159), .Z(n2787) );
  IV U2808 ( .A(n2787), .Z(n2723) );
  IV U2809 ( .A(n2699), .Z(n2700) );
  NOR U2810 ( .A(n2701), .B(n2700), .Z(n2705) );
  NOR U2811 ( .A(n2703), .B(n2702), .Z(n2704) );
  NOR U2812 ( .A(n2705), .B(n2704), .Z(n2792) );
  IV U2813 ( .A(n2792), .Z(n2721) );
  NOR U2814 ( .A(n2707), .B(n2706), .Z(n2711) );
  NOR U2815 ( .A(n2709), .B(n2708), .Z(n2710) );
  NOR U2816 ( .A(n2711), .B(n2710), .Z(n2801) );
  NOR U2817 ( .A(n88), .B(n162), .Z(n2799) );
  IV U2818 ( .A(n2799), .Z(n2720) );
  IV U2819 ( .A(n2712), .Z(n2713) );
  NOR U2820 ( .A(n2714), .B(n2713), .Z(n2718) );
  NOR U2821 ( .A(n2716), .B(n2715), .Z(n2717) );
  NOR U2822 ( .A(n2718), .B(n2717), .Z(n2806) );
  NOR U2823 ( .A(n164), .B(n106), .Z(n2804) );
  XOR U2824 ( .A(n2806), .B(n2804), .Z(n2808) );
  NOR U2825 ( .A(n166), .B(n105), .Z(n2719) );
  IV U2826 ( .A(n2719), .Z(n2807) );
  XOR U2827 ( .A(n2808), .B(n2807), .Z(n2798) );
  XOR U2828 ( .A(n2720), .B(n2798), .Z(n2800) );
  XOR U2829 ( .A(n2801), .B(n2800), .Z(n2793) );
  XOR U2830 ( .A(n2721), .B(n2793), .Z(n2795) );
  NOR U2831 ( .A(n107), .B(n160), .Z(n2722) );
  IV U2832 ( .A(n2722), .Z(n2794) );
  XOR U2833 ( .A(n2795), .B(n2794), .Z(n2786) );
  XOR U2834 ( .A(n2723), .B(n2786), .Z(n2788) );
  XOR U2835 ( .A(n2789), .B(n2788), .Z(n2781) );
  XOR U2836 ( .A(n2724), .B(n2781), .Z(n2783) );
  NOR U2837 ( .A(n108), .B(n157), .Z(n2725) );
  IV U2838 ( .A(n2725), .Z(n2782) );
  XOR U2839 ( .A(n2783), .B(n2782), .Z(n2774) );
  XOR U2840 ( .A(n2726), .B(n2774), .Z(n2776) );
  XOR U2841 ( .A(n2777), .B(n2776), .Z(n2769) );
  NOR U2842 ( .A(n110), .B(n152), .Z(n2767) );
  XOR U2843 ( .A(n2769), .B(n2767), .Z(n2770) );
  XOR U2844 ( .A(n2771), .B(n2770), .Z(n2761) );
  XOR U2845 ( .A(n2762), .B(n2761), .Z(n2727) );
  IV U2846 ( .A(n2727), .Z(n2763) );
  XOR U2847 ( .A(n2764), .B(n2763), .Z(n2818) );
  IV U2848 ( .A(n2728), .Z(n2729) );
  NOR U2849 ( .A(n2730), .B(n2729), .Z(n2734) );
  NOR U2850 ( .A(n2732), .B(n2731), .Z(n2733) );
  NOR U2851 ( .A(n2734), .B(n2733), .Z(n2816) );
  NOR U2852 ( .A(n111), .B(n149), .Z(n2814) );
  XOR U2853 ( .A(n2816), .B(n2814), .Z(n2817) );
  XOR U2854 ( .A(n2818), .B(n2817), .Z(n2755) );
  XOR U2855 ( .A(n2756), .B(n2755), .Z(n2735) );
  IV U2856 ( .A(n2735), .Z(n2757) );
  XOR U2857 ( .A(n2758), .B(n2757), .Z(n2824) );
  NOR U2858 ( .A(n112), .B(n144), .Z(n2822) );
  XOR U2859 ( .A(n2824), .B(n2822), .Z(n2825) );
  XOR U2860 ( .A(n2826), .B(n2825), .Z(n2749) );
  XOR U2861 ( .A(n2750), .B(n2749), .Z(n2736) );
  IV U2862 ( .A(n2736), .Z(n2751) );
  XOR U2863 ( .A(n2752), .B(n2751), .Z(n2832) );
  NOR U2864 ( .A(n113), .B(n140), .Z(n2830) );
  XOR U2865 ( .A(n2832), .B(n2830), .Z(n2833) );
  XOR U2866 ( .A(n2834), .B(n2833), .Z(n2743) );
  XOR U2867 ( .A(n2744), .B(n2743), .Z(n2737) );
  IV U2868 ( .A(n2737), .Z(n2745) );
  XOR U2869 ( .A(n2746), .B(n2745), .Z(n2954) );
  XOR U2870 ( .A(n2739), .B(n2738), .Z(n2953) );
  NOR U2871 ( .A(n2954), .B(n2953), .Z(n2740) );
  NOR U2872 ( .A(n2741), .B(n2740), .Z(n2839) );
  NOR U2873 ( .A(n82), .B(n136), .Z(n2838) );
  IV U2874 ( .A(n2838), .Z(n2742) );
  NOR U2875 ( .A(n2839), .B(n2742), .Z(n2841) );
  NOR U2876 ( .A(n2744), .B(n2743), .Z(n2748) );
  NOR U2877 ( .A(n2746), .B(n2745), .Z(n2747) );
  NOR U2878 ( .A(n2748), .B(n2747), .Z(n2845) );
  NOR U2879 ( .A(n114), .B(n138), .Z(n2843) );
  NOR U2880 ( .A(n2750), .B(n2749), .Z(n2754) );
  NOR U2881 ( .A(n2752), .B(n2751), .Z(n2753) );
  NOR U2882 ( .A(n2754), .B(n2753), .Z(n2858) );
  NOR U2883 ( .A(n113), .B(n142), .Z(n2856) );
  NOR U2884 ( .A(n2756), .B(n2755), .Z(n2760) );
  NOR U2885 ( .A(n2758), .B(n2757), .Z(n2759) );
  NOR U2886 ( .A(n2760), .B(n2759), .Z(n2871) );
  NOR U2887 ( .A(n112), .B(n146), .Z(n2869) );
  NOR U2888 ( .A(n2762), .B(n2761), .Z(n2766) );
  NOR U2889 ( .A(n2764), .B(n2763), .Z(n2765) );
  NOR U2890 ( .A(n2766), .B(n2765), .Z(n2878) );
  NOR U2891 ( .A(n111), .B(n151), .Z(n2876) );
  NOR U2892 ( .A(n86), .B(n152), .Z(n2885) );
  IV U2893 ( .A(n2767), .Z(n2768) );
  NOR U2894 ( .A(n2769), .B(n2768), .Z(n2773) );
  NOR U2895 ( .A(n2771), .B(n2770), .Z(n2772) );
  NOR U2896 ( .A(n2773), .B(n2772), .Z(n2881) );
  NOR U2897 ( .A(n2775), .B(n2774), .Z(n2779) );
  NOR U2898 ( .A(n2777), .B(n2776), .Z(n2778) );
  NOR U2899 ( .A(n2779), .B(n2778), .Z(n2893) );
  NOR U2900 ( .A(n110), .B(n154), .Z(n2890) );
  NOR U2901 ( .A(n2781), .B(n2780), .Z(n2785) );
  NOR U2902 ( .A(n2783), .B(n2782), .Z(n2784) );
  NOR U2903 ( .A(n2785), .B(n2784), .Z(n2896) );
  NOR U2904 ( .A(n2787), .B(n2786), .Z(n2791) );
  NOR U2905 ( .A(n2789), .B(n2788), .Z(n2790) );
  NOR U2906 ( .A(n2791), .B(n2790), .Z(n2907) );
  NOR U2907 ( .A(n108), .B(n159), .Z(n2905) );
  IV U2908 ( .A(n2905), .Z(n2813) );
  NOR U2909 ( .A(n2793), .B(n2792), .Z(n2797) );
  NOR U2910 ( .A(n2795), .B(n2794), .Z(n2796) );
  NOR U2911 ( .A(n2797), .B(n2796), .Z(n2914) );
  NOR U2912 ( .A(n2799), .B(n2798), .Z(n2803) );
  NOR U2913 ( .A(n2801), .B(n2800), .Z(n2802) );
  NOR U2914 ( .A(n2803), .B(n2802), .Z(n2920) );
  NOR U2915 ( .A(n107), .B(n162), .Z(n2918) );
  IV U2916 ( .A(n2918), .Z(n2812) );
  IV U2917 ( .A(n2804), .Z(n2805) );
  NOR U2918 ( .A(n2806), .B(n2805), .Z(n2810) );
  NOR U2919 ( .A(n2808), .B(n2807), .Z(n2809) );
  NOR U2920 ( .A(n2810), .B(n2809), .Z(n2925) );
  NOR U2921 ( .A(n164), .B(n88), .Z(n2923) );
  XOR U2922 ( .A(n2925), .B(n2923), .Z(n2927) );
  NOR U2923 ( .A(n166), .B(n106), .Z(n2811) );
  IV U2924 ( .A(n2811), .Z(n2926) );
  XOR U2925 ( .A(n2927), .B(n2926), .Z(n2917) );
  XOR U2926 ( .A(n2812), .B(n2917), .Z(n2919) );
  XOR U2927 ( .A(n2920), .B(n2919), .Z(n2912) );
  NOR U2928 ( .A(n87), .B(n160), .Z(n2910) );
  XOR U2929 ( .A(n2912), .B(n2910), .Z(n2913) );
  XOR U2930 ( .A(n2914), .B(n2913), .Z(n2904) );
  XOR U2931 ( .A(n2813), .B(n2904), .Z(n2906) );
  XOR U2932 ( .A(n2907), .B(n2906), .Z(n2897) );
  XOR U2933 ( .A(n2896), .B(n2897), .Z(n2898) );
  NOR U2934 ( .A(n109), .B(n157), .Z(n2899) );
  XOR U2935 ( .A(n2898), .B(n2899), .Z(n2889) );
  XOR U2936 ( .A(n2890), .B(n2889), .Z(n2891) );
  XOR U2937 ( .A(n2893), .B(n2891), .Z(n2882) );
  XOR U2938 ( .A(n2881), .B(n2882), .Z(n2884) );
  XOR U2939 ( .A(n2885), .B(n2884), .Z(n2874) );
  XOR U2940 ( .A(n2876), .B(n2874), .Z(n2877) );
  XOR U2941 ( .A(n2878), .B(n2877), .Z(n2941) );
  IV U2942 ( .A(n2814), .Z(n2815) );
  NOR U2943 ( .A(n2816), .B(n2815), .Z(n2820) );
  NOR U2944 ( .A(n2818), .B(n2817), .Z(n2819) );
  NOR U2945 ( .A(n2820), .B(n2819), .Z(n2939) );
  NOR U2946 ( .A(n85), .B(n149), .Z(n2937) );
  XOR U2947 ( .A(n2939), .B(n2937), .Z(n2940) );
  XOR U2948 ( .A(n2941), .B(n2940), .Z(n2868) );
  XOR U2949 ( .A(n2869), .B(n2868), .Z(n2821) );
  IV U2950 ( .A(n2821), .Z(n2870) );
  XOR U2951 ( .A(n2871), .B(n2870), .Z(n2865) );
  IV U2952 ( .A(n2822), .Z(n2823) );
  NOR U2953 ( .A(n2824), .B(n2823), .Z(n2828) );
  NOR U2954 ( .A(n2826), .B(n2825), .Z(n2827) );
  NOR U2955 ( .A(n2828), .B(n2827), .Z(n2863) );
  NOR U2956 ( .A(n84), .B(n144), .Z(n2861) );
  XOR U2957 ( .A(n2863), .B(n2861), .Z(n2864) );
  XOR U2958 ( .A(n2865), .B(n2864), .Z(n2855) );
  XOR U2959 ( .A(n2856), .B(n2855), .Z(n2829) );
  IV U2960 ( .A(n2829), .Z(n2857) );
  XOR U2961 ( .A(n2858), .B(n2857), .Z(n2852) );
  IV U2962 ( .A(n2830), .Z(n2831) );
  NOR U2963 ( .A(n2832), .B(n2831), .Z(n2836) );
  NOR U2964 ( .A(n2834), .B(n2833), .Z(n2835) );
  NOR U2965 ( .A(n2836), .B(n2835), .Z(n2850) );
  NOR U2966 ( .A(n83), .B(n140), .Z(n2848) );
  XOR U2967 ( .A(n2850), .B(n2848), .Z(n2851) );
  XOR U2968 ( .A(n2852), .B(n2851), .Z(n2842) );
  XOR U2969 ( .A(n2843), .B(n2842), .Z(n2837) );
  IV U2970 ( .A(n2837), .Z(n2844) );
  XOR U2971 ( .A(n2845), .B(n2844), .Z(n2952) );
  XOR U2972 ( .A(n2839), .B(n2838), .Z(n2951) );
  NOR U2973 ( .A(n2952), .B(n2951), .Z(n2840) );
  NOR U2974 ( .A(n2841), .B(n2840), .Z(n3306) );
  IV U2975 ( .A(n3306), .Z(n2949) );
  NOR U2976 ( .A(n2843), .B(n2842), .Z(n2847) );
  NOR U2977 ( .A(n2845), .B(n2844), .Z(n2846) );
  NOR U2978 ( .A(n2847), .B(n2846), .Z(n3208) );
  NOR U2979 ( .A(n82), .B(n138), .Z(n3206) );
  IV U2980 ( .A(n3206), .Z(n2948) );
  IV U2981 ( .A(n2848), .Z(n2849) );
  NOR U2982 ( .A(n2850), .B(n2849), .Z(n2854) );
  NOR U2983 ( .A(n2852), .B(n2851), .Z(n2853) );
  NOR U2984 ( .A(n2854), .B(n2853), .Z(n3302) );
  NOR U2985 ( .A(n2856), .B(n2855), .Z(n2860) );
  NOR U2986 ( .A(n2858), .B(n2857), .Z(n2859) );
  NOR U2987 ( .A(n2860), .B(n2859), .Z(n3214) );
  NOR U2988 ( .A(n83), .B(n142), .Z(n3212) );
  IV U2989 ( .A(n3212), .Z(n2947) );
  IV U2990 ( .A(n2861), .Z(n2862) );
  NOR U2991 ( .A(n2863), .B(n2862), .Z(n2867) );
  NOR U2992 ( .A(n2865), .B(n2864), .Z(n2866) );
  NOR U2993 ( .A(n2867), .B(n2866), .Z(n3217) );
  IV U2994 ( .A(n3217), .Z(n2945) );
  NOR U2995 ( .A(n2869), .B(n2868), .Z(n2873) );
  NOR U2996 ( .A(n2871), .B(n2870), .Z(n2872) );
  NOR U2997 ( .A(n2873), .B(n2872), .Z(n3226) );
  NOR U2998 ( .A(n84), .B(n146), .Z(n3224) );
  IV U2999 ( .A(n3224), .Z(n2944) );
  IV U3000 ( .A(n2874), .Z(n2875) );
  NOR U3001 ( .A(n2876), .B(n2875), .Z(n2880) );
  NOR U3002 ( .A(n2878), .B(n2877), .Z(n2879) );
  NOR U3003 ( .A(n2880), .B(n2879), .Z(n3239) );
  NOR U3004 ( .A(n85), .B(n151), .Z(n3237) );
  IV U3005 ( .A(n3237), .Z(n2936) );
  IV U3006 ( .A(n2881), .Z(n2883) );
  NOR U3007 ( .A(n2883), .B(n2882), .Z(n2887) );
  NOR U3008 ( .A(n2885), .B(n2884), .Z(n2886) );
  NOR U3009 ( .A(n2887), .B(n2886), .Z(n2888) );
  IV U3010 ( .A(n2888), .Z(n3288) );
  NOR U3011 ( .A(n2890), .B(n2889), .Z(n2895) );
  IV U3012 ( .A(n2891), .Z(n2892) );
  NOR U3013 ( .A(n2893), .B(n2892), .Z(n2894) );
  NOR U3014 ( .A(n2895), .B(n2894), .Z(n3245) );
  NOR U3015 ( .A(n86), .B(n154), .Z(n3243) );
  NOR U3016 ( .A(n2897), .B(n2896), .Z(n2903) );
  IV U3017 ( .A(n2898), .Z(n2901) );
  IV U3018 ( .A(n2899), .Z(n2900) );
  NOR U3019 ( .A(n2901), .B(n2900), .Z(n2902) );
  NOR U3020 ( .A(n2903), .B(n2902), .Z(n3280) );
  NOR U3021 ( .A(n2905), .B(n2904), .Z(n2909) );
  NOR U3022 ( .A(n2907), .B(n2906), .Z(n2908) );
  NOR U3023 ( .A(n2909), .B(n2908), .Z(n3251) );
  NOR U3024 ( .A(n109), .B(n159), .Z(n3249) );
  IV U3025 ( .A(n3249), .Z(n2934) );
  IV U3026 ( .A(n2910), .Z(n2911) );
  NOR U3027 ( .A(n2912), .B(n2911), .Z(n2916) );
  NOR U3028 ( .A(n2914), .B(n2913), .Z(n2915) );
  NOR U3029 ( .A(n2916), .B(n2915), .Z(n3254) );
  IV U3030 ( .A(n3254), .Z(n2932) );
  NOR U3031 ( .A(n2918), .B(n2917), .Z(n2922) );
  NOR U3032 ( .A(n2920), .B(n2919), .Z(n2921) );
  NOR U3033 ( .A(n2922), .B(n2921), .Z(n3263) );
  NOR U3034 ( .A(n87), .B(n162), .Z(n3261) );
  IV U3035 ( .A(n3261), .Z(n2931) );
  IV U3036 ( .A(n2923), .Z(n2924) );
  NOR U3037 ( .A(n2925), .B(n2924), .Z(n2929) );
  NOR U3038 ( .A(n2927), .B(n2926), .Z(n2928) );
  NOR U3039 ( .A(n2929), .B(n2928), .Z(n3268) );
  NOR U3040 ( .A(n164), .B(n107), .Z(n3266) );
  XOR U3041 ( .A(n3268), .B(n3266), .Z(n3270) );
  NOR U3042 ( .A(n166), .B(n88), .Z(n2930) );
  IV U3043 ( .A(n2930), .Z(n3269) );
  XOR U3044 ( .A(n3270), .B(n3269), .Z(n3260) );
  XOR U3045 ( .A(n2931), .B(n3260), .Z(n3262) );
  XOR U3046 ( .A(n3263), .B(n3262), .Z(n3255) );
  XOR U3047 ( .A(n2932), .B(n3255), .Z(n3257) );
  NOR U3048 ( .A(n108), .B(n160), .Z(n2933) );
  IV U3049 ( .A(n2933), .Z(n3256) );
  XOR U3050 ( .A(n3257), .B(n3256), .Z(n3248) );
  XOR U3051 ( .A(n2934), .B(n3248), .Z(n3250) );
  XOR U3052 ( .A(n3251), .B(n3250), .Z(n3278) );
  NOR U3053 ( .A(n110), .B(n157), .Z(n3276) );
  XOR U3054 ( .A(n3278), .B(n3276), .Z(n3279) );
  XOR U3055 ( .A(n3280), .B(n3279), .Z(n3242) );
  XOR U3056 ( .A(n3243), .B(n3242), .Z(n2935) );
  IV U3057 ( .A(n2935), .Z(n3244) );
  XOR U3058 ( .A(n3245), .B(n3244), .Z(n3286) );
  NOR U3059 ( .A(n111), .B(n152), .Z(n3284) );
  XOR U3060 ( .A(n3286), .B(n3284), .Z(n3287) );
  XOR U3061 ( .A(n3288), .B(n3287), .Z(n3236) );
  XOR U3062 ( .A(n2936), .B(n3236), .Z(n3238) );
  XOR U3063 ( .A(n3239), .B(n3238), .Z(n3233) );
  IV U3064 ( .A(n2937), .Z(n2938) );
  NOR U3065 ( .A(n2939), .B(n2938), .Z(n2943) );
  NOR U3066 ( .A(n2941), .B(n2940), .Z(n2942) );
  NOR U3067 ( .A(n2943), .B(n2942), .Z(n3231) );
  NOR U3068 ( .A(n112), .B(n149), .Z(n3229) );
  XOR U3069 ( .A(n3231), .B(n3229), .Z(n3232) );
  XOR U3070 ( .A(n3233), .B(n3232), .Z(n3223) );
  XOR U3071 ( .A(n2944), .B(n3223), .Z(n3225) );
  XOR U3072 ( .A(n3226), .B(n3225), .Z(n3218) );
  XOR U3073 ( .A(n2945), .B(n3218), .Z(n3220) );
  NOR U3074 ( .A(n113), .B(n144), .Z(n2946) );
  IV U3075 ( .A(n2946), .Z(n3219) );
  XOR U3076 ( .A(n3220), .B(n3219), .Z(n3211) );
  XOR U3077 ( .A(n2947), .B(n3211), .Z(n3213) );
  XOR U3078 ( .A(n3214), .B(n3213), .Z(n3300) );
  NOR U3079 ( .A(n114), .B(n140), .Z(n3298) );
  XOR U3080 ( .A(n3300), .B(n3298), .Z(n3301) );
  XOR U3081 ( .A(n3302), .B(n3301), .Z(n3205) );
  XOR U3082 ( .A(n2948), .B(n3205), .Z(n3207) );
  XOR U3083 ( .A(n3208), .B(n3207), .Z(n3307) );
  XOR U3084 ( .A(n2949), .B(n3307), .Z(n3309) );
  NOR U3085 ( .A(n115), .B(n136), .Z(n2950) );
  IV U3086 ( .A(n2950), .Z(n3308) );
  XOR U3087 ( .A(n3309), .B(n3308), .Z(n3201) );
  NOR U3088 ( .A(n3200), .B(n3201), .Z(n3204) );
  NOR U3089 ( .A(n115), .B(n134), .Z(n3196) );
  XOR U3090 ( .A(n2952), .B(n2951), .Z(n3195) );
  NOR U3091 ( .A(n3196), .B(n3195), .Z(n3199) );
  NOR U3092 ( .A(n82), .B(n134), .Z(n3191) );
  XOR U3093 ( .A(n2954), .B(n2953), .Z(n3190) );
  NOR U3094 ( .A(n3191), .B(n3190), .Z(n3194) );
  NOR U3095 ( .A(n114), .B(n134), .Z(n3186) );
  XOR U3096 ( .A(n2956), .B(n2955), .Z(n3185) );
  NOR U3097 ( .A(n3186), .B(n3185), .Z(n3189) );
  NOR U3098 ( .A(n83), .B(n134), .Z(n3181) );
  XOR U3099 ( .A(n2958), .B(n2957), .Z(n3180) );
  NOR U3100 ( .A(n3181), .B(n3180), .Z(n3184) );
  NOR U3101 ( .A(n113), .B(n134), .Z(n3176) );
  XOR U3102 ( .A(n2960), .B(n2959), .Z(n3175) );
  NOR U3103 ( .A(n3176), .B(n3175), .Z(n3179) );
  XOR U3104 ( .A(n2962), .B(n2961), .Z(n3171) );
  NOR U3105 ( .A(n84), .B(n134), .Z(n3170) );
  IV U3106 ( .A(n3170), .Z(n2963) );
  NOR U3107 ( .A(n3171), .B(n2963), .Z(n3173) );
  XOR U3108 ( .A(n2965), .B(n2964), .Z(n3166) );
  NOR U3109 ( .A(n112), .B(n134), .Z(n3167) );
  IV U3110 ( .A(n3167), .Z(n2966) );
  NOR U3111 ( .A(n3166), .B(n2966), .Z(n3169) );
  XOR U3112 ( .A(n2968), .B(n2967), .Z(n3162) );
  NOR U3113 ( .A(n85), .B(n134), .Z(n3163) );
  IV U3114 ( .A(n3163), .Z(n2969) );
  NOR U3115 ( .A(n3162), .B(n2969), .Z(n3165) );
  XOR U3116 ( .A(n2971), .B(n2970), .Z(n2974) );
  NOR U3117 ( .A(n111), .B(n134), .Z(n2973) );
  IV U3118 ( .A(n2973), .Z(n2972) );
  NOR U3119 ( .A(n2974), .B(n2972), .Z(n3161) );
  XOR U3120 ( .A(n2974), .B(n2973), .Z(n3519) );
  NOR U3121 ( .A(n86), .B(n134), .Z(n3154) );
  XOR U3122 ( .A(n2976), .B(n2975), .Z(n3155) );
  NOR U3123 ( .A(n3154), .B(n3155), .Z(n3158) );
  NOR U3124 ( .A(n110), .B(n134), .Z(n3150) );
  XOR U3125 ( .A(n2978), .B(n2977), .Z(n3149) );
  NOR U3126 ( .A(n3150), .B(n3149), .Z(n3153) );
  NOR U3127 ( .A(n109), .B(n134), .Z(n3145) );
  XOR U3128 ( .A(n2980), .B(n2979), .Z(n3144) );
  NOR U3129 ( .A(n3145), .B(n3144), .Z(n3148) );
  NOR U3130 ( .A(n108), .B(n134), .Z(n3140) );
  XOR U3131 ( .A(n2982), .B(n2981), .Z(n3139) );
  NOR U3132 ( .A(n3140), .B(n3139), .Z(n3143) );
  IV U3133 ( .A(n2983), .Z(n2985) );
  XOR U3134 ( .A(n2985), .B(n2984), .Z(n3134) );
  NOR U3135 ( .A(n87), .B(n134), .Z(n3135) );
  IV U3136 ( .A(n3135), .Z(n2986) );
  NOR U3137 ( .A(n3134), .B(n2986), .Z(n3137) );
  XOR U3138 ( .A(n2988), .B(n2987), .Z(n3130) );
  IV U3139 ( .A(n3130), .Z(n2990) );
  NOR U3140 ( .A(n107), .B(n134), .Z(n2989) );
  IV U3141 ( .A(n2989), .Z(n3131) );
  NOR U3142 ( .A(n2990), .B(n3131), .Z(n3133) );
  IV U3143 ( .A(n2991), .Z(n2993) );
  XOR U3144 ( .A(n2993), .B(n2992), .Z(n3126) );
  NOR U3145 ( .A(n88), .B(n134), .Z(n3127) );
  IV U3146 ( .A(n3127), .Z(n2994) );
  NOR U3147 ( .A(n3126), .B(n2994), .Z(n3129) );
  XOR U3148 ( .A(n2996), .B(n2995), .Z(n2997) );
  IV U3149 ( .A(n2997), .Z(n3122) );
  NOR U3150 ( .A(n106), .B(n134), .Z(n3123) );
  IV U3151 ( .A(n3123), .Z(n2998) );
  NOR U3152 ( .A(n3122), .B(n2998), .Z(n3125) );
  XOR U3153 ( .A(n3000), .B(n2999), .Z(n3001) );
  IV U3154 ( .A(n3001), .Z(n3118) );
  NOR U3155 ( .A(n105), .B(n134), .Z(n3119) );
  IV U3156 ( .A(n3119), .Z(n3002) );
  NOR U3157 ( .A(n3118), .B(n3002), .Z(n3121) );
  XOR U3158 ( .A(n3004), .B(n3003), .Z(n3005) );
  IV U3159 ( .A(n3005), .Z(n3114) );
  NOR U3160 ( .A(n104), .B(n134), .Z(n3115) );
  IV U3161 ( .A(n3115), .Z(n3006) );
  NOR U3162 ( .A(n3114), .B(n3006), .Z(n3117) );
  XOR U3163 ( .A(n3008), .B(n3007), .Z(n3009) );
  IV U3164 ( .A(n3009), .Z(n3110) );
  NOR U3165 ( .A(n89), .B(n134), .Z(n3111) );
  IV U3166 ( .A(n3111), .Z(n3010) );
  NOR U3167 ( .A(n3110), .B(n3010), .Z(n3113) );
  XOR U3168 ( .A(n3012), .B(n3011), .Z(n3013) );
  IV U3169 ( .A(n3013), .Z(n3106) );
  NOR U3170 ( .A(n103), .B(n134), .Z(n3107) );
  IV U3171 ( .A(n3107), .Z(n3014) );
  NOR U3172 ( .A(n3106), .B(n3014), .Z(n3109) );
  XOR U3173 ( .A(n3016), .B(n3015), .Z(n3017) );
  IV U3174 ( .A(n3017), .Z(n3102) );
  NOR U3175 ( .A(n90), .B(n134), .Z(n3103) );
  IV U3176 ( .A(n3103), .Z(n3018) );
  NOR U3177 ( .A(n3102), .B(n3018), .Z(n3105) );
  XOR U3178 ( .A(n3020), .B(n3019), .Z(n3021) );
  IV U3179 ( .A(n3021), .Z(n3098) );
  NOR U3180 ( .A(n102), .B(n134), .Z(n3099) );
  IV U3181 ( .A(n3099), .Z(n3022) );
  NOR U3182 ( .A(n3098), .B(n3022), .Z(n3101) );
  XOR U3183 ( .A(n3024), .B(n3023), .Z(n3025) );
  IV U3184 ( .A(n3025), .Z(n3094) );
  NOR U3185 ( .A(n101), .B(n134), .Z(n3095) );
  IV U3186 ( .A(n3095), .Z(n3026) );
  NOR U3187 ( .A(n3094), .B(n3026), .Z(n3097) );
  XOR U3188 ( .A(n3028), .B(n3027), .Z(n3029) );
  IV U3189 ( .A(n3029), .Z(n3090) );
  NOR U3190 ( .A(n100), .B(n134), .Z(n3091) );
  IV U3191 ( .A(n3091), .Z(n3030) );
  NOR U3192 ( .A(n3090), .B(n3030), .Z(n3093) );
  XOR U3193 ( .A(n3032), .B(n3031), .Z(n3033) );
  IV U3194 ( .A(n3033), .Z(n3086) );
  NOR U3195 ( .A(n99), .B(n134), .Z(n3087) );
  IV U3196 ( .A(n3087), .Z(n3034) );
  NOR U3197 ( .A(n3086), .B(n3034), .Z(n3089) );
  XOR U3198 ( .A(n3036), .B(n3035), .Z(n3037) );
  IV U3199 ( .A(n3037), .Z(n3082) );
  NOR U3200 ( .A(n98), .B(n134), .Z(n3083) );
  IV U3201 ( .A(n3083), .Z(n3038) );
  NOR U3202 ( .A(n3082), .B(n3038), .Z(n3085) );
  XOR U3203 ( .A(n3040), .B(n3039), .Z(n3041) );
  IV U3204 ( .A(n3041), .Z(n3078) );
  NOR U3205 ( .A(n91), .B(n134), .Z(n3079) );
  IV U3206 ( .A(n3079), .Z(n3042) );
  NOR U3207 ( .A(n3078), .B(n3042), .Z(n3081) );
  IV U3208 ( .A(n3043), .Z(n3045) );
  XOR U3209 ( .A(n3045), .B(n3044), .Z(n3074) );
  NOR U3210 ( .A(n97), .B(n134), .Z(n3075) );
  IV U3211 ( .A(n3075), .Z(n3046) );
  NOR U3212 ( .A(n3074), .B(n3046), .Z(n3077) );
  NOR U3213 ( .A(n96), .B(n134), .Z(n3071) );
  IV U3214 ( .A(n3071), .Z(n3050) );
  XOR U3215 ( .A(n3048), .B(n3047), .Z(n3049) );
  IV U3216 ( .A(n3049), .Z(n3070) );
  NOR U3217 ( .A(n3050), .B(n3070), .Z(n3073) );
  NOR U3218 ( .A(n93), .B(n134), .Z(n3819) );
  IV U3219 ( .A(n3819), .Z(n3052) );
  NOR U3220 ( .A(n136), .B(n168), .Z(n3055) );
  IV U3221 ( .A(n3055), .Z(n3051) );
  NOR U3222 ( .A(n3052), .B(n3051), .Z(n3405) );
  IV U3223 ( .A(n3405), .Z(n3053) );
  NOR U3224 ( .A(n3054), .B(n3053), .Z(n3062) );
  XOR U3225 ( .A(n3056), .B(n3055), .Z(n3057) );
  NOR U3226 ( .A(n3405), .B(n3057), .Z(n3058) );
  NOR U3227 ( .A(n3062), .B(n3058), .Z(n3059) );
  IV U3228 ( .A(n3059), .Z(n3418) );
  NOR U3229 ( .A(n94), .B(n134), .Z(n3417) );
  IV U3230 ( .A(n3417), .Z(n3060) );
  NOR U3231 ( .A(n3418), .B(n3060), .Z(n3061) );
  NOR U3232 ( .A(n3062), .B(n3061), .Z(n3064) );
  NOR U3233 ( .A(n95), .B(n134), .Z(n3065) );
  IV U3234 ( .A(n3065), .Z(n3063) );
  NOR U3235 ( .A(n3064), .B(n3063), .Z(n3069) );
  XOR U3236 ( .A(n3065), .B(n3064), .Z(n3398) );
  XOR U3237 ( .A(n3067), .B(n3066), .Z(n3399) );
  NOR U3238 ( .A(n3398), .B(n3399), .Z(n3068) );
  NOR U3239 ( .A(n3069), .B(n3068), .Z(n3394) );
  XOR U3240 ( .A(n3071), .B(n3070), .Z(n3395) );
  NOR U3241 ( .A(n3394), .B(n3395), .Z(n3072) );
  NOR U3242 ( .A(n3073), .B(n3072), .Z(n3390) );
  XOR U3243 ( .A(n3075), .B(n3074), .Z(n3391) );
  NOR U3244 ( .A(n3390), .B(n3391), .Z(n3076) );
  NOR U3245 ( .A(n3077), .B(n3076), .Z(n3386) );
  XOR U3246 ( .A(n3079), .B(n3078), .Z(n3387) );
  NOR U3247 ( .A(n3386), .B(n3387), .Z(n3080) );
  NOR U3248 ( .A(n3081), .B(n3080), .Z(n3382) );
  XOR U3249 ( .A(n3083), .B(n3082), .Z(n3383) );
  NOR U3250 ( .A(n3382), .B(n3383), .Z(n3084) );
  NOR U3251 ( .A(n3085), .B(n3084), .Z(n3378) );
  XOR U3252 ( .A(n3087), .B(n3086), .Z(n3379) );
  NOR U3253 ( .A(n3378), .B(n3379), .Z(n3088) );
  NOR U3254 ( .A(n3089), .B(n3088), .Z(n3374) );
  XOR U3255 ( .A(n3091), .B(n3090), .Z(n3375) );
  NOR U3256 ( .A(n3374), .B(n3375), .Z(n3092) );
  NOR U3257 ( .A(n3093), .B(n3092), .Z(n3370) );
  XOR U3258 ( .A(n3095), .B(n3094), .Z(n3371) );
  NOR U3259 ( .A(n3370), .B(n3371), .Z(n3096) );
  NOR U3260 ( .A(n3097), .B(n3096), .Z(n3366) );
  XOR U3261 ( .A(n3099), .B(n3098), .Z(n3367) );
  NOR U3262 ( .A(n3366), .B(n3367), .Z(n3100) );
  NOR U3263 ( .A(n3101), .B(n3100), .Z(n3362) );
  XOR U3264 ( .A(n3103), .B(n3102), .Z(n3363) );
  NOR U3265 ( .A(n3362), .B(n3363), .Z(n3104) );
  NOR U3266 ( .A(n3105), .B(n3104), .Z(n3358) );
  XOR U3267 ( .A(n3107), .B(n3106), .Z(n3359) );
  NOR U3268 ( .A(n3358), .B(n3359), .Z(n3108) );
  NOR U3269 ( .A(n3109), .B(n3108), .Z(n3354) );
  XOR U3270 ( .A(n3111), .B(n3110), .Z(n3355) );
  NOR U3271 ( .A(n3354), .B(n3355), .Z(n3112) );
  NOR U3272 ( .A(n3113), .B(n3112), .Z(n3350) );
  XOR U3273 ( .A(n3115), .B(n3114), .Z(n3351) );
  NOR U3274 ( .A(n3350), .B(n3351), .Z(n3116) );
  NOR U3275 ( .A(n3117), .B(n3116), .Z(n3346) );
  XOR U3276 ( .A(n3119), .B(n3118), .Z(n3347) );
  NOR U3277 ( .A(n3346), .B(n3347), .Z(n3120) );
  NOR U3278 ( .A(n3121), .B(n3120), .Z(n3342) );
  XOR U3279 ( .A(n3123), .B(n3122), .Z(n3343) );
  NOR U3280 ( .A(n3342), .B(n3343), .Z(n3124) );
  NOR U3281 ( .A(n3125), .B(n3124), .Z(n3338) );
  XOR U3282 ( .A(n3127), .B(n3126), .Z(n3339) );
  NOR U3283 ( .A(n3338), .B(n3339), .Z(n3128) );
  NOR U3284 ( .A(n3129), .B(n3128), .Z(n3486) );
  XOR U3285 ( .A(n3131), .B(n3130), .Z(n3485) );
  NOR U3286 ( .A(n3486), .B(n3485), .Z(n3132) );
  NOR U3287 ( .A(n3133), .B(n3132), .Z(n3334) );
  XOR U3288 ( .A(n3135), .B(n3134), .Z(n3335) );
  NOR U3289 ( .A(n3334), .B(n3335), .Z(n3136) );
  NOR U3290 ( .A(n3137), .B(n3136), .Z(n3138) );
  IV U3291 ( .A(n3138), .Z(n3332) );
  XOR U3292 ( .A(n3140), .B(n3139), .Z(n3141) );
  IV U3293 ( .A(n3141), .Z(n3331) );
  NOR U3294 ( .A(n3332), .B(n3331), .Z(n3142) );
  NOR U3295 ( .A(n3143), .B(n3142), .Z(n3329) );
  XOR U3296 ( .A(n3145), .B(n3144), .Z(n3146) );
  IV U3297 ( .A(n3146), .Z(n3328) );
  NOR U3298 ( .A(n3329), .B(n3328), .Z(n3147) );
  NOR U3299 ( .A(n3148), .B(n3147), .Z(n3507) );
  XOR U3300 ( .A(n3150), .B(n3149), .Z(n3151) );
  IV U3301 ( .A(n3151), .Z(n3506) );
  NOR U3302 ( .A(n3507), .B(n3506), .Z(n3152) );
  NOR U3303 ( .A(n3153), .B(n3152), .Z(n3326) );
  IV U3304 ( .A(n3154), .Z(n3156) );
  XOR U3305 ( .A(n3156), .B(n3155), .Z(n3325) );
  NOR U3306 ( .A(n3326), .B(n3325), .Z(n3157) );
  NOR U3307 ( .A(n3158), .B(n3157), .Z(n3520) );
  IV U3308 ( .A(n3520), .Z(n3159) );
  NOR U3309 ( .A(n3519), .B(n3159), .Z(n3160) );
  NOR U3310 ( .A(n3161), .B(n3160), .Z(n3321) );
  XOR U3311 ( .A(n3163), .B(n3162), .Z(n3322) );
  NOR U3312 ( .A(n3321), .B(n3322), .Z(n3164) );
  NOR U3313 ( .A(n3165), .B(n3164), .Z(n3531) );
  XOR U3314 ( .A(n3167), .B(n3166), .Z(n3530) );
  NOR U3315 ( .A(n3531), .B(n3530), .Z(n3168) );
  NOR U3316 ( .A(n3169), .B(n3168), .Z(n3537) );
  XOR U3317 ( .A(n3171), .B(n3170), .Z(n3536) );
  NOR U3318 ( .A(n3537), .B(n3536), .Z(n3172) );
  NOR U3319 ( .A(n3173), .B(n3172), .Z(n3174) );
  IV U3320 ( .A(n3174), .Z(n3545) );
  XOR U3321 ( .A(n3176), .B(n3175), .Z(n3177) );
  IV U3322 ( .A(n3177), .Z(n3544) );
  NOR U3323 ( .A(n3545), .B(n3544), .Z(n3178) );
  NOR U3324 ( .A(n3179), .B(n3178), .Z(n3552) );
  XOR U3325 ( .A(n3181), .B(n3180), .Z(n3182) );
  IV U3326 ( .A(n3182), .Z(n3551) );
  NOR U3327 ( .A(n3552), .B(n3551), .Z(n3183) );
  NOR U3328 ( .A(n3184), .B(n3183), .Z(n3319) );
  XOR U3329 ( .A(n3186), .B(n3185), .Z(n3187) );
  IV U3330 ( .A(n3187), .Z(n3318) );
  NOR U3331 ( .A(n3319), .B(n3318), .Z(n3188) );
  NOR U3332 ( .A(n3189), .B(n3188), .Z(n3316) );
  XOR U3333 ( .A(n3191), .B(n3190), .Z(n3192) );
  IV U3334 ( .A(n3192), .Z(n3315) );
  NOR U3335 ( .A(n3316), .B(n3315), .Z(n3193) );
  NOR U3336 ( .A(n3194), .B(n3193), .Z(n3567) );
  XOR U3337 ( .A(n3196), .B(n3195), .Z(n3197) );
  IV U3338 ( .A(n3197), .Z(n3566) );
  NOR U3339 ( .A(n3567), .B(n3566), .Z(n3198) );
  NOR U3340 ( .A(n3199), .B(n3198), .Z(n3314) );
  IV U3341 ( .A(n3200), .Z(n3202) );
  XOR U3342 ( .A(n3202), .B(n3201), .Z(n3313) );
  NOR U3343 ( .A(n3314), .B(n3313), .Z(n3203) );
  NOR U3344 ( .A(n3204), .B(n3203), .Z(n3587) );
  NOR U3345 ( .A(n116), .B(n134), .Z(n3585) );
  IV U3346 ( .A(n3585), .Z(n3312) );
  NOR U3347 ( .A(n3206), .B(n3205), .Z(n3210) );
  NOR U3348 ( .A(n3208), .B(n3207), .Z(n3209) );
  NOR U3349 ( .A(n3210), .B(n3209), .Z(n3600) );
  NOR U3350 ( .A(n115), .B(n138), .Z(n3598) );
  NOR U3351 ( .A(n3212), .B(n3211), .Z(n3216) );
  NOR U3352 ( .A(n3214), .B(n3213), .Z(n3215) );
  NOR U3353 ( .A(n3216), .B(n3215), .Z(n3613) );
  NOR U3354 ( .A(n114), .B(n142), .Z(n3611) );
  IV U3355 ( .A(n3611), .Z(n3297) );
  NOR U3356 ( .A(n3218), .B(n3217), .Z(n3222) );
  NOR U3357 ( .A(n3220), .B(n3219), .Z(n3221) );
  NOR U3358 ( .A(n3222), .B(n3221), .Z(n3616) );
  IV U3359 ( .A(n3616), .Z(n3295) );
  NOR U3360 ( .A(n3224), .B(n3223), .Z(n3228) );
  NOR U3361 ( .A(n3226), .B(n3225), .Z(n3227) );
  NOR U3362 ( .A(n3228), .B(n3227), .Z(n3625) );
  NOR U3363 ( .A(n113), .B(n146), .Z(n3623) );
  IV U3364 ( .A(n3623), .Z(n3294) );
  IV U3365 ( .A(n3229), .Z(n3230) );
  NOR U3366 ( .A(n3231), .B(n3230), .Z(n3235) );
  NOR U3367 ( .A(n3233), .B(n3232), .Z(n3234) );
  NOR U3368 ( .A(n3235), .B(n3234), .Z(n3628) );
  IV U3369 ( .A(n3628), .Z(n3292) );
  NOR U3370 ( .A(n3237), .B(n3236), .Z(n3241) );
  NOR U3371 ( .A(n3239), .B(n3238), .Z(n3240) );
  NOR U3372 ( .A(n3241), .B(n3240), .Z(n3637) );
  NOR U3373 ( .A(n112), .B(n151), .Z(n3635) );
  IV U3374 ( .A(n3635), .Z(n3291) );
  NOR U3375 ( .A(n3243), .B(n3242), .Z(n3247) );
  NOR U3376 ( .A(n3245), .B(n3244), .Z(n3246) );
  NOR U3377 ( .A(n3247), .B(n3246), .Z(n3650) );
  NOR U3378 ( .A(n111), .B(n154), .Z(n3648) );
  NOR U3379 ( .A(n3249), .B(n3248), .Z(n3253) );
  NOR U3380 ( .A(n3251), .B(n3250), .Z(n3252) );
  NOR U3381 ( .A(n3253), .B(n3252), .Z(n3656) );
  NOR U3382 ( .A(n110), .B(n159), .Z(n3654) );
  NOR U3383 ( .A(n3255), .B(n3254), .Z(n3259) );
  NOR U3384 ( .A(n3257), .B(n3256), .Z(n3258) );
  NOR U3385 ( .A(n3259), .B(n3258), .Z(n3677) );
  NOR U3386 ( .A(n3261), .B(n3260), .Z(n3265) );
  NOR U3387 ( .A(n3263), .B(n3262), .Z(n3264) );
  NOR U3388 ( .A(n3265), .B(n3264), .Z(n3662) );
  NOR U3389 ( .A(n108), .B(n162), .Z(n3660) );
  IV U3390 ( .A(n3660), .Z(n3274) );
  IV U3391 ( .A(n3266), .Z(n3267) );
  NOR U3392 ( .A(n3268), .B(n3267), .Z(n3272) );
  NOR U3393 ( .A(n3270), .B(n3269), .Z(n3271) );
  NOR U3394 ( .A(n3272), .B(n3271), .Z(n3667) );
  NOR U3395 ( .A(n164), .B(n87), .Z(n3665) );
  XOR U3396 ( .A(n3667), .B(n3665), .Z(n3669) );
  NOR U3397 ( .A(n166), .B(n107), .Z(n3273) );
  IV U3398 ( .A(n3273), .Z(n3668) );
  XOR U3399 ( .A(n3669), .B(n3668), .Z(n3659) );
  XOR U3400 ( .A(n3274), .B(n3659), .Z(n3661) );
  XOR U3401 ( .A(n3662), .B(n3661), .Z(n3675) );
  NOR U3402 ( .A(n109), .B(n160), .Z(n3673) );
  XOR U3403 ( .A(n3675), .B(n3673), .Z(n3676) );
  XOR U3404 ( .A(n3677), .B(n3676), .Z(n3653) );
  XOR U3405 ( .A(n3654), .B(n3653), .Z(n3275) );
  IV U3406 ( .A(n3275), .Z(n3655) );
  XOR U3407 ( .A(n3656), .B(n3655), .Z(n3684) );
  IV U3408 ( .A(n3276), .Z(n3277) );
  NOR U3409 ( .A(n3278), .B(n3277), .Z(n3282) );
  NOR U3410 ( .A(n3280), .B(n3279), .Z(n3281) );
  NOR U3411 ( .A(n3282), .B(n3281), .Z(n3682) );
  NOR U3412 ( .A(n86), .B(n157), .Z(n3680) );
  XOR U3413 ( .A(n3682), .B(n3680), .Z(n3683) );
  XOR U3414 ( .A(n3684), .B(n3683), .Z(n3647) );
  XOR U3415 ( .A(n3648), .B(n3647), .Z(n3283) );
  IV U3416 ( .A(n3283), .Z(n3649) );
  XOR U3417 ( .A(n3650), .B(n3649), .Z(n3644) );
  IV U3418 ( .A(n3284), .Z(n3285) );
  NOR U3419 ( .A(n3286), .B(n3285), .Z(n3290) );
  NOR U3420 ( .A(n3288), .B(n3287), .Z(n3289) );
  NOR U3421 ( .A(n3290), .B(n3289), .Z(n3642) );
  NOR U3422 ( .A(n85), .B(n152), .Z(n3640) );
  XOR U3423 ( .A(n3642), .B(n3640), .Z(n3643) );
  XOR U3424 ( .A(n3644), .B(n3643), .Z(n3634) );
  XOR U3425 ( .A(n3291), .B(n3634), .Z(n3636) );
  XOR U3426 ( .A(n3637), .B(n3636), .Z(n3629) );
  XOR U3427 ( .A(n3292), .B(n3629), .Z(n3631) );
  NOR U3428 ( .A(n84), .B(n149), .Z(n3293) );
  IV U3429 ( .A(n3293), .Z(n3630) );
  XOR U3430 ( .A(n3631), .B(n3630), .Z(n3622) );
  XOR U3431 ( .A(n3294), .B(n3622), .Z(n3624) );
  XOR U3432 ( .A(n3625), .B(n3624), .Z(n3617) );
  XOR U3433 ( .A(n3295), .B(n3617), .Z(n3619) );
  NOR U3434 ( .A(n83), .B(n144), .Z(n3296) );
  IV U3435 ( .A(n3296), .Z(n3618) );
  XOR U3436 ( .A(n3619), .B(n3618), .Z(n3610) );
  XOR U3437 ( .A(n3297), .B(n3610), .Z(n3612) );
  XOR U3438 ( .A(n3613), .B(n3612), .Z(n3607) );
  IV U3439 ( .A(n3298), .Z(n3299) );
  NOR U3440 ( .A(n3300), .B(n3299), .Z(n3304) );
  NOR U3441 ( .A(n3302), .B(n3301), .Z(n3303) );
  NOR U3442 ( .A(n3304), .B(n3303), .Z(n3605) );
  NOR U3443 ( .A(n82), .B(n140), .Z(n3603) );
  XOR U3444 ( .A(n3605), .B(n3603), .Z(n3606) );
  XOR U3445 ( .A(n3607), .B(n3606), .Z(n3597) );
  XOR U3446 ( .A(n3598), .B(n3597), .Z(n3305) );
  IV U3447 ( .A(n3305), .Z(n3599) );
  XOR U3448 ( .A(n3600), .B(n3599), .Z(n3594) );
  NOR U3449 ( .A(n3307), .B(n3306), .Z(n3311) );
  NOR U3450 ( .A(n3309), .B(n3308), .Z(n3310) );
  NOR U3451 ( .A(n3311), .B(n3310), .Z(n3592) );
  NOR U3452 ( .A(n81), .B(n136), .Z(n3590) );
  XOR U3453 ( .A(n3592), .B(n3590), .Z(n3593) );
  XOR U3454 ( .A(n3594), .B(n3593), .Z(n3584) );
  XOR U3455 ( .A(n3312), .B(n3584), .Z(n3586) );
  XOR U3456 ( .A(n3587), .B(n3586), .Z(n3579) );
  XOR U3457 ( .A(n3314), .B(n3313), .Z(n3573) );
  XOR U3458 ( .A(n3316), .B(n3315), .Z(n3562) );
  NOR U3459 ( .A(n115), .B(n132), .Z(n3561) );
  IV U3460 ( .A(n3561), .Z(n3317) );
  NOR U3461 ( .A(n3562), .B(n3317), .Z(n3564) );
  XOR U3462 ( .A(n3319), .B(n3318), .Z(n3558) );
  NOR U3463 ( .A(n82), .B(n132), .Z(n3557) );
  IV U3464 ( .A(n3557), .Z(n3320) );
  NOR U3465 ( .A(n3558), .B(n3320), .Z(n3560) );
  NOR U3466 ( .A(n113), .B(n132), .Z(n3539) );
  IV U3467 ( .A(n3321), .Z(n3323) );
  XOR U3468 ( .A(n3323), .B(n3322), .Z(n3523) );
  NOR U3469 ( .A(n112), .B(n132), .Z(n3524) );
  IV U3470 ( .A(n3524), .Z(n3324) );
  NOR U3471 ( .A(n3523), .B(n3324), .Z(n3526) );
  XOR U3472 ( .A(n3326), .B(n3325), .Z(n3513) );
  NOR U3473 ( .A(n111), .B(n132), .Z(n3512) );
  IV U3474 ( .A(n3512), .Z(n3327) );
  NOR U3475 ( .A(n3513), .B(n3327), .Z(n3515) );
  XOR U3476 ( .A(n3329), .B(n3328), .Z(n3502) );
  NOR U3477 ( .A(n110), .B(n132), .Z(n3501) );
  IV U3478 ( .A(n3501), .Z(n3330) );
  NOR U3479 ( .A(n3502), .B(n3330), .Z(n3504) );
  XOR U3480 ( .A(n3332), .B(n3331), .Z(n3498) );
  NOR U3481 ( .A(n109), .B(n132), .Z(n3497) );
  IV U3482 ( .A(n3497), .Z(n3333) );
  NOR U3483 ( .A(n3498), .B(n3333), .Z(n3500) );
  IV U3484 ( .A(n3334), .Z(n3336) );
  XOR U3485 ( .A(n3336), .B(n3335), .Z(n3493) );
  NOR U3486 ( .A(n108), .B(n132), .Z(n3494) );
  IV U3487 ( .A(n3494), .Z(n3337) );
  NOR U3488 ( .A(n3493), .B(n3337), .Z(n3496) );
  IV U3489 ( .A(n3338), .Z(n3340) );
  XOR U3490 ( .A(n3340), .B(n3339), .Z(n3481) );
  NOR U3491 ( .A(n107), .B(n132), .Z(n3482) );
  IV U3492 ( .A(n3482), .Z(n3341) );
  NOR U3493 ( .A(n3481), .B(n3341), .Z(n3484) );
  XOR U3494 ( .A(n3343), .B(n3342), .Z(n3344) );
  IV U3495 ( .A(n3344), .Z(n3477) );
  NOR U3496 ( .A(n88), .B(n132), .Z(n3478) );
  IV U3497 ( .A(n3478), .Z(n3345) );
  NOR U3498 ( .A(n3477), .B(n3345), .Z(n3480) );
  XOR U3499 ( .A(n3347), .B(n3346), .Z(n3348) );
  IV U3500 ( .A(n3348), .Z(n3473) );
  NOR U3501 ( .A(n106), .B(n132), .Z(n3474) );
  IV U3502 ( .A(n3474), .Z(n3349) );
  NOR U3503 ( .A(n3473), .B(n3349), .Z(n3476) );
  XOR U3504 ( .A(n3351), .B(n3350), .Z(n3352) );
  IV U3505 ( .A(n3352), .Z(n3469) );
  NOR U3506 ( .A(n105), .B(n132), .Z(n3470) );
  IV U3507 ( .A(n3470), .Z(n3353) );
  NOR U3508 ( .A(n3469), .B(n3353), .Z(n3472) );
  XOR U3509 ( .A(n3355), .B(n3354), .Z(n3356) );
  IV U3510 ( .A(n3356), .Z(n3465) );
  NOR U3511 ( .A(n104), .B(n132), .Z(n3466) );
  IV U3512 ( .A(n3466), .Z(n3357) );
  NOR U3513 ( .A(n3465), .B(n3357), .Z(n3468) );
  XOR U3514 ( .A(n3359), .B(n3358), .Z(n3360) );
  IV U3515 ( .A(n3360), .Z(n3461) );
  NOR U3516 ( .A(n89), .B(n132), .Z(n3462) );
  IV U3517 ( .A(n3462), .Z(n3361) );
  NOR U3518 ( .A(n3461), .B(n3361), .Z(n3464) );
  XOR U3519 ( .A(n3363), .B(n3362), .Z(n3364) );
  IV U3520 ( .A(n3364), .Z(n3457) );
  NOR U3521 ( .A(n103), .B(n132), .Z(n3458) );
  IV U3522 ( .A(n3458), .Z(n3365) );
  NOR U3523 ( .A(n3457), .B(n3365), .Z(n3460) );
  XOR U3524 ( .A(n3367), .B(n3366), .Z(n3368) );
  IV U3525 ( .A(n3368), .Z(n3453) );
  NOR U3526 ( .A(n90), .B(n132), .Z(n3454) );
  IV U3527 ( .A(n3454), .Z(n3369) );
  NOR U3528 ( .A(n3453), .B(n3369), .Z(n3456) );
  XOR U3529 ( .A(n3371), .B(n3370), .Z(n3372) );
  IV U3530 ( .A(n3372), .Z(n3449) );
  NOR U3531 ( .A(n102), .B(n132), .Z(n3450) );
  IV U3532 ( .A(n3450), .Z(n3373) );
  NOR U3533 ( .A(n3449), .B(n3373), .Z(n3452) );
  XOR U3534 ( .A(n3375), .B(n3374), .Z(n3376) );
  IV U3535 ( .A(n3376), .Z(n3445) );
  NOR U3536 ( .A(n101), .B(n132), .Z(n3446) );
  IV U3537 ( .A(n3446), .Z(n3377) );
  NOR U3538 ( .A(n3445), .B(n3377), .Z(n3448) );
  XOR U3539 ( .A(n3379), .B(n3378), .Z(n3380) );
  IV U3540 ( .A(n3380), .Z(n3441) );
  NOR U3541 ( .A(n100), .B(n132), .Z(n3442) );
  IV U3542 ( .A(n3442), .Z(n3381) );
  NOR U3543 ( .A(n3441), .B(n3381), .Z(n3444) );
  XOR U3544 ( .A(n3383), .B(n3382), .Z(n3384) );
  IV U3545 ( .A(n3384), .Z(n3437) );
  NOR U3546 ( .A(n99), .B(n132), .Z(n3438) );
  IV U3547 ( .A(n3438), .Z(n3385) );
  NOR U3548 ( .A(n3437), .B(n3385), .Z(n3440) );
  XOR U3549 ( .A(n3387), .B(n3386), .Z(n3388) );
  IV U3550 ( .A(n3388), .Z(n3433) );
  NOR U3551 ( .A(n98), .B(n132), .Z(n3434) );
  IV U3552 ( .A(n3434), .Z(n3389) );
  NOR U3553 ( .A(n3433), .B(n3389), .Z(n3436) );
  XOR U3554 ( .A(n3391), .B(n3390), .Z(n3392) );
  IV U3555 ( .A(n3392), .Z(n3429) );
  NOR U3556 ( .A(n91), .B(n132), .Z(n3430) );
  IV U3557 ( .A(n3430), .Z(n3393) );
  NOR U3558 ( .A(n3429), .B(n3393), .Z(n3432) );
  XOR U3559 ( .A(n3395), .B(n3394), .Z(n3396) );
  IV U3560 ( .A(n3396), .Z(n3425) );
  NOR U3561 ( .A(n97), .B(n132), .Z(n3426) );
  IV U3562 ( .A(n3426), .Z(n3397) );
  NOR U3563 ( .A(n3425), .B(n3397), .Z(n3428) );
  XOR U3564 ( .A(n3399), .B(n3398), .Z(n3400) );
  IV U3565 ( .A(n3400), .Z(n3421) );
  NOR U3566 ( .A(n96), .B(n132), .Z(n3422) );
  IV U3567 ( .A(n3422), .Z(n3401) );
  NOR U3568 ( .A(n3421), .B(n3401), .Z(n3424) );
  NOR U3569 ( .A(n93), .B(n132), .Z(n4221) );
  IV U3570 ( .A(n4221), .Z(n3403) );
  NOR U3571 ( .A(n134), .B(n168), .Z(n3406) );
  IV U3572 ( .A(n3406), .Z(n3402) );
  NOR U3573 ( .A(n3403), .B(n3402), .Z(n3817) );
  IV U3574 ( .A(n3817), .Z(n3404) );
  NOR U3575 ( .A(n3405), .B(n3404), .Z(n3413) );
  XOR U3576 ( .A(n3407), .B(n3406), .Z(n3408) );
  NOR U3577 ( .A(n3817), .B(n3408), .Z(n3409) );
  NOR U3578 ( .A(n3413), .B(n3409), .Z(n3410) );
  IV U3579 ( .A(n3410), .Z(n3830) );
  NOR U3580 ( .A(n94), .B(n132), .Z(n3829) );
  IV U3581 ( .A(n3829), .Z(n3411) );
  NOR U3582 ( .A(n3830), .B(n3411), .Z(n3412) );
  NOR U3583 ( .A(n3413), .B(n3412), .Z(n3416) );
  NOR U3584 ( .A(n95), .B(n132), .Z(n3415) );
  IV U3585 ( .A(n3415), .Z(n3414) );
  NOR U3586 ( .A(n3416), .B(n3414), .Z(n3420) );
  XOR U3587 ( .A(n3416), .B(n3415), .Z(n3810) );
  XOR U3588 ( .A(n3418), .B(n3417), .Z(n3811) );
  NOR U3589 ( .A(n3810), .B(n3811), .Z(n3419) );
  NOR U3590 ( .A(n3420), .B(n3419), .Z(n3806) );
  XOR U3591 ( .A(n3422), .B(n3421), .Z(n3807) );
  NOR U3592 ( .A(n3806), .B(n3807), .Z(n3423) );
  NOR U3593 ( .A(n3424), .B(n3423), .Z(n3802) );
  XOR U3594 ( .A(n3426), .B(n3425), .Z(n3803) );
  NOR U3595 ( .A(n3802), .B(n3803), .Z(n3427) );
  NOR U3596 ( .A(n3428), .B(n3427), .Z(n3798) );
  XOR U3597 ( .A(n3430), .B(n3429), .Z(n3799) );
  NOR U3598 ( .A(n3798), .B(n3799), .Z(n3431) );
  NOR U3599 ( .A(n3432), .B(n3431), .Z(n3794) );
  XOR U3600 ( .A(n3434), .B(n3433), .Z(n3795) );
  NOR U3601 ( .A(n3794), .B(n3795), .Z(n3435) );
  NOR U3602 ( .A(n3436), .B(n3435), .Z(n3790) );
  XOR U3603 ( .A(n3438), .B(n3437), .Z(n3791) );
  NOR U3604 ( .A(n3790), .B(n3791), .Z(n3439) );
  NOR U3605 ( .A(n3440), .B(n3439), .Z(n3786) );
  XOR U3606 ( .A(n3442), .B(n3441), .Z(n3787) );
  NOR U3607 ( .A(n3786), .B(n3787), .Z(n3443) );
  NOR U3608 ( .A(n3444), .B(n3443), .Z(n3782) );
  XOR U3609 ( .A(n3446), .B(n3445), .Z(n3783) );
  NOR U3610 ( .A(n3782), .B(n3783), .Z(n3447) );
  NOR U3611 ( .A(n3448), .B(n3447), .Z(n3778) );
  XOR U3612 ( .A(n3450), .B(n3449), .Z(n3779) );
  NOR U3613 ( .A(n3778), .B(n3779), .Z(n3451) );
  NOR U3614 ( .A(n3452), .B(n3451), .Z(n3774) );
  XOR U3615 ( .A(n3454), .B(n3453), .Z(n3775) );
  NOR U3616 ( .A(n3774), .B(n3775), .Z(n3455) );
  NOR U3617 ( .A(n3456), .B(n3455), .Z(n3770) );
  XOR U3618 ( .A(n3458), .B(n3457), .Z(n3771) );
  NOR U3619 ( .A(n3770), .B(n3771), .Z(n3459) );
  NOR U3620 ( .A(n3460), .B(n3459), .Z(n3766) );
  XOR U3621 ( .A(n3462), .B(n3461), .Z(n3767) );
  NOR U3622 ( .A(n3766), .B(n3767), .Z(n3463) );
  NOR U3623 ( .A(n3464), .B(n3463), .Z(n3762) );
  XOR U3624 ( .A(n3466), .B(n3465), .Z(n3763) );
  NOR U3625 ( .A(n3762), .B(n3763), .Z(n3467) );
  NOR U3626 ( .A(n3468), .B(n3467), .Z(n3758) );
  XOR U3627 ( .A(n3470), .B(n3469), .Z(n3759) );
  NOR U3628 ( .A(n3758), .B(n3759), .Z(n3471) );
  NOR U3629 ( .A(n3472), .B(n3471), .Z(n3754) );
  XOR U3630 ( .A(n3474), .B(n3473), .Z(n3755) );
  NOR U3631 ( .A(n3754), .B(n3755), .Z(n3475) );
  NOR U3632 ( .A(n3476), .B(n3475), .Z(n3750) );
  XOR U3633 ( .A(n3478), .B(n3477), .Z(n3751) );
  NOR U3634 ( .A(n3750), .B(n3751), .Z(n3479) );
  NOR U3635 ( .A(n3480), .B(n3479), .Z(n3746) );
  XOR U3636 ( .A(n3482), .B(n3481), .Z(n3747) );
  NOR U3637 ( .A(n3746), .B(n3747), .Z(n3483) );
  NOR U3638 ( .A(n3484), .B(n3483), .Z(n3489) );
  XOR U3639 ( .A(n3486), .B(n3485), .Z(n3488) );
  IV U3640 ( .A(n3488), .Z(n3487) );
  NOR U3641 ( .A(n3489), .B(n3487), .Z(n3492) );
  XOR U3642 ( .A(n3489), .B(n3488), .Z(n3743) );
  NOR U3643 ( .A(n87), .B(n132), .Z(n3744) );
  IV U3644 ( .A(n3744), .Z(n3490) );
  NOR U3645 ( .A(n3743), .B(n3490), .Z(n3491) );
  NOR U3646 ( .A(n3492), .B(n3491), .Z(n3739) );
  XOR U3647 ( .A(n3494), .B(n3493), .Z(n3740) );
  NOR U3648 ( .A(n3739), .B(n3740), .Z(n3495) );
  NOR U3649 ( .A(n3496), .B(n3495), .Z(n3735) );
  XOR U3650 ( .A(n3498), .B(n3497), .Z(n3736) );
  NOR U3651 ( .A(n3735), .B(n3736), .Z(n3499) );
  NOR U3652 ( .A(n3500), .B(n3499), .Z(n3734) );
  XOR U3653 ( .A(n3502), .B(n3501), .Z(n3733) );
  NOR U3654 ( .A(n3734), .B(n3733), .Z(n3503) );
  NOR U3655 ( .A(n3504), .B(n3503), .Z(n3509) );
  NOR U3656 ( .A(n86), .B(n132), .Z(n3508) );
  IV U3657 ( .A(n3508), .Z(n3505) );
  NOR U3658 ( .A(n3509), .B(n3505), .Z(n3511) );
  XOR U3659 ( .A(n3507), .B(n3506), .Z(n3732) );
  XOR U3660 ( .A(n3509), .B(n3508), .Z(n3731) );
  NOR U3661 ( .A(n3732), .B(n3731), .Z(n3510) );
  NOR U3662 ( .A(n3511), .B(n3510), .Z(n3730) );
  XOR U3663 ( .A(n3513), .B(n3512), .Z(n3729) );
  NOR U3664 ( .A(n3730), .B(n3729), .Z(n3514) );
  NOR U3665 ( .A(n3515), .B(n3514), .Z(n3518) );
  NOR U3666 ( .A(n85), .B(n132), .Z(n3517) );
  IV U3667 ( .A(n3517), .Z(n3516) );
  NOR U3668 ( .A(n3518), .B(n3516), .Z(n3522) );
  XOR U3669 ( .A(n3518), .B(n3517), .Z(n3728) );
  XOR U3670 ( .A(n3520), .B(n3519), .Z(n3727) );
  NOR U3671 ( .A(n3728), .B(n3727), .Z(n3521) );
  NOR U3672 ( .A(n3522), .B(n3521), .Z(n3722) );
  XOR U3673 ( .A(n3524), .B(n3523), .Z(n3721) );
  NOR U3674 ( .A(n3722), .B(n3721), .Z(n3525) );
  NOR U3675 ( .A(n3526), .B(n3525), .Z(n3529) );
  NOR U3676 ( .A(n84), .B(n132), .Z(n3528) );
  IV U3677 ( .A(n3528), .Z(n3527) );
  NOR U3678 ( .A(n3529), .B(n3527), .Z(n3534) );
  XOR U3679 ( .A(n3529), .B(n3528), .Z(n3718) );
  XOR U3680 ( .A(n3531), .B(n3530), .Z(n3719) );
  IV U3681 ( .A(n3719), .Z(n3532) );
  NOR U3682 ( .A(n3718), .B(n3532), .Z(n3533) );
  NOR U3683 ( .A(n3534), .B(n3533), .Z(n3538) );
  IV U3684 ( .A(n3538), .Z(n3535) );
  NOR U3685 ( .A(n3539), .B(n3535), .Z(n3541) );
  XOR U3686 ( .A(n3537), .B(n3536), .Z(n3716) );
  XOR U3687 ( .A(n3539), .B(n3538), .Z(n3715) );
  NOR U3688 ( .A(n3716), .B(n3715), .Z(n3540) );
  NOR U3689 ( .A(n3541), .B(n3540), .Z(n3542) );
  IV U3690 ( .A(n3542), .Z(n3547) );
  NOR U3691 ( .A(n83), .B(n132), .Z(n3546) );
  IV U3692 ( .A(n3546), .Z(n3543) );
  NOR U3693 ( .A(n3547), .B(n3543), .Z(n3549) );
  XOR U3694 ( .A(n3545), .B(n3544), .Z(n3712) );
  XOR U3695 ( .A(n3547), .B(n3546), .Z(n3711) );
  NOR U3696 ( .A(n3712), .B(n3711), .Z(n3548) );
  NOR U3697 ( .A(n3549), .B(n3548), .Z(n3554) );
  NOR U3698 ( .A(n114), .B(n132), .Z(n3553) );
  IV U3699 ( .A(n3553), .Z(n3550) );
  NOR U3700 ( .A(n3554), .B(n3550), .Z(n3556) );
  XOR U3701 ( .A(n3552), .B(n3551), .Z(n3710) );
  XOR U3702 ( .A(n3554), .B(n3553), .Z(n3709) );
  NOR U3703 ( .A(n3710), .B(n3709), .Z(n3555) );
  NOR U3704 ( .A(n3556), .B(n3555), .Z(n3708) );
  XOR U3705 ( .A(n3558), .B(n3557), .Z(n3707) );
  NOR U3706 ( .A(n3708), .B(n3707), .Z(n3559) );
  NOR U3707 ( .A(n3560), .B(n3559), .Z(n3706) );
  XOR U3708 ( .A(n3562), .B(n3561), .Z(n3705) );
  NOR U3709 ( .A(n3706), .B(n3705), .Z(n3563) );
  NOR U3710 ( .A(n3564), .B(n3563), .Z(n3569) );
  NOR U3711 ( .A(n81), .B(n132), .Z(n3568) );
  IV U3712 ( .A(n3568), .Z(n3565) );
  NOR U3713 ( .A(n3569), .B(n3565), .Z(n3571) );
  XOR U3714 ( .A(n3567), .B(n3566), .Z(n3704) );
  XOR U3715 ( .A(n3569), .B(n3568), .Z(n3703) );
  NOR U3716 ( .A(n3704), .B(n3703), .Z(n3570) );
  NOR U3717 ( .A(n3571), .B(n3570), .Z(n3572) );
  NOR U3718 ( .A(n3573), .B(n3572), .Z(n3577) );
  IV U3719 ( .A(n3572), .Z(n3574) );
  XOR U3720 ( .A(n3574), .B(n3573), .Z(n3702) );
  NOR U3721 ( .A(n116), .B(n132), .Z(n3575) );
  IV U3722 ( .A(n3575), .Z(n3701) );
  NOR U3723 ( .A(n3702), .B(n3701), .Z(n3576) );
  NOR U3724 ( .A(n3577), .B(n3576), .Z(n3578) );
  NOR U3725 ( .A(n3579), .B(n3578), .Z(n3583) );
  IV U3726 ( .A(n3578), .Z(n3580) );
  XOR U3727 ( .A(n3580), .B(n3579), .Z(n3700) );
  NOR U3728 ( .A(n80), .B(n132), .Z(n3581) );
  IV U3729 ( .A(n3581), .Z(n3699) );
  NOR U3730 ( .A(n3700), .B(n3699), .Z(n3582) );
  NOR U3731 ( .A(n3583), .B(n3582), .Z(n3989) );
  NOR U3732 ( .A(n3585), .B(n3584), .Z(n3589) );
  NOR U3733 ( .A(n3587), .B(n3586), .Z(n3588) );
  NOR U3734 ( .A(n3589), .B(n3588), .Z(n3995) );
  NOR U3735 ( .A(n80), .B(n134), .Z(n3993) );
  IV U3736 ( .A(n3590), .Z(n3591) );
  NOR U3737 ( .A(n3592), .B(n3591), .Z(n3596) );
  NOR U3738 ( .A(n3594), .B(n3593), .Z(n3595) );
  NOR U3739 ( .A(n3596), .B(n3595), .Z(n4099) );
  NOR U3740 ( .A(n3598), .B(n3597), .Z(n3602) );
  NOR U3741 ( .A(n3600), .B(n3599), .Z(n3601) );
  NOR U3742 ( .A(n3602), .B(n3601), .Z(n4001) );
  NOR U3743 ( .A(n81), .B(n138), .Z(n3999) );
  IV U3744 ( .A(n3999), .Z(n3697) );
  IV U3745 ( .A(n3603), .Z(n3604) );
  NOR U3746 ( .A(n3605), .B(n3604), .Z(n3609) );
  NOR U3747 ( .A(n3607), .B(n3606), .Z(n3608) );
  NOR U3748 ( .A(n3609), .B(n3608), .Z(n4004) );
  IV U3749 ( .A(n4004), .Z(n3695) );
  NOR U3750 ( .A(n3611), .B(n3610), .Z(n3615) );
  NOR U3751 ( .A(n3613), .B(n3612), .Z(n3614) );
  NOR U3752 ( .A(n3615), .B(n3614), .Z(n4013) );
  NOR U3753 ( .A(n82), .B(n142), .Z(n4011) );
  IV U3754 ( .A(n4011), .Z(n3694) );
  NOR U3755 ( .A(n3617), .B(n3616), .Z(n3621) );
  NOR U3756 ( .A(n3619), .B(n3618), .Z(n3620) );
  NOR U3757 ( .A(n3621), .B(n3620), .Z(n4016) );
  IV U3758 ( .A(n4016), .Z(n3692) );
  NOR U3759 ( .A(n3623), .B(n3622), .Z(n3627) );
  NOR U3760 ( .A(n3625), .B(n3624), .Z(n3626) );
  NOR U3761 ( .A(n3627), .B(n3626), .Z(n4025) );
  NOR U3762 ( .A(n83), .B(n146), .Z(n4023) );
  IV U3763 ( .A(n4023), .Z(n3691) );
  NOR U3764 ( .A(n3629), .B(n3628), .Z(n3633) );
  NOR U3765 ( .A(n3631), .B(n3630), .Z(n3632) );
  NOR U3766 ( .A(n3633), .B(n3632), .Z(n4087) );
  IV U3767 ( .A(n4087), .Z(n3689) );
  NOR U3768 ( .A(n3635), .B(n3634), .Z(n3639) );
  NOR U3769 ( .A(n3637), .B(n3636), .Z(n3638) );
  NOR U3770 ( .A(n3639), .B(n3638), .Z(n4031) );
  NOR U3771 ( .A(n84), .B(n151), .Z(n4029) );
  IV U3772 ( .A(n4029), .Z(n3688) );
  IV U3773 ( .A(n3640), .Z(n3641) );
  NOR U3774 ( .A(n3642), .B(n3641), .Z(n3646) );
  NOR U3775 ( .A(n3644), .B(n3643), .Z(n3645) );
  NOR U3776 ( .A(n3646), .B(n3645), .Z(n4084) );
  NOR U3777 ( .A(n3648), .B(n3647), .Z(n3652) );
  NOR U3778 ( .A(n3650), .B(n3649), .Z(n3651) );
  NOR U3779 ( .A(n3652), .B(n3651), .Z(n4037) );
  NOR U3780 ( .A(n85), .B(n154), .Z(n4035) );
  NOR U3781 ( .A(n3654), .B(n3653), .Z(n3658) );
  NOR U3782 ( .A(n3656), .B(n3655), .Z(n3657) );
  NOR U3783 ( .A(n3658), .B(n3657), .Z(n4051) );
  NOR U3784 ( .A(n86), .B(n159), .Z(n4049) );
  NOR U3785 ( .A(n3660), .B(n3659), .Z(n3664) );
  NOR U3786 ( .A(n3662), .B(n3661), .Z(n3663) );
  NOR U3787 ( .A(n3664), .B(n3663), .Z(n4058) );
  NOR U3788 ( .A(n109), .B(n162), .Z(n4055) );
  IV U3789 ( .A(n3665), .Z(n3666) );
  NOR U3790 ( .A(n3667), .B(n3666), .Z(n3671) );
  NOR U3791 ( .A(n3669), .B(n3668), .Z(n3670) );
  NOR U3792 ( .A(n3671), .B(n3670), .Z(n4063) );
  NOR U3793 ( .A(n164), .B(n108), .Z(n4061) );
  XOR U3794 ( .A(n4063), .B(n4061), .Z(n4065) );
  NOR U3795 ( .A(n166), .B(n87), .Z(n3672) );
  IV U3796 ( .A(n3672), .Z(n4064) );
  XOR U3797 ( .A(n4065), .B(n4064), .Z(n4054) );
  XOR U3798 ( .A(n4055), .B(n4054), .Z(n4056) );
  XOR U3799 ( .A(n4058), .B(n4056), .Z(n4073) );
  NOR U3800 ( .A(n110), .B(n160), .Z(n4072) );
  IV U3801 ( .A(n3673), .Z(n3674) );
  NOR U3802 ( .A(n3675), .B(n3674), .Z(n3679) );
  NOR U3803 ( .A(n3677), .B(n3676), .Z(n3678) );
  NOR U3804 ( .A(n3679), .B(n3678), .Z(n4070) );
  XOR U3805 ( .A(n4072), .B(n4070), .Z(n4074) );
  XOR U3806 ( .A(n4073), .B(n4074), .Z(n4047) );
  XOR U3807 ( .A(n4049), .B(n4047), .Z(n4050) );
  XOR U3808 ( .A(n4051), .B(n4050), .Z(n4044) );
  IV U3809 ( .A(n3680), .Z(n3681) );
  NOR U3810 ( .A(n3682), .B(n3681), .Z(n3686) );
  NOR U3811 ( .A(n3684), .B(n3683), .Z(n3685) );
  NOR U3812 ( .A(n3686), .B(n3685), .Z(n4042) );
  NOR U3813 ( .A(n111), .B(n157), .Z(n4040) );
  XOR U3814 ( .A(n4042), .B(n4040), .Z(n4043) );
  XOR U3815 ( .A(n4044), .B(n4043), .Z(n4034) );
  XOR U3816 ( .A(n4035), .B(n4034), .Z(n3687) );
  IV U3817 ( .A(n3687), .Z(n4036) );
  XOR U3818 ( .A(n4037), .B(n4036), .Z(n4082) );
  NOR U3819 ( .A(n112), .B(n152), .Z(n4080) );
  XOR U3820 ( .A(n4082), .B(n4080), .Z(n4083) );
  XOR U3821 ( .A(n4084), .B(n4083), .Z(n4028) );
  XOR U3822 ( .A(n3688), .B(n4028), .Z(n4030) );
  XOR U3823 ( .A(n4031), .B(n4030), .Z(n4088) );
  XOR U3824 ( .A(n3689), .B(n4088), .Z(n4090) );
  NOR U3825 ( .A(n113), .B(n149), .Z(n3690) );
  IV U3826 ( .A(n3690), .Z(n4089) );
  XOR U3827 ( .A(n4090), .B(n4089), .Z(n4022) );
  XOR U3828 ( .A(n3691), .B(n4022), .Z(n4024) );
  XOR U3829 ( .A(n4025), .B(n4024), .Z(n4017) );
  XOR U3830 ( .A(n3692), .B(n4017), .Z(n4019) );
  NOR U3831 ( .A(n114), .B(n144), .Z(n3693) );
  IV U3832 ( .A(n3693), .Z(n4018) );
  XOR U3833 ( .A(n4019), .B(n4018), .Z(n4010) );
  XOR U3834 ( .A(n3694), .B(n4010), .Z(n4012) );
  XOR U3835 ( .A(n4013), .B(n4012), .Z(n4005) );
  XOR U3836 ( .A(n3695), .B(n4005), .Z(n4007) );
  NOR U3837 ( .A(n115), .B(n140), .Z(n3696) );
  IV U3838 ( .A(n3696), .Z(n4006) );
  XOR U3839 ( .A(n4007), .B(n4006), .Z(n3998) );
  XOR U3840 ( .A(n3697), .B(n3998), .Z(n4000) );
  XOR U3841 ( .A(n4001), .B(n4000), .Z(n4097) );
  NOR U3842 ( .A(n116), .B(n136), .Z(n4095) );
  XOR U3843 ( .A(n4097), .B(n4095), .Z(n4098) );
  XOR U3844 ( .A(n4099), .B(n4098), .Z(n3992) );
  XOR U3845 ( .A(n3993), .B(n3992), .Z(n3698) );
  IV U3846 ( .A(n3698), .Z(n3994) );
  XOR U3847 ( .A(n3995), .B(n3994), .Z(n3987) );
  NOR U3848 ( .A(n117), .B(n132), .Z(n3985) );
  XOR U3849 ( .A(n3987), .B(n3985), .Z(n3988) );
  XOR U3850 ( .A(n3989), .B(n3988), .Z(n3980) );
  NOR U3851 ( .A(n3981), .B(n3980), .Z(n3984) );
  NOR U3852 ( .A(n117), .B(n130), .Z(n3975) );
  XOR U3853 ( .A(n3700), .B(n3699), .Z(n3976) );
  NOR U3854 ( .A(n3975), .B(n3976), .Z(n3979) );
  NOR U3855 ( .A(n80), .B(n130), .Z(n3970) );
  XOR U3856 ( .A(n3702), .B(n3701), .Z(n3971) );
  NOR U3857 ( .A(n3970), .B(n3971), .Z(n3974) );
  NOR U3858 ( .A(n116), .B(n130), .Z(n3966) );
  XOR U3859 ( .A(n3704), .B(n3703), .Z(n3965) );
  NOR U3860 ( .A(n3966), .B(n3965), .Z(n3969) );
  NOR U3861 ( .A(n81), .B(n130), .Z(n3961) );
  XOR U3862 ( .A(n3706), .B(n3705), .Z(n3960) );
  NOR U3863 ( .A(n3961), .B(n3960), .Z(n3964) );
  NOR U3864 ( .A(n115), .B(n130), .Z(n3956) );
  XOR U3865 ( .A(n3708), .B(n3707), .Z(n3955) );
  NOR U3866 ( .A(n3956), .B(n3955), .Z(n3959) );
  NOR U3867 ( .A(n82), .B(n130), .Z(n3951) );
  XOR U3868 ( .A(n3710), .B(n3709), .Z(n3950) );
  NOR U3869 ( .A(n3951), .B(n3950), .Z(n3954) );
  XOR U3870 ( .A(n3712), .B(n3711), .Z(n3713) );
  IV U3871 ( .A(n3713), .Z(n3945) );
  NOR U3872 ( .A(n114), .B(n130), .Z(n3946) );
  IV U3873 ( .A(n3946), .Z(n3714) );
  NOR U3874 ( .A(n3945), .B(n3714), .Z(n3948) );
  XOR U3875 ( .A(n3716), .B(n3715), .Z(n3942) );
  NOR U3876 ( .A(n83), .B(n130), .Z(n3941) );
  IV U3877 ( .A(n3941), .Z(n3717) );
  NOR U3878 ( .A(n3942), .B(n3717), .Z(n3944) );
  XOR U3879 ( .A(n3719), .B(n3718), .Z(n3937) );
  NOR U3880 ( .A(n113), .B(n130), .Z(n3938) );
  IV U3881 ( .A(n3938), .Z(n3720) );
  NOR U3882 ( .A(n3937), .B(n3720), .Z(n3940) );
  XOR U3883 ( .A(n3722), .B(n3721), .Z(n3725) );
  IV U3884 ( .A(n3725), .Z(n3724) );
  NOR U3885 ( .A(n84), .B(n130), .Z(n3723) );
  IV U3886 ( .A(n3723), .Z(n3726) );
  NOR U3887 ( .A(n3724), .B(n3726), .Z(n3936) );
  XOR U3888 ( .A(n3726), .B(n3725), .Z(n4129) );
  NOR U3889 ( .A(n112), .B(n130), .Z(n3930) );
  XOR U3890 ( .A(n3728), .B(n3727), .Z(n3929) );
  NOR U3891 ( .A(n3930), .B(n3929), .Z(n3933) );
  NOR U3892 ( .A(n85), .B(n130), .Z(n3925) );
  XOR U3893 ( .A(n3730), .B(n3729), .Z(n3924) );
  NOR U3894 ( .A(n3925), .B(n3924), .Z(n3928) );
  NOR U3895 ( .A(n111), .B(n130), .Z(n3920) );
  XOR U3896 ( .A(n3732), .B(n3731), .Z(n3919) );
  NOR U3897 ( .A(n3920), .B(n3919), .Z(n3923) );
  NOR U3898 ( .A(n86), .B(n130), .Z(n3915) );
  XOR U3899 ( .A(n3734), .B(n3733), .Z(n3914) );
  NOR U3900 ( .A(n3915), .B(n3914), .Z(n3918) );
  IV U3901 ( .A(n3735), .Z(n3737) );
  XOR U3902 ( .A(n3737), .B(n3736), .Z(n3909) );
  NOR U3903 ( .A(n110), .B(n130), .Z(n3910) );
  IV U3904 ( .A(n3910), .Z(n3738) );
  NOR U3905 ( .A(n3909), .B(n3738), .Z(n3912) );
  IV U3906 ( .A(n3739), .Z(n3741) );
  XOR U3907 ( .A(n3741), .B(n3740), .Z(n3905) );
  NOR U3908 ( .A(n109), .B(n130), .Z(n3906) );
  IV U3909 ( .A(n3906), .Z(n3742) );
  NOR U3910 ( .A(n3905), .B(n3742), .Z(n3908) );
  XOR U3911 ( .A(n3744), .B(n3743), .Z(n3901) );
  NOR U3912 ( .A(n108), .B(n130), .Z(n3902) );
  IV U3913 ( .A(n3902), .Z(n3745) );
  NOR U3914 ( .A(n3901), .B(n3745), .Z(n3904) );
  IV U3915 ( .A(n3746), .Z(n3748) );
  XOR U3916 ( .A(n3748), .B(n3747), .Z(n3897) );
  NOR U3917 ( .A(n87), .B(n130), .Z(n3898) );
  IV U3918 ( .A(n3898), .Z(n3749) );
  NOR U3919 ( .A(n3897), .B(n3749), .Z(n3900) );
  XOR U3920 ( .A(n3751), .B(n3750), .Z(n3752) );
  IV U3921 ( .A(n3752), .Z(n3893) );
  NOR U3922 ( .A(n107), .B(n130), .Z(n3894) );
  IV U3923 ( .A(n3894), .Z(n3753) );
  NOR U3924 ( .A(n3893), .B(n3753), .Z(n3896) );
  XOR U3925 ( .A(n3755), .B(n3754), .Z(n3756) );
  IV U3926 ( .A(n3756), .Z(n3889) );
  NOR U3927 ( .A(n88), .B(n130), .Z(n3890) );
  IV U3928 ( .A(n3890), .Z(n3757) );
  NOR U3929 ( .A(n3889), .B(n3757), .Z(n3892) );
  XOR U3930 ( .A(n3759), .B(n3758), .Z(n3760) );
  IV U3931 ( .A(n3760), .Z(n3885) );
  NOR U3932 ( .A(n106), .B(n130), .Z(n3886) );
  IV U3933 ( .A(n3886), .Z(n3761) );
  NOR U3934 ( .A(n3885), .B(n3761), .Z(n3888) );
  XOR U3935 ( .A(n3763), .B(n3762), .Z(n3764) );
  IV U3936 ( .A(n3764), .Z(n3881) );
  NOR U3937 ( .A(n105), .B(n130), .Z(n3882) );
  IV U3938 ( .A(n3882), .Z(n3765) );
  NOR U3939 ( .A(n3881), .B(n3765), .Z(n3884) );
  IV U3940 ( .A(n3766), .Z(n3768) );
  XOR U3941 ( .A(n3768), .B(n3767), .Z(n3877) );
  NOR U3942 ( .A(n104), .B(n130), .Z(n3878) );
  IV U3943 ( .A(n3878), .Z(n3769) );
  NOR U3944 ( .A(n3877), .B(n3769), .Z(n3880) );
  XOR U3945 ( .A(n3771), .B(n3770), .Z(n3772) );
  IV U3946 ( .A(n3772), .Z(n3873) );
  NOR U3947 ( .A(n89), .B(n130), .Z(n3874) );
  IV U3948 ( .A(n3874), .Z(n3773) );
  NOR U3949 ( .A(n3873), .B(n3773), .Z(n3876) );
  XOR U3950 ( .A(n3775), .B(n3774), .Z(n3776) );
  IV U3951 ( .A(n3776), .Z(n3869) );
  NOR U3952 ( .A(n103), .B(n130), .Z(n3870) );
  IV U3953 ( .A(n3870), .Z(n3777) );
  NOR U3954 ( .A(n3869), .B(n3777), .Z(n3872) );
  XOR U3955 ( .A(n3779), .B(n3778), .Z(n3780) );
  IV U3956 ( .A(n3780), .Z(n3865) );
  NOR U3957 ( .A(n90), .B(n130), .Z(n3866) );
  IV U3958 ( .A(n3866), .Z(n3781) );
  NOR U3959 ( .A(n3865), .B(n3781), .Z(n3868) );
  XOR U3960 ( .A(n3783), .B(n3782), .Z(n3784) );
  IV U3961 ( .A(n3784), .Z(n3861) );
  NOR U3962 ( .A(n102), .B(n130), .Z(n3862) );
  IV U3963 ( .A(n3862), .Z(n3785) );
  NOR U3964 ( .A(n3861), .B(n3785), .Z(n3864) );
  XOR U3965 ( .A(n3787), .B(n3786), .Z(n3788) );
  IV U3966 ( .A(n3788), .Z(n3857) );
  NOR U3967 ( .A(n101), .B(n130), .Z(n3858) );
  IV U3968 ( .A(n3858), .Z(n3789) );
  NOR U3969 ( .A(n3857), .B(n3789), .Z(n3860) );
  XOR U3970 ( .A(n3791), .B(n3790), .Z(n3792) );
  IV U3971 ( .A(n3792), .Z(n3853) );
  NOR U3972 ( .A(n100), .B(n130), .Z(n3854) );
  IV U3973 ( .A(n3854), .Z(n3793) );
  NOR U3974 ( .A(n3853), .B(n3793), .Z(n3856) );
  XOR U3975 ( .A(n3795), .B(n3794), .Z(n3796) );
  IV U3976 ( .A(n3796), .Z(n3849) );
  NOR U3977 ( .A(n99), .B(n130), .Z(n3850) );
  IV U3978 ( .A(n3850), .Z(n3797) );
  NOR U3979 ( .A(n3849), .B(n3797), .Z(n3852) );
  XOR U3980 ( .A(n3799), .B(n3798), .Z(n3800) );
  IV U3981 ( .A(n3800), .Z(n3845) );
  NOR U3982 ( .A(n98), .B(n130), .Z(n3846) );
  IV U3983 ( .A(n3846), .Z(n3801) );
  NOR U3984 ( .A(n3845), .B(n3801), .Z(n3848) );
  XOR U3985 ( .A(n3803), .B(n3802), .Z(n3804) );
  IV U3986 ( .A(n3804), .Z(n3841) );
  NOR U3987 ( .A(n91), .B(n130), .Z(n3842) );
  IV U3988 ( .A(n3842), .Z(n3805) );
  NOR U3989 ( .A(n3841), .B(n3805), .Z(n3844) );
  IV U3990 ( .A(n3806), .Z(n3808) );
  XOR U3991 ( .A(n3808), .B(n3807), .Z(n3837) );
  NOR U3992 ( .A(n97), .B(n130), .Z(n3838) );
  IV U3993 ( .A(n3838), .Z(n3809) );
  NOR U3994 ( .A(n3837), .B(n3809), .Z(n3840) );
  NOR U3995 ( .A(n96), .B(n130), .Z(n3834) );
  IV U3996 ( .A(n3834), .Z(n3813) );
  XOR U3997 ( .A(n3811), .B(n3810), .Z(n3812) );
  IV U3998 ( .A(n3812), .Z(n3833) );
  NOR U3999 ( .A(n3813), .B(n3833), .Z(n3836) );
  NOR U4000 ( .A(n93), .B(n130), .Z(n4532) );
  IV U4001 ( .A(n4532), .Z(n3815) );
  NOR U4002 ( .A(n132), .B(n168), .Z(n3818) );
  IV U4003 ( .A(n3818), .Z(n3814) );
  NOR U4004 ( .A(n3815), .B(n3814), .Z(n4219) );
  IV U4005 ( .A(n4219), .Z(n3816) );
  NOR U4006 ( .A(n3817), .B(n3816), .Z(n3825) );
  XOR U4007 ( .A(n3819), .B(n3818), .Z(n3820) );
  NOR U4008 ( .A(n4219), .B(n3820), .Z(n3821) );
  NOR U4009 ( .A(n3825), .B(n3821), .Z(n3822) );
  IV U4010 ( .A(n3822), .Z(n4232) );
  NOR U4011 ( .A(n94), .B(n130), .Z(n4231) );
  IV U4012 ( .A(n4231), .Z(n3823) );
  NOR U4013 ( .A(n4232), .B(n3823), .Z(n3824) );
  NOR U4014 ( .A(n3825), .B(n3824), .Z(n3828) );
  NOR U4015 ( .A(n95), .B(n130), .Z(n3827) );
  IV U4016 ( .A(n3827), .Z(n3826) );
  NOR U4017 ( .A(n3828), .B(n3826), .Z(n3832) );
  XOR U4018 ( .A(n3828), .B(n3827), .Z(n4212) );
  XOR U4019 ( .A(n3830), .B(n3829), .Z(n4213) );
  NOR U4020 ( .A(n4212), .B(n4213), .Z(n3831) );
  NOR U4021 ( .A(n3832), .B(n3831), .Z(n4208) );
  XOR U4022 ( .A(n3834), .B(n3833), .Z(n4209) );
  NOR U4023 ( .A(n4208), .B(n4209), .Z(n3835) );
  NOR U4024 ( .A(n3836), .B(n3835), .Z(n4204) );
  XOR U4025 ( .A(n3838), .B(n3837), .Z(n4205) );
  NOR U4026 ( .A(n4204), .B(n4205), .Z(n3839) );
  NOR U4027 ( .A(n3840), .B(n3839), .Z(n4200) );
  XOR U4028 ( .A(n3842), .B(n3841), .Z(n4201) );
  NOR U4029 ( .A(n4200), .B(n4201), .Z(n3843) );
  NOR U4030 ( .A(n3844), .B(n3843), .Z(n4196) );
  XOR U4031 ( .A(n3846), .B(n3845), .Z(n4197) );
  NOR U4032 ( .A(n4196), .B(n4197), .Z(n3847) );
  NOR U4033 ( .A(n3848), .B(n3847), .Z(n4192) );
  XOR U4034 ( .A(n3850), .B(n3849), .Z(n4193) );
  NOR U4035 ( .A(n4192), .B(n4193), .Z(n3851) );
  NOR U4036 ( .A(n3852), .B(n3851), .Z(n4188) );
  XOR U4037 ( .A(n3854), .B(n3853), .Z(n4189) );
  NOR U4038 ( .A(n4188), .B(n4189), .Z(n3855) );
  NOR U4039 ( .A(n3856), .B(n3855), .Z(n4184) );
  XOR U4040 ( .A(n3858), .B(n3857), .Z(n4185) );
  NOR U4041 ( .A(n4184), .B(n4185), .Z(n3859) );
  NOR U4042 ( .A(n3860), .B(n3859), .Z(n4180) );
  XOR U4043 ( .A(n3862), .B(n3861), .Z(n4181) );
  NOR U4044 ( .A(n4180), .B(n4181), .Z(n3863) );
  NOR U4045 ( .A(n3864), .B(n3863), .Z(n4176) );
  XOR U4046 ( .A(n3866), .B(n3865), .Z(n4177) );
  NOR U4047 ( .A(n4176), .B(n4177), .Z(n3867) );
  NOR U4048 ( .A(n3868), .B(n3867), .Z(n4172) );
  XOR U4049 ( .A(n3870), .B(n3869), .Z(n4173) );
  NOR U4050 ( .A(n4172), .B(n4173), .Z(n3871) );
  NOR U4051 ( .A(n3872), .B(n3871), .Z(n4168) );
  XOR U4052 ( .A(n3874), .B(n3873), .Z(n4169) );
  NOR U4053 ( .A(n4168), .B(n4169), .Z(n3875) );
  NOR U4054 ( .A(n3876), .B(n3875), .Z(n4164) );
  XOR U4055 ( .A(n3878), .B(n3877), .Z(n4165) );
  NOR U4056 ( .A(n4164), .B(n4165), .Z(n3879) );
  NOR U4057 ( .A(n3880), .B(n3879), .Z(n4160) );
  XOR U4058 ( .A(n3882), .B(n3881), .Z(n4161) );
  NOR U4059 ( .A(n4160), .B(n4161), .Z(n3883) );
  NOR U4060 ( .A(n3884), .B(n3883), .Z(n4156) );
  XOR U4061 ( .A(n3886), .B(n3885), .Z(n4157) );
  NOR U4062 ( .A(n4156), .B(n4157), .Z(n3887) );
  NOR U4063 ( .A(n3888), .B(n3887), .Z(n4152) );
  XOR U4064 ( .A(n3890), .B(n3889), .Z(n4153) );
  NOR U4065 ( .A(n4152), .B(n4153), .Z(n3891) );
  NOR U4066 ( .A(n3892), .B(n3891), .Z(n4148) );
  XOR U4067 ( .A(n3894), .B(n3893), .Z(n4149) );
  NOR U4068 ( .A(n4148), .B(n4149), .Z(n3895) );
  NOR U4069 ( .A(n3896), .B(n3895), .Z(n4144) );
  XOR U4070 ( .A(n3898), .B(n3897), .Z(n4145) );
  NOR U4071 ( .A(n4144), .B(n4145), .Z(n3899) );
  NOR U4072 ( .A(n3900), .B(n3899), .Z(n4309) );
  XOR U4073 ( .A(n3902), .B(n3901), .Z(n4308) );
  NOR U4074 ( .A(n4309), .B(n4308), .Z(n3903) );
  NOR U4075 ( .A(n3904), .B(n3903), .Z(n4140) );
  XOR U4076 ( .A(n3906), .B(n3905), .Z(n4141) );
  NOR U4077 ( .A(n4140), .B(n4141), .Z(n3907) );
  NOR U4078 ( .A(n3908), .B(n3907), .Z(n4136) );
  XOR U4079 ( .A(n3910), .B(n3909), .Z(n4137) );
  NOR U4080 ( .A(n4136), .B(n4137), .Z(n3911) );
  NOR U4081 ( .A(n3912), .B(n3911), .Z(n3913) );
  IV U4082 ( .A(n3913), .Z(n4134) );
  XOR U4083 ( .A(n3915), .B(n3914), .Z(n3916) );
  IV U4084 ( .A(n3916), .Z(n4133) );
  NOR U4085 ( .A(n4134), .B(n4133), .Z(n3917) );
  NOR U4086 ( .A(n3918), .B(n3917), .Z(n4329) );
  XOR U4087 ( .A(n3920), .B(n3919), .Z(n3921) );
  IV U4088 ( .A(n3921), .Z(n4328) );
  NOR U4089 ( .A(n4329), .B(n4328), .Z(n3922) );
  NOR U4090 ( .A(n3923), .B(n3922), .Z(n4335) );
  XOR U4091 ( .A(n3925), .B(n3924), .Z(n4334) );
  IV U4092 ( .A(n4334), .Z(n3926) );
  NOR U4093 ( .A(n4335), .B(n3926), .Z(n3927) );
  NOR U4094 ( .A(n3928), .B(n3927), .Z(n4131) );
  XOR U4095 ( .A(n3930), .B(n3929), .Z(n3931) );
  IV U4096 ( .A(n3931), .Z(n4130) );
  NOR U4097 ( .A(n4131), .B(n4130), .Z(n3932) );
  NOR U4098 ( .A(n3933), .B(n3932), .Z(n3934) );
  IV U4099 ( .A(n3934), .Z(n4128) );
  NOR U4100 ( .A(n4129), .B(n4128), .Z(n3935) );
  NOR U4101 ( .A(n3936), .B(n3935), .Z(n4124) );
  XOR U4102 ( .A(n3938), .B(n3937), .Z(n4125) );
  NOR U4103 ( .A(n4124), .B(n4125), .Z(n3939) );
  NOR U4104 ( .A(n3940), .B(n3939), .Z(n4120) );
  XOR U4105 ( .A(n3942), .B(n3941), .Z(n4121) );
  NOR U4106 ( .A(n4120), .B(n4121), .Z(n3943) );
  NOR U4107 ( .A(n3944), .B(n3943), .Z(n4116) );
  XOR U4108 ( .A(n3946), .B(n3945), .Z(n4117) );
  NOR U4109 ( .A(n4116), .B(n4117), .Z(n3947) );
  NOR U4110 ( .A(n3948), .B(n3947), .Z(n3949) );
  IV U4111 ( .A(n3949), .Z(n4114) );
  XOR U4112 ( .A(n3951), .B(n3950), .Z(n3952) );
  IV U4113 ( .A(n3952), .Z(n4113) );
  NOR U4114 ( .A(n4114), .B(n4113), .Z(n3953) );
  NOR U4115 ( .A(n3954), .B(n3953), .Z(n4372) );
  XOR U4116 ( .A(n3956), .B(n3955), .Z(n4371) );
  IV U4117 ( .A(n4371), .Z(n3957) );
  NOR U4118 ( .A(n4372), .B(n3957), .Z(n3958) );
  NOR U4119 ( .A(n3959), .B(n3958), .Z(n4111) );
  XOR U4120 ( .A(n3961), .B(n3960), .Z(n3962) );
  IV U4121 ( .A(n3962), .Z(n4110) );
  NOR U4122 ( .A(n4111), .B(n4110), .Z(n3963) );
  NOR U4123 ( .A(n3964), .B(n3963), .Z(n4108) );
  XOR U4124 ( .A(n3966), .B(n3965), .Z(n3967) );
  IV U4125 ( .A(n3967), .Z(n4107) );
  NOR U4126 ( .A(n4108), .B(n4107), .Z(n3968) );
  NOR U4127 ( .A(n3969), .B(n3968), .Z(n4386) );
  IV U4128 ( .A(n3970), .Z(n3972) );
  XOR U4129 ( .A(n3972), .B(n3971), .Z(n4385) );
  NOR U4130 ( .A(n4386), .B(n4385), .Z(n3973) );
  NOR U4131 ( .A(n3974), .B(n3973), .Z(n4105) );
  IV U4132 ( .A(n3975), .Z(n3977) );
  XOR U4133 ( .A(n3977), .B(n3976), .Z(n4104) );
  NOR U4134 ( .A(n4105), .B(n4104), .Z(n3978) );
  NOR U4135 ( .A(n3979), .B(n3978), .Z(n4397) );
  XOR U4136 ( .A(n3981), .B(n3980), .Z(n3982) );
  IV U4137 ( .A(n3982), .Z(n4396) );
  NOR U4138 ( .A(n4397), .B(n4396), .Z(n3983) );
  NOR U4139 ( .A(n3984), .B(n3983), .Z(n4720) );
  NOR U4140 ( .A(n119), .B(n130), .Z(n4718) );
  IV U4141 ( .A(n3985), .Z(n3986) );
  NOR U4142 ( .A(n3987), .B(n3986), .Z(n3991) );
  NOR U4143 ( .A(n3989), .B(n3988), .Z(n3990) );
  NOR U4144 ( .A(n3991), .B(n3990), .Z(n4841) );
  NOR U4145 ( .A(n3993), .B(n3992), .Z(n3997) );
  NOR U4146 ( .A(n3995), .B(n3994), .Z(n3996) );
  NOR U4147 ( .A(n3997), .B(n3996), .Z(n4726) );
  NOR U4148 ( .A(n117), .B(n134), .Z(n4724) );
  NOR U4149 ( .A(n3999), .B(n3998), .Z(n4003) );
  NOR U4150 ( .A(n4001), .B(n4000), .Z(n4002) );
  NOR U4151 ( .A(n4003), .B(n4002), .Z(n4732) );
  NOR U4152 ( .A(n116), .B(n138), .Z(n4730) );
  NOR U4153 ( .A(n4005), .B(n4004), .Z(n4009) );
  NOR U4154 ( .A(n4007), .B(n4006), .Z(n4008) );
  NOR U4155 ( .A(n4009), .B(n4008), .Z(n4826) );
  NOR U4156 ( .A(n4011), .B(n4010), .Z(n4015) );
  NOR U4157 ( .A(n4013), .B(n4012), .Z(n4014) );
  NOR U4158 ( .A(n4015), .B(n4014), .Z(n4738) );
  NOR U4159 ( .A(n115), .B(n142), .Z(n4736) );
  NOR U4160 ( .A(n4017), .B(n4016), .Z(n4021) );
  NOR U4161 ( .A(n4019), .B(n4018), .Z(n4020) );
  NOR U4162 ( .A(n4021), .B(n4020), .Z(n4819) );
  NOR U4163 ( .A(n4023), .B(n4022), .Z(n4027) );
  NOR U4164 ( .A(n4025), .B(n4024), .Z(n4026) );
  NOR U4165 ( .A(n4027), .B(n4026), .Z(n4745) );
  NOR U4166 ( .A(n114), .B(n146), .Z(n4743) );
  NOR U4167 ( .A(n4029), .B(n4028), .Z(n4033) );
  NOR U4168 ( .A(n4031), .B(n4030), .Z(n4032) );
  NOR U4169 ( .A(n4033), .B(n4032), .Z(n4752) );
  NOR U4170 ( .A(n113), .B(n151), .Z(n4749) );
  NOR U4171 ( .A(n4035), .B(n4034), .Z(n4039) );
  NOR U4172 ( .A(n4037), .B(n4036), .Z(n4038) );
  NOR U4173 ( .A(n4039), .B(n4038), .Z(n4765) );
  NOR U4174 ( .A(n112), .B(n154), .Z(n4763) );
  IV U4175 ( .A(n4040), .Z(n4041) );
  NOR U4176 ( .A(n4042), .B(n4041), .Z(n4046) );
  NOR U4177 ( .A(n4044), .B(n4043), .Z(n4045) );
  NOR U4178 ( .A(n4046), .B(n4045), .Z(n4801) );
  IV U4179 ( .A(n4047), .Z(n4048) );
  NOR U4180 ( .A(n4049), .B(n4048), .Z(n4053) );
  NOR U4181 ( .A(n4051), .B(n4050), .Z(n4052) );
  NOR U4182 ( .A(n4053), .B(n4052), .Z(n4771) );
  NOR U4183 ( .A(n111), .B(n159), .Z(n4769) );
  IV U4184 ( .A(n4769), .Z(n4078) );
  NOR U4185 ( .A(n4055), .B(n4054), .Z(n4060) );
  IV U4186 ( .A(n4056), .Z(n4057) );
  NOR U4187 ( .A(n4058), .B(n4057), .Z(n4059) );
  NOR U4188 ( .A(n4060), .B(n4059), .Z(n4777) );
  NOR U4189 ( .A(n110), .B(n162), .Z(n4775) );
  IV U4190 ( .A(n4775), .Z(n4069) );
  IV U4191 ( .A(n4061), .Z(n4062) );
  NOR U4192 ( .A(n4063), .B(n4062), .Z(n4067) );
  NOR U4193 ( .A(n4065), .B(n4064), .Z(n4066) );
  NOR U4194 ( .A(n4067), .B(n4066), .Z(n4782) );
  NOR U4195 ( .A(n164), .B(n109), .Z(n4780) );
  XOR U4196 ( .A(n4782), .B(n4780), .Z(n4784) );
  NOR U4197 ( .A(n166), .B(n108), .Z(n4068) );
  IV U4198 ( .A(n4068), .Z(n4783) );
  XOR U4199 ( .A(n4784), .B(n4783), .Z(n4774) );
  XOR U4200 ( .A(n4069), .B(n4774), .Z(n4776) );
  XOR U4201 ( .A(n4777), .B(n4776), .Z(n4791) );
  IV U4202 ( .A(n4070), .Z(n4071) );
  NOR U4203 ( .A(n4072), .B(n4071), .Z(n4076) );
  NOR U4204 ( .A(n4074), .B(n4073), .Z(n4075) );
  NOR U4205 ( .A(n4076), .B(n4075), .Z(n4789) );
  XOR U4206 ( .A(n4791), .B(n4789), .Z(n4793) );
  NOR U4207 ( .A(n86), .B(n160), .Z(n4077) );
  IV U4208 ( .A(n4077), .Z(n4792) );
  XOR U4209 ( .A(n4793), .B(n4792), .Z(n4768) );
  XOR U4210 ( .A(n4078), .B(n4768), .Z(n4770) );
  XOR U4211 ( .A(n4771), .B(n4770), .Z(n4799) );
  NOR U4212 ( .A(n85), .B(n157), .Z(n4797) );
  XOR U4213 ( .A(n4799), .B(n4797), .Z(n4800) );
  XOR U4214 ( .A(n4801), .B(n4800), .Z(n4762) );
  XOR U4215 ( .A(n4763), .B(n4762), .Z(n4079) );
  IV U4216 ( .A(n4079), .Z(n4764) );
  XOR U4217 ( .A(n4765), .B(n4764), .Z(n4759) );
  IV U4218 ( .A(n4080), .Z(n4081) );
  NOR U4219 ( .A(n4082), .B(n4081), .Z(n4086) );
  NOR U4220 ( .A(n4084), .B(n4083), .Z(n4085) );
  NOR U4221 ( .A(n4086), .B(n4085), .Z(n4757) );
  NOR U4222 ( .A(n84), .B(n152), .Z(n4755) );
  XOR U4223 ( .A(n4757), .B(n4755), .Z(n4758) );
  XOR U4224 ( .A(n4759), .B(n4758), .Z(n4748) );
  XOR U4225 ( .A(n4749), .B(n4748), .Z(n4750) );
  XOR U4226 ( .A(n4752), .B(n4750), .Z(n4809) );
  NOR U4227 ( .A(n83), .B(n149), .Z(n4808) );
  NOR U4228 ( .A(n4088), .B(n4087), .Z(n4092) );
  NOR U4229 ( .A(n4090), .B(n4089), .Z(n4091) );
  NOR U4230 ( .A(n4092), .B(n4091), .Z(n4806) );
  XOR U4231 ( .A(n4808), .B(n4806), .Z(n4810) );
  XOR U4232 ( .A(n4809), .B(n4810), .Z(n4741) );
  XOR U4233 ( .A(n4743), .B(n4741), .Z(n4744) );
  XOR U4234 ( .A(n4745), .B(n4744), .Z(n4817) );
  NOR U4235 ( .A(n82), .B(n144), .Z(n4815) );
  XOR U4236 ( .A(n4817), .B(n4815), .Z(n4818) );
  XOR U4237 ( .A(n4819), .B(n4818), .Z(n4735) );
  XOR U4238 ( .A(n4736), .B(n4735), .Z(n4093) );
  IV U4239 ( .A(n4093), .Z(n4737) );
  XOR U4240 ( .A(n4738), .B(n4737), .Z(n4824) );
  NOR U4241 ( .A(n81), .B(n140), .Z(n4822) );
  XOR U4242 ( .A(n4824), .B(n4822), .Z(n4825) );
  XOR U4243 ( .A(n4826), .B(n4825), .Z(n4729) );
  XOR U4244 ( .A(n4730), .B(n4729), .Z(n4094) );
  IV U4245 ( .A(n4094), .Z(n4731) );
  XOR U4246 ( .A(n4732), .B(n4731), .Z(n4833) );
  IV U4247 ( .A(n4095), .Z(n4096) );
  NOR U4248 ( .A(n4097), .B(n4096), .Z(n4101) );
  NOR U4249 ( .A(n4099), .B(n4098), .Z(n4100) );
  NOR U4250 ( .A(n4101), .B(n4100), .Z(n4831) );
  NOR U4251 ( .A(n80), .B(n136), .Z(n4829) );
  XOR U4252 ( .A(n4831), .B(n4829), .Z(n4832) );
  XOR U4253 ( .A(n4833), .B(n4832), .Z(n4723) );
  XOR U4254 ( .A(n4724), .B(n4723), .Z(n4102) );
  IV U4255 ( .A(n4102), .Z(n4725) );
  XOR U4256 ( .A(n4726), .B(n4725), .Z(n4839) );
  NOR U4257 ( .A(n79), .B(n132), .Z(n4837) );
  XOR U4258 ( .A(n4839), .B(n4837), .Z(n4840) );
  XOR U4259 ( .A(n4841), .B(n4840), .Z(n4717) );
  XOR U4260 ( .A(n4718), .B(n4717), .Z(n4103) );
  IV U4261 ( .A(n4103), .Z(n4719) );
  XOR U4262 ( .A(n4720), .B(n4719), .Z(n4714) );
  XOR U4263 ( .A(n4105), .B(n4104), .Z(n4392) );
  NOR U4264 ( .A(n79), .B(n129), .Z(n4391) );
  IV U4265 ( .A(n4391), .Z(n4106) );
  NOR U4266 ( .A(n4392), .B(n4106), .Z(n4394) );
  XOR U4267 ( .A(n4108), .B(n4107), .Z(n4381) );
  NOR U4268 ( .A(n80), .B(n129), .Z(n4380) );
  IV U4269 ( .A(n4380), .Z(n4109) );
  NOR U4270 ( .A(n4381), .B(n4109), .Z(n4383) );
  XOR U4271 ( .A(n4111), .B(n4110), .Z(n4377) );
  NOR U4272 ( .A(n116), .B(n129), .Z(n4376) );
  IV U4273 ( .A(n4376), .Z(n4112) );
  NOR U4274 ( .A(n4377), .B(n4112), .Z(n4379) );
  NOR U4275 ( .A(n81), .B(n129), .Z(n4370) );
  XOR U4276 ( .A(n4114), .B(n4113), .Z(n4365) );
  NOR U4277 ( .A(n115), .B(n129), .Z(n4364) );
  IV U4278 ( .A(n4364), .Z(n4115) );
  NOR U4279 ( .A(n4365), .B(n4115), .Z(n4367) );
  IV U4280 ( .A(n4116), .Z(n4118) );
  XOR U4281 ( .A(n4118), .B(n4117), .Z(n4360) );
  NOR U4282 ( .A(n82), .B(n129), .Z(n4361) );
  IV U4283 ( .A(n4361), .Z(n4119) );
  NOR U4284 ( .A(n4360), .B(n4119), .Z(n4363) );
  IV U4285 ( .A(n4120), .Z(n4122) );
  XOR U4286 ( .A(n4122), .B(n4121), .Z(n4356) );
  NOR U4287 ( .A(n114), .B(n129), .Z(n4357) );
  IV U4288 ( .A(n4357), .Z(n4123) );
  NOR U4289 ( .A(n4356), .B(n4123), .Z(n4359) );
  IV U4290 ( .A(n4124), .Z(n4126) );
  XOR U4291 ( .A(n4126), .B(n4125), .Z(n4351) );
  NOR U4292 ( .A(n83), .B(n129), .Z(n4352) );
  IV U4293 ( .A(n4352), .Z(n4127) );
  NOR U4294 ( .A(n4351), .B(n4127), .Z(n4355) );
  XOR U4295 ( .A(n4129), .B(n4128), .Z(n4348) );
  XOR U4296 ( .A(n4131), .B(n4130), .Z(n4343) );
  NOR U4297 ( .A(n84), .B(n129), .Z(n4342) );
  IV U4298 ( .A(n4342), .Z(n4132) );
  NOR U4299 ( .A(n4343), .B(n4132), .Z(n4345) );
  XOR U4300 ( .A(n4134), .B(n4133), .Z(n4324) );
  NOR U4301 ( .A(n111), .B(n129), .Z(n4323) );
  IV U4302 ( .A(n4323), .Z(n4135) );
  NOR U4303 ( .A(n4324), .B(n4135), .Z(n4326) );
  IV U4304 ( .A(n4136), .Z(n4138) );
  XOR U4305 ( .A(n4138), .B(n4137), .Z(n4319) );
  NOR U4306 ( .A(n86), .B(n129), .Z(n4320) );
  IV U4307 ( .A(n4320), .Z(n4139) );
  NOR U4308 ( .A(n4319), .B(n4139), .Z(n4322) );
  IV U4309 ( .A(n4140), .Z(n4142) );
  XOR U4310 ( .A(n4142), .B(n4141), .Z(n4315) );
  NOR U4311 ( .A(n110), .B(n129), .Z(n4316) );
  IV U4312 ( .A(n4316), .Z(n4143) );
  NOR U4313 ( .A(n4315), .B(n4143), .Z(n4318) );
  IV U4314 ( .A(n4144), .Z(n4146) );
  XOR U4315 ( .A(n4146), .B(n4145), .Z(n4303) );
  NOR U4316 ( .A(n108), .B(n129), .Z(n4304) );
  IV U4317 ( .A(n4304), .Z(n4147) );
  NOR U4318 ( .A(n4303), .B(n4147), .Z(n4306) );
  XOR U4319 ( .A(n4149), .B(n4148), .Z(n4150) );
  IV U4320 ( .A(n4150), .Z(n4299) );
  NOR U4321 ( .A(n87), .B(n129), .Z(n4300) );
  IV U4322 ( .A(n4300), .Z(n4151) );
  NOR U4323 ( .A(n4299), .B(n4151), .Z(n4302) );
  XOR U4324 ( .A(n4153), .B(n4152), .Z(n4154) );
  IV U4325 ( .A(n4154), .Z(n4295) );
  NOR U4326 ( .A(n107), .B(n129), .Z(n4296) );
  IV U4327 ( .A(n4296), .Z(n4155) );
  NOR U4328 ( .A(n4295), .B(n4155), .Z(n4298) );
  XOR U4329 ( .A(n4157), .B(n4156), .Z(n4158) );
  IV U4330 ( .A(n4158), .Z(n4291) );
  NOR U4331 ( .A(n88), .B(n129), .Z(n4292) );
  IV U4332 ( .A(n4292), .Z(n4159) );
  NOR U4333 ( .A(n4291), .B(n4159), .Z(n4294) );
  XOR U4334 ( .A(n4161), .B(n4160), .Z(n4162) );
  IV U4335 ( .A(n4162), .Z(n4287) );
  NOR U4336 ( .A(n106), .B(n129), .Z(n4288) );
  IV U4337 ( .A(n4288), .Z(n4163) );
  NOR U4338 ( .A(n4287), .B(n4163), .Z(n4290) );
  XOR U4339 ( .A(n4165), .B(n4164), .Z(n4166) );
  IV U4340 ( .A(n4166), .Z(n4283) );
  NOR U4341 ( .A(n105), .B(n129), .Z(n4284) );
  IV U4342 ( .A(n4284), .Z(n4167) );
  NOR U4343 ( .A(n4283), .B(n4167), .Z(n4286) );
  XOR U4344 ( .A(n4169), .B(n4168), .Z(n4170) );
  IV U4345 ( .A(n4170), .Z(n4279) );
  NOR U4346 ( .A(n104), .B(n129), .Z(n4280) );
  IV U4347 ( .A(n4280), .Z(n4171) );
  NOR U4348 ( .A(n4279), .B(n4171), .Z(n4282) );
  XOR U4349 ( .A(n4173), .B(n4172), .Z(n4174) );
  IV U4350 ( .A(n4174), .Z(n4275) );
  NOR U4351 ( .A(n89), .B(n129), .Z(n4276) );
  IV U4352 ( .A(n4276), .Z(n4175) );
  NOR U4353 ( .A(n4275), .B(n4175), .Z(n4278) );
  XOR U4354 ( .A(n4177), .B(n4176), .Z(n4178) );
  IV U4355 ( .A(n4178), .Z(n4271) );
  NOR U4356 ( .A(n103), .B(n129), .Z(n4272) );
  IV U4357 ( .A(n4272), .Z(n4179) );
  NOR U4358 ( .A(n4271), .B(n4179), .Z(n4274) );
  XOR U4359 ( .A(n4181), .B(n4180), .Z(n4182) );
  IV U4360 ( .A(n4182), .Z(n4267) );
  NOR U4361 ( .A(n90), .B(n129), .Z(n4268) );
  IV U4362 ( .A(n4268), .Z(n4183) );
  NOR U4363 ( .A(n4267), .B(n4183), .Z(n4270) );
  XOR U4364 ( .A(n4185), .B(n4184), .Z(n4186) );
  IV U4365 ( .A(n4186), .Z(n4263) );
  NOR U4366 ( .A(n102), .B(n129), .Z(n4264) );
  IV U4367 ( .A(n4264), .Z(n4187) );
  NOR U4368 ( .A(n4263), .B(n4187), .Z(n4266) );
  XOR U4369 ( .A(n4189), .B(n4188), .Z(n4190) );
  IV U4370 ( .A(n4190), .Z(n4259) );
  NOR U4371 ( .A(n101), .B(n129), .Z(n4260) );
  IV U4372 ( .A(n4260), .Z(n4191) );
  NOR U4373 ( .A(n4259), .B(n4191), .Z(n4262) );
  XOR U4374 ( .A(n4193), .B(n4192), .Z(n4194) );
  IV U4375 ( .A(n4194), .Z(n4255) );
  NOR U4376 ( .A(n100), .B(n129), .Z(n4256) );
  IV U4377 ( .A(n4256), .Z(n4195) );
  NOR U4378 ( .A(n4255), .B(n4195), .Z(n4258) );
  XOR U4379 ( .A(n4197), .B(n4196), .Z(n4198) );
  IV U4380 ( .A(n4198), .Z(n4251) );
  NOR U4381 ( .A(n99), .B(n129), .Z(n4252) );
  IV U4382 ( .A(n4252), .Z(n4199) );
  NOR U4383 ( .A(n4251), .B(n4199), .Z(n4254) );
  XOR U4384 ( .A(n4201), .B(n4200), .Z(n4202) );
  IV U4385 ( .A(n4202), .Z(n4247) );
  NOR U4386 ( .A(n98), .B(n129), .Z(n4248) );
  IV U4387 ( .A(n4248), .Z(n4203) );
  NOR U4388 ( .A(n4247), .B(n4203), .Z(n4250) );
  IV U4389 ( .A(n4204), .Z(n4206) );
  XOR U4390 ( .A(n4206), .B(n4205), .Z(n4243) );
  NOR U4391 ( .A(n91), .B(n129), .Z(n4244) );
  IV U4392 ( .A(n4244), .Z(n4207) );
  NOR U4393 ( .A(n4243), .B(n4207), .Z(n4246) );
  IV U4394 ( .A(n4208), .Z(n4210) );
  XOR U4395 ( .A(n4210), .B(n4209), .Z(n4239) );
  NOR U4396 ( .A(n97), .B(n129), .Z(n4240) );
  IV U4397 ( .A(n4240), .Z(n4211) );
  NOR U4398 ( .A(n4239), .B(n4211), .Z(n4242) );
  XOR U4399 ( .A(n4213), .B(n4212), .Z(n4214) );
  IV U4400 ( .A(n4214), .Z(n4235) );
  NOR U4401 ( .A(n96), .B(n129), .Z(n4236) );
  IV U4402 ( .A(n4236), .Z(n4215) );
  NOR U4403 ( .A(n4235), .B(n4215), .Z(n4238) );
  NOR U4404 ( .A(n93), .B(n129), .Z(n4968) );
  IV U4405 ( .A(n4968), .Z(n4217) );
  NOR U4406 ( .A(n130), .B(n168), .Z(n4220) );
  IV U4407 ( .A(n4220), .Z(n4216) );
  NOR U4408 ( .A(n4217), .B(n4216), .Z(n4530) );
  IV U4409 ( .A(n4530), .Z(n4218) );
  NOR U4410 ( .A(n4219), .B(n4218), .Z(n4227) );
  XOR U4411 ( .A(n4221), .B(n4220), .Z(n4222) );
  NOR U4412 ( .A(n4530), .B(n4222), .Z(n4223) );
  NOR U4413 ( .A(n4227), .B(n4223), .Z(n4224) );
  IV U4414 ( .A(n4224), .Z(n4543) );
  NOR U4415 ( .A(n94), .B(n129), .Z(n4542) );
  IV U4416 ( .A(n4542), .Z(n4225) );
  NOR U4417 ( .A(n4543), .B(n4225), .Z(n4226) );
  NOR U4418 ( .A(n4227), .B(n4226), .Z(n4230) );
  NOR U4419 ( .A(n95), .B(n129), .Z(n4229) );
  IV U4420 ( .A(n4229), .Z(n4228) );
  NOR U4421 ( .A(n4230), .B(n4228), .Z(n4234) );
  XOR U4422 ( .A(n4230), .B(n4229), .Z(n4523) );
  XOR U4423 ( .A(n4232), .B(n4231), .Z(n4524) );
  NOR U4424 ( .A(n4523), .B(n4524), .Z(n4233) );
  NOR U4425 ( .A(n4234), .B(n4233), .Z(n4519) );
  XOR U4426 ( .A(n4236), .B(n4235), .Z(n4520) );
  NOR U4427 ( .A(n4519), .B(n4520), .Z(n4237) );
  NOR U4428 ( .A(n4238), .B(n4237), .Z(n4515) );
  XOR U4429 ( .A(n4240), .B(n4239), .Z(n4516) );
  NOR U4430 ( .A(n4515), .B(n4516), .Z(n4241) );
  NOR U4431 ( .A(n4242), .B(n4241), .Z(n4511) );
  XOR U4432 ( .A(n4244), .B(n4243), .Z(n4512) );
  NOR U4433 ( .A(n4511), .B(n4512), .Z(n4245) );
  NOR U4434 ( .A(n4246), .B(n4245), .Z(n4507) );
  XOR U4435 ( .A(n4248), .B(n4247), .Z(n4508) );
  NOR U4436 ( .A(n4507), .B(n4508), .Z(n4249) );
  NOR U4437 ( .A(n4250), .B(n4249), .Z(n4503) );
  XOR U4438 ( .A(n4252), .B(n4251), .Z(n4504) );
  NOR U4439 ( .A(n4503), .B(n4504), .Z(n4253) );
  NOR U4440 ( .A(n4254), .B(n4253), .Z(n4499) );
  XOR U4441 ( .A(n4256), .B(n4255), .Z(n4500) );
  NOR U4442 ( .A(n4499), .B(n4500), .Z(n4257) );
  NOR U4443 ( .A(n4258), .B(n4257), .Z(n4495) );
  XOR U4444 ( .A(n4260), .B(n4259), .Z(n4496) );
  NOR U4445 ( .A(n4495), .B(n4496), .Z(n4261) );
  NOR U4446 ( .A(n4262), .B(n4261), .Z(n4491) );
  XOR U4447 ( .A(n4264), .B(n4263), .Z(n4492) );
  NOR U4448 ( .A(n4491), .B(n4492), .Z(n4265) );
  NOR U4449 ( .A(n4266), .B(n4265), .Z(n4487) );
  XOR U4450 ( .A(n4268), .B(n4267), .Z(n4488) );
  NOR U4451 ( .A(n4487), .B(n4488), .Z(n4269) );
  NOR U4452 ( .A(n4270), .B(n4269), .Z(n4483) );
  XOR U4453 ( .A(n4272), .B(n4271), .Z(n4484) );
  NOR U4454 ( .A(n4483), .B(n4484), .Z(n4273) );
  NOR U4455 ( .A(n4274), .B(n4273), .Z(n4479) );
  XOR U4456 ( .A(n4276), .B(n4275), .Z(n4480) );
  NOR U4457 ( .A(n4479), .B(n4480), .Z(n4277) );
  NOR U4458 ( .A(n4278), .B(n4277), .Z(n4475) );
  XOR U4459 ( .A(n4280), .B(n4279), .Z(n4476) );
  NOR U4460 ( .A(n4475), .B(n4476), .Z(n4281) );
  NOR U4461 ( .A(n4282), .B(n4281), .Z(n4471) );
  XOR U4462 ( .A(n4284), .B(n4283), .Z(n4472) );
  NOR U4463 ( .A(n4471), .B(n4472), .Z(n4285) );
  NOR U4464 ( .A(n4286), .B(n4285), .Z(n4467) );
  XOR U4465 ( .A(n4288), .B(n4287), .Z(n4468) );
  NOR U4466 ( .A(n4467), .B(n4468), .Z(n4289) );
  NOR U4467 ( .A(n4290), .B(n4289), .Z(n4463) );
  XOR U4468 ( .A(n4292), .B(n4291), .Z(n4464) );
  NOR U4469 ( .A(n4463), .B(n4464), .Z(n4293) );
  NOR U4470 ( .A(n4294), .B(n4293), .Z(n4459) );
  XOR U4471 ( .A(n4296), .B(n4295), .Z(n4460) );
  NOR U4472 ( .A(n4459), .B(n4460), .Z(n4297) );
  NOR U4473 ( .A(n4298), .B(n4297), .Z(n4455) );
  XOR U4474 ( .A(n4300), .B(n4299), .Z(n4456) );
  NOR U4475 ( .A(n4455), .B(n4456), .Z(n4301) );
  NOR U4476 ( .A(n4302), .B(n4301), .Z(n4451) );
  XOR U4477 ( .A(n4304), .B(n4303), .Z(n4452) );
  NOR U4478 ( .A(n4451), .B(n4452), .Z(n4305) );
  NOR U4479 ( .A(n4306), .B(n4305), .Z(n4311) );
  NOR U4480 ( .A(n109), .B(n129), .Z(n4310) );
  IV U4481 ( .A(n4310), .Z(n4307) );
  NOR U4482 ( .A(n4311), .B(n4307), .Z(n4314) );
  XOR U4483 ( .A(n4309), .B(n4308), .Z(n4449) );
  IV U4484 ( .A(n4449), .Z(n4312) );
  XOR U4485 ( .A(n4311), .B(n4310), .Z(n4448) );
  NOR U4486 ( .A(n4312), .B(n4448), .Z(n4313) );
  NOR U4487 ( .A(n4314), .B(n4313), .Z(n4447) );
  XOR U4488 ( .A(n4316), .B(n4315), .Z(n4446) );
  NOR U4489 ( .A(n4447), .B(n4446), .Z(n4317) );
  NOR U4490 ( .A(n4318), .B(n4317), .Z(n4445) );
  XOR U4491 ( .A(n4320), .B(n4319), .Z(n4444) );
  NOR U4492 ( .A(n4445), .B(n4444), .Z(n4321) );
  NOR U4493 ( .A(n4322), .B(n4321), .Z(n4443) );
  XOR U4494 ( .A(n4324), .B(n4323), .Z(n4442) );
  NOR U4495 ( .A(n4443), .B(n4442), .Z(n4325) );
  NOR U4496 ( .A(n4326), .B(n4325), .Z(n4331) );
  NOR U4497 ( .A(n85), .B(n129), .Z(n4330) );
  IV U4498 ( .A(n4330), .Z(n4327) );
  NOR U4499 ( .A(n4331), .B(n4327), .Z(n4333) );
  XOR U4500 ( .A(n4329), .B(n4328), .Z(n4441) );
  XOR U4501 ( .A(n4331), .B(n4330), .Z(n4440) );
  NOR U4502 ( .A(n4441), .B(n4440), .Z(n4332) );
  NOR U4503 ( .A(n4333), .B(n4332), .Z(n4338) );
  IV U4504 ( .A(n4338), .Z(n4336) );
  XOR U4505 ( .A(n4335), .B(n4334), .Z(n4337) );
  NOR U4506 ( .A(n4336), .B(n4337), .Z(n4340) );
  NOR U4507 ( .A(n112), .B(n129), .Z(n4438) );
  XOR U4508 ( .A(n4338), .B(n4337), .Z(n4437) );
  NOR U4509 ( .A(n4438), .B(n4437), .Z(n4339) );
  NOR U4510 ( .A(n4340), .B(n4339), .Z(n4341) );
  IV U4511 ( .A(n4341), .Z(n4436) );
  XOR U4512 ( .A(n4343), .B(n4342), .Z(n4435) );
  NOR U4513 ( .A(n4436), .B(n4435), .Z(n4344) );
  NOR U4514 ( .A(n4345), .B(n4344), .Z(n4347) );
  IV U4515 ( .A(n4347), .Z(n4346) );
  NOR U4516 ( .A(n4348), .B(n4346), .Z(n4350) );
  NOR U4517 ( .A(n113), .B(n129), .Z(n4433) );
  XOR U4518 ( .A(n4348), .B(n4347), .Z(n4432) );
  NOR U4519 ( .A(n4433), .B(n4432), .Z(n4349) );
  NOR U4520 ( .A(n4350), .B(n4349), .Z(n4428) );
  IV U4521 ( .A(n4428), .Z(n4353) );
  XOR U4522 ( .A(n4352), .B(n4351), .Z(n4427) );
  NOR U4523 ( .A(n4353), .B(n4427), .Z(n4354) );
  NOR U4524 ( .A(n4355), .B(n4354), .Z(n4424) );
  XOR U4525 ( .A(n4357), .B(n4356), .Z(n4423) );
  NOR U4526 ( .A(n4424), .B(n4423), .Z(n4358) );
  NOR U4527 ( .A(n4359), .B(n4358), .Z(n4419) );
  XOR U4528 ( .A(n4361), .B(n4360), .Z(n4420) );
  NOR U4529 ( .A(n4419), .B(n4420), .Z(n4362) );
  NOR U4530 ( .A(n4363), .B(n4362), .Z(n4415) );
  XOR U4531 ( .A(n4365), .B(n4364), .Z(n4416) );
  NOR U4532 ( .A(n4415), .B(n4416), .Z(n4366) );
  NOR U4533 ( .A(n4367), .B(n4366), .Z(n4369) );
  IV U4534 ( .A(n4369), .Z(n4368) );
  NOR U4535 ( .A(n4370), .B(n4368), .Z(n4374) );
  XOR U4536 ( .A(n4370), .B(n4369), .Z(n4412) );
  XOR U4537 ( .A(n4372), .B(n4371), .Z(n4413) );
  NOR U4538 ( .A(n4412), .B(n4413), .Z(n4373) );
  NOR U4539 ( .A(n4374), .B(n4373), .Z(n4375) );
  IV U4540 ( .A(n4375), .Z(n4411) );
  XOR U4541 ( .A(n4377), .B(n4376), .Z(n4410) );
  NOR U4542 ( .A(n4411), .B(n4410), .Z(n4378) );
  NOR U4543 ( .A(n4379), .B(n4378), .Z(n4409) );
  XOR U4544 ( .A(n4381), .B(n4380), .Z(n4408) );
  NOR U4545 ( .A(n4409), .B(n4408), .Z(n4382) );
  NOR U4546 ( .A(n4383), .B(n4382), .Z(n4388) );
  NOR U4547 ( .A(n117), .B(n129), .Z(n4387) );
  IV U4548 ( .A(n4387), .Z(n4384) );
  NOR U4549 ( .A(n4388), .B(n4384), .Z(n4390) );
  XOR U4550 ( .A(n4386), .B(n4385), .Z(n4407) );
  XOR U4551 ( .A(n4388), .B(n4387), .Z(n4406) );
  NOR U4552 ( .A(n4407), .B(n4406), .Z(n4389) );
  NOR U4553 ( .A(n4390), .B(n4389), .Z(n4405) );
  XOR U4554 ( .A(n4392), .B(n4391), .Z(n4404) );
  NOR U4555 ( .A(n4405), .B(n4404), .Z(n4393) );
  NOR U4556 ( .A(n4394), .B(n4393), .Z(n4399) );
  NOR U4557 ( .A(n119), .B(n129), .Z(n4398) );
  IV U4558 ( .A(n4398), .Z(n4395) );
  NOR U4559 ( .A(n4399), .B(n4395), .Z(n4401) );
  XOR U4560 ( .A(n4397), .B(n4396), .Z(n4403) );
  XOR U4561 ( .A(n4399), .B(n4398), .Z(n4402) );
  NOR U4562 ( .A(n4403), .B(n4402), .Z(n4400) );
  NOR U4563 ( .A(n4401), .B(n4400), .Z(n4712) );
  NOR U4564 ( .A(n120), .B(n129), .Z(n4710) );
  XOR U4565 ( .A(n4712), .B(n4710), .Z(n4713) );
  XOR U4566 ( .A(n4714), .B(n4713), .Z(n4705) );
  NOR U4567 ( .A(n4706), .B(n4705), .Z(n4709) );
  NOR U4568 ( .A(n120), .B(n127), .Z(n4700) );
  XOR U4569 ( .A(n4403), .B(n4402), .Z(n4701) );
  NOR U4570 ( .A(n4700), .B(n4701), .Z(n4704) );
  NOR U4571 ( .A(n119), .B(n127), .Z(n4696) );
  XOR U4572 ( .A(n4405), .B(n4404), .Z(n4695) );
  NOR U4573 ( .A(n4696), .B(n4695), .Z(n4699) );
  NOR U4574 ( .A(n79), .B(n127), .Z(n4691) );
  XOR U4575 ( .A(n4407), .B(n4406), .Z(n4690) );
  NOR U4576 ( .A(n4691), .B(n4690), .Z(n4694) );
  NOR U4577 ( .A(n117), .B(n127), .Z(n4685) );
  XOR U4578 ( .A(n4409), .B(n4408), .Z(n4686) );
  NOR U4579 ( .A(n4685), .B(n4686), .Z(n4689) );
  NOR U4580 ( .A(n80), .B(n127), .Z(n4681) );
  XOR U4581 ( .A(n4411), .B(n4410), .Z(n4680) );
  NOR U4582 ( .A(n4681), .B(n4680), .Z(n4684) );
  NOR U4583 ( .A(n116), .B(n127), .Z(n4677) );
  XOR U4584 ( .A(n4413), .B(n4412), .Z(n4676) );
  IV U4585 ( .A(n4676), .Z(n4414) );
  NOR U4586 ( .A(n4677), .B(n4414), .Z(n4679) );
  IV U4587 ( .A(n4415), .Z(n4417) );
  XOR U4588 ( .A(n4417), .B(n4416), .Z(n4671) );
  NOR U4589 ( .A(n81), .B(n127), .Z(n4672) );
  IV U4590 ( .A(n4672), .Z(n4418) );
  NOR U4591 ( .A(n4671), .B(n4418), .Z(n4674) );
  IV U4592 ( .A(n4419), .Z(n4421) );
  XOR U4593 ( .A(n4421), .B(n4420), .Z(n4667) );
  NOR U4594 ( .A(n115), .B(n127), .Z(n4668) );
  IV U4595 ( .A(n4668), .Z(n4422) );
  NOR U4596 ( .A(n4667), .B(n4422), .Z(n4670) );
  XOR U4597 ( .A(n4424), .B(n4423), .Z(n4663) );
  IV U4598 ( .A(n4663), .Z(n4426) );
  NOR U4599 ( .A(n82), .B(n127), .Z(n4425) );
  IV U4600 ( .A(n4425), .Z(n4664) );
  NOR U4601 ( .A(n4426), .B(n4664), .Z(n4666) );
  XOR U4602 ( .A(n4428), .B(n4427), .Z(n4430) );
  NOR U4603 ( .A(n114), .B(n127), .Z(n4431) );
  IV U4604 ( .A(n4431), .Z(n4429) );
  NOR U4605 ( .A(n4430), .B(n4429), .Z(n4662) );
  XOR U4606 ( .A(n4431), .B(n4430), .Z(n4859) );
  NOR U4607 ( .A(n83), .B(n127), .Z(n4657) );
  XOR U4608 ( .A(n4433), .B(n4432), .Z(n4656) );
  IV U4609 ( .A(n4656), .Z(n4434) );
  NOR U4610 ( .A(n4657), .B(n4434), .Z(n4659) );
  NOR U4611 ( .A(n113), .B(n127), .Z(n4651) );
  XOR U4612 ( .A(n4436), .B(n4435), .Z(n4652) );
  NOR U4613 ( .A(n4651), .B(n4652), .Z(n4655) );
  NOR U4614 ( .A(n84), .B(n127), .Z(n4648) );
  XOR U4615 ( .A(n4438), .B(n4437), .Z(n4647) );
  IV U4616 ( .A(n4647), .Z(n4439) );
  NOR U4617 ( .A(n4648), .B(n4439), .Z(n4650) );
  NOR U4618 ( .A(n112), .B(n127), .Z(n4643) );
  XOR U4619 ( .A(n4441), .B(n4440), .Z(n4642) );
  NOR U4620 ( .A(n4643), .B(n4642), .Z(n4646) );
  NOR U4621 ( .A(n85), .B(n127), .Z(n4638) );
  XOR U4622 ( .A(n4443), .B(n4442), .Z(n4637) );
  NOR U4623 ( .A(n4638), .B(n4637), .Z(n4641) );
  NOR U4624 ( .A(n111), .B(n127), .Z(n4633) );
  XOR U4625 ( .A(n4445), .B(n4444), .Z(n4632) );
  NOR U4626 ( .A(n4633), .B(n4632), .Z(n4636) );
  NOR U4627 ( .A(n86), .B(n127), .Z(n4628) );
  XOR U4628 ( .A(n4447), .B(n4446), .Z(n4627) );
  NOR U4629 ( .A(n4628), .B(n4627), .Z(n4631) );
  XOR U4630 ( .A(n4449), .B(n4448), .Z(n4622) );
  NOR U4631 ( .A(n110), .B(n127), .Z(n4623) );
  IV U4632 ( .A(n4623), .Z(n4450) );
  NOR U4633 ( .A(n4622), .B(n4450), .Z(n4625) );
  IV U4634 ( .A(n4451), .Z(n4453) );
  XOR U4635 ( .A(n4453), .B(n4452), .Z(n4618) );
  NOR U4636 ( .A(n109), .B(n127), .Z(n4619) );
  IV U4637 ( .A(n4619), .Z(n4454) );
  NOR U4638 ( .A(n4618), .B(n4454), .Z(n4621) );
  XOR U4639 ( .A(n4456), .B(n4455), .Z(n4457) );
  IV U4640 ( .A(n4457), .Z(n4614) );
  NOR U4641 ( .A(n108), .B(n127), .Z(n4615) );
  IV U4642 ( .A(n4615), .Z(n4458) );
  NOR U4643 ( .A(n4614), .B(n4458), .Z(n4617) );
  XOR U4644 ( .A(n4460), .B(n4459), .Z(n4461) );
  IV U4645 ( .A(n4461), .Z(n4610) );
  NOR U4646 ( .A(n87), .B(n127), .Z(n4611) );
  IV U4647 ( .A(n4611), .Z(n4462) );
  NOR U4648 ( .A(n4610), .B(n4462), .Z(n4613) );
  XOR U4649 ( .A(n4464), .B(n4463), .Z(n4465) );
  IV U4650 ( .A(n4465), .Z(n4606) );
  NOR U4651 ( .A(n107), .B(n127), .Z(n4607) );
  IV U4652 ( .A(n4607), .Z(n4466) );
  NOR U4653 ( .A(n4606), .B(n4466), .Z(n4609) );
  XOR U4654 ( .A(n4468), .B(n4467), .Z(n4469) );
  IV U4655 ( .A(n4469), .Z(n4602) );
  NOR U4656 ( .A(n88), .B(n127), .Z(n4603) );
  IV U4657 ( .A(n4603), .Z(n4470) );
  NOR U4658 ( .A(n4602), .B(n4470), .Z(n4605) );
  XOR U4659 ( .A(n4472), .B(n4471), .Z(n4473) );
  IV U4660 ( .A(n4473), .Z(n4598) );
  NOR U4661 ( .A(n106), .B(n127), .Z(n4599) );
  IV U4662 ( .A(n4599), .Z(n4474) );
  NOR U4663 ( .A(n4598), .B(n4474), .Z(n4601) );
  XOR U4664 ( .A(n4476), .B(n4475), .Z(n4477) );
  IV U4665 ( .A(n4477), .Z(n4594) );
  NOR U4666 ( .A(n105), .B(n127), .Z(n4595) );
  IV U4667 ( .A(n4595), .Z(n4478) );
  NOR U4668 ( .A(n4594), .B(n4478), .Z(n4597) );
  XOR U4669 ( .A(n4480), .B(n4479), .Z(n4481) );
  IV U4670 ( .A(n4481), .Z(n4590) );
  NOR U4671 ( .A(n104), .B(n127), .Z(n4591) );
  IV U4672 ( .A(n4591), .Z(n4482) );
  NOR U4673 ( .A(n4590), .B(n4482), .Z(n4593) );
  XOR U4674 ( .A(n4484), .B(n4483), .Z(n4485) );
  IV U4675 ( .A(n4485), .Z(n4586) );
  NOR U4676 ( .A(n89), .B(n127), .Z(n4587) );
  IV U4677 ( .A(n4587), .Z(n4486) );
  NOR U4678 ( .A(n4586), .B(n4486), .Z(n4589) );
  XOR U4679 ( .A(n4488), .B(n4487), .Z(n4489) );
  IV U4680 ( .A(n4489), .Z(n4582) );
  NOR U4681 ( .A(n103), .B(n127), .Z(n4583) );
  IV U4682 ( .A(n4583), .Z(n4490) );
  NOR U4683 ( .A(n4582), .B(n4490), .Z(n4585) );
  XOR U4684 ( .A(n4492), .B(n4491), .Z(n4493) );
  IV U4685 ( .A(n4493), .Z(n4578) );
  NOR U4686 ( .A(n90), .B(n127), .Z(n4579) );
  IV U4687 ( .A(n4579), .Z(n4494) );
  NOR U4688 ( .A(n4578), .B(n4494), .Z(n4581) );
  IV U4689 ( .A(n4495), .Z(n4497) );
  XOR U4690 ( .A(n4497), .B(n4496), .Z(n4574) );
  NOR U4691 ( .A(n102), .B(n127), .Z(n4575) );
  IV U4692 ( .A(n4575), .Z(n4498) );
  NOR U4693 ( .A(n4574), .B(n4498), .Z(n4577) );
  XOR U4694 ( .A(n4500), .B(n4499), .Z(n4501) );
  IV U4695 ( .A(n4501), .Z(n4570) );
  NOR U4696 ( .A(n101), .B(n127), .Z(n4571) );
  IV U4697 ( .A(n4571), .Z(n4502) );
  NOR U4698 ( .A(n4570), .B(n4502), .Z(n4573) );
  XOR U4699 ( .A(n4504), .B(n4503), .Z(n4505) );
  IV U4700 ( .A(n4505), .Z(n4566) );
  NOR U4701 ( .A(n100), .B(n127), .Z(n4567) );
  IV U4702 ( .A(n4567), .Z(n4506) );
  NOR U4703 ( .A(n4566), .B(n4506), .Z(n4569) );
  XOR U4704 ( .A(n4508), .B(n4507), .Z(n4509) );
  IV U4705 ( .A(n4509), .Z(n4562) );
  NOR U4706 ( .A(n99), .B(n127), .Z(n4563) );
  IV U4707 ( .A(n4563), .Z(n4510) );
  NOR U4708 ( .A(n4562), .B(n4510), .Z(n4565) );
  XOR U4709 ( .A(n4512), .B(n4511), .Z(n4513) );
  IV U4710 ( .A(n4513), .Z(n4558) );
  NOR U4711 ( .A(n98), .B(n127), .Z(n4559) );
  IV U4712 ( .A(n4559), .Z(n4514) );
  NOR U4713 ( .A(n4558), .B(n4514), .Z(n4561) );
  IV U4714 ( .A(n4515), .Z(n4517) );
  XOR U4715 ( .A(n4517), .B(n4516), .Z(n4554) );
  NOR U4716 ( .A(n91), .B(n127), .Z(n4555) );
  IV U4717 ( .A(n4555), .Z(n4518) );
  NOR U4718 ( .A(n4554), .B(n4518), .Z(n4557) );
  IV U4719 ( .A(n4519), .Z(n4521) );
  XOR U4720 ( .A(n4521), .B(n4520), .Z(n4550) );
  NOR U4721 ( .A(n97), .B(n127), .Z(n4551) );
  IV U4722 ( .A(n4551), .Z(n4522) );
  NOR U4723 ( .A(n4550), .B(n4522), .Z(n4553) );
  NOR U4724 ( .A(n96), .B(n127), .Z(n4547) );
  IV U4725 ( .A(n4547), .Z(n4526) );
  XOR U4726 ( .A(n4524), .B(n4523), .Z(n4525) );
  IV U4727 ( .A(n4525), .Z(n4546) );
  NOR U4728 ( .A(n4526), .B(n4546), .Z(n4549) );
  NOR U4729 ( .A(n93), .B(n127), .Z(n5446) );
  IV U4730 ( .A(n5446), .Z(n4528) );
  NOR U4731 ( .A(n129), .B(n168), .Z(n4531) );
  IV U4732 ( .A(n4531), .Z(n4527) );
  NOR U4733 ( .A(n4528), .B(n4527), .Z(n4966) );
  IV U4734 ( .A(n4966), .Z(n4529) );
  NOR U4735 ( .A(n4530), .B(n4529), .Z(n4538) );
  XOR U4736 ( .A(n4532), .B(n4531), .Z(n4533) );
  NOR U4737 ( .A(n4966), .B(n4533), .Z(n4534) );
  NOR U4738 ( .A(n4538), .B(n4534), .Z(n4535) );
  IV U4739 ( .A(n4535), .Z(n4979) );
  NOR U4740 ( .A(n94), .B(n127), .Z(n4978) );
  IV U4741 ( .A(n4978), .Z(n4536) );
  NOR U4742 ( .A(n4979), .B(n4536), .Z(n4537) );
  NOR U4743 ( .A(n4538), .B(n4537), .Z(n4541) );
  NOR U4744 ( .A(n95), .B(n127), .Z(n4540) );
  IV U4745 ( .A(n4540), .Z(n4539) );
  NOR U4746 ( .A(n4541), .B(n4539), .Z(n4545) );
  XOR U4747 ( .A(n4541), .B(n4540), .Z(n4959) );
  XOR U4748 ( .A(n4543), .B(n4542), .Z(n4960) );
  NOR U4749 ( .A(n4959), .B(n4960), .Z(n4544) );
  NOR U4750 ( .A(n4545), .B(n4544), .Z(n4956) );
  XOR U4751 ( .A(n4547), .B(n4546), .Z(n4955) );
  NOR U4752 ( .A(n4956), .B(n4955), .Z(n4548) );
  NOR U4753 ( .A(n4549), .B(n4548), .Z(n4951) );
  XOR U4754 ( .A(n4551), .B(n4550), .Z(n4952) );
  NOR U4755 ( .A(n4951), .B(n4952), .Z(n4552) );
  NOR U4756 ( .A(n4553), .B(n4552), .Z(n4948) );
  XOR U4757 ( .A(n4555), .B(n4554), .Z(n4947) );
  NOR U4758 ( .A(n4948), .B(n4947), .Z(n4556) );
  NOR U4759 ( .A(n4557), .B(n4556), .Z(n4943) );
  XOR U4760 ( .A(n4559), .B(n4558), .Z(n4944) );
  NOR U4761 ( .A(n4943), .B(n4944), .Z(n4560) );
  NOR U4762 ( .A(n4561), .B(n4560), .Z(n4939) );
  XOR U4763 ( .A(n4563), .B(n4562), .Z(n4940) );
  NOR U4764 ( .A(n4939), .B(n4940), .Z(n4564) );
  NOR U4765 ( .A(n4565), .B(n4564), .Z(n4935) );
  XOR U4766 ( .A(n4567), .B(n4566), .Z(n4936) );
  NOR U4767 ( .A(n4935), .B(n4936), .Z(n4568) );
  NOR U4768 ( .A(n4569), .B(n4568), .Z(n4931) );
  XOR U4769 ( .A(n4571), .B(n4570), .Z(n4932) );
  NOR U4770 ( .A(n4931), .B(n4932), .Z(n4572) );
  NOR U4771 ( .A(n4573), .B(n4572), .Z(n4927) );
  XOR U4772 ( .A(n4575), .B(n4574), .Z(n4928) );
  NOR U4773 ( .A(n4927), .B(n4928), .Z(n4576) );
  NOR U4774 ( .A(n4577), .B(n4576), .Z(n4923) );
  XOR U4775 ( .A(n4579), .B(n4578), .Z(n4924) );
  NOR U4776 ( .A(n4923), .B(n4924), .Z(n4580) );
  NOR U4777 ( .A(n4581), .B(n4580), .Z(n4919) );
  XOR U4778 ( .A(n4583), .B(n4582), .Z(n4920) );
  NOR U4779 ( .A(n4919), .B(n4920), .Z(n4584) );
  NOR U4780 ( .A(n4585), .B(n4584), .Z(n4915) );
  XOR U4781 ( .A(n4587), .B(n4586), .Z(n4916) );
  NOR U4782 ( .A(n4915), .B(n4916), .Z(n4588) );
  NOR U4783 ( .A(n4589), .B(n4588), .Z(n4911) );
  XOR U4784 ( .A(n4591), .B(n4590), .Z(n4912) );
  NOR U4785 ( .A(n4911), .B(n4912), .Z(n4592) );
  NOR U4786 ( .A(n4593), .B(n4592), .Z(n4907) );
  XOR U4787 ( .A(n4595), .B(n4594), .Z(n4908) );
  NOR U4788 ( .A(n4907), .B(n4908), .Z(n4596) );
  NOR U4789 ( .A(n4597), .B(n4596), .Z(n4903) );
  XOR U4790 ( .A(n4599), .B(n4598), .Z(n4904) );
  NOR U4791 ( .A(n4903), .B(n4904), .Z(n4600) );
  NOR U4792 ( .A(n4601), .B(n4600), .Z(n4899) );
  XOR U4793 ( .A(n4603), .B(n4602), .Z(n4900) );
  NOR U4794 ( .A(n4899), .B(n4900), .Z(n4604) );
  NOR U4795 ( .A(n4605), .B(n4604), .Z(n4895) );
  XOR U4796 ( .A(n4607), .B(n4606), .Z(n4896) );
  NOR U4797 ( .A(n4895), .B(n4896), .Z(n4608) );
  NOR U4798 ( .A(n4609), .B(n4608), .Z(n4891) );
  XOR U4799 ( .A(n4611), .B(n4610), .Z(n4892) );
  NOR U4800 ( .A(n4891), .B(n4892), .Z(n4612) );
  NOR U4801 ( .A(n4613), .B(n4612), .Z(n4887) );
  XOR U4802 ( .A(n4615), .B(n4614), .Z(n4888) );
  NOR U4803 ( .A(n4887), .B(n4888), .Z(n4616) );
  NOR U4804 ( .A(n4617), .B(n4616), .Z(n4883) );
  XOR U4805 ( .A(n4619), .B(n4618), .Z(n4884) );
  NOR U4806 ( .A(n4883), .B(n4884), .Z(n4620) );
  NOR U4807 ( .A(n4621), .B(n4620), .Z(n4879) );
  XOR U4808 ( .A(n4623), .B(n4622), .Z(n4880) );
  NOR U4809 ( .A(n4879), .B(n4880), .Z(n4624) );
  NOR U4810 ( .A(n4625), .B(n4624), .Z(n4626) );
  IV U4811 ( .A(n4626), .Z(n4877) );
  XOR U4812 ( .A(n4628), .B(n4627), .Z(n4629) );
  IV U4813 ( .A(n4629), .Z(n4876) );
  NOR U4814 ( .A(n4877), .B(n4876), .Z(n4630) );
  NOR U4815 ( .A(n4631), .B(n4630), .Z(n4874) );
  XOR U4816 ( .A(n4633), .B(n4632), .Z(n4634) );
  IV U4817 ( .A(n4634), .Z(n4873) );
  NOR U4818 ( .A(n4874), .B(n4873), .Z(n4635) );
  NOR U4819 ( .A(n4636), .B(n4635), .Z(n4871) );
  XOR U4820 ( .A(n4638), .B(n4637), .Z(n4639) );
  IV U4821 ( .A(n4639), .Z(n4870) );
  NOR U4822 ( .A(n4871), .B(n4870), .Z(n4640) );
  NOR U4823 ( .A(n4641), .B(n4640), .Z(n4868) );
  XOR U4824 ( .A(n4643), .B(n4642), .Z(n4644) );
  IV U4825 ( .A(n4644), .Z(n4867) );
  NOR U4826 ( .A(n4868), .B(n4867), .Z(n4645) );
  NOR U4827 ( .A(n4646), .B(n4645), .Z(n4866) );
  XOR U4828 ( .A(n4648), .B(n4647), .Z(n4865) );
  NOR U4829 ( .A(n4866), .B(n4865), .Z(n4649) );
  NOR U4830 ( .A(n4650), .B(n4649), .Z(n4863) );
  IV U4831 ( .A(n4651), .Z(n4653) );
  XOR U4832 ( .A(n4653), .B(n4652), .Z(n4862) );
  NOR U4833 ( .A(n4863), .B(n4862), .Z(n4654) );
  NOR U4834 ( .A(n4655), .B(n4654), .Z(n5094) );
  XOR U4835 ( .A(n4657), .B(n4656), .Z(n5093) );
  NOR U4836 ( .A(n5094), .B(n5093), .Z(n4658) );
  NOR U4837 ( .A(n4659), .B(n4658), .Z(n4860) );
  IV U4838 ( .A(n4860), .Z(n4660) );
  NOR U4839 ( .A(n4859), .B(n4660), .Z(n4661) );
  NOR U4840 ( .A(n4662), .B(n4661), .Z(n5107) );
  XOR U4841 ( .A(n4664), .B(n4663), .Z(n5106) );
  NOR U4842 ( .A(n5107), .B(n5106), .Z(n4665) );
  NOR U4843 ( .A(n4666), .B(n4665), .Z(n4855) );
  XOR U4844 ( .A(n4668), .B(n4667), .Z(n4854) );
  NOR U4845 ( .A(n4855), .B(n4854), .Z(n4669) );
  NOR U4846 ( .A(n4670), .B(n4669), .Z(n4850) );
  XOR U4847 ( .A(n4672), .B(n4671), .Z(n4851) );
  NOR U4848 ( .A(n4850), .B(n4851), .Z(n4673) );
  NOR U4849 ( .A(n4674), .B(n4673), .Z(n4675) );
  IV U4850 ( .A(n4675), .Z(n5121) );
  XOR U4851 ( .A(n4677), .B(n4676), .Z(n5120) );
  NOR U4852 ( .A(n5121), .B(n5120), .Z(n4678) );
  NOR U4853 ( .A(n4679), .B(n4678), .Z(n5130) );
  XOR U4854 ( .A(n4681), .B(n4680), .Z(n5129) );
  IV U4855 ( .A(n5129), .Z(n4682) );
  NOR U4856 ( .A(n5130), .B(n4682), .Z(n4683) );
  NOR U4857 ( .A(n4684), .B(n4683), .Z(n5136) );
  IV U4858 ( .A(n4685), .Z(n4687) );
  XOR U4859 ( .A(n4687), .B(n4686), .Z(n5135) );
  NOR U4860 ( .A(n5136), .B(n5135), .Z(n4688) );
  NOR U4861 ( .A(n4689), .B(n4688), .Z(n5143) );
  XOR U4862 ( .A(n4691), .B(n4690), .Z(n4692) );
  IV U4863 ( .A(n4692), .Z(n5142) );
  NOR U4864 ( .A(n5143), .B(n5142), .Z(n4693) );
  NOR U4865 ( .A(n4694), .B(n4693), .Z(n5150) );
  XOR U4866 ( .A(n4696), .B(n4695), .Z(n4697) );
  IV U4867 ( .A(n4697), .Z(n5149) );
  NOR U4868 ( .A(n5150), .B(n5149), .Z(n4698) );
  NOR U4869 ( .A(n4699), .B(n4698), .Z(n4849) );
  IV U4870 ( .A(n4700), .Z(n4702) );
  XOR U4871 ( .A(n4702), .B(n4701), .Z(n4848) );
  NOR U4872 ( .A(n4849), .B(n4848), .Z(n4703) );
  NOR U4873 ( .A(n4704), .B(n4703), .Z(n5163) );
  XOR U4874 ( .A(n4706), .B(n4705), .Z(n4707) );
  IV U4875 ( .A(n4707), .Z(n5162) );
  NOR U4876 ( .A(n5163), .B(n5162), .Z(n4708) );
  NOR U4877 ( .A(n4709), .B(n4708), .Z(n5177) );
  NOR U4878 ( .A(n125), .B(n127), .Z(n5175) );
  IV U4879 ( .A(n5175), .Z(n4847) );
  IV U4880 ( .A(n4710), .Z(n4711) );
  NOR U4881 ( .A(n4712), .B(n4711), .Z(n4716) );
  NOR U4882 ( .A(n4714), .B(n4713), .Z(n4715) );
  NOR U4883 ( .A(n4716), .B(n4715), .Z(n5311) );
  IV U4884 ( .A(n5311), .Z(n4845) );
  NOR U4885 ( .A(n4718), .B(n4717), .Z(n4722) );
  NOR U4886 ( .A(n4720), .B(n4719), .Z(n4721) );
  NOR U4887 ( .A(n4722), .B(n4721), .Z(n5183) );
  NOR U4888 ( .A(n120), .B(n130), .Z(n5181) );
  IV U4889 ( .A(n5181), .Z(n4844) );
  NOR U4890 ( .A(n4724), .B(n4723), .Z(n4728) );
  NOR U4891 ( .A(n4726), .B(n4725), .Z(n4727) );
  NOR U4892 ( .A(n4728), .B(n4727), .Z(n5196) );
  NOR U4893 ( .A(n79), .B(n134), .Z(n5194) );
  NOR U4894 ( .A(n4730), .B(n4729), .Z(n4734) );
  NOR U4895 ( .A(n4732), .B(n4731), .Z(n4733) );
  NOR U4896 ( .A(n4734), .B(n4733), .Z(n5210) );
  NOR U4897 ( .A(n80), .B(n138), .Z(n5208) );
  NOR U4898 ( .A(n4736), .B(n4735), .Z(n4740) );
  NOR U4899 ( .A(n4738), .B(n4737), .Z(n4739) );
  NOR U4900 ( .A(n4740), .B(n4739), .Z(n5217) );
  NOR U4901 ( .A(n81), .B(n142), .Z(n5214) );
  IV U4902 ( .A(n4741), .Z(n4742) );
  NOR U4903 ( .A(n4743), .B(n4742), .Z(n4747) );
  NOR U4904 ( .A(n4745), .B(n4744), .Z(n4746) );
  NOR U4905 ( .A(n4747), .B(n4746), .Z(n5223) );
  NOR U4906 ( .A(n82), .B(n146), .Z(n5221) );
  IV U4907 ( .A(n5221), .Z(n4814) );
  NOR U4908 ( .A(n4749), .B(n4748), .Z(n4754) );
  IV U4909 ( .A(n4750), .Z(n4751) );
  NOR U4910 ( .A(n4752), .B(n4751), .Z(n4753) );
  NOR U4911 ( .A(n4754), .B(n4753), .Z(n5236) );
  NOR U4912 ( .A(n83), .B(n151), .Z(n5234) );
  IV U4913 ( .A(n4755), .Z(n4756) );
  NOR U4914 ( .A(n4757), .B(n4756), .Z(n4761) );
  NOR U4915 ( .A(n4759), .B(n4758), .Z(n4760) );
  NOR U4916 ( .A(n4761), .B(n4760), .Z(n5243) );
  NOR U4917 ( .A(n4763), .B(n4762), .Z(n4767) );
  NOR U4918 ( .A(n4765), .B(n4764), .Z(n4766) );
  NOR U4919 ( .A(n4767), .B(n4766), .Z(n5249) );
  NOR U4920 ( .A(n84), .B(n154), .Z(n5247) );
  NOR U4921 ( .A(n4769), .B(n4768), .Z(n4773) );
  NOR U4922 ( .A(n4771), .B(n4770), .Z(n4772) );
  NOR U4923 ( .A(n4773), .B(n4772), .Z(n5262) );
  NOR U4924 ( .A(n85), .B(n159), .Z(n5260) );
  NOR U4925 ( .A(n4775), .B(n4774), .Z(n4779) );
  NOR U4926 ( .A(n4777), .B(n4776), .Z(n4778) );
  NOR U4927 ( .A(n4779), .B(n4778), .Z(n5275) );
  NOR U4928 ( .A(n86), .B(n162), .Z(n5273) );
  IV U4929 ( .A(n5273), .Z(n4788) );
  IV U4930 ( .A(n4780), .Z(n4781) );
  NOR U4931 ( .A(n4782), .B(n4781), .Z(n4786) );
  NOR U4932 ( .A(n4784), .B(n4783), .Z(n4785) );
  NOR U4933 ( .A(n4786), .B(n4785), .Z(n5280) );
  NOR U4934 ( .A(n164), .B(n110), .Z(n5278) );
  XOR U4935 ( .A(n5280), .B(n5278), .Z(n5282) );
  NOR U4936 ( .A(n166), .B(n109), .Z(n4787) );
  IV U4937 ( .A(n4787), .Z(n5281) );
  XOR U4938 ( .A(n5282), .B(n5281), .Z(n5272) );
  XOR U4939 ( .A(n4788), .B(n5272), .Z(n5274) );
  XOR U4940 ( .A(n5275), .B(n5274), .Z(n5269) );
  IV U4941 ( .A(n4789), .Z(n4790) );
  NOR U4942 ( .A(n4791), .B(n4790), .Z(n4795) );
  NOR U4943 ( .A(n4793), .B(n4792), .Z(n4794) );
  NOR U4944 ( .A(n4795), .B(n4794), .Z(n5267) );
  NOR U4945 ( .A(n111), .B(n160), .Z(n5265) );
  XOR U4946 ( .A(n5267), .B(n5265), .Z(n5268) );
  XOR U4947 ( .A(n5269), .B(n5268), .Z(n5259) );
  XOR U4948 ( .A(n5260), .B(n5259), .Z(n4796) );
  IV U4949 ( .A(n4796), .Z(n5261) );
  XOR U4950 ( .A(n5262), .B(n5261), .Z(n5256) );
  IV U4951 ( .A(n4797), .Z(n4798) );
  NOR U4952 ( .A(n4799), .B(n4798), .Z(n4803) );
  NOR U4953 ( .A(n4801), .B(n4800), .Z(n4802) );
  NOR U4954 ( .A(n4803), .B(n4802), .Z(n5254) );
  NOR U4955 ( .A(n112), .B(n157), .Z(n5252) );
  XOR U4956 ( .A(n5254), .B(n5252), .Z(n5255) );
  XOR U4957 ( .A(n5256), .B(n5255), .Z(n5246) );
  XOR U4958 ( .A(n5247), .B(n5246), .Z(n4804) );
  IV U4959 ( .A(n4804), .Z(n5248) );
  XOR U4960 ( .A(n5249), .B(n5248), .Z(n5241) );
  NOR U4961 ( .A(n113), .B(n152), .Z(n5239) );
  XOR U4962 ( .A(n5241), .B(n5239), .Z(n5242) );
  XOR U4963 ( .A(n5243), .B(n5242), .Z(n5233) );
  XOR U4964 ( .A(n5234), .B(n5233), .Z(n4805) );
  IV U4965 ( .A(n4805), .Z(n5235) );
  XOR U4966 ( .A(n5236), .B(n5235), .Z(n5228) );
  IV U4967 ( .A(n4806), .Z(n4807) );
  NOR U4968 ( .A(n4808), .B(n4807), .Z(n4812) );
  NOR U4969 ( .A(n4810), .B(n4809), .Z(n4811) );
  NOR U4970 ( .A(n4812), .B(n4811), .Z(n5226) );
  XOR U4971 ( .A(n5228), .B(n5226), .Z(n5230) );
  NOR U4972 ( .A(n114), .B(n149), .Z(n4813) );
  IV U4973 ( .A(n4813), .Z(n5229) );
  XOR U4974 ( .A(n5230), .B(n5229), .Z(n5220) );
  XOR U4975 ( .A(n4814), .B(n5220), .Z(n5222) );
  XOR U4976 ( .A(n5223), .B(n5222), .Z(n5297) );
  IV U4977 ( .A(n4815), .Z(n4816) );
  NOR U4978 ( .A(n4817), .B(n4816), .Z(n4821) );
  NOR U4979 ( .A(n4819), .B(n4818), .Z(n4820) );
  NOR U4980 ( .A(n4821), .B(n4820), .Z(n5295) );
  NOR U4981 ( .A(n115), .B(n144), .Z(n5293) );
  XOR U4982 ( .A(n5295), .B(n5293), .Z(n5296) );
  XOR U4983 ( .A(n5297), .B(n5296), .Z(n5213) );
  XOR U4984 ( .A(n5214), .B(n5213), .Z(n5215) );
  XOR U4985 ( .A(n5217), .B(n5215), .Z(n5304) );
  NOR U4986 ( .A(n116), .B(n140), .Z(n5303) );
  IV U4987 ( .A(n4822), .Z(n4823) );
  NOR U4988 ( .A(n4824), .B(n4823), .Z(n4828) );
  NOR U4989 ( .A(n4826), .B(n4825), .Z(n4827) );
  NOR U4990 ( .A(n4828), .B(n4827), .Z(n5301) );
  XOR U4991 ( .A(n5303), .B(n5301), .Z(n5305) );
  XOR U4992 ( .A(n5304), .B(n5305), .Z(n5206) );
  XOR U4993 ( .A(n5208), .B(n5206), .Z(n5209) );
  XOR U4994 ( .A(n5210), .B(n5209), .Z(n5203) );
  IV U4995 ( .A(n4829), .Z(n4830) );
  NOR U4996 ( .A(n4831), .B(n4830), .Z(n4835) );
  NOR U4997 ( .A(n4833), .B(n4832), .Z(n4834) );
  NOR U4998 ( .A(n4835), .B(n4834), .Z(n5201) );
  NOR U4999 ( .A(n117), .B(n136), .Z(n5199) );
  XOR U5000 ( .A(n5201), .B(n5199), .Z(n5202) );
  XOR U5001 ( .A(n5203), .B(n5202), .Z(n5193) );
  XOR U5002 ( .A(n5194), .B(n5193), .Z(n4836) );
  IV U5003 ( .A(n4836), .Z(n5195) );
  XOR U5004 ( .A(n5196), .B(n5195), .Z(n5190) );
  IV U5005 ( .A(n4837), .Z(n4838) );
  NOR U5006 ( .A(n4839), .B(n4838), .Z(n4843) );
  NOR U5007 ( .A(n4841), .B(n4840), .Z(n4842) );
  NOR U5008 ( .A(n4843), .B(n4842), .Z(n5188) );
  NOR U5009 ( .A(n119), .B(n132), .Z(n5186) );
  XOR U5010 ( .A(n5188), .B(n5186), .Z(n5189) );
  XOR U5011 ( .A(n5190), .B(n5189), .Z(n5180) );
  XOR U5012 ( .A(n4844), .B(n5180), .Z(n5182) );
  XOR U5013 ( .A(n5183), .B(n5182), .Z(n5312) );
  XOR U5014 ( .A(n4845), .B(n5312), .Z(n5314) );
  NOR U5015 ( .A(n123), .B(n129), .Z(n4846) );
  IV U5016 ( .A(n4846), .Z(n5313) );
  XOR U5017 ( .A(n5314), .B(n5313), .Z(n5174) );
  XOR U5018 ( .A(n4847), .B(n5174), .Z(n5176) );
  XOR U5019 ( .A(n5177), .B(n5176), .Z(n5169) );
  XOR U5020 ( .A(n4849), .B(n4848), .Z(n5156) );
  NOR U5021 ( .A(n117), .B(n124), .Z(n5128) );
  IV U5022 ( .A(n4850), .Z(n4852) );
  XOR U5023 ( .A(n4852), .B(n4851), .Z(n5114) );
  NOR U5024 ( .A(n116), .B(n124), .Z(n5115) );
  IV U5025 ( .A(n5115), .Z(n4853) );
  NOR U5026 ( .A(n5114), .B(n4853), .Z(n5118) );
  NOR U5027 ( .A(n81), .B(n124), .Z(n4857) );
  XOR U5028 ( .A(n4855), .B(n4854), .Z(n4856) );
  NOR U5029 ( .A(n4857), .B(n4856), .Z(n5113) );
  XOR U5030 ( .A(n4857), .B(n4856), .Z(n4858) );
  IV U5031 ( .A(n4858), .Z(n5340) );
  XOR U5032 ( .A(n4860), .B(n4859), .Z(n5099) );
  NOR U5033 ( .A(n82), .B(n124), .Z(n5100) );
  IV U5034 ( .A(n5100), .Z(n4861) );
  NOR U5035 ( .A(n5099), .B(n4861), .Z(n5102) );
  XOR U5036 ( .A(n4863), .B(n4862), .Z(n5089) );
  NOR U5037 ( .A(n83), .B(n124), .Z(n5088) );
  IV U5038 ( .A(n5088), .Z(n4864) );
  NOR U5039 ( .A(n5089), .B(n4864), .Z(n5091) );
  XOR U5040 ( .A(n4866), .B(n4865), .Z(n5083) );
  XOR U5041 ( .A(n4868), .B(n4867), .Z(n5079) );
  NOR U5042 ( .A(n84), .B(n124), .Z(n5078) );
  IV U5043 ( .A(n5078), .Z(n4869) );
  NOR U5044 ( .A(n5079), .B(n4869), .Z(n5081) );
  XOR U5045 ( .A(n4871), .B(n4870), .Z(n5075) );
  NOR U5046 ( .A(n112), .B(n124), .Z(n5074) );
  IV U5047 ( .A(n5074), .Z(n4872) );
  NOR U5048 ( .A(n5075), .B(n4872), .Z(n5077) );
  XOR U5049 ( .A(n4874), .B(n4873), .Z(n5071) );
  NOR U5050 ( .A(n85), .B(n124), .Z(n5070) );
  IV U5051 ( .A(n5070), .Z(n4875) );
  NOR U5052 ( .A(n5071), .B(n4875), .Z(n5073) );
  XOR U5053 ( .A(n4877), .B(n4876), .Z(n5067) );
  NOR U5054 ( .A(n111), .B(n124), .Z(n5066) );
  IV U5055 ( .A(n5066), .Z(n4878) );
  NOR U5056 ( .A(n5067), .B(n4878), .Z(n5069) );
  IV U5057 ( .A(n4879), .Z(n4881) );
  XOR U5058 ( .A(n4881), .B(n4880), .Z(n5062) );
  NOR U5059 ( .A(n86), .B(n124), .Z(n5063) );
  IV U5060 ( .A(n5063), .Z(n4882) );
  NOR U5061 ( .A(n5062), .B(n4882), .Z(n5065) );
  IV U5062 ( .A(n4883), .Z(n4885) );
  XOR U5063 ( .A(n4885), .B(n4884), .Z(n5058) );
  NOR U5064 ( .A(n110), .B(n124), .Z(n5059) );
  IV U5065 ( .A(n5059), .Z(n4886) );
  NOR U5066 ( .A(n5058), .B(n4886), .Z(n5061) );
  XOR U5067 ( .A(n4888), .B(n4887), .Z(n4889) );
  IV U5068 ( .A(n4889), .Z(n5054) );
  NOR U5069 ( .A(n109), .B(n124), .Z(n5055) );
  IV U5070 ( .A(n5055), .Z(n4890) );
  NOR U5071 ( .A(n5054), .B(n4890), .Z(n5057) );
  XOR U5072 ( .A(n4892), .B(n4891), .Z(n4893) );
  IV U5073 ( .A(n4893), .Z(n5050) );
  NOR U5074 ( .A(n108), .B(n124), .Z(n5051) );
  IV U5075 ( .A(n5051), .Z(n4894) );
  NOR U5076 ( .A(n5050), .B(n4894), .Z(n5053) );
  XOR U5077 ( .A(n4896), .B(n4895), .Z(n4897) );
  IV U5078 ( .A(n4897), .Z(n5046) );
  NOR U5079 ( .A(n87), .B(n124), .Z(n5047) );
  IV U5080 ( .A(n5047), .Z(n4898) );
  NOR U5081 ( .A(n5046), .B(n4898), .Z(n5049) );
  IV U5082 ( .A(n4899), .Z(n4901) );
  XOR U5083 ( .A(n4901), .B(n4900), .Z(n5042) );
  NOR U5084 ( .A(n107), .B(n124), .Z(n5043) );
  IV U5085 ( .A(n5043), .Z(n4902) );
  NOR U5086 ( .A(n5042), .B(n4902), .Z(n5045) );
  XOR U5087 ( .A(n4904), .B(n4903), .Z(n4905) );
  IV U5088 ( .A(n4905), .Z(n5038) );
  NOR U5089 ( .A(n88), .B(n124), .Z(n5039) );
  IV U5090 ( .A(n5039), .Z(n4906) );
  NOR U5091 ( .A(n5038), .B(n4906), .Z(n5041) );
  XOR U5092 ( .A(n4908), .B(n4907), .Z(n4909) );
  IV U5093 ( .A(n4909), .Z(n5034) );
  NOR U5094 ( .A(n106), .B(n124), .Z(n5035) );
  IV U5095 ( .A(n5035), .Z(n4910) );
  NOR U5096 ( .A(n5034), .B(n4910), .Z(n5037) );
  XOR U5097 ( .A(n4912), .B(n4911), .Z(n4913) );
  IV U5098 ( .A(n4913), .Z(n5030) );
  NOR U5099 ( .A(n105), .B(n124), .Z(n5031) );
  IV U5100 ( .A(n5031), .Z(n4914) );
  NOR U5101 ( .A(n5030), .B(n4914), .Z(n5033) );
  XOR U5102 ( .A(n4916), .B(n4915), .Z(n4917) );
  IV U5103 ( .A(n4917), .Z(n5026) );
  NOR U5104 ( .A(n104), .B(n124), .Z(n5027) );
  IV U5105 ( .A(n5027), .Z(n4918) );
  NOR U5106 ( .A(n5026), .B(n4918), .Z(n5029) );
  XOR U5107 ( .A(n4920), .B(n4919), .Z(n4921) );
  IV U5108 ( .A(n4921), .Z(n5022) );
  NOR U5109 ( .A(n89), .B(n124), .Z(n5023) );
  IV U5110 ( .A(n5023), .Z(n4922) );
  NOR U5111 ( .A(n5022), .B(n4922), .Z(n5025) );
  XOR U5112 ( .A(n4924), .B(n4923), .Z(n4925) );
  IV U5113 ( .A(n4925), .Z(n5018) );
  NOR U5114 ( .A(n103), .B(n124), .Z(n5019) );
  IV U5115 ( .A(n5019), .Z(n4926) );
  NOR U5116 ( .A(n5018), .B(n4926), .Z(n5021) );
  XOR U5117 ( .A(n4928), .B(n4927), .Z(n4929) );
  IV U5118 ( .A(n4929), .Z(n5014) );
  NOR U5119 ( .A(n90), .B(n124), .Z(n5015) );
  IV U5120 ( .A(n5015), .Z(n4930) );
  NOR U5121 ( .A(n5014), .B(n4930), .Z(n5017) );
  XOR U5122 ( .A(n4932), .B(n4931), .Z(n4933) );
  IV U5123 ( .A(n4933), .Z(n5010) );
  NOR U5124 ( .A(n102), .B(n124), .Z(n5011) );
  IV U5125 ( .A(n5011), .Z(n4934) );
  NOR U5126 ( .A(n5010), .B(n4934), .Z(n5013) );
  XOR U5127 ( .A(n4936), .B(n4935), .Z(n4937) );
  IV U5128 ( .A(n4937), .Z(n5006) );
  NOR U5129 ( .A(n101), .B(n124), .Z(n5007) );
  IV U5130 ( .A(n5007), .Z(n4938) );
  NOR U5131 ( .A(n5006), .B(n4938), .Z(n5009) );
  XOR U5132 ( .A(n4940), .B(n4939), .Z(n4941) );
  IV U5133 ( .A(n4941), .Z(n5002) );
  NOR U5134 ( .A(n100), .B(n124), .Z(n5003) );
  IV U5135 ( .A(n5003), .Z(n4942) );
  NOR U5136 ( .A(n5002), .B(n4942), .Z(n5005) );
  IV U5137 ( .A(n4943), .Z(n4945) );
  XOR U5138 ( .A(n4945), .B(n4944), .Z(n4998) );
  NOR U5139 ( .A(n99), .B(n124), .Z(n4999) );
  IV U5140 ( .A(n4999), .Z(n4946) );
  NOR U5141 ( .A(n4998), .B(n4946), .Z(n5001) );
  XOR U5142 ( .A(n4948), .B(n4947), .Z(n4994) );
  IV U5143 ( .A(n4994), .Z(n4950) );
  NOR U5144 ( .A(n98), .B(n124), .Z(n4949) );
  IV U5145 ( .A(n4949), .Z(n4995) );
  NOR U5146 ( .A(n4950), .B(n4995), .Z(n4997) );
  IV U5147 ( .A(n4951), .Z(n4953) );
  XOR U5148 ( .A(n4953), .B(n4952), .Z(n4990) );
  NOR U5149 ( .A(n91), .B(n124), .Z(n4991) );
  IV U5150 ( .A(n4991), .Z(n4954) );
  NOR U5151 ( .A(n4990), .B(n4954), .Z(n4993) );
  IV U5152 ( .A(n4955), .Z(n4957) );
  XOR U5153 ( .A(n4957), .B(n4956), .Z(n4986) );
  NOR U5154 ( .A(n97), .B(n124), .Z(n4987) );
  IV U5155 ( .A(n4987), .Z(n4958) );
  NOR U5156 ( .A(n4986), .B(n4958), .Z(n4989) );
  NOR U5157 ( .A(n96), .B(n124), .Z(n4983) );
  IV U5158 ( .A(n4983), .Z(n4962) );
  XOR U5159 ( .A(n4960), .B(n4959), .Z(n4961) );
  IV U5160 ( .A(n4961), .Z(n4982) );
  NOR U5161 ( .A(n4962), .B(n4982), .Z(n4985) );
  NOR U5162 ( .A(n93), .B(n124), .Z(n5962) );
  IV U5163 ( .A(n5962), .Z(n4964) );
  NOR U5164 ( .A(n127), .B(n168), .Z(n4967) );
  IV U5165 ( .A(n4967), .Z(n4963) );
  NOR U5166 ( .A(n4964), .B(n4963), .Z(n5444) );
  IV U5167 ( .A(n5444), .Z(n4965) );
  NOR U5168 ( .A(n4966), .B(n4965), .Z(n4974) );
  XOR U5169 ( .A(n4968), .B(n4967), .Z(n4969) );
  NOR U5170 ( .A(n5444), .B(n4969), .Z(n4970) );
  NOR U5171 ( .A(n4974), .B(n4970), .Z(n4971) );
  IV U5172 ( .A(n4971), .Z(n5457) );
  NOR U5173 ( .A(n94), .B(n124), .Z(n5456) );
  IV U5174 ( .A(n5456), .Z(n4972) );
  NOR U5175 ( .A(n5457), .B(n4972), .Z(n4973) );
  NOR U5176 ( .A(n4974), .B(n4973), .Z(n4977) );
  NOR U5177 ( .A(n95), .B(n124), .Z(n4976) );
  IV U5178 ( .A(n4976), .Z(n4975) );
  NOR U5179 ( .A(n4977), .B(n4975), .Z(n4981) );
  XOR U5180 ( .A(n4977), .B(n4976), .Z(n5437) );
  XOR U5181 ( .A(n4979), .B(n4978), .Z(n5438) );
  NOR U5182 ( .A(n5437), .B(n5438), .Z(n4980) );
  NOR U5183 ( .A(n4981), .B(n4980), .Z(n5433) );
  XOR U5184 ( .A(n4983), .B(n4982), .Z(n5434) );
  NOR U5185 ( .A(n5433), .B(n5434), .Z(n4984) );
  NOR U5186 ( .A(n4985), .B(n4984), .Z(n5432) );
  XOR U5187 ( .A(n4987), .B(n4986), .Z(n5431) );
  NOR U5188 ( .A(n5432), .B(n5431), .Z(n4988) );
  NOR U5189 ( .A(n4989), .B(n4988), .Z(n5474) );
  XOR U5190 ( .A(n4991), .B(n4990), .Z(n5475) );
  NOR U5191 ( .A(n5474), .B(n5475), .Z(n4992) );
  NOR U5192 ( .A(n4993), .B(n4992), .Z(n5430) );
  XOR U5193 ( .A(n4995), .B(n4994), .Z(n5429) );
  NOR U5194 ( .A(n5430), .B(n5429), .Z(n4996) );
  NOR U5195 ( .A(n4997), .B(n4996), .Z(n5487) );
  XOR U5196 ( .A(n4999), .B(n4998), .Z(n5488) );
  NOR U5197 ( .A(n5487), .B(n5488), .Z(n5000) );
  NOR U5198 ( .A(n5001), .B(n5000), .Z(n5425) );
  XOR U5199 ( .A(n5003), .B(n5002), .Z(n5426) );
  NOR U5200 ( .A(n5425), .B(n5426), .Z(n5004) );
  NOR U5201 ( .A(n5005), .B(n5004), .Z(n5421) );
  XOR U5202 ( .A(n5007), .B(n5006), .Z(n5422) );
  NOR U5203 ( .A(n5421), .B(n5422), .Z(n5008) );
  NOR U5204 ( .A(n5009), .B(n5008), .Z(n5417) );
  XOR U5205 ( .A(n5011), .B(n5010), .Z(n5418) );
  NOR U5206 ( .A(n5417), .B(n5418), .Z(n5012) );
  NOR U5207 ( .A(n5013), .B(n5012), .Z(n5413) );
  XOR U5208 ( .A(n5015), .B(n5014), .Z(n5414) );
  NOR U5209 ( .A(n5413), .B(n5414), .Z(n5016) );
  NOR U5210 ( .A(n5017), .B(n5016), .Z(n5409) );
  XOR U5211 ( .A(n5019), .B(n5018), .Z(n5410) );
  NOR U5212 ( .A(n5409), .B(n5410), .Z(n5020) );
  NOR U5213 ( .A(n5021), .B(n5020), .Z(n5405) );
  XOR U5214 ( .A(n5023), .B(n5022), .Z(n5406) );
  NOR U5215 ( .A(n5405), .B(n5406), .Z(n5024) );
  NOR U5216 ( .A(n5025), .B(n5024), .Z(n5401) );
  XOR U5217 ( .A(n5027), .B(n5026), .Z(n5402) );
  NOR U5218 ( .A(n5401), .B(n5402), .Z(n5028) );
  NOR U5219 ( .A(n5029), .B(n5028), .Z(n5397) );
  XOR U5220 ( .A(n5031), .B(n5030), .Z(n5398) );
  NOR U5221 ( .A(n5397), .B(n5398), .Z(n5032) );
  NOR U5222 ( .A(n5033), .B(n5032), .Z(n5393) );
  XOR U5223 ( .A(n5035), .B(n5034), .Z(n5394) );
  NOR U5224 ( .A(n5393), .B(n5394), .Z(n5036) );
  NOR U5225 ( .A(n5037), .B(n5036), .Z(n5389) );
  XOR U5226 ( .A(n5039), .B(n5038), .Z(n5390) );
  NOR U5227 ( .A(n5389), .B(n5390), .Z(n5040) );
  NOR U5228 ( .A(n5041), .B(n5040), .Z(n5385) );
  XOR U5229 ( .A(n5043), .B(n5042), .Z(n5386) );
  NOR U5230 ( .A(n5385), .B(n5386), .Z(n5044) );
  NOR U5231 ( .A(n5045), .B(n5044), .Z(n5381) );
  XOR U5232 ( .A(n5047), .B(n5046), .Z(n5382) );
  NOR U5233 ( .A(n5381), .B(n5382), .Z(n5048) );
  NOR U5234 ( .A(n5049), .B(n5048), .Z(n5377) );
  XOR U5235 ( .A(n5051), .B(n5050), .Z(n5378) );
  NOR U5236 ( .A(n5377), .B(n5378), .Z(n5052) );
  NOR U5237 ( .A(n5053), .B(n5052), .Z(n5373) );
  XOR U5238 ( .A(n5055), .B(n5054), .Z(n5374) );
  NOR U5239 ( .A(n5373), .B(n5374), .Z(n5056) );
  NOR U5240 ( .A(n5057), .B(n5056), .Z(n5369) );
  XOR U5241 ( .A(n5059), .B(n5058), .Z(n5370) );
  NOR U5242 ( .A(n5369), .B(n5370), .Z(n5060) );
  NOR U5243 ( .A(n5061), .B(n5060), .Z(n5365) );
  XOR U5244 ( .A(n5063), .B(n5062), .Z(n5366) );
  NOR U5245 ( .A(n5365), .B(n5366), .Z(n5064) );
  NOR U5246 ( .A(n5065), .B(n5064), .Z(n5361) );
  XOR U5247 ( .A(n5067), .B(n5066), .Z(n5362) );
  NOR U5248 ( .A(n5361), .B(n5362), .Z(n5068) );
  NOR U5249 ( .A(n5069), .B(n5068), .Z(n5360) );
  XOR U5250 ( .A(n5071), .B(n5070), .Z(n5359) );
  NOR U5251 ( .A(n5360), .B(n5359), .Z(n5072) );
  NOR U5252 ( .A(n5073), .B(n5072), .Z(n5358) );
  XOR U5253 ( .A(n5075), .B(n5074), .Z(n5357) );
  NOR U5254 ( .A(n5358), .B(n5357), .Z(n5076) );
  NOR U5255 ( .A(n5077), .B(n5076), .Z(n5356) );
  XOR U5256 ( .A(n5079), .B(n5078), .Z(n5355) );
  NOR U5257 ( .A(n5356), .B(n5355), .Z(n5080) );
  NOR U5258 ( .A(n5081), .B(n5080), .Z(n5082) );
  NOR U5259 ( .A(n5083), .B(n5082), .Z(n5087) );
  IV U5260 ( .A(n5082), .Z(n5084) );
  XOR U5261 ( .A(n5084), .B(n5083), .Z(n5354) );
  NOR U5262 ( .A(n113), .B(n124), .Z(n5085) );
  IV U5263 ( .A(n5085), .Z(n5353) );
  NOR U5264 ( .A(n5354), .B(n5353), .Z(n5086) );
  NOR U5265 ( .A(n5087), .B(n5086), .Z(n5352) );
  XOR U5266 ( .A(n5089), .B(n5088), .Z(n5351) );
  NOR U5267 ( .A(n5352), .B(n5351), .Z(n5090) );
  NOR U5268 ( .A(n5091), .B(n5090), .Z(n5096) );
  NOR U5269 ( .A(n114), .B(n124), .Z(n5095) );
  IV U5270 ( .A(n5095), .Z(n5092) );
  NOR U5271 ( .A(n5096), .B(n5092), .Z(n5098) );
  XOR U5272 ( .A(n5094), .B(n5093), .Z(n5350) );
  XOR U5273 ( .A(n5096), .B(n5095), .Z(n5349) );
  NOR U5274 ( .A(n5350), .B(n5349), .Z(n5097) );
  NOR U5275 ( .A(n5098), .B(n5097), .Z(n5348) );
  XOR U5276 ( .A(n5100), .B(n5099), .Z(n5347) );
  NOR U5277 ( .A(n5348), .B(n5347), .Z(n5101) );
  NOR U5278 ( .A(n5102), .B(n5101), .Z(n5105) );
  NOR U5279 ( .A(n115), .B(n124), .Z(n5104) );
  IV U5280 ( .A(n5104), .Z(n5103) );
  NOR U5281 ( .A(n5105), .B(n5103), .Z(n5110) );
  XOR U5282 ( .A(n5105), .B(n5104), .Z(n5342) );
  XOR U5283 ( .A(n5107), .B(n5106), .Z(n5343) );
  IV U5284 ( .A(n5343), .Z(n5108) );
  NOR U5285 ( .A(n5342), .B(n5108), .Z(n5109) );
  NOR U5286 ( .A(n5110), .B(n5109), .Z(n5111) );
  IV U5287 ( .A(n5111), .Z(n5339) );
  NOR U5288 ( .A(n5340), .B(n5339), .Z(n5112) );
  NOR U5289 ( .A(n5113), .B(n5112), .Z(n5337) );
  IV U5290 ( .A(n5337), .Z(n5116) );
  XOR U5291 ( .A(n5115), .B(n5114), .Z(n5336) );
  NOR U5292 ( .A(n5116), .B(n5336), .Z(n5117) );
  NOR U5293 ( .A(n5118), .B(n5117), .Z(n5123) );
  NOR U5294 ( .A(n80), .B(n124), .Z(n5122) );
  IV U5295 ( .A(n5122), .Z(n5119) );
  NOR U5296 ( .A(n5123), .B(n5119), .Z(n5125) );
  XOR U5297 ( .A(n5121), .B(n5120), .Z(n5335) );
  XOR U5298 ( .A(n5123), .B(n5122), .Z(n5334) );
  NOR U5299 ( .A(n5335), .B(n5334), .Z(n5124) );
  NOR U5300 ( .A(n5125), .B(n5124), .Z(n5127) );
  IV U5301 ( .A(n5127), .Z(n5126) );
  NOR U5302 ( .A(n5128), .B(n5126), .Z(n5132) );
  XOR U5303 ( .A(n5128), .B(n5127), .Z(n5331) );
  XOR U5304 ( .A(n5130), .B(n5129), .Z(n5332) );
  NOR U5305 ( .A(n5331), .B(n5332), .Z(n5131) );
  NOR U5306 ( .A(n5132), .B(n5131), .Z(n5133) );
  IV U5307 ( .A(n5133), .Z(n5138) );
  NOR U5308 ( .A(n79), .B(n124), .Z(n5137) );
  IV U5309 ( .A(n5137), .Z(n5134) );
  NOR U5310 ( .A(n5138), .B(n5134), .Z(n5140) );
  XOR U5311 ( .A(n5136), .B(n5135), .Z(n5329) );
  XOR U5312 ( .A(n5138), .B(n5137), .Z(n5330) );
  NOR U5313 ( .A(n5329), .B(n5330), .Z(n5139) );
  NOR U5314 ( .A(n5140), .B(n5139), .Z(n5145) );
  NOR U5315 ( .A(n119), .B(n124), .Z(n5144) );
  IV U5316 ( .A(n5144), .Z(n5141) );
  NOR U5317 ( .A(n5145), .B(n5141), .Z(n5147) );
  XOR U5318 ( .A(n5143), .B(n5142), .Z(n5328) );
  XOR U5319 ( .A(n5145), .B(n5144), .Z(n5327) );
  NOR U5320 ( .A(n5328), .B(n5327), .Z(n5146) );
  NOR U5321 ( .A(n5147), .B(n5146), .Z(n5152) );
  NOR U5322 ( .A(n120), .B(n124), .Z(n5151) );
  IV U5323 ( .A(n5151), .Z(n5148) );
  NOR U5324 ( .A(n5152), .B(n5148), .Z(n5154) );
  XOR U5325 ( .A(n5150), .B(n5149), .Z(n5326) );
  XOR U5326 ( .A(n5152), .B(n5151), .Z(n5325) );
  NOR U5327 ( .A(n5326), .B(n5325), .Z(n5153) );
  NOR U5328 ( .A(n5154), .B(n5153), .Z(n5155) );
  NOR U5329 ( .A(n5156), .B(n5155), .Z(n5160) );
  IV U5330 ( .A(n5155), .Z(n5157) );
  XOR U5331 ( .A(n5157), .B(n5156), .Z(n5324) );
  NOR U5332 ( .A(n123), .B(n124), .Z(n5158) );
  IV U5333 ( .A(n5158), .Z(n5323) );
  NOR U5334 ( .A(n5324), .B(n5323), .Z(n5159) );
  NOR U5335 ( .A(n5160), .B(n5159), .Z(n5165) );
  NOR U5336 ( .A(n125), .B(n124), .Z(n5164) );
  IV U5337 ( .A(n5164), .Z(n5161) );
  NOR U5338 ( .A(n5165), .B(n5161), .Z(n5167) );
  XOR U5339 ( .A(n5163), .B(n5162), .Z(n5322) );
  XOR U5340 ( .A(n5165), .B(n5164), .Z(n5321) );
  NOR U5341 ( .A(n5322), .B(n5321), .Z(n5166) );
  NOR U5342 ( .A(n5167), .B(n5166), .Z(n5168) );
  NOR U5343 ( .A(n5169), .B(n5168), .Z(n5173) );
  IV U5344 ( .A(n5168), .Z(n5170) );
  XOR U5345 ( .A(n5170), .B(n5169), .Z(n5320) );
  NOR U5346 ( .A(n126), .B(n124), .Z(n5171) );
  IV U5347 ( .A(n5171), .Z(n5319) );
  NOR U5348 ( .A(n5320), .B(n5319), .Z(n5172) );
  NOR U5349 ( .A(n5173), .B(n5172), .Z(n5655) );
  IV U5350 ( .A(n5655), .Z(n5317) );
  NOR U5351 ( .A(n5175), .B(n5174), .Z(n5179) );
  NOR U5352 ( .A(n5177), .B(n5176), .Z(n5178) );
  NOR U5353 ( .A(n5179), .B(n5178), .Z(n5665) );
  NOR U5354 ( .A(n126), .B(n127), .Z(n5663) );
  NOR U5355 ( .A(n5181), .B(n5180), .Z(n5185) );
  NOR U5356 ( .A(n5183), .B(n5182), .Z(n5184) );
  NOR U5357 ( .A(n5185), .B(n5184), .Z(n5680) );
  NOR U5358 ( .A(n123), .B(n130), .Z(n5677) );
  IV U5359 ( .A(n5186), .Z(n5187) );
  NOR U5360 ( .A(n5188), .B(n5187), .Z(n5192) );
  NOR U5361 ( .A(n5190), .B(n5189), .Z(n5191) );
  NOR U5362 ( .A(n5192), .B(n5191), .Z(n5683) );
  NOR U5363 ( .A(n5194), .B(n5193), .Z(n5198) );
  NOR U5364 ( .A(n5196), .B(n5195), .Z(n5197) );
  NOR U5365 ( .A(n5198), .B(n5197), .Z(n5694) );
  NOR U5366 ( .A(n119), .B(n134), .Z(n5692) );
  IV U5367 ( .A(n5692), .Z(n5310) );
  IV U5368 ( .A(n5199), .Z(n5200) );
  NOR U5369 ( .A(n5201), .B(n5200), .Z(n5205) );
  NOR U5370 ( .A(n5203), .B(n5202), .Z(n5204) );
  NOR U5371 ( .A(n5205), .B(n5204), .Z(n5701) );
  IV U5372 ( .A(n5206), .Z(n5207) );
  NOR U5373 ( .A(n5208), .B(n5207), .Z(n5212) );
  NOR U5374 ( .A(n5210), .B(n5209), .Z(n5211) );
  NOR U5375 ( .A(n5212), .B(n5211), .Z(n5707) );
  NOR U5376 ( .A(n117), .B(n138), .Z(n5705) );
  IV U5377 ( .A(n5705), .Z(n5309) );
  NOR U5378 ( .A(n5214), .B(n5213), .Z(n5219) );
  IV U5379 ( .A(n5215), .Z(n5216) );
  NOR U5380 ( .A(n5217), .B(n5216), .Z(n5218) );
  NOR U5381 ( .A(n5219), .B(n5218), .Z(n5720) );
  NOR U5382 ( .A(n116), .B(n142), .Z(n5718) );
  NOR U5383 ( .A(n5221), .B(n5220), .Z(n5225) );
  NOR U5384 ( .A(n5223), .B(n5222), .Z(n5224) );
  NOR U5385 ( .A(n5225), .B(n5224), .Z(n5727) );
  NOR U5386 ( .A(n115), .B(n146), .Z(n5725) );
  NOR U5387 ( .A(n82), .B(n149), .Z(n5793) );
  IV U5388 ( .A(n5226), .Z(n5227) );
  NOR U5389 ( .A(n5228), .B(n5227), .Z(n5232) );
  NOR U5390 ( .A(n5230), .B(n5229), .Z(n5231) );
  NOR U5391 ( .A(n5232), .B(n5231), .Z(n5789) );
  NOR U5392 ( .A(n5234), .B(n5233), .Z(n5238) );
  NOR U5393 ( .A(n5236), .B(n5235), .Z(n5237) );
  NOR U5394 ( .A(n5238), .B(n5237), .Z(n5734) );
  NOR U5395 ( .A(n114), .B(n151), .Z(n5731) );
  IV U5396 ( .A(n5239), .Z(n5240) );
  NOR U5397 ( .A(n5241), .B(n5240), .Z(n5245) );
  NOR U5398 ( .A(n5243), .B(n5242), .Z(n5244) );
  NOR U5399 ( .A(n5245), .B(n5244), .Z(n5737) );
  NOR U5400 ( .A(n5247), .B(n5246), .Z(n5251) );
  NOR U5401 ( .A(n5249), .B(n5248), .Z(n5250) );
  NOR U5402 ( .A(n5251), .B(n5250), .Z(n5748) );
  NOR U5403 ( .A(n113), .B(n154), .Z(n5746) );
  IV U5404 ( .A(n5746), .Z(n5292) );
  IV U5405 ( .A(n5252), .Z(n5253) );
  NOR U5406 ( .A(n5254), .B(n5253), .Z(n5258) );
  NOR U5407 ( .A(n5256), .B(n5255), .Z(n5257) );
  NOR U5408 ( .A(n5258), .B(n5257), .Z(n5751) );
  IV U5409 ( .A(n5751), .Z(n5290) );
  NOR U5410 ( .A(n5260), .B(n5259), .Z(n5264) );
  NOR U5411 ( .A(n5262), .B(n5261), .Z(n5263) );
  NOR U5412 ( .A(n5264), .B(n5263), .Z(n5760) );
  NOR U5413 ( .A(n112), .B(n159), .Z(n5758) );
  IV U5414 ( .A(n5758), .Z(n5289) );
  IV U5415 ( .A(n5265), .Z(n5266) );
  NOR U5416 ( .A(n5267), .B(n5266), .Z(n5271) );
  NOR U5417 ( .A(n5269), .B(n5268), .Z(n5270) );
  NOR U5418 ( .A(n5271), .B(n5270), .Z(n5778) );
  IV U5419 ( .A(n5778), .Z(n5287) );
  NOR U5420 ( .A(n5273), .B(n5272), .Z(n5277) );
  NOR U5421 ( .A(n5275), .B(n5274), .Z(n5276) );
  NOR U5422 ( .A(n5277), .B(n5276), .Z(n5766) );
  NOR U5423 ( .A(n111), .B(n162), .Z(n5764) );
  IV U5424 ( .A(n5764), .Z(n5286) );
  IV U5425 ( .A(n5278), .Z(n5279) );
  NOR U5426 ( .A(n5280), .B(n5279), .Z(n5284) );
  NOR U5427 ( .A(n5282), .B(n5281), .Z(n5283) );
  NOR U5428 ( .A(n5284), .B(n5283), .Z(n5771) );
  NOR U5429 ( .A(n164), .B(n86), .Z(n5769) );
  XOR U5430 ( .A(n5771), .B(n5769), .Z(n5773) );
  NOR U5431 ( .A(n166), .B(n110), .Z(n5285) );
  IV U5432 ( .A(n5285), .Z(n5772) );
  XOR U5433 ( .A(n5773), .B(n5772), .Z(n5763) );
  XOR U5434 ( .A(n5286), .B(n5763), .Z(n5765) );
  XOR U5435 ( .A(n5766), .B(n5765), .Z(n5779) );
  XOR U5436 ( .A(n5287), .B(n5779), .Z(n5781) );
  NOR U5437 ( .A(n85), .B(n160), .Z(n5288) );
  IV U5438 ( .A(n5288), .Z(n5780) );
  XOR U5439 ( .A(n5781), .B(n5780), .Z(n5757) );
  XOR U5440 ( .A(n5289), .B(n5757), .Z(n5759) );
  XOR U5441 ( .A(n5760), .B(n5759), .Z(n5752) );
  XOR U5442 ( .A(n5290), .B(n5752), .Z(n5754) );
  NOR U5443 ( .A(n84), .B(n157), .Z(n5291) );
  IV U5444 ( .A(n5291), .Z(n5753) );
  XOR U5445 ( .A(n5754), .B(n5753), .Z(n5745) );
  XOR U5446 ( .A(n5292), .B(n5745), .Z(n5747) );
  XOR U5447 ( .A(n5748), .B(n5747), .Z(n5738) );
  XOR U5448 ( .A(n5737), .B(n5738), .Z(n5739) );
  NOR U5449 ( .A(n83), .B(n152), .Z(n5740) );
  XOR U5450 ( .A(n5739), .B(n5740), .Z(n5730) );
  XOR U5451 ( .A(n5731), .B(n5730), .Z(n5732) );
  XOR U5452 ( .A(n5734), .B(n5732), .Z(n5790) );
  XOR U5453 ( .A(n5789), .B(n5790), .Z(n5792) );
  XOR U5454 ( .A(n5793), .B(n5792), .Z(n5723) );
  XOR U5455 ( .A(n5725), .B(n5723), .Z(n5726) );
  XOR U5456 ( .A(n5727), .B(n5726), .Z(n5802) );
  IV U5457 ( .A(n5293), .Z(n5294) );
  NOR U5458 ( .A(n5295), .B(n5294), .Z(n5299) );
  NOR U5459 ( .A(n5297), .B(n5296), .Z(n5298) );
  NOR U5460 ( .A(n5299), .B(n5298), .Z(n5800) );
  NOR U5461 ( .A(n81), .B(n144), .Z(n5798) );
  XOR U5462 ( .A(n5800), .B(n5798), .Z(n5801) );
  XOR U5463 ( .A(n5802), .B(n5801), .Z(n5717) );
  XOR U5464 ( .A(n5718), .B(n5717), .Z(n5300) );
  IV U5465 ( .A(n5300), .Z(n5719) );
  XOR U5466 ( .A(n5720), .B(n5719), .Z(n5712) );
  IV U5467 ( .A(n5301), .Z(n5302) );
  NOR U5468 ( .A(n5303), .B(n5302), .Z(n5307) );
  NOR U5469 ( .A(n5305), .B(n5304), .Z(n5306) );
  NOR U5470 ( .A(n5307), .B(n5306), .Z(n5710) );
  XOR U5471 ( .A(n5712), .B(n5710), .Z(n5714) );
  NOR U5472 ( .A(n80), .B(n140), .Z(n5308) );
  IV U5473 ( .A(n5308), .Z(n5713) );
  XOR U5474 ( .A(n5714), .B(n5713), .Z(n5704) );
  XOR U5475 ( .A(n5309), .B(n5704), .Z(n5706) );
  XOR U5476 ( .A(n5707), .B(n5706), .Z(n5699) );
  NOR U5477 ( .A(n79), .B(n136), .Z(n5697) );
  XOR U5478 ( .A(n5699), .B(n5697), .Z(n5700) );
  XOR U5479 ( .A(n5701), .B(n5700), .Z(n5691) );
  XOR U5480 ( .A(n5310), .B(n5691), .Z(n5693) );
  XOR U5481 ( .A(n5694), .B(n5693), .Z(n5684) );
  XOR U5482 ( .A(n5683), .B(n5684), .Z(n5685) );
  NOR U5483 ( .A(n120), .B(n132), .Z(n5686) );
  XOR U5484 ( .A(n5685), .B(n5686), .Z(n5676) );
  XOR U5485 ( .A(n5677), .B(n5676), .Z(n5678) );
  XOR U5486 ( .A(n5680), .B(n5678), .Z(n5671) );
  NOR U5487 ( .A(n125), .B(n129), .Z(n5670) );
  NOR U5488 ( .A(n5312), .B(n5311), .Z(n5316) );
  NOR U5489 ( .A(n5314), .B(n5313), .Z(n5315) );
  NOR U5490 ( .A(n5316), .B(n5315), .Z(n5668) );
  XOR U5491 ( .A(n5670), .B(n5668), .Z(n5672) );
  XOR U5492 ( .A(n5671), .B(n5672), .Z(n5661) );
  XOR U5493 ( .A(n5663), .B(n5661), .Z(n5664) );
  XOR U5494 ( .A(n5665), .B(n5664), .Z(n5656) );
  XOR U5495 ( .A(n5317), .B(n5656), .Z(n5658) );
  NOR U5496 ( .A(n128), .B(n124), .Z(n5318) );
  IV U5497 ( .A(n5318), .Z(n5657) );
  XOR U5498 ( .A(n5658), .B(n5657), .Z(n5650) );
  NOR U5499 ( .A(n5649), .B(n5650), .Z(n5653) );
  NOR U5500 ( .A(n128), .B(n122), .Z(n5644) );
  XOR U5501 ( .A(n5320), .B(n5319), .Z(n5645) );
  NOR U5502 ( .A(n5644), .B(n5645), .Z(n5648) );
  NOR U5503 ( .A(n126), .B(n122), .Z(n5640) );
  XOR U5504 ( .A(n5322), .B(n5321), .Z(n5639) );
  NOR U5505 ( .A(n5640), .B(n5639), .Z(n5643) );
  NOR U5506 ( .A(n125), .B(n122), .Z(n5634) );
  XOR U5507 ( .A(n5324), .B(n5323), .Z(n5635) );
  NOR U5508 ( .A(n5634), .B(n5635), .Z(n5638) );
  NOR U5509 ( .A(n123), .B(n122), .Z(n5630) );
  XOR U5510 ( .A(n5326), .B(n5325), .Z(n5629) );
  NOR U5511 ( .A(n5630), .B(n5629), .Z(n5633) );
  NOR U5512 ( .A(n120), .B(n122), .Z(n5625) );
  XOR U5513 ( .A(n5328), .B(n5327), .Z(n5624) );
  NOR U5514 ( .A(n5625), .B(n5624), .Z(n5628) );
  NOR U5515 ( .A(n119), .B(n122), .Z(n5619) );
  XOR U5516 ( .A(n5330), .B(n5329), .Z(n5620) );
  NOR U5517 ( .A(n5619), .B(n5620), .Z(n5623) );
  NOR U5518 ( .A(n79), .B(n122), .Z(n5616) );
  XOR U5519 ( .A(n5332), .B(n5331), .Z(n5615) );
  IV U5520 ( .A(n5615), .Z(n5333) );
  NOR U5521 ( .A(n5616), .B(n5333), .Z(n5618) );
  NOR U5522 ( .A(n117), .B(n122), .Z(n5611) );
  XOR U5523 ( .A(n5335), .B(n5334), .Z(n5610) );
  NOR U5524 ( .A(n5611), .B(n5610), .Z(n5614) );
  XOR U5525 ( .A(n5337), .B(n5336), .Z(n5605) );
  NOR U5526 ( .A(n80), .B(n122), .Z(n5606) );
  IV U5527 ( .A(n5606), .Z(n5338) );
  NOR U5528 ( .A(n5605), .B(n5338), .Z(n5608) );
  XOR U5529 ( .A(n5340), .B(n5339), .Z(n5602) );
  NOR U5530 ( .A(n116), .B(n122), .Z(n5601) );
  IV U5531 ( .A(n5601), .Z(n5341) );
  NOR U5532 ( .A(n5602), .B(n5341), .Z(n5604) );
  XOR U5533 ( .A(n5343), .B(n5342), .Z(n5345) );
  NOR U5534 ( .A(n81), .B(n122), .Z(n5346) );
  IV U5535 ( .A(n5346), .Z(n5344) );
  NOR U5536 ( .A(n5345), .B(n5344), .Z(n5600) );
  XOR U5537 ( .A(n5346), .B(n5345), .Z(n5844) );
  NOR U5538 ( .A(n115), .B(n122), .Z(n5594) );
  XOR U5539 ( .A(n5348), .B(n5347), .Z(n5593) );
  NOR U5540 ( .A(n5594), .B(n5593), .Z(n5597) );
  NOR U5541 ( .A(n82), .B(n122), .Z(n5589) );
  XOR U5542 ( .A(n5350), .B(n5349), .Z(n5588) );
  NOR U5543 ( .A(n5589), .B(n5588), .Z(n5592) );
  NOR U5544 ( .A(n114), .B(n122), .Z(n5584) );
  XOR U5545 ( .A(n5352), .B(n5351), .Z(n5583) );
  NOR U5546 ( .A(n5584), .B(n5583), .Z(n5587) );
  NOR U5547 ( .A(n83), .B(n122), .Z(n5578) );
  XOR U5548 ( .A(n5354), .B(n5353), .Z(n5579) );
  NOR U5549 ( .A(n5578), .B(n5579), .Z(n5582) );
  NOR U5550 ( .A(n113), .B(n122), .Z(n5574) );
  XOR U5551 ( .A(n5356), .B(n5355), .Z(n5573) );
  NOR U5552 ( .A(n5574), .B(n5573), .Z(n5577) );
  NOR U5553 ( .A(n84), .B(n122), .Z(n5569) );
  XOR U5554 ( .A(n5358), .B(n5357), .Z(n5568) );
  NOR U5555 ( .A(n5569), .B(n5568), .Z(n5572) );
  NOR U5556 ( .A(n112), .B(n122), .Z(n5564) );
  XOR U5557 ( .A(n5360), .B(n5359), .Z(n5563) );
  NOR U5558 ( .A(n5564), .B(n5563), .Z(n5567) );
  IV U5559 ( .A(n5361), .Z(n5363) );
  XOR U5560 ( .A(n5363), .B(n5362), .Z(n5558) );
  NOR U5561 ( .A(n85), .B(n122), .Z(n5559) );
  IV U5562 ( .A(n5559), .Z(n5364) );
  NOR U5563 ( .A(n5558), .B(n5364), .Z(n5561) );
  IV U5564 ( .A(n5365), .Z(n5367) );
  XOR U5565 ( .A(n5367), .B(n5366), .Z(n5554) );
  NOR U5566 ( .A(n111), .B(n122), .Z(n5555) );
  IV U5567 ( .A(n5555), .Z(n5368) );
  NOR U5568 ( .A(n5554), .B(n5368), .Z(n5557) );
  IV U5569 ( .A(n5369), .Z(n5371) );
  XOR U5570 ( .A(n5371), .B(n5370), .Z(n5550) );
  NOR U5571 ( .A(n86), .B(n122), .Z(n5551) );
  IV U5572 ( .A(n5551), .Z(n5372) );
  NOR U5573 ( .A(n5550), .B(n5372), .Z(n5553) );
  XOR U5574 ( .A(n5374), .B(n5373), .Z(n5375) );
  IV U5575 ( .A(n5375), .Z(n5546) );
  NOR U5576 ( .A(n110), .B(n122), .Z(n5547) );
  IV U5577 ( .A(n5547), .Z(n5376) );
  NOR U5578 ( .A(n5546), .B(n5376), .Z(n5549) );
  XOR U5579 ( .A(n5378), .B(n5377), .Z(n5379) );
  IV U5580 ( .A(n5379), .Z(n5542) );
  NOR U5581 ( .A(n109), .B(n122), .Z(n5543) );
  IV U5582 ( .A(n5543), .Z(n5380) );
  NOR U5583 ( .A(n5542), .B(n5380), .Z(n5545) );
  XOR U5584 ( .A(n5382), .B(n5381), .Z(n5383) );
  IV U5585 ( .A(n5383), .Z(n5538) );
  NOR U5586 ( .A(n108), .B(n122), .Z(n5539) );
  IV U5587 ( .A(n5539), .Z(n5384) );
  NOR U5588 ( .A(n5538), .B(n5384), .Z(n5541) );
  XOR U5589 ( .A(n5386), .B(n5385), .Z(n5387) );
  IV U5590 ( .A(n5387), .Z(n5534) );
  NOR U5591 ( .A(n87), .B(n122), .Z(n5535) );
  IV U5592 ( .A(n5535), .Z(n5388) );
  NOR U5593 ( .A(n5534), .B(n5388), .Z(n5537) );
  XOR U5594 ( .A(n5390), .B(n5389), .Z(n5391) );
  IV U5595 ( .A(n5391), .Z(n5530) );
  NOR U5596 ( .A(n107), .B(n122), .Z(n5531) );
  IV U5597 ( .A(n5531), .Z(n5392) );
  NOR U5598 ( .A(n5530), .B(n5392), .Z(n5533) );
  XOR U5599 ( .A(n5394), .B(n5393), .Z(n5395) );
  IV U5600 ( .A(n5395), .Z(n5526) );
  NOR U5601 ( .A(n88), .B(n122), .Z(n5527) );
  IV U5602 ( .A(n5527), .Z(n5396) );
  NOR U5603 ( .A(n5526), .B(n5396), .Z(n5529) );
  XOR U5604 ( .A(n5398), .B(n5397), .Z(n5399) );
  IV U5605 ( .A(n5399), .Z(n5522) );
  NOR U5606 ( .A(n106), .B(n122), .Z(n5523) );
  IV U5607 ( .A(n5523), .Z(n5400) );
  NOR U5608 ( .A(n5522), .B(n5400), .Z(n5525) );
  XOR U5609 ( .A(n5402), .B(n5401), .Z(n5403) );
  IV U5610 ( .A(n5403), .Z(n5518) );
  NOR U5611 ( .A(n105), .B(n122), .Z(n5519) );
  IV U5612 ( .A(n5519), .Z(n5404) );
  NOR U5613 ( .A(n5518), .B(n5404), .Z(n5521) );
  XOR U5614 ( .A(n5406), .B(n5405), .Z(n5407) );
  IV U5615 ( .A(n5407), .Z(n5514) );
  NOR U5616 ( .A(n104), .B(n122), .Z(n5515) );
  IV U5617 ( .A(n5515), .Z(n5408) );
  NOR U5618 ( .A(n5514), .B(n5408), .Z(n5517) );
  XOR U5619 ( .A(n5410), .B(n5409), .Z(n5411) );
  IV U5620 ( .A(n5411), .Z(n5510) );
  NOR U5621 ( .A(n89), .B(n122), .Z(n5511) );
  IV U5622 ( .A(n5511), .Z(n5412) );
  NOR U5623 ( .A(n5510), .B(n5412), .Z(n5513) );
  XOR U5624 ( .A(n5414), .B(n5413), .Z(n5415) );
  IV U5625 ( .A(n5415), .Z(n5506) );
  NOR U5626 ( .A(n103), .B(n122), .Z(n5507) );
  IV U5627 ( .A(n5507), .Z(n5416) );
  NOR U5628 ( .A(n5506), .B(n5416), .Z(n5509) );
  XOR U5629 ( .A(n5418), .B(n5417), .Z(n5419) );
  IV U5630 ( .A(n5419), .Z(n5502) );
  NOR U5631 ( .A(n90), .B(n122), .Z(n5503) );
  IV U5632 ( .A(n5503), .Z(n5420) );
  NOR U5633 ( .A(n5502), .B(n5420), .Z(n5505) );
  XOR U5634 ( .A(n5422), .B(n5421), .Z(n5423) );
  IV U5635 ( .A(n5423), .Z(n5498) );
  NOR U5636 ( .A(n102), .B(n122), .Z(n5499) );
  IV U5637 ( .A(n5499), .Z(n5424) );
  NOR U5638 ( .A(n5498), .B(n5424), .Z(n5501) );
  NOR U5639 ( .A(n101), .B(n122), .Z(n5495) );
  IV U5640 ( .A(n5495), .Z(n5428) );
  XOR U5641 ( .A(n5426), .B(n5425), .Z(n5427) );
  IV U5642 ( .A(n5427), .Z(n5494) );
  NOR U5643 ( .A(n5428), .B(n5494), .Z(n5497) );
  NOR U5644 ( .A(n99), .B(n122), .Z(n5482) );
  IV U5645 ( .A(n5482), .Z(n5999) );
  XOR U5646 ( .A(n5430), .B(n5429), .Z(n5481) );
  IV U5647 ( .A(n5481), .Z(n5998) );
  NOR U5648 ( .A(n5999), .B(n5998), .Z(n5485) );
  XOR U5649 ( .A(n5432), .B(n5431), .Z(n5469) );
  IV U5650 ( .A(n5469), .Z(n5941) );
  NOR U5651 ( .A(n91), .B(n122), .Z(n5468) );
  IV U5652 ( .A(n5468), .Z(n5940) );
  NOR U5653 ( .A(n5941), .B(n5940), .Z(n5472) );
  XOR U5654 ( .A(n5434), .B(n5433), .Z(n5435) );
  IV U5655 ( .A(n5435), .Z(n5464) );
  NOR U5656 ( .A(n97), .B(n122), .Z(n5465) );
  IV U5657 ( .A(n5465), .Z(n5436) );
  NOR U5658 ( .A(n5464), .B(n5436), .Z(n5467) );
  NOR U5659 ( .A(n96), .B(n122), .Z(n5461) );
  IV U5660 ( .A(n5461), .Z(n5440) );
  XOR U5661 ( .A(n5438), .B(n5437), .Z(n5439) );
  IV U5662 ( .A(n5439), .Z(n5460) );
  NOR U5663 ( .A(n5440), .B(n5460), .Z(n5463) );
  NOR U5664 ( .A(n93), .B(n122), .Z(n6490) );
  IV U5665 ( .A(n6490), .Z(n5442) );
  NOR U5666 ( .A(n124), .B(n168), .Z(n5445) );
  IV U5667 ( .A(n5445), .Z(n5441) );
  NOR U5668 ( .A(n5442), .B(n5441), .Z(n5960) );
  IV U5669 ( .A(n5960), .Z(n5443) );
  NOR U5670 ( .A(n5444), .B(n5443), .Z(n5452) );
  XOR U5671 ( .A(n5446), .B(n5445), .Z(n5447) );
  NOR U5672 ( .A(n5960), .B(n5447), .Z(n5448) );
  NOR U5673 ( .A(n5452), .B(n5448), .Z(n5449) );
  IV U5674 ( .A(n5449), .Z(n5973) );
  NOR U5675 ( .A(n94), .B(n122), .Z(n5972) );
  IV U5676 ( .A(n5972), .Z(n5450) );
  NOR U5677 ( .A(n5973), .B(n5450), .Z(n5451) );
  NOR U5678 ( .A(n5452), .B(n5451), .Z(n5455) );
  NOR U5679 ( .A(n95), .B(n122), .Z(n5454) );
  IV U5680 ( .A(n5454), .Z(n5453) );
  NOR U5681 ( .A(n5455), .B(n5453), .Z(n5459) );
  XOR U5682 ( .A(n5455), .B(n5454), .Z(n5953) );
  XOR U5683 ( .A(n5457), .B(n5456), .Z(n5954) );
  NOR U5684 ( .A(n5953), .B(n5954), .Z(n5458) );
  NOR U5685 ( .A(n5459), .B(n5458), .Z(n5949) );
  XOR U5686 ( .A(n5461), .B(n5460), .Z(n5950) );
  NOR U5687 ( .A(n5949), .B(n5950), .Z(n5462) );
  NOR U5688 ( .A(n5463), .B(n5462), .Z(n5946) );
  XOR U5689 ( .A(n5465), .B(n5464), .Z(n5945) );
  NOR U5690 ( .A(n5946), .B(n5945), .Z(n5466) );
  NOR U5691 ( .A(n5467), .B(n5466), .Z(n5943) );
  NOR U5692 ( .A(n5469), .B(n5468), .Z(n5470) );
  NOR U5693 ( .A(n5943), .B(n5470), .Z(n5471) );
  NOR U5694 ( .A(n5472), .B(n5471), .Z(n5478) );
  NOR U5695 ( .A(n98), .B(n122), .Z(n5477) );
  IV U5696 ( .A(n5477), .Z(n5473) );
  NOR U5697 ( .A(n5478), .B(n5473), .Z(n5480) );
  IV U5698 ( .A(n5474), .Z(n5476) );
  XOR U5699 ( .A(n5476), .B(n5475), .Z(n5937) );
  XOR U5700 ( .A(n5478), .B(n5477), .Z(n5936) );
  NOR U5701 ( .A(n5937), .B(n5936), .Z(n5479) );
  NOR U5702 ( .A(n5480), .B(n5479), .Z(n6001) );
  NOR U5703 ( .A(n5482), .B(n5481), .Z(n5483) );
  NOR U5704 ( .A(n6001), .B(n5483), .Z(n5484) );
  NOR U5705 ( .A(n5485), .B(n5484), .Z(n5491) );
  NOR U5706 ( .A(n100), .B(n122), .Z(n5490) );
  IV U5707 ( .A(n5490), .Z(n5486) );
  NOR U5708 ( .A(n5491), .B(n5486), .Z(n5493) );
  XOR U5709 ( .A(n5488), .B(n5487), .Z(n5489) );
  IV U5710 ( .A(n5489), .Z(n5933) );
  XOR U5711 ( .A(n5491), .B(n5490), .Z(n5932) );
  NOR U5712 ( .A(n5933), .B(n5932), .Z(n5492) );
  NOR U5713 ( .A(n5493), .B(n5492), .Z(n6012) );
  XOR U5714 ( .A(n5495), .B(n5494), .Z(n6013) );
  NOR U5715 ( .A(n6012), .B(n6013), .Z(n5496) );
  NOR U5716 ( .A(n5497), .B(n5496), .Z(n5929) );
  XOR U5717 ( .A(n5499), .B(n5498), .Z(n5930) );
  NOR U5718 ( .A(n5929), .B(n5930), .Z(n5500) );
  NOR U5719 ( .A(n5501), .B(n5500), .Z(n5924) );
  XOR U5720 ( .A(n5503), .B(n5502), .Z(n5925) );
  NOR U5721 ( .A(n5924), .B(n5925), .Z(n5504) );
  NOR U5722 ( .A(n5505), .B(n5504), .Z(n5920) );
  XOR U5723 ( .A(n5507), .B(n5506), .Z(n5921) );
  NOR U5724 ( .A(n5920), .B(n5921), .Z(n5508) );
  NOR U5725 ( .A(n5509), .B(n5508), .Z(n5917) );
  XOR U5726 ( .A(n5511), .B(n5510), .Z(n5916) );
  NOR U5727 ( .A(n5917), .B(n5916), .Z(n5512) );
  NOR U5728 ( .A(n5513), .B(n5512), .Z(n5913) );
  XOR U5729 ( .A(n5515), .B(n5514), .Z(n5912) );
  NOR U5730 ( .A(n5913), .B(n5912), .Z(n5516) );
  NOR U5731 ( .A(n5517), .B(n5516), .Z(n5908) );
  XOR U5732 ( .A(n5519), .B(n5518), .Z(n5909) );
  NOR U5733 ( .A(n5908), .B(n5909), .Z(n5520) );
  NOR U5734 ( .A(n5521), .B(n5520), .Z(n5904) );
  XOR U5735 ( .A(n5523), .B(n5522), .Z(n5905) );
  NOR U5736 ( .A(n5904), .B(n5905), .Z(n5524) );
  NOR U5737 ( .A(n5525), .B(n5524), .Z(n5900) );
  XOR U5738 ( .A(n5527), .B(n5526), .Z(n5901) );
  NOR U5739 ( .A(n5900), .B(n5901), .Z(n5528) );
  NOR U5740 ( .A(n5529), .B(n5528), .Z(n5896) );
  XOR U5741 ( .A(n5531), .B(n5530), .Z(n5897) );
  NOR U5742 ( .A(n5896), .B(n5897), .Z(n5532) );
  NOR U5743 ( .A(n5533), .B(n5532), .Z(n5892) );
  XOR U5744 ( .A(n5535), .B(n5534), .Z(n5893) );
  NOR U5745 ( .A(n5892), .B(n5893), .Z(n5536) );
  NOR U5746 ( .A(n5537), .B(n5536), .Z(n5888) );
  XOR U5747 ( .A(n5539), .B(n5538), .Z(n5889) );
  NOR U5748 ( .A(n5888), .B(n5889), .Z(n5540) );
  NOR U5749 ( .A(n5541), .B(n5540), .Z(n5884) );
  XOR U5750 ( .A(n5543), .B(n5542), .Z(n5885) );
  NOR U5751 ( .A(n5884), .B(n5885), .Z(n5544) );
  NOR U5752 ( .A(n5545), .B(n5544), .Z(n5880) );
  XOR U5753 ( .A(n5547), .B(n5546), .Z(n5881) );
  NOR U5754 ( .A(n5880), .B(n5881), .Z(n5548) );
  NOR U5755 ( .A(n5549), .B(n5548), .Z(n5876) );
  XOR U5756 ( .A(n5551), .B(n5550), .Z(n5877) );
  NOR U5757 ( .A(n5876), .B(n5877), .Z(n5552) );
  NOR U5758 ( .A(n5553), .B(n5552), .Z(n5872) );
  XOR U5759 ( .A(n5555), .B(n5554), .Z(n5873) );
  NOR U5760 ( .A(n5872), .B(n5873), .Z(n5556) );
  NOR U5761 ( .A(n5557), .B(n5556), .Z(n5868) );
  XOR U5762 ( .A(n5559), .B(n5558), .Z(n5869) );
  NOR U5763 ( .A(n5868), .B(n5869), .Z(n5560) );
  NOR U5764 ( .A(n5561), .B(n5560), .Z(n5562) );
  IV U5765 ( .A(n5562), .Z(n5866) );
  XOR U5766 ( .A(n5564), .B(n5563), .Z(n5565) );
  IV U5767 ( .A(n5565), .Z(n5865) );
  NOR U5768 ( .A(n5866), .B(n5865), .Z(n5566) );
  NOR U5769 ( .A(n5567), .B(n5566), .Z(n5863) );
  XOR U5770 ( .A(n5569), .B(n5568), .Z(n5570) );
  IV U5771 ( .A(n5570), .Z(n5862) );
  NOR U5772 ( .A(n5863), .B(n5862), .Z(n5571) );
  NOR U5773 ( .A(n5572), .B(n5571), .Z(n5860) );
  XOR U5774 ( .A(n5574), .B(n5573), .Z(n5575) );
  IV U5775 ( .A(n5575), .Z(n5859) );
  NOR U5776 ( .A(n5860), .B(n5859), .Z(n5576) );
  NOR U5777 ( .A(n5577), .B(n5576), .Z(n5857) );
  IV U5778 ( .A(n5578), .Z(n5580) );
  XOR U5779 ( .A(n5580), .B(n5579), .Z(n5856) );
  NOR U5780 ( .A(n5857), .B(n5856), .Z(n5581) );
  NOR U5781 ( .A(n5582), .B(n5581), .Z(n5854) );
  XOR U5782 ( .A(n5584), .B(n5583), .Z(n5585) );
  IV U5783 ( .A(n5585), .Z(n5853) );
  NOR U5784 ( .A(n5854), .B(n5853), .Z(n5586) );
  NOR U5785 ( .A(n5587), .B(n5586), .Z(n5851) );
  XOR U5786 ( .A(n5589), .B(n5588), .Z(n5590) );
  IV U5787 ( .A(n5590), .Z(n5850) );
  NOR U5788 ( .A(n5851), .B(n5850), .Z(n5591) );
  NOR U5789 ( .A(n5592), .B(n5591), .Z(n5848) );
  XOR U5790 ( .A(n5594), .B(n5593), .Z(n5595) );
  IV U5791 ( .A(n5595), .Z(n5847) );
  NOR U5792 ( .A(n5848), .B(n5847), .Z(n5596) );
  NOR U5793 ( .A(n5597), .B(n5596), .Z(n5845) );
  IV U5794 ( .A(n5845), .Z(n5598) );
  NOR U5795 ( .A(n5844), .B(n5598), .Z(n5599) );
  NOR U5796 ( .A(n5600), .B(n5599), .Z(n5840) );
  XOR U5797 ( .A(n5602), .B(n5601), .Z(n5841) );
  NOR U5798 ( .A(n5840), .B(n5841), .Z(n5603) );
  NOR U5799 ( .A(n5604), .B(n5603), .Z(n5836) );
  XOR U5800 ( .A(n5606), .B(n5605), .Z(n5837) );
  NOR U5801 ( .A(n5836), .B(n5837), .Z(n5607) );
  NOR U5802 ( .A(n5608), .B(n5607), .Z(n5609) );
  IV U5803 ( .A(n5609), .Z(n5834) );
  XOR U5804 ( .A(n5611), .B(n5610), .Z(n5612) );
  IV U5805 ( .A(n5612), .Z(n5833) );
  NOR U5806 ( .A(n5834), .B(n5833), .Z(n5613) );
  NOR U5807 ( .A(n5614), .B(n5613), .Z(n5831) );
  XOR U5808 ( .A(n5616), .B(n5615), .Z(n5830) );
  NOR U5809 ( .A(n5831), .B(n5830), .Z(n5617) );
  NOR U5810 ( .A(n5618), .B(n5617), .Z(n5828) );
  IV U5811 ( .A(n5619), .Z(n5621) );
  XOR U5812 ( .A(n5621), .B(n5620), .Z(n5827) );
  NOR U5813 ( .A(n5828), .B(n5827), .Z(n5622) );
  NOR U5814 ( .A(n5623), .B(n5622), .Z(n5825) );
  XOR U5815 ( .A(n5625), .B(n5624), .Z(n5626) );
  IV U5816 ( .A(n5626), .Z(n5824) );
  NOR U5817 ( .A(n5825), .B(n5824), .Z(n5627) );
  NOR U5818 ( .A(n5628), .B(n5627), .Z(n5822) );
  XOR U5819 ( .A(n5630), .B(n5629), .Z(n5631) );
  IV U5820 ( .A(n5631), .Z(n5821) );
  NOR U5821 ( .A(n5822), .B(n5821), .Z(n5632) );
  NOR U5822 ( .A(n5633), .B(n5632), .Z(n5819) );
  IV U5823 ( .A(n5634), .Z(n5636) );
  XOR U5824 ( .A(n5636), .B(n5635), .Z(n5818) );
  NOR U5825 ( .A(n5819), .B(n5818), .Z(n5637) );
  NOR U5826 ( .A(n5638), .B(n5637), .Z(n5816) );
  XOR U5827 ( .A(n5640), .B(n5639), .Z(n5641) );
  IV U5828 ( .A(n5641), .Z(n5815) );
  NOR U5829 ( .A(n5816), .B(n5815), .Z(n5642) );
  NOR U5830 ( .A(n5643), .B(n5642), .Z(n5813) );
  IV U5831 ( .A(n5644), .Z(n5646) );
  XOR U5832 ( .A(n5646), .B(n5645), .Z(n5812) );
  NOR U5833 ( .A(n5813), .B(n5812), .Z(n5647) );
  NOR U5834 ( .A(n5648), .B(n5647), .Z(n5810) );
  IV U5835 ( .A(n5649), .Z(n5651) );
  XOR U5836 ( .A(n5651), .B(n5650), .Z(n5809) );
  NOR U5837 ( .A(n5810), .B(n5809), .Z(n5652) );
  NOR U5838 ( .A(n5653), .B(n5652), .Z(n6167) );
  NOR U5839 ( .A(n133), .B(n122), .Z(n6164) );
  NOR U5840 ( .A(n131), .B(n124), .Z(n5654) );
  IV U5841 ( .A(n5654), .Z(n6176) );
  NOR U5842 ( .A(n5656), .B(n5655), .Z(n5660) );
  NOR U5843 ( .A(n5658), .B(n5657), .Z(n5659) );
  NOR U5844 ( .A(n5660), .B(n5659), .Z(n6173) );
  IV U5845 ( .A(n5661), .Z(n5662) );
  NOR U5846 ( .A(n5663), .B(n5662), .Z(n5667) );
  NOR U5847 ( .A(n5665), .B(n5664), .Z(n5666) );
  NOR U5848 ( .A(n5667), .B(n5666), .Z(n6183) );
  NOR U5849 ( .A(n128), .B(n127), .Z(n6181) );
  IV U5850 ( .A(n6181), .Z(n5807) );
  IV U5851 ( .A(n5668), .Z(n5669) );
  NOR U5852 ( .A(n5670), .B(n5669), .Z(n5674) );
  NOR U5853 ( .A(n5672), .B(n5671), .Z(n5673) );
  NOR U5854 ( .A(n5674), .B(n5673), .Z(n5675) );
  IV U5855 ( .A(n5675), .Z(n6320) );
  NOR U5856 ( .A(n5677), .B(n5676), .Z(n5682) );
  IV U5857 ( .A(n5678), .Z(n5679) );
  NOR U5858 ( .A(n5680), .B(n5679), .Z(n5681) );
  NOR U5859 ( .A(n5682), .B(n5681), .Z(n6190) );
  NOR U5860 ( .A(n125), .B(n130), .Z(n6188) );
  NOR U5861 ( .A(n123), .B(n132), .Z(n6197) );
  NOR U5862 ( .A(n5684), .B(n5683), .Z(n5690) );
  IV U5863 ( .A(n5685), .Z(n5688) );
  IV U5864 ( .A(n5686), .Z(n5687) );
  NOR U5865 ( .A(n5688), .B(n5687), .Z(n5689) );
  NOR U5866 ( .A(n5690), .B(n5689), .Z(n6193) );
  NOR U5867 ( .A(n5692), .B(n5691), .Z(n5696) );
  NOR U5868 ( .A(n5694), .B(n5693), .Z(n5695) );
  NOR U5869 ( .A(n5696), .B(n5695), .Z(n6205) );
  NOR U5870 ( .A(n120), .B(n134), .Z(n6202) );
  IV U5871 ( .A(n5697), .Z(n5698) );
  NOR U5872 ( .A(n5699), .B(n5698), .Z(n5703) );
  NOR U5873 ( .A(n5701), .B(n5700), .Z(n5702) );
  NOR U5874 ( .A(n5703), .B(n5702), .Z(n6306) );
  NOR U5875 ( .A(n5705), .B(n5704), .Z(n5709) );
  NOR U5876 ( .A(n5707), .B(n5706), .Z(n5708) );
  NOR U5877 ( .A(n5709), .B(n5708), .Z(n6211) );
  NOR U5878 ( .A(n79), .B(n138), .Z(n6209) );
  IV U5879 ( .A(n6209), .Z(n5806) );
  IV U5880 ( .A(n5710), .Z(n5711) );
  NOR U5881 ( .A(n5712), .B(n5711), .Z(n5716) );
  NOR U5882 ( .A(n5714), .B(n5713), .Z(n5715) );
  NOR U5883 ( .A(n5716), .B(n5715), .Z(n6216) );
  NOR U5884 ( .A(n117), .B(n140), .Z(n6215) );
  NOR U5885 ( .A(n5718), .B(n5717), .Z(n5722) );
  NOR U5886 ( .A(n5720), .B(n5719), .Z(n5721) );
  NOR U5887 ( .A(n5722), .B(n5721), .Z(n6226) );
  NOR U5888 ( .A(n80), .B(n142), .Z(n6223) );
  IV U5889 ( .A(n5723), .Z(n5724) );
  NOR U5890 ( .A(n5725), .B(n5724), .Z(n5729) );
  NOR U5891 ( .A(n5727), .B(n5726), .Z(n5728) );
  NOR U5892 ( .A(n5729), .B(n5728), .Z(n6239) );
  NOR U5893 ( .A(n81), .B(n146), .Z(n6237) );
  IV U5894 ( .A(n6237), .Z(n5797) );
  NOR U5895 ( .A(n5731), .B(n5730), .Z(n5736) );
  IV U5896 ( .A(n5732), .Z(n5733) );
  NOR U5897 ( .A(n5734), .B(n5733), .Z(n5735) );
  NOR U5898 ( .A(n5736), .B(n5735), .Z(n6252) );
  NOR U5899 ( .A(n82), .B(n151), .Z(n6250) );
  NOR U5900 ( .A(n5738), .B(n5737), .Z(n5744) );
  IV U5901 ( .A(n5739), .Z(n5742) );
  IV U5902 ( .A(n5740), .Z(n5741) );
  NOR U5903 ( .A(n5742), .B(n5741), .Z(n5743) );
  NOR U5904 ( .A(n5744), .B(n5743), .Z(n6259) );
  NOR U5905 ( .A(n5746), .B(n5745), .Z(n5750) );
  NOR U5906 ( .A(n5748), .B(n5747), .Z(n5749) );
  NOR U5907 ( .A(n5750), .B(n5749), .Z(n6265) );
  NOR U5908 ( .A(n83), .B(n154), .Z(n6263) );
  IV U5909 ( .A(n6263), .Z(n5787) );
  NOR U5910 ( .A(n5752), .B(n5751), .Z(n5756) );
  NOR U5911 ( .A(n5754), .B(n5753), .Z(n5755) );
  NOR U5912 ( .A(n5756), .B(n5755), .Z(n6297) );
  IV U5913 ( .A(n6297), .Z(n5785) );
  NOR U5914 ( .A(n5758), .B(n5757), .Z(n5762) );
  NOR U5915 ( .A(n5760), .B(n5759), .Z(n5761) );
  NOR U5916 ( .A(n5762), .B(n5761), .Z(n6271) );
  NOR U5917 ( .A(n84), .B(n159), .Z(n6269) );
  IV U5918 ( .A(n6269), .Z(n5784) );
  NOR U5919 ( .A(n5764), .B(n5763), .Z(n5768) );
  NOR U5920 ( .A(n5766), .B(n5765), .Z(n5767) );
  NOR U5921 ( .A(n5768), .B(n5767), .Z(n6277) );
  NOR U5922 ( .A(n85), .B(n162), .Z(n6275) );
  IV U5923 ( .A(n6275), .Z(n5777) );
  IV U5924 ( .A(n5769), .Z(n5770) );
  NOR U5925 ( .A(n5771), .B(n5770), .Z(n5775) );
  NOR U5926 ( .A(n5773), .B(n5772), .Z(n5774) );
  NOR U5927 ( .A(n5775), .B(n5774), .Z(n6282) );
  NOR U5928 ( .A(n164), .B(n111), .Z(n6280) );
  XOR U5929 ( .A(n6282), .B(n6280), .Z(n6284) );
  NOR U5930 ( .A(n166), .B(n86), .Z(n5776) );
  IV U5931 ( .A(n5776), .Z(n6283) );
  XOR U5932 ( .A(n6284), .B(n6283), .Z(n6274) );
  XOR U5933 ( .A(n5777), .B(n6274), .Z(n6276) );
  XOR U5934 ( .A(n6277), .B(n6276), .Z(n6293) );
  NOR U5935 ( .A(n5779), .B(n5778), .Z(n5783) );
  NOR U5936 ( .A(n5781), .B(n5780), .Z(n5782) );
  NOR U5937 ( .A(n5783), .B(n5782), .Z(n6291) );
  NOR U5938 ( .A(n112), .B(n160), .Z(n6289) );
  XOR U5939 ( .A(n6291), .B(n6289), .Z(n6292) );
  XOR U5940 ( .A(n6293), .B(n6292), .Z(n6268) );
  XOR U5941 ( .A(n5784), .B(n6268), .Z(n6270) );
  XOR U5942 ( .A(n6271), .B(n6270), .Z(n6298) );
  XOR U5943 ( .A(n5785), .B(n6298), .Z(n6300) );
  NOR U5944 ( .A(n113), .B(n157), .Z(n5786) );
  IV U5945 ( .A(n5786), .Z(n6299) );
  XOR U5946 ( .A(n6300), .B(n6299), .Z(n6262) );
  XOR U5947 ( .A(n5787), .B(n6262), .Z(n6264) );
  XOR U5948 ( .A(n6265), .B(n6264), .Z(n6257) );
  NOR U5949 ( .A(n114), .B(n152), .Z(n6255) );
  XOR U5950 ( .A(n6257), .B(n6255), .Z(n6258) );
  XOR U5951 ( .A(n6259), .B(n6258), .Z(n6249) );
  XOR U5952 ( .A(n6250), .B(n6249), .Z(n5788) );
  IV U5953 ( .A(n5788), .Z(n6251) );
  XOR U5954 ( .A(n6252), .B(n6251), .Z(n6244) );
  NOR U5955 ( .A(n115), .B(n149), .Z(n6242) );
  XOR U5956 ( .A(n6244), .B(n6242), .Z(n6246) );
  IV U5957 ( .A(n5789), .Z(n5791) );
  NOR U5958 ( .A(n5791), .B(n5790), .Z(n5795) );
  NOR U5959 ( .A(n5793), .B(n5792), .Z(n5794) );
  NOR U5960 ( .A(n5795), .B(n5794), .Z(n5796) );
  IV U5961 ( .A(n5796), .Z(n6245) );
  XOR U5962 ( .A(n6246), .B(n6245), .Z(n6236) );
  XOR U5963 ( .A(n5797), .B(n6236), .Z(n6238) );
  XOR U5964 ( .A(n6239), .B(n6238), .Z(n6233) );
  IV U5965 ( .A(n5798), .Z(n5799) );
  NOR U5966 ( .A(n5800), .B(n5799), .Z(n5804) );
  NOR U5967 ( .A(n5802), .B(n5801), .Z(n5803) );
  NOR U5968 ( .A(n5804), .B(n5803), .Z(n6231) );
  NOR U5969 ( .A(n116), .B(n144), .Z(n6229) );
  XOR U5970 ( .A(n6231), .B(n6229), .Z(n6232) );
  XOR U5971 ( .A(n6233), .B(n6232), .Z(n6222) );
  XOR U5972 ( .A(n6223), .B(n6222), .Z(n6224) );
  XOR U5973 ( .A(n6226), .B(n6224), .Z(n6214) );
  XOR U5974 ( .A(n6215), .B(n6214), .Z(n5805) );
  IV U5975 ( .A(n5805), .Z(n6217) );
  XOR U5976 ( .A(n6216), .B(n6217), .Z(n6208) );
  XOR U5977 ( .A(n5806), .B(n6208), .Z(n6210) );
  XOR U5978 ( .A(n6211), .B(n6210), .Z(n6307) );
  XOR U5979 ( .A(n6306), .B(n6307), .Z(n6308) );
  NOR U5980 ( .A(n119), .B(n136), .Z(n6309) );
  XOR U5981 ( .A(n6308), .B(n6309), .Z(n6201) );
  XOR U5982 ( .A(n6202), .B(n6201), .Z(n6203) );
  XOR U5983 ( .A(n6205), .B(n6203), .Z(n6194) );
  XOR U5984 ( .A(n6193), .B(n6194), .Z(n6196) );
  XOR U5985 ( .A(n6197), .B(n6196), .Z(n6186) );
  XOR U5986 ( .A(n6188), .B(n6186), .Z(n6189) );
  XOR U5987 ( .A(n6190), .B(n6189), .Z(n6318) );
  NOR U5988 ( .A(n126), .B(n129), .Z(n6316) );
  XOR U5989 ( .A(n6318), .B(n6316), .Z(n6319) );
  XOR U5990 ( .A(n6320), .B(n6319), .Z(n6180) );
  XOR U5991 ( .A(n5807), .B(n6180), .Z(n6182) );
  XOR U5992 ( .A(n6183), .B(n6182), .Z(n6174) );
  XOR U5993 ( .A(n6173), .B(n6174), .Z(n6175) );
  XOR U5994 ( .A(n6176), .B(n6175), .Z(n6166) );
  XOR U5995 ( .A(n6164), .B(n6166), .Z(n6169) );
  XOR U5996 ( .A(n6167), .B(n6169), .Z(n6160) );
  NOR U5997 ( .A(n135), .B(n121), .Z(n6161) );
  IV U5998 ( .A(n6161), .Z(n5808) );
  NOR U5999 ( .A(n6160), .B(n5808), .Z(n6163) );
  XOR U6000 ( .A(n5810), .B(n5809), .Z(n6157) );
  NOR U6001 ( .A(n133), .B(n121), .Z(n6156) );
  IV U6002 ( .A(n6156), .Z(n5811) );
  NOR U6003 ( .A(n6157), .B(n5811), .Z(n6159) );
  XOR U6004 ( .A(n5813), .B(n5812), .Z(n6153) );
  NOR U6005 ( .A(n131), .B(n121), .Z(n6152) );
  IV U6006 ( .A(n6152), .Z(n5814) );
  NOR U6007 ( .A(n6153), .B(n5814), .Z(n6155) );
  XOR U6008 ( .A(n5816), .B(n5815), .Z(n6149) );
  NOR U6009 ( .A(n128), .B(n121), .Z(n6148) );
  IV U6010 ( .A(n6148), .Z(n5817) );
  NOR U6011 ( .A(n6149), .B(n5817), .Z(n6151) );
  XOR U6012 ( .A(n5819), .B(n5818), .Z(n6145) );
  NOR U6013 ( .A(n126), .B(n121), .Z(n6144) );
  IV U6014 ( .A(n6144), .Z(n5820) );
  NOR U6015 ( .A(n6145), .B(n5820), .Z(n6147) );
  XOR U6016 ( .A(n5822), .B(n5821), .Z(n6141) );
  NOR U6017 ( .A(n125), .B(n121), .Z(n6140) );
  IV U6018 ( .A(n6140), .Z(n5823) );
  NOR U6019 ( .A(n6141), .B(n5823), .Z(n6143) );
  XOR U6020 ( .A(n5825), .B(n5824), .Z(n6137) );
  NOR U6021 ( .A(n123), .B(n121), .Z(n6136) );
  IV U6022 ( .A(n6136), .Z(n5826) );
  NOR U6023 ( .A(n6137), .B(n5826), .Z(n6139) );
  XOR U6024 ( .A(n5828), .B(n5827), .Z(n6133) );
  NOR U6025 ( .A(n120), .B(n121), .Z(n6132) );
  IV U6026 ( .A(n6132), .Z(n5829) );
  NOR U6027 ( .A(n6133), .B(n5829), .Z(n6135) );
  XOR U6028 ( .A(n5831), .B(n5830), .Z(n6129) );
  NOR U6029 ( .A(n119), .B(n121), .Z(n6128) );
  IV U6030 ( .A(n6128), .Z(n5832) );
  NOR U6031 ( .A(n6129), .B(n5832), .Z(n6131) );
  XOR U6032 ( .A(n5834), .B(n5833), .Z(n6125) );
  NOR U6033 ( .A(n79), .B(n121), .Z(n6124) );
  IV U6034 ( .A(n6124), .Z(n5835) );
  NOR U6035 ( .A(n6125), .B(n5835), .Z(n6127) );
  IV U6036 ( .A(n5836), .Z(n5838) );
  XOR U6037 ( .A(n5838), .B(n5837), .Z(n6120) );
  NOR U6038 ( .A(n117), .B(n121), .Z(n6121) );
  IV U6039 ( .A(n6121), .Z(n5839) );
  NOR U6040 ( .A(n6120), .B(n5839), .Z(n6123) );
  IV U6041 ( .A(n5840), .Z(n5842) );
  XOR U6042 ( .A(n5842), .B(n5841), .Z(n6116) );
  NOR U6043 ( .A(n80), .B(n121), .Z(n6117) );
  IV U6044 ( .A(n6117), .Z(n5843) );
  NOR U6045 ( .A(n6116), .B(n5843), .Z(n6119) );
  XOR U6046 ( .A(n5845), .B(n5844), .Z(n6112) );
  NOR U6047 ( .A(n116), .B(n121), .Z(n6113) );
  IV U6048 ( .A(n6113), .Z(n5846) );
  NOR U6049 ( .A(n6112), .B(n5846), .Z(n6115) );
  XOR U6050 ( .A(n5848), .B(n5847), .Z(n6109) );
  NOR U6051 ( .A(n81), .B(n121), .Z(n6108) );
  IV U6052 ( .A(n6108), .Z(n5849) );
  NOR U6053 ( .A(n6109), .B(n5849), .Z(n6111) );
  XOR U6054 ( .A(n5851), .B(n5850), .Z(n6105) );
  NOR U6055 ( .A(n115), .B(n121), .Z(n6104) );
  IV U6056 ( .A(n6104), .Z(n5852) );
  NOR U6057 ( .A(n6105), .B(n5852), .Z(n6107) );
  XOR U6058 ( .A(n5854), .B(n5853), .Z(n6101) );
  NOR U6059 ( .A(n82), .B(n121), .Z(n6100) );
  IV U6060 ( .A(n6100), .Z(n5855) );
  NOR U6061 ( .A(n6101), .B(n5855), .Z(n6103) );
  XOR U6062 ( .A(n5857), .B(n5856), .Z(n6097) );
  NOR U6063 ( .A(n114), .B(n121), .Z(n6096) );
  IV U6064 ( .A(n6096), .Z(n5858) );
  NOR U6065 ( .A(n6097), .B(n5858), .Z(n6099) );
  XOR U6066 ( .A(n5860), .B(n5859), .Z(n6093) );
  NOR U6067 ( .A(n83), .B(n121), .Z(n6092) );
  IV U6068 ( .A(n6092), .Z(n5861) );
  NOR U6069 ( .A(n6093), .B(n5861), .Z(n6095) );
  XOR U6070 ( .A(n5863), .B(n5862), .Z(n6089) );
  NOR U6071 ( .A(n113), .B(n121), .Z(n6088) );
  IV U6072 ( .A(n6088), .Z(n5864) );
  NOR U6073 ( .A(n6089), .B(n5864), .Z(n6091) );
  XOR U6074 ( .A(n5866), .B(n5865), .Z(n6085) );
  NOR U6075 ( .A(n84), .B(n121), .Z(n6084) );
  IV U6076 ( .A(n6084), .Z(n5867) );
  NOR U6077 ( .A(n6085), .B(n5867), .Z(n6087) );
  IV U6078 ( .A(n5868), .Z(n5870) );
  XOR U6079 ( .A(n5870), .B(n5869), .Z(n6080) );
  NOR U6080 ( .A(n112), .B(n121), .Z(n6081) );
  IV U6081 ( .A(n6081), .Z(n5871) );
  NOR U6082 ( .A(n6080), .B(n5871), .Z(n6083) );
  IV U6083 ( .A(n5872), .Z(n5874) );
  XOR U6084 ( .A(n5874), .B(n5873), .Z(n6076) );
  NOR U6085 ( .A(n85), .B(n121), .Z(n6077) );
  IV U6086 ( .A(n6077), .Z(n5875) );
  NOR U6087 ( .A(n6076), .B(n5875), .Z(n6079) );
  IV U6088 ( .A(n5876), .Z(n5878) );
  XOR U6089 ( .A(n5878), .B(n5877), .Z(n6072) );
  NOR U6090 ( .A(n111), .B(n121), .Z(n6073) );
  IV U6091 ( .A(n6073), .Z(n5879) );
  NOR U6092 ( .A(n6072), .B(n5879), .Z(n6075) );
  XOR U6093 ( .A(n5881), .B(n5880), .Z(n5882) );
  IV U6094 ( .A(n5882), .Z(n6068) );
  NOR U6095 ( .A(n86), .B(n121), .Z(n6069) );
  IV U6096 ( .A(n6069), .Z(n5883) );
  NOR U6097 ( .A(n6068), .B(n5883), .Z(n6071) );
  XOR U6098 ( .A(n5885), .B(n5884), .Z(n5886) );
  IV U6099 ( .A(n5886), .Z(n6064) );
  NOR U6100 ( .A(n110), .B(n121), .Z(n6065) );
  IV U6101 ( .A(n6065), .Z(n5887) );
  NOR U6102 ( .A(n6064), .B(n5887), .Z(n6067) );
  XOR U6103 ( .A(n5889), .B(n5888), .Z(n5890) );
  IV U6104 ( .A(n5890), .Z(n6060) );
  NOR U6105 ( .A(n109), .B(n121), .Z(n6061) );
  IV U6106 ( .A(n6061), .Z(n5891) );
  NOR U6107 ( .A(n6060), .B(n5891), .Z(n6063) );
  IV U6108 ( .A(n5892), .Z(n5894) );
  XOR U6109 ( .A(n5894), .B(n5893), .Z(n6056) );
  NOR U6110 ( .A(n108), .B(n121), .Z(n6057) );
  IV U6111 ( .A(n6057), .Z(n5895) );
  NOR U6112 ( .A(n6056), .B(n5895), .Z(n6059) );
  XOR U6113 ( .A(n5897), .B(n5896), .Z(n5898) );
  IV U6114 ( .A(n5898), .Z(n6052) );
  NOR U6115 ( .A(n87), .B(n121), .Z(n6053) );
  IV U6116 ( .A(n6053), .Z(n5899) );
  NOR U6117 ( .A(n6052), .B(n5899), .Z(n6055) );
  XOR U6118 ( .A(n5901), .B(n5900), .Z(n5902) );
  IV U6119 ( .A(n5902), .Z(n6048) );
  NOR U6120 ( .A(n107), .B(n121), .Z(n6049) );
  IV U6121 ( .A(n6049), .Z(n5903) );
  NOR U6122 ( .A(n6048), .B(n5903), .Z(n6051) );
  XOR U6123 ( .A(n5905), .B(n5904), .Z(n5906) );
  IV U6124 ( .A(n5906), .Z(n6044) );
  NOR U6125 ( .A(n88), .B(n121), .Z(n6045) );
  IV U6126 ( .A(n6045), .Z(n5907) );
  NOR U6127 ( .A(n6044), .B(n5907), .Z(n6047) );
  XOR U6128 ( .A(n5909), .B(n5908), .Z(n5910) );
  IV U6129 ( .A(n5910), .Z(n6040) );
  NOR U6130 ( .A(n106), .B(n121), .Z(n6041) );
  IV U6131 ( .A(n6041), .Z(n5911) );
  NOR U6132 ( .A(n6040), .B(n5911), .Z(n6043) );
  IV U6133 ( .A(n5912), .Z(n5914) );
  XOR U6134 ( .A(n5914), .B(n5913), .Z(n6036) );
  NOR U6135 ( .A(n105), .B(n121), .Z(n6037) );
  IV U6136 ( .A(n6037), .Z(n5915) );
  NOR U6137 ( .A(n6036), .B(n5915), .Z(n6039) );
  IV U6138 ( .A(n5916), .Z(n5918) );
  XOR U6139 ( .A(n5918), .B(n5917), .Z(n6032) );
  NOR U6140 ( .A(n104), .B(n121), .Z(n6033) );
  IV U6141 ( .A(n6033), .Z(n5919) );
  NOR U6142 ( .A(n6032), .B(n5919), .Z(n6035) );
  XOR U6143 ( .A(n5921), .B(n5920), .Z(n5922) );
  IV U6144 ( .A(n5922), .Z(n6028) );
  NOR U6145 ( .A(n89), .B(n121), .Z(n6029) );
  IV U6146 ( .A(n6029), .Z(n5923) );
  NOR U6147 ( .A(n6028), .B(n5923), .Z(n6031) );
  XOR U6148 ( .A(n5925), .B(n5924), .Z(n5926) );
  IV U6149 ( .A(n5926), .Z(n6024) );
  NOR U6150 ( .A(n103), .B(n121), .Z(n6025) );
  IV U6151 ( .A(n6025), .Z(n5927) );
  NOR U6152 ( .A(n6024), .B(n5927), .Z(n6027) );
  NOR U6153 ( .A(n90), .B(n121), .Z(n5928) );
  IV U6154 ( .A(n5928), .Z(n6020) );
  XOR U6155 ( .A(n5930), .B(n5929), .Z(n5931) );
  IV U6156 ( .A(n5931), .Z(n6019) );
  NOR U6157 ( .A(n6020), .B(n6019), .Z(n6023) );
  XOR U6158 ( .A(n5933), .B(n5932), .Z(n5934) );
  NOR U6159 ( .A(n101), .B(n121), .Z(n5935) );
  NOR U6160 ( .A(n5934), .B(n5935), .Z(n6009) );
  IV U6161 ( .A(n5934), .Z(n6541) );
  IV U6162 ( .A(n5935), .Z(n6540) );
  NOR U6163 ( .A(n6541), .B(n6540), .Z(n6007) );
  XOR U6164 ( .A(n5937), .B(n5936), .Z(n5938) );
  NOR U6165 ( .A(n99), .B(n121), .Z(n5939) );
  NOR U6166 ( .A(n5938), .B(n5939), .Z(n5995) );
  IV U6167 ( .A(n5938), .Z(n6465) );
  IV U6168 ( .A(n5939), .Z(n6464) );
  NOR U6169 ( .A(n6465), .B(n6464), .Z(n5993) );
  XOR U6170 ( .A(n5941), .B(n5940), .Z(n5942) );
  XOR U6171 ( .A(n5943), .B(n5942), .Z(n5989) );
  NOR U6172 ( .A(n98), .B(n121), .Z(n5988) );
  IV U6173 ( .A(n5988), .Z(n5944) );
  NOR U6174 ( .A(n5989), .B(n5944), .Z(n5991) );
  XOR U6175 ( .A(n5946), .B(n5945), .Z(n5984) );
  IV U6176 ( .A(n5984), .Z(n5948) );
  NOR U6177 ( .A(n91), .B(n121), .Z(n5947) );
  IV U6178 ( .A(n5947), .Z(n5985) );
  NOR U6179 ( .A(n5948), .B(n5985), .Z(n5987) );
  IV U6180 ( .A(n5949), .Z(n5951) );
  XOR U6181 ( .A(n5951), .B(n5950), .Z(n5980) );
  NOR U6182 ( .A(n97), .B(n121), .Z(n5981) );
  IV U6183 ( .A(n5981), .Z(n5952) );
  NOR U6184 ( .A(n5980), .B(n5952), .Z(n5983) );
  NOR U6185 ( .A(n96), .B(n121), .Z(n5977) );
  IV U6186 ( .A(n5977), .Z(n5956) );
  XOR U6187 ( .A(n5954), .B(n5953), .Z(n5955) );
  IV U6188 ( .A(n5955), .Z(n5976) );
  NOR U6189 ( .A(n5956), .B(n5976), .Z(n5979) );
  NOR U6190 ( .A(n93), .B(n121), .Z(n7045) );
  IV U6191 ( .A(n7045), .Z(n5958) );
  NOR U6192 ( .A(n122), .B(n168), .Z(n5961) );
  IV U6193 ( .A(n5961), .Z(n5957) );
  NOR U6194 ( .A(n5958), .B(n5957), .Z(n6488) );
  IV U6195 ( .A(n6488), .Z(n5959) );
  NOR U6196 ( .A(n5960), .B(n5959), .Z(n5968) );
  XOR U6197 ( .A(n5962), .B(n5961), .Z(n5963) );
  NOR U6198 ( .A(n6488), .B(n5963), .Z(n5964) );
  NOR U6199 ( .A(n5968), .B(n5964), .Z(n5965) );
  IV U6200 ( .A(n5965), .Z(n6502) );
  NOR U6201 ( .A(n94), .B(n121), .Z(n6501) );
  IV U6202 ( .A(n6501), .Z(n5966) );
  NOR U6203 ( .A(n6502), .B(n5966), .Z(n5967) );
  NOR U6204 ( .A(n5968), .B(n5967), .Z(n5971) );
  NOR U6205 ( .A(n95), .B(n121), .Z(n5970) );
  IV U6206 ( .A(n5970), .Z(n5969) );
  NOR U6207 ( .A(n5971), .B(n5969), .Z(n5975) );
  XOR U6208 ( .A(n5971), .B(n5970), .Z(n6481) );
  XOR U6209 ( .A(n5973), .B(n5972), .Z(n6482) );
  NOR U6210 ( .A(n6481), .B(n6482), .Z(n5974) );
  NOR U6211 ( .A(n5975), .B(n5974), .Z(n6478) );
  XOR U6212 ( .A(n5977), .B(n5976), .Z(n6477) );
  NOR U6213 ( .A(n6478), .B(n6477), .Z(n5978) );
  NOR U6214 ( .A(n5979), .B(n5978), .Z(n6474) );
  XOR U6215 ( .A(n5981), .B(n5980), .Z(n6473) );
  NOR U6216 ( .A(n6474), .B(n6473), .Z(n5982) );
  NOR U6217 ( .A(n5983), .B(n5982), .Z(n6522) );
  XOR U6218 ( .A(n5985), .B(n5984), .Z(n6521) );
  NOR U6219 ( .A(n6522), .B(n6521), .Z(n5986) );
  NOR U6220 ( .A(n5987), .B(n5986), .Z(n6471) );
  XOR U6221 ( .A(n5989), .B(n5988), .Z(n6470) );
  NOR U6222 ( .A(n6471), .B(n6470), .Z(n5990) );
  NOR U6223 ( .A(n5991), .B(n5990), .Z(n6467) );
  IV U6224 ( .A(n6467), .Z(n5992) );
  NOR U6225 ( .A(n5993), .B(n5992), .Z(n5994) );
  NOR U6226 ( .A(n5995), .B(n5994), .Z(n5996) );
  IV U6227 ( .A(n5996), .Z(n6003) );
  NOR U6228 ( .A(n100), .B(n121), .Z(n6002) );
  IV U6229 ( .A(n6002), .Z(n5997) );
  NOR U6230 ( .A(n6003), .B(n5997), .Z(n6005) );
  XOR U6231 ( .A(n5999), .B(n5998), .Z(n6000) );
  XOR U6232 ( .A(n6001), .B(n6000), .Z(n6460) );
  XOR U6233 ( .A(n6003), .B(n6002), .Z(n6461) );
  NOR U6234 ( .A(n6460), .B(n6461), .Z(n6004) );
  NOR U6235 ( .A(n6005), .B(n6004), .Z(n6543) );
  IV U6236 ( .A(n6543), .Z(n6006) );
  NOR U6237 ( .A(n6007), .B(n6006), .Z(n6008) );
  NOR U6238 ( .A(n6009), .B(n6008), .Z(n6010) );
  IV U6239 ( .A(n6010), .Z(n6015) );
  NOR U6240 ( .A(n102), .B(n121), .Z(n6014) );
  IV U6241 ( .A(n6014), .Z(n6011) );
  NOR U6242 ( .A(n6015), .B(n6011), .Z(n6018) );
  XOR U6243 ( .A(n6013), .B(n6012), .Z(n6457) );
  IV U6244 ( .A(n6457), .Z(n6016) );
  XOR U6245 ( .A(n6015), .B(n6014), .Z(n6458) );
  NOR U6246 ( .A(n6016), .B(n6458), .Z(n6017) );
  NOR U6247 ( .A(n6018), .B(n6017), .Z(n6553) );
  XOR U6248 ( .A(n6020), .B(n6019), .Z(n6554) );
  IV U6249 ( .A(n6554), .Z(n6021) );
  NOR U6250 ( .A(n6553), .B(n6021), .Z(n6022) );
  NOR U6251 ( .A(n6023), .B(n6022), .Z(n6453) );
  XOR U6252 ( .A(n6025), .B(n6024), .Z(n6454) );
  NOR U6253 ( .A(n6453), .B(n6454), .Z(n6026) );
  NOR U6254 ( .A(n6027), .B(n6026), .Z(n6449) );
  XOR U6255 ( .A(n6029), .B(n6028), .Z(n6450) );
  NOR U6256 ( .A(n6449), .B(n6450), .Z(n6030) );
  NOR U6257 ( .A(n6031), .B(n6030), .Z(n6447) );
  XOR U6258 ( .A(n6033), .B(n6032), .Z(n6448) );
  NOR U6259 ( .A(n6447), .B(n6448), .Z(n6034) );
  NOR U6260 ( .A(n6035), .B(n6034), .Z(n6574) );
  XOR U6261 ( .A(n6037), .B(n6036), .Z(n6573) );
  NOR U6262 ( .A(n6574), .B(n6573), .Z(n6038) );
  NOR U6263 ( .A(n6039), .B(n6038), .Z(n6443) );
  XOR U6264 ( .A(n6041), .B(n6040), .Z(n6444) );
  NOR U6265 ( .A(n6443), .B(n6444), .Z(n6042) );
  NOR U6266 ( .A(n6043), .B(n6042), .Z(n6440) );
  XOR U6267 ( .A(n6045), .B(n6044), .Z(n6439) );
  NOR U6268 ( .A(n6440), .B(n6439), .Z(n6046) );
  NOR U6269 ( .A(n6047), .B(n6046), .Z(n6435) );
  XOR U6270 ( .A(n6049), .B(n6048), .Z(n6436) );
  NOR U6271 ( .A(n6435), .B(n6436), .Z(n6050) );
  NOR U6272 ( .A(n6051), .B(n6050), .Z(n6431) );
  XOR U6273 ( .A(n6053), .B(n6052), .Z(n6432) );
  NOR U6274 ( .A(n6431), .B(n6432), .Z(n6054) );
  NOR U6275 ( .A(n6055), .B(n6054), .Z(n6427) );
  XOR U6276 ( .A(n6057), .B(n6056), .Z(n6428) );
  NOR U6277 ( .A(n6427), .B(n6428), .Z(n6058) );
  NOR U6278 ( .A(n6059), .B(n6058), .Z(n6423) );
  XOR U6279 ( .A(n6061), .B(n6060), .Z(n6424) );
  NOR U6280 ( .A(n6423), .B(n6424), .Z(n6062) );
  NOR U6281 ( .A(n6063), .B(n6062), .Z(n6419) );
  XOR U6282 ( .A(n6065), .B(n6064), .Z(n6420) );
  NOR U6283 ( .A(n6419), .B(n6420), .Z(n6066) );
  NOR U6284 ( .A(n6067), .B(n6066), .Z(n6415) );
  XOR U6285 ( .A(n6069), .B(n6068), .Z(n6416) );
  NOR U6286 ( .A(n6415), .B(n6416), .Z(n6070) );
  NOR U6287 ( .A(n6071), .B(n6070), .Z(n6411) );
  XOR U6288 ( .A(n6073), .B(n6072), .Z(n6412) );
  NOR U6289 ( .A(n6411), .B(n6412), .Z(n6074) );
  NOR U6290 ( .A(n6075), .B(n6074), .Z(n6407) );
  XOR U6291 ( .A(n6077), .B(n6076), .Z(n6408) );
  NOR U6292 ( .A(n6407), .B(n6408), .Z(n6078) );
  NOR U6293 ( .A(n6079), .B(n6078), .Z(n6403) );
  XOR U6294 ( .A(n6081), .B(n6080), .Z(n6404) );
  NOR U6295 ( .A(n6403), .B(n6404), .Z(n6082) );
  NOR U6296 ( .A(n6083), .B(n6082), .Z(n6399) );
  XOR U6297 ( .A(n6085), .B(n6084), .Z(n6400) );
  NOR U6298 ( .A(n6399), .B(n6400), .Z(n6086) );
  NOR U6299 ( .A(n6087), .B(n6086), .Z(n6395) );
  XOR U6300 ( .A(n6089), .B(n6088), .Z(n6396) );
  NOR U6301 ( .A(n6395), .B(n6396), .Z(n6090) );
  NOR U6302 ( .A(n6091), .B(n6090), .Z(n6391) );
  XOR U6303 ( .A(n6093), .B(n6092), .Z(n6392) );
  NOR U6304 ( .A(n6391), .B(n6392), .Z(n6094) );
  NOR U6305 ( .A(n6095), .B(n6094), .Z(n6387) );
  XOR U6306 ( .A(n6097), .B(n6096), .Z(n6388) );
  NOR U6307 ( .A(n6387), .B(n6388), .Z(n6098) );
  NOR U6308 ( .A(n6099), .B(n6098), .Z(n6383) );
  XOR U6309 ( .A(n6101), .B(n6100), .Z(n6384) );
  NOR U6310 ( .A(n6383), .B(n6384), .Z(n6102) );
  NOR U6311 ( .A(n6103), .B(n6102), .Z(n6379) );
  XOR U6312 ( .A(n6105), .B(n6104), .Z(n6380) );
  NOR U6313 ( .A(n6379), .B(n6380), .Z(n6106) );
  NOR U6314 ( .A(n6107), .B(n6106), .Z(n6375) );
  XOR U6315 ( .A(n6109), .B(n6108), .Z(n6376) );
  NOR U6316 ( .A(n6375), .B(n6376), .Z(n6110) );
  NOR U6317 ( .A(n6111), .B(n6110), .Z(n6371) );
  XOR U6318 ( .A(n6113), .B(n6112), .Z(n6372) );
  NOR U6319 ( .A(n6371), .B(n6372), .Z(n6114) );
  NOR U6320 ( .A(n6115), .B(n6114), .Z(n6367) );
  XOR U6321 ( .A(n6117), .B(n6116), .Z(n6368) );
  NOR U6322 ( .A(n6367), .B(n6368), .Z(n6118) );
  NOR U6323 ( .A(n6119), .B(n6118), .Z(n6363) );
  XOR U6324 ( .A(n6121), .B(n6120), .Z(n6364) );
  NOR U6325 ( .A(n6363), .B(n6364), .Z(n6122) );
  NOR U6326 ( .A(n6123), .B(n6122), .Z(n6359) );
  XOR U6327 ( .A(n6125), .B(n6124), .Z(n6360) );
  NOR U6328 ( .A(n6359), .B(n6360), .Z(n6126) );
  NOR U6329 ( .A(n6127), .B(n6126), .Z(n6355) );
  XOR U6330 ( .A(n6129), .B(n6128), .Z(n6356) );
  NOR U6331 ( .A(n6355), .B(n6356), .Z(n6130) );
  NOR U6332 ( .A(n6131), .B(n6130), .Z(n6351) );
  XOR U6333 ( .A(n6133), .B(n6132), .Z(n6352) );
  NOR U6334 ( .A(n6351), .B(n6352), .Z(n6134) );
  NOR U6335 ( .A(n6135), .B(n6134), .Z(n6350) );
  XOR U6336 ( .A(n6137), .B(n6136), .Z(n6349) );
  NOR U6337 ( .A(n6350), .B(n6349), .Z(n6138) );
  NOR U6338 ( .A(n6139), .B(n6138), .Z(n6343) );
  XOR U6339 ( .A(n6141), .B(n6140), .Z(n6344) );
  NOR U6340 ( .A(n6343), .B(n6344), .Z(n6142) );
  NOR U6341 ( .A(n6143), .B(n6142), .Z(n6342) );
  XOR U6342 ( .A(n6145), .B(n6144), .Z(n6341) );
  NOR U6343 ( .A(n6342), .B(n6341), .Z(n6146) );
  NOR U6344 ( .A(n6147), .B(n6146), .Z(n6335) );
  XOR U6345 ( .A(n6149), .B(n6148), .Z(n6336) );
  NOR U6346 ( .A(n6335), .B(n6336), .Z(n6150) );
  NOR U6347 ( .A(n6151), .B(n6150), .Z(n6331) );
  XOR U6348 ( .A(n6153), .B(n6152), .Z(n6332) );
  NOR U6349 ( .A(n6331), .B(n6332), .Z(n6154) );
  NOR U6350 ( .A(n6155), .B(n6154), .Z(n6327) );
  XOR U6351 ( .A(n6157), .B(n6156), .Z(n6328) );
  NOR U6352 ( .A(n6327), .B(n6328), .Z(n6158) );
  NOR U6353 ( .A(n6159), .B(n6158), .Z(n6323) );
  XOR U6354 ( .A(n6161), .B(n6160), .Z(n6324) );
  NOR U6355 ( .A(n6323), .B(n6324), .Z(n6162) );
  NOR U6356 ( .A(n6163), .B(n6162), .Z(n6716) );
  IV U6357 ( .A(n6164), .Z(n6165) );
  NOR U6358 ( .A(n6166), .B(n6165), .Z(n6171) );
  IV U6359 ( .A(n6167), .Z(n6168) );
  NOR U6360 ( .A(n6169), .B(n6168), .Z(n6170) );
  NOR U6361 ( .A(n6171), .B(n6170), .Z(n6172) );
  IV U6362 ( .A(n6172), .Z(n6723) );
  NOR U6363 ( .A(n135), .B(n122), .Z(n6721) );
  NOR U6364 ( .A(n133), .B(n124), .Z(n6730) );
  NOR U6365 ( .A(n6174), .B(n6173), .Z(n6179) );
  IV U6366 ( .A(n6175), .Z(n6177) );
  NOR U6367 ( .A(n6177), .B(n6176), .Z(n6178) );
  NOR U6368 ( .A(n6179), .B(n6178), .Z(n6726) );
  NOR U6369 ( .A(n6181), .B(n6180), .Z(n6185) );
  NOR U6370 ( .A(n6183), .B(n6182), .Z(n6184) );
  NOR U6371 ( .A(n6185), .B(n6184), .Z(n6738) );
  NOR U6372 ( .A(n131), .B(n127), .Z(n6735) );
  IV U6373 ( .A(n6186), .Z(n6187) );
  NOR U6374 ( .A(n6188), .B(n6187), .Z(n6192) );
  NOR U6375 ( .A(n6190), .B(n6189), .Z(n6191) );
  NOR U6376 ( .A(n6192), .B(n6191), .Z(n6751) );
  NOR U6377 ( .A(n126), .B(n130), .Z(n6749) );
  IV U6378 ( .A(n6749), .Z(n6315) );
  IV U6379 ( .A(n6193), .Z(n6195) );
  NOR U6380 ( .A(n6195), .B(n6194), .Z(n6199) );
  NOR U6381 ( .A(n6197), .B(n6196), .Z(n6198) );
  NOR U6382 ( .A(n6199), .B(n6198), .Z(n6200) );
  IV U6383 ( .A(n6200), .Z(n6874) );
  NOR U6384 ( .A(n125), .B(n132), .Z(n6872) );
  XOR U6385 ( .A(n6874), .B(n6872), .Z(n6875) );
  NOR U6386 ( .A(n6202), .B(n6201), .Z(n6207) );
  IV U6387 ( .A(n6203), .Z(n6204) );
  NOR U6388 ( .A(n6205), .B(n6204), .Z(n6206) );
  NOR U6389 ( .A(n6207), .B(n6206), .Z(n6757) );
  NOR U6390 ( .A(n123), .B(n134), .Z(n6755) );
  IV U6391 ( .A(n6755), .Z(n6314) );
  NOR U6392 ( .A(n6209), .B(n6208), .Z(n6213) );
  NOR U6393 ( .A(n6211), .B(n6210), .Z(n6212) );
  NOR U6394 ( .A(n6213), .B(n6212), .Z(n6770) );
  NOR U6395 ( .A(n119), .B(n138), .Z(n6768) );
  IV U6396 ( .A(n6768), .Z(n6305) );
  NOR U6397 ( .A(n6215), .B(n6214), .Z(n6220) );
  IV U6398 ( .A(n6216), .Z(n6218) );
  NOR U6399 ( .A(n6218), .B(n6217), .Z(n6219) );
  NOR U6400 ( .A(n6220), .B(n6219), .Z(n6221) );
  IV U6401 ( .A(n6221), .Z(n6775) );
  NOR U6402 ( .A(n79), .B(n140), .Z(n6773) );
  XOR U6403 ( .A(n6775), .B(n6773), .Z(n6776) );
  NOR U6404 ( .A(n6223), .B(n6222), .Z(n6228) );
  IV U6405 ( .A(n6224), .Z(n6225) );
  NOR U6406 ( .A(n6226), .B(n6225), .Z(n6227) );
  NOR U6407 ( .A(n6228), .B(n6227), .Z(n6783) );
  NOR U6408 ( .A(n117), .B(n142), .Z(n6781) );
  IV U6409 ( .A(n6781), .Z(n6304) );
  IV U6410 ( .A(n6229), .Z(n6230) );
  NOR U6411 ( .A(n6231), .B(n6230), .Z(n6235) );
  NOR U6412 ( .A(n6233), .B(n6232), .Z(n6234) );
  NOR U6413 ( .A(n6235), .B(n6234), .Z(n6790) );
  NOR U6414 ( .A(n6237), .B(n6236), .Z(n6241) );
  NOR U6415 ( .A(n6239), .B(n6238), .Z(n6240) );
  NOR U6416 ( .A(n6241), .B(n6240), .Z(n6797) );
  NOR U6417 ( .A(n116), .B(n146), .Z(n6795) );
  NOR U6418 ( .A(n81), .B(n149), .Z(n6804) );
  IV U6419 ( .A(n6242), .Z(n6243) );
  NOR U6420 ( .A(n6244), .B(n6243), .Z(n6248) );
  NOR U6421 ( .A(n6246), .B(n6245), .Z(n6247) );
  NOR U6422 ( .A(n6248), .B(n6247), .Z(n6800) );
  NOR U6423 ( .A(n6250), .B(n6249), .Z(n6254) );
  NOR U6424 ( .A(n6252), .B(n6251), .Z(n6253) );
  NOR U6425 ( .A(n6254), .B(n6253), .Z(n6812) );
  NOR U6426 ( .A(n115), .B(n151), .Z(n6810) );
  NOR U6427 ( .A(n82), .B(n152), .Z(n6819) );
  IV U6428 ( .A(n6255), .Z(n6256) );
  NOR U6429 ( .A(n6257), .B(n6256), .Z(n6261) );
  NOR U6430 ( .A(n6259), .B(n6258), .Z(n6260) );
  NOR U6431 ( .A(n6261), .B(n6260), .Z(n6815) );
  NOR U6432 ( .A(n6263), .B(n6262), .Z(n6267) );
  NOR U6433 ( .A(n6265), .B(n6264), .Z(n6266) );
  NOR U6434 ( .A(n6267), .B(n6266), .Z(n6827) );
  NOR U6435 ( .A(n114), .B(n154), .Z(n6824) );
  NOR U6436 ( .A(n6269), .B(n6268), .Z(n6273) );
  NOR U6437 ( .A(n6271), .B(n6270), .Z(n6272) );
  NOR U6438 ( .A(n6273), .B(n6272), .Z(n6833) );
  NOR U6439 ( .A(n113), .B(n159), .Z(n6831) );
  NOR U6440 ( .A(n6275), .B(n6274), .Z(n6279) );
  NOR U6441 ( .A(n6277), .B(n6276), .Z(n6278) );
  NOR U6442 ( .A(n6279), .B(n6278), .Z(n6839) );
  NOR U6443 ( .A(n112), .B(n162), .Z(n6837) );
  IV U6444 ( .A(n6837), .Z(n6288) );
  IV U6445 ( .A(n6280), .Z(n6281) );
  NOR U6446 ( .A(n6282), .B(n6281), .Z(n6286) );
  NOR U6447 ( .A(n6284), .B(n6283), .Z(n6285) );
  NOR U6448 ( .A(n6286), .B(n6285), .Z(n6844) );
  NOR U6449 ( .A(n164), .B(n85), .Z(n6842) );
  XOR U6450 ( .A(n6844), .B(n6842), .Z(n6846) );
  NOR U6451 ( .A(n166), .B(n111), .Z(n6287) );
  IV U6452 ( .A(n6287), .Z(n6845) );
  XOR U6453 ( .A(n6846), .B(n6845), .Z(n6836) );
  XOR U6454 ( .A(n6288), .B(n6836), .Z(n6838) );
  XOR U6455 ( .A(n6839), .B(n6838), .Z(n6855) );
  IV U6456 ( .A(n6289), .Z(n6290) );
  NOR U6457 ( .A(n6291), .B(n6290), .Z(n6295) );
  NOR U6458 ( .A(n6293), .B(n6292), .Z(n6294) );
  NOR U6459 ( .A(n6295), .B(n6294), .Z(n6853) );
  NOR U6460 ( .A(n84), .B(n160), .Z(n6851) );
  XOR U6461 ( .A(n6853), .B(n6851), .Z(n6854) );
  XOR U6462 ( .A(n6855), .B(n6854), .Z(n6830) );
  XOR U6463 ( .A(n6831), .B(n6830), .Z(n6296) );
  IV U6464 ( .A(n6296), .Z(n6832) );
  XOR U6465 ( .A(n6833), .B(n6832), .Z(n6863) );
  NOR U6466 ( .A(n6298), .B(n6297), .Z(n6302) );
  NOR U6467 ( .A(n6300), .B(n6299), .Z(n6301) );
  NOR U6468 ( .A(n6302), .B(n6301), .Z(n6861) );
  NOR U6469 ( .A(n83), .B(n157), .Z(n6859) );
  XOR U6470 ( .A(n6861), .B(n6859), .Z(n6862) );
  XOR U6471 ( .A(n6863), .B(n6862), .Z(n6823) );
  XOR U6472 ( .A(n6824), .B(n6823), .Z(n6825) );
  XOR U6473 ( .A(n6827), .B(n6825), .Z(n6816) );
  XOR U6474 ( .A(n6815), .B(n6816), .Z(n6818) );
  XOR U6475 ( .A(n6819), .B(n6818), .Z(n6808) );
  XOR U6476 ( .A(n6810), .B(n6808), .Z(n6811) );
  XOR U6477 ( .A(n6812), .B(n6811), .Z(n6303) );
  IV U6478 ( .A(n6303), .Z(n6801) );
  XOR U6479 ( .A(n6800), .B(n6801), .Z(n6803) );
  XOR U6480 ( .A(n6804), .B(n6803), .Z(n6793) );
  XOR U6481 ( .A(n6795), .B(n6793), .Z(n6796) );
  XOR U6482 ( .A(n6797), .B(n6796), .Z(n6788) );
  NOR U6483 ( .A(n80), .B(n144), .Z(n6786) );
  XOR U6484 ( .A(n6788), .B(n6786), .Z(n6789) );
  XOR U6485 ( .A(n6790), .B(n6789), .Z(n6780) );
  XOR U6486 ( .A(n6304), .B(n6780), .Z(n6782) );
  XOR U6487 ( .A(n6783), .B(n6782), .Z(n6777) );
  XOR U6488 ( .A(n6776), .B(n6777), .Z(n6767) );
  XOR U6489 ( .A(n6305), .B(n6767), .Z(n6769) );
  XOR U6490 ( .A(n6770), .B(n6769), .Z(n6764) );
  NOR U6491 ( .A(n6307), .B(n6306), .Z(n6313) );
  IV U6492 ( .A(n6308), .Z(n6311) );
  IV U6493 ( .A(n6309), .Z(n6310) );
  NOR U6494 ( .A(n6311), .B(n6310), .Z(n6312) );
  NOR U6495 ( .A(n6313), .B(n6312), .Z(n6762) );
  NOR U6496 ( .A(n120), .B(n136), .Z(n6760) );
  XOR U6497 ( .A(n6762), .B(n6760), .Z(n6763) );
  XOR U6498 ( .A(n6764), .B(n6763), .Z(n6754) );
  XOR U6499 ( .A(n6314), .B(n6754), .Z(n6756) );
  XOR U6500 ( .A(n6757), .B(n6756), .Z(n6876) );
  XOR U6501 ( .A(n6875), .B(n6876), .Z(n6748) );
  XOR U6502 ( .A(n6315), .B(n6748), .Z(n6750) );
  XOR U6503 ( .A(n6751), .B(n6750), .Z(n6745) );
  IV U6504 ( .A(n6316), .Z(n6317) );
  NOR U6505 ( .A(n6318), .B(n6317), .Z(n6322) );
  NOR U6506 ( .A(n6320), .B(n6319), .Z(n6321) );
  NOR U6507 ( .A(n6322), .B(n6321), .Z(n6743) );
  NOR U6508 ( .A(n128), .B(n129), .Z(n6741) );
  XOR U6509 ( .A(n6743), .B(n6741), .Z(n6744) );
  XOR U6510 ( .A(n6745), .B(n6744), .Z(n6734) );
  XOR U6511 ( .A(n6735), .B(n6734), .Z(n6736) );
  XOR U6512 ( .A(n6738), .B(n6736), .Z(n6727) );
  XOR U6513 ( .A(n6726), .B(n6727), .Z(n6729) );
  XOR U6514 ( .A(n6730), .B(n6729), .Z(n6719) );
  XOR U6515 ( .A(n6721), .B(n6719), .Z(n6722) );
  XOR U6516 ( .A(n6723), .B(n6722), .Z(n6714) );
  NOR U6517 ( .A(n137), .B(n121), .Z(n6712) );
  XOR U6518 ( .A(n6714), .B(n6712), .Z(n6715) );
  XOR U6519 ( .A(n6716), .B(n6715), .Z(n6707) );
  NOR U6520 ( .A(n6708), .B(n6707), .Z(n6711) );
  IV U6521 ( .A(n6323), .Z(n6325) );
  XOR U6522 ( .A(n6325), .B(n6324), .Z(n6702) );
  NOR U6523 ( .A(n137), .B(n118), .Z(n6703) );
  IV U6524 ( .A(n6703), .Z(n6326) );
  NOR U6525 ( .A(n6702), .B(n6326), .Z(n6705) );
  IV U6526 ( .A(n6327), .Z(n6329) );
  XOR U6527 ( .A(n6329), .B(n6328), .Z(n6698) );
  NOR U6528 ( .A(n135), .B(n118), .Z(n6699) );
  IV U6529 ( .A(n6699), .Z(n6330) );
  NOR U6530 ( .A(n6698), .B(n6330), .Z(n6701) );
  IV U6531 ( .A(n6331), .Z(n6333) );
  XOR U6532 ( .A(n6333), .B(n6332), .Z(n6694) );
  NOR U6533 ( .A(n133), .B(n118), .Z(n6695) );
  IV U6534 ( .A(n6695), .Z(n6334) );
  NOR U6535 ( .A(n6694), .B(n6334), .Z(n6697) );
  IV U6536 ( .A(n6335), .Z(n6337) );
  XOR U6537 ( .A(n6337), .B(n6336), .Z(n6339) );
  NOR U6538 ( .A(n131), .B(n118), .Z(n6340) );
  IV U6539 ( .A(n6340), .Z(n6338) );
  NOR U6540 ( .A(n6339), .B(n6338), .Z(n6693) );
  XOR U6541 ( .A(n6340), .B(n6339), .Z(n6899) );
  NOR U6542 ( .A(n128), .B(n118), .Z(n6687) );
  XOR U6543 ( .A(n6342), .B(n6341), .Z(n6686) );
  NOR U6544 ( .A(n6687), .B(n6686), .Z(n6690) );
  IV U6545 ( .A(n6343), .Z(n6345) );
  XOR U6546 ( .A(n6345), .B(n6344), .Z(n6347) );
  NOR U6547 ( .A(n126), .B(n118), .Z(n6348) );
  IV U6548 ( .A(n6348), .Z(n6346) );
  NOR U6549 ( .A(n6347), .B(n6346), .Z(n6684) );
  XOR U6550 ( .A(n6348), .B(n6347), .Z(n6905) );
  NOR U6551 ( .A(n125), .B(n118), .Z(n6678) );
  XOR U6552 ( .A(n6350), .B(n6349), .Z(n6677) );
  NOR U6553 ( .A(n6678), .B(n6677), .Z(n6681) );
  IV U6554 ( .A(n6351), .Z(n6353) );
  XOR U6555 ( .A(n6353), .B(n6352), .Z(n6672) );
  NOR U6556 ( .A(n123), .B(n118), .Z(n6673) );
  IV U6557 ( .A(n6673), .Z(n6354) );
  NOR U6558 ( .A(n6672), .B(n6354), .Z(n6675) );
  IV U6559 ( .A(n6355), .Z(n6357) );
  XOR U6560 ( .A(n6357), .B(n6356), .Z(n6668) );
  NOR U6561 ( .A(n120), .B(n118), .Z(n6669) );
  IV U6562 ( .A(n6669), .Z(n6358) );
  NOR U6563 ( .A(n6668), .B(n6358), .Z(n6671) );
  IV U6564 ( .A(n6359), .Z(n6361) );
  XOR U6565 ( .A(n6361), .B(n6360), .Z(n6664) );
  NOR U6566 ( .A(n119), .B(n118), .Z(n6665) );
  IV U6567 ( .A(n6665), .Z(n6362) );
  NOR U6568 ( .A(n6664), .B(n6362), .Z(n6667) );
  IV U6569 ( .A(n6363), .Z(n6365) );
  XOR U6570 ( .A(n6365), .B(n6364), .Z(n6660) );
  NOR U6571 ( .A(n79), .B(n118), .Z(n6661) );
  IV U6572 ( .A(n6661), .Z(n6366) );
  NOR U6573 ( .A(n6660), .B(n6366), .Z(n6663) );
  IV U6574 ( .A(n6367), .Z(n6369) );
  XOR U6575 ( .A(n6369), .B(n6368), .Z(n6656) );
  NOR U6576 ( .A(n117), .B(n118), .Z(n6657) );
  IV U6577 ( .A(n6657), .Z(n6370) );
  NOR U6578 ( .A(n6656), .B(n6370), .Z(n6659) );
  IV U6579 ( .A(n6371), .Z(n6373) );
  XOR U6580 ( .A(n6373), .B(n6372), .Z(n6652) );
  NOR U6581 ( .A(n80), .B(n118), .Z(n6653) );
  IV U6582 ( .A(n6653), .Z(n6374) );
  NOR U6583 ( .A(n6652), .B(n6374), .Z(n6655) );
  IV U6584 ( .A(n6375), .Z(n6377) );
  XOR U6585 ( .A(n6377), .B(n6376), .Z(n6648) );
  NOR U6586 ( .A(n116), .B(n118), .Z(n6649) );
  IV U6587 ( .A(n6649), .Z(n6378) );
  NOR U6588 ( .A(n6648), .B(n6378), .Z(n6651) );
  IV U6589 ( .A(n6379), .Z(n6381) );
  XOR U6590 ( .A(n6381), .B(n6380), .Z(n6644) );
  NOR U6591 ( .A(n81), .B(n118), .Z(n6645) );
  IV U6592 ( .A(n6645), .Z(n6382) );
  NOR U6593 ( .A(n6644), .B(n6382), .Z(n6647) );
  IV U6594 ( .A(n6383), .Z(n6385) );
  XOR U6595 ( .A(n6385), .B(n6384), .Z(n6640) );
  NOR U6596 ( .A(n115), .B(n118), .Z(n6641) );
  IV U6597 ( .A(n6641), .Z(n6386) );
  NOR U6598 ( .A(n6640), .B(n6386), .Z(n6643) );
  IV U6599 ( .A(n6387), .Z(n6389) );
  XOR U6600 ( .A(n6389), .B(n6388), .Z(n6636) );
  NOR U6601 ( .A(n82), .B(n118), .Z(n6637) );
  IV U6602 ( .A(n6637), .Z(n6390) );
  NOR U6603 ( .A(n6636), .B(n6390), .Z(n6639) );
  IV U6604 ( .A(n6391), .Z(n6393) );
  XOR U6605 ( .A(n6393), .B(n6392), .Z(n6632) );
  NOR U6606 ( .A(n114), .B(n118), .Z(n6633) );
  IV U6607 ( .A(n6633), .Z(n6394) );
  NOR U6608 ( .A(n6632), .B(n6394), .Z(n6635) );
  IV U6609 ( .A(n6395), .Z(n6397) );
  XOR U6610 ( .A(n6397), .B(n6396), .Z(n6628) );
  NOR U6611 ( .A(n83), .B(n118), .Z(n6629) );
  IV U6612 ( .A(n6629), .Z(n6398) );
  NOR U6613 ( .A(n6628), .B(n6398), .Z(n6631) );
  IV U6614 ( .A(n6399), .Z(n6401) );
  XOR U6615 ( .A(n6401), .B(n6400), .Z(n6624) );
  NOR U6616 ( .A(n113), .B(n118), .Z(n6625) );
  IV U6617 ( .A(n6625), .Z(n6402) );
  NOR U6618 ( .A(n6624), .B(n6402), .Z(n6627) );
  IV U6619 ( .A(n6403), .Z(n6405) );
  XOR U6620 ( .A(n6405), .B(n6404), .Z(n6620) );
  NOR U6621 ( .A(n84), .B(n118), .Z(n6621) );
  IV U6622 ( .A(n6621), .Z(n6406) );
  NOR U6623 ( .A(n6620), .B(n6406), .Z(n6623) );
  IV U6624 ( .A(n6407), .Z(n6409) );
  XOR U6625 ( .A(n6409), .B(n6408), .Z(n6616) );
  NOR U6626 ( .A(n112), .B(n118), .Z(n6617) );
  IV U6627 ( .A(n6617), .Z(n6410) );
  NOR U6628 ( .A(n6616), .B(n6410), .Z(n6619) );
  IV U6629 ( .A(n6411), .Z(n6413) );
  XOR U6630 ( .A(n6413), .B(n6412), .Z(n6612) );
  NOR U6631 ( .A(n85), .B(n118), .Z(n6613) );
  IV U6632 ( .A(n6613), .Z(n6414) );
  NOR U6633 ( .A(n6612), .B(n6414), .Z(n6615) );
  XOR U6634 ( .A(n6416), .B(n6415), .Z(n6417) );
  IV U6635 ( .A(n6417), .Z(n6608) );
  NOR U6636 ( .A(n111), .B(n118), .Z(n6609) );
  IV U6637 ( .A(n6609), .Z(n6418) );
  NOR U6638 ( .A(n6608), .B(n6418), .Z(n6611) );
  XOR U6639 ( .A(n6420), .B(n6419), .Z(n6421) );
  IV U6640 ( .A(n6421), .Z(n6604) );
  NOR U6641 ( .A(n86), .B(n118), .Z(n6605) );
  IV U6642 ( .A(n6605), .Z(n6422) );
  NOR U6643 ( .A(n6604), .B(n6422), .Z(n6607) );
  XOR U6644 ( .A(n6424), .B(n6423), .Z(n6425) );
  IV U6645 ( .A(n6425), .Z(n6600) );
  NOR U6646 ( .A(n110), .B(n118), .Z(n6601) );
  IV U6647 ( .A(n6601), .Z(n6426) );
  NOR U6648 ( .A(n6600), .B(n6426), .Z(n6603) );
  XOR U6649 ( .A(n6428), .B(n6427), .Z(n6429) );
  IV U6650 ( .A(n6429), .Z(n6596) );
  NOR U6651 ( .A(n109), .B(n118), .Z(n6597) );
  IV U6652 ( .A(n6597), .Z(n6430) );
  NOR U6653 ( .A(n6596), .B(n6430), .Z(n6599) );
  XOR U6654 ( .A(n6432), .B(n6431), .Z(n6433) );
  IV U6655 ( .A(n6433), .Z(n6592) );
  NOR U6656 ( .A(n108), .B(n118), .Z(n6593) );
  IV U6657 ( .A(n6593), .Z(n6434) );
  NOR U6658 ( .A(n6592), .B(n6434), .Z(n6595) );
  XOR U6659 ( .A(n6436), .B(n6435), .Z(n6437) );
  IV U6660 ( .A(n6437), .Z(n6588) );
  NOR U6661 ( .A(n87), .B(n118), .Z(n6589) );
  IV U6662 ( .A(n6589), .Z(n6438) );
  NOR U6663 ( .A(n6588), .B(n6438), .Z(n6591) );
  IV U6664 ( .A(n6439), .Z(n6441) );
  XOR U6665 ( .A(n6441), .B(n6440), .Z(n6584) );
  NOR U6666 ( .A(n107), .B(n118), .Z(n6585) );
  IV U6667 ( .A(n6585), .Z(n6442) );
  NOR U6668 ( .A(n6584), .B(n6442), .Z(n6587) );
  NOR U6669 ( .A(n88), .B(n118), .Z(n6581) );
  IV U6670 ( .A(n6581), .Z(n6446) );
  XOR U6671 ( .A(n6444), .B(n6443), .Z(n6445) );
  IV U6672 ( .A(n6445), .Z(n6580) );
  NOR U6673 ( .A(n6446), .B(n6580), .Z(n6583) );
  XOR U6674 ( .A(n6448), .B(n6447), .Z(n6568) );
  IV U6675 ( .A(n6568), .Z(n7005) );
  NOR U6676 ( .A(n105), .B(n118), .Z(n6567) );
  IV U6677 ( .A(n6567), .Z(n7004) );
  NOR U6678 ( .A(n7005), .B(n7004), .Z(n6571) );
  XOR U6679 ( .A(n6450), .B(n6449), .Z(n6451) );
  IV U6680 ( .A(n6451), .Z(n6563) );
  NOR U6681 ( .A(n104), .B(n118), .Z(n6564) );
  IV U6682 ( .A(n6564), .Z(n6452) );
  NOR U6683 ( .A(n6563), .B(n6452), .Z(n6566) );
  NOR U6684 ( .A(n89), .B(n118), .Z(n6560) );
  IV U6685 ( .A(n6560), .Z(n6456) );
  XOR U6686 ( .A(n6454), .B(n6453), .Z(n6455) );
  IV U6687 ( .A(n6455), .Z(n6559) );
  NOR U6688 ( .A(n6456), .B(n6559), .Z(n6562) );
  NOR U6689 ( .A(n90), .B(n118), .Z(n6549) );
  IV U6690 ( .A(n6549), .Z(n6459) );
  XOR U6691 ( .A(n6458), .B(n6457), .Z(n6548) );
  NOR U6692 ( .A(n6459), .B(n6548), .Z(n6551) );
  XOR U6693 ( .A(n6461), .B(n6460), .Z(n6462) );
  NOR U6694 ( .A(n101), .B(n118), .Z(n6463) );
  NOR U6695 ( .A(n6462), .B(n6463), .Z(n6537) );
  IV U6696 ( .A(n6462), .Z(n7018) );
  IV U6697 ( .A(n6463), .Z(n7017) );
  NOR U6698 ( .A(n7018), .B(n7017), .Z(n6535) );
  XOR U6699 ( .A(n6465), .B(n6464), .Z(n6466) );
  XOR U6700 ( .A(n6467), .B(n6466), .Z(n6531) );
  NOR U6701 ( .A(n100), .B(n118), .Z(n6530) );
  IV U6702 ( .A(n6530), .Z(n6468) );
  NOR U6703 ( .A(n6531), .B(n6468), .Z(n6533) );
  NOR U6704 ( .A(n99), .B(n118), .Z(n6469) );
  IV U6705 ( .A(n6469), .Z(n6527) );
  XOR U6706 ( .A(n6471), .B(n6470), .Z(n6526) );
  IV U6707 ( .A(n6526), .Z(n6472) );
  NOR U6708 ( .A(n6527), .B(n6472), .Z(n6529) );
  XOR U6709 ( .A(n6474), .B(n6473), .Z(n6475) );
  NOR U6710 ( .A(n91), .B(n118), .Z(n6476) );
  NOR U6711 ( .A(n6475), .B(n6476), .Z(n6516) );
  IV U6712 ( .A(n6475), .Z(n7072) );
  IV U6713 ( .A(n6476), .Z(n7071) );
  NOR U6714 ( .A(n7072), .B(n7071), .Z(n6514) );
  IV U6715 ( .A(n6477), .Z(n6479) );
  XOR U6716 ( .A(n6479), .B(n6478), .Z(n6509) );
  NOR U6717 ( .A(n97), .B(n118), .Z(n6510) );
  IV U6718 ( .A(n6510), .Z(n6480) );
  NOR U6719 ( .A(n6509), .B(n6480), .Z(n6512) );
  XOR U6720 ( .A(n6482), .B(n6481), .Z(n6483) );
  IV U6721 ( .A(n6483), .Z(n6505) );
  NOR U6722 ( .A(n96), .B(n118), .Z(n6506) );
  IV U6723 ( .A(n6506), .Z(n6484) );
  NOR U6724 ( .A(n6505), .B(n6484), .Z(n6508) );
  NOR U6725 ( .A(n93), .B(n118), .Z(n7556) );
  IV U6726 ( .A(n7556), .Z(n6486) );
  NOR U6727 ( .A(n121), .B(n168), .Z(n6489) );
  IV U6728 ( .A(n6489), .Z(n6485) );
  NOR U6729 ( .A(n6486), .B(n6485), .Z(n6492) );
  IV U6730 ( .A(n6492), .Z(n6487) );
  NOR U6731 ( .A(n6488), .B(n6487), .Z(n6497) );
  XOR U6732 ( .A(n6490), .B(n6489), .Z(n6491) );
  NOR U6733 ( .A(n6492), .B(n6491), .Z(n6493) );
  NOR U6734 ( .A(n6497), .B(n6493), .Z(n6494) );
  IV U6735 ( .A(n6494), .Z(n7054) );
  NOR U6736 ( .A(n94), .B(n118), .Z(n7053) );
  IV U6737 ( .A(n7053), .Z(n6495) );
  NOR U6738 ( .A(n7054), .B(n6495), .Z(n6496) );
  NOR U6739 ( .A(n6497), .B(n6496), .Z(n6500) );
  NOR U6740 ( .A(n95), .B(n118), .Z(n6499) );
  IV U6741 ( .A(n6499), .Z(n6498) );
  NOR U6742 ( .A(n6500), .B(n6498), .Z(n6504) );
  XOR U6743 ( .A(n6500), .B(n6499), .Z(n7034) );
  XOR U6744 ( .A(n6502), .B(n6501), .Z(n7035) );
  NOR U6745 ( .A(n7034), .B(n7035), .Z(n6503) );
  NOR U6746 ( .A(n6504), .B(n6503), .Z(n7030) );
  XOR U6747 ( .A(n6506), .B(n6505), .Z(n7031) );
  NOR U6748 ( .A(n7030), .B(n7031), .Z(n6507) );
  NOR U6749 ( .A(n6508), .B(n6507), .Z(n7029) );
  XOR U6750 ( .A(n6510), .B(n6509), .Z(n7028) );
  NOR U6751 ( .A(n7029), .B(n7028), .Z(n6511) );
  NOR U6752 ( .A(n6512), .B(n6511), .Z(n7074) );
  IV U6753 ( .A(n7074), .Z(n6513) );
  NOR U6754 ( .A(n6514), .B(n6513), .Z(n6515) );
  NOR U6755 ( .A(n6516), .B(n6515), .Z(n6517) );
  IV U6756 ( .A(n6517), .Z(n6520) );
  NOR U6757 ( .A(n98), .B(n118), .Z(n6519) );
  IV U6758 ( .A(n6519), .Z(n6518) );
  NOR U6759 ( .A(n6520), .B(n6518), .Z(n6525) );
  XOR U6760 ( .A(n6520), .B(n6519), .Z(n7025) );
  XOR U6761 ( .A(n6522), .B(n6521), .Z(n6523) );
  IV U6762 ( .A(n6523), .Z(n7024) );
  NOR U6763 ( .A(n7025), .B(n7024), .Z(n6524) );
  NOR U6764 ( .A(n6525), .B(n6524), .Z(n7086) );
  XOR U6765 ( .A(n6527), .B(n6526), .Z(n7085) );
  NOR U6766 ( .A(n7086), .B(n7085), .Z(n6528) );
  NOR U6767 ( .A(n6529), .B(n6528), .Z(n7023) );
  XOR U6768 ( .A(n6531), .B(n6530), .Z(n7022) );
  NOR U6769 ( .A(n7023), .B(n7022), .Z(n6532) );
  NOR U6770 ( .A(n6533), .B(n6532), .Z(n7020) );
  IV U6771 ( .A(n7020), .Z(n6534) );
  NOR U6772 ( .A(n6535), .B(n6534), .Z(n6536) );
  NOR U6773 ( .A(n6537), .B(n6536), .Z(n6538) );
  IV U6774 ( .A(n6538), .Z(n6545) );
  NOR U6775 ( .A(n102), .B(n118), .Z(n6544) );
  IV U6776 ( .A(n6544), .Z(n6539) );
  NOR U6777 ( .A(n6545), .B(n6539), .Z(n6547) );
  XOR U6778 ( .A(n6541), .B(n6540), .Z(n6542) );
  XOR U6779 ( .A(n6543), .B(n6542), .Z(n7013) );
  XOR U6780 ( .A(n6545), .B(n6544), .Z(n7014) );
  NOR U6781 ( .A(n7013), .B(n7014), .Z(n6546) );
  NOR U6782 ( .A(n6547), .B(n6546), .Z(n7110) );
  XOR U6783 ( .A(n6549), .B(n6548), .Z(n7109) );
  NOR U6784 ( .A(n7110), .B(n7109), .Z(n6550) );
  NOR U6785 ( .A(n6551), .B(n6550), .Z(n6556) );
  NOR U6786 ( .A(n103), .B(n118), .Z(n6555) );
  IV U6787 ( .A(n6555), .Z(n6552) );
  NOR U6788 ( .A(n6556), .B(n6552), .Z(n6558) );
  XOR U6789 ( .A(n6554), .B(n6553), .Z(n7118) );
  XOR U6790 ( .A(n6556), .B(n6555), .Z(n7117) );
  NOR U6791 ( .A(n7118), .B(n7117), .Z(n6557) );
  NOR U6792 ( .A(n6558), .B(n6557), .Z(n7126) );
  XOR U6793 ( .A(n6560), .B(n6559), .Z(n7125) );
  NOR U6794 ( .A(n7126), .B(n7125), .Z(n6561) );
  NOR U6795 ( .A(n6562), .B(n6561), .Z(n7010) );
  XOR U6796 ( .A(n6564), .B(n6563), .Z(n7009) );
  NOR U6797 ( .A(n7010), .B(n7009), .Z(n6565) );
  NOR U6798 ( .A(n6566), .B(n6565), .Z(n7007) );
  NOR U6799 ( .A(n6568), .B(n6567), .Z(n6569) );
  NOR U6800 ( .A(n7007), .B(n6569), .Z(n6570) );
  NOR U6801 ( .A(n6571), .B(n6570), .Z(n6576) );
  NOR U6802 ( .A(n106), .B(n118), .Z(n6577) );
  IV U6803 ( .A(n6577), .Z(n6572) );
  NOR U6804 ( .A(n6576), .B(n6572), .Z(n6579) );
  XOR U6805 ( .A(n6574), .B(n6573), .Z(n6575) );
  IV U6806 ( .A(n6575), .Z(n7001) );
  XOR U6807 ( .A(n6577), .B(n6576), .Z(n7000) );
  NOR U6808 ( .A(n7001), .B(n7000), .Z(n6578) );
  NOR U6809 ( .A(n6579), .B(n6578), .Z(n7146) );
  XOR U6810 ( .A(n6581), .B(n6580), .Z(n7147) );
  NOR U6811 ( .A(n7146), .B(n7147), .Z(n6582) );
  NOR U6812 ( .A(n6583), .B(n6582), .Z(n7152) );
  XOR U6813 ( .A(n6585), .B(n6584), .Z(n7153) );
  NOR U6814 ( .A(n7152), .B(n7153), .Z(n6586) );
  NOR U6815 ( .A(n6587), .B(n6586), .Z(n6997) );
  XOR U6816 ( .A(n6589), .B(n6588), .Z(n6996) );
  NOR U6817 ( .A(n6997), .B(n6996), .Z(n6590) );
  NOR U6818 ( .A(n6591), .B(n6590), .Z(n6992) );
  XOR U6819 ( .A(n6593), .B(n6592), .Z(n6993) );
  NOR U6820 ( .A(n6992), .B(n6993), .Z(n6594) );
  NOR U6821 ( .A(n6595), .B(n6594), .Z(n6989) );
  XOR U6822 ( .A(n6597), .B(n6596), .Z(n6988) );
  NOR U6823 ( .A(n6989), .B(n6988), .Z(n6598) );
  NOR U6824 ( .A(n6599), .B(n6598), .Z(n6984) );
  XOR U6825 ( .A(n6601), .B(n6600), .Z(n6985) );
  NOR U6826 ( .A(n6984), .B(n6985), .Z(n6602) );
  NOR U6827 ( .A(n6603), .B(n6602), .Z(n6980) );
  XOR U6828 ( .A(n6605), .B(n6604), .Z(n6981) );
  NOR U6829 ( .A(n6980), .B(n6981), .Z(n6606) );
  NOR U6830 ( .A(n6607), .B(n6606), .Z(n6976) );
  XOR U6831 ( .A(n6609), .B(n6608), .Z(n6975) );
  NOR U6832 ( .A(n6976), .B(n6975), .Z(n6610) );
  NOR U6833 ( .A(n6611), .B(n6610), .Z(n6972) );
  XOR U6834 ( .A(n6613), .B(n6612), .Z(n6971) );
  NOR U6835 ( .A(n6972), .B(n6971), .Z(n6614) );
  NOR U6836 ( .A(n6615), .B(n6614), .Z(n6967) );
  XOR U6837 ( .A(n6617), .B(n6616), .Z(n6968) );
  NOR U6838 ( .A(n6967), .B(n6968), .Z(n6618) );
  NOR U6839 ( .A(n6619), .B(n6618), .Z(n6963) );
  XOR U6840 ( .A(n6621), .B(n6620), .Z(n6964) );
  NOR U6841 ( .A(n6963), .B(n6964), .Z(n6622) );
  NOR U6842 ( .A(n6623), .B(n6622), .Z(n6959) );
  XOR U6843 ( .A(n6625), .B(n6624), .Z(n6960) );
  NOR U6844 ( .A(n6959), .B(n6960), .Z(n6626) );
  NOR U6845 ( .A(n6627), .B(n6626), .Z(n6956) );
  XOR U6846 ( .A(n6629), .B(n6628), .Z(n6955) );
  NOR U6847 ( .A(n6956), .B(n6955), .Z(n6630) );
  NOR U6848 ( .A(n6631), .B(n6630), .Z(n6951) );
  XOR U6849 ( .A(n6633), .B(n6632), .Z(n6952) );
  NOR U6850 ( .A(n6951), .B(n6952), .Z(n6634) );
  NOR U6851 ( .A(n6635), .B(n6634), .Z(n6947) );
  XOR U6852 ( .A(n6637), .B(n6636), .Z(n6948) );
  NOR U6853 ( .A(n6947), .B(n6948), .Z(n6638) );
  NOR U6854 ( .A(n6639), .B(n6638), .Z(n6943) );
  XOR U6855 ( .A(n6641), .B(n6640), .Z(n6944) );
  NOR U6856 ( .A(n6943), .B(n6944), .Z(n6642) );
  NOR U6857 ( .A(n6643), .B(n6642), .Z(n6939) );
  XOR U6858 ( .A(n6645), .B(n6644), .Z(n6940) );
  NOR U6859 ( .A(n6939), .B(n6940), .Z(n6646) );
  NOR U6860 ( .A(n6647), .B(n6646), .Z(n6935) );
  XOR U6861 ( .A(n6649), .B(n6648), .Z(n6936) );
  NOR U6862 ( .A(n6935), .B(n6936), .Z(n6650) );
  NOR U6863 ( .A(n6651), .B(n6650), .Z(n6931) );
  XOR U6864 ( .A(n6653), .B(n6652), .Z(n6932) );
  NOR U6865 ( .A(n6931), .B(n6932), .Z(n6654) );
  NOR U6866 ( .A(n6655), .B(n6654), .Z(n6928) );
  XOR U6867 ( .A(n6657), .B(n6656), .Z(n6927) );
  NOR U6868 ( .A(n6928), .B(n6927), .Z(n6658) );
  NOR U6869 ( .A(n6659), .B(n6658), .Z(n6923) );
  XOR U6870 ( .A(n6661), .B(n6660), .Z(n6924) );
  NOR U6871 ( .A(n6923), .B(n6924), .Z(n6662) );
  NOR U6872 ( .A(n6663), .B(n6662), .Z(n6919) );
  XOR U6873 ( .A(n6665), .B(n6664), .Z(n6920) );
  NOR U6874 ( .A(n6919), .B(n6920), .Z(n6666) );
  NOR U6875 ( .A(n6667), .B(n6666), .Z(n6916) );
  XOR U6876 ( .A(n6669), .B(n6668), .Z(n6915) );
  NOR U6877 ( .A(n6916), .B(n6915), .Z(n6670) );
  NOR U6878 ( .A(n6671), .B(n6670), .Z(n6912) );
  XOR U6879 ( .A(n6673), .B(n6672), .Z(n6911) );
  NOR U6880 ( .A(n6912), .B(n6911), .Z(n6674) );
  NOR U6881 ( .A(n6675), .B(n6674), .Z(n6676) );
  IV U6882 ( .A(n6676), .Z(n6909) );
  XOR U6883 ( .A(n6678), .B(n6677), .Z(n6679) );
  IV U6884 ( .A(n6679), .Z(n6908) );
  NOR U6885 ( .A(n6909), .B(n6908), .Z(n6680) );
  NOR U6886 ( .A(n6681), .B(n6680), .Z(n6906) );
  IV U6887 ( .A(n6906), .Z(n6682) );
  NOR U6888 ( .A(n6905), .B(n6682), .Z(n6683) );
  NOR U6889 ( .A(n6684), .B(n6683), .Z(n6685) );
  IV U6890 ( .A(n6685), .Z(n6903) );
  XOR U6891 ( .A(n6687), .B(n6686), .Z(n6688) );
  IV U6892 ( .A(n6688), .Z(n6902) );
  NOR U6893 ( .A(n6903), .B(n6902), .Z(n6689) );
  NOR U6894 ( .A(n6690), .B(n6689), .Z(n6900) );
  IV U6895 ( .A(n6900), .Z(n6691) );
  NOR U6896 ( .A(n6899), .B(n6691), .Z(n6692) );
  NOR U6897 ( .A(n6693), .B(n6692), .Z(n6896) );
  XOR U6898 ( .A(n6695), .B(n6694), .Z(n6895) );
  NOR U6899 ( .A(n6896), .B(n6895), .Z(n6696) );
  NOR U6900 ( .A(n6697), .B(n6696), .Z(n6892) );
  XOR U6901 ( .A(n6699), .B(n6698), .Z(n6891) );
  NOR U6902 ( .A(n6892), .B(n6891), .Z(n6700) );
  NOR U6903 ( .A(n6701), .B(n6700), .Z(n6888) );
  XOR U6904 ( .A(n6703), .B(n6702), .Z(n6887) );
  NOR U6905 ( .A(n6888), .B(n6887), .Z(n6704) );
  NOR U6906 ( .A(n6705), .B(n6704), .Z(n6706) );
  IV U6907 ( .A(n6706), .Z(n6885) );
  XOR U6908 ( .A(n6708), .B(n6707), .Z(n6709) );
  IV U6909 ( .A(n6709), .Z(n6884) );
  NOR U6910 ( .A(n6885), .B(n6884), .Z(n6710) );
  NOR U6911 ( .A(n6711), .B(n6710), .Z(n7449) );
  NOR U6912 ( .A(n141), .B(n118), .Z(n7446) );
  IV U6913 ( .A(n6712), .Z(n6713) );
  NOR U6914 ( .A(n6714), .B(n6713), .Z(n6718) );
  NOR U6915 ( .A(n6716), .B(n6715), .Z(n6717) );
  NOR U6916 ( .A(n6718), .B(n6717), .Z(n7287) );
  IV U6917 ( .A(n7287), .Z(n6882) );
  IV U6918 ( .A(n6719), .Z(n6720) );
  NOR U6919 ( .A(n6721), .B(n6720), .Z(n6725) );
  NOR U6920 ( .A(n6723), .B(n6722), .Z(n6724) );
  NOR U6921 ( .A(n6725), .B(n6724), .Z(n7293) );
  NOR U6922 ( .A(n137), .B(n122), .Z(n7291) );
  IV U6923 ( .A(n7291), .Z(n6881) );
  IV U6924 ( .A(n6726), .Z(n6728) );
  NOR U6925 ( .A(n6728), .B(n6727), .Z(n6732) );
  NOR U6926 ( .A(n6730), .B(n6729), .Z(n6731) );
  NOR U6927 ( .A(n6732), .B(n6731), .Z(n6733) );
  IV U6928 ( .A(n6733), .Z(n7300) );
  NOR U6929 ( .A(n6735), .B(n6734), .Z(n6740) );
  IV U6930 ( .A(n6736), .Z(n6737) );
  NOR U6931 ( .A(n6738), .B(n6737), .Z(n6739) );
  NOR U6932 ( .A(n6740), .B(n6739), .Z(n7306) );
  NOR U6933 ( .A(n133), .B(n127), .Z(n7304) );
  IV U6934 ( .A(n6741), .Z(n6742) );
  NOR U6935 ( .A(n6743), .B(n6742), .Z(n6747) );
  NOR U6936 ( .A(n6745), .B(n6744), .Z(n6746) );
  NOR U6937 ( .A(n6747), .B(n6746), .Z(n7313) );
  NOR U6938 ( .A(n6749), .B(n6748), .Z(n6753) );
  NOR U6939 ( .A(n6751), .B(n6750), .Z(n6752) );
  NOR U6940 ( .A(n6753), .B(n6752), .Z(n7319) );
  NOR U6941 ( .A(n128), .B(n130), .Z(n7317) );
  NOR U6942 ( .A(n6755), .B(n6754), .Z(n6759) );
  NOR U6943 ( .A(n6757), .B(n6756), .Z(n6758) );
  NOR U6944 ( .A(n6759), .B(n6758), .Z(n7332) );
  NOR U6945 ( .A(n125), .B(n134), .Z(n7330) );
  IV U6946 ( .A(n6760), .Z(n6761) );
  NOR U6947 ( .A(n6762), .B(n6761), .Z(n6766) );
  NOR U6948 ( .A(n6764), .B(n6763), .Z(n6765) );
  NOR U6949 ( .A(n6766), .B(n6765), .Z(n7339) );
  NOR U6950 ( .A(n6768), .B(n6767), .Z(n6772) );
  NOR U6951 ( .A(n6770), .B(n6769), .Z(n6771) );
  NOR U6952 ( .A(n6772), .B(n6771), .Z(n7345) );
  NOR U6953 ( .A(n120), .B(n138), .Z(n7343) );
  IV U6954 ( .A(n7343), .Z(n6870) );
  IV U6955 ( .A(n6773), .Z(n6774) );
  NOR U6956 ( .A(n6775), .B(n6774), .Z(n6779) );
  NOR U6957 ( .A(n6777), .B(n6776), .Z(n6778) );
  NOR U6958 ( .A(n6779), .B(n6778), .Z(n7350) );
  NOR U6959 ( .A(n119), .B(n140), .Z(n7349) );
  NOR U6960 ( .A(n6781), .B(n6780), .Z(n6785) );
  NOR U6961 ( .A(n6783), .B(n6782), .Z(n6784) );
  NOR U6962 ( .A(n6785), .B(n6784), .Z(n7360) );
  NOR U6963 ( .A(n79), .B(n142), .Z(n7357) );
  IV U6964 ( .A(n6786), .Z(n6787) );
  NOR U6965 ( .A(n6788), .B(n6787), .Z(n6792) );
  NOR U6966 ( .A(n6790), .B(n6789), .Z(n6791) );
  NOR U6967 ( .A(n6792), .B(n6791), .Z(n7438) );
  IV U6968 ( .A(n6793), .Z(n6794) );
  NOR U6969 ( .A(n6795), .B(n6794), .Z(n6799) );
  NOR U6970 ( .A(n6797), .B(n6796), .Z(n6798) );
  NOR U6971 ( .A(n6799), .B(n6798), .Z(n7366) );
  NOR U6972 ( .A(n80), .B(n146), .Z(n7364) );
  IV U6973 ( .A(n7364), .Z(n6868) );
  IV U6974 ( .A(n6800), .Z(n6802) );
  NOR U6975 ( .A(n6802), .B(n6801), .Z(n6806) );
  NOR U6976 ( .A(n6804), .B(n6803), .Z(n6805) );
  NOR U6977 ( .A(n6806), .B(n6805), .Z(n6807) );
  IV U6978 ( .A(n6807), .Z(n7430) );
  IV U6979 ( .A(n6808), .Z(n6809) );
  NOR U6980 ( .A(n6810), .B(n6809), .Z(n6814) );
  NOR U6981 ( .A(n6812), .B(n6811), .Z(n6813) );
  NOR U6982 ( .A(n6814), .B(n6813), .Z(n7372) );
  NOR U6983 ( .A(n81), .B(n151), .Z(n7370) );
  IV U6984 ( .A(n7370), .Z(n6867) );
  IV U6985 ( .A(n6815), .Z(n6817) );
  NOR U6986 ( .A(n6817), .B(n6816), .Z(n6821) );
  NOR U6987 ( .A(n6819), .B(n6818), .Z(n6820) );
  NOR U6988 ( .A(n6821), .B(n6820), .Z(n6822) );
  IV U6989 ( .A(n6822), .Z(n7420) );
  NOR U6990 ( .A(n115), .B(n152), .Z(n7418) );
  XOR U6991 ( .A(n7420), .B(n7418), .Z(n7421) );
  NOR U6992 ( .A(n6824), .B(n6823), .Z(n6829) );
  IV U6993 ( .A(n6825), .Z(n6826) );
  NOR U6994 ( .A(n6827), .B(n6826), .Z(n6828) );
  NOR U6995 ( .A(n6829), .B(n6828), .Z(n7378) );
  NOR U6996 ( .A(n82), .B(n154), .Z(n7376) );
  IV U6997 ( .A(n7376), .Z(n6866) );
  NOR U6998 ( .A(n6831), .B(n6830), .Z(n6835) );
  NOR U6999 ( .A(n6833), .B(n6832), .Z(n6834) );
  NOR U7000 ( .A(n6835), .B(n6834), .Z(n7391) );
  NOR U7001 ( .A(n83), .B(n159), .Z(n7389) );
  NOR U7002 ( .A(n6837), .B(n6836), .Z(n6841) );
  NOR U7003 ( .A(n6839), .B(n6838), .Z(n6840) );
  NOR U7004 ( .A(n6841), .B(n6840), .Z(n7397) );
  NOR U7005 ( .A(n84), .B(n162), .Z(n7395) );
  IV U7006 ( .A(n7395), .Z(n6850) );
  IV U7007 ( .A(n6842), .Z(n6843) );
  NOR U7008 ( .A(n6844), .B(n6843), .Z(n6848) );
  NOR U7009 ( .A(n6846), .B(n6845), .Z(n6847) );
  NOR U7010 ( .A(n6848), .B(n6847), .Z(n7402) );
  NOR U7011 ( .A(n164), .B(n112), .Z(n7400) );
  XOR U7012 ( .A(n7402), .B(n7400), .Z(n7404) );
  NOR U7013 ( .A(n166), .B(n85), .Z(n6849) );
  IV U7014 ( .A(n6849), .Z(n7403) );
  XOR U7015 ( .A(n7404), .B(n7403), .Z(n7394) );
  XOR U7016 ( .A(n6850), .B(n7394), .Z(n7396) );
  XOR U7017 ( .A(n7397), .B(n7396), .Z(n7413) );
  IV U7018 ( .A(n6851), .Z(n6852) );
  NOR U7019 ( .A(n6853), .B(n6852), .Z(n6857) );
  NOR U7020 ( .A(n6855), .B(n6854), .Z(n6856) );
  NOR U7021 ( .A(n6857), .B(n6856), .Z(n7411) );
  NOR U7022 ( .A(n113), .B(n160), .Z(n7409) );
  XOR U7023 ( .A(n7411), .B(n7409), .Z(n7412) );
  XOR U7024 ( .A(n7413), .B(n7412), .Z(n7388) );
  XOR U7025 ( .A(n7389), .B(n7388), .Z(n6858) );
  IV U7026 ( .A(n6858), .Z(n7390) );
  XOR U7027 ( .A(n7391), .B(n7390), .Z(n7385) );
  IV U7028 ( .A(n6859), .Z(n6860) );
  NOR U7029 ( .A(n6861), .B(n6860), .Z(n6865) );
  NOR U7030 ( .A(n6863), .B(n6862), .Z(n6864) );
  NOR U7031 ( .A(n6865), .B(n6864), .Z(n7383) );
  NOR U7032 ( .A(n114), .B(n157), .Z(n7381) );
  XOR U7033 ( .A(n7383), .B(n7381), .Z(n7384) );
  XOR U7034 ( .A(n7385), .B(n7384), .Z(n7375) );
  XOR U7035 ( .A(n6866), .B(n7375), .Z(n7377) );
  XOR U7036 ( .A(n7378), .B(n7377), .Z(n7422) );
  XOR U7037 ( .A(n7421), .B(n7422), .Z(n7369) );
  XOR U7038 ( .A(n6867), .B(n7369), .Z(n7371) );
  XOR U7039 ( .A(n7372), .B(n7371), .Z(n7428) );
  NOR U7040 ( .A(n116), .B(n149), .Z(n7426) );
  XOR U7041 ( .A(n7428), .B(n7426), .Z(n7429) );
  XOR U7042 ( .A(n7430), .B(n7429), .Z(n7363) );
  XOR U7043 ( .A(n6868), .B(n7363), .Z(n7365) );
  XOR U7044 ( .A(n7366), .B(n7365), .Z(n7436) );
  NOR U7045 ( .A(n117), .B(n144), .Z(n7434) );
  XOR U7046 ( .A(n7436), .B(n7434), .Z(n7437) );
  XOR U7047 ( .A(n7438), .B(n7437), .Z(n7356) );
  XOR U7048 ( .A(n7357), .B(n7356), .Z(n7358) );
  XOR U7049 ( .A(n7360), .B(n7358), .Z(n7348) );
  XOR U7050 ( .A(n7349), .B(n7348), .Z(n6869) );
  IV U7051 ( .A(n6869), .Z(n7351) );
  XOR U7052 ( .A(n7350), .B(n7351), .Z(n7342) );
  XOR U7053 ( .A(n6870), .B(n7342), .Z(n7344) );
  XOR U7054 ( .A(n7345), .B(n7344), .Z(n7337) );
  NOR U7055 ( .A(n123), .B(n136), .Z(n7335) );
  XOR U7056 ( .A(n7337), .B(n7335), .Z(n7338) );
  XOR U7057 ( .A(n7339), .B(n7338), .Z(n7329) );
  XOR U7058 ( .A(n7330), .B(n7329), .Z(n6871) );
  IV U7059 ( .A(n6871), .Z(n7331) );
  XOR U7060 ( .A(n7332), .B(n7331), .Z(n7326) );
  IV U7061 ( .A(n6872), .Z(n6873) );
  NOR U7062 ( .A(n6874), .B(n6873), .Z(n6878) );
  NOR U7063 ( .A(n6876), .B(n6875), .Z(n6877) );
  NOR U7064 ( .A(n6878), .B(n6877), .Z(n7324) );
  NOR U7065 ( .A(n126), .B(n132), .Z(n7322) );
  XOR U7066 ( .A(n7324), .B(n7322), .Z(n7325) );
  XOR U7067 ( .A(n7326), .B(n7325), .Z(n7316) );
  XOR U7068 ( .A(n7317), .B(n7316), .Z(n6879) );
  IV U7069 ( .A(n6879), .Z(n7318) );
  XOR U7070 ( .A(n7319), .B(n7318), .Z(n7311) );
  NOR U7071 ( .A(n131), .B(n129), .Z(n7309) );
  XOR U7072 ( .A(n7311), .B(n7309), .Z(n7312) );
  XOR U7073 ( .A(n7313), .B(n7312), .Z(n7303) );
  XOR U7074 ( .A(n7304), .B(n7303), .Z(n6880) );
  IV U7075 ( .A(n6880), .Z(n7305) );
  XOR U7076 ( .A(n7306), .B(n7305), .Z(n7298) );
  NOR U7077 ( .A(n135), .B(n124), .Z(n7296) );
  XOR U7078 ( .A(n7298), .B(n7296), .Z(n7299) );
  XOR U7079 ( .A(n7300), .B(n7299), .Z(n7290) );
  XOR U7080 ( .A(n6881), .B(n7290), .Z(n7292) );
  XOR U7081 ( .A(n7293), .B(n7292), .Z(n7285) );
  NOR U7082 ( .A(n139), .B(n121), .Z(n7283) );
  XOR U7083 ( .A(n7285), .B(n7283), .Z(n7286) );
  XOR U7084 ( .A(n6882), .B(n7286), .Z(n7448) );
  XOR U7085 ( .A(n7446), .B(n7448), .Z(n7451) );
  XOR U7086 ( .A(n7449), .B(n7451), .Z(n7279) );
  NOR U7087 ( .A(n143), .B(n43), .Z(n7280) );
  IV U7088 ( .A(n7280), .Z(n6883) );
  NOR U7089 ( .A(n7279), .B(n6883), .Z(n7282) );
  XOR U7090 ( .A(n6885), .B(n6884), .Z(n7276) );
  NOR U7091 ( .A(n141), .B(n43), .Z(n7275) );
  IV U7092 ( .A(n7275), .Z(n6886) );
  NOR U7093 ( .A(n7276), .B(n6886), .Z(n7278) );
  XOR U7094 ( .A(n6888), .B(n6887), .Z(n7271) );
  IV U7095 ( .A(n7271), .Z(n6890) );
  NOR U7096 ( .A(n139), .B(n43), .Z(n6889) );
  IV U7097 ( .A(n6889), .Z(n7272) );
  NOR U7098 ( .A(n6890), .B(n7272), .Z(n7274) );
  XOR U7099 ( .A(n6892), .B(n6891), .Z(n7267) );
  IV U7100 ( .A(n7267), .Z(n6894) );
  NOR U7101 ( .A(n137), .B(n43), .Z(n6893) );
  IV U7102 ( .A(n6893), .Z(n7268) );
  NOR U7103 ( .A(n6894), .B(n7268), .Z(n7270) );
  XOR U7104 ( .A(n6896), .B(n6895), .Z(n7263) );
  IV U7105 ( .A(n7263), .Z(n6898) );
  NOR U7106 ( .A(n135), .B(n43), .Z(n6897) );
  IV U7107 ( .A(n6897), .Z(n7264) );
  NOR U7108 ( .A(n6898), .B(n7264), .Z(n7266) );
  XOR U7109 ( .A(n6900), .B(n6899), .Z(n7259) );
  NOR U7110 ( .A(n133), .B(n43), .Z(n7260) );
  IV U7111 ( .A(n7260), .Z(n6901) );
  NOR U7112 ( .A(n7259), .B(n6901), .Z(n7262) );
  XOR U7113 ( .A(n6903), .B(n6902), .Z(n7256) );
  NOR U7114 ( .A(n131), .B(n43), .Z(n7255) );
  IV U7115 ( .A(n7255), .Z(n6904) );
  NOR U7116 ( .A(n7256), .B(n6904), .Z(n7258) );
  XOR U7117 ( .A(n6906), .B(n6905), .Z(n7251) );
  NOR U7118 ( .A(n128), .B(n43), .Z(n7252) );
  IV U7119 ( .A(n7252), .Z(n6907) );
  NOR U7120 ( .A(n7251), .B(n6907), .Z(n7254) );
  XOR U7121 ( .A(n6909), .B(n6908), .Z(n7248) );
  NOR U7122 ( .A(n126), .B(n43), .Z(n7247) );
  IV U7123 ( .A(n7247), .Z(n6910) );
  NOR U7124 ( .A(n7248), .B(n6910), .Z(n7250) );
  XOR U7125 ( .A(n6912), .B(n6911), .Z(n7243) );
  IV U7126 ( .A(n7243), .Z(n6914) );
  NOR U7127 ( .A(n125), .B(n43), .Z(n6913) );
  IV U7128 ( .A(n6913), .Z(n7244) );
  NOR U7129 ( .A(n6914), .B(n7244), .Z(n7246) );
  XOR U7130 ( .A(n6916), .B(n6915), .Z(n7239) );
  IV U7131 ( .A(n7239), .Z(n6918) );
  NOR U7132 ( .A(n123), .B(n43), .Z(n6917) );
  IV U7133 ( .A(n6917), .Z(n7240) );
  NOR U7134 ( .A(n6918), .B(n7240), .Z(n7242) );
  IV U7135 ( .A(n6919), .Z(n6921) );
  XOR U7136 ( .A(n6921), .B(n6920), .Z(n7235) );
  NOR U7137 ( .A(n120), .B(n43), .Z(n7236) );
  IV U7138 ( .A(n7236), .Z(n6922) );
  NOR U7139 ( .A(n7235), .B(n6922), .Z(n7238) );
  IV U7140 ( .A(n6923), .Z(n6925) );
  XOR U7141 ( .A(n6925), .B(n6924), .Z(n7231) );
  NOR U7142 ( .A(n119), .B(n43), .Z(n7232) );
  IV U7143 ( .A(n7232), .Z(n6926) );
  NOR U7144 ( .A(n7231), .B(n6926), .Z(n7234) );
  XOR U7145 ( .A(n6928), .B(n6927), .Z(n7227) );
  IV U7146 ( .A(n7227), .Z(n6930) );
  NOR U7147 ( .A(n79), .B(n43), .Z(n6929) );
  IV U7148 ( .A(n6929), .Z(n7228) );
  NOR U7149 ( .A(n6930), .B(n7228), .Z(n7230) );
  IV U7150 ( .A(n6931), .Z(n6933) );
  XOR U7151 ( .A(n6933), .B(n6932), .Z(n7223) );
  NOR U7152 ( .A(n117), .B(n43), .Z(n7224) );
  IV U7153 ( .A(n7224), .Z(n6934) );
  NOR U7154 ( .A(n7223), .B(n6934), .Z(n7226) );
  IV U7155 ( .A(n6935), .Z(n6937) );
  XOR U7156 ( .A(n6937), .B(n6936), .Z(n7219) );
  NOR U7157 ( .A(n80), .B(n43), .Z(n7220) );
  IV U7158 ( .A(n7220), .Z(n6938) );
  NOR U7159 ( .A(n7219), .B(n6938), .Z(n7222) );
  IV U7160 ( .A(n6939), .Z(n6941) );
  XOR U7161 ( .A(n6941), .B(n6940), .Z(n7215) );
  NOR U7162 ( .A(n116), .B(n43), .Z(n7216) );
  IV U7163 ( .A(n7216), .Z(n6942) );
  NOR U7164 ( .A(n7215), .B(n6942), .Z(n7218) );
  IV U7165 ( .A(n6943), .Z(n6945) );
  XOR U7166 ( .A(n6945), .B(n6944), .Z(n7211) );
  NOR U7167 ( .A(n81), .B(n43), .Z(n7212) );
  IV U7168 ( .A(n7212), .Z(n6946) );
  NOR U7169 ( .A(n7211), .B(n6946), .Z(n7214) );
  IV U7170 ( .A(n6947), .Z(n6949) );
  XOR U7171 ( .A(n6949), .B(n6948), .Z(n7207) );
  NOR U7172 ( .A(n115), .B(n43), .Z(n7208) );
  IV U7173 ( .A(n7208), .Z(n6950) );
  NOR U7174 ( .A(n7207), .B(n6950), .Z(n7210) );
  IV U7175 ( .A(n6951), .Z(n6953) );
  XOR U7176 ( .A(n6953), .B(n6952), .Z(n7203) );
  NOR U7177 ( .A(n82), .B(n43), .Z(n7204) );
  IV U7178 ( .A(n7204), .Z(n6954) );
  NOR U7179 ( .A(n7203), .B(n6954), .Z(n7206) );
  XOR U7180 ( .A(n6956), .B(n6955), .Z(n7199) );
  IV U7181 ( .A(n7199), .Z(n6958) );
  NOR U7182 ( .A(n114), .B(n43), .Z(n6957) );
  IV U7183 ( .A(n6957), .Z(n7200) );
  NOR U7184 ( .A(n6958), .B(n7200), .Z(n7202) );
  IV U7185 ( .A(n6959), .Z(n6961) );
  XOR U7186 ( .A(n6961), .B(n6960), .Z(n7195) );
  NOR U7187 ( .A(n83), .B(n43), .Z(n7196) );
  IV U7188 ( .A(n7196), .Z(n6962) );
  NOR U7189 ( .A(n7195), .B(n6962), .Z(n7198) );
  IV U7190 ( .A(n6963), .Z(n6965) );
  XOR U7191 ( .A(n6965), .B(n6964), .Z(n7191) );
  NOR U7192 ( .A(n113), .B(n43), .Z(n7192) );
  IV U7193 ( .A(n7192), .Z(n6966) );
  NOR U7194 ( .A(n7191), .B(n6966), .Z(n7194) );
  IV U7195 ( .A(n6967), .Z(n6969) );
  XOR U7196 ( .A(n6969), .B(n6968), .Z(n7187) );
  NOR U7197 ( .A(n84), .B(n43), .Z(n7188) );
  IV U7198 ( .A(n7188), .Z(n6970) );
  NOR U7199 ( .A(n7187), .B(n6970), .Z(n7190) );
  XOR U7200 ( .A(n6972), .B(n6971), .Z(n7183) );
  IV U7201 ( .A(n7183), .Z(n6974) );
  NOR U7202 ( .A(n112), .B(n43), .Z(n6973) );
  IV U7203 ( .A(n6973), .Z(n7184) );
  NOR U7204 ( .A(n6974), .B(n7184), .Z(n7186) );
  XOR U7205 ( .A(n6976), .B(n6975), .Z(n6977) );
  NOR U7206 ( .A(n85), .B(n43), .Z(n6978) );
  NOR U7207 ( .A(n6977), .B(n6978), .Z(n7181) );
  XOR U7208 ( .A(n6978), .B(n6977), .Z(n6979) );
  IV U7209 ( .A(n6979), .Z(n7705) );
  XOR U7210 ( .A(n6981), .B(n6980), .Z(n6982) );
  IV U7211 ( .A(n6982), .Z(n7175) );
  NOR U7212 ( .A(n111), .B(n43), .Z(n7176) );
  IV U7213 ( .A(n7176), .Z(n6983) );
  NOR U7214 ( .A(n7175), .B(n6983), .Z(n7178) );
  XOR U7215 ( .A(n6985), .B(n6984), .Z(n6986) );
  IV U7216 ( .A(n6986), .Z(n7171) );
  NOR U7217 ( .A(n86), .B(n43), .Z(n7172) );
  IV U7218 ( .A(n7172), .Z(n6987) );
  NOR U7219 ( .A(n7171), .B(n6987), .Z(n7174) );
  IV U7220 ( .A(n6988), .Z(n6990) );
  XOR U7221 ( .A(n6990), .B(n6989), .Z(n7167) );
  NOR U7222 ( .A(n110), .B(n43), .Z(n7168) );
  IV U7223 ( .A(n7168), .Z(n6991) );
  NOR U7224 ( .A(n7167), .B(n6991), .Z(n7170) );
  XOR U7225 ( .A(n6993), .B(n6992), .Z(n6994) );
  IV U7226 ( .A(n6994), .Z(n7163) );
  NOR U7227 ( .A(n109), .B(n43), .Z(n7164) );
  IV U7228 ( .A(n7164), .Z(n6995) );
  NOR U7229 ( .A(n7163), .B(n6995), .Z(n7166) );
  IV U7230 ( .A(n6996), .Z(n6998) );
  XOR U7231 ( .A(n6998), .B(n6997), .Z(n7159) );
  NOR U7232 ( .A(n108), .B(n43), .Z(n7160) );
  IV U7233 ( .A(n7160), .Z(n6999) );
  NOR U7234 ( .A(n7159), .B(n6999), .Z(n7162) );
  XOR U7235 ( .A(n7001), .B(n7000), .Z(n7003) );
  IV U7236 ( .A(n7003), .Z(n7657) );
  NOR U7237 ( .A(n88), .B(n43), .Z(n7002) );
  IV U7238 ( .A(n7002), .Z(n7656) );
  NOR U7239 ( .A(n7657), .B(n7656), .Z(n7142) );
  NOR U7240 ( .A(n7003), .B(n7002), .Z(n7140) );
  XOR U7241 ( .A(n7005), .B(n7004), .Z(n7006) );
  XOR U7242 ( .A(n7007), .B(n7006), .Z(n7137) );
  NOR U7243 ( .A(n106), .B(n43), .Z(n7136) );
  IV U7244 ( .A(n7136), .Z(n7008) );
  NOR U7245 ( .A(n7137), .B(n7008), .Z(n7139) );
  IV U7246 ( .A(n7009), .Z(n7011) );
  XOR U7247 ( .A(n7011), .B(n7010), .Z(n7132) );
  NOR U7248 ( .A(n105), .B(n43), .Z(n7133) );
  IV U7249 ( .A(n7133), .Z(n7012) );
  NOR U7250 ( .A(n7132), .B(n7012), .Z(n7135) );
  NOR U7251 ( .A(n89), .B(n43), .Z(n7120) );
  XOR U7252 ( .A(n7014), .B(n7013), .Z(n7015) );
  NOR U7253 ( .A(n90), .B(n43), .Z(n7016) );
  NOR U7254 ( .A(n7015), .B(n7016), .Z(n7106) );
  IV U7255 ( .A(n7015), .Z(n7623) );
  IV U7256 ( .A(n7016), .Z(n7622) );
  NOR U7257 ( .A(n7623), .B(n7622), .Z(n7104) );
  XOR U7258 ( .A(n7018), .B(n7017), .Z(n7019) );
  XOR U7259 ( .A(n7020), .B(n7019), .Z(n7100) );
  NOR U7260 ( .A(n102), .B(n43), .Z(n7099) );
  IV U7261 ( .A(n7099), .Z(n7021) );
  NOR U7262 ( .A(n7100), .B(n7021), .Z(n7102) );
  XOR U7263 ( .A(n7023), .B(n7022), .Z(n7093) );
  NOR U7264 ( .A(n101), .B(n43), .Z(n7094) );
  NOR U7265 ( .A(n7093), .B(n7094), .Z(n7097) );
  XOR U7266 ( .A(n7025), .B(n7024), .Z(n7026) );
  NOR U7267 ( .A(n99), .B(n43), .Z(n7027) );
  NOR U7268 ( .A(n7026), .B(n7027), .Z(n7082) );
  IV U7269 ( .A(n7026), .Z(n7597) );
  IV U7270 ( .A(n7027), .Z(n7596) );
  NOR U7271 ( .A(n7597), .B(n7596), .Z(n7080) );
  XOR U7272 ( .A(n7029), .B(n7028), .Z(n7066) );
  IV U7273 ( .A(n7066), .Z(n7583) );
  NOR U7274 ( .A(n91), .B(n43), .Z(n7065) );
  IV U7275 ( .A(n7065), .Z(n7582) );
  NOR U7276 ( .A(n7583), .B(n7582), .Z(n7069) );
  IV U7277 ( .A(n7030), .Z(n7032) );
  XOR U7278 ( .A(n7032), .B(n7031), .Z(n7061) );
  NOR U7279 ( .A(n97), .B(n43), .Z(n7062) );
  IV U7280 ( .A(n7062), .Z(n7033) );
  NOR U7281 ( .A(n7061), .B(n7033), .Z(n7064) );
  XOR U7282 ( .A(n7035), .B(n7034), .Z(n7036) );
  IV U7283 ( .A(n7036), .Z(n7057) );
  NOR U7284 ( .A(n96), .B(n43), .Z(n7058) );
  IV U7285 ( .A(n7058), .Z(n7037) );
  NOR U7286 ( .A(n7057), .B(n7037), .Z(n7060) );
  NOR U7287 ( .A(n93), .B(n43), .Z(n7963) );
  IV U7288 ( .A(n7963), .Z(n7038) );
  NOR U7289 ( .A(n118), .B(n168), .Z(n7046) );
  IV U7290 ( .A(n7046), .Z(n7041) );
  NOR U7291 ( .A(n7038), .B(n7041), .Z(n7039) );
  IV U7292 ( .A(n7039), .Z(n7040) );
  NOR U7293 ( .A(n94), .B(n7040), .Z(n7049) );
  NOR U7294 ( .A(n7041), .B(n93), .Z(n7042) );
  XOR U7295 ( .A(n94), .B(n7042), .Z(n7043) );
  NOR U7296 ( .A(n43), .B(n7043), .Z(n7044) );
  IV U7297 ( .A(n7044), .Z(n7562) );
  XOR U7298 ( .A(n7046), .B(n7045), .Z(n7561) );
  IV U7299 ( .A(n7561), .Z(n7047) );
  NOR U7300 ( .A(n7562), .B(n7047), .Z(n7048) );
  NOR U7301 ( .A(n7049), .B(n7048), .Z(n7052) );
  NOR U7302 ( .A(n95), .B(n43), .Z(n7051) );
  IV U7303 ( .A(n7051), .Z(n7050) );
  NOR U7304 ( .A(n7052), .B(n7050), .Z(n7056) );
  XOR U7305 ( .A(n7052), .B(n7051), .Z(n7545) );
  XOR U7306 ( .A(n7054), .B(n7053), .Z(n7546) );
  NOR U7307 ( .A(n7545), .B(n7546), .Z(n7055) );
  NOR U7308 ( .A(n7056), .B(n7055), .Z(n7541) );
  XOR U7309 ( .A(n7058), .B(n7057), .Z(n7542) );
  NOR U7310 ( .A(n7541), .B(n7542), .Z(n7059) );
  NOR U7311 ( .A(n7060), .B(n7059), .Z(n7539) );
  XOR U7312 ( .A(n7062), .B(n7061), .Z(n7538) );
  NOR U7313 ( .A(n7539), .B(n7538), .Z(n7063) );
  NOR U7314 ( .A(n7064), .B(n7063), .Z(n7585) );
  NOR U7315 ( .A(n7066), .B(n7065), .Z(n7067) );
  NOR U7316 ( .A(n7585), .B(n7067), .Z(n7068) );
  NOR U7317 ( .A(n7069), .B(n7068), .Z(n7076) );
  NOR U7318 ( .A(n98), .B(n43), .Z(n7075) );
  IV U7319 ( .A(n7075), .Z(n7070) );
  NOR U7320 ( .A(n7076), .B(n7070), .Z(n7078) );
  XOR U7321 ( .A(n7072), .B(n7071), .Z(n7073) );
  XOR U7322 ( .A(n7074), .B(n7073), .Z(n7536) );
  XOR U7323 ( .A(n7076), .B(n7075), .Z(n7535) );
  NOR U7324 ( .A(n7536), .B(n7535), .Z(n7077) );
  NOR U7325 ( .A(n7078), .B(n7077), .Z(n7599) );
  IV U7326 ( .A(n7599), .Z(n7079) );
  NOR U7327 ( .A(n7080), .B(n7079), .Z(n7081) );
  NOR U7328 ( .A(n7082), .B(n7081), .Z(n7089) );
  IV U7329 ( .A(n7089), .Z(n7084) );
  NOR U7330 ( .A(n100), .B(n43), .Z(n7083) );
  IV U7331 ( .A(n7083), .Z(n7088) );
  NOR U7332 ( .A(n7084), .B(n7088), .Z(n7091) );
  IV U7333 ( .A(n7085), .Z(n7087) );
  XOR U7334 ( .A(n7087), .B(n7086), .Z(n7532) );
  XOR U7335 ( .A(n7089), .B(n7088), .Z(n7531) );
  NOR U7336 ( .A(n7532), .B(n7531), .Z(n7090) );
  NOR U7337 ( .A(n7091), .B(n7090), .Z(n7092) );
  IV U7338 ( .A(n7092), .Z(n7611) );
  XOR U7339 ( .A(n7094), .B(n7093), .Z(n7095) );
  IV U7340 ( .A(n7095), .Z(n7610) );
  NOR U7341 ( .A(n7611), .B(n7610), .Z(n7096) );
  NOR U7342 ( .A(n7097), .B(n7096), .Z(n7098) );
  IV U7343 ( .A(n7098), .Z(n7530) );
  XOR U7344 ( .A(n7100), .B(n7099), .Z(n7529) );
  NOR U7345 ( .A(n7530), .B(n7529), .Z(n7101) );
  NOR U7346 ( .A(n7102), .B(n7101), .Z(n7625) );
  IV U7347 ( .A(n7625), .Z(n7103) );
  NOR U7348 ( .A(n7104), .B(n7103), .Z(n7105) );
  NOR U7349 ( .A(n7106), .B(n7105), .Z(n7112) );
  IV U7350 ( .A(n7112), .Z(n7108) );
  NOR U7351 ( .A(n103), .B(n43), .Z(n7107) );
  IV U7352 ( .A(n7107), .Z(n7111) );
  NOR U7353 ( .A(n7108), .B(n7111), .Z(n7115) );
  XOR U7354 ( .A(n7110), .B(n7109), .Z(n7527) );
  IV U7355 ( .A(n7527), .Z(n7113) );
  XOR U7356 ( .A(n7112), .B(n7111), .Z(n7526) );
  NOR U7357 ( .A(n7113), .B(n7526), .Z(n7114) );
  NOR U7358 ( .A(n7115), .B(n7114), .Z(n7119) );
  IV U7359 ( .A(n7119), .Z(n7116) );
  NOR U7360 ( .A(n7120), .B(n7116), .Z(n7122) );
  XOR U7361 ( .A(n7118), .B(n7117), .Z(n7632) );
  XOR U7362 ( .A(n7120), .B(n7119), .Z(n7631) );
  NOR U7363 ( .A(n7632), .B(n7631), .Z(n7121) );
  NOR U7364 ( .A(n7122), .B(n7121), .Z(n7123) );
  IV U7365 ( .A(n7123), .Z(n7128) );
  NOR U7366 ( .A(n104), .B(n43), .Z(n7127) );
  IV U7367 ( .A(n7127), .Z(n7124) );
  NOR U7368 ( .A(n7128), .B(n7124), .Z(n7131) );
  XOR U7369 ( .A(n7126), .B(n7125), .Z(n7523) );
  IV U7370 ( .A(n7523), .Z(n7129) );
  XOR U7371 ( .A(n7128), .B(n7127), .Z(n7524) );
  NOR U7372 ( .A(n7129), .B(n7524), .Z(n7130) );
  NOR U7373 ( .A(n7131), .B(n7130), .Z(n7643) );
  XOR U7374 ( .A(n7133), .B(n7132), .Z(n7644) );
  NOR U7375 ( .A(n7643), .B(n7644), .Z(n7134) );
  NOR U7376 ( .A(n7135), .B(n7134), .Z(n7519) );
  XOR U7377 ( .A(n7137), .B(n7136), .Z(n7520) );
  NOR U7378 ( .A(n7519), .B(n7520), .Z(n7138) );
  NOR U7379 ( .A(n7139), .B(n7138), .Z(n7659) );
  NOR U7380 ( .A(n7140), .B(n7659), .Z(n7141) );
  NOR U7381 ( .A(n7142), .B(n7141), .Z(n7144) );
  NOR U7382 ( .A(n107), .B(n43), .Z(n7145) );
  IV U7383 ( .A(n7145), .Z(n7143) );
  NOR U7384 ( .A(n7144), .B(n7143), .Z(n7150) );
  XOR U7385 ( .A(n7145), .B(n7144), .Z(n7516) );
  XOR U7386 ( .A(n7147), .B(n7146), .Z(n7148) );
  IV U7387 ( .A(n7148), .Z(n7515) );
  NOR U7388 ( .A(n7516), .B(n7515), .Z(n7149) );
  NOR U7389 ( .A(n7150), .B(n7149), .Z(n7155) );
  NOR U7390 ( .A(n87), .B(n43), .Z(n7154) );
  IV U7391 ( .A(n7154), .Z(n7151) );
  NOR U7392 ( .A(n7155), .B(n7151), .Z(n7158) );
  XOR U7393 ( .A(n7153), .B(n7152), .Z(n7671) );
  IV U7394 ( .A(n7671), .Z(n7156) );
  XOR U7395 ( .A(n7155), .B(n7154), .Z(n7670) );
  NOR U7396 ( .A(n7156), .B(n7670), .Z(n7157) );
  NOR U7397 ( .A(n7158), .B(n7157), .Z(n7511) );
  XOR U7398 ( .A(n7160), .B(n7159), .Z(n7512) );
  NOR U7399 ( .A(n7511), .B(n7512), .Z(n7161) );
  NOR U7400 ( .A(n7162), .B(n7161), .Z(n7680) );
  XOR U7401 ( .A(n7164), .B(n7163), .Z(n7681) );
  NOR U7402 ( .A(n7680), .B(n7681), .Z(n7165) );
  NOR U7403 ( .A(n7166), .B(n7165), .Z(n7509) );
  XOR U7404 ( .A(n7168), .B(n7167), .Z(n7510) );
  NOR U7405 ( .A(n7509), .B(n7510), .Z(n7169) );
  NOR U7406 ( .A(n7170), .B(n7169), .Z(n7693) );
  XOR U7407 ( .A(n7172), .B(n7171), .Z(n7694) );
  NOR U7408 ( .A(n7693), .B(n7694), .Z(n7173) );
  NOR U7409 ( .A(n7174), .B(n7173), .Z(n7506) );
  XOR U7410 ( .A(n7176), .B(n7175), .Z(n7505) );
  NOR U7411 ( .A(n7506), .B(n7505), .Z(n7177) );
  NOR U7412 ( .A(n7178), .B(n7177), .Z(n7179) );
  IV U7413 ( .A(n7179), .Z(n7704) );
  NOR U7414 ( .A(n7705), .B(n7704), .Z(n7180) );
  NOR U7415 ( .A(n7181), .B(n7180), .Z(n7182) );
  IV U7416 ( .A(n7182), .Z(n7712) );
  XOR U7417 ( .A(n7184), .B(n7183), .Z(n7711) );
  NOR U7418 ( .A(n7712), .B(n7711), .Z(n7185) );
  NOR U7419 ( .A(n7186), .B(n7185), .Z(n7717) );
  XOR U7420 ( .A(n7188), .B(n7187), .Z(n7716) );
  NOR U7421 ( .A(n7717), .B(n7716), .Z(n7189) );
  NOR U7422 ( .A(n7190), .B(n7189), .Z(n7499) );
  XOR U7423 ( .A(n7192), .B(n7191), .Z(n7500) );
  NOR U7424 ( .A(n7499), .B(n7500), .Z(n7193) );
  NOR U7425 ( .A(n7194), .B(n7193), .Z(n7495) );
  XOR U7426 ( .A(n7196), .B(n7195), .Z(n7496) );
  NOR U7427 ( .A(n7495), .B(n7496), .Z(n7197) );
  NOR U7428 ( .A(n7198), .B(n7197), .Z(n7734) );
  XOR U7429 ( .A(n7200), .B(n7199), .Z(n7733) );
  NOR U7430 ( .A(n7734), .B(n7733), .Z(n7201) );
  NOR U7431 ( .A(n7202), .B(n7201), .Z(n7491) );
  XOR U7432 ( .A(n7204), .B(n7203), .Z(n7492) );
  NOR U7433 ( .A(n7491), .B(n7492), .Z(n7205) );
  NOR U7434 ( .A(n7206), .B(n7205), .Z(n7487) );
  XOR U7435 ( .A(n7208), .B(n7207), .Z(n7488) );
  NOR U7436 ( .A(n7487), .B(n7488), .Z(n7209) );
  NOR U7437 ( .A(n7210), .B(n7209), .Z(n7483) );
  XOR U7438 ( .A(n7212), .B(n7211), .Z(n7484) );
  NOR U7439 ( .A(n7483), .B(n7484), .Z(n7213) );
  NOR U7440 ( .A(n7214), .B(n7213), .Z(n7479) );
  XOR U7441 ( .A(n7216), .B(n7215), .Z(n7480) );
  NOR U7442 ( .A(n7479), .B(n7480), .Z(n7217) );
  NOR U7443 ( .A(n7218), .B(n7217), .Z(n7476) );
  XOR U7444 ( .A(n7220), .B(n7219), .Z(n7475) );
  NOR U7445 ( .A(n7476), .B(n7475), .Z(n7221) );
  NOR U7446 ( .A(n7222), .B(n7221), .Z(n7472) );
  XOR U7447 ( .A(n7224), .B(n7223), .Z(n7471) );
  NOR U7448 ( .A(n7472), .B(n7471), .Z(n7225) );
  NOR U7449 ( .A(n7226), .B(n7225), .Z(n7766) );
  XOR U7450 ( .A(n7228), .B(n7227), .Z(n7765) );
  NOR U7451 ( .A(n7766), .B(n7765), .Z(n7229) );
  NOR U7452 ( .A(n7230), .B(n7229), .Z(n7468) );
  XOR U7453 ( .A(n7232), .B(n7231), .Z(n7467) );
  NOR U7454 ( .A(n7468), .B(n7467), .Z(n7233) );
  NOR U7455 ( .A(n7234), .B(n7233), .Z(n7464) );
  XOR U7456 ( .A(n7236), .B(n7235), .Z(n7463) );
  NOR U7457 ( .A(n7464), .B(n7463), .Z(n7237) );
  NOR U7458 ( .A(n7238), .B(n7237), .Z(n7782) );
  XOR U7459 ( .A(n7240), .B(n7239), .Z(n7781) );
  NOR U7460 ( .A(n7782), .B(n7781), .Z(n7241) );
  NOR U7461 ( .A(n7242), .B(n7241), .Z(n7788) );
  XOR U7462 ( .A(n7244), .B(n7243), .Z(n7787) );
  NOR U7463 ( .A(n7788), .B(n7787), .Z(n7245) );
  NOR U7464 ( .A(n7246), .B(n7245), .Z(n7460) );
  XOR U7465 ( .A(n7248), .B(n7247), .Z(n7459) );
  NOR U7466 ( .A(n7460), .B(n7459), .Z(n7249) );
  NOR U7467 ( .A(n7250), .B(n7249), .Z(n7800) );
  XOR U7468 ( .A(n7252), .B(n7251), .Z(n7799) );
  NOR U7469 ( .A(n7800), .B(n7799), .Z(n7253) );
  NOR U7470 ( .A(n7254), .B(n7253), .Z(n7808) );
  XOR U7471 ( .A(n7256), .B(n7255), .Z(n7807) );
  NOR U7472 ( .A(n7808), .B(n7807), .Z(n7257) );
  NOR U7473 ( .A(n7258), .B(n7257), .Z(n7816) );
  XOR U7474 ( .A(n7260), .B(n7259), .Z(n7815) );
  NOR U7475 ( .A(n7816), .B(n7815), .Z(n7261) );
  NOR U7476 ( .A(n7262), .B(n7261), .Z(n7824) );
  XOR U7477 ( .A(n7264), .B(n7263), .Z(n7823) );
  NOR U7478 ( .A(n7824), .B(n7823), .Z(n7265) );
  NOR U7479 ( .A(n7266), .B(n7265), .Z(n7832) );
  XOR U7480 ( .A(n7268), .B(n7267), .Z(n7831) );
  NOR U7481 ( .A(n7832), .B(n7831), .Z(n7269) );
  NOR U7482 ( .A(n7270), .B(n7269), .Z(n7840) );
  XOR U7483 ( .A(n7272), .B(n7271), .Z(n7839) );
  NOR U7484 ( .A(n7840), .B(n7839), .Z(n7273) );
  NOR U7485 ( .A(n7274), .B(n7273), .Z(n7456) );
  XOR U7486 ( .A(n7276), .B(n7275), .Z(n7455) );
  NOR U7487 ( .A(n7456), .B(n7455), .Z(n7277) );
  NOR U7488 ( .A(n7278), .B(n7277), .Z(n7852) );
  XOR U7489 ( .A(n7280), .B(n7279), .Z(n7851) );
  NOR U7490 ( .A(n7852), .B(n7851), .Z(n7281) );
  NOR U7491 ( .A(n7282), .B(n7281), .Z(n8300) );
  NOR U7492 ( .A(n143), .B(n118), .Z(n8305) );
  IV U7493 ( .A(n7283), .Z(n7284) );
  NOR U7494 ( .A(n7285), .B(n7284), .Z(n7289) );
  NOR U7495 ( .A(n7287), .B(n7286), .Z(n7288) );
  NOR U7496 ( .A(n7289), .B(n7288), .Z(n8314) );
  NOR U7497 ( .A(n7291), .B(n7290), .Z(n7295) );
  NOR U7498 ( .A(n7293), .B(n7292), .Z(n7294) );
  NOR U7499 ( .A(n7295), .B(n7294), .Z(n8321) );
  NOR U7500 ( .A(n139), .B(n122), .Z(n8319) );
  NOR U7501 ( .A(n137), .B(n124), .Z(n8328) );
  IV U7502 ( .A(n7296), .Z(n7297) );
  NOR U7503 ( .A(n7298), .B(n7297), .Z(n7302) );
  NOR U7504 ( .A(n7300), .B(n7299), .Z(n7301) );
  NOR U7505 ( .A(n7302), .B(n7301), .Z(n8324) );
  NOR U7506 ( .A(n7304), .B(n7303), .Z(n7308) );
  NOR U7507 ( .A(n7306), .B(n7305), .Z(n7307) );
  NOR U7508 ( .A(n7308), .B(n7307), .Z(n8336) );
  NOR U7509 ( .A(n135), .B(n127), .Z(n8333) );
  IV U7510 ( .A(n7309), .Z(n7310) );
  NOR U7511 ( .A(n7311), .B(n7310), .Z(n7315) );
  NOR U7512 ( .A(n7313), .B(n7312), .Z(n7314) );
  NOR U7513 ( .A(n7315), .B(n7314), .Z(n8339) );
  NOR U7514 ( .A(n7317), .B(n7316), .Z(n7321) );
  NOR U7515 ( .A(n7319), .B(n7318), .Z(n7320) );
  NOR U7516 ( .A(n7321), .B(n7320), .Z(n8350) );
  NOR U7517 ( .A(n131), .B(n130), .Z(n8348) );
  IV U7518 ( .A(n8348), .Z(n7444) );
  IV U7519 ( .A(n7322), .Z(n7323) );
  NOR U7520 ( .A(n7324), .B(n7323), .Z(n7328) );
  NOR U7521 ( .A(n7326), .B(n7325), .Z(n7327) );
  NOR U7522 ( .A(n7328), .B(n7327), .Z(n8355) );
  NOR U7523 ( .A(n128), .B(n132), .Z(n8354) );
  NOR U7524 ( .A(n7330), .B(n7329), .Z(n7334) );
  NOR U7525 ( .A(n7332), .B(n7331), .Z(n7333) );
  NOR U7526 ( .A(n7334), .B(n7333), .Z(n8365) );
  NOR U7527 ( .A(n126), .B(n134), .Z(n8362) );
  IV U7528 ( .A(n7335), .Z(n7336) );
  NOR U7529 ( .A(n7337), .B(n7336), .Z(n7341) );
  NOR U7530 ( .A(n7339), .B(n7338), .Z(n7340) );
  NOR U7531 ( .A(n7341), .B(n7340), .Z(n8370) );
  NOR U7532 ( .A(n125), .B(n136), .Z(n8369) );
  NOR U7533 ( .A(n7343), .B(n7342), .Z(n7347) );
  NOR U7534 ( .A(n7345), .B(n7344), .Z(n7346) );
  NOR U7535 ( .A(n7347), .B(n7346), .Z(n8380) );
  NOR U7536 ( .A(n123), .B(n138), .Z(n8377) );
  NOR U7537 ( .A(n7349), .B(n7348), .Z(n7354) );
  IV U7538 ( .A(n7350), .Z(n7352) );
  NOR U7539 ( .A(n7352), .B(n7351), .Z(n7353) );
  NOR U7540 ( .A(n7354), .B(n7353), .Z(n7355) );
  IV U7541 ( .A(n7355), .Z(n8385) );
  NOR U7542 ( .A(n120), .B(n140), .Z(n8383) );
  XOR U7543 ( .A(n8385), .B(n8383), .Z(n8386) );
  NOR U7544 ( .A(n7357), .B(n7356), .Z(n7362) );
  IV U7545 ( .A(n7358), .Z(n7359) );
  NOR U7546 ( .A(n7360), .B(n7359), .Z(n7361) );
  NOR U7547 ( .A(n7362), .B(n7361), .Z(n8393) );
  NOR U7548 ( .A(n119), .B(n142), .Z(n8391) );
  IV U7549 ( .A(n8391), .Z(n7441) );
  NOR U7550 ( .A(n7364), .B(n7363), .Z(n7368) );
  NOR U7551 ( .A(n7366), .B(n7365), .Z(n7367) );
  NOR U7552 ( .A(n7368), .B(n7367), .Z(n8406) );
  NOR U7553 ( .A(n117), .B(n146), .Z(n8404) );
  NOR U7554 ( .A(n7370), .B(n7369), .Z(n7374) );
  NOR U7555 ( .A(n7372), .B(n7371), .Z(n7373) );
  NOR U7556 ( .A(n7374), .B(n7373), .Z(n8419) );
  NOR U7557 ( .A(n116), .B(n151), .Z(n8417) );
  NOR U7558 ( .A(n7376), .B(n7375), .Z(n7380) );
  NOR U7559 ( .A(n7378), .B(n7377), .Z(n7379) );
  NOR U7560 ( .A(n7380), .B(n7379), .Z(n8425) );
  NOR U7561 ( .A(n115), .B(n154), .Z(n8423) );
  IV U7562 ( .A(n7381), .Z(n7382) );
  NOR U7563 ( .A(n7383), .B(n7382), .Z(n7387) );
  NOR U7564 ( .A(n7385), .B(n7384), .Z(n7386) );
  NOR U7565 ( .A(n7387), .B(n7386), .Z(n8432) );
  NOR U7566 ( .A(n7389), .B(n7388), .Z(n7393) );
  NOR U7567 ( .A(n7391), .B(n7390), .Z(n7392) );
  NOR U7568 ( .A(n7393), .B(n7392), .Z(n8438) );
  NOR U7569 ( .A(n114), .B(n159), .Z(n8436) );
  NOR U7570 ( .A(n7395), .B(n7394), .Z(n7399) );
  NOR U7571 ( .A(n7397), .B(n7396), .Z(n7398) );
  NOR U7572 ( .A(n7399), .B(n7398), .Z(n8444) );
  NOR U7573 ( .A(n113), .B(n162), .Z(n8442) );
  IV U7574 ( .A(n8442), .Z(n7408) );
  IV U7575 ( .A(n7400), .Z(n7401) );
  NOR U7576 ( .A(n7402), .B(n7401), .Z(n7406) );
  NOR U7577 ( .A(n7404), .B(n7403), .Z(n7405) );
  NOR U7578 ( .A(n7406), .B(n7405), .Z(n8449) );
  NOR U7579 ( .A(n164), .B(n84), .Z(n8447) );
  XOR U7580 ( .A(n8449), .B(n8447), .Z(n8451) );
  NOR U7581 ( .A(n166), .B(n112), .Z(n7407) );
  IV U7582 ( .A(n7407), .Z(n8450) );
  XOR U7583 ( .A(n8451), .B(n8450), .Z(n8441) );
  XOR U7584 ( .A(n7408), .B(n8441), .Z(n8443) );
  XOR U7585 ( .A(n8444), .B(n8443), .Z(n8460) );
  IV U7586 ( .A(n7409), .Z(n7410) );
  NOR U7587 ( .A(n7411), .B(n7410), .Z(n7415) );
  NOR U7588 ( .A(n7413), .B(n7412), .Z(n7414) );
  NOR U7589 ( .A(n7415), .B(n7414), .Z(n8458) );
  NOR U7590 ( .A(n83), .B(n160), .Z(n8456) );
  XOR U7591 ( .A(n8458), .B(n8456), .Z(n8459) );
  XOR U7592 ( .A(n8460), .B(n8459), .Z(n8435) );
  XOR U7593 ( .A(n8436), .B(n8435), .Z(n7416) );
  IV U7594 ( .A(n7416), .Z(n8437) );
  XOR U7595 ( .A(n8438), .B(n8437), .Z(n8430) );
  NOR U7596 ( .A(n82), .B(n157), .Z(n8428) );
  XOR U7597 ( .A(n8430), .B(n8428), .Z(n8431) );
  XOR U7598 ( .A(n8432), .B(n8431), .Z(n8422) );
  XOR U7599 ( .A(n8423), .B(n8422), .Z(n7417) );
  IV U7600 ( .A(n7417), .Z(n8424) );
  XOR U7601 ( .A(n8425), .B(n8424), .Z(n8469) );
  IV U7602 ( .A(n7418), .Z(n7419) );
  NOR U7603 ( .A(n7420), .B(n7419), .Z(n7424) );
  NOR U7604 ( .A(n7422), .B(n7421), .Z(n7423) );
  NOR U7605 ( .A(n7424), .B(n7423), .Z(n8467) );
  NOR U7606 ( .A(n81), .B(n152), .Z(n8465) );
  XOR U7607 ( .A(n8467), .B(n8465), .Z(n8468) );
  XOR U7608 ( .A(n8469), .B(n8468), .Z(n8416) );
  XOR U7609 ( .A(n8417), .B(n8416), .Z(n7425) );
  IV U7610 ( .A(n7425), .Z(n8418) );
  XOR U7611 ( .A(n8419), .B(n8418), .Z(n8413) );
  IV U7612 ( .A(n7426), .Z(n7427) );
  NOR U7613 ( .A(n7428), .B(n7427), .Z(n7432) );
  NOR U7614 ( .A(n7430), .B(n7429), .Z(n7431) );
  NOR U7615 ( .A(n7432), .B(n7431), .Z(n8411) );
  NOR U7616 ( .A(n80), .B(n149), .Z(n8409) );
  XOR U7617 ( .A(n8411), .B(n8409), .Z(n8412) );
  XOR U7618 ( .A(n8413), .B(n8412), .Z(n8403) );
  XOR U7619 ( .A(n8404), .B(n8403), .Z(n7433) );
  IV U7620 ( .A(n7433), .Z(n8405) );
  XOR U7621 ( .A(n8406), .B(n8405), .Z(n8400) );
  IV U7622 ( .A(n7434), .Z(n7435) );
  NOR U7623 ( .A(n7436), .B(n7435), .Z(n7440) );
  NOR U7624 ( .A(n7438), .B(n7437), .Z(n7439) );
  NOR U7625 ( .A(n7440), .B(n7439), .Z(n8398) );
  NOR U7626 ( .A(n79), .B(n144), .Z(n8396) );
  XOR U7627 ( .A(n8398), .B(n8396), .Z(n8399) );
  XOR U7628 ( .A(n8400), .B(n8399), .Z(n8390) );
  XOR U7629 ( .A(n7441), .B(n8390), .Z(n8392) );
  XOR U7630 ( .A(n8393), .B(n8392), .Z(n8387) );
  XOR U7631 ( .A(n8386), .B(n8387), .Z(n8376) );
  XOR U7632 ( .A(n8377), .B(n8376), .Z(n8378) );
  XOR U7633 ( .A(n8380), .B(n8378), .Z(n8368) );
  XOR U7634 ( .A(n8369), .B(n8368), .Z(n7442) );
  IV U7635 ( .A(n7442), .Z(n8371) );
  XOR U7636 ( .A(n8370), .B(n8371), .Z(n8361) );
  XOR U7637 ( .A(n8362), .B(n8361), .Z(n8363) );
  XOR U7638 ( .A(n8365), .B(n8363), .Z(n8353) );
  XOR U7639 ( .A(n8354), .B(n8353), .Z(n7443) );
  IV U7640 ( .A(n7443), .Z(n8357) );
  XOR U7641 ( .A(n8355), .B(n8357), .Z(n8347) );
  XOR U7642 ( .A(n7444), .B(n8347), .Z(n8349) );
  XOR U7643 ( .A(n8350), .B(n8349), .Z(n8340) );
  XOR U7644 ( .A(n8339), .B(n8340), .Z(n8341) );
  NOR U7645 ( .A(n133), .B(n129), .Z(n8342) );
  XOR U7646 ( .A(n8341), .B(n8342), .Z(n8332) );
  XOR U7647 ( .A(n8333), .B(n8332), .Z(n8334) );
  XOR U7648 ( .A(n8336), .B(n8334), .Z(n8325) );
  XOR U7649 ( .A(n8324), .B(n8325), .Z(n8327) );
  XOR U7650 ( .A(n8328), .B(n8327), .Z(n8317) );
  XOR U7651 ( .A(n8319), .B(n8317), .Z(n8320) );
  XOR U7652 ( .A(n8321), .B(n8320), .Z(n8312) );
  NOR U7653 ( .A(n141), .B(n121), .Z(n8310) );
  XOR U7654 ( .A(n8312), .B(n8310), .Z(n8313) );
  XOR U7655 ( .A(n8314), .B(n8313), .Z(n8304) );
  XOR U7656 ( .A(n8305), .B(n8304), .Z(n7445) );
  IV U7657 ( .A(n7445), .Z(n8307) );
  IV U7658 ( .A(n7446), .Z(n7447) );
  NOR U7659 ( .A(n7448), .B(n7447), .Z(n7453) );
  IV U7660 ( .A(n7449), .Z(n7450) );
  NOR U7661 ( .A(n7451), .B(n7450), .Z(n7452) );
  NOR U7662 ( .A(n7453), .B(n7452), .Z(n7454) );
  IV U7663 ( .A(n7454), .Z(n8306) );
  XOR U7664 ( .A(n8307), .B(n8306), .Z(n8298) );
  NOR U7665 ( .A(n145), .B(n43), .Z(n8296) );
  XOR U7666 ( .A(n8298), .B(n8296), .Z(n8299) );
  XOR U7667 ( .A(n8300), .B(n8299), .Z(n8291) );
  XOR U7668 ( .A(n7456), .B(n7455), .Z(n7846) );
  IV U7669 ( .A(n7846), .Z(n7458) );
  NOR U7670 ( .A(n143), .B(n42), .Z(n7457) );
  IV U7671 ( .A(n7457), .Z(n7847) );
  NOR U7672 ( .A(n7458), .B(n7847), .Z(n7849) );
  XOR U7673 ( .A(n7460), .B(n7459), .Z(n7794) );
  IV U7674 ( .A(n7794), .Z(n7462) );
  NOR U7675 ( .A(n128), .B(n42), .Z(n7461) );
  IV U7676 ( .A(n7461), .Z(n7795) );
  NOR U7677 ( .A(n7462), .B(n7795), .Z(n7797) );
  XOR U7678 ( .A(n7464), .B(n7463), .Z(n7774) );
  IV U7679 ( .A(n7774), .Z(n7466) );
  NOR U7680 ( .A(n123), .B(n42), .Z(n7465) );
  IV U7681 ( .A(n7465), .Z(n7775) );
  NOR U7682 ( .A(n7466), .B(n7775), .Z(n7777) );
  XOR U7683 ( .A(n7468), .B(n7467), .Z(n7770) );
  IV U7684 ( .A(n7770), .Z(n7470) );
  NOR U7685 ( .A(n120), .B(n42), .Z(n7469) );
  IV U7686 ( .A(n7469), .Z(n7771) );
  NOR U7687 ( .A(n7470), .B(n7771), .Z(n7773) );
  XOR U7688 ( .A(n7472), .B(n7471), .Z(n7758) );
  IV U7689 ( .A(n7758), .Z(n7474) );
  NOR U7690 ( .A(n79), .B(n42), .Z(n7473) );
  IV U7691 ( .A(n7473), .Z(n7759) );
  NOR U7692 ( .A(n7474), .B(n7759), .Z(n7761) );
  XOR U7693 ( .A(n7476), .B(n7475), .Z(n7754) );
  IV U7694 ( .A(n7754), .Z(n7478) );
  NOR U7695 ( .A(n117), .B(n42), .Z(n7477) );
  IV U7696 ( .A(n7477), .Z(n7755) );
  NOR U7697 ( .A(n7478), .B(n7755), .Z(n7757) );
  IV U7698 ( .A(n7479), .Z(n7481) );
  XOR U7699 ( .A(n7481), .B(n7480), .Z(n7750) );
  NOR U7700 ( .A(n80), .B(n42), .Z(n7751) );
  IV U7701 ( .A(n7751), .Z(n7482) );
  NOR U7702 ( .A(n7750), .B(n7482), .Z(n7753) );
  IV U7703 ( .A(n7483), .Z(n7485) );
  XOR U7704 ( .A(n7485), .B(n7484), .Z(n7746) );
  NOR U7705 ( .A(n116), .B(n42), .Z(n7747) );
  IV U7706 ( .A(n7747), .Z(n7486) );
  NOR U7707 ( .A(n7746), .B(n7486), .Z(n7749) );
  IV U7708 ( .A(n7487), .Z(n7489) );
  XOR U7709 ( .A(n7489), .B(n7488), .Z(n7742) );
  NOR U7710 ( .A(n81), .B(n42), .Z(n7743) );
  IV U7711 ( .A(n7743), .Z(n7490) );
  NOR U7712 ( .A(n7742), .B(n7490), .Z(n7745) );
  IV U7713 ( .A(n7491), .Z(n7493) );
  XOR U7714 ( .A(n7493), .B(n7492), .Z(n7738) );
  NOR U7715 ( .A(n115), .B(n42), .Z(n7739) );
  IV U7716 ( .A(n7739), .Z(n7494) );
  NOR U7717 ( .A(n7738), .B(n7494), .Z(n7741) );
  IV U7718 ( .A(n7495), .Z(n7497) );
  XOR U7719 ( .A(n7497), .B(n7496), .Z(n7726) );
  NOR U7720 ( .A(n114), .B(n42), .Z(n7727) );
  IV U7721 ( .A(n7727), .Z(n7498) );
  NOR U7722 ( .A(n7726), .B(n7498), .Z(n7729) );
  IV U7723 ( .A(n7499), .Z(n7501) );
  XOR U7724 ( .A(n7501), .B(n7500), .Z(n7503) );
  NOR U7725 ( .A(n83), .B(n42), .Z(n7504) );
  IV U7726 ( .A(n7504), .Z(n7502) );
  NOR U7727 ( .A(n7503), .B(n7502), .Z(n7725) );
  XOR U7728 ( .A(n7504), .B(n7503), .Z(n8127) );
  NOR U7729 ( .A(n113), .B(n42), .Z(n7719) );
  NOR U7730 ( .A(n84), .B(n42), .Z(n7709) );
  XOR U7731 ( .A(n7506), .B(n7505), .Z(n7507) );
  NOR U7732 ( .A(n85), .B(n42), .Z(n7508) );
  NOR U7733 ( .A(n7507), .B(n7508), .Z(n7701) );
  IV U7734 ( .A(n7507), .Z(n8100) );
  IV U7735 ( .A(n7508), .Z(n8099) );
  NOR U7736 ( .A(n8100), .B(n8099), .Z(n7699) );
  XOR U7737 ( .A(n7510), .B(n7509), .Z(n7686) );
  IV U7738 ( .A(n7686), .Z(n8086) );
  NOR U7739 ( .A(n86), .B(n42), .Z(n7685) );
  IV U7740 ( .A(n7685), .Z(n8085) );
  NOR U7741 ( .A(n8086), .B(n8085), .Z(n7689) );
  XOR U7742 ( .A(n7512), .B(n7511), .Z(n7514) );
  IV U7743 ( .A(n7514), .Z(n8075) );
  NOR U7744 ( .A(n109), .B(n42), .Z(n7513) );
  IV U7745 ( .A(n7513), .Z(n8074) );
  NOR U7746 ( .A(n8075), .B(n8074), .Z(n7676) );
  NOR U7747 ( .A(n7514), .B(n7513), .Z(n7674) );
  XOR U7748 ( .A(n7516), .B(n7515), .Z(n7517) );
  NOR U7749 ( .A(n87), .B(n42), .Z(n7518) );
  NOR U7750 ( .A(n7517), .B(n7518), .Z(n7665) );
  IV U7751 ( .A(n7517), .Z(n7900) );
  IV U7752 ( .A(n7518), .Z(n7899) );
  NOR U7753 ( .A(n7900), .B(n7899), .Z(n7663) );
  NOR U7754 ( .A(n88), .B(n42), .Z(n7522) );
  IV U7755 ( .A(n7522), .Z(n8052) );
  XOR U7756 ( .A(n7520), .B(n7519), .Z(n7521) );
  IV U7757 ( .A(n7521), .Z(n8051) );
  NOR U7758 ( .A(n8052), .B(n8051), .Z(n7652) );
  NOR U7759 ( .A(n7522), .B(n7521), .Z(n7650) );
  XOR U7760 ( .A(n7524), .B(n7523), .Z(n7637) );
  NOR U7761 ( .A(n105), .B(n42), .Z(n7525) );
  IV U7762 ( .A(n7525), .Z(n7638) );
  NOR U7763 ( .A(n7637), .B(n7638), .Z(n7641) );
  XOR U7764 ( .A(n7527), .B(n7526), .Z(n7916) );
  NOR U7765 ( .A(n89), .B(n42), .Z(n7528) );
  IV U7766 ( .A(n7528), .Z(n7915) );
  XOR U7767 ( .A(n7530), .B(n7529), .Z(n7617) );
  IV U7768 ( .A(n7617), .Z(n8017) );
  NOR U7769 ( .A(n90), .B(n42), .Z(n7616) );
  IV U7770 ( .A(n7616), .Z(n8016) );
  NOR U7771 ( .A(n8017), .B(n8016), .Z(n7620) );
  NOR U7772 ( .A(n102), .B(n42), .Z(n7613) );
  IV U7773 ( .A(n7613), .Z(n7609) );
  NOR U7774 ( .A(n101), .B(n42), .Z(n7533) );
  XOR U7775 ( .A(n7532), .B(n7531), .Z(n7534) );
  NOR U7776 ( .A(n7533), .B(n7534), .Z(n7607) );
  IV U7777 ( .A(n7533), .Z(n7925) );
  IV U7778 ( .A(n7534), .Z(n7924) );
  NOR U7779 ( .A(n7925), .B(n7924), .Z(n7605) );
  XOR U7780 ( .A(n7536), .B(n7535), .Z(n7591) );
  IV U7781 ( .A(n7591), .Z(n7934) );
  NOR U7782 ( .A(n99), .B(n42), .Z(n7590) );
  IV U7783 ( .A(n7590), .Z(n7933) );
  NOR U7784 ( .A(n7934), .B(n7933), .Z(n7594) );
  NOR U7785 ( .A(n91), .B(n42), .Z(n7537) );
  IV U7786 ( .A(n7537), .Z(n7578) );
  XOR U7787 ( .A(n7539), .B(n7538), .Z(n7577) );
  IV U7788 ( .A(n7577), .Z(n7540) );
  NOR U7789 ( .A(n7578), .B(n7540), .Z(n7580) );
  XOR U7790 ( .A(n7542), .B(n7541), .Z(n7543) );
  IV U7791 ( .A(n7543), .Z(n7573) );
  NOR U7792 ( .A(n97), .B(n42), .Z(n7574) );
  IV U7793 ( .A(n7574), .Z(n7544) );
  NOR U7794 ( .A(n7573), .B(n7544), .Z(n7576) );
  XOR U7795 ( .A(n7546), .B(n7545), .Z(n7547) );
  IV U7796 ( .A(n7547), .Z(n7569) );
  NOR U7797 ( .A(n96), .B(n42), .Z(n7570) );
  IV U7798 ( .A(n7570), .Z(n7548) );
  NOR U7799 ( .A(n7569), .B(n7548), .Z(n7572) );
  NOR U7800 ( .A(n93), .B(n42), .Z(n10507) );
  IV U7801 ( .A(n10507), .Z(n7549) );
  NOR U7802 ( .A(n43), .B(n168), .Z(n7557) );
  IV U7803 ( .A(n7557), .Z(n7552) );
  NOR U7804 ( .A(n7549), .B(n7552), .Z(n7550) );
  IV U7805 ( .A(n7550), .Z(n7551) );
  NOR U7806 ( .A(n94), .B(n7551), .Z(n7560) );
  NOR U7807 ( .A(n7552), .B(n93), .Z(n7553) );
  XOR U7808 ( .A(n94), .B(n7553), .Z(n7554) );
  NOR U7809 ( .A(n42), .B(n7554), .Z(n7555) );
  IV U7810 ( .A(n7555), .Z(n7954) );
  XOR U7811 ( .A(n7557), .B(n7556), .Z(n7953) );
  IV U7812 ( .A(n7953), .Z(n7558) );
  NOR U7813 ( .A(n7954), .B(n7558), .Z(n7559) );
  NOR U7814 ( .A(n7560), .B(n7559), .Z(n7563) );
  XOR U7815 ( .A(n7562), .B(n7561), .Z(n7564) );
  NOR U7816 ( .A(n7563), .B(n7564), .Z(n7568) );
  IV U7817 ( .A(n7563), .Z(n7565) );
  XOR U7818 ( .A(n7565), .B(n7564), .Z(n7950) );
  NOR U7819 ( .A(n95), .B(n42), .Z(n7951) );
  IV U7820 ( .A(n7951), .Z(n7566) );
  NOR U7821 ( .A(n7950), .B(n7566), .Z(n7567) );
  NOR U7822 ( .A(n7568), .B(n7567), .Z(n7946) );
  XOR U7823 ( .A(n7570), .B(n7569), .Z(n7947) );
  NOR U7824 ( .A(n7946), .B(n7947), .Z(n7571) );
  NOR U7825 ( .A(n7572), .B(n7571), .Z(n7943) );
  XOR U7826 ( .A(n7574), .B(n7573), .Z(n7942) );
  NOR U7827 ( .A(n7943), .B(n7942), .Z(n7575) );
  NOR U7828 ( .A(n7576), .B(n7575), .Z(n7987) );
  XOR U7829 ( .A(n7578), .B(n7577), .Z(n7986) );
  NOR U7830 ( .A(n7987), .B(n7986), .Z(n7579) );
  NOR U7831 ( .A(n7580), .B(n7579), .Z(n7587) );
  NOR U7832 ( .A(n98), .B(n42), .Z(n7586) );
  IV U7833 ( .A(n7586), .Z(n7581) );
  NOR U7834 ( .A(n7587), .B(n7581), .Z(n7589) );
  XOR U7835 ( .A(n7583), .B(n7582), .Z(n7584) );
  XOR U7836 ( .A(n7585), .B(n7584), .Z(n7940) );
  XOR U7837 ( .A(n7587), .B(n7586), .Z(n7939) );
  NOR U7838 ( .A(n7940), .B(n7939), .Z(n7588) );
  NOR U7839 ( .A(n7589), .B(n7588), .Z(n7936) );
  NOR U7840 ( .A(n7591), .B(n7590), .Z(n7592) );
  NOR U7841 ( .A(n7936), .B(n7592), .Z(n7593) );
  NOR U7842 ( .A(n7594), .B(n7593), .Z(n7601) );
  NOR U7843 ( .A(n100), .B(n42), .Z(n7600) );
  IV U7844 ( .A(n7600), .Z(n7595) );
  NOR U7845 ( .A(n7601), .B(n7595), .Z(n7603) );
  XOR U7846 ( .A(n7597), .B(n7596), .Z(n7598) );
  XOR U7847 ( .A(n7599), .B(n7598), .Z(n7930) );
  XOR U7848 ( .A(n7601), .B(n7600), .Z(n7929) );
  NOR U7849 ( .A(n7930), .B(n7929), .Z(n7602) );
  NOR U7850 ( .A(n7603), .B(n7602), .Z(n7927) );
  IV U7851 ( .A(n7927), .Z(n7604) );
  NOR U7852 ( .A(n7605), .B(n7604), .Z(n7606) );
  NOR U7853 ( .A(n7607), .B(n7606), .Z(n7608) );
  IV U7854 ( .A(n7608), .Z(n7612) );
  NOR U7855 ( .A(n7609), .B(n7612), .Z(n7615) );
  XOR U7856 ( .A(n7611), .B(n7610), .Z(n7922) );
  XOR U7857 ( .A(n7613), .B(n7612), .Z(n7923) );
  NOR U7858 ( .A(n7922), .B(n7923), .Z(n7614) );
  NOR U7859 ( .A(n7615), .B(n7614), .Z(n8019) );
  NOR U7860 ( .A(n7617), .B(n7616), .Z(n7618) );
  NOR U7861 ( .A(n8019), .B(n7618), .Z(n7619) );
  NOR U7862 ( .A(n7620), .B(n7619), .Z(n7627) );
  NOR U7863 ( .A(n103), .B(n42), .Z(n7626) );
  IV U7864 ( .A(n7626), .Z(n7621) );
  NOR U7865 ( .A(n7627), .B(n7621), .Z(n7629) );
  XOR U7866 ( .A(n7623), .B(n7622), .Z(n7624) );
  XOR U7867 ( .A(n7625), .B(n7624), .Z(n7921) );
  XOR U7868 ( .A(n7627), .B(n7626), .Z(n7920) );
  NOR U7869 ( .A(n7921), .B(n7920), .Z(n7628) );
  NOR U7870 ( .A(n7629), .B(n7628), .Z(n7918) );
  NOR U7871 ( .A(n104), .B(n42), .Z(n7633) );
  IV U7872 ( .A(n7633), .Z(n7630) );
  NOR U7873 ( .A(n7634), .B(n7630), .Z(n7636) );
  XOR U7874 ( .A(n7632), .B(n7631), .Z(n7911) );
  XOR U7875 ( .A(n7634), .B(n7633), .Z(n7912) );
  NOR U7876 ( .A(n7911), .B(n7912), .Z(n7635) );
  NOR U7877 ( .A(n7636), .B(n7635), .Z(n8040) );
  XOR U7878 ( .A(n7638), .B(n7637), .Z(n8041) );
  IV U7879 ( .A(n8041), .Z(n7639) );
  NOR U7880 ( .A(n8040), .B(n7639), .Z(n7640) );
  NOR U7881 ( .A(n7641), .B(n7640), .Z(n7646) );
  NOR U7882 ( .A(n106), .B(n42), .Z(n7645) );
  IV U7883 ( .A(n7645), .Z(n7642) );
  NOR U7884 ( .A(n7646), .B(n7642), .Z(n7649) );
  XOR U7885 ( .A(n7644), .B(n7643), .Z(n7909) );
  IV U7886 ( .A(n7909), .Z(n7647) );
  XOR U7887 ( .A(n7646), .B(n7645), .Z(n7908) );
  NOR U7888 ( .A(n7647), .B(n7908), .Z(n7648) );
  NOR U7889 ( .A(n7649), .B(n7648), .Z(n8054) );
  NOR U7890 ( .A(n7650), .B(n8054), .Z(n7651) );
  NOR U7891 ( .A(n7652), .B(n7651), .Z(n7655) );
  NOR U7892 ( .A(n107), .B(n42), .Z(n7654) );
  IV U7893 ( .A(n7654), .Z(n7653) );
  NOR U7894 ( .A(n7655), .B(n7653), .Z(n7661) );
  XOR U7895 ( .A(n7655), .B(n7654), .Z(n7905) );
  XOR U7896 ( .A(n7657), .B(n7656), .Z(n7658) );
  XOR U7897 ( .A(n7659), .B(n7658), .Z(n7906) );
  NOR U7898 ( .A(n7905), .B(n7906), .Z(n7660) );
  NOR U7899 ( .A(n7661), .B(n7660), .Z(n7902) );
  IV U7900 ( .A(n7902), .Z(n7662) );
  NOR U7901 ( .A(n7663), .B(n7662), .Z(n7664) );
  NOR U7902 ( .A(n7665), .B(n7664), .Z(n7666) );
  IV U7903 ( .A(n7666), .Z(n7669) );
  NOR U7904 ( .A(n108), .B(n42), .Z(n7668) );
  IV U7905 ( .A(n7668), .Z(n7667) );
  NOR U7906 ( .A(n7669), .B(n7667), .Z(n7673) );
  XOR U7907 ( .A(n7669), .B(n7668), .Z(n7896) );
  XOR U7908 ( .A(n7671), .B(n7670), .Z(n7895) );
  NOR U7909 ( .A(n7896), .B(n7895), .Z(n7672) );
  NOR U7910 ( .A(n7673), .B(n7672), .Z(n8077) );
  NOR U7911 ( .A(n7674), .B(n8077), .Z(n7675) );
  NOR U7912 ( .A(n7676), .B(n7675), .Z(n7679) );
  NOR U7913 ( .A(n110), .B(n42), .Z(n7678) );
  IV U7914 ( .A(n7678), .Z(n7677) );
  NOR U7915 ( .A(n7679), .B(n7677), .Z(n7684) );
  XOR U7916 ( .A(n7679), .B(n7678), .Z(n7892) );
  XOR U7917 ( .A(n7681), .B(n7680), .Z(n7682) );
  IV U7918 ( .A(n7682), .Z(n7891) );
  NOR U7919 ( .A(n7892), .B(n7891), .Z(n7683) );
  NOR U7920 ( .A(n7684), .B(n7683), .Z(n8088) );
  NOR U7921 ( .A(n7686), .B(n7685), .Z(n7687) );
  NOR U7922 ( .A(n8088), .B(n7687), .Z(n7688) );
  NOR U7923 ( .A(n7689), .B(n7688), .Z(n7692) );
  NOR U7924 ( .A(n111), .B(n42), .Z(n7691) );
  IV U7925 ( .A(n7691), .Z(n7690) );
  NOR U7926 ( .A(n7692), .B(n7690), .Z(n7697) );
  XOR U7927 ( .A(n7692), .B(n7691), .Z(n7887) );
  XOR U7928 ( .A(n7694), .B(n7693), .Z(n7695) );
  IV U7929 ( .A(n7695), .Z(n7886) );
  NOR U7930 ( .A(n7887), .B(n7886), .Z(n7696) );
  NOR U7931 ( .A(n7697), .B(n7696), .Z(n8102) );
  IV U7932 ( .A(n8102), .Z(n7698) );
  NOR U7933 ( .A(n7699), .B(n7698), .Z(n7700) );
  NOR U7934 ( .A(n7701), .B(n7700), .Z(n7703) );
  IV U7935 ( .A(n7703), .Z(n7882) );
  NOR U7936 ( .A(n112), .B(n42), .Z(n7702) );
  IV U7937 ( .A(n7702), .Z(n7881) );
  NOR U7938 ( .A(n7882), .B(n7881), .Z(n7708) );
  NOR U7939 ( .A(n7703), .B(n7702), .Z(n7706) );
  XOR U7940 ( .A(n7705), .B(n7704), .Z(n7884) );
  NOR U7941 ( .A(n7706), .B(n7884), .Z(n7707) );
  NOR U7942 ( .A(n7708), .B(n7707), .Z(n7710) );
  IV U7943 ( .A(n7710), .Z(n8111) );
  NOR U7944 ( .A(n7709), .B(n8111), .Z(n7715) );
  IV U7945 ( .A(n7709), .Z(n8112) );
  NOR U7946 ( .A(n7710), .B(n8112), .Z(n7713) );
  XOR U7947 ( .A(n7712), .B(n7711), .Z(n8114) );
  NOR U7948 ( .A(n7713), .B(n8114), .Z(n7714) );
  NOR U7949 ( .A(n7715), .B(n7714), .Z(n7718) );
  NOR U7950 ( .A(n7719), .B(n7718), .Z(n7722) );
  XOR U7951 ( .A(n7717), .B(n7716), .Z(n7877) );
  XOR U7952 ( .A(n7719), .B(n7718), .Z(n7878) );
  IV U7953 ( .A(n7878), .Z(n7720) );
  NOR U7954 ( .A(n7877), .B(n7720), .Z(n7721) );
  NOR U7955 ( .A(n7722), .B(n7721), .Z(n7723) );
  IV U7956 ( .A(n7723), .Z(n8126) );
  NOR U7957 ( .A(n8127), .B(n8126), .Z(n7724) );
  NOR U7958 ( .A(n7725), .B(n7724), .Z(n8134) );
  XOR U7959 ( .A(n7727), .B(n7726), .Z(n8133) );
  NOR U7960 ( .A(n8134), .B(n8133), .Z(n7728) );
  NOR U7961 ( .A(n7729), .B(n7728), .Z(n7732) );
  NOR U7962 ( .A(n82), .B(n42), .Z(n7731) );
  IV U7963 ( .A(n7731), .Z(n7730) );
  NOR U7964 ( .A(n7732), .B(n7730), .Z(n7737) );
  XOR U7965 ( .A(n7732), .B(n7731), .Z(n8140) );
  XOR U7966 ( .A(n7734), .B(n7733), .Z(n8141) );
  IV U7967 ( .A(n8141), .Z(n7735) );
  NOR U7968 ( .A(n8140), .B(n7735), .Z(n7736) );
  NOR U7969 ( .A(n7737), .B(n7736), .Z(n8151) );
  XOR U7970 ( .A(n7739), .B(n7738), .Z(n8150) );
  NOR U7971 ( .A(n8151), .B(n8150), .Z(n7740) );
  NOR U7972 ( .A(n7741), .B(n7740), .Z(n8156) );
  XOR U7973 ( .A(n7743), .B(n7742), .Z(n8155) );
  NOR U7974 ( .A(n8156), .B(n8155), .Z(n7744) );
  NOR U7975 ( .A(n7745), .B(n7744), .Z(n8163) );
  XOR U7976 ( .A(n7747), .B(n7746), .Z(n8162) );
  NOR U7977 ( .A(n8163), .B(n8162), .Z(n7748) );
  NOR U7978 ( .A(n7749), .B(n7748), .Z(n8174) );
  XOR U7979 ( .A(n7751), .B(n7750), .Z(n8173) );
  NOR U7980 ( .A(n8174), .B(n8173), .Z(n7752) );
  NOR U7981 ( .A(n7753), .B(n7752), .Z(n8182) );
  XOR U7982 ( .A(n7755), .B(n7754), .Z(n8181) );
  NOR U7983 ( .A(n8182), .B(n8181), .Z(n7756) );
  NOR U7984 ( .A(n7757), .B(n7756), .Z(n8189) );
  XOR U7985 ( .A(n7759), .B(n7758), .Z(n8190) );
  NOR U7986 ( .A(n8189), .B(n8190), .Z(n7760) );
  NOR U7987 ( .A(n7761), .B(n7760), .Z(n7764) );
  NOR U7988 ( .A(n119), .B(n42), .Z(n7763) );
  IV U7989 ( .A(n7763), .Z(n7762) );
  NOR U7990 ( .A(n7764), .B(n7762), .Z(n7769) );
  XOR U7991 ( .A(n7764), .B(n7763), .Z(n8197) );
  XOR U7992 ( .A(n7766), .B(n7765), .Z(n8198) );
  IV U7993 ( .A(n8198), .Z(n7767) );
  NOR U7994 ( .A(n8197), .B(n7767), .Z(n7768) );
  NOR U7995 ( .A(n7769), .B(n7768), .Z(n8205) );
  XOR U7996 ( .A(n7771), .B(n7770), .Z(n8204) );
  NOR U7997 ( .A(n8205), .B(n8204), .Z(n7772) );
  NOR U7998 ( .A(n7773), .B(n7772), .Z(n8213) );
  XOR U7999 ( .A(n7775), .B(n7774), .Z(n8212) );
  NOR U8000 ( .A(n8213), .B(n8212), .Z(n7776) );
  NOR U8001 ( .A(n7777), .B(n7776), .Z(n7780) );
  NOR U8002 ( .A(n125), .B(n42), .Z(n7779) );
  IV U8003 ( .A(n7779), .Z(n7778) );
  NOR U8004 ( .A(n7780), .B(n7778), .Z(n7785) );
  XOR U8005 ( .A(n7780), .B(n7779), .Z(n8217) );
  XOR U8006 ( .A(n7782), .B(n7781), .Z(n8218) );
  IV U8007 ( .A(n8218), .Z(n7783) );
  NOR U8008 ( .A(n8217), .B(n7783), .Z(n7784) );
  NOR U8009 ( .A(n7785), .B(n7784), .Z(n7790) );
  NOR U8010 ( .A(n126), .B(n42), .Z(n7789) );
  IV U8011 ( .A(n7789), .Z(n7786) );
  NOR U8012 ( .A(n7790), .B(n7786), .Z(n7793) );
  XOR U8013 ( .A(n7788), .B(n7787), .Z(n7875) );
  IV U8014 ( .A(n7875), .Z(n7791) );
  XOR U8015 ( .A(n7790), .B(n7789), .Z(n7874) );
  NOR U8016 ( .A(n7791), .B(n7874), .Z(n7792) );
  NOR U8017 ( .A(n7793), .B(n7792), .Z(n8233) );
  XOR U8018 ( .A(n7795), .B(n7794), .Z(n8232) );
  NOR U8019 ( .A(n8233), .B(n8232), .Z(n7796) );
  NOR U8020 ( .A(n7797), .B(n7796), .Z(n7802) );
  NOR U8021 ( .A(n131), .B(n42), .Z(n7801) );
  IV U8022 ( .A(n7801), .Z(n7798) );
  NOR U8023 ( .A(n7802), .B(n7798), .Z(n7805) );
  XOR U8024 ( .A(n7800), .B(n7799), .Z(n8238) );
  IV U8025 ( .A(n8238), .Z(n7803) );
  XOR U8026 ( .A(n7802), .B(n7801), .Z(n8237) );
  NOR U8027 ( .A(n7803), .B(n8237), .Z(n7804) );
  NOR U8028 ( .A(n7805), .B(n7804), .Z(n7810) );
  NOR U8029 ( .A(n133), .B(n42), .Z(n7809) );
  IV U8030 ( .A(n7809), .Z(n7806) );
  NOR U8031 ( .A(n7810), .B(n7806), .Z(n7813) );
  XOR U8032 ( .A(n7808), .B(n7807), .Z(n7872) );
  IV U8033 ( .A(n7872), .Z(n7811) );
  XOR U8034 ( .A(n7810), .B(n7809), .Z(n7871) );
  NOR U8035 ( .A(n7811), .B(n7871), .Z(n7812) );
  NOR U8036 ( .A(n7813), .B(n7812), .Z(n7818) );
  NOR U8037 ( .A(n135), .B(n42), .Z(n7817) );
  IV U8038 ( .A(n7817), .Z(n7814) );
  NOR U8039 ( .A(n7818), .B(n7814), .Z(n7821) );
  XOR U8040 ( .A(n7816), .B(n7815), .Z(n7869) );
  IV U8041 ( .A(n7869), .Z(n7819) );
  XOR U8042 ( .A(n7818), .B(n7817), .Z(n7868) );
  NOR U8043 ( .A(n7819), .B(n7868), .Z(n7820) );
  NOR U8044 ( .A(n7821), .B(n7820), .Z(n7826) );
  NOR U8045 ( .A(n137), .B(n42), .Z(n7825) );
  IV U8046 ( .A(n7825), .Z(n7822) );
  NOR U8047 ( .A(n7826), .B(n7822), .Z(n7829) );
  XOR U8048 ( .A(n7824), .B(n7823), .Z(n7866) );
  IV U8049 ( .A(n7866), .Z(n7827) );
  XOR U8050 ( .A(n7826), .B(n7825), .Z(n7865) );
  NOR U8051 ( .A(n7827), .B(n7865), .Z(n7828) );
  NOR U8052 ( .A(n7829), .B(n7828), .Z(n7834) );
  NOR U8053 ( .A(n139), .B(n42), .Z(n7833) );
  IV U8054 ( .A(n7833), .Z(n7830) );
  NOR U8055 ( .A(n7834), .B(n7830), .Z(n7837) );
  XOR U8056 ( .A(n7832), .B(n7831), .Z(n7863) );
  IV U8057 ( .A(n7863), .Z(n7835) );
  XOR U8058 ( .A(n7834), .B(n7833), .Z(n7862) );
  NOR U8059 ( .A(n7835), .B(n7862), .Z(n7836) );
  NOR U8060 ( .A(n7837), .B(n7836), .Z(n7842) );
  NOR U8061 ( .A(n141), .B(n42), .Z(n7841) );
  IV U8062 ( .A(n7841), .Z(n7838) );
  NOR U8063 ( .A(n7842), .B(n7838), .Z(n7845) );
  XOR U8064 ( .A(n7840), .B(n7839), .Z(n7860) );
  IV U8065 ( .A(n7860), .Z(n7843) );
  XOR U8066 ( .A(n7842), .B(n7841), .Z(n7859) );
  NOR U8067 ( .A(n7843), .B(n7859), .Z(n7844) );
  NOR U8068 ( .A(n7845), .B(n7844), .Z(n8269) );
  XOR U8069 ( .A(n7847), .B(n7846), .Z(n8268) );
  NOR U8070 ( .A(n8269), .B(n8268), .Z(n7848) );
  NOR U8071 ( .A(n7849), .B(n7848), .Z(n7854) );
  NOR U8072 ( .A(n145), .B(n42), .Z(n7853) );
  IV U8073 ( .A(n7853), .Z(n7850) );
  NOR U8074 ( .A(n7854), .B(n7850), .Z(n7857) );
  XOR U8075 ( .A(n7852), .B(n7851), .Z(n8274) );
  IV U8076 ( .A(n8274), .Z(n7855) );
  XOR U8077 ( .A(n7854), .B(n7853), .Z(n8273) );
  NOR U8078 ( .A(n7855), .B(n8273), .Z(n7856) );
  NOR U8079 ( .A(n7857), .B(n7856), .Z(n8290) );
  NOR U8080 ( .A(n147), .B(n42), .Z(n8288) );
  XOR U8081 ( .A(n8290), .B(n8288), .Z(n8293) );
  XOR U8082 ( .A(n8291), .B(n8293), .Z(n8281) );
  NOR U8083 ( .A(n148), .B(n44), .Z(n8282) );
  IV U8084 ( .A(n8282), .Z(n7858) );
  NOR U8085 ( .A(n8281), .B(n7858), .Z(n8284) );
  XOR U8086 ( .A(n7860), .B(n7859), .Z(n8261) );
  NOR U8087 ( .A(n143), .B(n44), .Z(n8262) );
  IV U8088 ( .A(n8262), .Z(n7861) );
  NOR U8089 ( .A(n8261), .B(n7861), .Z(n8264) );
  XOR U8090 ( .A(n7863), .B(n7862), .Z(n8257) );
  NOR U8091 ( .A(n141), .B(n44), .Z(n8258) );
  IV U8092 ( .A(n8258), .Z(n7864) );
  NOR U8093 ( .A(n8257), .B(n7864), .Z(n8260) );
  XOR U8094 ( .A(n7866), .B(n7865), .Z(n8253) );
  NOR U8095 ( .A(n139), .B(n44), .Z(n8254) );
  IV U8096 ( .A(n8254), .Z(n7867) );
  NOR U8097 ( .A(n8253), .B(n7867), .Z(n8256) );
  XOR U8098 ( .A(n7869), .B(n7868), .Z(n8249) );
  NOR U8099 ( .A(n137), .B(n44), .Z(n8250) );
  IV U8100 ( .A(n8250), .Z(n7870) );
  NOR U8101 ( .A(n8249), .B(n7870), .Z(n8252) );
  XOR U8102 ( .A(n7872), .B(n7871), .Z(n8245) );
  NOR U8103 ( .A(n135), .B(n44), .Z(n8246) );
  IV U8104 ( .A(n8246), .Z(n7873) );
  NOR U8105 ( .A(n8245), .B(n7873), .Z(n8248) );
  XOR U8106 ( .A(n7875), .B(n7874), .Z(n8225) );
  NOR U8107 ( .A(n128), .B(n44), .Z(n8226) );
  IV U8108 ( .A(n8226), .Z(n7876) );
  NOR U8109 ( .A(n8225), .B(n7876), .Z(n8228) );
  NOR U8110 ( .A(n80), .B(n44), .Z(n8165) );
  NOR U8111 ( .A(n116), .B(n44), .Z(n8157) );
  NOR U8112 ( .A(n81), .B(n44), .Z(n8148) );
  NOR U8113 ( .A(n114), .B(n44), .Z(n8124) );
  XOR U8114 ( .A(n7878), .B(n7877), .Z(n10679) );
  IV U8115 ( .A(n10679), .Z(n7880) );
  NOR U8116 ( .A(n83), .B(n44), .Z(n10677) );
  IV U8117 ( .A(n10677), .Z(n7879) );
  NOR U8118 ( .A(n7880), .B(n7879), .Z(n8123) );
  NOR U8119 ( .A(n10677), .B(n10679), .Z(n8121) );
  XOR U8120 ( .A(n7882), .B(n7881), .Z(n7883) );
  XOR U8121 ( .A(n7884), .B(n7883), .Z(n8108) );
  NOR U8122 ( .A(n84), .B(n44), .Z(n8107) );
  IV U8123 ( .A(n8107), .Z(n7885) );
  NOR U8124 ( .A(n8108), .B(n7885), .Z(n8110) );
  NOR U8125 ( .A(n112), .B(n44), .Z(n8104) );
  IV U8126 ( .A(n8104), .Z(n8098) );
  XOR U8127 ( .A(n7887), .B(n7886), .Z(n7888) );
  NOR U8128 ( .A(n85), .B(n44), .Z(n7889) );
  NOR U8129 ( .A(n7888), .B(n7889), .Z(n8096) );
  IV U8130 ( .A(n7888), .Z(n10647) );
  IV U8131 ( .A(n7889), .Z(n10646) );
  NOR U8132 ( .A(n10647), .B(n10646), .Z(n8094) );
  NOR U8133 ( .A(n111), .B(n44), .Z(n7890) );
  IV U8134 ( .A(n7890), .Z(n8090) );
  NOR U8135 ( .A(n86), .B(n44), .Z(n7893) );
  XOR U8136 ( .A(n7892), .B(n7891), .Z(n7894) );
  NOR U8137 ( .A(n7893), .B(n7894), .Z(n8083) );
  IV U8138 ( .A(n7893), .Z(n10634) );
  IV U8139 ( .A(n7894), .Z(n10633) );
  NOR U8140 ( .A(n10634), .B(n10633), .Z(n8081) );
  XOR U8141 ( .A(n7896), .B(n7895), .Z(n7897) );
  IV U8142 ( .A(n7897), .Z(n8067) );
  NOR U8143 ( .A(n109), .B(n44), .Z(n8068) );
  IV U8144 ( .A(n8068), .Z(n7898) );
  NOR U8145 ( .A(n8067), .B(n7898), .Z(n8070) );
  XOR U8146 ( .A(n7900), .B(n7899), .Z(n7901) );
  XOR U8147 ( .A(n7902), .B(n7901), .Z(n8064) );
  NOR U8148 ( .A(n108), .B(n44), .Z(n8063) );
  IV U8149 ( .A(n8063), .Z(n7903) );
  NOR U8150 ( .A(n8064), .B(n7903), .Z(n8066) );
  NOR U8151 ( .A(n87), .B(n44), .Z(n7904) );
  IV U8152 ( .A(n7904), .Z(n8060) );
  XOR U8153 ( .A(n7906), .B(n7905), .Z(n8059) );
  IV U8154 ( .A(n8059), .Z(n7907) );
  NOR U8155 ( .A(n8060), .B(n7907), .Z(n8062) );
  XOR U8156 ( .A(n7909), .B(n7908), .Z(n8046) );
  NOR U8157 ( .A(n88), .B(n44), .Z(n8047) );
  IV U8158 ( .A(n8047), .Z(n7910) );
  NOR U8159 ( .A(n8046), .B(n7910), .Z(n8049) );
  IV U8160 ( .A(n7911), .Z(n7913) );
  XOR U8161 ( .A(n7913), .B(n7912), .Z(n8035) );
  NOR U8162 ( .A(n105), .B(n44), .Z(n8036) );
  IV U8163 ( .A(n8036), .Z(n7914) );
  NOR U8164 ( .A(n8035), .B(n7914), .Z(n8038) );
  XOR U8165 ( .A(n7916), .B(n7915), .Z(n7917) );
  XOR U8166 ( .A(n7918), .B(n7917), .Z(n8032) );
  NOR U8167 ( .A(n104), .B(n44), .Z(n8031) );
  IV U8168 ( .A(n8031), .Z(n7919) );
  NOR U8169 ( .A(n8032), .B(n7919), .Z(n8034) );
  XOR U8170 ( .A(n7921), .B(n7920), .Z(n8025) );
  NOR U8171 ( .A(n89), .B(n44), .Z(n8026) );
  NOR U8172 ( .A(n8025), .B(n8026), .Z(n8029) );
  XOR U8173 ( .A(n7923), .B(n7922), .Z(n8011) );
  IV U8174 ( .A(n8011), .Z(n10466) );
  NOR U8175 ( .A(n90), .B(n44), .Z(n8010) );
  IV U8176 ( .A(n8010), .Z(n10465) );
  NOR U8177 ( .A(n10466), .B(n10465), .Z(n8014) );
  XOR U8178 ( .A(n7925), .B(n7924), .Z(n7926) );
  XOR U8179 ( .A(n7927), .B(n7926), .Z(n8007) );
  NOR U8180 ( .A(n102), .B(n44), .Z(n8006) );
  IV U8181 ( .A(n8006), .Z(n7928) );
  NOR U8182 ( .A(n8007), .B(n7928), .Z(n8009) );
  XOR U8183 ( .A(n7930), .B(n7929), .Z(n7931) );
  NOR U8184 ( .A(n101), .B(n44), .Z(n7932) );
  NOR U8185 ( .A(n7931), .B(n7932), .Z(n8004) );
  XOR U8186 ( .A(n7932), .B(n7931), .Z(n10472) );
  IV U8187 ( .A(n10472), .Z(n8002) );
  XOR U8188 ( .A(n7934), .B(n7933), .Z(n7935) );
  XOR U8189 ( .A(n7936), .B(n7935), .Z(n7998) );
  NOR U8190 ( .A(n100), .B(n44), .Z(n7997) );
  IV U8191 ( .A(n7997), .Z(n7937) );
  NOR U8192 ( .A(n7998), .B(n7937), .Z(n8000) );
  NOR U8193 ( .A(n99), .B(n44), .Z(n7938) );
  IV U8194 ( .A(n7938), .Z(n7994) );
  XOR U8195 ( .A(n7940), .B(n7939), .Z(n7993) );
  IV U8196 ( .A(n7993), .Z(n7941) );
  NOR U8197 ( .A(n7994), .B(n7941), .Z(n7996) );
  XOR U8198 ( .A(n7943), .B(n7942), .Z(n7944) );
  NOR U8199 ( .A(n91), .B(n44), .Z(n7945) );
  NOR U8200 ( .A(n7944), .B(n7945), .Z(n7983) );
  IV U8201 ( .A(n7944), .Z(n10485) );
  IV U8202 ( .A(n7945), .Z(n10484) );
  NOR U8203 ( .A(n10485), .B(n10484), .Z(n7981) );
  IV U8204 ( .A(n7946), .Z(n7948) );
  XOR U8205 ( .A(n7948), .B(n7947), .Z(n7976) );
  NOR U8206 ( .A(n97), .B(n44), .Z(n7977) );
  IV U8207 ( .A(n7977), .Z(n7949) );
  NOR U8208 ( .A(n7976), .B(n7949), .Z(n7979) );
  XOR U8209 ( .A(n7951), .B(n7950), .Z(n7972) );
  NOR U8210 ( .A(n96), .B(n44), .Z(n7973) );
  IV U8211 ( .A(n7973), .Z(n7952) );
  NOR U8212 ( .A(n7972), .B(n7952), .Z(n7975) );
  XOR U8213 ( .A(n7954), .B(n7953), .Z(n7968) );
  NOR U8214 ( .A(n95), .B(n44), .Z(n7969) );
  IV U8215 ( .A(n7969), .Z(n7955) );
  NOR U8216 ( .A(n7968), .B(n7955), .Z(n7971) );
  NOR U8217 ( .A(n93), .B(n44), .Z(n11001) );
  IV U8218 ( .A(n11001), .Z(n7956) );
  NOR U8219 ( .A(n42), .B(n168), .Z(n7964) );
  IV U8220 ( .A(n7964), .Z(n7959) );
  NOR U8221 ( .A(n7956), .B(n7959), .Z(n7957) );
  IV U8222 ( .A(n7957), .Z(n7958) );
  NOR U8223 ( .A(n94), .B(n7958), .Z(n7967) );
  NOR U8224 ( .A(n7959), .B(n93), .Z(n7960) );
  XOR U8225 ( .A(n94), .B(n7960), .Z(n7961) );
  NOR U8226 ( .A(n44), .B(n7961), .Z(n7962) );
  IV U8227 ( .A(n7962), .Z(n10498) );
  XOR U8228 ( .A(n7964), .B(n7963), .Z(n10497) );
  IV U8229 ( .A(n10497), .Z(n7965) );
  NOR U8230 ( .A(n10498), .B(n7965), .Z(n7966) );
  NOR U8231 ( .A(n7967), .B(n7966), .Z(n10493) );
  XOR U8232 ( .A(n7969), .B(n7968), .Z(n10494) );
  NOR U8233 ( .A(n10493), .B(n10494), .Z(n7970) );
  NOR U8234 ( .A(n7971), .B(n7970), .Z(n10524) );
  XOR U8235 ( .A(n7973), .B(n7972), .Z(n10523) );
  NOR U8236 ( .A(n10524), .B(n10523), .Z(n7974) );
  NOR U8237 ( .A(n7975), .B(n7974), .Z(n10489) );
  XOR U8238 ( .A(n7977), .B(n7976), .Z(n10490) );
  NOR U8239 ( .A(n10489), .B(n10490), .Z(n7978) );
  NOR U8240 ( .A(n7979), .B(n7978), .Z(n10487) );
  IV U8241 ( .A(n10487), .Z(n7980) );
  NOR U8242 ( .A(n7981), .B(n7980), .Z(n7982) );
  NOR U8243 ( .A(n7983), .B(n7982), .Z(n7990) );
  IV U8244 ( .A(n7990), .Z(n7985) );
  NOR U8245 ( .A(n98), .B(n44), .Z(n7984) );
  IV U8246 ( .A(n7984), .Z(n7989) );
  NOR U8247 ( .A(n7985), .B(n7989), .Z(n7992) );
  IV U8248 ( .A(n7986), .Z(n7988) );
  XOR U8249 ( .A(n7988), .B(n7987), .Z(n10481) );
  XOR U8250 ( .A(n7990), .B(n7989), .Z(n10480) );
  NOR U8251 ( .A(n10481), .B(n10480), .Z(n7991) );
  NOR U8252 ( .A(n7992), .B(n7991), .Z(n10542) );
  XOR U8253 ( .A(n7994), .B(n7993), .Z(n10543) );
  NOR U8254 ( .A(n10542), .B(n10543), .Z(n7995) );
  NOR U8255 ( .A(n7996), .B(n7995), .Z(n10476) );
  XOR U8256 ( .A(n7998), .B(n7997), .Z(n10475) );
  NOR U8257 ( .A(n10476), .B(n10475), .Z(n7999) );
  NOR U8258 ( .A(n8000), .B(n7999), .Z(n10473) );
  IV U8259 ( .A(n10473), .Z(n8001) );
  NOR U8260 ( .A(n8002), .B(n8001), .Z(n8003) );
  NOR U8261 ( .A(n8004), .B(n8003), .Z(n8005) );
  IV U8262 ( .A(n8005), .Z(n10471) );
  XOR U8263 ( .A(n8007), .B(n8006), .Z(n10470) );
  NOR U8264 ( .A(n10471), .B(n10470), .Z(n8008) );
  NOR U8265 ( .A(n8009), .B(n8008), .Z(n10468) );
  NOR U8266 ( .A(n8011), .B(n8010), .Z(n8012) );
  NOR U8267 ( .A(n10468), .B(n8012), .Z(n8013) );
  NOR U8268 ( .A(n8014), .B(n8013), .Z(n8020) );
  NOR U8269 ( .A(n103), .B(n44), .Z(n8021) );
  IV U8270 ( .A(n8021), .Z(n8015) );
  NOR U8271 ( .A(n8020), .B(n8015), .Z(n8023) );
  XOR U8272 ( .A(n8017), .B(n8016), .Z(n8018) );
  XOR U8273 ( .A(n8019), .B(n8018), .Z(n10464) );
  XOR U8274 ( .A(n8021), .B(n8020), .Z(n10463) );
  NOR U8275 ( .A(n10464), .B(n10463), .Z(n8022) );
  NOR U8276 ( .A(n8023), .B(n8022), .Z(n8024) );
  IV U8277 ( .A(n8024), .Z(n10573) );
  XOR U8278 ( .A(n8026), .B(n8025), .Z(n8027) );
  IV U8279 ( .A(n8027), .Z(n10572) );
  NOR U8280 ( .A(n10573), .B(n10572), .Z(n8028) );
  NOR U8281 ( .A(n8029), .B(n8028), .Z(n8030) );
  IV U8282 ( .A(n8030), .Z(n10462) );
  XOR U8283 ( .A(n8032), .B(n8031), .Z(n10461) );
  NOR U8284 ( .A(n10462), .B(n10461), .Z(n8033) );
  NOR U8285 ( .A(n8034), .B(n8033), .Z(n10460) );
  XOR U8286 ( .A(n8036), .B(n8035), .Z(n10459) );
  NOR U8287 ( .A(n10460), .B(n10459), .Z(n8037) );
  NOR U8288 ( .A(n8038), .B(n8037), .Z(n8043) );
  NOR U8289 ( .A(n106), .B(n44), .Z(n8042) );
  IV U8290 ( .A(n8042), .Z(n8039) );
  NOR U8291 ( .A(n8043), .B(n8039), .Z(n8045) );
  XOR U8292 ( .A(n8041), .B(n8040), .Z(n10458) );
  XOR U8293 ( .A(n8043), .B(n8042), .Z(n10457) );
  NOR U8294 ( .A(n10458), .B(n10457), .Z(n8044) );
  NOR U8295 ( .A(n8045), .B(n8044), .Z(n10596) );
  XOR U8296 ( .A(n8047), .B(n8046), .Z(n10597) );
  NOR U8297 ( .A(n10596), .B(n10597), .Z(n8048) );
  NOR U8298 ( .A(n8049), .B(n8048), .Z(n8055) );
  NOR U8299 ( .A(n107), .B(n44), .Z(n8056) );
  IV U8300 ( .A(n8056), .Z(n8050) );
  NOR U8301 ( .A(n8055), .B(n8050), .Z(n8058) );
  XOR U8302 ( .A(n8052), .B(n8051), .Z(n8053) );
  XOR U8303 ( .A(n8054), .B(n8053), .Z(n10454) );
  XOR U8304 ( .A(n8056), .B(n8055), .Z(n10453) );
  NOR U8305 ( .A(n10454), .B(n10453), .Z(n8057) );
  NOR U8306 ( .A(n8058), .B(n8057), .Z(n10611) );
  XOR U8307 ( .A(n8060), .B(n8059), .Z(n10612) );
  NOR U8308 ( .A(n10611), .B(n10612), .Z(n8061) );
  NOR U8309 ( .A(n8062), .B(n8061), .Z(n10452) );
  XOR U8310 ( .A(n8064), .B(n8063), .Z(n10451) );
  NOR U8311 ( .A(n10452), .B(n10451), .Z(n8065) );
  NOR U8312 ( .A(n8066), .B(n8065), .Z(n10450) );
  XOR U8313 ( .A(n8068), .B(n8067), .Z(n10449) );
  NOR U8314 ( .A(n10450), .B(n10449), .Z(n8069) );
  NOR U8315 ( .A(n8070), .B(n8069), .Z(n8072) );
  NOR U8316 ( .A(n110), .B(n44), .Z(n8073) );
  IV U8317 ( .A(n8073), .Z(n8071) );
  NOR U8318 ( .A(n8072), .B(n8071), .Z(n8079) );
  XOR U8319 ( .A(n8073), .B(n8072), .Z(n10448) );
  XOR U8320 ( .A(n8075), .B(n8074), .Z(n8076) );
  XOR U8321 ( .A(n8077), .B(n8076), .Z(n10447) );
  NOR U8322 ( .A(n10448), .B(n10447), .Z(n8078) );
  NOR U8323 ( .A(n8079), .B(n8078), .Z(n10636) );
  IV U8324 ( .A(n10636), .Z(n8080) );
  NOR U8325 ( .A(n8081), .B(n8080), .Z(n8082) );
  NOR U8326 ( .A(n8083), .B(n8082), .Z(n8089) );
  IV U8327 ( .A(n8089), .Z(n8084) );
  NOR U8328 ( .A(n8090), .B(n8084), .Z(n8092) );
  XOR U8329 ( .A(n8086), .B(n8085), .Z(n8087) );
  XOR U8330 ( .A(n8088), .B(n8087), .Z(n10443) );
  XOR U8331 ( .A(n8090), .B(n8089), .Z(n10442) );
  NOR U8332 ( .A(n10443), .B(n10442), .Z(n8091) );
  NOR U8333 ( .A(n8092), .B(n8091), .Z(n10649) );
  IV U8334 ( .A(n10649), .Z(n8093) );
  NOR U8335 ( .A(n8094), .B(n8093), .Z(n8095) );
  NOR U8336 ( .A(n8096), .B(n8095), .Z(n8097) );
  IV U8337 ( .A(n8097), .Z(n8103) );
  NOR U8338 ( .A(n8098), .B(n8103), .Z(n8106) );
  XOR U8339 ( .A(n8100), .B(n8099), .Z(n8101) );
  XOR U8340 ( .A(n8102), .B(n8101), .Z(n10440) );
  XOR U8341 ( .A(n8104), .B(n8103), .Z(n10439) );
  NOR U8342 ( .A(n10440), .B(n10439), .Z(n8105) );
  NOR U8343 ( .A(n8106), .B(n8105), .Z(n10662) );
  XOR U8344 ( .A(n8108), .B(n8107), .Z(n10663) );
  NOR U8345 ( .A(n10662), .B(n10663), .Z(n8109) );
  NOR U8346 ( .A(n8110), .B(n8109), .Z(n8115) );
  XOR U8347 ( .A(n8112), .B(n8111), .Z(n8113) );
  XOR U8348 ( .A(n8114), .B(n8113), .Z(n10669) );
  NOR U8349 ( .A(n8115), .B(n10669), .Z(n8120) );
  IV U8350 ( .A(n10669), .Z(n8116) );
  IV U8351 ( .A(n8115), .Z(n10668) );
  NOR U8352 ( .A(n8116), .B(n10668), .Z(n8118) );
  NOR U8353 ( .A(n113), .B(n44), .Z(n10671) );
  IV U8354 ( .A(n10671), .Z(n8117) );
  NOR U8355 ( .A(n8118), .B(n8117), .Z(n8119) );
  NOR U8356 ( .A(n8120), .B(n8119), .Z(n10676) );
  NOR U8357 ( .A(n8121), .B(n10676), .Z(n8122) );
  NOR U8358 ( .A(n8123), .B(n8122), .Z(n8125) );
  IV U8359 ( .A(n8125), .Z(n10433) );
  NOR U8360 ( .A(n8124), .B(n10433), .Z(n8130) );
  IV U8361 ( .A(n8124), .Z(n10434) );
  NOR U8362 ( .A(n8125), .B(n10434), .Z(n8128) );
  XOR U8363 ( .A(n8127), .B(n8126), .Z(n10436) );
  NOR U8364 ( .A(n8128), .B(n10436), .Z(n8129) );
  NOR U8365 ( .A(n8130), .B(n8129), .Z(n8131) );
  IV U8366 ( .A(n8131), .Z(n8136) );
  NOR U8367 ( .A(n82), .B(n44), .Z(n8135) );
  IV U8368 ( .A(n8135), .Z(n8132) );
  NOR U8369 ( .A(n8136), .B(n8132), .Z(n8139) );
  XOR U8370 ( .A(n8134), .B(n8133), .Z(n10690) );
  IV U8371 ( .A(n10690), .Z(n8137) );
  XOR U8372 ( .A(n8136), .B(n8135), .Z(n10691) );
  NOR U8373 ( .A(n8137), .B(n10691), .Z(n8138) );
  NOR U8374 ( .A(n8139), .B(n8138), .Z(n8143) );
  XOR U8375 ( .A(n8141), .B(n8140), .Z(n8142) );
  NOR U8376 ( .A(n8143), .B(n8142), .Z(n8147) );
  XOR U8377 ( .A(n8143), .B(n8142), .Z(n8144) );
  IV U8378 ( .A(n8144), .Z(n10701) );
  NOR U8379 ( .A(n115), .B(n44), .Z(n10702) );
  IV U8380 ( .A(n10702), .Z(n8145) );
  NOR U8381 ( .A(n10701), .B(n8145), .Z(n8146) );
  NOR U8382 ( .A(n8147), .B(n8146), .Z(n8149) );
  IV U8383 ( .A(n8149), .Z(n10706) );
  NOR U8384 ( .A(n8148), .B(n10706), .Z(n8154) );
  IV U8385 ( .A(n8148), .Z(n10707) );
  NOR U8386 ( .A(n8149), .B(n10707), .Z(n8152) );
  XOR U8387 ( .A(n8151), .B(n8150), .Z(n10709) );
  NOR U8388 ( .A(n8152), .B(n10709), .Z(n8153) );
  NOR U8389 ( .A(n8154), .B(n8153), .Z(n8158) );
  NOR U8390 ( .A(n8157), .B(n8158), .Z(n8161) );
  XOR U8391 ( .A(n8156), .B(n8155), .Z(n10431) );
  IV U8392 ( .A(n8157), .Z(n8159) );
  XOR U8393 ( .A(n8159), .B(n8158), .Z(n10432) );
  NOR U8394 ( .A(n10431), .B(n10432), .Z(n8160) );
  NOR U8395 ( .A(n8161), .B(n8160), .Z(n8164) );
  NOR U8396 ( .A(n8165), .B(n8164), .Z(n8168) );
  XOR U8397 ( .A(n8163), .B(n8162), .Z(n10723) );
  XOR U8398 ( .A(n8165), .B(n8164), .Z(n10722) );
  IV U8399 ( .A(n10722), .Z(n8166) );
  NOR U8400 ( .A(n10723), .B(n8166), .Z(n8167) );
  NOR U8401 ( .A(n8168), .B(n8167), .Z(n8169) );
  IV U8402 ( .A(n8169), .Z(n8172) );
  NOR U8403 ( .A(n117), .B(n44), .Z(n8171) );
  IV U8404 ( .A(n8171), .Z(n8170) );
  NOR U8405 ( .A(n8172), .B(n8170), .Z(n8177) );
  XOR U8406 ( .A(n8172), .B(n8171), .Z(n10730) );
  XOR U8407 ( .A(n8174), .B(n8173), .Z(n10729) );
  IV U8408 ( .A(n10729), .Z(n8175) );
  NOR U8409 ( .A(n10730), .B(n8175), .Z(n8176) );
  NOR U8410 ( .A(n8177), .B(n8176), .Z(n8180) );
  NOR U8411 ( .A(n79), .B(n44), .Z(n8179) );
  IV U8412 ( .A(n8179), .Z(n8178) );
  NOR U8413 ( .A(n8180), .B(n8178), .Z(n8185) );
  XOR U8414 ( .A(n8180), .B(n8179), .Z(n10735) );
  XOR U8415 ( .A(n8182), .B(n8181), .Z(n10736) );
  IV U8416 ( .A(n10736), .Z(n8183) );
  NOR U8417 ( .A(n10735), .B(n8183), .Z(n8184) );
  NOR U8418 ( .A(n8185), .B(n8184), .Z(n8188) );
  NOR U8419 ( .A(n119), .B(n44), .Z(n8187) );
  IV U8420 ( .A(n8187), .Z(n8186) );
  NOR U8421 ( .A(n8188), .B(n8186), .Z(n8193) );
  XOR U8422 ( .A(n8188), .B(n8187), .Z(n10744) );
  IV U8423 ( .A(n8189), .Z(n8191) );
  XOR U8424 ( .A(n8191), .B(n8190), .Z(n10745) );
  NOR U8425 ( .A(n10744), .B(n10745), .Z(n8192) );
  NOR U8426 ( .A(n8193), .B(n8192), .Z(n8196) );
  NOR U8427 ( .A(n120), .B(n44), .Z(n8195) );
  IV U8428 ( .A(n8195), .Z(n8194) );
  NOR U8429 ( .A(n8196), .B(n8194), .Z(n8200) );
  XOR U8430 ( .A(n8196), .B(n8195), .Z(n10754) );
  XOR U8431 ( .A(n8198), .B(n8197), .Z(n10755) );
  NOR U8432 ( .A(n10754), .B(n10755), .Z(n8199) );
  NOR U8433 ( .A(n8200), .B(n8199), .Z(n8203) );
  NOR U8434 ( .A(n123), .B(n44), .Z(n8202) );
  IV U8435 ( .A(n8202), .Z(n8201) );
  NOR U8436 ( .A(n8203), .B(n8201), .Z(n8208) );
  XOR U8437 ( .A(n8203), .B(n8202), .Z(n10762) );
  XOR U8438 ( .A(n8205), .B(n8204), .Z(n10763) );
  IV U8439 ( .A(n10763), .Z(n8206) );
  NOR U8440 ( .A(n10762), .B(n8206), .Z(n8207) );
  NOR U8441 ( .A(n8208), .B(n8207), .Z(n8211) );
  NOR U8442 ( .A(n125), .B(n44), .Z(n8210) );
  IV U8443 ( .A(n8210), .Z(n8209) );
  NOR U8444 ( .A(n8211), .B(n8209), .Z(n8216) );
  XOR U8445 ( .A(n8211), .B(n8210), .Z(n10766) );
  XOR U8446 ( .A(n8213), .B(n8212), .Z(n10767) );
  IV U8447 ( .A(n10767), .Z(n8214) );
  NOR U8448 ( .A(n10766), .B(n8214), .Z(n8215) );
  NOR U8449 ( .A(n8216), .B(n8215), .Z(n8220) );
  XOR U8450 ( .A(n8218), .B(n8217), .Z(n8219) );
  NOR U8451 ( .A(n8220), .B(n8219), .Z(n8224) );
  XOR U8452 ( .A(n8220), .B(n8219), .Z(n10428) );
  IV U8453 ( .A(n10428), .Z(n8222) );
  NOR U8454 ( .A(n126), .B(n44), .Z(n10427) );
  IV U8455 ( .A(n10427), .Z(n8221) );
  NOR U8456 ( .A(n8222), .B(n8221), .Z(n8223) );
  NOR U8457 ( .A(n8224), .B(n8223), .Z(n10778) );
  XOR U8458 ( .A(n8226), .B(n8225), .Z(n10779) );
  NOR U8459 ( .A(n10778), .B(n10779), .Z(n8227) );
  NOR U8460 ( .A(n8228), .B(n8227), .Z(n8231) );
  NOR U8461 ( .A(n131), .B(n44), .Z(n8230) );
  IV U8462 ( .A(n8230), .Z(n8229) );
  NOR U8463 ( .A(n8231), .B(n8229), .Z(n8236) );
  XOR U8464 ( .A(n8231), .B(n8230), .Z(n10424) );
  XOR U8465 ( .A(n8233), .B(n8232), .Z(n10425) );
  IV U8466 ( .A(n10425), .Z(n8234) );
  NOR U8467 ( .A(n10424), .B(n8234), .Z(n8235) );
  NOR U8468 ( .A(n8236), .B(n8235), .Z(n8240) );
  XOR U8469 ( .A(n8238), .B(n8237), .Z(n8239) );
  NOR U8470 ( .A(n8240), .B(n8239), .Z(n8244) );
  XOR U8471 ( .A(n8240), .B(n8239), .Z(n8241) );
  IV U8472 ( .A(n8241), .Z(n10794) );
  NOR U8473 ( .A(n133), .B(n44), .Z(n10795) );
  IV U8474 ( .A(n10795), .Z(n8242) );
  NOR U8475 ( .A(n10794), .B(n8242), .Z(n8243) );
  NOR U8476 ( .A(n8244), .B(n8243), .Z(n10799) );
  XOR U8477 ( .A(n8246), .B(n8245), .Z(n10798) );
  NOR U8478 ( .A(n10799), .B(n10798), .Z(n8247) );
  NOR U8479 ( .A(n8248), .B(n8247), .Z(n10807) );
  XOR U8480 ( .A(n8250), .B(n8249), .Z(n10806) );
  NOR U8481 ( .A(n10807), .B(n10806), .Z(n8251) );
  NOR U8482 ( .A(n8252), .B(n8251), .Z(n10815) );
  XOR U8483 ( .A(n8254), .B(n8253), .Z(n10814) );
  NOR U8484 ( .A(n10815), .B(n10814), .Z(n8255) );
  NOR U8485 ( .A(n8256), .B(n8255), .Z(n10823) );
  XOR U8486 ( .A(n8258), .B(n8257), .Z(n10822) );
  NOR U8487 ( .A(n10823), .B(n10822), .Z(n8259) );
  NOR U8488 ( .A(n8260), .B(n8259), .Z(n10831) );
  XOR U8489 ( .A(n8262), .B(n8261), .Z(n10830) );
  NOR U8490 ( .A(n10831), .B(n10830), .Z(n8263) );
  NOR U8491 ( .A(n8264), .B(n8263), .Z(n8267) );
  NOR U8492 ( .A(n145), .B(n44), .Z(n8266) );
  IV U8493 ( .A(n8266), .Z(n8265) );
  NOR U8494 ( .A(n8267), .B(n8265), .Z(n8272) );
  XOR U8495 ( .A(n8267), .B(n8266), .Z(n10421) );
  XOR U8496 ( .A(n8269), .B(n8268), .Z(n10422) );
  IV U8497 ( .A(n10422), .Z(n8270) );
  NOR U8498 ( .A(n10421), .B(n8270), .Z(n8271) );
  NOR U8499 ( .A(n8272), .B(n8271), .Z(n8276) );
  XOR U8500 ( .A(n8274), .B(n8273), .Z(n8275) );
  NOR U8501 ( .A(n8276), .B(n8275), .Z(n8280) );
  XOR U8502 ( .A(n8276), .B(n8275), .Z(n8277) );
  IV U8503 ( .A(n8277), .Z(n10845) );
  NOR U8504 ( .A(n147), .B(n44), .Z(n10846) );
  IV U8505 ( .A(n10846), .Z(n8278) );
  NOR U8506 ( .A(n10845), .B(n8278), .Z(n8279) );
  NOR U8507 ( .A(n8280), .B(n8279), .Z(n10850) );
  XOR U8508 ( .A(n8282), .B(n8281), .Z(n10849) );
  NOR U8509 ( .A(n10850), .B(n10849), .Z(n8283) );
  NOR U8510 ( .A(n8284), .B(n8283), .Z(n8287) );
  NOR U8511 ( .A(n150), .B(n44), .Z(n8286) );
  IV U8512 ( .A(n8286), .Z(n8285) );
  NOR U8513 ( .A(n8287), .B(n8285), .Z(n8485) );
  XOR U8514 ( .A(n8287), .B(n8286), .Z(n10418) );
  IV U8515 ( .A(n8288), .Z(n8289) );
  NOR U8516 ( .A(n8290), .B(n8289), .Z(n8295) );
  IV U8517 ( .A(n8291), .Z(n8292) );
  NOR U8518 ( .A(n8293), .B(n8292), .Z(n8294) );
  NOR U8519 ( .A(n8295), .B(n8294), .Z(n8491) );
  IV U8520 ( .A(n8296), .Z(n8297) );
  NOR U8521 ( .A(n8298), .B(n8297), .Z(n8302) );
  NOR U8522 ( .A(n8300), .B(n8299), .Z(n8301) );
  NOR U8523 ( .A(n8302), .B(n8301), .Z(n8303) );
  IV U8524 ( .A(n8303), .Z(n8497) );
  NOR U8525 ( .A(n147), .B(n43), .Z(n8495) );
  NOR U8526 ( .A(n8305), .B(n8304), .Z(n8309) );
  NOR U8527 ( .A(n8307), .B(n8306), .Z(n8308) );
  NOR U8528 ( .A(n8309), .B(n8308), .Z(n8504) );
  NOR U8529 ( .A(n145), .B(n118), .Z(n8501) );
  IV U8530 ( .A(n8310), .Z(n8311) );
  NOR U8531 ( .A(n8312), .B(n8311), .Z(n8316) );
  NOR U8532 ( .A(n8314), .B(n8313), .Z(n8315) );
  NOR U8533 ( .A(n8316), .B(n8315), .Z(n8511) );
  IV U8534 ( .A(n8317), .Z(n8318) );
  NOR U8535 ( .A(n8319), .B(n8318), .Z(n8323) );
  NOR U8536 ( .A(n8321), .B(n8320), .Z(n8322) );
  NOR U8537 ( .A(n8323), .B(n8322), .Z(n8517) );
  NOR U8538 ( .A(n141), .B(n122), .Z(n8515) );
  IV U8539 ( .A(n8515), .Z(n8481) );
  IV U8540 ( .A(n8324), .Z(n8326) );
  NOR U8541 ( .A(n8326), .B(n8325), .Z(n8330) );
  NOR U8542 ( .A(n8328), .B(n8327), .Z(n8329) );
  NOR U8543 ( .A(n8330), .B(n8329), .Z(n8331) );
  IV U8544 ( .A(n8331), .Z(n8660) );
  NOR U8545 ( .A(n139), .B(n124), .Z(n8658) );
  XOR U8546 ( .A(n8660), .B(n8658), .Z(n8661) );
  NOR U8547 ( .A(n8333), .B(n8332), .Z(n8338) );
  IV U8548 ( .A(n8334), .Z(n8335) );
  NOR U8549 ( .A(n8336), .B(n8335), .Z(n8337) );
  NOR U8550 ( .A(n8338), .B(n8337), .Z(n8523) );
  NOR U8551 ( .A(n137), .B(n127), .Z(n8521) );
  IV U8552 ( .A(n8521), .Z(n8480) );
  NOR U8553 ( .A(n8340), .B(n8339), .Z(n8346) );
  IV U8554 ( .A(n8341), .Z(n8344) );
  IV U8555 ( .A(n8342), .Z(n8343) );
  NOR U8556 ( .A(n8344), .B(n8343), .Z(n8345) );
  NOR U8557 ( .A(n8346), .B(n8345), .Z(n8652) );
  IV U8558 ( .A(n8652), .Z(n8478) );
  NOR U8559 ( .A(n8348), .B(n8347), .Z(n8352) );
  NOR U8560 ( .A(n8350), .B(n8349), .Z(n8351) );
  NOR U8561 ( .A(n8352), .B(n8351), .Z(n8529) );
  NOR U8562 ( .A(n133), .B(n130), .Z(n8527) );
  IV U8563 ( .A(n8527), .Z(n8477) );
  NOR U8564 ( .A(n8354), .B(n8353), .Z(n8359) );
  IV U8565 ( .A(n8355), .Z(n8356) );
  NOR U8566 ( .A(n8357), .B(n8356), .Z(n8358) );
  NOR U8567 ( .A(n8359), .B(n8358), .Z(n8360) );
  IV U8568 ( .A(n8360), .Z(n8534) );
  NOR U8569 ( .A(n131), .B(n132), .Z(n8532) );
  XOR U8570 ( .A(n8534), .B(n8532), .Z(n8535) );
  NOR U8571 ( .A(n8362), .B(n8361), .Z(n8367) );
  IV U8572 ( .A(n8363), .Z(n8364) );
  NOR U8573 ( .A(n8365), .B(n8364), .Z(n8366) );
  NOR U8574 ( .A(n8367), .B(n8366), .Z(n8542) );
  NOR U8575 ( .A(n128), .B(n134), .Z(n8540) );
  IV U8576 ( .A(n8540), .Z(n8476) );
  NOR U8577 ( .A(n8369), .B(n8368), .Z(n8374) );
  IV U8578 ( .A(n8370), .Z(n8372) );
  NOR U8579 ( .A(n8372), .B(n8371), .Z(n8373) );
  NOR U8580 ( .A(n8374), .B(n8373), .Z(n8375) );
  IV U8581 ( .A(n8375), .Z(n8547) );
  NOR U8582 ( .A(n126), .B(n136), .Z(n8545) );
  XOR U8583 ( .A(n8547), .B(n8545), .Z(n8548) );
  NOR U8584 ( .A(n8377), .B(n8376), .Z(n8382) );
  IV U8585 ( .A(n8378), .Z(n8379) );
  NOR U8586 ( .A(n8380), .B(n8379), .Z(n8381) );
  NOR U8587 ( .A(n8382), .B(n8381), .Z(n8555) );
  NOR U8588 ( .A(n125), .B(n138), .Z(n8553) );
  IV U8589 ( .A(n8553), .Z(n8475) );
  IV U8590 ( .A(n8383), .Z(n8384) );
  NOR U8591 ( .A(n8385), .B(n8384), .Z(n8389) );
  NOR U8592 ( .A(n8387), .B(n8386), .Z(n8388) );
  NOR U8593 ( .A(n8389), .B(n8388), .Z(n8560) );
  NOR U8594 ( .A(n123), .B(n140), .Z(n8559) );
  NOR U8595 ( .A(n8391), .B(n8390), .Z(n8395) );
  NOR U8596 ( .A(n8393), .B(n8392), .Z(n8394) );
  NOR U8597 ( .A(n8395), .B(n8394), .Z(n8570) );
  NOR U8598 ( .A(n120), .B(n142), .Z(n8567) );
  IV U8599 ( .A(n8396), .Z(n8397) );
  NOR U8600 ( .A(n8398), .B(n8397), .Z(n8402) );
  NOR U8601 ( .A(n8400), .B(n8399), .Z(n8401) );
  NOR U8602 ( .A(n8402), .B(n8401), .Z(n8648) );
  NOR U8603 ( .A(n8404), .B(n8403), .Z(n8408) );
  NOR U8604 ( .A(n8406), .B(n8405), .Z(n8407) );
  NOR U8605 ( .A(n8408), .B(n8407), .Z(n8576) );
  NOR U8606 ( .A(n79), .B(n146), .Z(n8574) );
  IV U8607 ( .A(n8409), .Z(n8410) );
  NOR U8608 ( .A(n8411), .B(n8410), .Z(n8415) );
  NOR U8609 ( .A(n8413), .B(n8412), .Z(n8414) );
  NOR U8610 ( .A(n8415), .B(n8414), .Z(n8640) );
  NOR U8611 ( .A(n8417), .B(n8416), .Z(n8421) );
  NOR U8612 ( .A(n8419), .B(n8418), .Z(n8420) );
  NOR U8613 ( .A(n8421), .B(n8420), .Z(n8582) );
  NOR U8614 ( .A(n80), .B(n151), .Z(n8580) );
  NOR U8615 ( .A(n8423), .B(n8422), .Z(n8427) );
  NOR U8616 ( .A(n8425), .B(n8424), .Z(n8426) );
  NOR U8617 ( .A(n8427), .B(n8426), .Z(n8595) );
  NOR U8618 ( .A(n81), .B(n154), .Z(n8593) );
  IV U8619 ( .A(n8428), .Z(n8429) );
  NOR U8620 ( .A(n8430), .B(n8429), .Z(n8434) );
  NOR U8621 ( .A(n8432), .B(n8431), .Z(n8433) );
  NOR U8622 ( .A(n8434), .B(n8433), .Z(n8602) );
  NOR U8623 ( .A(n8436), .B(n8435), .Z(n8440) );
  NOR U8624 ( .A(n8438), .B(n8437), .Z(n8439) );
  NOR U8625 ( .A(n8440), .B(n8439), .Z(n8608) );
  NOR U8626 ( .A(n82), .B(n159), .Z(n8606) );
  NOR U8627 ( .A(n8442), .B(n8441), .Z(n8446) );
  NOR U8628 ( .A(n8444), .B(n8443), .Z(n8445) );
  NOR U8629 ( .A(n8446), .B(n8445), .Z(n8621) );
  NOR U8630 ( .A(n83), .B(n162), .Z(n8619) );
  IV U8631 ( .A(n8619), .Z(n8455) );
  IV U8632 ( .A(n8447), .Z(n8448) );
  NOR U8633 ( .A(n8449), .B(n8448), .Z(n8453) );
  NOR U8634 ( .A(n8451), .B(n8450), .Z(n8452) );
  NOR U8635 ( .A(n8453), .B(n8452), .Z(n8626) );
  NOR U8636 ( .A(n164), .B(n113), .Z(n8624) );
  XOR U8637 ( .A(n8626), .B(n8624), .Z(n8628) );
  NOR U8638 ( .A(n166), .B(n84), .Z(n8454) );
  IV U8639 ( .A(n8454), .Z(n8627) );
  XOR U8640 ( .A(n8628), .B(n8627), .Z(n8618) );
  XOR U8641 ( .A(n8455), .B(n8618), .Z(n8620) );
  XOR U8642 ( .A(n8621), .B(n8620), .Z(n8615) );
  IV U8643 ( .A(n8456), .Z(n8457) );
  NOR U8644 ( .A(n8458), .B(n8457), .Z(n8462) );
  NOR U8645 ( .A(n8460), .B(n8459), .Z(n8461) );
  NOR U8646 ( .A(n8462), .B(n8461), .Z(n8613) );
  NOR U8647 ( .A(n114), .B(n160), .Z(n8611) );
  XOR U8648 ( .A(n8613), .B(n8611), .Z(n8614) );
  XOR U8649 ( .A(n8615), .B(n8614), .Z(n8605) );
  XOR U8650 ( .A(n8606), .B(n8605), .Z(n8463) );
  IV U8651 ( .A(n8463), .Z(n8607) );
  XOR U8652 ( .A(n8608), .B(n8607), .Z(n8600) );
  NOR U8653 ( .A(n115), .B(n157), .Z(n8598) );
  XOR U8654 ( .A(n8600), .B(n8598), .Z(n8601) );
  XOR U8655 ( .A(n8602), .B(n8601), .Z(n8592) );
  XOR U8656 ( .A(n8593), .B(n8592), .Z(n8464) );
  IV U8657 ( .A(n8464), .Z(n8594) );
  XOR U8658 ( .A(n8595), .B(n8594), .Z(n8589) );
  IV U8659 ( .A(n8465), .Z(n8466) );
  NOR U8660 ( .A(n8467), .B(n8466), .Z(n8471) );
  NOR U8661 ( .A(n8469), .B(n8468), .Z(n8470) );
  NOR U8662 ( .A(n8471), .B(n8470), .Z(n8587) );
  NOR U8663 ( .A(n116), .B(n152), .Z(n8585) );
  XOR U8664 ( .A(n8587), .B(n8585), .Z(n8588) );
  XOR U8665 ( .A(n8589), .B(n8588), .Z(n8579) );
  XOR U8666 ( .A(n8580), .B(n8579), .Z(n8472) );
  IV U8667 ( .A(n8472), .Z(n8581) );
  XOR U8668 ( .A(n8582), .B(n8581), .Z(n8638) );
  NOR U8669 ( .A(n117), .B(n149), .Z(n8636) );
  XOR U8670 ( .A(n8638), .B(n8636), .Z(n8639) );
  XOR U8671 ( .A(n8640), .B(n8639), .Z(n8573) );
  XOR U8672 ( .A(n8574), .B(n8573), .Z(n8473) );
  IV U8673 ( .A(n8473), .Z(n8575) );
  XOR U8674 ( .A(n8576), .B(n8575), .Z(n8646) );
  NOR U8675 ( .A(n119), .B(n144), .Z(n8644) );
  XOR U8676 ( .A(n8646), .B(n8644), .Z(n8647) );
  XOR U8677 ( .A(n8648), .B(n8647), .Z(n8566) );
  XOR U8678 ( .A(n8567), .B(n8566), .Z(n8568) );
  XOR U8679 ( .A(n8570), .B(n8568), .Z(n8558) );
  XOR U8680 ( .A(n8559), .B(n8558), .Z(n8474) );
  IV U8681 ( .A(n8474), .Z(n8561) );
  XOR U8682 ( .A(n8560), .B(n8561), .Z(n8552) );
  XOR U8683 ( .A(n8475), .B(n8552), .Z(n8554) );
  XOR U8684 ( .A(n8555), .B(n8554), .Z(n8549) );
  XOR U8685 ( .A(n8548), .B(n8549), .Z(n8539) );
  XOR U8686 ( .A(n8476), .B(n8539), .Z(n8541) );
  XOR U8687 ( .A(n8542), .B(n8541), .Z(n8536) );
  XOR U8688 ( .A(n8535), .B(n8536), .Z(n8526) );
  XOR U8689 ( .A(n8477), .B(n8526), .Z(n8528) );
  XOR U8690 ( .A(n8529), .B(n8528), .Z(n8653) );
  XOR U8691 ( .A(n8478), .B(n8653), .Z(n8655) );
  NOR U8692 ( .A(n135), .B(n129), .Z(n8479) );
  IV U8693 ( .A(n8479), .Z(n8654) );
  XOR U8694 ( .A(n8655), .B(n8654), .Z(n8520) );
  XOR U8695 ( .A(n8480), .B(n8520), .Z(n8522) );
  XOR U8696 ( .A(n8523), .B(n8522), .Z(n8662) );
  XOR U8697 ( .A(n8661), .B(n8662), .Z(n8514) );
  XOR U8698 ( .A(n8481), .B(n8514), .Z(n8516) );
  XOR U8699 ( .A(n8517), .B(n8516), .Z(n8509) );
  NOR U8700 ( .A(n143), .B(n121), .Z(n8507) );
  XOR U8701 ( .A(n8509), .B(n8507), .Z(n8510) );
  XOR U8702 ( .A(n8511), .B(n8510), .Z(n8500) );
  XOR U8703 ( .A(n8501), .B(n8500), .Z(n8502) );
  XOR U8704 ( .A(n8504), .B(n8502), .Z(n8494) );
  XOR U8705 ( .A(n8495), .B(n8494), .Z(n8482) );
  IV U8706 ( .A(n8482), .Z(n8496) );
  XOR U8707 ( .A(n8497), .B(n8496), .Z(n8489) );
  NOR U8708 ( .A(n148), .B(n42), .Z(n8487) );
  XOR U8709 ( .A(n8489), .B(n8487), .Z(n8490) );
  XOR U8710 ( .A(n8491), .B(n8490), .Z(n10419) );
  IV U8711 ( .A(n10419), .Z(n8483) );
  NOR U8712 ( .A(n10418), .B(n8483), .Z(n8484) );
  NOR U8713 ( .A(n8485), .B(n8484), .Z(n8668) );
  NOR U8714 ( .A(n153), .B(n44), .Z(n8667) );
  IV U8715 ( .A(n8667), .Z(n8486) );
  NOR U8716 ( .A(n8668), .B(n8486), .Z(n8671) );
  IV U8717 ( .A(n8487), .Z(n8488) );
  NOR U8718 ( .A(n8489), .B(n8488), .Z(n8493) );
  NOR U8719 ( .A(n8491), .B(n8490), .Z(n8492) );
  NOR U8720 ( .A(n8493), .B(n8492), .Z(n8865) );
  NOR U8721 ( .A(n150), .B(n42), .Z(n8861) );
  NOR U8722 ( .A(n8495), .B(n8494), .Z(n8499) );
  NOR U8723 ( .A(n8497), .B(n8496), .Z(n8498) );
  NOR U8724 ( .A(n8499), .B(n8498), .Z(n8675) );
  NOR U8725 ( .A(n8501), .B(n8500), .Z(n8506) );
  IV U8726 ( .A(n8502), .Z(n8503) );
  NOR U8727 ( .A(n8504), .B(n8503), .Z(n8505) );
  NOR U8728 ( .A(n8506), .B(n8505), .Z(n8684) );
  NOR U8729 ( .A(n147), .B(n118), .Z(n8682) );
  IV U8730 ( .A(n8507), .Z(n8508) );
  NOR U8731 ( .A(n8509), .B(n8508), .Z(n8513) );
  NOR U8732 ( .A(n8511), .B(n8510), .Z(n8512) );
  NOR U8733 ( .A(n8513), .B(n8512), .Z(n8693) );
  NOR U8734 ( .A(n8515), .B(n8514), .Z(n8519) );
  NOR U8735 ( .A(n8517), .B(n8516), .Z(n8518) );
  NOR U8736 ( .A(n8519), .B(n8518), .Z(n8699) );
  NOR U8737 ( .A(n143), .B(n122), .Z(n8697) );
  NOR U8738 ( .A(n8521), .B(n8520), .Z(n8525) );
  NOR U8739 ( .A(n8523), .B(n8522), .Z(n8524) );
  NOR U8740 ( .A(n8525), .B(n8524), .Z(n8706) );
  NOR U8741 ( .A(n139), .B(n127), .Z(n8704) );
  NOR U8742 ( .A(n8527), .B(n8526), .Z(n8531) );
  NOR U8743 ( .A(n8529), .B(n8528), .Z(n8530) );
  NOR U8744 ( .A(n8531), .B(n8530), .Z(n8721) );
  NOR U8745 ( .A(n135), .B(n130), .Z(n8718) );
  IV U8746 ( .A(n8532), .Z(n8533) );
  NOR U8747 ( .A(n8534), .B(n8533), .Z(n8538) );
  NOR U8748 ( .A(n8536), .B(n8535), .Z(n8537) );
  NOR U8749 ( .A(n8538), .B(n8537), .Z(n8724) );
  NOR U8750 ( .A(n8540), .B(n8539), .Z(n8544) );
  NOR U8751 ( .A(n8542), .B(n8541), .Z(n8543) );
  NOR U8752 ( .A(n8544), .B(n8543), .Z(n8736) );
  NOR U8753 ( .A(n131), .B(n134), .Z(n8734) );
  NOR U8754 ( .A(n128), .B(n136), .Z(n8743) );
  IV U8755 ( .A(n8545), .Z(n8546) );
  NOR U8756 ( .A(n8547), .B(n8546), .Z(n8551) );
  NOR U8757 ( .A(n8549), .B(n8548), .Z(n8550) );
  NOR U8758 ( .A(n8551), .B(n8550), .Z(n8739) );
  NOR U8759 ( .A(n8553), .B(n8552), .Z(n8557) );
  NOR U8760 ( .A(n8555), .B(n8554), .Z(n8556) );
  NOR U8761 ( .A(n8557), .B(n8556), .Z(n8751) );
  NOR U8762 ( .A(n126), .B(n138), .Z(n8748) );
  NOR U8763 ( .A(n8559), .B(n8558), .Z(n8564) );
  IV U8764 ( .A(n8560), .Z(n8562) );
  NOR U8765 ( .A(n8562), .B(n8561), .Z(n8563) );
  NOR U8766 ( .A(n8564), .B(n8563), .Z(n8565) );
  IV U8767 ( .A(n8565), .Z(n8840) );
  NOR U8768 ( .A(n125), .B(n140), .Z(n8838) );
  XOR U8769 ( .A(n8840), .B(n8838), .Z(n8841) );
  NOR U8770 ( .A(n8567), .B(n8566), .Z(n8572) );
  IV U8771 ( .A(n8568), .Z(n8569) );
  NOR U8772 ( .A(n8570), .B(n8569), .Z(n8571) );
  NOR U8773 ( .A(n8572), .B(n8571), .Z(n8757) );
  NOR U8774 ( .A(n123), .B(n142), .Z(n8755) );
  IV U8775 ( .A(n8755), .Z(n8651) );
  NOR U8776 ( .A(n8574), .B(n8573), .Z(n8578) );
  NOR U8777 ( .A(n8576), .B(n8575), .Z(n8577) );
  NOR U8778 ( .A(n8578), .B(n8577), .Z(n8763) );
  NOR U8779 ( .A(n119), .B(n146), .Z(n8761) );
  NOR U8780 ( .A(n8580), .B(n8579), .Z(n8584) );
  NOR U8781 ( .A(n8582), .B(n8581), .Z(n8583) );
  NOR U8782 ( .A(n8584), .B(n8583), .Z(n8769) );
  NOR U8783 ( .A(n117), .B(n151), .Z(n8767) );
  IV U8784 ( .A(n8585), .Z(n8586) );
  NOR U8785 ( .A(n8587), .B(n8586), .Z(n8591) );
  NOR U8786 ( .A(n8589), .B(n8588), .Z(n8590) );
  NOR U8787 ( .A(n8591), .B(n8590), .Z(n8819) );
  NOR U8788 ( .A(n8593), .B(n8592), .Z(n8597) );
  NOR U8789 ( .A(n8595), .B(n8594), .Z(n8596) );
  NOR U8790 ( .A(n8597), .B(n8596), .Z(n8775) );
  NOR U8791 ( .A(n116), .B(n154), .Z(n8773) );
  IV U8792 ( .A(n8598), .Z(n8599) );
  NOR U8793 ( .A(n8600), .B(n8599), .Z(n8604) );
  NOR U8794 ( .A(n8602), .B(n8601), .Z(n8603) );
  NOR U8795 ( .A(n8604), .B(n8603), .Z(n8782) );
  NOR U8796 ( .A(n8606), .B(n8605), .Z(n8610) );
  NOR U8797 ( .A(n8608), .B(n8607), .Z(n8609) );
  NOR U8798 ( .A(n8610), .B(n8609), .Z(n8788) );
  NOR U8799 ( .A(n115), .B(n159), .Z(n8786) );
  IV U8800 ( .A(n8611), .Z(n8612) );
  NOR U8801 ( .A(n8613), .B(n8612), .Z(n8617) );
  NOR U8802 ( .A(n8615), .B(n8614), .Z(n8616) );
  NOR U8803 ( .A(n8617), .B(n8616), .Z(n8795) );
  NOR U8804 ( .A(n8619), .B(n8618), .Z(n8623) );
  NOR U8805 ( .A(n8621), .B(n8620), .Z(n8622) );
  NOR U8806 ( .A(n8623), .B(n8622), .Z(n8801) );
  NOR U8807 ( .A(n114), .B(n162), .Z(n8799) );
  IV U8808 ( .A(n8799), .Z(n8632) );
  IV U8809 ( .A(n8624), .Z(n8625) );
  NOR U8810 ( .A(n8626), .B(n8625), .Z(n8630) );
  NOR U8811 ( .A(n8628), .B(n8627), .Z(n8629) );
  NOR U8812 ( .A(n8630), .B(n8629), .Z(n8806) );
  NOR U8813 ( .A(n164), .B(n83), .Z(n8804) );
  XOR U8814 ( .A(n8806), .B(n8804), .Z(n8808) );
  NOR U8815 ( .A(n166), .B(n113), .Z(n8631) );
  IV U8816 ( .A(n8631), .Z(n8807) );
  XOR U8817 ( .A(n8808), .B(n8807), .Z(n8798) );
  XOR U8818 ( .A(n8632), .B(n8798), .Z(n8800) );
  XOR U8819 ( .A(n8801), .B(n8800), .Z(n8793) );
  NOR U8820 ( .A(n82), .B(n160), .Z(n8791) );
  XOR U8821 ( .A(n8793), .B(n8791), .Z(n8794) );
  XOR U8822 ( .A(n8795), .B(n8794), .Z(n8785) );
  XOR U8823 ( .A(n8786), .B(n8785), .Z(n8633) );
  IV U8824 ( .A(n8633), .Z(n8787) );
  XOR U8825 ( .A(n8788), .B(n8787), .Z(n8780) );
  NOR U8826 ( .A(n81), .B(n157), .Z(n8778) );
  XOR U8827 ( .A(n8780), .B(n8778), .Z(n8781) );
  XOR U8828 ( .A(n8782), .B(n8781), .Z(n8772) );
  XOR U8829 ( .A(n8773), .B(n8772), .Z(n8634) );
  IV U8830 ( .A(n8634), .Z(n8774) );
  XOR U8831 ( .A(n8775), .B(n8774), .Z(n8817) );
  NOR U8832 ( .A(n80), .B(n152), .Z(n8815) );
  XOR U8833 ( .A(n8817), .B(n8815), .Z(n8818) );
  XOR U8834 ( .A(n8819), .B(n8818), .Z(n8766) );
  XOR U8835 ( .A(n8767), .B(n8766), .Z(n8635) );
  IV U8836 ( .A(n8635), .Z(n8768) );
  XOR U8837 ( .A(n8769), .B(n8768), .Z(n8827) );
  IV U8838 ( .A(n8636), .Z(n8637) );
  NOR U8839 ( .A(n8638), .B(n8637), .Z(n8642) );
  NOR U8840 ( .A(n8640), .B(n8639), .Z(n8641) );
  NOR U8841 ( .A(n8642), .B(n8641), .Z(n8825) );
  NOR U8842 ( .A(n79), .B(n149), .Z(n8823) );
  XOR U8843 ( .A(n8825), .B(n8823), .Z(n8826) );
  XOR U8844 ( .A(n8827), .B(n8826), .Z(n8760) );
  XOR U8845 ( .A(n8761), .B(n8760), .Z(n8643) );
  IV U8846 ( .A(n8643), .Z(n8762) );
  XOR U8847 ( .A(n8763), .B(n8762), .Z(n8835) );
  IV U8848 ( .A(n8644), .Z(n8645) );
  NOR U8849 ( .A(n8646), .B(n8645), .Z(n8650) );
  NOR U8850 ( .A(n8648), .B(n8647), .Z(n8649) );
  NOR U8851 ( .A(n8650), .B(n8649), .Z(n8833) );
  NOR U8852 ( .A(n120), .B(n144), .Z(n8831) );
  XOR U8853 ( .A(n8833), .B(n8831), .Z(n8834) );
  XOR U8854 ( .A(n8835), .B(n8834), .Z(n8754) );
  XOR U8855 ( .A(n8651), .B(n8754), .Z(n8756) );
  XOR U8856 ( .A(n8757), .B(n8756), .Z(n8842) );
  XOR U8857 ( .A(n8841), .B(n8842), .Z(n8747) );
  XOR U8858 ( .A(n8748), .B(n8747), .Z(n8749) );
  XOR U8859 ( .A(n8751), .B(n8749), .Z(n8740) );
  XOR U8860 ( .A(n8739), .B(n8740), .Z(n8742) );
  XOR U8861 ( .A(n8743), .B(n8742), .Z(n8732) );
  XOR U8862 ( .A(n8734), .B(n8732), .Z(n8735) );
  XOR U8863 ( .A(n8736), .B(n8735), .Z(n8725) );
  XOR U8864 ( .A(n8724), .B(n8725), .Z(n8726) );
  NOR U8865 ( .A(n133), .B(n132), .Z(n8727) );
  XOR U8866 ( .A(n8726), .B(n8727), .Z(n8717) );
  XOR U8867 ( .A(n8718), .B(n8717), .Z(n8719) );
  XOR U8868 ( .A(n8721), .B(n8719), .Z(n8712) );
  NOR U8869 ( .A(n137), .B(n129), .Z(n8711) );
  NOR U8870 ( .A(n8653), .B(n8652), .Z(n8657) );
  NOR U8871 ( .A(n8655), .B(n8654), .Z(n8656) );
  NOR U8872 ( .A(n8657), .B(n8656), .Z(n8709) );
  XOR U8873 ( .A(n8711), .B(n8709), .Z(n8713) );
  XOR U8874 ( .A(n8712), .B(n8713), .Z(n8702) );
  XOR U8875 ( .A(n8704), .B(n8702), .Z(n8705) );
  XOR U8876 ( .A(n8706), .B(n8705), .Z(n8853) );
  NOR U8877 ( .A(n141), .B(n124), .Z(n8852) );
  IV U8878 ( .A(n8658), .Z(n8659) );
  NOR U8879 ( .A(n8660), .B(n8659), .Z(n8664) );
  NOR U8880 ( .A(n8662), .B(n8661), .Z(n8663) );
  NOR U8881 ( .A(n8664), .B(n8663), .Z(n8850) );
  XOR U8882 ( .A(n8852), .B(n8850), .Z(n8855) );
  XOR U8883 ( .A(n8853), .B(n8855), .Z(n8696) );
  XOR U8884 ( .A(n8697), .B(n8696), .Z(n8665) );
  IV U8885 ( .A(n8665), .Z(n8698) );
  XOR U8886 ( .A(n8699), .B(n8698), .Z(n8691) );
  NOR U8887 ( .A(n145), .B(n121), .Z(n8689) );
  XOR U8888 ( .A(n8691), .B(n8689), .Z(n8692) );
  XOR U8889 ( .A(n8693), .B(n8692), .Z(n8681) );
  XOR U8890 ( .A(n8682), .B(n8681), .Z(n8666) );
  IV U8891 ( .A(n8666), .Z(n8683) );
  XOR U8892 ( .A(n8684), .B(n8683), .Z(n8674) );
  NOR U8893 ( .A(n148), .B(n43), .Z(n8672) );
  XOR U8894 ( .A(n8674), .B(n8672), .Z(n8677) );
  XOR U8895 ( .A(n8675), .B(n8677), .Z(n8863) );
  XOR U8896 ( .A(n8861), .B(n8863), .Z(n8864) );
  XOR U8897 ( .A(n8865), .B(n8864), .Z(n10862) );
  IV U8898 ( .A(n10862), .Z(n8669) );
  XOR U8899 ( .A(n8668), .B(n8667), .Z(n10861) );
  NOR U8900 ( .A(n8669), .B(n10861), .Z(n8670) );
  NOR U8901 ( .A(n8671), .B(n8670), .Z(n8870) );
  IV U8902 ( .A(n8672), .Z(n8673) );
  NOR U8903 ( .A(n8674), .B(n8673), .Z(n8679) );
  IV U8904 ( .A(n8675), .Z(n8676) );
  NOR U8905 ( .A(n8677), .B(n8676), .Z(n8678) );
  NOR U8906 ( .A(n8679), .B(n8678), .Z(n8680) );
  IV U8907 ( .A(n8680), .Z(n8887) );
  NOR U8908 ( .A(n150), .B(n43), .Z(n8885) );
  NOR U8909 ( .A(n8682), .B(n8681), .Z(n8686) );
  NOR U8910 ( .A(n8684), .B(n8683), .Z(n8685) );
  NOR U8911 ( .A(n8686), .B(n8685), .Z(n8687) );
  IV U8912 ( .A(n8687), .Z(n8894) );
  NOR U8913 ( .A(n148), .B(n118), .Z(n8688) );
  IV U8914 ( .A(n8688), .Z(n8891) );
  IV U8915 ( .A(n8689), .Z(n8690) );
  NOR U8916 ( .A(n8691), .B(n8690), .Z(n8695) );
  NOR U8917 ( .A(n8693), .B(n8692), .Z(n8694) );
  NOR U8918 ( .A(n8695), .B(n8694), .Z(n8901) );
  NOR U8919 ( .A(n8697), .B(n8696), .Z(n8701) );
  NOR U8920 ( .A(n8699), .B(n8698), .Z(n8700) );
  NOR U8921 ( .A(n8701), .B(n8700), .Z(n8907) );
  NOR U8922 ( .A(n145), .B(n122), .Z(n8905) );
  IV U8923 ( .A(n8905), .Z(n8859) );
  IV U8924 ( .A(n8702), .Z(n8703) );
  NOR U8925 ( .A(n8704), .B(n8703), .Z(n8708) );
  NOR U8926 ( .A(n8706), .B(n8705), .Z(n8707) );
  NOR U8927 ( .A(n8708), .B(n8707), .Z(n8920) );
  NOR U8928 ( .A(n141), .B(n127), .Z(n8918) );
  IV U8929 ( .A(n8918), .Z(n8849) );
  IV U8930 ( .A(n8709), .Z(n8710) );
  NOR U8931 ( .A(n8711), .B(n8710), .Z(n8715) );
  NOR U8932 ( .A(n8713), .B(n8712), .Z(n8714) );
  NOR U8933 ( .A(n8715), .B(n8714), .Z(n8716) );
  IV U8934 ( .A(n8716), .Z(n9060) );
  NOR U8935 ( .A(n8718), .B(n8717), .Z(n8723) );
  IV U8936 ( .A(n8719), .Z(n8720) );
  NOR U8937 ( .A(n8721), .B(n8720), .Z(n8722) );
  NOR U8938 ( .A(n8723), .B(n8722), .Z(n8926) );
  NOR U8939 ( .A(n137), .B(n130), .Z(n8924) );
  IV U8940 ( .A(n8924), .Z(n8848) );
  NOR U8941 ( .A(n8725), .B(n8724), .Z(n8731) );
  IV U8942 ( .A(n8726), .Z(n8729) );
  IV U8943 ( .A(n8727), .Z(n8728) );
  NOR U8944 ( .A(n8729), .B(n8728), .Z(n8730) );
  NOR U8945 ( .A(n8731), .B(n8730), .Z(n8929) );
  IV U8946 ( .A(n8929), .Z(n8846) );
  IV U8947 ( .A(n8732), .Z(n8733) );
  NOR U8948 ( .A(n8734), .B(n8733), .Z(n8738) );
  NOR U8949 ( .A(n8736), .B(n8735), .Z(n8737) );
  NOR U8950 ( .A(n8738), .B(n8737), .Z(n8938) );
  NOR U8951 ( .A(n133), .B(n134), .Z(n8936) );
  IV U8952 ( .A(n8936), .Z(n8845) );
  IV U8953 ( .A(n8739), .Z(n8741) );
  NOR U8954 ( .A(n8741), .B(n8740), .Z(n8745) );
  NOR U8955 ( .A(n8743), .B(n8742), .Z(n8744) );
  NOR U8956 ( .A(n8745), .B(n8744), .Z(n8746) );
  IV U8957 ( .A(n8746), .Z(n8943) );
  NOR U8958 ( .A(n131), .B(n136), .Z(n8941) );
  XOR U8959 ( .A(n8943), .B(n8941), .Z(n8944) );
  NOR U8960 ( .A(n8748), .B(n8747), .Z(n8753) );
  IV U8961 ( .A(n8749), .Z(n8750) );
  NOR U8962 ( .A(n8751), .B(n8750), .Z(n8752) );
  NOR U8963 ( .A(n8753), .B(n8752), .Z(n8952) );
  NOR U8964 ( .A(n128), .B(n138), .Z(n8950) );
  NOR U8965 ( .A(n8755), .B(n8754), .Z(n8759) );
  NOR U8966 ( .A(n8757), .B(n8756), .Z(n8758) );
  NOR U8967 ( .A(n8759), .B(n8758), .Z(n8967) );
  NOR U8968 ( .A(n125), .B(n142), .Z(n8964) );
  NOR U8969 ( .A(n8761), .B(n8760), .Z(n8765) );
  NOR U8970 ( .A(n8763), .B(n8762), .Z(n8764) );
  NOR U8971 ( .A(n8765), .B(n8764), .Z(n8973) );
  NOR U8972 ( .A(n120), .B(n146), .Z(n8971) );
  NOR U8973 ( .A(n8767), .B(n8766), .Z(n8771) );
  NOR U8974 ( .A(n8769), .B(n8768), .Z(n8770) );
  NOR U8975 ( .A(n8771), .B(n8770), .Z(n8986) );
  NOR U8976 ( .A(n79), .B(n151), .Z(n8984) );
  NOR U8977 ( .A(n8773), .B(n8772), .Z(n8777) );
  NOR U8978 ( .A(n8775), .B(n8774), .Z(n8776) );
  NOR U8979 ( .A(n8777), .B(n8776), .Z(n8999) );
  NOR U8980 ( .A(n80), .B(n154), .Z(n8997) );
  IV U8981 ( .A(n8778), .Z(n8779) );
  NOR U8982 ( .A(n8780), .B(n8779), .Z(n8784) );
  NOR U8983 ( .A(n8782), .B(n8781), .Z(n8783) );
  NOR U8984 ( .A(n8784), .B(n8783), .Z(n9006) );
  NOR U8985 ( .A(n8786), .B(n8785), .Z(n8790) );
  NOR U8986 ( .A(n8788), .B(n8787), .Z(n8789) );
  NOR U8987 ( .A(n8790), .B(n8789), .Z(n9012) );
  NOR U8988 ( .A(n81), .B(n159), .Z(n9010) );
  IV U8989 ( .A(n8791), .Z(n8792) );
  NOR U8990 ( .A(n8793), .B(n8792), .Z(n8797) );
  NOR U8991 ( .A(n8795), .B(n8794), .Z(n8796) );
  NOR U8992 ( .A(n8797), .B(n8796), .Z(n9019) );
  NOR U8993 ( .A(n8799), .B(n8798), .Z(n8803) );
  NOR U8994 ( .A(n8801), .B(n8800), .Z(n8802) );
  NOR U8995 ( .A(n8803), .B(n8802), .Z(n9025) );
  NOR U8996 ( .A(n82), .B(n162), .Z(n9023) );
  IV U8997 ( .A(n9023), .Z(n8812) );
  IV U8998 ( .A(n8804), .Z(n8805) );
  NOR U8999 ( .A(n8806), .B(n8805), .Z(n8810) );
  NOR U9000 ( .A(n8808), .B(n8807), .Z(n8809) );
  NOR U9001 ( .A(n8810), .B(n8809), .Z(n9030) );
  NOR U9002 ( .A(n164), .B(n114), .Z(n9028) );
  XOR U9003 ( .A(n9030), .B(n9028), .Z(n9032) );
  NOR U9004 ( .A(n166), .B(n83), .Z(n8811) );
  IV U9005 ( .A(n8811), .Z(n9031) );
  XOR U9006 ( .A(n9032), .B(n9031), .Z(n9022) );
  XOR U9007 ( .A(n8812), .B(n9022), .Z(n9024) );
  XOR U9008 ( .A(n9025), .B(n9024), .Z(n9017) );
  NOR U9009 ( .A(n115), .B(n160), .Z(n9015) );
  XOR U9010 ( .A(n9017), .B(n9015), .Z(n9018) );
  XOR U9011 ( .A(n9019), .B(n9018), .Z(n9009) );
  XOR U9012 ( .A(n9010), .B(n9009), .Z(n8813) );
  IV U9013 ( .A(n8813), .Z(n9011) );
  XOR U9014 ( .A(n9012), .B(n9011), .Z(n9004) );
  NOR U9015 ( .A(n116), .B(n157), .Z(n9002) );
  XOR U9016 ( .A(n9004), .B(n9002), .Z(n9005) );
  XOR U9017 ( .A(n9006), .B(n9005), .Z(n8996) );
  XOR U9018 ( .A(n8997), .B(n8996), .Z(n8814) );
  IV U9019 ( .A(n8814), .Z(n8998) );
  XOR U9020 ( .A(n8999), .B(n8998), .Z(n8993) );
  IV U9021 ( .A(n8815), .Z(n8816) );
  NOR U9022 ( .A(n8817), .B(n8816), .Z(n8821) );
  NOR U9023 ( .A(n8819), .B(n8818), .Z(n8820) );
  NOR U9024 ( .A(n8821), .B(n8820), .Z(n8991) );
  NOR U9025 ( .A(n117), .B(n152), .Z(n8989) );
  XOR U9026 ( .A(n8991), .B(n8989), .Z(n8992) );
  XOR U9027 ( .A(n8993), .B(n8992), .Z(n8983) );
  XOR U9028 ( .A(n8984), .B(n8983), .Z(n8822) );
  IV U9029 ( .A(n8822), .Z(n8985) );
  XOR U9030 ( .A(n8986), .B(n8985), .Z(n8980) );
  IV U9031 ( .A(n8823), .Z(n8824) );
  NOR U9032 ( .A(n8825), .B(n8824), .Z(n8829) );
  NOR U9033 ( .A(n8827), .B(n8826), .Z(n8828) );
  NOR U9034 ( .A(n8829), .B(n8828), .Z(n8978) );
  NOR U9035 ( .A(n119), .B(n149), .Z(n8976) );
  XOR U9036 ( .A(n8978), .B(n8976), .Z(n8979) );
  XOR U9037 ( .A(n8980), .B(n8979), .Z(n8970) );
  XOR U9038 ( .A(n8971), .B(n8970), .Z(n8830) );
  IV U9039 ( .A(n8830), .Z(n8972) );
  XOR U9040 ( .A(n8973), .B(n8972), .Z(n9047) );
  IV U9041 ( .A(n8831), .Z(n8832) );
  NOR U9042 ( .A(n8833), .B(n8832), .Z(n8837) );
  NOR U9043 ( .A(n8835), .B(n8834), .Z(n8836) );
  NOR U9044 ( .A(n8837), .B(n8836), .Z(n9045) );
  NOR U9045 ( .A(n123), .B(n144), .Z(n9043) );
  XOR U9046 ( .A(n9045), .B(n9043), .Z(n9046) );
  XOR U9047 ( .A(n9047), .B(n9046), .Z(n8963) );
  XOR U9048 ( .A(n8964), .B(n8963), .Z(n8965) );
  XOR U9049 ( .A(n8967), .B(n8965), .Z(n8958) );
  NOR U9050 ( .A(n126), .B(n140), .Z(n8957) );
  IV U9051 ( .A(n8838), .Z(n8839) );
  NOR U9052 ( .A(n8840), .B(n8839), .Z(n8844) );
  NOR U9053 ( .A(n8842), .B(n8841), .Z(n8843) );
  NOR U9054 ( .A(n8844), .B(n8843), .Z(n8955) );
  XOR U9055 ( .A(n8957), .B(n8955), .Z(n8959) );
  XOR U9056 ( .A(n8958), .B(n8959), .Z(n8948) );
  XOR U9057 ( .A(n8950), .B(n8948), .Z(n8951) );
  XOR U9058 ( .A(n8952), .B(n8951), .Z(n8945) );
  XOR U9059 ( .A(n8944), .B(n8945), .Z(n8935) );
  XOR U9060 ( .A(n8845), .B(n8935), .Z(n8937) );
  XOR U9061 ( .A(n8938), .B(n8937), .Z(n8930) );
  XOR U9062 ( .A(n8846), .B(n8930), .Z(n8932) );
  NOR U9063 ( .A(n135), .B(n132), .Z(n8847) );
  IV U9064 ( .A(n8847), .Z(n8931) );
  XOR U9065 ( .A(n8932), .B(n8931), .Z(n8923) );
  XOR U9066 ( .A(n8848), .B(n8923), .Z(n8925) );
  XOR U9067 ( .A(n8926), .B(n8925), .Z(n9058) );
  NOR U9068 ( .A(n139), .B(n129), .Z(n9056) );
  XOR U9069 ( .A(n9058), .B(n9056), .Z(n9059) );
  XOR U9070 ( .A(n9060), .B(n9059), .Z(n8917) );
  XOR U9071 ( .A(n8849), .B(n8917), .Z(n8919) );
  XOR U9072 ( .A(n8920), .B(n8919), .Z(n8912) );
  IV U9073 ( .A(n8850), .Z(n8851) );
  NOR U9074 ( .A(n8852), .B(n8851), .Z(n8857) );
  IV U9075 ( .A(n8853), .Z(n8854) );
  NOR U9076 ( .A(n8855), .B(n8854), .Z(n8856) );
  NOR U9077 ( .A(n8857), .B(n8856), .Z(n8910) );
  XOR U9078 ( .A(n8912), .B(n8910), .Z(n8914) );
  NOR U9079 ( .A(n143), .B(n124), .Z(n8858) );
  IV U9080 ( .A(n8858), .Z(n8913) );
  XOR U9081 ( .A(n8914), .B(n8913), .Z(n8904) );
  XOR U9082 ( .A(n8859), .B(n8904), .Z(n8906) );
  XOR U9083 ( .A(n8907), .B(n8906), .Z(n8899) );
  NOR U9084 ( .A(n147), .B(n121), .Z(n8897) );
  XOR U9085 ( .A(n8899), .B(n8897), .Z(n8900) );
  XOR U9086 ( .A(n8901), .B(n8900), .Z(n8890) );
  XOR U9087 ( .A(n8891), .B(n8890), .Z(n8893) );
  XOR U9088 ( .A(n8894), .B(n8893), .Z(n8884) );
  XOR U9089 ( .A(n8885), .B(n8884), .Z(n8860) );
  IV U9090 ( .A(n8860), .Z(n8886) );
  XOR U9091 ( .A(n8887), .B(n8886), .Z(n8881) );
  IV U9092 ( .A(n8861), .Z(n8862) );
  NOR U9093 ( .A(n8863), .B(n8862), .Z(n8867) );
  NOR U9094 ( .A(n8865), .B(n8864), .Z(n8866) );
  NOR U9095 ( .A(n8867), .B(n8866), .Z(n8879) );
  NOR U9096 ( .A(n153), .B(n42), .Z(n8877) );
  XOR U9097 ( .A(n8879), .B(n8877), .Z(n8880) );
  XOR U9098 ( .A(n8881), .B(n8880), .Z(n8869) );
  IV U9099 ( .A(n8869), .Z(n8868) );
  NOR U9100 ( .A(n8870), .B(n8868), .Z(n8873) );
  XOR U9101 ( .A(n8870), .B(n8869), .Z(n10415) );
  NOR U9102 ( .A(n155), .B(n44), .Z(n10416) );
  IV U9103 ( .A(n10416), .Z(n8871) );
  NOR U9104 ( .A(n10415), .B(n8871), .Z(n8872) );
  NOR U9105 ( .A(n8873), .B(n8872), .Z(n8876) );
  NOR U9106 ( .A(n156), .B(n44), .Z(n8875) );
  IV U9107 ( .A(n8875), .Z(n8874) );
  NOR U9108 ( .A(n8876), .B(n8874), .Z(n9071) );
  XOR U9109 ( .A(n8876), .B(n8875), .Z(n10876) );
  IV U9110 ( .A(n8877), .Z(n8878) );
  NOR U9111 ( .A(n8879), .B(n8878), .Z(n8883) );
  NOR U9112 ( .A(n8881), .B(n8880), .Z(n8882) );
  NOR U9113 ( .A(n8883), .B(n8882), .Z(n9079) );
  NOR U9114 ( .A(n8885), .B(n8884), .Z(n8889) );
  NOR U9115 ( .A(n8887), .B(n8886), .Z(n8888) );
  NOR U9116 ( .A(n8889), .B(n8888), .Z(n9085) );
  NOR U9117 ( .A(n153), .B(n43), .Z(n9083) );
  IV U9118 ( .A(n8890), .Z(n8892) );
  NOR U9119 ( .A(n8892), .B(n8891), .Z(n8896) );
  NOR U9120 ( .A(n8894), .B(n8893), .Z(n8895) );
  NOR U9121 ( .A(n8896), .B(n8895), .Z(n9092) );
  NOR U9122 ( .A(n150), .B(n118), .Z(n9088) );
  IV U9123 ( .A(n8897), .Z(n8898) );
  NOR U9124 ( .A(n8899), .B(n8898), .Z(n8903) );
  NOR U9125 ( .A(n8901), .B(n8900), .Z(n8902) );
  NOR U9126 ( .A(n8903), .B(n8902), .Z(n9099) );
  IV U9127 ( .A(n9099), .Z(n9067) );
  NOR U9128 ( .A(n8905), .B(n8904), .Z(n8909) );
  NOR U9129 ( .A(n8907), .B(n8906), .Z(n8908) );
  NOR U9130 ( .A(n8909), .B(n8908), .Z(n9105) );
  NOR U9131 ( .A(n147), .B(n122), .Z(n9103) );
  IV U9132 ( .A(n9103), .Z(n9066) );
  IV U9133 ( .A(n8910), .Z(n8911) );
  NOR U9134 ( .A(n8912), .B(n8911), .Z(n8916) );
  NOR U9135 ( .A(n8914), .B(n8913), .Z(n8915) );
  NOR U9136 ( .A(n8916), .B(n8915), .Z(n9108) );
  IV U9137 ( .A(n9108), .Z(n9064) );
  NOR U9138 ( .A(n8918), .B(n8917), .Z(n8922) );
  NOR U9139 ( .A(n8920), .B(n8919), .Z(n8921) );
  NOR U9140 ( .A(n8922), .B(n8921), .Z(n9117) );
  NOR U9141 ( .A(n143), .B(n127), .Z(n9115) );
  IV U9142 ( .A(n9115), .Z(n9063) );
  NOR U9143 ( .A(n8924), .B(n8923), .Z(n8928) );
  NOR U9144 ( .A(n8926), .B(n8925), .Z(n8927) );
  NOR U9145 ( .A(n8928), .B(n8927), .Z(n9123) );
  NOR U9146 ( .A(n139), .B(n130), .Z(n9121) );
  IV U9147 ( .A(n9121), .Z(n9055) );
  NOR U9148 ( .A(n8930), .B(n8929), .Z(n8934) );
  NOR U9149 ( .A(n8932), .B(n8931), .Z(n8933) );
  NOR U9150 ( .A(n8934), .B(n8933), .Z(n9126) );
  IV U9151 ( .A(n9126), .Z(n9053) );
  NOR U9152 ( .A(n8936), .B(n8935), .Z(n8940) );
  NOR U9153 ( .A(n8938), .B(n8937), .Z(n8939) );
  NOR U9154 ( .A(n8940), .B(n8939), .Z(n9135) );
  NOR U9155 ( .A(n135), .B(n134), .Z(n9133) );
  IV U9156 ( .A(n9133), .Z(n9052) );
  IV U9157 ( .A(n8941), .Z(n8942) );
  NOR U9158 ( .A(n8943), .B(n8942), .Z(n8947) );
  NOR U9159 ( .A(n8945), .B(n8944), .Z(n8946) );
  NOR U9160 ( .A(n8947), .B(n8946), .Z(n9142) );
  IV U9161 ( .A(n8948), .Z(n8949) );
  NOR U9162 ( .A(n8950), .B(n8949), .Z(n8954) );
  NOR U9163 ( .A(n8952), .B(n8951), .Z(n8953) );
  NOR U9164 ( .A(n8954), .B(n8953), .Z(n9148) );
  NOR U9165 ( .A(n131), .B(n138), .Z(n9146) );
  IV U9166 ( .A(n9146), .Z(n9051) );
  IV U9167 ( .A(n8955), .Z(n8956) );
  NOR U9168 ( .A(n8957), .B(n8956), .Z(n8961) );
  NOR U9169 ( .A(n8959), .B(n8958), .Z(n8960) );
  NOR U9170 ( .A(n8961), .B(n8960), .Z(n8962) );
  IV U9171 ( .A(n8962), .Z(n9239) );
  NOR U9172 ( .A(n8964), .B(n8963), .Z(n8969) );
  IV U9173 ( .A(n8965), .Z(n8966) );
  NOR U9174 ( .A(n8967), .B(n8966), .Z(n8968) );
  NOR U9175 ( .A(n8969), .B(n8968), .Z(n9154) );
  NOR U9176 ( .A(n126), .B(n142), .Z(n9152) );
  NOR U9177 ( .A(n8971), .B(n8970), .Z(n8975) );
  NOR U9178 ( .A(n8973), .B(n8972), .Z(n8974) );
  NOR U9179 ( .A(n8975), .B(n8974), .Z(n9160) );
  NOR U9180 ( .A(n123), .B(n146), .Z(n9158) );
  IV U9181 ( .A(n8976), .Z(n8977) );
  NOR U9182 ( .A(n8978), .B(n8977), .Z(n8982) );
  NOR U9183 ( .A(n8980), .B(n8979), .Z(n8981) );
  NOR U9184 ( .A(n8982), .B(n8981), .Z(n9223) );
  NOR U9185 ( .A(n8984), .B(n8983), .Z(n8988) );
  NOR U9186 ( .A(n8986), .B(n8985), .Z(n8987) );
  NOR U9187 ( .A(n8988), .B(n8987), .Z(n9166) );
  NOR U9188 ( .A(n119), .B(n151), .Z(n9164) );
  IV U9189 ( .A(n9164), .Z(n9041) );
  IV U9190 ( .A(n8989), .Z(n8990) );
  NOR U9191 ( .A(n8991), .B(n8990), .Z(n8995) );
  NOR U9192 ( .A(n8993), .B(n8992), .Z(n8994) );
  NOR U9193 ( .A(n8995), .B(n8994), .Z(n9169) );
  IV U9194 ( .A(n9169), .Z(n9039) );
  NOR U9195 ( .A(n8997), .B(n8996), .Z(n9001) );
  NOR U9196 ( .A(n8999), .B(n8998), .Z(n9000) );
  NOR U9197 ( .A(n9001), .B(n9000), .Z(n9178) );
  NOR U9198 ( .A(n117), .B(n154), .Z(n9176) );
  IV U9199 ( .A(n9176), .Z(n9038) );
  IV U9200 ( .A(n9002), .Z(n9003) );
  NOR U9201 ( .A(n9004), .B(n9003), .Z(n9008) );
  NOR U9202 ( .A(n9006), .B(n9005), .Z(n9007) );
  NOR U9203 ( .A(n9008), .B(n9007), .Z(n9185) );
  NOR U9204 ( .A(n9010), .B(n9009), .Z(n9014) );
  NOR U9205 ( .A(n9012), .B(n9011), .Z(n9013) );
  NOR U9206 ( .A(n9014), .B(n9013), .Z(n9191) );
  NOR U9207 ( .A(n116), .B(n159), .Z(n9189) );
  IV U9208 ( .A(n9015), .Z(n9016) );
  NOR U9209 ( .A(n9017), .B(n9016), .Z(n9021) );
  NOR U9210 ( .A(n9019), .B(n9018), .Z(n9020) );
  NOR U9211 ( .A(n9021), .B(n9020), .Z(n9213) );
  NOR U9212 ( .A(n9023), .B(n9022), .Z(n9027) );
  NOR U9213 ( .A(n9025), .B(n9024), .Z(n9026) );
  NOR U9214 ( .A(n9027), .B(n9026), .Z(n9197) );
  NOR U9215 ( .A(n115), .B(n162), .Z(n9195) );
  IV U9216 ( .A(n9195), .Z(n9036) );
  IV U9217 ( .A(n9028), .Z(n9029) );
  NOR U9218 ( .A(n9030), .B(n9029), .Z(n9034) );
  NOR U9219 ( .A(n9032), .B(n9031), .Z(n9033) );
  NOR U9220 ( .A(n9034), .B(n9033), .Z(n9202) );
  NOR U9221 ( .A(n164), .B(n82), .Z(n9200) );
  XOR U9222 ( .A(n9202), .B(n9200), .Z(n9204) );
  NOR U9223 ( .A(n166), .B(n114), .Z(n9035) );
  IV U9224 ( .A(n9035), .Z(n9203) );
  XOR U9225 ( .A(n9204), .B(n9203), .Z(n9194) );
  XOR U9226 ( .A(n9036), .B(n9194), .Z(n9196) );
  XOR U9227 ( .A(n9197), .B(n9196), .Z(n9211) );
  NOR U9228 ( .A(n81), .B(n160), .Z(n9209) );
  XOR U9229 ( .A(n9211), .B(n9209), .Z(n9212) );
  XOR U9230 ( .A(n9213), .B(n9212), .Z(n9188) );
  XOR U9231 ( .A(n9189), .B(n9188), .Z(n9037) );
  IV U9232 ( .A(n9037), .Z(n9190) );
  XOR U9233 ( .A(n9191), .B(n9190), .Z(n9183) );
  NOR U9234 ( .A(n80), .B(n157), .Z(n9181) );
  XOR U9235 ( .A(n9183), .B(n9181), .Z(n9184) );
  XOR U9236 ( .A(n9185), .B(n9184), .Z(n9175) );
  XOR U9237 ( .A(n9038), .B(n9175), .Z(n9177) );
  XOR U9238 ( .A(n9178), .B(n9177), .Z(n9170) );
  XOR U9239 ( .A(n9039), .B(n9170), .Z(n9172) );
  NOR U9240 ( .A(n79), .B(n152), .Z(n9040) );
  IV U9241 ( .A(n9040), .Z(n9171) );
  XOR U9242 ( .A(n9172), .B(n9171), .Z(n9163) );
  XOR U9243 ( .A(n9041), .B(n9163), .Z(n9165) );
  XOR U9244 ( .A(n9166), .B(n9165), .Z(n9221) );
  NOR U9245 ( .A(n120), .B(n149), .Z(n9219) );
  XOR U9246 ( .A(n9221), .B(n9219), .Z(n9222) );
  XOR U9247 ( .A(n9223), .B(n9222), .Z(n9157) );
  XOR U9248 ( .A(n9158), .B(n9157), .Z(n9042) );
  IV U9249 ( .A(n9042), .Z(n9159) );
  XOR U9250 ( .A(n9160), .B(n9159), .Z(n9231) );
  IV U9251 ( .A(n9043), .Z(n9044) );
  NOR U9252 ( .A(n9045), .B(n9044), .Z(n9049) );
  NOR U9253 ( .A(n9047), .B(n9046), .Z(n9048) );
  NOR U9254 ( .A(n9049), .B(n9048), .Z(n9229) );
  NOR U9255 ( .A(n125), .B(n144), .Z(n9227) );
  XOR U9256 ( .A(n9229), .B(n9227), .Z(n9230) );
  XOR U9257 ( .A(n9231), .B(n9230), .Z(n9151) );
  XOR U9258 ( .A(n9152), .B(n9151), .Z(n9050) );
  IV U9259 ( .A(n9050), .Z(n9153) );
  XOR U9260 ( .A(n9154), .B(n9153), .Z(n9237) );
  NOR U9261 ( .A(n128), .B(n140), .Z(n9235) );
  XOR U9262 ( .A(n9237), .B(n9235), .Z(n9238) );
  XOR U9263 ( .A(n9239), .B(n9238), .Z(n9145) );
  XOR U9264 ( .A(n9051), .B(n9145), .Z(n9147) );
  XOR U9265 ( .A(n9148), .B(n9147), .Z(n9140) );
  NOR U9266 ( .A(n133), .B(n136), .Z(n9138) );
  XOR U9267 ( .A(n9140), .B(n9138), .Z(n9141) );
  XOR U9268 ( .A(n9142), .B(n9141), .Z(n9132) );
  XOR U9269 ( .A(n9052), .B(n9132), .Z(n9134) );
  XOR U9270 ( .A(n9135), .B(n9134), .Z(n9127) );
  XOR U9271 ( .A(n9053), .B(n9127), .Z(n9129) );
  NOR U9272 ( .A(n137), .B(n132), .Z(n9054) );
  IV U9273 ( .A(n9054), .Z(n9128) );
  XOR U9274 ( .A(n9129), .B(n9128), .Z(n9120) );
  XOR U9275 ( .A(n9055), .B(n9120), .Z(n9122) );
  XOR U9276 ( .A(n9123), .B(n9122), .Z(n9251) );
  IV U9277 ( .A(n9056), .Z(n9057) );
  NOR U9278 ( .A(n9058), .B(n9057), .Z(n9062) );
  NOR U9279 ( .A(n9060), .B(n9059), .Z(n9061) );
  NOR U9280 ( .A(n9062), .B(n9061), .Z(n9249) );
  NOR U9281 ( .A(n141), .B(n129), .Z(n9247) );
  XOR U9282 ( .A(n9249), .B(n9247), .Z(n9250) );
  XOR U9283 ( .A(n9251), .B(n9250), .Z(n9114) );
  XOR U9284 ( .A(n9063), .B(n9114), .Z(n9116) );
  XOR U9285 ( .A(n9117), .B(n9116), .Z(n9109) );
  XOR U9286 ( .A(n9064), .B(n9109), .Z(n9111) );
  NOR U9287 ( .A(n145), .B(n124), .Z(n9065) );
  IV U9288 ( .A(n9065), .Z(n9110) );
  XOR U9289 ( .A(n9111), .B(n9110), .Z(n9102) );
  XOR U9290 ( .A(n9066), .B(n9102), .Z(n9104) );
  XOR U9291 ( .A(n9105), .B(n9104), .Z(n9097) );
  NOR U9292 ( .A(n148), .B(n121), .Z(n9095) );
  XOR U9293 ( .A(n9097), .B(n9095), .Z(n9098) );
  XOR U9294 ( .A(n9067), .B(n9098), .Z(n9090) );
  XOR U9295 ( .A(n9088), .B(n9090), .Z(n9091) );
  XOR U9296 ( .A(n9092), .B(n9091), .Z(n9082) );
  XOR U9297 ( .A(n9083), .B(n9082), .Z(n9068) );
  IV U9298 ( .A(n9068), .Z(n9084) );
  XOR U9299 ( .A(n9085), .B(n9084), .Z(n9077) );
  NOR U9300 ( .A(n155), .B(n42), .Z(n9075) );
  XOR U9301 ( .A(n9077), .B(n9075), .Z(n9078) );
  XOR U9302 ( .A(n9079), .B(n9078), .Z(n10877) );
  IV U9303 ( .A(n10877), .Z(n9069) );
  NOR U9304 ( .A(n10876), .B(n9069), .Z(n9070) );
  NOR U9305 ( .A(n9071), .B(n9070), .Z(n9074) );
  NOR U9306 ( .A(n158), .B(n44), .Z(n9073) );
  IV U9307 ( .A(n9073), .Z(n9072) );
  NOR U9308 ( .A(n9074), .B(n9072), .Z(n9258) );
  XOR U9309 ( .A(n9074), .B(n9073), .Z(n10880) );
  IV U9310 ( .A(n9075), .Z(n9076) );
  NOR U9311 ( .A(n9077), .B(n9076), .Z(n9081) );
  NOR U9312 ( .A(n9079), .B(n9078), .Z(n9080) );
  NOR U9313 ( .A(n9081), .B(n9080), .Z(n9263) );
  NOR U9314 ( .A(n156), .B(n42), .Z(n9259) );
  NOR U9315 ( .A(n9083), .B(n9082), .Z(n9087) );
  NOR U9316 ( .A(n9085), .B(n9084), .Z(n9086) );
  NOR U9317 ( .A(n9087), .B(n9086), .Z(n9269) );
  NOR U9318 ( .A(n155), .B(n43), .Z(n9266) );
  IV U9319 ( .A(n9088), .Z(n9089) );
  NOR U9320 ( .A(n9090), .B(n9089), .Z(n9094) );
  NOR U9321 ( .A(n9092), .B(n9091), .Z(n9093) );
  NOR U9322 ( .A(n9094), .B(n9093), .Z(n9279) );
  IV U9323 ( .A(n9279), .Z(n9255) );
  NOR U9324 ( .A(n153), .B(n118), .Z(n9275) );
  IV U9325 ( .A(n9095), .Z(n9096) );
  NOR U9326 ( .A(n9097), .B(n9096), .Z(n9101) );
  NOR U9327 ( .A(n9099), .B(n9098), .Z(n9100) );
  NOR U9328 ( .A(n9101), .B(n9100), .Z(n9286) );
  IV U9329 ( .A(n9286), .Z(n9254) );
  NOR U9330 ( .A(n9103), .B(n9102), .Z(n9107) );
  NOR U9331 ( .A(n9105), .B(n9104), .Z(n9106) );
  NOR U9332 ( .A(n9107), .B(n9106), .Z(n9293) );
  NOR U9333 ( .A(n148), .B(n122), .Z(n9291) );
  NOR U9334 ( .A(n147), .B(n124), .Z(n9449) );
  NOR U9335 ( .A(n9109), .B(n9108), .Z(n9113) );
  NOR U9336 ( .A(n9111), .B(n9110), .Z(n9112) );
  NOR U9337 ( .A(n9113), .B(n9112), .Z(n9445) );
  NOR U9338 ( .A(n9115), .B(n9114), .Z(n9119) );
  NOR U9339 ( .A(n9117), .B(n9116), .Z(n9118) );
  NOR U9340 ( .A(n9119), .B(n9118), .Z(n9300) );
  NOR U9341 ( .A(n145), .B(n127), .Z(n9297) );
  NOR U9342 ( .A(n9121), .B(n9120), .Z(n9125) );
  NOR U9343 ( .A(n9123), .B(n9122), .Z(n9124) );
  NOR U9344 ( .A(n9125), .B(n9124), .Z(n9306) );
  NOR U9345 ( .A(n141), .B(n130), .Z(n9304) );
  IV U9346 ( .A(n9304), .Z(n9246) );
  NOR U9347 ( .A(n9127), .B(n9126), .Z(n9131) );
  NOR U9348 ( .A(n9129), .B(n9128), .Z(n9130) );
  NOR U9349 ( .A(n9131), .B(n9130), .Z(n9309) );
  IV U9350 ( .A(n9309), .Z(n9244) );
  NOR U9351 ( .A(n9133), .B(n9132), .Z(n9137) );
  NOR U9352 ( .A(n9135), .B(n9134), .Z(n9136) );
  NOR U9353 ( .A(n9137), .B(n9136), .Z(n9318) );
  NOR U9354 ( .A(n137), .B(n134), .Z(n9316) );
  IV U9355 ( .A(n9316), .Z(n9243) );
  IV U9356 ( .A(n9138), .Z(n9139) );
  NOR U9357 ( .A(n9140), .B(n9139), .Z(n9144) );
  NOR U9358 ( .A(n9142), .B(n9141), .Z(n9143) );
  NOR U9359 ( .A(n9144), .B(n9143), .Z(n9325) );
  NOR U9360 ( .A(n9146), .B(n9145), .Z(n9150) );
  NOR U9361 ( .A(n9148), .B(n9147), .Z(n9149) );
  NOR U9362 ( .A(n9150), .B(n9149), .Z(n9331) );
  NOR U9363 ( .A(n133), .B(n138), .Z(n9329) );
  NOR U9364 ( .A(n9152), .B(n9151), .Z(n9156) );
  NOR U9365 ( .A(n9154), .B(n9153), .Z(n9155) );
  NOR U9366 ( .A(n9156), .B(n9155), .Z(n9344) );
  NOR U9367 ( .A(n128), .B(n142), .Z(n9342) );
  NOR U9368 ( .A(n9158), .B(n9157), .Z(n9162) );
  NOR U9369 ( .A(n9160), .B(n9159), .Z(n9161) );
  NOR U9370 ( .A(n9162), .B(n9161), .Z(n9350) );
  NOR U9371 ( .A(n125), .B(n146), .Z(n9348) );
  NOR U9372 ( .A(n9164), .B(n9163), .Z(n9168) );
  NOR U9373 ( .A(n9166), .B(n9165), .Z(n9167) );
  NOR U9374 ( .A(n9168), .B(n9167), .Z(n9363) );
  NOR U9375 ( .A(n120), .B(n151), .Z(n9361) );
  NOR U9376 ( .A(n9170), .B(n9169), .Z(n9174) );
  NOR U9377 ( .A(n9172), .B(n9171), .Z(n9173) );
  NOR U9378 ( .A(n9174), .B(n9173), .Z(n9370) );
  NOR U9379 ( .A(n9176), .B(n9175), .Z(n9180) );
  NOR U9380 ( .A(n9178), .B(n9177), .Z(n9179) );
  NOR U9381 ( .A(n9180), .B(n9179), .Z(n9376) );
  NOR U9382 ( .A(n79), .B(n154), .Z(n9374) );
  IV U9383 ( .A(n9181), .Z(n9182) );
  NOR U9384 ( .A(n9183), .B(n9182), .Z(n9187) );
  NOR U9385 ( .A(n9185), .B(n9184), .Z(n9186) );
  NOR U9386 ( .A(n9187), .B(n9186), .Z(n9383) );
  NOR U9387 ( .A(n9189), .B(n9188), .Z(n9193) );
  NOR U9388 ( .A(n9191), .B(n9190), .Z(n9192) );
  NOR U9389 ( .A(n9193), .B(n9192), .Z(n9389) );
  NOR U9390 ( .A(n80), .B(n159), .Z(n9387) );
  NOR U9391 ( .A(n9195), .B(n9194), .Z(n9199) );
  NOR U9392 ( .A(n9197), .B(n9196), .Z(n9198) );
  NOR U9393 ( .A(n9199), .B(n9198), .Z(n9402) );
  NOR U9394 ( .A(n81), .B(n162), .Z(n9400) );
  IV U9395 ( .A(n9400), .Z(n9208) );
  IV U9396 ( .A(n9200), .Z(n9201) );
  NOR U9397 ( .A(n9202), .B(n9201), .Z(n9206) );
  NOR U9398 ( .A(n9204), .B(n9203), .Z(n9205) );
  NOR U9399 ( .A(n9206), .B(n9205), .Z(n9407) );
  NOR U9400 ( .A(n164), .B(n115), .Z(n9405) );
  XOR U9401 ( .A(n9407), .B(n9405), .Z(n9409) );
  NOR U9402 ( .A(n166), .B(n82), .Z(n9207) );
  IV U9403 ( .A(n9207), .Z(n9408) );
  XOR U9404 ( .A(n9409), .B(n9408), .Z(n9399) );
  XOR U9405 ( .A(n9208), .B(n9399), .Z(n9401) );
  XOR U9406 ( .A(n9402), .B(n9401), .Z(n9396) );
  IV U9407 ( .A(n9209), .Z(n9210) );
  NOR U9408 ( .A(n9211), .B(n9210), .Z(n9215) );
  NOR U9409 ( .A(n9213), .B(n9212), .Z(n9214) );
  NOR U9410 ( .A(n9215), .B(n9214), .Z(n9394) );
  NOR U9411 ( .A(n116), .B(n160), .Z(n9392) );
  XOR U9412 ( .A(n9394), .B(n9392), .Z(n9395) );
  XOR U9413 ( .A(n9396), .B(n9395), .Z(n9386) );
  XOR U9414 ( .A(n9387), .B(n9386), .Z(n9216) );
  IV U9415 ( .A(n9216), .Z(n9388) );
  XOR U9416 ( .A(n9389), .B(n9388), .Z(n9381) );
  NOR U9417 ( .A(n117), .B(n157), .Z(n9379) );
  XOR U9418 ( .A(n9381), .B(n9379), .Z(n9382) );
  XOR U9419 ( .A(n9383), .B(n9382), .Z(n9373) );
  XOR U9420 ( .A(n9374), .B(n9373), .Z(n9217) );
  IV U9421 ( .A(n9217), .Z(n9375) );
  XOR U9422 ( .A(n9376), .B(n9375), .Z(n9368) );
  NOR U9423 ( .A(n119), .B(n152), .Z(n9366) );
  XOR U9424 ( .A(n9368), .B(n9366), .Z(n9369) );
  XOR U9425 ( .A(n9370), .B(n9369), .Z(n9360) );
  XOR U9426 ( .A(n9361), .B(n9360), .Z(n9218) );
  IV U9427 ( .A(n9218), .Z(n9362) );
  XOR U9428 ( .A(n9363), .B(n9362), .Z(n9357) );
  IV U9429 ( .A(n9219), .Z(n9220) );
  NOR U9430 ( .A(n9221), .B(n9220), .Z(n9225) );
  NOR U9431 ( .A(n9223), .B(n9222), .Z(n9224) );
  NOR U9432 ( .A(n9225), .B(n9224), .Z(n9355) );
  NOR U9433 ( .A(n123), .B(n149), .Z(n9353) );
  XOR U9434 ( .A(n9355), .B(n9353), .Z(n9356) );
  XOR U9435 ( .A(n9357), .B(n9356), .Z(n9347) );
  XOR U9436 ( .A(n9348), .B(n9347), .Z(n9226) );
  IV U9437 ( .A(n9226), .Z(n9349) );
  XOR U9438 ( .A(n9350), .B(n9349), .Z(n9426) );
  IV U9439 ( .A(n9227), .Z(n9228) );
  NOR U9440 ( .A(n9229), .B(n9228), .Z(n9233) );
  NOR U9441 ( .A(n9231), .B(n9230), .Z(n9232) );
  NOR U9442 ( .A(n9233), .B(n9232), .Z(n9424) );
  NOR U9443 ( .A(n126), .B(n144), .Z(n9422) );
  XOR U9444 ( .A(n9424), .B(n9422), .Z(n9425) );
  XOR U9445 ( .A(n9426), .B(n9425), .Z(n9341) );
  XOR U9446 ( .A(n9342), .B(n9341), .Z(n9234) );
  IV U9447 ( .A(n9234), .Z(n9343) );
  XOR U9448 ( .A(n9344), .B(n9343), .Z(n9338) );
  IV U9449 ( .A(n9235), .Z(n9236) );
  NOR U9450 ( .A(n9237), .B(n9236), .Z(n9241) );
  NOR U9451 ( .A(n9239), .B(n9238), .Z(n9240) );
  NOR U9452 ( .A(n9241), .B(n9240), .Z(n9336) );
  NOR U9453 ( .A(n131), .B(n140), .Z(n9334) );
  XOR U9454 ( .A(n9336), .B(n9334), .Z(n9337) );
  XOR U9455 ( .A(n9338), .B(n9337), .Z(n9328) );
  XOR U9456 ( .A(n9329), .B(n9328), .Z(n9242) );
  IV U9457 ( .A(n9242), .Z(n9330) );
  XOR U9458 ( .A(n9331), .B(n9330), .Z(n9323) );
  NOR U9459 ( .A(n135), .B(n136), .Z(n9321) );
  XOR U9460 ( .A(n9323), .B(n9321), .Z(n9324) );
  XOR U9461 ( .A(n9325), .B(n9324), .Z(n9315) );
  XOR U9462 ( .A(n9243), .B(n9315), .Z(n9317) );
  XOR U9463 ( .A(n9318), .B(n9317), .Z(n9310) );
  XOR U9464 ( .A(n9244), .B(n9310), .Z(n9312) );
  NOR U9465 ( .A(n139), .B(n132), .Z(n9245) );
  IV U9466 ( .A(n9245), .Z(n9311) );
  XOR U9467 ( .A(n9312), .B(n9311), .Z(n9303) );
  XOR U9468 ( .A(n9246), .B(n9303), .Z(n9305) );
  XOR U9469 ( .A(n9306), .B(n9305), .Z(n9441) );
  IV U9470 ( .A(n9247), .Z(n9248) );
  NOR U9471 ( .A(n9249), .B(n9248), .Z(n9253) );
  NOR U9472 ( .A(n9251), .B(n9250), .Z(n9252) );
  NOR U9473 ( .A(n9253), .B(n9252), .Z(n9439) );
  NOR U9474 ( .A(n143), .B(n129), .Z(n9437) );
  XOR U9475 ( .A(n9439), .B(n9437), .Z(n9440) );
  XOR U9476 ( .A(n9441), .B(n9440), .Z(n9296) );
  XOR U9477 ( .A(n9297), .B(n9296), .Z(n9298) );
  XOR U9478 ( .A(n9300), .B(n9298), .Z(n9446) );
  XOR U9479 ( .A(n9445), .B(n9446), .Z(n9448) );
  XOR U9480 ( .A(n9449), .B(n9448), .Z(n9289) );
  XOR U9481 ( .A(n9291), .B(n9289), .Z(n9292) );
  XOR U9482 ( .A(n9293), .B(n9292), .Z(n9284) );
  NOR U9483 ( .A(n150), .B(n121), .Z(n9282) );
  XOR U9484 ( .A(n9284), .B(n9282), .Z(n9285) );
  XOR U9485 ( .A(n9254), .B(n9285), .Z(n9277) );
  XOR U9486 ( .A(n9275), .B(n9277), .Z(n9278) );
  XOR U9487 ( .A(n9255), .B(n9278), .Z(n9268) );
  XOR U9488 ( .A(n9266), .B(n9268), .Z(n9270) );
  XOR U9489 ( .A(n9269), .B(n9270), .Z(n9261) );
  XOR U9490 ( .A(n9259), .B(n9261), .Z(n9262) );
  XOR U9491 ( .A(n9263), .B(n9262), .Z(n10881) );
  IV U9492 ( .A(n10881), .Z(n9256) );
  NOR U9493 ( .A(n10880), .B(n9256), .Z(n9257) );
  NOR U9494 ( .A(n9258), .B(n9257), .Z(n9458) );
  IV U9495 ( .A(n9259), .Z(n9260) );
  NOR U9496 ( .A(n9261), .B(n9260), .Z(n9265) );
  NOR U9497 ( .A(n9263), .B(n9262), .Z(n9264) );
  NOR U9498 ( .A(n9265), .B(n9264), .Z(n9469) );
  IV U9499 ( .A(n9266), .Z(n9267) );
  NOR U9500 ( .A(n9268), .B(n9267), .Z(n9273) );
  IV U9501 ( .A(n9269), .Z(n9271) );
  NOR U9502 ( .A(n9271), .B(n9270), .Z(n9272) );
  NOR U9503 ( .A(n9273), .B(n9272), .Z(n9274) );
  IV U9504 ( .A(n9274), .Z(n9475) );
  NOR U9505 ( .A(n156), .B(n43), .Z(n9473) );
  IV U9506 ( .A(n9275), .Z(n9276) );
  NOR U9507 ( .A(n9277), .B(n9276), .Z(n9281) );
  NOR U9508 ( .A(n9279), .B(n9278), .Z(n9280) );
  NOR U9509 ( .A(n9281), .B(n9280), .Z(n9482) );
  NOR U9510 ( .A(n155), .B(n118), .Z(n9478) );
  IV U9511 ( .A(n9282), .Z(n9283) );
  NOR U9512 ( .A(n9284), .B(n9283), .Z(n9288) );
  NOR U9513 ( .A(n9286), .B(n9285), .Z(n9287) );
  NOR U9514 ( .A(n9288), .B(n9287), .Z(n9490) );
  IV U9515 ( .A(n9490), .Z(n9454) );
  IV U9516 ( .A(n9289), .Z(n9290) );
  NOR U9517 ( .A(n9291), .B(n9290), .Z(n9295) );
  NOR U9518 ( .A(n9293), .B(n9292), .Z(n9294) );
  NOR U9519 ( .A(n9295), .B(n9294), .Z(n9496) );
  NOR U9520 ( .A(n150), .B(n122), .Z(n9494) );
  IV U9521 ( .A(n9494), .Z(n9453) );
  NOR U9522 ( .A(n9297), .B(n9296), .Z(n9302) );
  IV U9523 ( .A(n9298), .Z(n9299) );
  NOR U9524 ( .A(n9300), .B(n9299), .Z(n9301) );
  NOR U9525 ( .A(n9302), .B(n9301), .Z(n9509) );
  NOR U9526 ( .A(n147), .B(n127), .Z(n9507) );
  NOR U9527 ( .A(n9304), .B(n9303), .Z(n9308) );
  NOR U9528 ( .A(n9306), .B(n9305), .Z(n9307) );
  NOR U9529 ( .A(n9308), .B(n9307), .Z(n9515) );
  NOR U9530 ( .A(n143), .B(n130), .Z(n9513) );
  IV U9531 ( .A(n9513), .Z(n9436) );
  NOR U9532 ( .A(n9310), .B(n9309), .Z(n9314) );
  NOR U9533 ( .A(n9312), .B(n9311), .Z(n9313) );
  NOR U9534 ( .A(n9314), .B(n9313), .Z(n9627) );
  IV U9535 ( .A(n9627), .Z(n9434) );
  NOR U9536 ( .A(n9316), .B(n9315), .Z(n9320) );
  NOR U9537 ( .A(n9318), .B(n9317), .Z(n9319) );
  NOR U9538 ( .A(n9320), .B(n9319), .Z(n9521) );
  NOR U9539 ( .A(n139), .B(n134), .Z(n9519) );
  IV U9540 ( .A(n9519), .Z(n9433) );
  IV U9541 ( .A(n9321), .Z(n9322) );
  NOR U9542 ( .A(n9323), .B(n9322), .Z(n9327) );
  NOR U9543 ( .A(n9325), .B(n9324), .Z(n9326) );
  NOR U9544 ( .A(n9327), .B(n9326), .Z(n9624) );
  NOR U9545 ( .A(n9329), .B(n9328), .Z(n9333) );
  NOR U9546 ( .A(n9331), .B(n9330), .Z(n9332) );
  NOR U9547 ( .A(n9333), .B(n9332), .Z(n9527) );
  NOR U9548 ( .A(n135), .B(n138), .Z(n9525) );
  IV U9549 ( .A(n9525), .Z(n9432) );
  IV U9550 ( .A(n9334), .Z(n9335) );
  NOR U9551 ( .A(n9336), .B(n9335), .Z(n9340) );
  NOR U9552 ( .A(n9338), .B(n9337), .Z(n9339) );
  NOR U9553 ( .A(n9340), .B(n9339), .Z(n9530) );
  IV U9554 ( .A(n9530), .Z(n9430) );
  NOR U9555 ( .A(n9342), .B(n9341), .Z(n9346) );
  NOR U9556 ( .A(n9344), .B(n9343), .Z(n9345) );
  NOR U9557 ( .A(n9346), .B(n9345), .Z(n9539) );
  NOR U9558 ( .A(n131), .B(n142), .Z(n9537) );
  IV U9559 ( .A(n9537), .Z(n9429) );
  NOR U9560 ( .A(n9348), .B(n9347), .Z(n9352) );
  NOR U9561 ( .A(n9350), .B(n9349), .Z(n9351) );
  NOR U9562 ( .A(n9352), .B(n9351), .Z(n9552) );
  NOR U9563 ( .A(n126), .B(n146), .Z(n9550) );
  IV U9564 ( .A(n9550), .Z(n9421) );
  IV U9565 ( .A(n9353), .Z(n9354) );
  NOR U9566 ( .A(n9355), .B(n9354), .Z(n9359) );
  NOR U9567 ( .A(n9357), .B(n9356), .Z(n9358) );
  NOR U9568 ( .A(n9359), .B(n9358), .Z(n9555) );
  IV U9569 ( .A(n9555), .Z(n9419) );
  NOR U9570 ( .A(n9361), .B(n9360), .Z(n9365) );
  NOR U9571 ( .A(n9363), .B(n9362), .Z(n9364) );
  NOR U9572 ( .A(n9365), .B(n9364), .Z(n9564) );
  NOR U9573 ( .A(n123), .B(n151), .Z(n9562) );
  IV U9574 ( .A(n9562), .Z(n9418) );
  IV U9575 ( .A(n9366), .Z(n9367) );
  NOR U9576 ( .A(n9368), .B(n9367), .Z(n9372) );
  NOR U9577 ( .A(n9370), .B(n9369), .Z(n9371) );
  NOR U9578 ( .A(n9372), .B(n9371), .Z(n9569) );
  NOR U9579 ( .A(n120), .B(n152), .Z(n9568) );
  NOR U9580 ( .A(n9374), .B(n9373), .Z(n9378) );
  NOR U9581 ( .A(n9376), .B(n9375), .Z(n9377) );
  NOR U9582 ( .A(n9378), .B(n9377), .Z(n9579) );
  NOR U9583 ( .A(n119), .B(n154), .Z(n9576) );
  IV U9584 ( .A(n9379), .Z(n9380) );
  NOR U9585 ( .A(n9381), .B(n9380), .Z(n9385) );
  NOR U9586 ( .A(n9383), .B(n9382), .Z(n9384) );
  NOR U9587 ( .A(n9385), .B(n9384), .Z(n9614) );
  NOR U9588 ( .A(n9387), .B(n9386), .Z(n9391) );
  NOR U9589 ( .A(n9389), .B(n9388), .Z(n9390) );
  NOR U9590 ( .A(n9391), .B(n9390), .Z(n9585) );
  NOR U9591 ( .A(n117), .B(n159), .Z(n9583) );
  IV U9592 ( .A(n9583), .Z(n9416) );
  IV U9593 ( .A(n9392), .Z(n9393) );
  NOR U9594 ( .A(n9394), .B(n9393), .Z(n9398) );
  NOR U9595 ( .A(n9396), .B(n9395), .Z(n9397) );
  NOR U9596 ( .A(n9398), .B(n9397), .Z(n9588) );
  IV U9597 ( .A(n9588), .Z(n9414) );
  NOR U9598 ( .A(n9400), .B(n9399), .Z(n9404) );
  NOR U9599 ( .A(n9402), .B(n9401), .Z(n9403) );
  NOR U9600 ( .A(n9404), .B(n9403), .Z(n9597) );
  NOR U9601 ( .A(n116), .B(n162), .Z(n9595) );
  IV U9602 ( .A(n9595), .Z(n9413) );
  IV U9603 ( .A(n9405), .Z(n9406) );
  NOR U9604 ( .A(n9407), .B(n9406), .Z(n9411) );
  NOR U9605 ( .A(n9409), .B(n9408), .Z(n9410) );
  NOR U9606 ( .A(n9411), .B(n9410), .Z(n9602) );
  NOR U9607 ( .A(n164), .B(n81), .Z(n9600) );
  XOR U9608 ( .A(n9602), .B(n9600), .Z(n9604) );
  NOR U9609 ( .A(n166), .B(n115), .Z(n9412) );
  IV U9610 ( .A(n9412), .Z(n9603) );
  XOR U9611 ( .A(n9604), .B(n9603), .Z(n9594) );
  XOR U9612 ( .A(n9413), .B(n9594), .Z(n9596) );
  XOR U9613 ( .A(n9597), .B(n9596), .Z(n9589) );
  XOR U9614 ( .A(n9414), .B(n9589), .Z(n9591) );
  NOR U9615 ( .A(n80), .B(n160), .Z(n9415) );
  IV U9616 ( .A(n9415), .Z(n9590) );
  XOR U9617 ( .A(n9591), .B(n9590), .Z(n9582) );
  XOR U9618 ( .A(n9416), .B(n9582), .Z(n9584) );
  XOR U9619 ( .A(n9585), .B(n9584), .Z(n9612) );
  NOR U9620 ( .A(n79), .B(n157), .Z(n9610) );
  XOR U9621 ( .A(n9612), .B(n9610), .Z(n9613) );
  XOR U9622 ( .A(n9614), .B(n9613), .Z(n9575) );
  XOR U9623 ( .A(n9576), .B(n9575), .Z(n9577) );
  XOR U9624 ( .A(n9579), .B(n9577), .Z(n9567) );
  XOR U9625 ( .A(n9568), .B(n9567), .Z(n9417) );
  IV U9626 ( .A(n9417), .Z(n9570) );
  XOR U9627 ( .A(n9569), .B(n9570), .Z(n9561) );
  XOR U9628 ( .A(n9418), .B(n9561), .Z(n9563) );
  XOR U9629 ( .A(n9564), .B(n9563), .Z(n9556) );
  XOR U9630 ( .A(n9419), .B(n9556), .Z(n9558) );
  NOR U9631 ( .A(n125), .B(n149), .Z(n9420) );
  IV U9632 ( .A(n9420), .Z(n9557) );
  XOR U9633 ( .A(n9558), .B(n9557), .Z(n9549) );
  XOR U9634 ( .A(n9421), .B(n9549), .Z(n9551) );
  XOR U9635 ( .A(n9552), .B(n9551), .Z(n9546) );
  IV U9636 ( .A(n9422), .Z(n9423) );
  NOR U9637 ( .A(n9424), .B(n9423), .Z(n9428) );
  NOR U9638 ( .A(n9426), .B(n9425), .Z(n9427) );
  NOR U9639 ( .A(n9428), .B(n9427), .Z(n9544) );
  NOR U9640 ( .A(n128), .B(n144), .Z(n9542) );
  XOR U9641 ( .A(n9544), .B(n9542), .Z(n9545) );
  XOR U9642 ( .A(n9546), .B(n9545), .Z(n9536) );
  XOR U9643 ( .A(n9429), .B(n9536), .Z(n9538) );
  XOR U9644 ( .A(n9539), .B(n9538), .Z(n9531) );
  XOR U9645 ( .A(n9430), .B(n9531), .Z(n9533) );
  NOR U9646 ( .A(n133), .B(n140), .Z(n9431) );
  IV U9647 ( .A(n9431), .Z(n9532) );
  XOR U9648 ( .A(n9533), .B(n9532), .Z(n9524) );
  XOR U9649 ( .A(n9432), .B(n9524), .Z(n9526) );
  XOR U9650 ( .A(n9527), .B(n9526), .Z(n9622) );
  NOR U9651 ( .A(n137), .B(n136), .Z(n9620) );
  XOR U9652 ( .A(n9622), .B(n9620), .Z(n9623) );
  XOR U9653 ( .A(n9624), .B(n9623), .Z(n9518) );
  XOR U9654 ( .A(n9433), .B(n9518), .Z(n9520) );
  XOR U9655 ( .A(n9521), .B(n9520), .Z(n9628) );
  XOR U9656 ( .A(n9434), .B(n9628), .Z(n9630) );
  NOR U9657 ( .A(n141), .B(n132), .Z(n9435) );
  IV U9658 ( .A(n9435), .Z(n9629) );
  XOR U9659 ( .A(n9630), .B(n9629), .Z(n9512) );
  XOR U9660 ( .A(n9436), .B(n9512), .Z(n9514) );
  XOR U9661 ( .A(n9515), .B(n9514), .Z(n9637) );
  IV U9662 ( .A(n9437), .Z(n9438) );
  NOR U9663 ( .A(n9439), .B(n9438), .Z(n9443) );
  NOR U9664 ( .A(n9441), .B(n9440), .Z(n9442) );
  NOR U9665 ( .A(n9443), .B(n9442), .Z(n9635) );
  NOR U9666 ( .A(n145), .B(n129), .Z(n9633) );
  XOR U9667 ( .A(n9635), .B(n9633), .Z(n9636) );
  XOR U9668 ( .A(n9637), .B(n9636), .Z(n9506) );
  XOR U9669 ( .A(n9507), .B(n9506), .Z(n9444) );
  IV U9670 ( .A(n9444), .Z(n9508) );
  XOR U9671 ( .A(n9509), .B(n9508), .Z(n9501) );
  IV U9672 ( .A(n9445), .Z(n9447) );
  NOR U9673 ( .A(n9447), .B(n9446), .Z(n9451) );
  NOR U9674 ( .A(n9449), .B(n9448), .Z(n9450) );
  NOR U9675 ( .A(n9451), .B(n9450), .Z(n9499) );
  XOR U9676 ( .A(n9501), .B(n9499), .Z(n9503) );
  NOR U9677 ( .A(n148), .B(n124), .Z(n9452) );
  IV U9678 ( .A(n9452), .Z(n9502) );
  XOR U9679 ( .A(n9503), .B(n9502), .Z(n9493) );
  XOR U9680 ( .A(n9453), .B(n9493), .Z(n9495) );
  XOR U9681 ( .A(n9496), .B(n9495), .Z(n9488) );
  NOR U9682 ( .A(n153), .B(n121), .Z(n9486) );
  XOR U9683 ( .A(n9488), .B(n9486), .Z(n9489) );
  XOR U9684 ( .A(n9454), .B(n9489), .Z(n9480) );
  XOR U9685 ( .A(n9478), .B(n9480), .Z(n9481) );
  XOR U9686 ( .A(n9482), .B(n9481), .Z(n9472) );
  XOR U9687 ( .A(n9473), .B(n9472), .Z(n9455) );
  IV U9688 ( .A(n9455), .Z(n9474) );
  XOR U9689 ( .A(n9475), .B(n9474), .Z(n9467) );
  NOR U9690 ( .A(n158), .B(n42), .Z(n9465) );
  XOR U9691 ( .A(n9467), .B(n9465), .Z(n9468) );
  XOR U9692 ( .A(n9469), .B(n9468), .Z(n9457) );
  IV U9693 ( .A(n9457), .Z(n9456) );
  NOR U9694 ( .A(n9458), .B(n9456), .Z(n9461) );
  XOR U9695 ( .A(n9458), .B(n9457), .Z(n10890) );
  NOR U9696 ( .A(n161), .B(n44), .Z(n9459) );
  IV U9697 ( .A(n9459), .Z(n10889) );
  NOR U9698 ( .A(n10890), .B(n10889), .Z(n9460) );
  NOR U9699 ( .A(n9461), .B(n9460), .Z(n9464) );
  NOR U9700 ( .A(n163), .B(n44), .Z(n9463) );
  IV U9701 ( .A(n9463), .Z(n9462) );
  NOR U9702 ( .A(n9464), .B(n9462), .Z(n9643) );
  XOR U9703 ( .A(n9464), .B(n9463), .Z(n10897) );
  IV U9704 ( .A(n9465), .Z(n9466) );
  NOR U9705 ( .A(n9467), .B(n9466), .Z(n9471) );
  NOR U9706 ( .A(n9469), .B(n9468), .Z(n9470) );
  NOR U9707 ( .A(n9471), .B(n9470), .Z(n9834) );
  NOR U9708 ( .A(n161), .B(n42), .Z(n9830) );
  NOR U9709 ( .A(n9473), .B(n9472), .Z(n9477) );
  NOR U9710 ( .A(n9475), .B(n9474), .Z(n9476) );
  NOR U9711 ( .A(n9477), .B(n9476), .Z(n9648) );
  IV U9712 ( .A(n9478), .Z(n9479) );
  NOR U9713 ( .A(n9480), .B(n9479), .Z(n9484) );
  NOR U9714 ( .A(n9482), .B(n9481), .Z(n9483) );
  NOR U9715 ( .A(n9484), .B(n9483), .Z(n9485) );
  IV U9716 ( .A(n9485), .Z(n9656) );
  NOR U9717 ( .A(n156), .B(n118), .Z(n9654) );
  IV U9718 ( .A(n9486), .Z(n9487) );
  NOR U9719 ( .A(n9488), .B(n9487), .Z(n9492) );
  NOR U9720 ( .A(n9490), .B(n9489), .Z(n9491) );
  NOR U9721 ( .A(n9492), .B(n9491), .Z(n9663) );
  NOR U9722 ( .A(n9494), .B(n9493), .Z(n9498) );
  NOR U9723 ( .A(n9496), .B(n9495), .Z(n9497) );
  NOR U9724 ( .A(n9498), .B(n9497), .Z(n9670) );
  NOR U9725 ( .A(n153), .B(n122), .Z(n9668) );
  NOR U9726 ( .A(n150), .B(n124), .Z(n9823) );
  IV U9727 ( .A(n9499), .Z(n9500) );
  NOR U9728 ( .A(n9501), .B(n9500), .Z(n9505) );
  NOR U9729 ( .A(n9503), .B(n9502), .Z(n9504) );
  NOR U9730 ( .A(n9505), .B(n9504), .Z(n9819) );
  NOR U9731 ( .A(n9507), .B(n9506), .Z(n9511) );
  NOR U9732 ( .A(n9509), .B(n9508), .Z(n9510) );
  NOR U9733 ( .A(n9511), .B(n9510), .Z(n9677) );
  NOR U9734 ( .A(n148), .B(n127), .Z(n9674) );
  NOR U9735 ( .A(n9513), .B(n9512), .Z(n9517) );
  NOR U9736 ( .A(n9515), .B(n9514), .Z(n9516) );
  NOR U9737 ( .A(n9517), .B(n9516), .Z(n9684) );
  NOR U9738 ( .A(n145), .B(n130), .Z(n9682) );
  NOR U9739 ( .A(n9519), .B(n9518), .Z(n9523) );
  NOR U9740 ( .A(n9521), .B(n9520), .Z(n9522) );
  NOR U9741 ( .A(n9523), .B(n9522), .Z(n9691) );
  NOR U9742 ( .A(n141), .B(n134), .Z(n9688) );
  NOR U9743 ( .A(n9525), .B(n9524), .Z(n9529) );
  NOR U9744 ( .A(n9527), .B(n9526), .Z(n9528) );
  NOR U9745 ( .A(n9529), .B(n9528), .Z(n9704) );
  NOR U9746 ( .A(n137), .B(n138), .Z(n9702) );
  NOR U9747 ( .A(n9531), .B(n9530), .Z(n9535) );
  NOR U9748 ( .A(n9533), .B(n9532), .Z(n9534) );
  NOR U9749 ( .A(n9535), .B(n9534), .Z(n9798) );
  NOR U9750 ( .A(n9537), .B(n9536), .Z(n9541) );
  NOR U9751 ( .A(n9539), .B(n9538), .Z(n9540) );
  NOR U9752 ( .A(n9541), .B(n9540), .Z(n9710) );
  NOR U9753 ( .A(n133), .B(n142), .Z(n9708) );
  IV U9754 ( .A(n9542), .Z(n9543) );
  NOR U9755 ( .A(n9544), .B(n9543), .Z(n9548) );
  NOR U9756 ( .A(n9546), .B(n9545), .Z(n9547) );
  NOR U9757 ( .A(n9548), .B(n9547), .Z(n9791) );
  NOR U9758 ( .A(n9550), .B(n9549), .Z(n9554) );
  NOR U9759 ( .A(n9552), .B(n9551), .Z(n9553) );
  NOR U9760 ( .A(n9554), .B(n9553), .Z(n9717) );
  NOR U9761 ( .A(n128), .B(n146), .Z(n9715) );
  NOR U9762 ( .A(n126), .B(n149), .Z(n9782) );
  NOR U9763 ( .A(n9556), .B(n9555), .Z(n9560) );
  NOR U9764 ( .A(n9558), .B(n9557), .Z(n9559) );
  NOR U9765 ( .A(n9560), .B(n9559), .Z(n9778) );
  NOR U9766 ( .A(n9562), .B(n9561), .Z(n9566) );
  NOR U9767 ( .A(n9564), .B(n9563), .Z(n9565) );
  NOR U9768 ( .A(n9566), .B(n9565), .Z(n9724) );
  NOR U9769 ( .A(n125), .B(n151), .Z(n9721) );
  NOR U9770 ( .A(n9568), .B(n9567), .Z(n9573) );
  IV U9771 ( .A(n9569), .Z(n9571) );
  NOR U9772 ( .A(n9571), .B(n9570), .Z(n9572) );
  NOR U9773 ( .A(n9573), .B(n9572), .Z(n9574) );
  IV U9774 ( .A(n9574), .Z(n9729) );
  NOR U9775 ( .A(n123), .B(n152), .Z(n9727) );
  XOR U9776 ( .A(n9729), .B(n9727), .Z(n9730) );
  NOR U9777 ( .A(n9576), .B(n9575), .Z(n9581) );
  IV U9778 ( .A(n9577), .Z(n9578) );
  NOR U9779 ( .A(n9579), .B(n9578), .Z(n9580) );
  NOR U9780 ( .A(n9581), .B(n9580), .Z(n9737) );
  NOR U9781 ( .A(n120), .B(n154), .Z(n9735) );
  IV U9782 ( .A(n9735), .Z(n9617) );
  NOR U9783 ( .A(n9583), .B(n9582), .Z(n9587) );
  NOR U9784 ( .A(n9585), .B(n9584), .Z(n9586) );
  NOR U9785 ( .A(n9587), .B(n9586), .Z(n9743) );
  NOR U9786 ( .A(n79), .B(n159), .Z(n9741) );
  NOR U9787 ( .A(n9589), .B(n9588), .Z(n9593) );
  NOR U9788 ( .A(n9591), .B(n9590), .Z(n9592) );
  NOR U9789 ( .A(n9593), .B(n9592), .Z(n9765) );
  NOR U9790 ( .A(n9595), .B(n9594), .Z(n9599) );
  NOR U9791 ( .A(n9597), .B(n9596), .Z(n9598) );
  NOR U9792 ( .A(n9599), .B(n9598), .Z(n9749) );
  NOR U9793 ( .A(n80), .B(n162), .Z(n9747) );
  IV U9794 ( .A(n9747), .Z(n9608) );
  IV U9795 ( .A(n9600), .Z(n9601) );
  NOR U9796 ( .A(n9602), .B(n9601), .Z(n9606) );
  NOR U9797 ( .A(n9604), .B(n9603), .Z(n9605) );
  NOR U9798 ( .A(n9606), .B(n9605), .Z(n9754) );
  NOR U9799 ( .A(n164), .B(n116), .Z(n9752) );
  XOR U9800 ( .A(n9754), .B(n9752), .Z(n9756) );
  NOR U9801 ( .A(n166), .B(n81), .Z(n9607) );
  IV U9802 ( .A(n9607), .Z(n9755) );
  XOR U9803 ( .A(n9756), .B(n9755), .Z(n9746) );
  XOR U9804 ( .A(n9608), .B(n9746), .Z(n9748) );
  XOR U9805 ( .A(n9749), .B(n9748), .Z(n9763) );
  NOR U9806 ( .A(n117), .B(n160), .Z(n9761) );
  XOR U9807 ( .A(n9763), .B(n9761), .Z(n9764) );
  XOR U9808 ( .A(n9765), .B(n9764), .Z(n9740) );
  XOR U9809 ( .A(n9741), .B(n9740), .Z(n9609) );
  IV U9810 ( .A(n9609), .Z(n9742) );
  XOR U9811 ( .A(n9743), .B(n9742), .Z(n9773) );
  IV U9812 ( .A(n9610), .Z(n9611) );
  NOR U9813 ( .A(n9612), .B(n9611), .Z(n9616) );
  NOR U9814 ( .A(n9614), .B(n9613), .Z(n9615) );
  NOR U9815 ( .A(n9616), .B(n9615), .Z(n9771) );
  NOR U9816 ( .A(n119), .B(n157), .Z(n9769) );
  XOR U9817 ( .A(n9771), .B(n9769), .Z(n9772) );
  XOR U9818 ( .A(n9773), .B(n9772), .Z(n9734) );
  XOR U9819 ( .A(n9617), .B(n9734), .Z(n9736) );
  XOR U9820 ( .A(n9737), .B(n9736), .Z(n9731) );
  XOR U9821 ( .A(n9730), .B(n9731), .Z(n9720) );
  XOR U9822 ( .A(n9721), .B(n9720), .Z(n9722) );
  XOR U9823 ( .A(n9724), .B(n9722), .Z(n9779) );
  XOR U9824 ( .A(n9778), .B(n9779), .Z(n9781) );
  XOR U9825 ( .A(n9782), .B(n9781), .Z(n9713) );
  XOR U9826 ( .A(n9715), .B(n9713), .Z(n9716) );
  XOR U9827 ( .A(n9717), .B(n9716), .Z(n9789) );
  NOR U9828 ( .A(n131), .B(n144), .Z(n9787) );
  XOR U9829 ( .A(n9789), .B(n9787), .Z(n9790) );
  XOR U9830 ( .A(n9791), .B(n9790), .Z(n9707) );
  XOR U9831 ( .A(n9708), .B(n9707), .Z(n9618) );
  IV U9832 ( .A(n9618), .Z(n9709) );
  XOR U9833 ( .A(n9710), .B(n9709), .Z(n9796) );
  NOR U9834 ( .A(n135), .B(n140), .Z(n9794) );
  XOR U9835 ( .A(n9796), .B(n9794), .Z(n9797) );
  XOR U9836 ( .A(n9798), .B(n9797), .Z(n9701) );
  XOR U9837 ( .A(n9702), .B(n9701), .Z(n9619) );
  IV U9838 ( .A(n9619), .Z(n9703) );
  XOR U9839 ( .A(n9704), .B(n9703), .Z(n9698) );
  IV U9840 ( .A(n9620), .Z(n9621) );
  NOR U9841 ( .A(n9622), .B(n9621), .Z(n9626) );
  NOR U9842 ( .A(n9624), .B(n9623), .Z(n9625) );
  NOR U9843 ( .A(n9626), .B(n9625), .Z(n9696) );
  NOR U9844 ( .A(n139), .B(n136), .Z(n9694) );
  XOR U9845 ( .A(n9696), .B(n9694), .Z(n9697) );
  XOR U9846 ( .A(n9698), .B(n9697), .Z(n9687) );
  XOR U9847 ( .A(n9688), .B(n9687), .Z(n9689) );
  XOR U9848 ( .A(n9691), .B(n9689), .Z(n9805) );
  NOR U9849 ( .A(n143), .B(n132), .Z(n9804) );
  NOR U9850 ( .A(n9628), .B(n9627), .Z(n9632) );
  NOR U9851 ( .A(n9630), .B(n9629), .Z(n9631) );
  NOR U9852 ( .A(n9632), .B(n9631), .Z(n9802) );
  XOR U9853 ( .A(n9804), .B(n9802), .Z(n9806) );
  XOR U9854 ( .A(n9805), .B(n9806), .Z(n9680) );
  XOR U9855 ( .A(n9682), .B(n9680), .Z(n9683) );
  XOR U9856 ( .A(n9684), .B(n9683), .Z(n9815) );
  IV U9857 ( .A(n9633), .Z(n9634) );
  NOR U9858 ( .A(n9635), .B(n9634), .Z(n9639) );
  NOR U9859 ( .A(n9637), .B(n9636), .Z(n9638) );
  NOR U9860 ( .A(n9639), .B(n9638), .Z(n9813) );
  NOR U9861 ( .A(n147), .B(n129), .Z(n9811) );
  XOR U9862 ( .A(n9813), .B(n9811), .Z(n9814) );
  XOR U9863 ( .A(n9815), .B(n9814), .Z(n9673) );
  XOR U9864 ( .A(n9674), .B(n9673), .Z(n9675) );
  XOR U9865 ( .A(n9677), .B(n9675), .Z(n9820) );
  XOR U9866 ( .A(n9819), .B(n9820), .Z(n9822) );
  XOR U9867 ( .A(n9823), .B(n9822), .Z(n9666) );
  XOR U9868 ( .A(n9668), .B(n9666), .Z(n9669) );
  XOR U9869 ( .A(n9670), .B(n9669), .Z(n9661) );
  NOR U9870 ( .A(n155), .B(n121), .Z(n9659) );
  XOR U9871 ( .A(n9661), .B(n9659), .Z(n9662) );
  XOR U9872 ( .A(n9663), .B(n9662), .Z(n9653) );
  XOR U9873 ( .A(n9654), .B(n9653), .Z(n9640) );
  IV U9874 ( .A(n9640), .Z(n9655) );
  XOR U9875 ( .A(n9656), .B(n9655), .Z(n9647) );
  NOR U9876 ( .A(n158), .B(n43), .Z(n9645) );
  XOR U9877 ( .A(n9647), .B(n9645), .Z(n9650) );
  XOR U9878 ( .A(n9648), .B(n9650), .Z(n9832) );
  XOR U9879 ( .A(n9830), .B(n9832), .Z(n9833) );
  XOR U9880 ( .A(n9834), .B(n9833), .Z(n10896) );
  IV U9881 ( .A(n10896), .Z(n9641) );
  NOR U9882 ( .A(n10897), .B(n9641), .Z(n9642) );
  NOR U9883 ( .A(n9643), .B(n9642), .Z(n9839) );
  NOR U9884 ( .A(n165), .B(n44), .Z(n9838) );
  IV U9885 ( .A(n9838), .Z(n9644) );
  NOR U9886 ( .A(n9839), .B(n9644), .Z(n9841) );
  NOR U9887 ( .A(n163), .B(n42), .Z(n9843) );
  IV U9888 ( .A(n9645), .Z(n9646) );
  NOR U9889 ( .A(n9647), .B(n9646), .Z(n9652) );
  IV U9890 ( .A(n9648), .Z(n9649) );
  NOR U9891 ( .A(n9650), .B(n9649), .Z(n9651) );
  NOR U9892 ( .A(n9652), .B(n9651), .Z(n9852) );
  NOR U9893 ( .A(n161), .B(n43), .Z(n9848) );
  NOR U9894 ( .A(n9654), .B(n9653), .Z(n9658) );
  NOR U9895 ( .A(n9656), .B(n9655), .Z(n9657) );
  NOR U9896 ( .A(n9658), .B(n9657), .Z(n9859) );
  NOR U9897 ( .A(n158), .B(n118), .Z(n9856) );
  IV U9898 ( .A(n9659), .Z(n9660) );
  NOR U9899 ( .A(n9661), .B(n9660), .Z(n9665) );
  NOR U9900 ( .A(n9663), .B(n9662), .Z(n9664) );
  NOR U9901 ( .A(n9665), .B(n9664), .Z(n9868) );
  IV U9902 ( .A(n9868), .Z(n9828) );
  IV U9903 ( .A(n9666), .Z(n9667) );
  NOR U9904 ( .A(n9668), .B(n9667), .Z(n9672) );
  NOR U9905 ( .A(n9670), .B(n9669), .Z(n9671) );
  NOR U9906 ( .A(n9672), .B(n9671), .Z(n9874) );
  NOR U9907 ( .A(n155), .B(n122), .Z(n9872) );
  IV U9908 ( .A(n9872), .Z(n9827) );
  NOR U9909 ( .A(n9674), .B(n9673), .Z(n9679) );
  IV U9910 ( .A(n9675), .Z(n9676) );
  NOR U9911 ( .A(n9677), .B(n9676), .Z(n9678) );
  NOR U9912 ( .A(n9679), .B(n9678), .Z(n9880) );
  NOR U9913 ( .A(n150), .B(n127), .Z(n9878) );
  IV U9914 ( .A(n9680), .Z(n9681) );
  NOR U9915 ( .A(n9682), .B(n9681), .Z(n9686) );
  NOR U9916 ( .A(n9684), .B(n9683), .Z(n9685) );
  NOR U9917 ( .A(n9686), .B(n9685), .Z(n9893) );
  NOR U9918 ( .A(n147), .B(n130), .Z(n9891) );
  IV U9919 ( .A(n9891), .Z(n9810) );
  NOR U9920 ( .A(n9688), .B(n9687), .Z(n9693) );
  IV U9921 ( .A(n9689), .Z(n9690) );
  NOR U9922 ( .A(n9691), .B(n9690), .Z(n9692) );
  NOR U9923 ( .A(n9693), .B(n9692), .Z(n9906) );
  NOR U9924 ( .A(n143), .B(n134), .Z(n9904) );
  IV U9925 ( .A(n9694), .Z(n9695) );
  NOR U9926 ( .A(n9696), .B(n9695), .Z(n9700) );
  NOR U9927 ( .A(n9698), .B(n9697), .Z(n9699) );
  NOR U9928 ( .A(n9700), .B(n9699), .Z(n10019) );
  NOR U9929 ( .A(n9702), .B(n9701), .Z(n9706) );
  NOR U9930 ( .A(n9704), .B(n9703), .Z(n9705) );
  NOR U9931 ( .A(n9706), .B(n9705), .Z(n9913) );
  NOR U9932 ( .A(n139), .B(n138), .Z(n9911) );
  NOR U9933 ( .A(n9708), .B(n9707), .Z(n9712) );
  NOR U9934 ( .A(n9710), .B(n9709), .Z(n9711) );
  NOR U9935 ( .A(n9712), .B(n9711), .Z(n9920) );
  NOR U9936 ( .A(n135), .B(n142), .Z(n9917) );
  IV U9937 ( .A(n9713), .Z(n9714) );
  NOR U9938 ( .A(n9715), .B(n9714), .Z(n9719) );
  NOR U9939 ( .A(n9717), .B(n9716), .Z(n9718) );
  NOR U9940 ( .A(n9719), .B(n9718), .Z(n9933) );
  NOR U9941 ( .A(n131), .B(n146), .Z(n9931) );
  IV U9942 ( .A(n9931), .Z(n9786) );
  NOR U9943 ( .A(n9721), .B(n9720), .Z(n9726) );
  IV U9944 ( .A(n9722), .Z(n9723) );
  NOR U9945 ( .A(n9724), .B(n9723), .Z(n9725) );
  NOR U9946 ( .A(n9726), .B(n9725), .Z(n9946) );
  NOR U9947 ( .A(n126), .B(n151), .Z(n9944) );
  IV U9948 ( .A(n9944), .Z(n9777) );
  IV U9949 ( .A(n9727), .Z(n9728) );
  NOR U9950 ( .A(n9729), .B(n9728), .Z(n9733) );
  NOR U9951 ( .A(n9731), .B(n9730), .Z(n9732) );
  NOR U9952 ( .A(n9733), .B(n9732), .Z(n9997) );
  NOR U9953 ( .A(n125), .B(n152), .Z(n9996) );
  NOR U9954 ( .A(n9735), .B(n9734), .Z(n9739) );
  NOR U9955 ( .A(n9737), .B(n9736), .Z(n9738) );
  NOR U9956 ( .A(n9739), .B(n9738), .Z(n9953) );
  NOR U9957 ( .A(n123), .B(n154), .Z(n9950) );
  NOR U9958 ( .A(n9741), .B(n9740), .Z(n9745) );
  NOR U9959 ( .A(n9743), .B(n9742), .Z(n9744) );
  NOR U9960 ( .A(n9745), .B(n9744), .Z(n9959) );
  NOR U9961 ( .A(n119), .B(n159), .Z(n9957) );
  NOR U9962 ( .A(n9747), .B(n9746), .Z(n9751) );
  NOR U9963 ( .A(n9749), .B(n9748), .Z(n9750) );
  NOR U9964 ( .A(n9751), .B(n9750), .Z(n9972) );
  NOR U9965 ( .A(n117), .B(n162), .Z(n9970) );
  IV U9966 ( .A(n9970), .Z(n9760) );
  IV U9967 ( .A(n9752), .Z(n9753) );
  NOR U9968 ( .A(n9754), .B(n9753), .Z(n9758) );
  NOR U9969 ( .A(n9756), .B(n9755), .Z(n9757) );
  NOR U9970 ( .A(n9758), .B(n9757), .Z(n9977) );
  NOR U9971 ( .A(n164), .B(n80), .Z(n9975) );
  XOR U9972 ( .A(n9977), .B(n9975), .Z(n9979) );
  NOR U9973 ( .A(n166), .B(n116), .Z(n9759) );
  IV U9974 ( .A(n9759), .Z(n9978) );
  XOR U9975 ( .A(n9979), .B(n9978), .Z(n9969) );
  XOR U9976 ( .A(n9760), .B(n9969), .Z(n9971) );
  XOR U9977 ( .A(n9972), .B(n9971), .Z(n9966) );
  IV U9978 ( .A(n9761), .Z(n9762) );
  NOR U9979 ( .A(n9763), .B(n9762), .Z(n9767) );
  NOR U9980 ( .A(n9765), .B(n9764), .Z(n9766) );
  NOR U9981 ( .A(n9767), .B(n9766), .Z(n9964) );
  NOR U9982 ( .A(n79), .B(n160), .Z(n9962) );
  XOR U9983 ( .A(n9964), .B(n9962), .Z(n9965) );
  XOR U9984 ( .A(n9966), .B(n9965), .Z(n9956) );
  XOR U9985 ( .A(n9957), .B(n9956), .Z(n9768) );
  IV U9986 ( .A(n9768), .Z(n9958) );
  XOR U9987 ( .A(n9959), .B(n9958), .Z(n9991) );
  IV U9988 ( .A(n9769), .Z(n9770) );
  NOR U9989 ( .A(n9771), .B(n9770), .Z(n9775) );
  NOR U9990 ( .A(n9773), .B(n9772), .Z(n9774) );
  NOR U9991 ( .A(n9775), .B(n9774), .Z(n9989) );
  NOR U9992 ( .A(n120), .B(n157), .Z(n9987) );
  XOR U9993 ( .A(n9989), .B(n9987), .Z(n9990) );
  XOR U9994 ( .A(n9991), .B(n9990), .Z(n9949) );
  XOR U9995 ( .A(n9950), .B(n9949), .Z(n9951) );
  XOR U9996 ( .A(n9953), .B(n9951), .Z(n9995) );
  XOR U9997 ( .A(n9996), .B(n9995), .Z(n9776) );
  IV U9998 ( .A(n9776), .Z(n9998) );
  XOR U9999 ( .A(n9997), .B(n9998), .Z(n9943) );
  XOR U10000 ( .A(n9777), .B(n9943), .Z(n9945) );
  XOR U10001 ( .A(n9946), .B(n9945), .Z(n9938) );
  IV U10002 ( .A(n9778), .Z(n9780) );
  NOR U10003 ( .A(n9780), .B(n9779), .Z(n9784) );
  NOR U10004 ( .A(n9782), .B(n9781), .Z(n9783) );
  NOR U10005 ( .A(n9784), .B(n9783), .Z(n9936) );
  XOR U10006 ( .A(n9938), .B(n9936), .Z(n9940) );
  NOR U10007 ( .A(n128), .B(n149), .Z(n9785) );
  IV U10008 ( .A(n9785), .Z(n9939) );
  XOR U10009 ( .A(n9940), .B(n9939), .Z(n9930) );
  XOR U10010 ( .A(n9786), .B(n9930), .Z(n9932) );
  XOR U10011 ( .A(n9933), .B(n9932), .Z(n9927) );
  IV U10012 ( .A(n9787), .Z(n9788) );
  NOR U10013 ( .A(n9789), .B(n9788), .Z(n9793) );
  NOR U10014 ( .A(n9791), .B(n9790), .Z(n9792) );
  NOR U10015 ( .A(n9793), .B(n9792), .Z(n9925) );
  NOR U10016 ( .A(n133), .B(n144), .Z(n9923) );
  XOR U10017 ( .A(n9925), .B(n9923), .Z(n9926) );
  XOR U10018 ( .A(n9927), .B(n9926), .Z(n9916) );
  XOR U10019 ( .A(n9917), .B(n9916), .Z(n9918) );
  XOR U10020 ( .A(n9920), .B(n9918), .Z(n10009) );
  NOR U10021 ( .A(n137), .B(n140), .Z(n10008) );
  IV U10022 ( .A(n9794), .Z(n9795) );
  NOR U10023 ( .A(n9796), .B(n9795), .Z(n9800) );
  NOR U10024 ( .A(n9798), .B(n9797), .Z(n9799) );
  NOR U10025 ( .A(n9800), .B(n9799), .Z(n10006) );
  XOR U10026 ( .A(n10008), .B(n10006), .Z(n10010) );
  XOR U10027 ( .A(n10009), .B(n10010), .Z(n9909) );
  XOR U10028 ( .A(n9911), .B(n9909), .Z(n9912) );
  XOR U10029 ( .A(n9913), .B(n9912), .Z(n10017) );
  NOR U10030 ( .A(n141), .B(n136), .Z(n10015) );
  XOR U10031 ( .A(n10017), .B(n10015), .Z(n10018) );
  XOR U10032 ( .A(n10019), .B(n10018), .Z(n9903) );
  XOR U10033 ( .A(n9904), .B(n9903), .Z(n9801) );
  IV U10034 ( .A(n9801), .Z(n9905) );
  XOR U10035 ( .A(n9906), .B(n9905), .Z(n9898) );
  IV U10036 ( .A(n9802), .Z(n9803) );
  NOR U10037 ( .A(n9804), .B(n9803), .Z(n9808) );
  NOR U10038 ( .A(n9806), .B(n9805), .Z(n9807) );
  NOR U10039 ( .A(n9808), .B(n9807), .Z(n9896) );
  XOR U10040 ( .A(n9898), .B(n9896), .Z(n9900) );
  NOR U10041 ( .A(n145), .B(n132), .Z(n9809) );
  IV U10042 ( .A(n9809), .Z(n9899) );
  XOR U10043 ( .A(n9900), .B(n9899), .Z(n9890) );
  XOR U10044 ( .A(n9810), .B(n9890), .Z(n9892) );
  XOR U10045 ( .A(n9893), .B(n9892), .Z(n9887) );
  IV U10046 ( .A(n9811), .Z(n9812) );
  NOR U10047 ( .A(n9813), .B(n9812), .Z(n9817) );
  NOR U10048 ( .A(n9815), .B(n9814), .Z(n9816) );
  NOR U10049 ( .A(n9817), .B(n9816), .Z(n9885) );
  NOR U10050 ( .A(n148), .B(n129), .Z(n9883) );
  XOR U10051 ( .A(n9885), .B(n9883), .Z(n9886) );
  XOR U10052 ( .A(n9887), .B(n9886), .Z(n9877) );
  XOR U10053 ( .A(n9878), .B(n9877), .Z(n9818) );
  IV U10054 ( .A(n9818), .Z(n9879) );
  XOR U10055 ( .A(n9880), .B(n9879), .Z(n10029) );
  NOR U10056 ( .A(n153), .B(n124), .Z(n10027) );
  XOR U10057 ( .A(n10029), .B(n10027), .Z(n10031) );
  IV U10058 ( .A(n9819), .Z(n9821) );
  NOR U10059 ( .A(n9821), .B(n9820), .Z(n9825) );
  NOR U10060 ( .A(n9823), .B(n9822), .Z(n9824) );
  NOR U10061 ( .A(n9825), .B(n9824), .Z(n9826) );
  IV U10062 ( .A(n9826), .Z(n10030) );
  XOR U10063 ( .A(n10031), .B(n10030), .Z(n9871) );
  XOR U10064 ( .A(n9827), .B(n9871), .Z(n9873) );
  XOR U10065 ( .A(n9874), .B(n9873), .Z(n9866) );
  NOR U10066 ( .A(n156), .B(n121), .Z(n9864) );
  XOR U10067 ( .A(n9866), .B(n9864), .Z(n9867) );
  XOR U10068 ( .A(n9828), .B(n9867), .Z(n9858) );
  XOR U10069 ( .A(n9856), .B(n9858), .Z(n9861) );
  XOR U10070 ( .A(n9859), .B(n9861), .Z(n9850) );
  XOR U10071 ( .A(n9848), .B(n9850), .Z(n9851) );
  XOR U10072 ( .A(n9852), .B(n9851), .Z(n9842) );
  XOR U10073 ( .A(n9843), .B(n9842), .Z(n9829) );
  IV U10074 ( .A(n9829), .Z(n9845) );
  IV U10075 ( .A(n9830), .Z(n9831) );
  NOR U10076 ( .A(n9832), .B(n9831), .Z(n9836) );
  NOR U10077 ( .A(n9834), .B(n9833), .Z(n9835) );
  NOR U10078 ( .A(n9836), .B(n9835), .Z(n9837) );
  IV U10079 ( .A(n9837), .Z(n9844) );
  XOR U10080 ( .A(n9845), .B(n9844), .Z(n11384) );
  XOR U10081 ( .A(n9839), .B(n9838), .Z(n11383) );
  NOR U10082 ( .A(n11384), .B(n11383), .Z(n9840) );
  NOR U10083 ( .A(n9841), .B(n9840), .Z(n10037) );
  NOR U10084 ( .A(n9843), .B(n9842), .Z(n9847) );
  NOR U10085 ( .A(n9845), .B(n9844), .Z(n9846) );
  NOR U10086 ( .A(n9847), .B(n9846), .Z(n10046) );
  IV U10087 ( .A(n9848), .Z(n9849) );
  NOR U10088 ( .A(n9850), .B(n9849), .Z(n9854) );
  NOR U10089 ( .A(n9852), .B(n9851), .Z(n9853) );
  NOR U10090 ( .A(n9854), .B(n9853), .Z(n9855) );
  IV U10091 ( .A(n9855), .Z(n10054) );
  NOR U10092 ( .A(n163), .B(n43), .Z(n10052) );
  IV U10093 ( .A(n9856), .Z(n9857) );
  NOR U10094 ( .A(n9858), .B(n9857), .Z(n9863) );
  IV U10095 ( .A(n9859), .Z(n9860) );
  NOR U10096 ( .A(n9861), .B(n9860), .Z(n9862) );
  NOR U10097 ( .A(n9863), .B(n9862), .Z(n10061) );
  NOR U10098 ( .A(n161), .B(n118), .Z(n10057) );
  IV U10099 ( .A(n9864), .Z(n9865) );
  NOR U10100 ( .A(n9866), .B(n9865), .Z(n9870) );
  NOR U10101 ( .A(n9868), .B(n9867), .Z(n9869) );
  NOR U10102 ( .A(n9870), .B(n9869), .Z(n10068) );
  IV U10103 ( .A(n10068), .Z(n10035) );
  NOR U10104 ( .A(n9872), .B(n9871), .Z(n9876) );
  NOR U10105 ( .A(n9874), .B(n9873), .Z(n9875) );
  NOR U10106 ( .A(n9876), .B(n9875), .Z(n10074) );
  NOR U10107 ( .A(n156), .B(n122), .Z(n10072) );
  NOR U10108 ( .A(n9878), .B(n9877), .Z(n9882) );
  NOR U10109 ( .A(n9880), .B(n9879), .Z(n9881) );
  NOR U10110 ( .A(n9882), .B(n9881), .Z(n10087) );
  NOR U10111 ( .A(n153), .B(n127), .Z(n10085) );
  IV U10112 ( .A(n9883), .Z(n9884) );
  NOR U10113 ( .A(n9885), .B(n9884), .Z(n9889) );
  NOR U10114 ( .A(n9887), .B(n9886), .Z(n9888) );
  NOR U10115 ( .A(n9889), .B(n9888), .Z(n10217) );
  NOR U10116 ( .A(n9891), .B(n9890), .Z(n9895) );
  NOR U10117 ( .A(n9893), .B(n9892), .Z(n9894) );
  NOR U10118 ( .A(n9895), .B(n9894), .Z(n10093) );
  NOR U10119 ( .A(n148), .B(n130), .Z(n10091) );
  IV U10120 ( .A(n10091), .Z(n10025) );
  IV U10121 ( .A(n9896), .Z(n9897) );
  NOR U10122 ( .A(n9898), .B(n9897), .Z(n9902) );
  NOR U10123 ( .A(n9900), .B(n9899), .Z(n9901) );
  NOR U10124 ( .A(n9902), .B(n9901), .Z(n10206) );
  IV U10125 ( .A(n10206), .Z(n10023) );
  NOR U10126 ( .A(n9904), .B(n9903), .Z(n9908) );
  NOR U10127 ( .A(n9906), .B(n9905), .Z(n9907) );
  NOR U10128 ( .A(n9908), .B(n9907), .Z(n10099) );
  NOR U10129 ( .A(n145), .B(n134), .Z(n10097) );
  IV U10130 ( .A(n10097), .Z(n10022) );
  IV U10131 ( .A(n9909), .Z(n9910) );
  NOR U10132 ( .A(n9911), .B(n9910), .Z(n9915) );
  NOR U10133 ( .A(n9913), .B(n9912), .Z(n9914) );
  NOR U10134 ( .A(n9915), .B(n9914), .Z(n10105) );
  NOR U10135 ( .A(n141), .B(n138), .Z(n10103) );
  IV U10136 ( .A(n10103), .Z(n10014) );
  NOR U10137 ( .A(n9917), .B(n9916), .Z(n9922) );
  IV U10138 ( .A(n9918), .Z(n9919) );
  NOR U10139 ( .A(n9920), .B(n9919), .Z(n9921) );
  NOR U10140 ( .A(n9922), .B(n9921), .Z(n10111) );
  NOR U10141 ( .A(n137), .B(n142), .Z(n10109) );
  IV U10142 ( .A(n10109), .Z(n10005) );
  IV U10143 ( .A(n9923), .Z(n9924) );
  NOR U10144 ( .A(n9925), .B(n9924), .Z(n9929) );
  NOR U10145 ( .A(n9927), .B(n9926), .Z(n9928) );
  NOR U10146 ( .A(n9929), .B(n9928), .Z(n10114) );
  IV U10147 ( .A(n10114), .Z(n10003) );
  NOR U10148 ( .A(n9931), .B(n9930), .Z(n9935) );
  NOR U10149 ( .A(n9933), .B(n9932), .Z(n9934) );
  NOR U10150 ( .A(n9935), .B(n9934), .Z(n10124) );
  NOR U10151 ( .A(n133), .B(n146), .Z(n10122) );
  NOR U10152 ( .A(n131), .B(n149), .Z(n10131) );
  IV U10153 ( .A(n9936), .Z(n9937) );
  NOR U10154 ( .A(n9938), .B(n9937), .Z(n9942) );
  NOR U10155 ( .A(n9940), .B(n9939), .Z(n9941) );
  NOR U10156 ( .A(n9942), .B(n9941), .Z(n10127) );
  NOR U10157 ( .A(n9944), .B(n9943), .Z(n9948) );
  NOR U10158 ( .A(n9946), .B(n9945), .Z(n9947) );
  NOR U10159 ( .A(n9948), .B(n9947), .Z(n10138) );
  NOR U10160 ( .A(n128), .B(n151), .Z(n10135) );
  NOR U10161 ( .A(n9950), .B(n9949), .Z(n9955) );
  IV U10162 ( .A(n9951), .Z(n9952) );
  NOR U10163 ( .A(n9953), .B(n9952), .Z(n9954) );
  NOR U10164 ( .A(n9955), .B(n9954), .Z(n10144) );
  NOR U10165 ( .A(n125), .B(n154), .Z(n10142) );
  NOR U10166 ( .A(n9957), .B(n9956), .Z(n9961) );
  NOR U10167 ( .A(n9959), .B(n9958), .Z(n9960) );
  NOR U10168 ( .A(n9961), .B(n9960), .Z(n10150) );
  NOR U10169 ( .A(n120), .B(n159), .Z(n10148) );
  IV U10170 ( .A(n10148), .Z(n9986) );
  IV U10171 ( .A(n9962), .Z(n9963) );
  NOR U10172 ( .A(n9964), .B(n9963), .Z(n9968) );
  NOR U10173 ( .A(n9966), .B(n9965), .Z(n9967) );
  NOR U10174 ( .A(n9968), .B(n9967), .Z(n10168) );
  IV U10175 ( .A(n10168), .Z(n9984) );
  NOR U10176 ( .A(n9970), .B(n9969), .Z(n9974) );
  NOR U10177 ( .A(n9972), .B(n9971), .Z(n9973) );
  NOR U10178 ( .A(n9974), .B(n9973), .Z(n10156) );
  NOR U10179 ( .A(n79), .B(n162), .Z(n10154) );
  IV U10180 ( .A(n10154), .Z(n9983) );
  IV U10181 ( .A(n9975), .Z(n9976) );
  NOR U10182 ( .A(n9977), .B(n9976), .Z(n9981) );
  NOR U10183 ( .A(n9979), .B(n9978), .Z(n9980) );
  NOR U10184 ( .A(n9981), .B(n9980), .Z(n10161) );
  NOR U10185 ( .A(n164), .B(n117), .Z(n10159) );
  XOR U10186 ( .A(n10161), .B(n10159), .Z(n10163) );
  NOR U10187 ( .A(n166), .B(n80), .Z(n9982) );
  IV U10188 ( .A(n9982), .Z(n10162) );
  XOR U10189 ( .A(n10163), .B(n10162), .Z(n10153) );
  XOR U10190 ( .A(n9983), .B(n10153), .Z(n10155) );
  XOR U10191 ( .A(n10156), .B(n10155), .Z(n10169) );
  XOR U10192 ( .A(n9984), .B(n10169), .Z(n10171) );
  NOR U10193 ( .A(n119), .B(n160), .Z(n9985) );
  IV U10194 ( .A(n9985), .Z(n10170) );
  XOR U10195 ( .A(n10171), .B(n10170), .Z(n10147) );
  XOR U10196 ( .A(n9986), .B(n10147), .Z(n10149) );
  XOR U10197 ( .A(n10150), .B(n10149), .Z(n10179) );
  IV U10198 ( .A(n9987), .Z(n9988) );
  NOR U10199 ( .A(n9989), .B(n9988), .Z(n9993) );
  NOR U10200 ( .A(n9991), .B(n9990), .Z(n9992) );
  NOR U10201 ( .A(n9993), .B(n9992), .Z(n10177) );
  NOR U10202 ( .A(n123), .B(n157), .Z(n10175) );
  XOR U10203 ( .A(n10177), .B(n10175), .Z(n10178) );
  XOR U10204 ( .A(n10179), .B(n10178), .Z(n10141) );
  XOR U10205 ( .A(n10142), .B(n10141), .Z(n9994) );
  IV U10206 ( .A(n9994), .Z(n10143) );
  XOR U10207 ( .A(n10144), .B(n10143), .Z(n10185) );
  NOR U10208 ( .A(n9996), .B(n9995), .Z(n10001) );
  IV U10209 ( .A(n9997), .Z(n9999) );
  NOR U10210 ( .A(n9999), .B(n9998), .Z(n10000) );
  NOR U10211 ( .A(n10001), .B(n10000), .Z(n10183) );
  XOR U10212 ( .A(n10185), .B(n10183), .Z(n10187) );
  NOR U10213 ( .A(n126), .B(n152), .Z(n10002) );
  IV U10214 ( .A(n10002), .Z(n10186) );
  XOR U10215 ( .A(n10187), .B(n10186), .Z(n10134) );
  XOR U10216 ( .A(n10135), .B(n10134), .Z(n10136) );
  XOR U10217 ( .A(n10138), .B(n10136), .Z(n10128) );
  XOR U10218 ( .A(n10127), .B(n10128), .Z(n10130) );
  XOR U10219 ( .A(n10131), .B(n10130), .Z(n10120) );
  XOR U10220 ( .A(n10122), .B(n10120), .Z(n10123) );
  XOR U10221 ( .A(n10124), .B(n10123), .Z(n10115) );
  XOR U10222 ( .A(n10003), .B(n10115), .Z(n10117) );
  NOR U10223 ( .A(n135), .B(n144), .Z(n10004) );
  IV U10224 ( .A(n10004), .Z(n10116) );
  XOR U10225 ( .A(n10117), .B(n10116), .Z(n10108) );
  XOR U10226 ( .A(n10005), .B(n10108), .Z(n10110) );
  XOR U10227 ( .A(n10111), .B(n10110), .Z(n10192) );
  IV U10228 ( .A(n10006), .Z(n10007) );
  NOR U10229 ( .A(n10008), .B(n10007), .Z(n10012) );
  NOR U10230 ( .A(n10010), .B(n10009), .Z(n10011) );
  NOR U10231 ( .A(n10012), .B(n10011), .Z(n10190) );
  XOR U10232 ( .A(n10192), .B(n10190), .Z(n10194) );
  NOR U10233 ( .A(n139), .B(n140), .Z(n10013) );
  IV U10234 ( .A(n10013), .Z(n10193) );
  XOR U10235 ( .A(n10194), .B(n10193), .Z(n10102) );
  XOR U10236 ( .A(n10014), .B(n10102), .Z(n10104) );
  XOR U10237 ( .A(n10105), .B(n10104), .Z(n10202) );
  IV U10238 ( .A(n10015), .Z(n10016) );
  NOR U10239 ( .A(n10017), .B(n10016), .Z(n10021) );
  NOR U10240 ( .A(n10019), .B(n10018), .Z(n10020) );
  NOR U10241 ( .A(n10021), .B(n10020), .Z(n10200) );
  NOR U10242 ( .A(n143), .B(n136), .Z(n10198) );
  XOR U10243 ( .A(n10200), .B(n10198), .Z(n10201) );
  XOR U10244 ( .A(n10202), .B(n10201), .Z(n10096) );
  XOR U10245 ( .A(n10022), .B(n10096), .Z(n10098) );
  XOR U10246 ( .A(n10099), .B(n10098), .Z(n10207) );
  XOR U10247 ( .A(n10023), .B(n10207), .Z(n10209) );
  NOR U10248 ( .A(n147), .B(n132), .Z(n10024) );
  IV U10249 ( .A(n10024), .Z(n10208) );
  XOR U10250 ( .A(n10209), .B(n10208), .Z(n10090) );
  XOR U10251 ( .A(n10025), .B(n10090), .Z(n10092) );
  XOR U10252 ( .A(n10093), .B(n10092), .Z(n10215) );
  NOR U10253 ( .A(n150), .B(n129), .Z(n10213) );
  XOR U10254 ( .A(n10215), .B(n10213), .Z(n10216) );
  XOR U10255 ( .A(n10217), .B(n10216), .Z(n10084) );
  XOR U10256 ( .A(n10085), .B(n10084), .Z(n10026) );
  IV U10257 ( .A(n10026), .Z(n10086) );
  XOR U10258 ( .A(n10087), .B(n10086), .Z(n10081) );
  IV U10259 ( .A(n10027), .Z(n10028) );
  NOR U10260 ( .A(n10029), .B(n10028), .Z(n10033) );
  NOR U10261 ( .A(n10031), .B(n10030), .Z(n10032) );
  NOR U10262 ( .A(n10033), .B(n10032), .Z(n10079) );
  NOR U10263 ( .A(n155), .B(n124), .Z(n10077) );
  XOR U10264 ( .A(n10079), .B(n10077), .Z(n10080) );
  XOR U10265 ( .A(n10081), .B(n10080), .Z(n10071) );
  XOR U10266 ( .A(n10072), .B(n10071), .Z(n10034) );
  IV U10267 ( .A(n10034), .Z(n10073) );
  XOR U10268 ( .A(n10074), .B(n10073), .Z(n10066) );
  NOR U10269 ( .A(n158), .B(n121), .Z(n10064) );
  XOR U10270 ( .A(n10066), .B(n10064), .Z(n10067) );
  XOR U10271 ( .A(n10035), .B(n10067), .Z(n10059) );
  XOR U10272 ( .A(n10057), .B(n10059), .Z(n10060) );
  XOR U10273 ( .A(n10061), .B(n10060), .Z(n10051) );
  XOR U10274 ( .A(n10052), .B(n10051), .Z(n10036) );
  IV U10275 ( .A(n10036), .Z(n10053) );
  XOR U10276 ( .A(n10054), .B(n10053), .Z(n10045) );
  NOR U10277 ( .A(n165), .B(n42), .Z(n10043) );
  XOR U10278 ( .A(n10045), .B(n10043), .Z(n10048) );
  XOR U10279 ( .A(n10046), .B(n10048), .Z(n10038) );
  NOR U10280 ( .A(n10037), .B(n10038), .Z(n10042) );
  IV U10281 ( .A(n10037), .Z(n10039) );
  XOR U10282 ( .A(n10039), .B(n10038), .Z(n11904) );
  NOR U10283 ( .A(n167), .B(n44), .Z(n11905) );
  IV U10284 ( .A(n11905), .Z(n10040) );
  NOR U10285 ( .A(n11904), .B(n10040), .Z(n10041) );
  NOR U10286 ( .A(n10042), .B(n10041), .Z(n28634) );
  IV U10287 ( .A(n10043), .Z(n10044) );
  NOR U10288 ( .A(n10045), .B(n10044), .Z(n10050) );
  IV U10289 ( .A(n10046), .Z(n10047) );
  NOR U10290 ( .A(n10048), .B(n10047), .Z(n10049) );
  NOR U10291 ( .A(n10050), .B(n10049), .Z(n10231) );
  NOR U10292 ( .A(n167), .B(n42), .Z(n10227) );
  NOR U10293 ( .A(n10052), .B(n10051), .Z(n10056) );
  NOR U10294 ( .A(n10054), .B(n10053), .Z(n10055) );
  NOR U10295 ( .A(n10056), .B(n10055), .Z(n10409) );
  NOR U10296 ( .A(n165), .B(n43), .Z(n10406) );
  IV U10297 ( .A(n10057), .Z(n10058) );
  NOR U10298 ( .A(n10059), .B(n10058), .Z(n10063) );
  NOR U10299 ( .A(n10061), .B(n10060), .Z(n10062) );
  NOR U10300 ( .A(n10063), .B(n10062), .Z(n10238) );
  IV U10301 ( .A(n10238), .Z(n10225) );
  NOR U10302 ( .A(n163), .B(n118), .Z(n10234) );
  IV U10303 ( .A(n10064), .Z(n10065) );
  NOR U10304 ( .A(n10066), .B(n10065), .Z(n10070) );
  NOR U10305 ( .A(n10068), .B(n10067), .Z(n10069) );
  NOR U10306 ( .A(n10070), .B(n10069), .Z(n10402) );
  IV U10307 ( .A(n10402), .Z(n10224) );
  NOR U10308 ( .A(n10072), .B(n10071), .Z(n10076) );
  NOR U10309 ( .A(n10074), .B(n10073), .Z(n10075) );
  NOR U10310 ( .A(n10076), .B(n10075), .Z(n10244) );
  NOR U10311 ( .A(n158), .B(n122), .Z(n10242) );
  IV U10312 ( .A(n10242), .Z(n10223) );
  IV U10313 ( .A(n10077), .Z(n10078) );
  NOR U10314 ( .A(n10079), .B(n10078), .Z(n10083) );
  NOR U10315 ( .A(n10081), .B(n10080), .Z(n10082) );
  NOR U10316 ( .A(n10083), .B(n10082), .Z(n10391) );
  IV U10317 ( .A(n10391), .Z(n10221) );
  NOR U10318 ( .A(n10085), .B(n10084), .Z(n10089) );
  NOR U10319 ( .A(n10087), .B(n10086), .Z(n10088) );
  NOR U10320 ( .A(n10089), .B(n10088), .Z(n10250) );
  NOR U10321 ( .A(n155), .B(n127), .Z(n10248) );
  IV U10322 ( .A(n10248), .Z(n10220) );
  NOR U10323 ( .A(n10091), .B(n10090), .Z(n10095) );
  NOR U10324 ( .A(n10093), .B(n10092), .Z(n10094) );
  NOR U10325 ( .A(n10095), .B(n10094), .Z(n10256) );
  NOR U10326 ( .A(n150), .B(n130), .Z(n10254) );
  NOR U10327 ( .A(n10097), .B(n10096), .Z(n10101) );
  NOR U10328 ( .A(n10099), .B(n10098), .Z(n10100) );
  NOR U10329 ( .A(n10101), .B(n10100), .Z(n10262) );
  NOR U10330 ( .A(n147), .B(n134), .Z(n10260) );
  NOR U10331 ( .A(n10103), .B(n10102), .Z(n10107) );
  NOR U10332 ( .A(n10105), .B(n10104), .Z(n10106) );
  NOR U10333 ( .A(n10107), .B(n10106), .Z(n10268) );
  NOR U10334 ( .A(n143), .B(n138), .Z(n10266) );
  NOR U10335 ( .A(n10109), .B(n10108), .Z(n10113) );
  NOR U10336 ( .A(n10111), .B(n10110), .Z(n10112) );
  NOR U10337 ( .A(n10113), .B(n10112), .Z(n10275) );
  NOR U10338 ( .A(n139), .B(n142), .Z(n10273) );
  NOR U10339 ( .A(n137), .B(n144), .Z(n10282) );
  NOR U10340 ( .A(n10115), .B(n10114), .Z(n10119) );
  NOR U10341 ( .A(n10117), .B(n10116), .Z(n10118) );
  NOR U10342 ( .A(n10119), .B(n10118), .Z(n10278) );
  IV U10343 ( .A(n10120), .Z(n10121) );
  NOR U10344 ( .A(n10122), .B(n10121), .Z(n10126) );
  NOR U10345 ( .A(n10124), .B(n10123), .Z(n10125) );
  NOR U10346 ( .A(n10126), .B(n10125), .Z(n10290) );
  NOR U10347 ( .A(n135), .B(n146), .Z(n10287) );
  NOR U10348 ( .A(n133), .B(n149), .Z(n10297) );
  IV U10349 ( .A(n10127), .Z(n10129) );
  NOR U10350 ( .A(n10129), .B(n10128), .Z(n10133) );
  NOR U10351 ( .A(n10131), .B(n10130), .Z(n10132) );
  NOR U10352 ( .A(n10133), .B(n10132), .Z(n10294) );
  NOR U10353 ( .A(n10135), .B(n10134), .Z(n10140) );
  IV U10354 ( .A(n10136), .Z(n10137) );
  NOR U10355 ( .A(n10138), .B(n10137), .Z(n10139) );
  NOR U10356 ( .A(n10140), .B(n10139), .Z(n10305) );
  NOR U10357 ( .A(n131), .B(n151), .Z(n10302) );
  NOR U10358 ( .A(n10142), .B(n10141), .Z(n10146) );
  NOR U10359 ( .A(n10144), .B(n10143), .Z(n10145) );
  NOR U10360 ( .A(n10146), .B(n10145), .Z(n10311) );
  NOR U10361 ( .A(n126), .B(n154), .Z(n10309) );
  NOR U10362 ( .A(n10148), .B(n10147), .Z(n10152) );
  NOR U10363 ( .A(n10150), .B(n10149), .Z(n10151) );
  NOR U10364 ( .A(n10152), .B(n10151), .Z(n10317) );
  NOR U10365 ( .A(n123), .B(n159), .Z(n10315) );
  NOR U10366 ( .A(n10154), .B(n10153), .Z(n10158) );
  NOR U10367 ( .A(n10156), .B(n10155), .Z(n10157) );
  NOR U10368 ( .A(n10158), .B(n10157), .Z(n10323) );
  NOR U10369 ( .A(n119), .B(n162), .Z(n10321) );
  IV U10370 ( .A(n10321), .Z(n10167) );
  IV U10371 ( .A(n10159), .Z(n10160) );
  NOR U10372 ( .A(n10161), .B(n10160), .Z(n10165) );
  NOR U10373 ( .A(n10163), .B(n10162), .Z(n10164) );
  NOR U10374 ( .A(n10165), .B(n10164), .Z(n10328) );
  NOR U10375 ( .A(n164), .B(n79), .Z(n10326) );
  XOR U10376 ( .A(n10328), .B(n10326), .Z(n10330) );
  NOR U10377 ( .A(n166), .B(n117), .Z(n10166) );
  IV U10378 ( .A(n10166), .Z(n10329) );
  XOR U10379 ( .A(n10330), .B(n10329), .Z(n10320) );
  XOR U10380 ( .A(n10167), .B(n10320), .Z(n10322) );
  XOR U10381 ( .A(n10323), .B(n10322), .Z(n10339) );
  NOR U10382 ( .A(n10169), .B(n10168), .Z(n10173) );
  NOR U10383 ( .A(n10171), .B(n10170), .Z(n10172) );
  NOR U10384 ( .A(n10173), .B(n10172), .Z(n10337) );
  NOR U10385 ( .A(n120), .B(n160), .Z(n10335) );
  XOR U10386 ( .A(n10337), .B(n10335), .Z(n10338) );
  XOR U10387 ( .A(n10339), .B(n10338), .Z(n10314) );
  XOR U10388 ( .A(n10315), .B(n10314), .Z(n10174) );
  IV U10389 ( .A(n10174), .Z(n10316) );
  XOR U10390 ( .A(n10317), .B(n10316), .Z(n10347) );
  IV U10391 ( .A(n10175), .Z(n10176) );
  NOR U10392 ( .A(n10177), .B(n10176), .Z(n10181) );
  NOR U10393 ( .A(n10179), .B(n10178), .Z(n10180) );
  NOR U10394 ( .A(n10181), .B(n10180), .Z(n10345) );
  NOR U10395 ( .A(n125), .B(n157), .Z(n10343) );
  XOR U10396 ( .A(n10345), .B(n10343), .Z(n10346) );
  XOR U10397 ( .A(n10347), .B(n10346), .Z(n10308) );
  XOR U10398 ( .A(n10309), .B(n10308), .Z(n10182) );
  IV U10399 ( .A(n10182), .Z(n10310) );
  XOR U10400 ( .A(n10311), .B(n10310), .Z(n10355) );
  IV U10401 ( .A(n10183), .Z(n10184) );
  NOR U10402 ( .A(n10185), .B(n10184), .Z(n10189) );
  NOR U10403 ( .A(n10187), .B(n10186), .Z(n10188) );
  NOR U10404 ( .A(n10189), .B(n10188), .Z(n10353) );
  NOR U10405 ( .A(n128), .B(n152), .Z(n10351) );
  XOR U10406 ( .A(n10353), .B(n10351), .Z(n10354) );
  XOR U10407 ( .A(n10355), .B(n10354), .Z(n10301) );
  XOR U10408 ( .A(n10302), .B(n10301), .Z(n10303) );
  XOR U10409 ( .A(n10305), .B(n10303), .Z(n10293) );
  XOR U10410 ( .A(n10294), .B(n10293), .Z(n10295) );
  XOR U10411 ( .A(n10297), .B(n10295), .Z(n10286) );
  XOR U10412 ( .A(n10287), .B(n10286), .Z(n10288) );
  XOR U10413 ( .A(n10290), .B(n10288), .Z(n10279) );
  XOR U10414 ( .A(n10278), .B(n10279), .Z(n10281) );
  XOR U10415 ( .A(n10282), .B(n10281), .Z(n10271) );
  XOR U10416 ( .A(n10273), .B(n10271), .Z(n10274) );
  XOR U10417 ( .A(n10275), .B(n10274), .Z(n10363) );
  IV U10418 ( .A(n10190), .Z(n10191) );
  NOR U10419 ( .A(n10192), .B(n10191), .Z(n10196) );
  NOR U10420 ( .A(n10194), .B(n10193), .Z(n10195) );
  NOR U10421 ( .A(n10196), .B(n10195), .Z(n10361) );
  NOR U10422 ( .A(n141), .B(n140), .Z(n10359) );
  XOR U10423 ( .A(n10361), .B(n10359), .Z(n10362) );
  XOR U10424 ( .A(n10363), .B(n10362), .Z(n10265) );
  XOR U10425 ( .A(n10266), .B(n10265), .Z(n10197) );
  IV U10426 ( .A(n10197), .Z(n10267) );
  XOR U10427 ( .A(n10268), .B(n10267), .Z(n10371) );
  IV U10428 ( .A(n10198), .Z(n10199) );
  NOR U10429 ( .A(n10200), .B(n10199), .Z(n10204) );
  NOR U10430 ( .A(n10202), .B(n10201), .Z(n10203) );
  NOR U10431 ( .A(n10204), .B(n10203), .Z(n10369) );
  NOR U10432 ( .A(n145), .B(n136), .Z(n10367) );
  XOR U10433 ( .A(n10369), .B(n10367), .Z(n10370) );
  XOR U10434 ( .A(n10371), .B(n10370), .Z(n10259) );
  XOR U10435 ( .A(n10260), .B(n10259), .Z(n10205) );
  IV U10436 ( .A(n10205), .Z(n10261) );
  XOR U10437 ( .A(n10262), .B(n10261), .Z(n10379) );
  NOR U10438 ( .A(n10207), .B(n10206), .Z(n10211) );
  NOR U10439 ( .A(n10209), .B(n10208), .Z(n10210) );
  NOR U10440 ( .A(n10211), .B(n10210), .Z(n10377) );
  NOR U10441 ( .A(n148), .B(n132), .Z(n10375) );
  XOR U10442 ( .A(n10377), .B(n10375), .Z(n10378) );
  XOR U10443 ( .A(n10379), .B(n10378), .Z(n10253) );
  XOR U10444 ( .A(n10254), .B(n10253), .Z(n10212) );
  IV U10445 ( .A(n10212), .Z(n10255) );
  XOR U10446 ( .A(n10256), .B(n10255), .Z(n10387) );
  IV U10447 ( .A(n10213), .Z(n10214) );
  NOR U10448 ( .A(n10215), .B(n10214), .Z(n10219) );
  NOR U10449 ( .A(n10217), .B(n10216), .Z(n10218) );
  NOR U10450 ( .A(n10219), .B(n10218), .Z(n10385) );
  NOR U10451 ( .A(n153), .B(n129), .Z(n10383) );
  XOR U10452 ( .A(n10385), .B(n10383), .Z(n10386) );
  XOR U10453 ( .A(n10387), .B(n10386), .Z(n10247) );
  XOR U10454 ( .A(n10220), .B(n10247), .Z(n10249) );
  XOR U10455 ( .A(n10250), .B(n10249), .Z(n10392) );
  XOR U10456 ( .A(n10221), .B(n10392), .Z(n10394) );
  NOR U10457 ( .A(n156), .B(n124), .Z(n10222) );
  IV U10458 ( .A(n10222), .Z(n10393) );
  XOR U10459 ( .A(n10394), .B(n10393), .Z(n10241) );
  XOR U10460 ( .A(n10223), .B(n10241), .Z(n10243) );
  XOR U10461 ( .A(n10244), .B(n10243), .Z(n10400) );
  NOR U10462 ( .A(n161), .B(n121), .Z(n10398) );
  XOR U10463 ( .A(n10400), .B(n10398), .Z(n10401) );
  XOR U10464 ( .A(n10224), .B(n10401), .Z(n10236) );
  XOR U10465 ( .A(n10234), .B(n10236), .Z(n10237) );
  XOR U10466 ( .A(n10225), .B(n10237), .Z(n10408) );
  XOR U10467 ( .A(n10406), .B(n10408), .Z(n10410) );
  XOR U10468 ( .A(n10409), .B(n10410), .Z(n10229) );
  XOR U10469 ( .A(n10227), .B(n10229), .Z(n10230) );
  XOR U10470 ( .A(n10231), .B(n10230), .Z(n10226) );
  IV U10471 ( .A(n10226), .Z(n28633) );
  NOR U10472 ( .A(n28634), .B(n28633), .Z(n31686) );
  IV U10473 ( .A(n31686), .Z(n10414) );
  IV U10474 ( .A(n10227), .Z(n10228) );
  NOR U10475 ( .A(n10229), .B(n10228), .Z(n10233) );
  NOR U10476 ( .A(n10231), .B(n10230), .Z(n10232) );
  NOR U10477 ( .A(n10233), .B(n10232), .Z(n28650) );
  IV U10478 ( .A(n10234), .Z(n10235) );
  NOR U10479 ( .A(n10236), .B(n10235), .Z(n10240) );
  NOR U10480 ( .A(n10238), .B(n10237), .Z(n10239) );
  NOR U10481 ( .A(n10240), .B(n10239), .Z(n28663) );
  NOR U10482 ( .A(n165), .B(n118), .Z(n28659) );
  NOR U10483 ( .A(n10242), .B(n10241), .Z(n10246) );
  NOR U10484 ( .A(n10244), .B(n10243), .Z(n10245) );
  NOR U10485 ( .A(n10246), .B(n10245), .Z(n28669) );
  NOR U10486 ( .A(n161), .B(n122), .Z(n28666) );
  NOR U10487 ( .A(n10248), .B(n10247), .Z(n10252) );
  NOR U10488 ( .A(n10250), .B(n10249), .Z(n10251) );
  NOR U10489 ( .A(n10252), .B(n10251), .Z(n28677) );
  NOR U10490 ( .A(n156), .B(n127), .Z(n28674) );
  NOR U10491 ( .A(n10254), .B(n10253), .Z(n10258) );
  NOR U10492 ( .A(n10256), .B(n10255), .Z(n10257) );
  NOR U10493 ( .A(n10258), .B(n10257), .Z(n28685) );
  NOR U10494 ( .A(n153), .B(n130), .Z(n28682) );
  NOR U10495 ( .A(n10260), .B(n10259), .Z(n10264) );
  NOR U10496 ( .A(n10262), .B(n10261), .Z(n10263) );
  NOR U10497 ( .A(n10264), .B(n10263), .Z(n28693) );
  NOR U10498 ( .A(n148), .B(n134), .Z(n28690) );
  NOR U10499 ( .A(n10266), .B(n10265), .Z(n10270) );
  NOR U10500 ( .A(n10268), .B(n10267), .Z(n10269) );
  NOR U10501 ( .A(n10270), .B(n10269), .Z(n28701) );
  NOR U10502 ( .A(n145), .B(n138), .Z(n28698) );
  IV U10503 ( .A(n10271), .Z(n10272) );
  NOR U10504 ( .A(n10273), .B(n10272), .Z(n10277) );
  NOR U10505 ( .A(n10275), .B(n10274), .Z(n10276) );
  NOR U10506 ( .A(n10277), .B(n10276), .Z(n28788) );
  NOR U10507 ( .A(n139), .B(n144), .Z(n28707) );
  IV U10508 ( .A(n10278), .Z(n10280) );
  NOR U10509 ( .A(n10280), .B(n10279), .Z(n10284) );
  NOR U10510 ( .A(n10282), .B(n10281), .Z(n10283) );
  NOR U10511 ( .A(n10284), .B(n10283), .Z(n28706) );
  XOR U10512 ( .A(n28707), .B(n28706), .Z(n10285) );
  IV U10513 ( .A(n10285), .Z(n28709) );
  NOR U10514 ( .A(n10287), .B(n10286), .Z(n10292) );
  IV U10515 ( .A(n10288), .Z(n10289) );
  NOR U10516 ( .A(n10290), .B(n10289), .Z(n10291) );
  NOR U10517 ( .A(n10292), .B(n10291), .Z(n28717) );
  NOR U10518 ( .A(n137), .B(n146), .Z(n28714) );
  NOR U10519 ( .A(n10294), .B(n10293), .Z(n10299) );
  IV U10520 ( .A(n10295), .Z(n10296) );
  NOR U10521 ( .A(n10297), .B(n10296), .Z(n10298) );
  NOR U10522 ( .A(n10299), .B(n10298), .Z(n10300) );
  IV U10523 ( .A(n10300), .Z(n28779) );
  NOR U10524 ( .A(n135), .B(n149), .Z(n28777) );
  XOR U10525 ( .A(n28779), .B(n28777), .Z(n28781) );
  NOR U10526 ( .A(n10302), .B(n10301), .Z(n10307) );
  IV U10527 ( .A(n10303), .Z(n10304) );
  NOR U10528 ( .A(n10305), .B(n10304), .Z(n10306) );
  NOR U10529 ( .A(n10307), .B(n10306), .Z(n28723) );
  NOR U10530 ( .A(n133), .B(n151), .Z(n28720) );
  NOR U10531 ( .A(n10309), .B(n10308), .Z(n10313) );
  NOR U10532 ( .A(n10311), .B(n10310), .Z(n10312) );
  NOR U10533 ( .A(n10313), .B(n10312), .Z(n28731) );
  NOR U10534 ( .A(n128), .B(n154), .Z(n28728) );
  NOR U10535 ( .A(n10315), .B(n10314), .Z(n10319) );
  NOR U10536 ( .A(n10317), .B(n10316), .Z(n10318) );
  NOR U10537 ( .A(n10319), .B(n10318), .Z(n28739) );
  NOR U10538 ( .A(n125), .B(n159), .Z(n28737) );
  IV U10539 ( .A(n28737), .Z(n10342) );
  NOR U10540 ( .A(n10321), .B(n10320), .Z(n10325) );
  NOR U10541 ( .A(n10323), .B(n10322), .Z(n10324) );
  NOR U10542 ( .A(n10325), .B(n10324), .Z(n28745) );
  NOR U10543 ( .A(n120), .B(n162), .Z(n28743) );
  IV U10544 ( .A(n28743), .Z(n10334) );
  NOR U10545 ( .A(n164), .B(n119), .Z(n28748) );
  IV U10546 ( .A(n10326), .Z(n10327) );
  NOR U10547 ( .A(n10328), .B(n10327), .Z(n10332) );
  NOR U10548 ( .A(n10330), .B(n10329), .Z(n10331) );
  NOR U10549 ( .A(n10332), .B(n10331), .Z(n28749) );
  XOR U10550 ( .A(n28748), .B(n28749), .Z(n28751) );
  NOR U10551 ( .A(n166), .B(n79), .Z(n10333) );
  IV U10552 ( .A(n10333), .Z(n28750) );
  XOR U10553 ( .A(n28751), .B(n28750), .Z(n28742) );
  XOR U10554 ( .A(n10334), .B(n28742), .Z(n28744) );
  XOR U10555 ( .A(n28745), .B(n28744), .Z(n28759) );
  IV U10556 ( .A(n10335), .Z(n10336) );
  NOR U10557 ( .A(n10337), .B(n10336), .Z(n10341) );
  NOR U10558 ( .A(n10339), .B(n10338), .Z(n10340) );
  NOR U10559 ( .A(n10341), .B(n10340), .Z(n28757) );
  NOR U10560 ( .A(n123), .B(n160), .Z(n28755) );
  XOR U10561 ( .A(n28757), .B(n28755), .Z(n28758) );
  XOR U10562 ( .A(n28759), .B(n28758), .Z(n28736) );
  XOR U10563 ( .A(n10342), .B(n28736), .Z(n28738) );
  XOR U10564 ( .A(n28739), .B(n28738), .Z(n28767) );
  IV U10565 ( .A(n28767), .Z(n10350) );
  IV U10566 ( .A(n10343), .Z(n10344) );
  NOR U10567 ( .A(n10345), .B(n10344), .Z(n10349) );
  NOR U10568 ( .A(n10347), .B(n10346), .Z(n10348) );
  NOR U10569 ( .A(n10349), .B(n10348), .Z(n28765) );
  NOR U10570 ( .A(n126), .B(n157), .Z(n28763) );
  XOR U10571 ( .A(n28765), .B(n28763), .Z(n28766) );
  XOR U10572 ( .A(n10350), .B(n28766), .Z(n28730) );
  XOR U10573 ( .A(n28728), .B(n28730), .Z(n28732) );
  XOR U10574 ( .A(n28731), .B(n28732), .Z(n28773) );
  IV U10575 ( .A(n10351), .Z(n10352) );
  NOR U10576 ( .A(n10353), .B(n10352), .Z(n10357) );
  NOR U10577 ( .A(n10355), .B(n10354), .Z(n10356) );
  NOR U10578 ( .A(n10357), .B(n10356), .Z(n28772) );
  NOR U10579 ( .A(n131), .B(n152), .Z(n28770) );
  XOR U10580 ( .A(n28772), .B(n28770), .Z(n28774) );
  XOR U10581 ( .A(n28773), .B(n28774), .Z(n10358) );
  IV U10582 ( .A(n10358), .Z(n28722) );
  XOR U10583 ( .A(n28720), .B(n28722), .Z(n28725) );
  XOR U10584 ( .A(n28723), .B(n28725), .Z(n28780) );
  XOR U10585 ( .A(n28781), .B(n28780), .Z(n28713) );
  XOR U10586 ( .A(n28714), .B(n28713), .Z(n28715) );
  XOR U10587 ( .A(n28717), .B(n28715), .Z(n28708) );
  XOR U10588 ( .A(n28709), .B(n28708), .Z(n28787) );
  NOR U10589 ( .A(n141), .B(n142), .Z(n28785) );
  XOR U10590 ( .A(n28787), .B(n28785), .Z(n28790) );
  XOR U10591 ( .A(n28788), .B(n28790), .Z(n28797) );
  IV U10592 ( .A(n10359), .Z(n10360) );
  NOR U10593 ( .A(n10361), .B(n10360), .Z(n10365) );
  NOR U10594 ( .A(n10363), .B(n10362), .Z(n10364) );
  NOR U10595 ( .A(n10365), .B(n10364), .Z(n28795) );
  NOR U10596 ( .A(n143), .B(n140), .Z(n28793) );
  XOR U10597 ( .A(n28795), .B(n28793), .Z(n28796) );
  XOR U10598 ( .A(n28797), .B(n28796), .Z(n10366) );
  IV U10599 ( .A(n10366), .Z(n28700) );
  XOR U10600 ( .A(n28698), .B(n28700), .Z(n28703) );
  XOR U10601 ( .A(n28701), .B(n28703), .Z(n28803) );
  IV U10602 ( .A(n10367), .Z(n10368) );
  NOR U10603 ( .A(n10369), .B(n10368), .Z(n10373) );
  NOR U10604 ( .A(n10371), .B(n10370), .Z(n10372) );
  NOR U10605 ( .A(n10373), .B(n10372), .Z(n28802) );
  NOR U10606 ( .A(n147), .B(n136), .Z(n28800) );
  XOR U10607 ( .A(n28802), .B(n28800), .Z(n28804) );
  XOR U10608 ( .A(n28803), .B(n28804), .Z(n10374) );
  IV U10609 ( .A(n10374), .Z(n28692) );
  XOR U10610 ( .A(n28690), .B(n28692), .Z(n28695) );
  XOR U10611 ( .A(n28693), .B(n28695), .Z(n28811) );
  IV U10612 ( .A(n10375), .Z(n10376) );
  NOR U10613 ( .A(n10377), .B(n10376), .Z(n10381) );
  NOR U10614 ( .A(n10379), .B(n10378), .Z(n10380) );
  NOR U10615 ( .A(n10381), .B(n10380), .Z(n28809) );
  NOR U10616 ( .A(n150), .B(n132), .Z(n28807) );
  XOR U10617 ( .A(n28809), .B(n28807), .Z(n28810) );
  XOR U10618 ( .A(n28811), .B(n28810), .Z(n10382) );
  IV U10619 ( .A(n10382), .Z(n28684) );
  XOR U10620 ( .A(n28682), .B(n28684), .Z(n28687) );
  XOR U10621 ( .A(n28685), .B(n28687), .Z(n28818) );
  IV U10622 ( .A(n10383), .Z(n10384) );
  NOR U10623 ( .A(n10385), .B(n10384), .Z(n10389) );
  NOR U10624 ( .A(n10387), .B(n10386), .Z(n10388) );
  NOR U10625 ( .A(n10389), .B(n10388), .Z(n28816) );
  NOR U10626 ( .A(n155), .B(n129), .Z(n28814) );
  XOR U10627 ( .A(n28816), .B(n28814), .Z(n28817) );
  XOR U10628 ( .A(n28818), .B(n28817), .Z(n10390) );
  IV U10629 ( .A(n10390), .Z(n28676) );
  XOR U10630 ( .A(n28674), .B(n28676), .Z(n28679) );
  XOR U10631 ( .A(n28677), .B(n28679), .Z(n28825) );
  NOR U10632 ( .A(n10392), .B(n10391), .Z(n10396) );
  NOR U10633 ( .A(n10394), .B(n10393), .Z(n10395) );
  NOR U10634 ( .A(n10396), .B(n10395), .Z(n28823) );
  NOR U10635 ( .A(n158), .B(n124), .Z(n28821) );
  XOR U10636 ( .A(n28823), .B(n28821), .Z(n28824) );
  XOR U10637 ( .A(n28825), .B(n28824), .Z(n10397) );
  IV U10638 ( .A(n10397), .Z(n28668) );
  XOR U10639 ( .A(n28666), .B(n28668), .Z(n28671) );
  XOR U10640 ( .A(n28669), .B(n28671), .Z(n28831) );
  IV U10641 ( .A(n28831), .Z(n10405) );
  IV U10642 ( .A(n10398), .Z(n10399) );
  NOR U10643 ( .A(n10400), .B(n10399), .Z(n10404) );
  NOR U10644 ( .A(n10402), .B(n10401), .Z(n10403) );
  NOR U10645 ( .A(n10404), .B(n10403), .Z(n28830) );
  NOR U10646 ( .A(n163), .B(n121), .Z(n28828) );
  XOR U10647 ( .A(n28830), .B(n28828), .Z(n28832) );
  XOR U10648 ( .A(n10405), .B(n28832), .Z(n28661) );
  XOR U10649 ( .A(n28659), .B(n28661), .Z(n28662) );
  XOR U10650 ( .A(n28663), .B(n28662), .Z(n28654) );
  IV U10651 ( .A(n10406), .Z(n10407) );
  NOR U10652 ( .A(n10408), .B(n10407), .Z(n10413) );
  IV U10653 ( .A(n10409), .Z(n10411) );
  NOR U10654 ( .A(n10411), .B(n10410), .Z(n10412) );
  NOR U10655 ( .A(n10413), .B(n10412), .Z(n28653) );
  NOR U10656 ( .A(n167), .B(n43), .Z(n28651) );
  XOR U10657 ( .A(n28653), .B(n28651), .Z(n28656) );
  XOR U10658 ( .A(n28654), .B(n28656), .Z(n28649) );
  XOR U10659 ( .A(n28650), .B(n28649), .Z(n28640) );
  IV U10660 ( .A(n28640), .Z(n31685) );
  NOR U10661 ( .A(n10414), .B(n31685), .Z(n28648) );
  NOR U10662 ( .A(n163), .B(n45), .Z(n10892) );
  XOR U10663 ( .A(n10416), .B(n10415), .Z(n10869) );
  NOR U10664 ( .A(n156), .B(n45), .Z(n10870) );
  IV U10665 ( .A(n10870), .Z(n10417) );
  NOR U10666 ( .A(n10869), .B(n10417), .Z(n10872) );
  XOR U10667 ( .A(n10419), .B(n10418), .Z(n10857) );
  NOR U10668 ( .A(n153), .B(n45), .Z(n10858) );
  IV U10669 ( .A(n10858), .Z(n10420) );
  NOR U10670 ( .A(n10857), .B(n10420), .Z(n10860) );
  XOR U10671 ( .A(n10422), .B(n10421), .Z(n10838) );
  NOR U10672 ( .A(n147), .B(n45), .Z(n10839) );
  IV U10673 ( .A(n10839), .Z(n10423) );
  NOR U10674 ( .A(n10838), .B(n10423), .Z(n10841) );
  XOR U10675 ( .A(n10425), .B(n10424), .Z(n10787) );
  NOR U10676 ( .A(n133), .B(n45), .Z(n10788) );
  IV U10677 ( .A(n10788), .Z(n10426) );
  NOR U10678 ( .A(n10787), .B(n10426), .Z(n10790) );
  NOR U10679 ( .A(n128), .B(n45), .Z(n10430) );
  XOR U10680 ( .A(n10428), .B(n10427), .Z(n10429) );
  NOR U10681 ( .A(n10430), .B(n10429), .Z(n10777) );
  XOR U10682 ( .A(n10430), .B(n10429), .Z(n11254) );
  IV U10683 ( .A(n11254), .Z(n10775) );
  NOR U10684 ( .A(n117), .B(n45), .Z(n10720) );
  XOR U10685 ( .A(n10432), .B(n10431), .Z(n10714) );
  NOR U10686 ( .A(n82), .B(n45), .Z(n10438) );
  XOR U10687 ( .A(n10434), .B(n10433), .Z(n10435) );
  XOR U10688 ( .A(n10436), .B(n10435), .Z(n11170) );
  IV U10689 ( .A(n11170), .Z(n10437) );
  NOR U10690 ( .A(n10438), .B(n10437), .Z(n10689) );
  IV U10691 ( .A(n10438), .Z(n11171) );
  NOR U10692 ( .A(n11171), .B(n11170), .Z(n10687) );
  XOR U10693 ( .A(n10440), .B(n10439), .Z(n10655) );
  IV U10694 ( .A(n10655), .Z(n11141) );
  NOR U10695 ( .A(n84), .B(n45), .Z(n10654) );
  IV U10696 ( .A(n10654), .Z(n11140) );
  NOR U10697 ( .A(n11141), .B(n11140), .Z(n10658) );
  NOR U10698 ( .A(n112), .B(n45), .Z(n10441) );
  IV U10699 ( .A(n10441), .Z(n10651) );
  NOR U10700 ( .A(n85), .B(n45), .Z(n10444) );
  XOR U10701 ( .A(n10443), .B(n10442), .Z(n10445) );
  NOR U10702 ( .A(n10444), .B(n10445), .Z(n10644) );
  IV U10703 ( .A(n10444), .Z(n11127) );
  IV U10704 ( .A(n10445), .Z(n11126) );
  NOR U10705 ( .A(n11127), .B(n11126), .Z(n10642) );
  NOR U10706 ( .A(n111), .B(n45), .Z(n10446) );
  IV U10707 ( .A(n10446), .Z(n10638) );
  NOR U10708 ( .A(n86), .B(n45), .Z(n10627) );
  XOR U10709 ( .A(n10448), .B(n10447), .Z(n10628) );
  NOR U10710 ( .A(n10627), .B(n10628), .Z(n10631) );
  XOR U10711 ( .A(n10450), .B(n10449), .Z(n10622) );
  NOR U10712 ( .A(n110), .B(n45), .Z(n10623) );
  NOR U10713 ( .A(n10622), .B(n10623), .Z(n10626) );
  NOR U10714 ( .A(n109), .B(n45), .Z(n10618) );
  XOR U10715 ( .A(n10452), .B(n10451), .Z(n10617) );
  NOR U10716 ( .A(n10618), .B(n10617), .Z(n10621) );
  XOR U10717 ( .A(n10454), .B(n10453), .Z(n10455) );
  NOR U10718 ( .A(n87), .B(n45), .Z(n10456) );
  NOR U10719 ( .A(n10455), .B(n10456), .Z(n10606) );
  IV U10720 ( .A(n10455), .Z(n11090) );
  IV U10721 ( .A(n10456), .Z(n11089) );
  NOR U10722 ( .A(n11090), .B(n11089), .Z(n10604) );
  NOR U10723 ( .A(n88), .B(n45), .Z(n10590) );
  XOR U10724 ( .A(n10458), .B(n10457), .Z(n10589) );
  NOR U10725 ( .A(n10590), .B(n10589), .Z(n10593) );
  NOR U10726 ( .A(n106), .B(n45), .Z(n10585) );
  XOR U10727 ( .A(n10460), .B(n10459), .Z(n10584) );
  NOR U10728 ( .A(n10585), .B(n10584), .Z(n10588) );
  NOR U10729 ( .A(n105), .B(n45), .Z(n10580) );
  XOR U10730 ( .A(n10462), .B(n10461), .Z(n10579) );
  NOR U10731 ( .A(n10580), .B(n10579), .Z(n10583) );
  XOR U10732 ( .A(n10464), .B(n10463), .Z(n10567) );
  IV U10733 ( .A(n10567), .Z(n10952) );
  NOR U10734 ( .A(n89), .B(n45), .Z(n10566) );
  IV U10735 ( .A(n10566), .Z(n10951) );
  NOR U10736 ( .A(n10952), .B(n10951), .Z(n10570) );
  XOR U10737 ( .A(n10466), .B(n10465), .Z(n10467) );
  XOR U10738 ( .A(n10468), .B(n10467), .Z(n10562) );
  NOR U10739 ( .A(n103), .B(n45), .Z(n10561) );
  IV U10740 ( .A(n10561), .Z(n10469) );
  NOR U10741 ( .A(n10562), .B(n10469), .Z(n10565) );
  NOR U10742 ( .A(n90), .B(n45), .Z(n10556) );
  XOR U10743 ( .A(n10471), .B(n10470), .Z(n10557) );
  NOR U10744 ( .A(n10556), .B(n10557), .Z(n10560) );
  NOR U10745 ( .A(n102), .B(n45), .Z(n10552) );
  XOR U10746 ( .A(n10473), .B(n10472), .Z(n10553) );
  IV U10747 ( .A(n10553), .Z(n10474) );
  NOR U10748 ( .A(n10552), .B(n10474), .Z(n10555) );
  NOR U10749 ( .A(n101), .B(n45), .Z(n10478) );
  XOR U10750 ( .A(n10476), .B(n10475), .Z(n10477) );
  NOR U10751 ( .A(n10478), .B(n10477), .Z(n10551) );
  XOR U10752 ( .A(n10478), .B(n10477), .Z(n10479) );
  IV U10753 ( .A(n10479), .Z(n11042) );
  NOR U10754 ( .A(n99), .B(n45), .Z(n10482) );
  XOR U10755 ( .A(n10481), .B(n10480), .Z(n10972) );
  NOR U10756 ( .A(n10482), .B(n10972), .Z(n10539) );
  IV U10757 ( .A(n10482), .Z(n10970) );
  IV U10758 ( .A(n10972), .Z(n10483) );
  NOR U10759 ( .A(n10970), .B(n10483), .Z(n10537) );
  XOR U10760 ( .A(n10485), .B(n10484), .Z(n10486) );
  XOR U10761 ( .A(n10487), .B(n10486), .Z(n10533) );
  NOR U10762 ( .A(n98), .B(n45), .Z(n10532) );
  IV U10763 ( .A(n10532), .Z(n10488) );
  NOR U10764 ( .A(n10533), .B(n10488), .Z(n10535) );
  IV U10765 ( .A(n10489), .Z(n10491) );
  XOR U10766 ( .A(n10491), .B(n10490), .Z(n10528) );
  NOR U10767 ( .A(n91), .B(n45), .Z(n10529) );
  IV U10768 ( .A(n10529), .Z(n10492) );
  NOR U10769 ( .A(n10528), .B(n10492), .Z(n10531) );
  IV U10770 ( .A(n10493), .Z(n10495) );
  XOR U10771 ( .A(n10495), .B(n10494), .Z(n10516) );
  NOR U10772 ( .A(n96), .B(n45), .Z(n10517) );
  IV U10773 ( .A(n10517), .Z(n10496) );
  NOR U10774 ( .A(n10516), .B(n10496), .Z(n10519) );
  NOR U10775 ( .A(n95), .B(n45), .Z(n10513) );
  IV U10776 ( .A(n10513), .Z(n10499) );
  XOR U10777 ( .A(n10498), .B(n10497), .Z(n10512) );
  NOR U10778 ( .A(n10499), .B(n10512), .Z(n10515) );
  NOR U10779 ( .A(n93), .B(n45), .Z(n11491) );
  IV U10780 ( .A(n11491), .Z(n10500) );
  NOR U10781 ( .A(n44), .B(n168), .Z(n10508) );
  IV U10782 ( .A(n10508), .Z(n10503) );
  NOR U10783 ( .A(n10500), .B(n10503), .Z(n10501) );
  IV U10784 ( .A(n10501), .Z(n10502) );
  NOR U10785 ( .A(n94), .B(n10502), .Z(n10511) );
  NOR U10786 ( .A(n10503), .B(n93), .Z(n10504) );
  XOR U10787 ( .A(n94), .B(n10504), .Z(n10505) );
  NOR U10788 ( .A(n45), .B(n10505), .Z(n10506) );
  IV U10789 ( .A(n10506), .Z(n10992) );
  XOR U10790 ( .A(n10508), .B(n10507), .Z(n10991) );
  IV U10791 ( .A(n10991), .Z(n10509) );
  NOR U10792 ( .A(n10992), .B(n10509), .Z(n10510) );
  NOR U10793 ( .A(n10511), .B(n10510), .Z(n10987) );
  XOR U10794 ( .A(n10513), .B(n10512), .Z(n10988) );
  NOR U10795 ( .A(n10987), .B(n10988), .Z(n10514) );
  NOR U10796 ( .A(n10515), .B(n10514), .Z(n10983) );
  XOR U10797 ( .A(n10517), .B(n10516), .Z(n10984) );
  NOR U10798 ( .A(n10983), .B(n10984), .Z(n10518) );
  NOR U10799 ( .A(n10519), .B(n10518), .Z(n10522) );
  NOR U10800 ( .A(n97), .B(n45), .Z(n10521) );
  IV U10801 ( .A(n10521), .Z(n10520) );
  NOR U10802 ( .A(n10522), .B(n10520), .Z(n10527) );
  XOR U10803 ( .A(n10522), .B(n10521), .Z(n10980) );
  XOR U10804 ( .A(n10524), .B(n10523), .Z(n10981) );
  IV U10805 ( .A(n10981), .Z(n10525) );
  NOR U10806 ( .A(n10980), .B(n10525), .Z(n10526) );
  NOR U10807 ( .A(n10527), .B(n10526), .Z(n10976) );
  XOR U10808 ( .A(n10529), .B(n10528), .Z(n10977) );
  NOR U10809 ( .A(n10976), .B(n10977), .Z(n10530) );
  NOR U10810 ( .A(n10531), .B(n10530), .Z(n10975) );
  XOR U10811 ( .A(n10533), .B(n10532), .Z(n10974) );
  NOR U10812 ( .A(n10975), .B(n10974), .Z(n10534) );
  NOR U10813 ( .A(n10535), .B(n10534), .Z(n10536) );
  IV U10814 ( .A(n10536), .Z(n10969) );
  NOR U10815 ( .A(n10537), .B(n10969), .Z(n10538) );
  NOR U10816 ( .A(n10539), .B(n10538), .Z(n10546) );
  IV U10817 ( .A(n10546), .Z(n10541) );
  NOR U10818 ( .A(n100), .B(n45), .Z(n10540) );
  IV U10819 ( .A(n10540), .Z(n10545) );
  NOR U10820 ( .A(n10541), .B(n10545), .Z(n10548) );
  XOR U10821 ( .A(n10543), .B(n10542), .Z(n10544) );
  IV U10822 ( .A(n10544), .Z(n10965) );
  XOR U10823 ( .A(n10546), .B(n10545), .Z(n10966) );
  NOR U10824 ( .A(n10965), .B(n10966), .Z(n10547) );
  NOR U10825 ( .A(n10548), .B(n10547), .Z(n10549) );
  IV U10826 ( .A(n10549), .Z(n11041) );
  NOR U10827 ( .A(n11042), .B(n11041), .Z(n10550) );
  NOR U10828 ( .A(n10551), .B(n10550), .Z(n10963) );
  XOR U10829 ( .A(n10553), .B(n10552), .Z(n10962) );
  NOR U10830 ( .A(n10963), .B(n10962), .Z(n10554) );
  NOR U10831 ( .A(n10555), .B(n10554), .Z(n10960) );
  IV U10832 ( .A(n10556), .Z(n10558) );
  XOR U10833 ( .A(n10558), .B(n10557), .Z(n10959) );
  NOR U10834 ( .A(n10960), .B(n10959), .Z(n10559) );
  NOR U10835 ( .A(n10560), .B(n10559), .Z(n10957) );
  IV U10836 ( .A(n10957), .Z(n10563) );
  XOR U10837 ( .A(n10562), .B(n10561), .Z(n10956) );
  NOR U10838 ( .A(n10563), .B(n10956), .Z(n10564) );
  NOR U10839 ( .A(n10565), .B(n10564), .Z(n10954) );
  NOR U10840 ( .A(n10567), .B(n10566), .Z(n10568) );
  NOR U10841 ( .A(n10954), .B(n10568), .Z(n10569) );
  NOR U10842 ( .A(n10570), .B(n10569), .Z(n10575) );
  NOR U10843 ( .A(n104), .B(n45), .Z(n10574) );
  IV U10844 ( .A(n10574), .Z(n10571) );
  NOR U10845 ( .A(n10575), .B(n10571), .Z(n10577) );
  XOR U10846 ( .A(n10573), .B(n10572), .Z(n10950) );
  XOR U10847 ( .A(n10575), .B(n10574), .Z(n10949) );
  NOR U10848 ( .A(n10950), .B(n10949), .Z(n10576) );
  NOR U10849 ( .A(n10577), .B(n10576), .Z(n10578) );
  IV U10850 ( .A(n10578), .Z(n11070) );
  XOR U10851 ( .A(n10580), .B(n10579), .Z(n10581) );
  IV U10852 ( .A(n10581), .Z(n11069) );
  NOR U10853 ( .A(n11070), .B(n11069), .Z(n10582) );
  NOR U10854 ( .A(n10583), .B(n10582), .Z(n10946) );
  XOR U10855 ( .A(n10585), .B(n10584), .Z(n10945) );
  IV U10856 ( .A(n10945), .Z(n10586) );
  NOR U10857 ( .A(n10946), .B(n10586), .Z(n10587) );
  NOR U10858 ( .A(n10588), .B(n10587), .Z(n11079) );
  XOR U10859 ( .A(n10590), .B(n10589), .Z(n11080) );
  IV U10860 ( .A(n11080), .Z(n10591) );
  NOR U10861 ( .A(n11079), .B(n10591), .Z(n10592) );
  NOR U10862 ( .A(n10593), .B(n10592), .Z(n10594) );
  IV U10863 ( .A(n10594), .Z(n10599) );
  NOR U10864 ( .A(n107), .B(n45), .Z(n10598) );
  IV U10865 ( .A(n10598), .Z(n10595) );
  NOR U10866 ( .A(n10599), .B(n10595), .Z(n10602) );
  XOR U10867 ( .A(n10597), .B(n10596), .Z(n10940) );
  IV U10868 ( .A(n10940), .Z(n10600) );
  XOR U10869 ( .A(n10599), .B(n10598), .Z(n10941) );
  NOR U10870 ( .A(n10600), .B(n10941), .Z(n10601) );
  NOR U10871 ( .A(n10602), .B(n10601), .Z(n11092) );
  IV U10872 ( .A(n11092), .Z(n10603) );
  NOR U10873 ( .A(n10604), .B(n10603), .Z(n10605) );
  NOR U10874 ( .A(n10606), .B(n10605), .Z(n10610) );
  IV U10875 ( .A(n10610), .Z(n10608) );
  NOR U10876 ( .A(n108), .B(n45), .Z(n10607) );
  IV U10877 ( .A(n10607), .Z(n10609) );
  NOR U10878 ( .A(n10608), .B(n10609), .Z(n10615) );
  XOR U10879 ( .A(n10610), .B(n10609), .Z(n10939) );
  XOR U10880 ( .A(n10612), .B(n10611), .Z(n10613) );
  IV U10881 ( .A(n10613), .Z(n10938) );
  NOR U10882 ( .A(n10939), .B(n10938), .Z(n10614) );
  NOR U10883 ( .A(n10615), .B(n10614), .Z(n10616) );
  IV U10884 ( .A(n10616), .Z(n11104) );
  XOR U10885 ( .A(n10618), .B(n10617), .Z(n10619) );
  IV U10886 ( .A(n10619), .Z(n11103) );
  NOR U10887 ( .A(n11104), .B(n11103), .Z(n10620) );
  NOR U10888 ( .A(n10621), .B(n10620), .Z(n10934) );
  XOR U10889 ( .A(n10623), .B(n10622), .Z(n10624) );
  IV U10890 ( .A(n10624), .Z(n10935) );
  NOR U10891 ( .A(n10934), .B(n10935), .Z(n10625) );
  NOR U10892 ( .A(n10626), .B(n10625), .Z(n11116) );
  IV U10893 ( .A(n10627), .Z(n11114) );
  IV U10894 ( .A(n10628), .Z(n11113) );
  NOR U10895 ( .A(n11114), .B(n11113), .Z(n10629) );
  NOR U10896 ( .A(n11116), .B(n10629), .Z(n10630) );
  NOR U10897 ( .A(n10631), .B(n10630), .Z(n10637) );
  IV U10898 ( .A(n10637), .Z(n10632) );
  NOR U10899 ( .A(n10638), .B(n10632), .Z(n10640) );
  XOR U10900 ( .A(n10634), .B(n10633), .Z(n10635) );
  XOR U10901 ( .A(n10636), .B(n10635), .Z(n10930) );
  XOR U10902 ( .A(n10638), .B(n10637), .Z(n10931) );
  NOR U10903 ( .A(n10930), .B(n10931), .Z(n10639) );
  NOR U10904 ( .A(n10640), .B(n10639), .Z(n11129) );
  IV U10905 ( .A(n11129), .Z(n10641) );
  NOR U10906 ( .A(n10642), .B(n10641), .Z(n10643) );
  NOR U10907 ( .A(n10644), .B(n10643), .Z(n10650) );
  IV U10908 ( .A(n10650), .Z(n10645) );
  NOR U10909 ( .A(n10651), .B(n10645), .Z(n10653) );
  XOR U10910 ( .A(n10647), .B(n10646), .Z(n10648) );
  XOR U10911 ( .A(n10649), .B(n10648), .Z(n10925) );
  XOR U10912 ( .A(n10651), .B(n10650), .Z(n10926) );
  NOR U10913 ( .A(n10925), .B(n10926), .Z(n10652) );
  NOR U10914 ( .A(n10653), .B(n10652), .Z(n11143) );
  NOR U10915 ( .A(n10655), .B(n10654), .Z(n10656) );
  NOR U10916 ( .A(n11143), .B(n10656), .Z(n10657) );
  NOR U10917 ( .A(n10658), .B(n10657), .Z(n10661) );
  NOR U10918 ( .A(n113), .B(n45), .Z(n10660) );
  IV U10919 ( .A(n10660), .Z(n10659) );
  NOR U10920 ( .A(n10661), .B(n10659), .Z(n10666) );
  XOR U10921 ( .A(n10661), .B(n10660), .Z(n11148) );
  XOR U10922 ( .A(n10663), .B(n10662), .Z(n10664) );
  IV U10923 ( .A(n10664), .Z(n11149) );
  NOR U10924 ( .A(n11148), .B(n11149), .Z(n10665) );
  NOR U10925 ( .A(n10666), .B(n10665), .Z(n10673) );
  NOR U10926 ( .A(n83), .B(n45), .Z(n10672) );
  IV U10927 ( .A(n10672), .Z(n10667) );
  NOR U10928 ( .A(n10673), .B(n10667), .Z(n10675) );
  XOR U10929 ( .A(n10669), .B(n10668), .Z(n10670) );
  XOR U10930 ( .A(n10671), .B(n10670), .Z(n10924) );
  XOR U10931 ( .A(n10673), .B(n10672), .Z(n10923) );
  NOR U10932 ( .A(n10924), .B(n10923), .Z(n10674) );
  NOR U10933 ( .A(n10675), .B(n10674), .Z(n10680) );
  XOR U10934 ( .A(n10677), .B(n10676), .Z(n10678) );
  XOR U10935 ( .A(n10679), .B(n10678), .Z(n10681) );
  NOR U10936 ( .A(n10680), .B(n10681), .Z(n10685) );
  IV U10937 ( .A(n10680), .Z(n10682) );
  XOR U10938 ( .A(n10682), .B(n10681), .Z(n11163) );
  NOR U10939 ( .A(n114), .B(n45), .Z(n11164) );
  IV U10940 ( .A(n11164), .Z(n10683) );
  NOR U10941 ( .A(n11163), .B(n10683), .Z(n10684) );
  NOR U10942 ( .A(n10685), .B(n10684), .Z(n11173) );
  IV U10943 ( .A(n11173), .Z(n10686) );
  NOR U10944 ( .A(n10687), .B(n10686), .Z(n10688) );
  NOR U10945 ( .A(n10689), .B(n10688), .Z(n10694) );
  IV U10946 ( .A(n10694), .Z(n10692) );
  XOR U10947 ( .A(n10691), .B(n10690), .Z(n10693) );
  NOR U10948 ( .A(n10692), .B(n10693), .Z(n10697) );
  XOR U10949 ( .A(n10694), .B(n10693), .Z(n11180) );
  NOR U10950 ( .A(n115), .B(n45), .Z(n10695) );
  IV U10951 ( .A(n10695), .Z(n11179) );
  NOR U10952 ( .A(n11180), .B(n11179), .Z(n10696) );
  NOR U10953 ( .A(n10697), .B(n10696), .Z(n10700) );
  NOR U10954 ( .A(n81), .B(n45), .Z(n10699) );
  IV U10955 ( .A(n10699), .Z(n10698) );
  NOR U10956 ( .A(n10700), .B(n10698), .Z(n10704) );
  XOR U10957 ( .A(n10700), .B(n10699), .Z(n11188) );
  XOR U10958 ( .A(n10702), .B(n10701), .Z(n11189) );
  NOR U10959 ( .A(n11188), .B(n11189), .Z(n10703) );
  NOR U10960 ( .A(n10704), .B(n10703), .Z(n10711) );
  NOR U10961 ( .A(n116), .B(n45), .Z(n10710) );
  IV U10962 ( .A(n10710), .Z(n10705) );
  NOR U10963 ( .A(n10711), .B(n10705), .Z(n10713) );
  XOR U10964 ( .A(n10707), .B(n10706), .Z(n10708) );
  XOR U10965 ( .A(n10709), .B(n10708), .Z(n11194) );
  XOR U10966 ( .A(n10711), .B(n10710), .Z(n11193) );
  NOR U10967 ( .A(n11194), .B(n11193), .Z(n10712) );
  NOR U10968 ( .A(n10713), .B(n10712), .Z(n10715) );
  NOR U10969 ( .A(n10714), .B(n10715), .Z(n10719) );
  XOR U10970 ( .A(n10715), .B(n10714), .Z(n10716) );
  IV U10971 ( .A(n10716), .Z(n11203) );
  NOR U10972 ( .A(n80), .B(n45), .Z(n10717) );
  IV U10973 ( .A(n10717), .Z(n11202) );
  NOR U10974 ( .A(n11203), .B(n11202), .Z(n10718) );
  NOR U10975 ( .A(n10719), .B(n10718), .Z(n10721) );
  IV U10976 ( .A(n10721), .Z(n11208) );
  NOR U10977 ( .A(n10720), .B(n11208), .Z(n10726) );
  IV U10978 ( .A(n10720), .Z(n11209) );
  NOR U10979 ( .A(n10721), .B(n11209), .Z(n10724) );
  XOR U10980 ( .A(n10723), .B(n10722), .Z(n11211) );
  NOR U10981 ( .A(n10724), .B(n11211), .Z(n10725) );
  NOR U10982 ( .A(n10726), .B(n10725), .Z(n10727) );
  IV U10983 ( .A(n10727), .Z(n10732) );
  NOR U10984 ( .A(n79), .B(n45), .Z(n10731) );
  IV U10985 ( .A(n10731), .Z(n10728) );
  NOR U10986 ( .A(n10732), .B(n10728), .Z(n10734) );
  XOR U10987 ( .A(n10730), .B(n10729), .Z(n10919) );
  XOR U10988 ( .A(n10732), .B(n10731), .Z(n10920) );
  NOR U10989 ( .A(n10919), .B(n10920), .Z(n10733) );
  NOR U10990 ( .A(n10734), .B(n10733), .Z(n10738) );
  XOR U10991 ( .A(n10736), .B(n10735), .Z(n10737) );
  NOR U10992 ( .A(n10738), .B(n10737), .Z(n10742) );
  XOR U10993 ( .A(n10738), .B(n10737), .Z(n10739) );
  IV U10994 ( .A(n10739), .Z(n10916) );
  NOR U10995 ( .A(n119), .B(n45), .Z(n10917) );
  IV U10996 ( .A(n10917), .Z(n10740) );
  NOR U10997 ( .A(n10916), .B(n10740), .Z(n10741) );
  NOR U10998 ( .A(n10742), .B(n10741), .Z(n10747) );
  NOR U10999 ( .A(n120), .B(n45), .Z(n10746) );
  IV U11000 ( .A(n10746), .Z(n10743) );
  NOR U11001 ( .A(n10747), .B(n10743), .Z(n10750) );
  XOR U11002 ( .A(n10745), .B(n10744), .Z(n10914) );
  IV U11003 ( .A(n10914), .Z(n10748) );
  XOR U11004 ( .A(n10747), .B(n10746), .Z(n10913) );
  NOR U11005 ( .A(n10748), .B(n10913), .Z(n10749) );
  NOR U11006 ( .A(n10750), .B(n10749), .Z(n10753) );
  NOR U11007 ( .A(n123), .B(n45), .Z(n10752) );
  IV U11008 ( .A(n10752), .Z(n10751) );
  NOR U11009 ( .A(n10753), .B(n10751), .Z(n10758) );
  XOR U11010 ( .A(n10753), .B(n10752), .Z(n11233) );
  XOR U11011 ( .A(n10755), .B(n10754), .Z(n11234) );
  IV U11012 ( .A(n11234), .Z(n10756) );
  NOR U11013 ( .A(n11233), .B(n10756), .Z(n10757) );
  NOR U11014 ( .A(n10758), .B(n10757), .Z(n10761) );
  NOR U11015 ( .A(n125), .B(n45), .Z(n10760) );
  IV U11016 ( .A(n10760), .Z(n10759) );
  NOR U11017 ( .A(n10761), .B(n10759), .Z(n10765) );
  XOR U11018 ( .A(n10761), .B(n10760), .Z(n11237) );
  XOR U11019 ( .A(n10763), .B(n10762), .Z(n11238) );
  NOR U11020 ( .A(n11237), .B(n11238), .Z(n10764) );
  NOR U11021 ( .A(n10765), .B(n10764), .Z(n10769) );
  XOR U11022 ( .A(n10767), .B(n10766), .Z(n10768) );
  NOR U11023 ( .A(n10769), .B(n10768), .Z(n10773) );
  XOR U11024 ( .A(n10769), .B(n10768), .Z(n10770) );
  IV U11025 ( .A(n10770), .Z(n11248) );
  NOR U11026 ( .A(n126), .B(n45), .Z(n11249) );
  IV U11027 ( .A(n11249), .Z(n10771) );
  NOR U11028 ( .A(n11248), .B(n10771), .Z(n10772) );
  NOR U11029 ( .A(n10773), .B(n10772), .Z(n11253) );
  IV U11030 ( .A(n11253), .Z(n10774) );
  NOR U11031 ( .A(n10775), .B(n10774), .Z(n10776) );
  NOR U11032 ( .A(n10777), .B(n10776), .Z(n10783) );
  IV U11033 ( .A(n10783), .Z(n10781) );
  IV U11034 ( .A(n10778), .Z(n10780) );
  XOR U11035 ( .A(n10780), .B(n10779), .Z(n10782) );
  NOR U11036 ( .A(n10781), .B(n10782), .Z(n10786) );
  XOR U11037 ( .A(n10783), .B(n10782), .Z(n11262) );
  NOR U11038 ( .A(n131), .B(n45), .Z(n11263) );
  IV U11039 ( .A(n11263), .Z(n10784) );
  NOR U11040 ( .A(n11262), .B(n10784), .Z(n10785) );
  NOR U11041 ( .A(n10786), .B(n10785), .Z(n11270) );
  XOR U11042 ( .A(n10788), .B(n10787), .Z(n11269) );
  NOR U11043 ( .A(n11270), .B(n11269), .Z(n10789) );
  NOR U11044 ( .A(n10790), .B(n10789), .Z(n10793) );
  NOR U11045 ( .A(n135), .B(n45), .Z(n10792) );
  IV U11046 ( .A(n10792), .Z(n10791) );
  NOR U11047 ( .A(n10793), .B(n10791), .Z(n10797) );
  XOR U11048 ( .A(n10793), .B(n10792), .Z(n11274) );
  XOR U11049 ( .A(n10795), .B(n10794), .Z(n11275) );
  NOR U11050 ( .A(n11274), .B(n11275), .Z(n10796) );
  NOR U11051 ( .A(n10797), .B(n10796), .Z(n10802) );
  XOR U11052 ( .A(n10799), .B(n10798), .Z(n10801) );
  IV U11053 ( .A(n10801), .Z(n10800) );
  NOR U11054 ( .A(n10802), .B(n10800), .Z(n10805) );
  XOR U11055 ( .A(n10802), .B(n10801), .Z(n10910) );
  NOR U11056 ( .A(n137), .B(n45), .Z(n10911) );
  IV U11057 ( .A(n10911), .Z(n10803) );
  NOR U11058 ( .A(n10910), .B(n10803), .Z(n10804) );
  NOR U11059 ( .A(n10805), .B(n10804), .Z(n10810) );
  XOR U11060 ( .A(n10807), .B(n10806), .Z(n10809) );
  IV U11061 ( .A(n10809), .Z(n10808) );
  NOR U11062 ( .A(n10810), .B(n10808), .Z(n10813) );
  XOR U11063 ( .A(n10810), .B(n10809), .Z(n11286) );
  NOR U11064 ( .A(n139), .B(n45), .Z(n11287) );
  IV U11065 ( .A(n11287), .Z(n10811) );
  NOR U11066 ( .A(n11286), .B(n10811), .Z(n10812) );
  NOR U11067 ( .A(n10813), .B(n10812), .Z(n10818) );
  XOR U11068 ( .A(n10815), .B(n10814), .Z(n10817) );
  IV U11069 ( .A(n10817), .Z(n10816) );
  NOR U11070 ( .A(n10818), .B(n10816), .Z(n10821) );
  XOR U11071 ( .A(n10818), .B(n10817), .Z(n10907) );
  NOR U11072 ( .A(n141), .B(n45), .Z(n10908) );
  IV U11073 ( .A(n10908), .Z(n10819) );
  NOR U11074 ( .A(n10907), .B(n10819), .Z(n10820) );
  NOR U11075 ( .A(n10821), .B(n10820), .Z(n10826) );
  XOR U11076 ( .A(n10823), .B(n10822), .Z(n10825) );
  IV U11077 ( .A(n10825), .Z(n10824) );
  NOR U11078 ( .A(n10826), .B(n10824), .Z(n10829) );
  XOR U11079 ( .A(n10826), .B(n10825), .Z(n10904) );
  NOR U11080 ( .A(n143), .B(n45), .Z(n10905) );
  IV U11081 ( .A(n10905), .Z(n10827) );
  NOR U11082 ( .A(n10904), .B(n10827), .Z(n10828) );
  NOR U11083 ( .A(n10829), .B(n10828), .Z(n10834) );
  XOR U11084 ( .A(n10831), .B(n10830), .Z(n10833) );
  IV U11085 ( .A(n10833), .Z(n10832) );
  NOR U11086 ( .A(n10834), .B(n10832), .Z(n10837) );
  XOR U11087 ( .A(n10834), .B(n10833), .Z(n10901) );
  NOR U11088 ( .A(n145), .B(n45), .Z(n10902) );
  IV U11089 ( .A(n10902), .Z(n10835) );
  NOR U11090 ( .A(n10901), .B(n10835), .Z(n10836) );
  NOR U11091 ( .A(n10837), .B(n10836), .Z(n11307) );
  XOR U11092 ( .A(n10839), .B(n10838), .Z(n11306) );
  NOR U11093 ( .A(n11307), .B(n11306), .Z(n10840) );
  NOR U11094 ( .A(n10841), .B(n10840), .Z(n10844) );
  NOR U11095 ( .A(n148), .B(n45), .Z(n10843) );
  IV U11096 ( .A(n10843), .Z(n10842) );
  NOR U11097 ( .A(n10844), .B(n10842), .Z(n10848) );
  XOR U11098 ( .A(n10844), .B(n10843), .Z(n11314) );
  XOR U11099 ( .A(n10846), .B(n10845), .Z(n11315) );
  NOR U11100 ( .A(n11314), .B(n11315), .Z(n10847) );
  NOR U11101 ( .A(n10848), .B(n10847), .Z(n10853) );
  XOR U11102 ( .A(n10850), .B(n10849), .Z(n10852) );
  IV U11103 ( .A(n10852), .Z(n10851) );
  NOR U11104 ( .A(n10853), .B(n10851), .Z(n10856) );
  XOR U11105 ( .A(n10853), .B(n10852), .Z(n10898) );
  NOR U11106 ( .A(n150), .B(n45), .Z(n10899) );
  IV U11107 ( .A(n10899), .Z(n10854) );
  NOR U11108 ( .A(n10898), .B(n10854), .Z(n10855) );
  NOR U11109 ( .A(n10856), .B(n10855), .Z(n11330) );
  XOR U11110 ( .A(n10858), .B(n10857), .Z(n11329) );
  NOR U11111 ( .A(n11330), .B(n11329), .Z(n10859) );
  NOR U11112 ( .A(n10860), .B(n10859), .Z(n10864) );
  XOR U11113 ( .A(n10862), .B(n10861), .Z(n10863) );
  NOR U11114 ( .A(n10864), .B(n10863), .Z(n10868) );
  XOR U11115 ( .A(n10864), .B(n10863), .Z(n10865) );
  IV U11116 ( .A(n10865), .Z(n11337) );
  NOR U11117 ( .A(n155), .B(n45), .Z(n11338) );
  IV U11118 ( .A(n11338), .Z(n10866) );
  NOR U11119 ( .A(n11337), .B(n10866), .Z(n10867) );
  NOR U11120 ( .A(n10868), .B(n10867), .Z(n11343) );
  XOR U11121 ( .A(n10870), .B(n10869), .Z(n11342) );
  NOR U11122 ( .A(n11343), .B(n11342), .Z(n10871) );
  NOR U11123 ( .A(n10872), .B(n10871), .Z(n10875) );
  NOR U11124 ( .A(n158), .B(n45), .Z(n10874) );
  IV U11125 ( .A(n10874), .Z(n10873) );
  NOR U11126 ( .A(n10875), .B(n10873), .Z(n10879) );
  XOR U11127 ( .A(n10875), .B(n10874), .Z(n11349) );
  XOR U11128 ( .A(n10877), .B(n10876), .Z(n11350) );
  NOR U11129 ( .A(n11349), .B(n11350), .Z(n10878) );
  NOR U11130 ( .A(n10879), .B(n10878), .Z(n10883) );
  XOR U11131 ( .A(n10881), .B(n10880), .Z(n10882) );
  NOR U11132 ( .A(n10883), .B(n10882), .Z(n10887) );
  XOR U11133 ( .A(n10883), .B(n10882), .Z(n10884) );
  IV U11134 ( .A(n10884), .Z(n11360) );
  NOR U11135 ( .A(n161), .B(n45), .Z(n11361) );
  IV U11136 ( .A(n11361), .Z(n10885) );
  NOR U11137 ( .A(n11360), .B(n10885), .Z(n10886) );
  NOR U11138 ( .A(n10887), .B(n10886), .Z(n10891) );
  IV U11139 ( .A(n10891), .Z(n10888) );
  NOR U11140 ( .A(n10892), .B(n10888), .Z(n10894) );
  XOR U11141 ( .A(n10890), .B(n10889), .Z(n11366) );
  XOR U11142 ( .A(n10892), .B(n10891), .Z(n11365) );
  NOR U11143 ( .A(n11366), .B(n11365), .Z(n10893) );
  NOR U11144 ( .A(n10894), .B(n10893), .Z(n11376) );
  NOR U11145 ( .A(n165), .B(n45), .Z(n10895) );
  IV U11146 ( .A(n10895), .Z(n11377) );
  XOR U11147 ( .A(n11376), .B(n11377), .Z(n11380) );
  XOR U11148 ( .A(n10897), .B(n10896), .Z(n11379) );
  XOR U11149 ( .A(n11380), .B(n11379), .Z(n11373) );
  XOR U11150 ( .A(n10899), .B(n10898), .Z(n11322) );
  NOR U11151 ( .A(n153), .B(n46), .Z(n11323) );
  IV U11152 ( .A(n11323), .Z(n10900) );
  NOR U11153 ( .A(n11322), .B(n10900), .Z(n11325) );
  XOR U11154 ( .A(n10902), .B(n10901), .Z(n11302) );
  NOR U11155 ( .A(n147), .B(n46), .Z(n11303) );
  IV U11156 ( .A(n11303), .Z(n10903) );
  NOR U11157 ( .A(n11302), .B(n10903), .Z(n11305) );
  XOR U11158 ( .A(n10905), .B(n10904), .Z(n11298) );
  NOR U11159 ( .A(n145), .B(n46), .Z(n11299) );
  IV U11160 ( .A(n11299), .Z(n10906) );
  NOR U11161 ( .A(n11298), .B(n10906), .Z(n11301) );
  XOR U11162 ( .A(n10908), .B(n10907), .Z(n11294) );
  NOR U11163 ( .A(n143), .B(n46), .Z(n11295) );
  IV U11164 ( .A(n11295), .Z(n10909) );
  NOR U11165 ( .A(n11294), .B(n10909), .Z(n11297) );
  XOR U11166 ( .A(n10911), .B(n10910), .Z(n11282) );
  NOR U11167 ( .A(n139), .B(n46), .Z(n11283) );
  IV U11168 ( .A(n11283), .Z(n10912) );
  NOR U11169 ( .A(n11282), .B(n10912), .Z(n11285) );
  XOR U11170 ( .A(n10914), .B(n10913), .Z(n11226) );
  NOR U11171 ( .A(n123), .B(n46), .Z(n11227) );
  IV U11172 ( .A(n11227), .Z(n10915) );
  NOR U11173 ( .A(n11226), .B(n10915), .Z(n11229) );
  XOR U11174 ( .A(n10917), .B(n10916), .Z(n11222) );
  NOR U11175 ( .A(n120), .B(n46), .Z(n11223) );
  IV U11176 ( .A(n11223), .Z(n10918) );
  NOR U11177 ( .A(n11222), .B(n10918), .Z(n11225) );
  XOR U11178 ( .A(n10920), .B(n10919), .Z(n10921) );
  IV U11179 ( .A(n10921), .Z(n11217) );
  NOR U11180 ( .A(n119), .B(n46), .Z(n11218) );
  IV U11181 ( .A(n11218), .Z(n10922) );
  NOR U11182 ( .A(n11217), .B(n10922), .Z(n11221) );
  NOR U11183 ( .A(n117), .B(n46), .Z(n11205) );
  NOR U11184 ( .A(n81), .B(n46), .Z(n11177) );
  XOR U11185 ( .A(n10924), .B(n10923), .Z(n11157) );
  NOR U11186 ( .A(n84), .B(n46), .Z(n10927) );
  XOR U11187 ( .A(n10926), .B(n10925), .Z(n10928) );
  NOR U11188 ( .A(n10927), .B(n10928), .Z(n11137) );
  IV U11189 ( .A(n10927), .Z(n11635) );
  IV U11190 ( .A(n10928), .Z(n11634) );
  NOR U11191 ( .A(n11635), .B(n11634), .Z(n11135) );
  NOR U11192 ( .A(n112), .B(n46), .Z(n10929) );
  IV U11193 ( .A(n10929), .Z(n11131) );
  NOR U11194 ( .A(n85), .B(n46), .Z(n11624) );
  XOR U11195 ( .A(n10931), .B(n10930), .Z(n10932) );
  NOR U11196 ( .A(n11624), .B(n10932), .Z(n11124) );
  IV U11197 ( .A(n11624), .Z(n10933) );
  IV U11198 ( .A(n10932), .Z(n11626) );
  NOR U11199 ( .A(n10933), .B(n11626), .Z(n11122) );
  NOR U11200 ( .A(n111), .B(n46), .Z(n11118) );
  NOR U11201 ( .A(n86), .B(n46), .Z(n10936) );
  XOR U11202 ( .A(n10935), .B(n10934), .Z(n10937) );
  IV U11203 ( .A(n10937), .Z(n11612) );
  NOR U11204 ( .A(n10936), .B(n11612), .Z(n11112) );
  IV U11205 ( .A(n10936), .Z(n11610) );
  NOR U11206 ( .A(n10937), .B(n11610), .Z(n11110) );
  XOR U11207 ( .A(n10939), .B(n10938), .Z(n11098) );
  IV U11208 ( .A(n11098), .Z(n11596) );
  NOR U11209 ( .A(n109), .B(n46), .Z(n11097) );
  IV U11210 ( .A(n11097), .Z(n11595) );
  NOR U11211 ( .A(n11596), .B(n11595), .Z(n11101) );
  XOR U11212 ( .A(n10941), .B(n10940), .Z(n10943) );
  NOR U11213 ( .A(n87), .B(n46), .Z(n10944) );
  IV U11214 ( .A(n10944), .Z(n10942) );
  NOR U11215 ( .A(n10943), .B(n10942), .Z(n11087) );
  XOR U11216 ( .A(n10944), .B(n10943), .Z(n11583) );
  NOR U11217 ( .A(n107), .B(n46), .Z(n11081) );
  XOR U11218 ( .A(n10946), .B(n10945), .Z(n11573) );
  IV U11219 ( .A(n11573), .Z(n10948) );
  NOR U11220 ( .A(n88), .B(n46), .Z(n11571) );
  IV U11221 ( .A(n11571), .Z(n10947) );
  NOR U11222 ( .A(n10948), .B(n10947), .Z(n11077) );
  XOR U11223 ( .A(n10950), .B(n10949), .Z(n11064) );
  IV U11224 ( .A(n11064), .Z(n11432) );
  NOR U11225 ( .A(n105), .B(n46), .Z(n11063) );
  IV U11226 ( .A(n11063), .Z(n11431) );
  NOR U11227 ( .A(n11432), .B(n11431), .Z(n11067) );
  XOR U11228 ( .A(n10952), .B(n10951), .Z(n10953) );
  XOR U11229 ( .A(n10954), .B(n10953), .Z(n11060) );
  NOR U11230 ( .A(n104), .B(n46), .Z(n11059) );
  IV U11231 ( .A(n11059), .Z(n10955) );
  NOR U11232 ( .A(n11060), .B(n10955), .Z(n11062) );
  XOR U11233 ( .A(n10957), .B(n10956), .Z(n11055) );
  NOR U11234 ( .A(n89), .B(n46), .Z(n11056) );
  IV U11235 ( .A(n11056), .Z(n10958) );
  NOR U11236 ( .A(n11055), .B(n10958), .Z(n11058) );
  XOR U11237 ( .A(n10960), .B(n10959), .Z(n11052) );
  NOR U11238 ( .A(n103), .B(n46), .Z(n11051) );
  IV U11239 ( .A(n11051), .Z(n10961) );
  NOR U11240 ( .A(n11052), .B(n10961), .Z(n11054) );
  XOR U11241 ( .A(n10963), .B(n10962), .Z(n11048) );
  NOR U11242 ( .A(n90), .B(n46), .Z(n11047) );
  IV U11243 ( .A(n11047), .Z(n10964) );
  NOR U11244 ( .A(n11048), .B(n10964), .Z(n11050) );
  NOR U11245 ( .A(n101), .B(n46), .Z(n10968) );
  IV U11246 ( .A(n10968), .Z(n11451) );
  XOR U11247 ( .A(n10966), .B(n10965), .Z(n10967) );
  IV U11248 ( .A(n10967), .Z(n11453) );
  NOR U11249 ( .A(n11451), .B(n11453), .Z(n11039) );
  NOR U11250 ( .A(n10968), .B(n10967), .Z(n11037) );
  NOR U11251 ( .A(n100), .B(n46), .Z(n11032) );
  XOR U11252 ( .A(n10970), .B(n10969), .Z(n10971) );
  XOR U11253 ( .A(n10972), .B(n10971), .Z(n11033) );
  IV U11254 ( .A(n11033), .Z(n10973) );
  NOR U11255 ( .A(n11032), .B(n10973), .Z(n11035) );
  NOR U11256 ( .A(n99), .B(n46), .Z(n11028) );
  XOR U11257 ( .A(n10975), .B(n10974), .Z(n11027) );
  NOR U11258 ( .A(n11028), .B(n11027), .Z(n11031) );
  IV U11259 ( .A(n10976), .Z(n10978) );
  XOR U11260 ( .A(n10978), .B(n10977), .Z(n11022) );
  NOR U11261 ( .A(n98), .B(n46), .Z(n11023) );
  IV U11262 ( .A(n11023), .Z(n10979) );
  NOR U11263 ( .A(n11022), .B(n10979), .Z(n11025) );
  XOR U11264 ( .A(n10981), .B(n10980), .Z(n11018) );
  NOR U11265 ( .A(n91), .B(n46), .Z(n11019) );
  IV U11266 ( .A(n11019), .Z(n10982) );
  NOR U11267 ( .A(n11018), .B(n10982), .Z(n11021) );
  IV U11268 ( .A(n10983), .Z(n10985) );
  XOR U11269 ( .A(n10985), .B(n10984), .Z(n11014) );
  NOR U11270 ( .A(n97), .B(n46), .Z(n11015) );
  IV U11271 ( .A(n11015), .Z(n10986) );
  NOR U11272 ( .A(n11014), .B(n10986), .Z(n11017) );
  IV U11273 ( .A(n10987), .Z(n10989) );
  XOR U11274 ( .A(n10989), .B(n10988), .Z(n11010) );
  NOR U11275 ( .A(n96), .B(n46), .Z(n11011) );
  IV U11276 ( .A(n11011), .Z(n10990) );
  NOR U11277 ( .A(n11010), .B(n10990), .Z(n11013) );
  NOR U11278 ( .A(n95), .B(n46), .Z(n11007) );
  IV U11279 ( .A(n11007), .Z(n10993) );
  XOR U11280 ( .A(n10992), .B(n10991), .Z(n11006) );
  NOR U11281 ( .A(n10993), .B(n11006), .Z(n11009) );
  NOR U11282 ( .A(n93), .B(n46), .Z(n12053) );
  IV U11283 ( .A(n12053), .Z(n10994) );
  NOR U11284 ( .A(n45), .B(n168), .Z(n11002) );
  IV U11285 ( .A(n11002), .Z(n10997) );
  NOR U11286 ( .A(n10994), .B(n10997), .Z(n10995) );
  IV U11287 ( .A(n10995), .Z(n10996) );
  NOR U11288 ( .A(n94), .B(n10996), .Z(n11005) );
  NOR U11289 ( .A(n10997), .B(n93), .Z(n10998) );
  XOR U11290 ( .A(n94), .B(n10998), .Z(n10999) );
  NOR U11291 ( .A(n46), .B(n10999), .Z(n11000) );
  IV U11292 ( .A(n11000), .Z(n11482) );
  XOR U11293 ( .A(n11002), .B(n11001), .Z(n11481) );
  IV U11294 ( .A(n11481), .Z(n11003) );
  NOR U11295 ( .A(n11482), .B(n11003), .Z(n11004) );
  NOR U11296 ( .A(n11005), .B(n11004), .Z(n11477) );
  XOR U11297 ( .A(n11007), .B(n11006), .Z(n11478) );
  NOR U11298 ( .A(n11477), .B(n11478), .Z(n11008) );
  NOR U11299 ( .A(n11009), .B(n11008), .Z(n11473) );
  XOR U11300 ( .A(n11011), .B(n11010), .Z(n11474) );
  NOR U11301 ( .A(n11473), .B(n11474), .Z(n11012) );
  NOR U11302 ( .A(n11013), .B(n11012), .Z(n11469) );
  XOR U11303 ( .A(n11015), .B(n11014), .Z(n11470) );
  NOR U11304 ( .A(n11469), .B(n11470), .Z(n11016) );
  NOR U11305 ( .A(n11017), .B(n11016), .Z(n11465) );
  XOR U11306 ( .A(n11019), .B(n11018), .Z(n11466) );
  NOR U11307 ( .A(n11465), .B(n11466), .Z(n11020) );
  NOR U11308 ( .A(n11021), .B(n11020), .Z(n11461) );
  XOR U11309 ( .A(n11023), .B(n11022), .Z(n11462) );
  NOR U11310 ( .A(n11461), .B(n11462), .Z(n11024) );
  NOR U11311 ( .A(n11025), .B(n11024), .Z(n11026) );
  IV U11312 ( .A(n11026), .Z(n11459) );
  XOR U11313 ( .A(n11028), .B(n11027), .Z(n11029) );
  IV U11314 ( .A(n11029), .Z(n11458) );
  NOR U11315 ( .A(n11459), .B(n11458), .Z(n11030) );
  NOR U11316 ( .A(n11031), .B(n11030), .Z(n11456) );
  XOR U11317 ( .A(n11033), .B(n11032), .Z(n11455) );
  NOR U11318 ( .A(n11456), .B(n11455), .Z(n11034) );
  NOR U11319 ( .A(n11035), .B(n11034), .Z(n11036) );
  IV U11320 ( .A(n11036), .Z(n11450) );
  NOR U11321 ( .A(n11037), .B(n11450), .Z(n11038) );
  NOR U11322 ( .A(n11039), .B(n11038), .Z(n11044) );
  NOR U11323 ( .A(n102), .B(n46), .Z(n11043) );
  IV U11324 ( .A(n11043), .Z(n11040) );
  NOR U11325 ( .A(n11044), .B(n11040), .Z(n11046) );
  XOR U11326 ( .A(n11042), .B(n11041), .Z(n11447) );
  XOR U11327 ( .A(n11044), .B(n11043), .Z(n11446) );
  NOR U11328 ( .A(n11447), .B(n11446), .Z(n11045) );
  NOR U11329 ( .A(n11046), .B(n11045), .Z(n11538) );
  XOR U11330 ( .A(n11048), .B(n11047), .Z(n11539) );
  NOR U11331 ( .A(n11538), .B(n11539), .Z(n11049) );
  NOR U11332 ( .A(n11050), .B(n11049), .Z(n11442) );
  XOR U11333 ( .A(n11052), .B(n11051), .Z(n11443) );
  NOR U11334 ( .A(n11442), .B(n11443), .Z(n11053) );
  NOR U11335 ( .A(n11054), .B(n11053), .Z(n11438) );
  XOR U11336 ( .A(n11056), .B(n11055), .Z(n11439) );
  NOR U11337 ( .A(n11438), .B(n11439), .Z(n11057) );
  NOR U11338 ( .A(n11058), .B(n11057), .Z(n11437) );
  XOR U11339 ( .A(n11060), .B(n11059), .Z(n11436) );
  NOR U11340 ( .A(n11437), .B(n11436), .Z(n11061) );
  NOR U11341 ( .A(n11062), .B(n11061), .Z(n11434) );
  NOR U11342 ( .A(n11064), .B(n11063), .Z(n11065) );
  NOR U11343 ( .A(n11434), .B(n11065), .Z(n11066) );
  NOR U11344 ( .A(n11067), .B(n11066), .Z(n11072) );
  NOR U11345 ( .A(n106), .B(n46), .Z(n11071) );
  IV U11346 ( .A(n11071), .Z(n11068) );
  NOR U11347 ( .A(n11072), .B(n11068), .Z(n11074) );
  XOR U11348 ( .A(n11070), .B(n11069), .Z(n11430) );
  XOR U11349 ( .A(n11072), .B(n11071), .Z(n11429) );
  NOR U11350 ( .A(n11430), .B(n11429), .Z(n11073) );
  NOR U11351 ( .A(n11074), .B(n11073), .Z(n11570) );
  NOR U11352 ( .A(n11571), .B(n11573), .Z(n11075) );
  NOR U11353 ( .A(n11570), .B(n11075), .Z(n11076) );
  NOR U11354 ( .A(n11077), .B(n11076), .Z(n11082) );
  IV U11355 ( .A(n11082), .Z(n11078) );
  NOR U11356 ( .A(n11081), .B(n11078), .Z(n11084) );
  XOR U11357 ( .A(n11080), .B(n11079), .Z(n11426) );
  XOR U11358 ( .A(n11082), .B(n11081), .Z(n11425) );
  NOR U11359 ( .A(n11426), .B(n11425), .Z(n11083) );
  NOR U11360 ( .A(n11084), .B(n11083), .Z(n11584) );
  IV U11361 ( .A(n11584), .Z(n11085) );
  NOR U11362 ( .A(n11583), .B(n11085), .Z(n11086) );
  NOR U11363 ( .A(n11087), .B(n11086), .Z(n11094) );
  NOR U11364 ( .A(n108), .B(n46), .Z(n11093) );
  IV U11365 ( .A(n11093), .Z(n11088) );
  NOR U11366 ( .A(n11094), .B(n11088), .Z(n11096) );
  XOR U11367 ( .A(n11090), .B(n11089), .Z(n11091) );
  XOR U11368 ( .A(n11092), .B(n11091), .Z(n11421) );
  XOR U11369 ( .A(n11094), .B(n11093), .Z(n11420) );
  NOR U11370 ( .A(n11421), .B(n11420), .Z(n11095) );
  NOR U11371 ( .A(n11096), .B(n11095), .Z(n11598) );
  NOR U11372 ( .A(n11098), .B(n11097), .Z(n11099) );
  NOR U11373 ( .A(n11598), .B(n11099), .Z(n11100) );
  NOR U11374 ( .A(n11101), .B(n11100), .Z(n11105) );
  NOR U11375 ( .A(n110), .B(n46), .Z(n11106) );
  IV U11376 ( .A(n11106), .Z(n11102) );
  NOR U11377 ( .A(n11105), .B(n11102), .Z(n11108) );
  XOR U11378 ( .A(n11104), .B(n11103), .Z(n11418) );
  XOR U11379 ( .A(n11106), .B(n11105), .Z(n11419) );
  NOR U11380 ( .A(n11418), .B(n11419), .Z(n11107) );
  NOR U11381 ( .A(n11108), .B(n11107), .Z(n11109) );
  IV U11382 ( .A(n11109), .Z(n11609) );
  NOR U11383 ( .A(n11110), .B(n11609), .Z(n11111) );
  NOR U11384 ( .A(n11112), .B(n11111), .Z(n11117) );
  NOR U11385 ( .A(n11118), .B(n11117), .Z(n11121) );
  XOR U11386 ( .A(n11114), .B(n11113), .Z(n11115) );
  XOR U11387 ( .A(n11116), .B(n11115), .Z(n11414) );
  XOR U11388 ( .A(n11118), .B(n11117), .Z(n11415) );
  IV U11389 ( .A(n11415), .Z(n11119) );
  NOR U11390 ( .A(n11414), .B(n11119), .Z(n11120) );
  NOR U11391 ( .A(n11121), .B(n11120), .Z(n11623) );
  NOR U11392 ( .A(n11122), .B(n11623), .Z(n11123) );
  NOR U11393 ( .A(n11124), .B(n11123), .Z(n11130) );
  IV U11394 ( .A(n11130), .Z(n11125) );
  NOR U11395 ( .A(n11131), .B(n11125), .Z(n11133) );
  XOR U11396 ( .A(n11127), .B(n11126), .Z(n11128) );
  XOR U11397 ( .A(n11129), .B(n11128), .Z(n11410) );
  XOR U11398 ( .A(n11131), .B(n11130), .Z(n11411) );
  NOR U11399 ( .A(n11410), .B(n11411), .Z(n11132) );
  NOR U11400 ( .A(n11133), .B(n11132), .Z(n11637) );
  IV U11401 ( .A(n11637), .Z(n11134) );
  NOR U11402 ( .A(n11135), .B(n11134), .Z(n11136) );
  NOR U11403 ( .A(n11137), .B(n11136), .Z(n11138) );
  IV U11404 ( .A(n11138), .Z(n11145) );
  NOR U11405 ( .A(n113), .B(n46), .Z(n11144) );
  IV U11406 ( .A(n11144), .Z(n11139) );
  NOR U11407 ( .A(n11145), .B(n11139), .Z(n11147) );
  XOR U11408 ( .A(n11141), .B(n11140), .Z(n11142) );
  XOR U11409 ( .A(n11143), .B(n11142), .Z(n11404) );
  XOR U11410 ( .A(n11145), .B(n11144), .Z(n11405) );
  NOR U11411 ( .A(n11404), .B(n11405), .Z(n11146) );
  NOR U11412 ( .A(n11147), .B(n11146), .Z(n11151) );
  XOR U11413 ( .A(n11149), .B(n11148), .Z(n11152) );
  IV U11414 ( .A(n11152), .Z(n11150) );
  NOR U11415 ( .A(n11151), .B(n11150), .Z(n11155) );
  NOR U11416 ( .A(n83), .B(n46), .Z(n11648) );
  IV U11417 ( .A(n11648), .Z(n11153) );
  XOR U11418 ( .A(n11152), .B(n11151), .Z(n11647) );
  NOR U11419 ( .A(n11153), .B(n11647), .Z(n11154) );
  NOR U11420 ( .A(n11155), .B(n11154), .Z(n11656) );
  IV U11421 ( .A(n11656), .Z(n11156) );
  NOR U11422 ( .A(n11157), .B(n11156), .Z(n11160) );
  IV U11423 ( .A(n11157), .Z(n11658) );
  NOR U11424 ( .A(n11656), .B(n11658), .Z(n11158) );
  NOR U11425 ( .A(n114), .B(n46), .Z(n11655) );
  NOR U11426 ( .A(n11158), .B(n11655), .Z(n11159) );
  NOR U11427 ( .A(n11160), .B(n11159), .Z(n11162) );
  IV U11428 ( .A(n11162), .Z(n11665) );
  NOR U11429 ( .A(n82), .B(n46), .Z(n11161) );
  IV U11430 ( .A(n11161), .Z(n11664) );
  NOR U11431 ( .A(n11665), .B(n11664), .Z(n11167) );
  NOR U11432 ( .A(n11162), .B(n11161), .Z(n11165) );
  XOR U11433 ( .A(n11164), .B(n11163), .Z(n11667) );
  NOR U11434 ( .A(n11165), .B(n11667), .Z(n11166) );
  NOR U11435 ( .A(n11167), .B(n11166), .Z(n11168) );
  NOR U11436 ( .A(n115), .B(n46), .Z(n11169) );
  IV U11437 ( .A(n11169), .Z(n11400) );
  NOR U11438 ( .A(n11168), .B(n11400), .Z(n11176) );
  IV U11439 ( .A(n11168), .Z(n11401) );
  NOR U11440 ( .A(n11169), .B(n11401), .Z(n11174) );
  XOR U11441 ( .A(n11171), .B(n11170), .Z(n11172) );
  XOR U11442 ( .A(n11173), .B(n11172), .Z(n11403) );
  NOR U11443 ( .A(n11174), .B(n11403), .Z(n11175) );
  NOR U11444 ( .A(n11176), .B(n11175), .Z(n11178) );
  IV U11445 ( .A(n11178), .Z(n11680) );
  NOR U11446 ( .A(n11177), .B(n11680), .Z(n11183) );
  IV U11447 ( .A(n11177), .Z(n11681) );
  NOR U11448 ( .A(n11178), .B(n11681), .Z(n11181) );
  XOR U11449 ( .A(n11180), .B(n11179), .Z(n11683) );
  NOR U11450 ( .A(n11181), .B(n11683), .Z(n11182) );
  NOR U11451 ( .A(n11183), .B(n11182), .Z(n11187) );
  IV U11452 ( .A(n11187), .Z(n11185) );
  NOR U11453 ( .A(n116), .B(n46), .Z(n11184) );
  IV U11454 ( .A(n11184), .Z(n11186) );
  NOR U11455 ( .A(n11185), .B(n11186), .Z(n11192) );
  XOR U11456 ( .A(n11187), .B(n11186), .Z(n11688) );
  XOR U11457 ( .A(n11189), .B(n11188), .Z(n11687) );
  IV U11458 ( .A(n11687), .Z(n11190) );
  NOR U11459 ( .A(n11688), .B(n11190), .Z(n11191) );
  NOR U11460 ( .A(n11192), .B(n11191), .Z(n11197) );
  XOR U11461 ( .A(n11194), .B(n11193), .Z(n11196) );
  IV U11462 ( .A(n11196), .Z(n11195) );
  NOR U11463 ( .A(n11197), .B(n11195), .Z(n11200) );
  XOR U11464 ( .A(n11197), .B(n11196), .Z(n11397) );
  NOR U11465 ( .A(n80), .B(n46), .Z(n11396) );
  IV U11466 ( .A(n11396), .Z(n11198) );
  NOR U11467 ( .A(n11397), .B(n11198), .Z(n11199) );
  NOR U11468 ( .A(n11200), .B(n11199), .Z(n11204) );
  IV U11469 ( .A(n11204), .Z(n11201) );
  NOR U11470 ( .A(n11205), .B(n11201), .Z(n11207) );
  XOR U11471 ( .A(n11203), .B(n11202), .Z(n11702) );
  XOR U11472 ( .A(n11205), .B(n11204), .Z(n11701) );
  NOR U11473 ( .A(n11702), .B(n11701), .Z(n11206) );
  NOR U11474 ( .A(n11207), .B(n11206), .Z(n11213) );
  XOR U11475 ( .A(n11209), .B(n11208), .Z(n11210) );
  XOR U11476 ( .A(n11211), .B(n11210), .Z(n11214) );
  IV U11477 ( .A(n11214), .Z(n11212) );
  NOR U11478 ( .A(n11213), .B(n11212), .Z(n11216) );
  NOR U11479 ( .A(n79), .B(n46), .Z(n11709) );
  XOR U11480 ( .A(n11214), .B(n11213), .Z(n11708) );
  NOR U11481 ( .A(n11709), .B(n11708), .Z(n11215) );
  NOR U11482 ( .A(n11216), .B(n11215), .Z(n11715) );
  IV U11483 ( .A(n11715), .Z(n11219) );
  XOR U11484 ( .A(n11218), .B(n11217), .Z(n11714) );
  NOR U11485 ( .A(n11219), .B(n11714), .Z(n11220) );
  NOR U11486 ( .A(n11221), .B(n11220), .Z(n11726) );
  XOR U11487 ( .A(n11223), .B(n11222), .Z(n11725) );
  NOR U11488 ( .A(n11726), .B(n11725), .Z(n11224) );
  NOR U11489 ( .A(n11225), .B(n11224), .Z(n11734) );
  XOR U11490 ( .A(n11227), .B(n11226), .Z(n11733) );
  NOR U11491 ( .A(n11734), .B(n11733), .Z(n11228) );
  NOR U11492 ( .A(n11229), .B(n11228), .Z(n11232) );
  NOR U11493 ( .A(n125), .B(n46), .Z(n11231) );
  IV U11494 ( .A(n11231), .Z(n11230) );
  NOR U11495 ( .A(n11232), .B(n11230), .Z(n11236) );
  XOR U11496 ( .A(n11232), .B(n11231), .Z(n11393) );
  XOR U11497 ( .A(n11234), .B(n11233), .Z(n11392) );
  NOR U11498 ( .A(n11393), .B(n11392), .Z(n11235) );
  NOR U11499 ( .A(n11236), .B(n11235), .Z(n11241) );
  XOR U11500 ( .A(n11238), .B(n11237), .Z(n11240) );
  IV U11501 ( .A(n11240), .Z(n11239) );
  NOR U11502 ( .A(n11241), .B(n11239), .Z(n11244) );
  XOR U11503 ( .A(n11241), .B(n11240), .Z(n11745) );
  NOR U11504 ( .A(n126), .B(n46), .Z(n11746) );
  IV U11505 ( .A(n11746), .Z(n11242) );
  NOR U11506 ( .A(n11745), .B(n11242), .Z(n11243) );
  NOR U11507 ( .A(n11244), .B(n11243), .Z(n11247) );
  NOR U11508 ( .A(n128), .B(n46), .Z(n11246) );
  IV U11509 ( .A(n11246), .Z(n11245) );
  NOR U11510 ( .A(n11247), .B(n11245), .Z(n11251) );
  XOR U11511 ( .A(n11247), .B(n11246), .Z(n11752) );
  XOR U11512 ( .A(n11249), .B(n11248), .Z(n11753) );
  NOR U11513 ( .A(n11752), .B(n11753), .Z(n11250) );
  NOR U11514 ( .A(n11251), .B(n11250), .Z(n11256) );
  NOR U11515 ( .A(n131), .B(n46), .Z(n11255) );
  IV U11516 ( .A(n11255), .Z(n11252) );
  NOR U11517 ( .A(n11256), .B(n11252), .Z(n11258) );
  XOR U11518 ( .A(n11254), .B(n11253), .Z(n11758) );
  XOR U11519 ( .A(n11256), .B(n11255), .Z(n11757) );
  NOR U11520 ( .A(n11758), .B(n11757), .Z(n11257) );
  NOR U11521 ( .A(n11258), .B(n11257), .Z(n11261) );
  NOR U11522 ( .A(n133), .B(n46), .Z(n11260) );
  IV U11523 ( .A(n11260), .Z(n11259) );
  NOR U11524 ( .A(n11261), .B(n11259), .Z(n11265) );
  XOR U11525 ( .A(n11261), .B(n11260), .Z(n11768) );
  XOR U11526 ( .A(n11263), .B(n11262), .Z(n11769) );
  NOR U11527 ( .A(n11768), .B(n11769), .Z(n11264) );
  NOR U11528 ( .A(n11265), .B(n11264), .Z(n11268) );
  NOR U11529 ( .A(n135), .B(n46), .Z(n11267) );
  IV U11530 ( .A(n11267), .Z(n11266) );
  NOR U11531 ( .A(n11268), .B(n11266), .Z(n11273) );
  XOR U11532 ( .A(n11268), .B(n11267), .Z(n11773) );
  XOR U11533 ( .A(n11270), .B(n11269), .Z(n11774) );
  IV U11534 ( .A(n11774), .Z(n11271) );
  NOR U11535 ( .A(n11773), .B(n11271), .Z(n11272) );
  NOR U11536 ( .A(n11273), .B(n11272), .Z(n11278) );
  XOR U11537 ( .A(n11275), .B(n11274), .Z(n11277) );
  IV U11538 ( .A(n11277), .Z(n11276) );
  NOR U11539 ( .A(n11278), .B(n11276), .Z(n11281) );
  XOR U11540 ( .A(n11278), .B(n11277), .Z(n11781) );
  NOR U11541 ( .A(n137), .B(n46), .Z(n11782) );
  IV U11542 ( .A(n11782), .Z(n11279) );
  NOR U11543 ( .A(n11781), .B(n11279), .Z(n11280) );
  NOR U11544 ( .A(n11281), .B(n11280), .Z(n11793) );
  XOR U11545 ( .A(n11283), .B(n11282), .Z(n11792) );
  NOR U11546 ( .A(n11793), .B(n11792), .Z(n11284) );
  NOR U11547 ( .A(n11285), .B(n11284), .Z(n11288) );
  XOR U11548 ( .A(n11287), .B(n11286), .Z(n11289) );
  NOR U11549 ( .A(n11288), .B(n11289), .Z(n11293) );
  IV U11550 ( .A(n11288), .Z(n11290) );
  XOR U11551 ( .A(n11290), .B(n11289), .Z(n11800) );
  NOR U11552 ( .A(n141), .B(n46), .Z(n11801) );
  IV U11553 ( .A(n11801), .Z(n11291) );
  NOR U11554 ( .A(n11800), .B(n11291), .Z(n11292) );
  NOR U11555 ( .A(n11293), .B(n11292), .Z(n11805) );
  XOR U11556 ( .A(n11295), .B(n11294), .Z(n11804) );
  NOR U11557 ( .A(n11805), .B(n11804), .Z(n11296) );
  NOR U11558 ( .A(n11297), .B(n11296), .Z(n11813) );
  XOR U11559 ( .A(n11299), .B(n11298), .Z(n11812) );
  NOR U11560 ( .A(n11813), .B(n11812), .Z(n11300) );
  NOR U11561 ( .A(n11301), .B(n11300), .Z(n11821) );
  XOR U11562 ( .A(n11303), .B(n11302), .Z(n11820) );
  NOR U11563 ( .A(n11821), .B(n11820), .Z(n11304) );
  NOR U11564 ( .A(n11305), .B(n11304), .Z(n11310) );
  XOR U11565 ( .A(n11307), .B(n11306), .Z(n11309) );
  IV U11566 ( .A(n11309), .Z(n11308) );
  NOR U11567 ( .A(n11310), .B(n11308), .Z(n11313) );
  XOR U11568 ( .A(n11310), .B(n11309), .Z(n11389) );
  NOR U11569 ( .A(n148), .B(n46), .Z(n11390) );
  IV U11570 ( .A(n11390), .Z(n11311) );
  NOR U11571 ( .A(n11389), .B(n11311), .Z(n11312) );
  NOR U11572 ( .A(n11313), .B(n11312), .Z(n11318) );
  XOR U11573 ( .A(n11315), .B(n11314), .Z(n11317) );
  IV U11574 ( .A(n11317), .Z(n11316) );
  NOR U11575 ( .A(n11318), .B(n11316), .Z(n11321) );
  XOR U11576 ( .A(n11318), .B(n11317), .Z(n11835) );
  NOR U11577 ( .A(n150), .B(n46), .Z(n11836) );
  IV U11578 ( .A(n11836), .Z(n11319) );
  NOR U11579 ( .A(n11835), .B(n11319), .Z(n11320) );
  NOR U11580 ( .A(n11321), .B(n11320), .Z(n11843) );
  XOR U11581 ( .A(n11323), .B(n11322), .Z(n11842) );
  NOR U11582 ( .A(n11843), .B(n11842), .Z(n11324) );
  NOR U11583 ( .A(n11325), .B(n11324), .Z(n11328) );
  NOR U11584 ( .A(n155), .B(n46), .Z(n11327) );
  IV U11585 ( .A(n11327), .Z(n11326) );
  NOR U11586 ( .A(n11328), .B(n11326), .Z(n11333) );
  XOR U11587 ( .A(n11328), .B(n11327), .Z(n11847) );
  XOR U11588 ( .A(n11330), .B(n11329), .Z(n11848) );
  IV U11589 ( .A(n11848), .Z(n11331) );
  NOR U11590 ( .A(n11847), .B(n11331), .Z(n11332) );
  NOR U11591 ( .A(n11333), .B(n11332), .Z(n11336) );
  NOR U11592 ( .A(n156), .B(n46), .Z(n11335) );
  IV U11593 ( .A(n11335), .Z(n11334) );
  NOR U11594 ( .A(n11336), .B(n11334), .Z(n11340) );
  XOR U11595 ( .A(n11336), .B(n11335), .Z(n11858) );
  XOR U11596 ( .A(n11338), .B(n11337), .Z(n11859) );
  NOR U11597 ( .A(n11858), .B(n11859), .Z(n11339) );
  NOR U11598 ( .A(n11340), .B(n11339), .Z(n11345) );
  NOR U11599 ( .A(n158), .B(n46), .Z(n11344) );
  IV U11600 ( .A(n11344), .Z(n11341) );
  NOR U11601 ( .A(n11345), .B(n11341), .Z(n11348) );
  XOR U11602 ( .A(n11343), .B(n11342), .Z(n11864) );
  IV U11603 ( .A(n11864), .Z(n11346) );
  XOR U11604 ( .A(n11345), .B(n11344), .Z(n11863) );
  NOR U11605 ( .A(n11346), .B(n11863), .Z(n11347) );
  NOR U11606 ( .A(n11348), .B(n11347), .Z(n11353) );
  XOR U11607 ( .A(n11350), .B(n11349), .Z(n11352) );
  IV U11608 ( .A(n11352), .Z(n11351) );
  NOR U11609 ( .A(n11353), .B(n11351), .Z(n11356) );
  XOR U11610 ( .A(n11353), .B(n11352), .Z(n11386) );
  NOR U11611 ( .A(n161), .B(n46), .Z(n11387) );
  IV U11612 ( .A(n11387), .Z(n11354) );
  NOR U11613 ( .A(n11386), .B(n11354), .Z(n11355) );
  NOR U11614 ( .A(n11356), .B(n11355), .Z(n11359) );
  NOR U11615 ( .A(n163), .B(n46), .Z(n11358) );
  IV U11616 ( .A(n11358), .Z(n11357) );
  NOR U11617 ( .A(n11359), .B(n11357), .Z(n11363) );
  XOR U11618 ( .A(n11359), .B(n11358), .Z(n11876) );
  XOR U11619 ( .A(n11361), .B(n11360), .Z(n11877) );
  NOR U11620 ( .A(n11876), .B(n11877), .Z(n11362) );
  NOR U11621 ( .A(n11363), .B(n11362), .Z(n11368) );
  NOR U11622 ( .A(n165), .B(n46), .Z(n11367) );
  IV U11623 ( .A(n11367), .Z(n11364) );
  NOR U11624 ( .A(n11368), .B(n11364), .Z(n11370) );
  XOR U11625 ( .A(n11366), .B(n11365), .Z(n11884) );
  XOR U11626 ( .A(n11368), .B(n11367), .Z(n11883) );
  NOR U11627 ( .A(n11884), .B(n11883), .Z(n11369) );
  NOR U11628 ( .A(n11370), .B(n11369), .Z(n11372) );
  IV U11629 ( .A(n11372), .Z(n11371) );
  NOR U11630 ( .A(n11373), .B(n11371), .Z(n11375) );
  NOR U11631 ( .A(n167), .B(n46), .Z(n11892) );
  XOR U11632 ( .A(n11373), .B(n11372), .Z(n11891) );
  NOR U11633 ( .A(n11892), .B(n11891), .Z(n11374) );
  NOR U11634 ( .A(n11375), .B(n11374), .Z(n11894) );
  IV U11635 ( .A(n11894), .Z(n11385) );
  NOR U11636 ( .A(n167), .B(n45), .Z(n11899) );
  IV U11637 ( .A(n11376), .Z(n11378) );
  NOR U11638 ( .A(n11378), .B(n11377), .Z(n11382) );
  NOR U11639 ( .A(n11380), .B(n11379), .Z(n11381) );
  NOR U11640 ( .A(n11382), .B(n11381), .Z(n11898) );
  XOR U11641 ( .A(n11384), .B(n11383), .Z(n11896) );
  XOR U11642 ( .A(n11898), .B(n11896), .Z(n11901) );
  XOR U11643 ( .A(n11899), .B(n11901), .Z(n11893) );
  NOR U11644 ( .A(n11385), .B(n11893), .Z(n31664) );
  XOR U11645 ( .A(n11387), .B(n11386), .Z(n11871) );
  NOR U11646 ( .A(n163), .B(n47), .Z(n11872) );
  IV U11647 ( .A(n11872), .Z(n11388) );
  NOR U11648 ( .A(n11871), .B(n11388), .Z(n11874) );
  XOR U11649 ( .A(n11390), .B(n11389), .Z(n11828) );
  NOR U11650 ( .A(n150), .B(n47), .Z(n11829) );
  IV U11651 ( .A(n11829), .Z(n11391) );
  NOR U11652 ( .A(n11828), .B(n11391), .Z(n11831) );
  IV U11653 ( .A(n11392), .Z(n11394) );
  XOR U11654 ( .A(n11394), .B(n11393), .Z(n11738) );
  NOR U11655 ( .A(n126), .B(n47), .Z(n11739) );
  IV U11656 ( .A(n11739), .Z(n11395) );
  NOR U11657 ( .A(n11738), .B(n11395), .Z(n11741) );
  NOR U11658 ( .A(n117), .B(n47), .Z(n11399) );
  XOR U11659 ( .A(n11397), .B(n11396), .Z(n12255) );
  IV U11660 ( .A(n12255), .Z(n11398) );
  NOR U11661 ( .A(n11399), .B(n11398), .Z(n11698) );
  IV U11662 ( .A(n11399), .Z(n12256) );
  NOR U11663 ( .A(n12256), .B(n12255), .Z(n11696) );
  XOR U11664 ( .A(n11401), .B(n11400), .Z(n11402) );
  XOR U11665 ( .A(n11403), .B(n11402), .Z(n12235) );
  IV U11666 ( .A(n12235), .Z(n11672) );
  NOR U11667 ( .A(n82), .B(n47), .Z(n11653) );
  XOR U11668 ( .A(n11405), .B(n11404), .Z(n11407) );
  NOR U11669 ( .A(n83), .B(n47), .Z(n11406) );
  NOR U11670 ( .A(n11407), .B(n11406), .Z(n11644) );
  IV U11671 ( .A(n11406), .Z(n11408) );
  XOR U11672 ( .A(n11408), .B(n11407), .Z(n12208) );
  NOR U11673 ( .A(n113), .B(n47), .Z(n11409) );
  IV U11674 ( .A(n11409), .Z(n11639) );
  XOR U11675 ( .A(n11411), .B(n11410), .Z(n11412) );
  NOR U11676 ( .A(n84), .B(n47), .Z(n11413) );
  NOR U11677 ( .A(n11412), .B(n11413), .Z(n11632) );
  IV U11678 ( .A(n11412), .Z(n11961) );
  IV U11679 ( .A(n11413), .Z(n11960) );
  NOR U11680 ( .A(n11961), .B(n11960), .Z(n11630) );
  XOR U11681 ( .A(n11415), .B(n11414), .Z(n12190) );
  IV U11682 ( .A(n12190), .Z(n11417) );
  NOR U11683 ( .A(n85), .B(n47), .Z(n12188) );
  IV U11684 ( .A(n12188), .Z(n11416) );
  NOR U11685 ( .A(n11417), .B(n11416), .Z(n11619) );
  NOR U11686 ( .A(n12188), .B(n12190), .Z(n11617) );
  XOR U11687 ( .A(n11419), .B(n11418), .Z(n11604) );
  IV U11688 ( .A(n11604), .Z(n12174) );
  NOR U11689 ( .A(n86), .B(n47), .Z(n11603) );
  IV U11690 ( .A(n11603), .Z(n12173) );
  NOR U11691 ( .A(n12174), .B(n12173), .Z(n11607) );
  XOR U11692 ( .A(n11421), .B(n11420), .Z(n11422) );
  NOR U11693 ( .A(n109), .B(n47), .Z(n11423) );
  NOR U11694 ( .A(n11422), .B(n11423), .Z(n11592) );
  IV U11695 ( .A(n11422), .Z(n11980) );
  IV U11696 ( .A(n11423), .Z(n11979) );
  NOR U11697 ( .A(n11980), .B(n11979), .Z(n11590) );
  NOR U11698 ( .A(n108), .B(n47), .Z(n11424) );
  IV U11699 ( .A(n11424), .Z(n11586) );
  NOR U11700 ( .A(n87), .B(n47), .Z(n11427) );
  XOR U11701 ( .A(n11426), .B(n11425), .Z(n11428) );
  IV U11702 ( .A(n11428), .Z(n12154) );
  NOR U11703 ( .A(n11427), .B(n12154), .Z(n11581) );
  IV U11704 ( .A(n11427), .Z(n12152) );
  NOR U11705 ( .A(n11428), .B(n12152), .Z(n11579) );
  XOR U11706 ( .A(n11430), .B(n11429), .Z(n11565) );
  IV U11707 ( .A(n11565), .Z(n11993) );
  NOR U11708 ( .A(n88), .B(n47), .Z(n11564) );
  IV U11709 ( .A(n11564), .Z(n11992) );
  NOR U11710 ( .A(n11993), .B(n11992), .Z(n11568) );
  XOR U11711 ( .A(n11432), .B(n11431), .Z(n11433) );
  XOR U11712 ( .A(n11434), .B(n11433), .Z(n11561) );
  NOR U11713 ( .A(n106), .B(n47), .Z(n11560) );
  IV U11714 ( .A(n11560), .Z(n11435) );
  NOR U11715 ( .A(n11561), .B(n11435), .Z(n11563) );
  NOR U11716 ( .A(n105), .B(n47), .Z(n11555) );
  XOR U11717 ( .A(n11437), .B(n11436), .Z(n11554) );
  NOR U11718 ( .A(n11555), .B(n11554), .Z(n11558) );
  XOR U11719 ( .A(n11439), .B(n11438), .Z(n11440) );
  IV U11720 ( .A(n11440), .Z(n11549) );
  NOR U11721 ( .A(n104), .B(n47), .Z(n11550) );
  IV U11722 ( .A(n11550), .Z(n11441) );
  NOR U11723 ( .A(n11549), .B(n11441), .Z(n11552) );
  NOR U11724 ( .A(n89), .B(n47), .Z(n11546) );
  IV U11725 ( .A(n11546), .Z(n11445) );
  IV U11726 ( .A(n11442), .Z(n11444) );
  XOR U11727 ( .A(n11444), .B(n11443), .Z(n11545) );
  NOR U11728 ( .A(n11445), .B(n11545), .Z(n11548) );
  NOR U11729 ( .A(n90), .B(n47), .Z(n11448) );
  XOR U11730 ( .A(n11447), .B(n11446), .Z(n11449) );
  NOR U11731 ( .A(n11448), .B(n11449), .Z(n11535) );
  IV U11732 ( .A(n11448), .Z(n12007) );
  IV U11733 ( .A(n11449), .Z(n12006) );
  NOR U11734 ( .A(n12007), .B(n12006), .Z(n11533) );
  XOR U11735 ( .A(n11451), .B(n11450), .Z(n11452) );
  XOR U11736 ( .A(n11453), .B(n11452), .Z(n11528) );
  NOR U11737 ( .A(n102), .B(n47), .Z(n11529) );
  IV U11738 ( .A(n11529), .Z(n11454) );
  NOR U11739 ( .A(n11528), .B(n11454), .Z(n11531) );
  XOR U11740 ( .A(n11456), .B(n11455), .Z(n11525) );
  NOR U11741 ( .A(n101), .B(n47), .Z(n11524) );
  IV U11742 ( .A(n11524), .Z(n11457) );
  NOR U11743 ( .A(n11525), .B(n11457), .Z(n11527) );
  XOR U11744 ( .A(n11459), .B(n11458), .Z(n11521) );
  NOR U11745 ( .A(n100), .B(n47), .Z(n11520) );
  IV U11746 ( .A(n11520), .Z(n11460) );
  NOR U11747 ( .A(n11521), .B(n11460), .Z(n11523) );
  IV U11748 ( .A(n11461), .Z(n11463) );
  XOR U11749 ( .A(n11463), .B(n11462), .Z(n11516) );
  NOR U11750 ( .A(n99), .B(n47), .Z(n11517) );
  IV U11751 ( .A(n11517), .Z(n11464) );
  NOR U11752 ( .A(n11516), .B(n11464), .Z(n11519) );
  IV U11753 ( .A(n11465), .Z(n11467) );
  XOR U11754 ( .A(n11467), .B(n11466), .Z(n11512) );
  NOR U11755 ( .A(n98), .B(n47), .Z(n11513) );
  IV U11756 ( .A(n11513), .Z(n11468) );
  NOR U11757 ( .A(n11512), .B(n11468), .Z(n11515) );
  IV U11758 ( .A(n11469), .Z(n11471) );
  XOR U11759 ( .A(n11471), .B(n11470), .Z(n11508) );
  NOR U11760 ( .A(n91), .B(n47), .Z(n11509) );
  IV U11761 ( .A(n11509), .Z(n11472) );
  NOR U11762 ( .A(n11508), .B(n11472), .Z(n11511) );
  IV U11763 ( .A(n11473), .Z(n11475) );
  XOR U11764 ( .A(n11475), .B(n11474), .Z(n11504) );
  NOR U11765 ( .A(n97), .B(n47), .Z(n11505) );
  IV U11766 ( .A(n11505), .Z(n11476) );
  NOR U11767 ( .A(n11504), .B(n11476), .Z(n11507) );
  IV U11768 ( .A(n11477), .Z(n11479) );
  XOR U11769 ( .A(n11479), .B(n11478), .Z(n11500) );
  NOR U11770 ( .A(n96), .B(n47), .Z(n11501) );
  IV U11771 ( .A(n11501), .Z(n11480) );
  NOR U11772 ( .A(n11500), .B(n11480), .Z(n11503) );
  NOR U11773 ( .A(n95), .B(n47), .Z(n11497) );
  IV U11774 ( .A(n11497), .Z(n11483) );
  XOR U11775 ( .A(n11482), .B(n11481), .Z(n11496) );
  NOR U11776 ( .A(n11483), .B(n11496), .Z(n11499) );
  NOR U11777 ( .A(n93), .B(n47), .Z(n12558) );
  IV U11778 ( .A(n12558), .Z(n11484) );
  NOR U11779 ( .A(n46), .B(n168), .Z(n11492) );
  IV U11780 ( .A(n11492), .Z(n11487) );
  NOR U11781 ( .A(n11484), .B(n11487), .Z(n11485) );
  IV U11782 ( .A(n11485), .Z(n11486) );
  NOR U11783 ( .A(n94), .B(n11486), .Z(n11495) );
  NOR U11784 ( .A(n11487), .B(n93), .Z(n11488) );
  XOR U11785 ( .A(n94), .B(n11488), .Z(n11489) );
  NOR U11786 ( .A(n47), .B(n11489), .Z(n11490) );
  IV U11787 ( .A(n11490), .Z(n12044) );
  XOR U11788 ( .A(n11492), .B(n11491), .Z(n12043) );
  IV U11789 ( .A(n12043), .Z(n11493) );
  NOR U11790 ( .A(n12044), .B(n11493), .Z(n11494) );
  NOR U11791 ( .A(n11495), .B(n11494), .Z(n12040) );
  XOR U11792 ( .A(n11497), .B(n11496), .Z(n12039) );
  NOR U11793 ( .A(n12040), .B(n12039), .Z(n11498) );
  NOR U11794 ( .A(n11499), .B(n11498), .Z(n12035) );
  XOR U11795 ( .A(n11501), .B(n11500), .Z(n12036) );
  NOR U11796 ( .A(n12035), .B(n12036), .Z(n11502) );
  NOR U11797 ( .A(n11503), .B(n11502), .Z(n12031) );
  XOR U11798 ( .A(n11505), .B(n11504), .Z(n12032) );
  NOR U11799 ( .A(n12031), .B(n12032), .Z(n11506) );
  NOR U11800 ( .A(n11507), .B(n11506), .Z(n12027) );
  XOR U11801 ( .A(n11509), .B(n11508), .Z(n12028) );
  NOR U11802 ( .A(n12027), .B(n12028), .Z(n11510) );
  NOR U11803 ( .A(n11511), .B(n11510), .Z(n12023) );
  XOR U11804 ( .A(n11513), .B(n11512), .Z(n12024) );
  NOR U11805 ( .A(n12023), .B(n12024), .Z(n11514) );
  NOR U11806 ( .A(n11515), .B(n11514), .Z(n12019) );
  XOR U11807 ( .A(n11517), .B(n11516), .Z(n12020) );
  NOR U11808 ( .A(n12019), .B(n12020), .Z(n11518) );
  NOR U11809 ( .A(n11519), .B(n11518), .Z(n12018) );
  XOR U11810 ( .A(n11521), .B(n11520), .Z(n12017) );
  NOR U11811 ( .A(n12018), .B(n12017), .Z(n11522) );
  NOR U11812 ( .A(n11523), .B(n11522), .Z(n12013) );
  XOR U11813 ( .A(n11525), .B(n11524), .Z(n12014) );
  NOR U11814 ( .A(n12013), .B(n12014), .Z(n11526) );
  NOR U11815 ( .A(n11527), .B(n11526), .Z(n12012) );
  XOR U11816 ( .A(n11529), .B(n11528), .Z(n12011) );
  NOR U11817 ( .A(n12012), .B(n12011), .Z(n11530) );
  NOR U11818 ( .A(n11531), .B(n11530), .Z(n12009) );
  IV U11819 ( .A(n12009), .Z(n11532) );
  NOR U11820 ( .A(n11533), .B(n11532), .Z(n11534) );
  NOR U11821 ( .A(n11535), .B(n11534), .Z(n11542) );
  IV U11822 ( .A(n11542), .Z(n11537) );
  NOR U11823 ( .A(n103), .B(n47), .Z(n11536) );
  IV U11824 ( .A(n11536), .Z(n11541) );
  NOR U11825 ( .A(n11537), .B(n11541), .Z(n11544) );
  IV U11826 ( .A(n11538), .Z(n11540) );
  XOR U11827 ( .A(n11540), .B(n11539), .Z(n12005) );
  XOR U11828 ( .A(n11542), .B(n11541), .Z(n12004) );
  NOR U11829 ( .A(n12005), .B(n12004), .Z(n11543) );
  NOR U11830 ( .A(n11544), .B(n11543), .Z(n12116) );
  XOR U11831 ( .A(n11546), .B(n11545), .Z(n12117) );
  NOR U11832 ( .A(n12116), .B(n12117), .Z(n11547) );
  NOR U11833 ( .A(n11548), .B(n11547), .Z(n12003) );
  XOR U11834 ( .A(n11550), .B(n11549), .Z(n12002) );
  NOR U11835 ( .A(n12003), .B(n12002), .Z(n11551) );
  NOR U11836 ( .A(n11552), .B(n11551), .Z(n11553) );
  IV U11837 ( .A(n11553), .Z(n12000) );
  XOR U11838 ( .A(n11555), .B(n11554), .Z(n11556) );
  IV U11839 ( .A(n11556), .Z(n11999) );
  NOR U11840 ( .A(n12000), .B(n11999), .Z(n11557) );
  NOR U11841 ( .A(n11558), .B(n11557), .Z(n11559) );
  IV U11842 ( .A(n11559), .Z(n11998) );
  XOR U11843 ( .A(n11561), .B(n11560), .Z(n11997) );
  NOR U11844 ( .A(n11998), .B(n11997), .Z(n11562) );
  NOR U11845 ( .A(n11563), .B(n11562), .Z(n11995) );
  NOR U11846 ( .A(n11565), .B(n11564), .Z(n11566) );
  NOR U11847 ( .A(n11995), .B(n11566), .Z(n11567) );
  NOR U11848 ( .A(n11568), .B(n11567), .Z(n11575) );
  NOR U11849 ( .A(n107), .B(n47), .Z(n11574) );
  IV U11850 ( .A(n11574), .Z(n11569) );
  NOR U11851 ( .A(n11575), .B(n11569), .Z(n11577) );
  XOR U11852 ( .A(n11571), .B(n11570), .Z(n11572) );
  XOR U11853 ( .A(n11573), .B(n11572), .Z(n11989) );
  XOR U11854 ( .A(n11575), .B(n11574), .Z(n11988) );
  NOR U11855 ( .A(n11989), .B(n11988), .Z(n11576) );
  NOR U11856 ( .A(n11577), .B(n11576), .Z(n11578) );
  IV U11857 ( .A(n11578), .Z(n12151) );
  NOR U11858 ( .A(n11579), .B(n12151), .Z(n11580) );
  NOR U11859 ( .A(n11581), .B(n11580), .Z(n11585) );
  IV U11860 ( .A(n11585), .Z(n11582) );
  NOR U11861 ( .A(n11586), .B(n11582), .Z(n11588) );
  XOR U11862 ( .A(n11584), .B(n11583), .Z(n11984) );
  XOR U11863 ( .A(n11586), .B(n11585), .Z(n11985) );
  NOR U11864 ( .A(n11984), .B(n11985), .Z(n11587) );
  NOR U11865 ( .A(n11588), .B(n11587), .Z(n11982) );
  IV U11866 ( .A(n11982), .Z(n11589) );
  NOR U11867 ( .A(n11590), .B(n11589), .Z(n11591) );
  NOR U11868 ( .A(n11592), .B(n11591), .Z(n11593) );
  IV U11869 ( .A(n11593), .Z(n11600) );
  NOR U11870 ( .A(n110), .B(n47), .Z(n11599) );
  IV U11871 ( .A(n11599), .Z(n11594) );
  NOR U11872 ( .A(n11600), .B(n11594), .Z(n11602) );
  XOR U11873 ( .A(n11596), .B(n11595), .Z(n11597) );
  XOR U11874 ( .A(n11598), .B(n11597), .Z(n11975) );
  XOR U11875 ( .A(n11600), .B(n11599), .Z(n11976) );
  NOR U11876 ( .A(n11975), .B(n11976), .Z(n11601) );
  NOR U11877 ( .A(n11602), .B(n11601), .Z(n12176) );
  NOR U11878 ( .A(n11604), .B(n11603), .Z(n11605) );
  NOR U11879 ( .A(n12176), .B(n11605), .Z(n11606) );
  NOR U11880 ( .A(n11607), .B(n11606), .Z(n11614) );
  NOR U11881 ( .A(n111), .B(n47), .Z(n11613) );
  IV U11882 ( .A(n11613), .Z(n11608) );
  NOR U11883 ( .A(n11614), .B(n11608), .Z(n11616) );
  XOR U11884 ( .A(n11610), .B(n11609), .Z(n11611) );
  XOR U11885 ( .A(n11612), .B(n11611), .Z(n11972) );
  XOR U11886 ( .A(n11614), .B(n11613), .Z(n11971) );
  NOR U11887 ( .A(n11972), .B(n11971), .Z(n11615) );
  NOR U11888 ( .A(n11616), .B(n11615), .Z(n12187) );
  NOR U11889 ( .A(n11617), .B(n12187), .Z(n11618) );
  NOR U11890 ( .A(n11619), .B(n11618), .Z(n11622) );
  NOR U11891 ( .A(n112), .B(n47), .Z(n11621) );
  IV U11892 ( .A(n11621), .Z(n11620) );
  NOR U11893 ( .A(n11622), .B(n11620), .Z(n11628) );
  XOR U11894 ( .A(n11622), .B(n11621), .Z(n11968) );
  XOR U11895 ( .A(n11624), .B(n11623), .Z(n11625) );
  XOR U11896 ( .A(n11626), .B(n11625), .Z(n11967) );
  NOR U11897 ( .A(n11968), .B(n11967), .Z(n11627) );
  NOR U11898 ( .A(n11628), .B(n11627), .Z(n11963) );
  IV U11899 ( .A(n11963), .Z(n11629) );
  NOR U11900 ( .A(n11630), .B(n11629), .Z(n11631) );
  NOR U11901 ( .A(n11632), .B(n11631), .Z(n11638) );
  IV U11902 ( .A(n11638), .Z(n11633) );
  NOR U11903 ( .A(n11639), .B(n11633), .Z(n11641) );
  XOR U11904 ( .A(n11635), .B(n11634), .Z(n11636) );
  XOR U11905 ( .A(n11637), .B(n11636), .Z(n11956) );
  XOR U11906 ( .A(n11639), .B(n11638), .Z(n11957) );
  NOR U11907 ( .A(n11956), .B(n11957), .Z(n11640) );
  NOR U11908 ( .A(n11641), .B(n11640), .Z(n11642) );
  IV U11909 ( .A(n11642), .Z(n12207) );
  NOR U11910 ( .A(n12208), .B(n12207), .Z(n11643) );
  NOR U11911 ( .A(n11644), .B(n11643), .Z(n11645) );
  IV U11912 ( .A(n11645), .Z(n11650) );
  NOR U11913 ( .A(n114), .B(n47), .Z(n11649) );
  IV U11914 ( .A(n11649), .Z(n11646) );
  NOR U11915 ( .A(n11650), .B(n11646), .Z(n11652) );
  XOR U11916 ( .A(n11648), .B(n11647), .Z(n11952) );
  XOR U11917 ( .A(n11650), .B(n11649), .Z(n11953) );
  NOR U11918 ( .A(n11952), .B(n11953), .Z(n11651) );
  NOR U11919 ( .A(n11652), .B(n11651), .Z(n11654) );
  IV U11920 ( .A(n11654), .Z(n12218) );
  NOR U11921 ( .A(n11653), .B(n12218), .Z(n11661) );
  IV U11922 ( .A(n11653), .Z(n12219) );
  NOR U11923 ( .A(n11654), .B(n12219), .Z(n11659) );
  XOR U11924 ( .A(n11656), .B(n11655), .Z(n11657) );
  XOR U11925 ( .A(n11658), .B(n11657), .Z(n12221) );
  NOR U11926 ( .A(n11659), .B(n12221), .Z(n11660) );
  NOR U11927 ( .A(n11661), .B(n11660), .Z(n11669) );
  IV U11928 ( .A(n11669), .Z(n11663) );
  NOR U11929 ( .A(n115), .B(n47), .Z(n11662) );
  IV U11930 ( .A(n11662), .Z(n11668) );
  NOR U11931 ( .A(n11663), .B(n11668), .Z(n11671) );
  XOR U11932 ( .A(n11665), .B(n11664), .Z(n11666) );
  XOR U11933 ( .A(n11667), .B(n11666), .Z(n11947) );
  XOR U11934 ( .A(n11669), .B(n11668), .Z(n11948) );
  NOR U11935 ( .A(n11947), .B(n11948), .Z(n11670) );
  NOR U11936 ( .A(n11671), .B(n11670), .Z(n11673) );
  NOR U11937 ( .A(n11672), .B(n11673), .Z(n11677) );
  IV U11938 ( .A(n11673), .Z(n12233) );
  NOR U11939 ( .A(n12235), .B(n12233), .Z(n11675) );
  NOR U11940 ( .A(n81), .B(n47), .Z(n11674) );
  IV U11941 ( .A(n11674), .Z(n12232) );
  NOR U11942 ( .A(n11675), .B(n12232), .Z(n11676) );
  NOR U11943 ( .A(n11677), .B(n11676), .Z(n11678) );
  NOR U11944 ( .A(n116), .B(n47), .Z(n11679) );
  IV U11945 ( .A(n11679), .Z(n12240) );
  NOR U11946 ( .A(n11678), .B(n12240), .Z(n11686) );
  IV U11947 ( .A(n11678), .Z(n12241) );
  NOR U11948 ( .A(n11679), .B(n12241), .Z(n11684) );
  XOR U11949 ( .A(n11681), .B(n11680), .Z(n11682) );
  XOR U11950 ( .A(n11683), .B(n11682), .Z(n12243) );
  NOR U11951 ( .A(n11684), .B(n12243), .Z(n11685) );
  NOR U11952 ( .A(n11686), .B(n11685), .Z(n11689) );
  XOR U11953 ( .A(n11688), .B(n11687), .Z(n11690) );
  NOR U11954 ( .A(n11689), .B(n11690), .Z(n11694) );
  IV U11955 ( .A(n11689), .Z(n11691) );
  XOR U11956 ( .A(n11691), .B(n11690), .Z(n11944) );
  NOR U11957 ( .A(n80), .B(n47), .Z(n11945) );
  IV U11958 ( .A(n11945), .Z(n11692) );
  NOR U11959 ( .A(n11944), .B(n11692), .Z(n11693) );
  NOR U11960 ( .A(n11694), .B(n11693), .Z(n12258) );
  IV U11961 ( .A(n12258), .Z(n11695) );
  NOR U11962 ( .A(n11696), .B(n11695), .Z(n11697) );
  NOR U11963 ( .A(n11698), .B(n11697), .Z(n11704) );
  IV U11964 ( .A(n11704), .Z(n11700) );
  NOR U11965 ( .A(n79), .B(n47), .Z(n11699) );
  IV U11966 ( .A(n11699), .Z(n11703) );
  NOR U11967 ( .A(n11700), .B(n11703), .Z(n11706) );
  XOR U11968 ( .A(n11702), .B(n11701), .Z(n12264) );
  XOR U11969 ( .A(n11704), .B(n11703), .Z(n12263) );
  NOR U11970 ( .A(n12264), .B(n12263), .Z(n11705) );
  NOR U11971 ( .A(n11706), .B(n11705), .Z(n11711) );
  NOR U11972 ( .A(n119), .B(n47), .Z(n11710) );
  IV U11973 ( .A(n11710), .Z(n11707) );
  NOR U11974 ( .A(n11711), .B(n11707), .Z(n11713) );
  XOR U11975 ( .A(n11709), .B(n11708), .Z(n11941) );
  XOR U11976 ( .A(n11711), .B(n11710), .Z(n11940) );
  NOR U11977 ( .A(n11941), .B(n11940), .Z(n11712) );
  NOR U11978 ( .A(n11713), .B(n11712), .Z(n11716) );
  XOR U11979 ( .A(n11715), .B(n11714), .Z(n11717) );
  NOR U11980 ( .A(n11716), .B(n11717), .Z(n11721) );
  IV U11981 ( .A(n11716), .Z(n11718) );
  XOR U11982 ( .A(n11718), .B(n11717), .Z(n11937) );
  NOR U11983 ( .A(n120), .B(n47), .Z(n11938) );
  IV U11984 ( .A(n11938), .Z(n11719) );
  NOR U11985 ( .A(n11937), .B(n11719), .Z(n11720) );
  NOR U11986 ( .A(n11721), .B(n11720), .Z(n11724) );
  NOR U11987 ( .A(n123), .B(n47), .Z(n11723) );
  IV U11988 ( .A(n11723), .Z(n11722) );
  NOR U11989 ( .A(n11724), .B(n11722), .Z(n11729) );
  XOR U11990 ( .A(n11724), .B(n11723), .Z(n12279) );
  XOR U11991 ( .A(n11726), .B(n11725), .Z(n12280) );
  IV U11992 ( .A(n12280), .Z(n11727) );
  NOR U11993 ( .A(n12279), .B(n11727), .Z(n11728) );
  NOR U11994 ( .A(n11729), .B(n11728), .Z(n11732) );
  NOR U11995 ( .A(n125), .B(n47), .Z(n11731) );
  IV U11996 ( .A(n11731), .Z(n11730) );
  NOR U11997 ( .A(n11732), .B(n11730), .Z(n11737) );
  XOR U11998 ( .A(n11732), .B(n11731), .Z(n11934) );
  XOR U11999 ( .A(n11734), .B(n11733), .Z(n11935) );
  IV U12000 ( .A(n11935), .Z(n11735) );
  NOR U12001 ( .A(n11934), .B(n11735), .Z(n11736) );
  NOR U12002 ( .A(n11737), .B(n11736), .Z(n12293) );
  XOR U12003 ( .A(n11739), .B(n11738), .Z(n12292) );
  NOR U12004 ( .A(n12293), .B(n12292), .Z(n11740) );
  NOR U12005 ( .A(n11741), .B(n11740), .Z(n11744) );
  NOR U12006 ( .A(n128), .B(n47), .Z(n11743) );
  IV U12007 ( .A(n11743), .Z(n11742) );
  NOR U12008 ( .A(n11744), .B(n11742), .Z(n11748) );
  XOR U12009 ( .A(n11744), .B(n11743), .Z(n12299) );
  XOR U12010 ( .A(n11746), .B(n11745), .Z(n12300) );
  NOR U12011 ( .A(n12299), .B(n12300), .Z(n11747) );
  NOR U12012 ( .A(n11748), .B(n11747), .Z(n11751) );
  NOR U12013 ( .A(n131), .B(n47), .Z(n11750) );
  IV U12014 ( .A(n11750), .Z(n11749) );
  NOR U12015 ( .A(n11751), .B(n11749), .Z(n11756) );
  XOR U12016 ( .A(n11751), .B(n11750), .Z(n11931) );
  XOR U12017 ( .A(n11753), .B(n11752), .Z(n11932) );
  IV U12018 ( .A(n11932), .Z(n11754) );
  NOR U12019 ( .A(n11931), .B(n11754), .Z(n11755) );
  NOR U12020 ( .A(n11756), .B(n11755), .Z(n11761) );
  XOR U12021 ( .A(n11758), .B(n11757), .Z(n11760) );
  IV U12022 ( .A(n11760), .Z(n11759) );
  NOR U12023 ( .A(n11761), .B(n11759), .Z(n11764) );
  XOR U12024 ( .A(n11761), .B(n11760), .Z(n12314) );
  NOR U12025 ( .A(n133), .B(n47), .Z(n12315) );
  IV U12026 ( .A(n12315), .Z(n11762) );
  NOR U12027 ( .A(n12314), .B(n11762), .Z(n11763) );
  NOR U12028 ( .A(n11764), .B(n11763), .Z(n11767) );
  NOR U12029 ( .A(n135), .B(n47), .Z(n11766) );
  IV U12030 ( .A(n11766), .Z(n11765) );
  NOR U12031 ( .A(n11767), .B(n11765), .Z(n11772) );
  XOR U12032 ( .A(n11767), .B(n11766), .Z(n12318) );
  XOR U12033 ( .A(n11769), .B(n11768), .Z(n12319) );
  IV U12034 ( .A(n12319), .Z(n11770) );
  NOR U12035 ( .A(n12318), .B(n11770), .Z(n11771) );
  NOR U12036 ( .A(n11772), .B(n11771), .Z(n11776) );
  XOR U12037 ( .A(n11774), .B(n11773), .Z(n11775) );
  NOR U12038 ( .A(n11776), .B(n11775), .Z(n11780) );
  XOR U12039 ( .A(n11776), .B(n11775), .Z(n11777) );
  IV U12040 ( .A(n11777), .Z(n11928) );
  NOR U12041 ( .A(n137), .B(n47), .Z(n11929) );
  IV U12042 ( .A(n11929), .Z(n11778) );
  NOR U12043 ( .A(n11928), .B(n11778), .Z(n11779) );
  NOR U12044 ( .A(n11780), .B(n11779), .Z(n11783) );
  XOR U12045 ( .A(n11782), .B(n11781), .Z(n11784) );
  NOR U12046 ( .A(n11783), .B(n11784), .Z(n11788) );
  IV U12047 ( .A(n11783), .Z(n11785) );
  XOR U12048 ( .A(n11785), .B(n11784), .Z(n11925) );
  NOR U12049 ( .A(n139), .B(n47), .Z(n11926) );
  IV U12050 ( .A(n11926), .Z(n11786) );
  NOR U12051 ( .A(n11925), .B(n11786), .Z(n11787) );
  NOR U12052 ( .A(n11788), .B(n11787), .Z(n11791) );
  NOR U12053 ( .A(n141), .B(n47), .Z(n11790) );
  IV U12054 ( .A(n11790), .Z(n11789) );
  NOR U12055 ( .A(n11791), .B(n11789), .Z(n11796) );
  XOR U12056 ( .A(n11791), .B(n11790), .Z(n12334) );
  XOR U12057 ( .A(n11793), .B(n11792), .Z(n12335) );
  IV U12058 ( .A(n12335), .Z(n11794) );
  NOR U12059 ( .A(n12334), .B(n11794), .Z(n11795) );
  NOR U12060 ( .A(n11796), .B(n11795), .Z(n11799) );
  NOR U12061 ( .A(n143), .B(n47), .Z(n11798) );
  IV U12062 ( .A(n11798), .Z(n11797) );
  NOR U12063 ( .A(n11799), .B(n11797), .Z(n11803) );
  XOR U12064 ( .A(n11799), .B(n11798), .Z(n11922) );
  XOR U12065 ( .A(n11801), .B(n11800), .Z(n11921) );
  NOR U12066 ( .A(n11922), .B(n11921), .Z(n11802) );
  NOR U12067 ( .A(n11803), .B(n11802), .Z(n11808) );
  XOR U12068 ( .A(n11805), .B(n11804), .Z(n11807) );
  IV U12069 ( .A(n11807), .Z(n11806) );
  NOR U12070 ( .A(n11808), .B(n11806), .Z(n11811) );
  XOR U12071 ( .A(n11808), .B(n11807), .Z(n11918) );
  NOR U12072 ( .A(n145), .B(n47), .Z(n11919) );
  IV U12073 ( .A(n11919), .Z(n11809) );
  NOR U12074 ( .A(n11918), .B(n11809), .Z(n11810) );
  NOR U12075 ( .A(n11811), .B(n11810), .Z(n11816) );
  XOR U12076 ( .A(n11813), .B(n11812), .Z(n11815) );
  IV U12077 ( .A(n11815), .Z(n11814) );
  NOR U12078 ( .A(n11816), .B(n11814), .Z(n11819) );
  XOR U12079 ( .A(n11816), .B(n11815), .Z(n12350) );
  NOR U12080 ( .A(n147), .B(n47), .Z(n12351) );
  IV U12081 ( .A(n12351), .Z(n11817) );
  NOR U12082 ( .A(n12350), .B(n11817), .Z(n11818) );
  NOR U12083 ( .A(n11819), .B(n11818), .Z(n11824) );
  XOR U12084 ( .A(n11821), .B(n11820), .Z(n11823) );
  IV U12085 ( .A(n11823), .Z(n11822) );
  NOR U12086 ( .A(n11824), .B(n11822), .Z(n11827) );
  XOR U12087 ( .A(n11824), .B(n11823), .Z(n11915) );
  NOR U12088 ( .A(n148), .B(n47), .Z(n11916) );
  IV U12089 ( .A(n11916), .Z(n11825) );
  NOR U12090 ( .A(n11915), .B(n11825), .Z(n11826) );
  NOR U12091 ( .A(n11827), .B(n11826), .Z(n12366) );
  XOR U12092 ( .A(n11829), .B(n11828), .Z(n12365) );
  NOR U12093 ( .A(n12366), .B(n12365), .Z(n11830) );
  NOR U12094 ( .A(n11831), .B(n11830), .Z(n11834) );
  NOR U12095 ( .A(n153), .B(n47), .Z(n11833) );
  IV U12096 ( .A(n11833), .Z(n11832) );
  NOR U12097 ( .A(n11834), .B(n11832), .Z(n11838) );
  XOR U12098 ( .A(n11834), .B(n11833), .Z(n12370) );
  XOR U12099 ( .A(n11836), .B(n11835), .Z(n12371) );
  NOR U12100 ( .A(n12370), .B(n12371), .Z(n11837) );
  NOR U12101 ( .A(n11838), .B(n11837), .Z(n11841) );
  NOR U12102 ( .A(n155), .B(n47), .Z(n11840) );
  IV U12103 ( .A(n11840), .Z(n11839) );
  NOR U12104 ( .A(n11841), .B(n11839), .Z(n11846) );
  XOR U12105 ( .A(n11841), .B(n11840), .Z(n11912) );
  XOR U12106 ( .A(n11843), .B(n11842), .Z(n11913) );
  IV U12107 ( .A(n11913), .Z(n11844) );
  NOR U12108 ( .A(n11912), .B(n11844), .Z(n11845) );
  NOR U12109 ( .A(n11846), .B(n11845), .Z(n11850) );
  XOR U12110 ( .A(n11848), .B(n11847), .Z(n11849) );
  NOR U12111 ( .A(n11850), .B(n11849), .Z(n11854) );
  XOR U12112 ( .A(n11850), .B(n11849), .Z(n11851) );
  IV U12113 ( .A(n11851), .Z(n12385) );
  NOR U12114 ( .A(n156), .B(n47), .Z(n12386) );
  IV U12115 ( .A(n12386), .Z(n11852) );
  NOR U12116 ( .A(n12385), .B(n11852), .Z(n11853) );
  NOR U12117 ( .A(n11854), .B(n11853), .Z(n11857) );
  NOR U12118 ( .A(n158), .B(n47), .Z(n11856) );
  IV U12119 ( .A(n11856), .Z(n11855) );
  NOR U12120 ( .A(n11857), .B(n11855), .Z(n11862) );
  XOR U12121 ( .A(n11857), .B(n11856), .Z(n12389) );
  XOR U12122 ( .A(n11859), .B(n11858), .Z(n12390) );
  IV U12123 ( .A(n12390), .Z(n11860) );
  NOR U12124 ( .A(n12389), .B(n11860), .Z(n11861) );
  NOR U12125 ( .A(n11862), .B(n11861), .Z(n11866) );
  XOR U12126 ( .A(n11864), .B(n11863), .Z(n11865) );
  NOR U12127 ( .A(n11866), .B(n11865), .Z(n11870) );
  XOR U12128 ( .A(n11866), .B(n11865), .Z(n11867) );
  IV U12129 ( .A(n11867), .Z(n11909) );
  NOR U12130 ( .A(n161), .B(n47), .Z(n11910) );
  IV U12131 ( .A(n11910), .Z(n11868) );
  NOR U12132 ( .A(n11909), .B(n11868), .Z(n11869) );
  NOR U12133 ( .A(n11870), .B(n11869), .Z(n12402) );
  XOR U12134 ( .A(n11872), .B(n11871), .Z(n12401) );
  NOR U12135 ( .A(n12402), .B(n12401), .Z(n11873) );
  NOR U12136 ( .A(n11874), .B(n11873), .Z(n11879) );
  NOR U12137 ( .A(n165), .B(n47), .Z(n11878) );
  IV U12138 ( .A(n11878), .Z(n11875) );
  NOR U12139 ( .A(n11879), .B(n11875), .Z(n11882) );
  XOR U12140 ( .A(n11877), .B(n11876), .Z(n12410) );
  IV U12141 ( .A(n12410), .Z(n11880) );
  XOR U12142 ( .A(n11879), .B(n11878), .Z(n12409) );
  NOR U12143 ( .A(n11880), .B(n12409), .Z(n11881) );
  NOR U12144 ( .A(n11882), .B(n11881), .Z(n11887) );
  XOR U12145 ( .A(n11884), .B(n11883), .Z(n11886) );
  IV U12146 ( .A(n11886), .Z(n11885) );
  NOR U12147 ( .A(n11887), .B(n11885), .Z(n11890) );
  XOR U12148 ( .A(n11887), .B(n11886), .Z(n12417) );
  NOR U12149 ( .A(n167), .B(n47), .Z(n12418) );
  IV U12150 ( .A(n12418), .Z(n11888) );
  NOR U12151 ( .A(n12417), .B(n11888), .Z(n11889) );
  NOR U12152 ( .A(n11890), .B(n11889), .Z(n12420) );
  XOR U12153 ( .A(n11892), .B(n11891), .Z(n12419) );
  NOR U12154 ( .A(n12420), .B(n12419), .Z(n11908) );
  IV U12155 ( .A(n11908), .Z(n31669) );
  XOR U12156 ( .A(n11894), .B(n11893), .Z(n31661) );
  NOR U12157 ( .A(n31669), .B(n31661), .Z(n11895) );
  NOR U12158 ( .A(n31664), .B(n11895), .Z(n31670) );
  IV U12159 ( .A(n11896), .Z(n11897) );
  NOR U12160 ( .A(n11898), .B(n11897), .Z(n11903) );
  IV U12161 ( .A(n11899), .Z(n11900) );
  NOR U12162 ( .A(n11901), .B(n11900), .Z(n11902) );
  NOR U12163 ( .A(n11903), .B(n11902), .Z(n28632) );
  XOR U12164 ( .A(n11905), .B(n11904), .Z(n28631) );
  XOR U12165 ( .A(n28632), .B(n28631), .Z(n11906) );
  IV U12166 ( .A(n11906), .Z(n31676) );
  NOR U12167 ( .A(n31670), .B(n31676), .Z(n28639) );
  NOR U12168 ( .A(n31664), .B(n11906), .Z(n28630) );
  IV U12169 ( .A(n31661), .Z(n11907) );
  NOR U12170 ( .A(n11908), .B(n11907), .Z(n28628) );
  XOR U12171 ( .A(n11910), .B(n11909), .Z(n12397) );
  NOR U12172 ( .A(n163), .B(n48), .Z(n12398) );
  IV U12173 ( .A(n12398), .Z(n11911) );
  NOR U12174 ( .A(n12397), .B(n11911), .Z(n12400) );
  XOR U12175 ( .A(n11913), .B(n11912), .Z(n12378) );
  NOR U12176 ( .A(n156), .B(n48), .Z(n12379) );
  IV U12177 ( .A(n12379), .Z(n11914) );
  NOR U12178 ( .A(n12378), .B(n11914), .Z(n12381) );
  XOR U12179 ( .A(n11916), .B(n11915), .Z(n12358) );
  NOR U12180 ( .A(n150), .B(n48), .Z(n12359) );
  IV U12181 ( .A(n12359), .Z(n11917) );
  NOR U12182 ( .A(n12358), .B(n11917), .Z(n12361) );
  XOR U12183 ( .A(n11919), .B(n11918), .Z(n12346) );
  NOR U12184 ( .A(n147), .B(n48), .Z(n12347) );
  IV U12185 ( .A(n12347), .Z(n11920) );
  NOR U12186 ( .A(n12346), .B(n11920), .Z(n12349) );
  IV U12187 ( .A(n11921), .Z(n11923) );
  XOR U12188 ( .A(n11923), .B(n11922), .Z(n12342) );
  NOR U12189 ( .A(n145), .B(n48), .Z(n12343) );
  IV U12190 ( .A(n12343), .Z(n11924) );
  NOR U12191 ( .A(n12342), .B(n11924), .Z(n12345) );
  XOR U12192 ( .A(n11926), .B(n11925), .Z(n12330) );
  NOR U12193 ( .A(n141), .B(n48), .Z(n12331) );
  IV U12194 ( .A(n12331), .Z(n11927) );
  NOR U12195 ( .A(n12330), .B(n11927), .Z(n12333) );
  XOR U12196 ( .A(n11929), .B(n11928), .Z(n12326) );
  NOR U12197 ( .A(n139), .B(n48), .Z(n12327) );
  IV U12198 ( .A(n12327), .Z(n11930) );
  NOR U12199 ( .A(n12326), .B(n11930), .Z(n12329) );
  XOR U12200 ( .A(n11932), .B(n11931), .Z(n12307) );
  NOR U12201 ( .A(n133), .B(n48), .Z(n12308) );
  IV U12202 ( .A(n12308), .Z(n11933) );
  NOR U12203 ( .A(n12307), .B(n11933), .Z(n12310) );
  XOR U12204 ( .A(n11935), .B(n11934), .Z(n12287) );
  NOR U12205 ( .A(n126), .B(n48), .Z(n12288) );
  IV U12206 ( .A(n12288), .Z(n11936) );
  NOR U12207 ( .A(n12287), .B(n11936), .Z(n12290) );
  XOR U12208 ( .A(n11938), .B(n11937), .Z(n12275) );
  NOR U12209 ( .A(n123), .B(n48), .Z(n12276) );
  IV U12210 ( .A(n12276), .Z(n11939) );
  NOR U12211 ( .A(n12275), .B(n11939), .Z(n12278) );
  XOR U12212 ( .A(n11941), .B(n11940), .Z(n12271) );
  IV U12213 ( .A(n12271), .Z(n11943) );
  NOR U12214 ( .A(n120), .B(n48), .Z(n11942) );
  IV U12215 ( .A(n11942), .Z(n12272) );
  NOR U12216 ( .A(n11943), .B(n12272), .Z(n12274) );
  XOR U12217 ( .A(n11945), .B(n11944), .Z(n12250) );
  NOR U12218 ( .A(n117), .B(n48), .Z(n12251) );
  IV U12219 ( .A(n12251), .Z(n11946) );
  NOR U12220 ( .A(n12250), .B(n11946), .Z(n12253) );
  XOR U12221 ( .A(n11948), .B(n11947), .Z(n11950) );
  IV U12222 ( .A(n11950), .Z(n12715) );
  NOR U12223 ( .A(n81), .B(n48), .Z(n11949) );
  IV U12224 ( .A(n11949), .Z(n12714) );
  NOR U12225 ( .A(n12715), .B(n12714), .Z(n12230) );
  NOR U12226 ( .A(n11950), .B(n11949), .Z(n12228) );
  NOR U12227 ( .A(n82), .B(n48), .Z(n11951) );
  IV U12228 ( .A(n11951), .Z(n12214) );
  XOR U12229 ( .A(n11953), .B(n11952), .Z(n11954) );
  IV U12230 ( .A(n11954), .Z(n12213) );
  NOR U12231 ( .A(n12214), .B(n12213), .Z(n12217) );
  NOR U12232 ( .A(n114), .B(n48), .Z(n11955) );
  IV U12233 ( .A(n11955), .Z(n12210) );
  XOR U12234 ( .A(n11957), .B(n11956), .Z(n11958) );
  NOR U12235 ( .A(n83), .B(n48), .Z(n11959) );
  NOR U12236 ( .A(n11958), .B(n11959), .Z(n12205) );
  IV U12237 ( .A(n11958), .Z(n12461) );
  IV U12238 ( .A(n11959), .Z(n12460) );
  NOR U12239 ( .A(n12461), .B(n12460), .Z(n12203) );
  XOR U12240 ( .A(n11961), .B(n11960), .Z(n11962) );
  XOR U12241 ( .A(n11963), .B(n11962), .Z(n11966) );
  NOR U12242 ( .A(n113), .B(n48), .Z(n11965) );
  IV U12243 ( .A(n11965), .Z(n11964) );
  NOR U12244 ( .A(n11966), .B(n11964), .Z(n12201) );
  XOR U12245 ( .A(n11966), .B(n11965), .Z(n12465) );
  XOR U12246 ( .A(n11968), .B(n11967), .Z(n11969) );
  NOR U12247 ( .A(n84), .B(n48), .Z(n11970) );
  NOR U12248 ( .A(n11969), .B(n11970), .Z(n12198) );
  XOR U12249 ( .A(n11970), .B(n11969), .Z(n12683) );
  IV U12250 ( .A(n12683), .Z(n12196) );
  XOR U12251 ( .A(n11972), .B(n11971), .Z(n11973) );
  NOR U12252 ( .A(n85), .B(n48), .Z(n11974) );
  NOR U12253 ( .A(n11973), .B(n11974), .Z(n12184) );
  IV U12254 ( .A(n11973), .Z(n12669) );
  IV U12255 ( .A(n11974), .Z(n12668) );
  NOR U12256 ( .A(n12669), .B(n12668), .Z(n12182) );
  NOR U12257 ( .A(n111), .B(n48), .Z(n12178) );
  IV U12258 ( .A(n12178), .Z(n12172) );
  XOR U12259 ( .A(n11976), .B(n11975), .Z(n11977) );
  NOR U12260 ( .A(n86), .B(n48), .Z(n11978) );
  NOR U12261 ( .A(n11977), .B(n11978), .Z(n12170) );
  IV U12262 ( .A(n11977), .Z(n12475) );
  IV U12263 ( .A(n11978), .Z(n12474) );
  NOR U12264 ( .A(n12475), .B(n12474), .Z(n12168) );
  XOR U12265 ( .A(n11980), .B(n11979), .Z(n11981) );
  XOR U12266 ( .A(n11982), .B(n11981), .Z(n12164) );
  NOR U12267 ( .A(n110), .B(n48), .Z(n12163) );
  IV U12268 ( .A(n12163), .Z(n11983) );
  NOR U12269 ( .A(n12164), .B(n11983), .Z(n12166) );
  NOR U12270 ( .A(n109), .B(n48), .Z(n12160) );
  IV U12271 ( .A(n12160), .Z(n11987) );
  XOR U12272 ( .A(n11985), .B(n11984), .Z(n11986) );
  IV U12273 ( .A(n11986), .Z(n12159) );
  NOR U12274 ( .A(n11987), .B(n12159), .Z(n12162) );
  XOR U12275 ( .A(n11989), .B(n11988), .Z(n11990) );
  NOR U12276 ( .A(n87), .B(n48), .Z(n11991) );
  NOR U12277 ( .A(n11990), .B(n11991), .Z(n12148) );
  IV U12278 ( .A(n11990), .Z(n12492) );
  IV U12279 ( .A(n11991), .Z(n12491) );
  NOR U12280 ( .A(n12492), .B(n12491), .Z(n12146) );
  XOR U12281 ( .A(n11993), .B(n11992), .Z(n11994) );
  XOR U12282 ( .A(n11995), .B(n11994), .Z(n12141) );
  NOR U12283 ( .A(n107), .B(n48), .Z(n12140) );
  IV U12284 ( .A(n12140), .Z(n11996) );
  NOR U12285 ( .A(n12141), .B(n11996), .Z(n12144) );
  NOR U12286 ( .A(n88), .B(n48), .Z(n12134) );
  XOR U12287 ( .A(n11998), .B(n11997), .Z(n12135) );
  NOR U12288 ( .A(n12134), .B(n12135), .Z(n12139) );
  XOR U12289 ( .A(n12000), .B(n11999), .Z(n12130) );
  NOR U12290 ( .A(n106), .B(n48), .Z(n12129) );
  IV U12291 ( .A(n12129), .Z(n12001) );
  NOR U12292 ( .A(n12130), .B(n12001), .Z(n12133) );
  NOR U12293 ( .A(n105), .B(n48), .Z(n12125) );
  XOR U12294 ( .A(n12003), .B(n12002), .Z(n12124) );
  NOR U12295 ( .A(n12125), .B(n12124), .Z(n12128) );
  NOR U12296 ( .A(n104), .B(n48), .Z(n12120) );
  IV U12297 ( .A(n12120), .Z(n12115) );
  NOR U12298 ( .A(n89), .B(n48), .Z(n12110) );
  XOR U12299 ( .A(n12005), .B(n12004), .Z(n12109) );
  NOR U12300 ( .A(n12110), .B(n12109), .Z(n12113) );
  XOR U12301 ( .A(n12007), .B(n12006), .Z(n12008) );
  XOR U12302 ( .A(n12009), .B(n12008), .Z(n12104) );
  NOR U12303 ( .A(n103), .B(n48), .Z(n12103) );
  IV U12304 ( .A(n12103), .Z(n12010) );
  NOR U12305 ( .A(n12104), .B(n12010), .Z(n12107) );
  NOR U12306 ( .A(n90), .B(n48), .Z(n12099) );
  XOR U12307 ( .A(n12012), .B(n12011), .Z(n12098) );
  NOR U12308 ( .A(n12099), .B(n12098), .Z(n12102) );
  IV U12309 ( .A(n12013), .Z(n12015) );
  XOR U12310 ( .A(n12015), .B(n12014), .Z(n12092) );
  NOR U12311 ( .A(n102), .B(n48), .Z(n12093) );
  IV U12312 ( .A(n12093), .Z(n12016) );
  NOR U12313 ( .A(n12092), .B(n12016), .Z(n12096) );
  NOR U12314 ( .A(n101), .B(n48), .Z(n12088) );
  XOR U12315 ( .A(n12018), .B(n12017), .Z(n12087) );
  NOR U12316 ( .A(n12088), .B(n12087), .Z(n12091) );
  IV U12317 ( .A(n12019), .Z(n12021) );
  XOR U12318 ( .A(n12021), .B(n12020), .Z(n12082) );
  NOR U12319 ( .A(n100), .B(n48), .Z(n12083) );
  IV U12320 ( .A(n12083), .Z(n12022) );
  NOR U12321 ( .A(n12082), .B(n12022), .Z(n12085) );
  IV U12322 ( .A(n12023), .Z(n12025) );
  XOR U12323 ( .A(n12025), .B(n12024), .Z(n12078) );
  NOR U12324 ( .A(n99), .B(n48), .Z(n12079) );
  IV U12325 ( .A(n12079), .Z(n12026) );
  NOR U12326 ( .A(n12078), .B(n12026), .Z(n12081) );
  IV U12327 ( .A(n12027), .Z(n12029) );
  XOR U12328 ( .A(n12029), .B(n12028), .Z(n12074) );
  NOR U12329 ( .A(n98), .B(n48), .Z(n12075) );
  IV U12330 ( .A(n12075), .Z(n12030) );
  NOR U12331 ( .A(n12074), .B(n12030), .Z(n12077) );
  IV U12332 ( .A(n12031), .Z(n12033) );
  XOR U12333 ( .A(n12033), .B(n12032), .Z(n12070) );
  NOR U12334 ( .A(n91), .B(n48), .Z(n12071) );
  IV U12335 ( .A(n12071), .Z(n12034) );
  NOR U12336 ( .A(n12070), .B(n12034), .Z(n12073) );
  IV U12337 ( .A(n12035), .Z(n12037) );
  XOR U12338 ( .A(n12037), .B(n12036), .Z(n12066) );
  NOR U12339 ( .A(n97), .B(n48), .Z(n12067) );
  IV U12340 ( .A(n12067), .Z(n12038) );
  NOR U12341 ( .A(n12066), .B(n12038), .Z(n12069) );
  XOR U12342 ( .A(n12040), .B(n12039), .Z(n12062) );
  IV U12343 ( .A(n12062), .Z(n12042) );
  NOR U12344 ( .A(n96), .B(n48), .Z(n12041) );
  IV U12345 ( .A(n12041), .Z(n12063) );
  NOR U12346 ( .A(n12042), .B(n12063), .Z(n12065) );
  NOR U12347 ( .A(n95), .B(n48), .Z(n12059) );
  IV U12348 ( .A(n12059), .Z(n12045) );
  XOR U12349 ( .A(n12044), .B(n12043), .Z(n12058) );
  NOR U12350 ( .A(n12045), .B(n12058), .Z(n12061) );
  NOR U12351 ( .A(n48), .B(n93), .Z(n13017) );
  IV U12352 ( .A(n13017), .Z(n12046) );
  NOR U12353 ( .A(n47), .B(n168), .Z(n12054) );
  IV U12354 ( .A(n12054), .Z(n12049) );
  NOR U12355 ( .A(n12046), .B(n12049), .Z(n12047) );
  IV U12356 ( .A(n12047), .Z(n12048) );
  NOR U12357 ( .A(n94), .B(n12048), .Z(n12057) );
  NOR U12358 ( .A(n12049), .B(n93), .Z(n12050) );
  XOR U12359 ( .A(n94), .B(n12050), .Z(n12051) );
  NOR U12360 ( .A(n48), .B(n12051), .Z(n12052) );
  IV U12361 ( .A(n12052), .Z(n12549) );
  XOR U12362 ( .A(n12054), .B(n12053), .Z(n12548) );
  IV U12363 ( .A(n12548), .Z(n12055) );
  NOR U12364 ( .A(n12549), .B(n12055), .Z(n12056) );
  NOR U12365 ( .A(n12057), .B(n12056), .Z(n12545) );
  XOR U12366 ( .A(n12059), .B(n12058), .Z(n12544) );
  NOR U12367 ( .A(n12545), .B(n12544), .Z(n12060) );
  NOR U12368 ( .A(n12061), .B(n12060), .Z(n12575) );
  XOR U12369 ( .A(n12063), .B(n12062), .Z(n12574) );
  NOR U12370 ( .A(n12575), .B(n12574), .Z(n12064) );
  NOR U12371 ( .A(n12065), .B(n12064), .Z(n12540) );
  XOR U12372 ( .A(n12067), .B(n12066), .Z(n12541) );
  NOR U12373 ( .A(n12540), .B(n12541), .Z(n12068) );
  NOR U12374 ( .A(n12069), .B(n12068), .Z(n12536) );
  XOR U12375 ( .A(n12071), .B(n12070), .Z(n12537) );
  NOR U12376 ( .A(n12536), .B(n12537), .Z(n12072) );
  NOR U12377 ( .A(n12073), .B(n12072), .Z(n12532) );
  XOR U12378 ( .A(n12075), .B(n12074), .Z(n12533) );
  NOR U12379 ( .A(n12532), .B(n12533), .Z(n12076) );
  NOR U12380 ( .A(n12077), .B(n12076), .Z(n12528) );
  XOR U12381 ( .A(n12079), .B(n12078), .Z(n12529) );
  NOR U12382 ( .A(n12528), .B(n12529), .Z(n12080) );
  NOR U12383 ( .A(n12081), .B(n12080), .Z(n12524) );
  XOR U12384 ( .A(n12083), .B(n12082), .Z(n12525) );
  NOR U12385 ( .A(n12524), .B(n12525), .Z(n12084) );
  NOR U12386 ( .A(n12085), .B(n12084), .Z(n12086) );
  IV U12387 ( .A(n12086), .Z(n12522) );
  XOR U12388 ( .A(n12088), .B(n12087), .Z(n12089) );
  IV U12389 ( .A(n12089), .Z(n12521) );
  NOR U12390 ( .A(n12522), .B(n12521), .Z(n12090) );
  NOR U12391 ( .A(n12091), .B(n12090), .Z(n12519) );
  IV U12392 ( .A(n12519), .Z(n12094) );
  XOR U12393 ( .A(n12093), .B(n12092), .Z(n12518) );
  NOR U12394 ( .A(n12094), .B(n12518), .Z(n12095) );
  NOR U12395 ( .A(n12096), .B(n12095), .Z(n12097) );
  IV U12396 ( .A(n12097), .Z(n12516) );
  XOR U12397 ( .A(n12099), .B(n12098), .Z(n12100) );
  IV U12398 ( .A(n12100), .Z(n12515) );
  NOR U12399 ( .A(n12516), .B(n12515), .Z(n12101) );
  NOR U12400 ( .A(n12102), .B(n12101), .Z(n12513) );
  IV U12401 ( .A(n12513), .Z(n12105) );
  XOR U12402 ( .A(n12104), .B(n12103), .Z(n12512) );
  NOR U12403 ( .A(n12105), .B(n12512), .Z(n12106) );
  NOR U12404 ( .A(n12107), .B(n12106), .Z(n12108) );
  IV U12405 ( .A(n12108), .Z(n12510) );
  XOR U12406 ( .A(n12110), .B(n12109), .Z(n12111) );
  IV U12407 ( .A(n12111), .Z(n12509) );
  NOR U12408 ( .A(n12510), .B(n12509), .Z(n12112) );
  NOR U12409 ( .A(n12113), .B(n12112), .Z(n12114) );
  IV U12410 ( .A(n12114), .Z(n12119) );
  NOR U12411 ( .A(n12115), .B(n12119), .Z(n12122) );
  XOR U12412 ( .A(n12117), .B(n12116), .Z(n12118) );
  IV U12413 ( .A(n12118), .Z(n12507) );
  XOR U12414 ( .A(n12120), .B(n12119), .Z(n12508) );
  NOR U12415 ( .A(n12507), .B(n12508), .Z(n12121) );
  NOR U12416 ( .A(n12122), .B(n12121), .Z(n12123) );
  IV U12417 ( .A(n12123), .Z(n12626) );
  XOR U12418 ( .A(n12125), .B(n12124), .Z(n12126) );
  IV U12419 ( .A(n12126), .Z(n12625) );
  NOR U12420 ( .A(n12626), .B(n12625), .Z(n12127) );
  NOR U12421 ( .A(n12128), .B(n12127), .Z(n12505) );
  IV U12422 ( .A(n12505), .Z(n12131) );
  XOR U12423 ( .A(n12130), .B(n12129), .Z(n12504) );
  NOR U12424 ( .A(n12131), .B(n12504), .Z(n12132) );
  NOR U12425 ( .A(n12133), .B(n12132), .Z(n12500) );
  IV U12426 ( .A(n12500), .Z(n12137) );
  IV U12427 ( .A(n12134), .Z(n12136) );
  XOR U12428 ( .A(n12136), .B(n12135), .Z(n12499) );
  NOR U12429 ( .A(n12137), .B(n12499), .Z(n12138) );
  NOR U12430 ( .A(n12139), .B(n12138), .Z(n12496) );
  IV U12431 ( .A(n12496), .Z(n12142) );
  XOR U12432 ( .A(n12141), .B(n12140), .Z(n12495) );
  NOR U12433 ( .A(n12142), .B(n12495), .Z(n12143) );
  NOR U12434 ( .A(n12144), .B(n12143), .Z(n12494) );
  IV U12435 ( .A(n12494), .Z(n12145) );
  NOR U12436 ( .A(n12146), .B(n12145), .Z(n12147) );
  NOR U12437 ( .A(n12148), .B(n12147), .Z(n12149) );
  IV U12438 ( .A(n12149), .Z(n12156) );
  NOR U12439 ( .A(n108), .B(n48), .Z(n12155) );
  IV U12440 ( .A(n12155), .Z(n12150) );
  NOR U12441 ( .A(n12156), .B(n12150), .Z(n12158) );
  XOR U12442 ( .A(n12152), .B(n12151), .Z(n12153) );
  XOR U12443 ( .A(n12154), .B(n12153), .Z(n12489) );
  XOR U12444 ( .A(n12156), .B(n12155), .Z(n12490) );
  NOR U12445 ( .A(n12489), .B(n12490), .Z(n12157) );
  NOR U12446 ( .A(n12158), .B(n12157), .Z(n12483) );
  XOR U12447 ( .A(n12160), .B(n12159), .Z(n12484) );
  NOR U12448 ( .A(n12483), .B(n12484), .Z(n12161) );
  NOR U12449 ( .A(n12162), .B(n12161), .Z(n12479) );
  XOR U12450 ( .A(n12164), .B(n12163), .Z(n12480) );
  NOR U12451 ( .A(n12479), .B(n12480), .Z(n12165) );
  NOR U12452 ( .A(n12166), .B(n12165), .Z(n12477) );
  IV U12453 ( .A(n12477), .Z(n12167) );
  NOR U12454 ( .A(n12168), .B(n12167), .Z(n12169) );
  NOR U12455 ( .A(n12170), .B(n12169), .Z(n12171) );
  IV U12456 ( .A(n12171), .Z(n12177) );
  NOR U12457 ( .A(n12172), .B(n12177), .Z(n12180) );
  XOR U12458 ( .A(n12174), .B(n12173), .Z(n12175) );
  XOR U12459 ( .A(n12176), .B(n12175), .Z(n12471) );
  XOR U12460 ( .A(n12178), .B(n12177), .Z(n12470) );
  NOR U12461 ( .A(n12471), .B(n12470), .Z(n12179) );
  NOR U12462 ( .A(n12180), .B(n12179), .Z(n12671) );
  IV U12463 ( .A(n12671), .Z(n12181) );
  NOR U12464 ( .A(n12182), .B(n12181), .Z(n12183) );
  NOR U12465 ( .A(n12184), .B(n12183), .Z(n12192) );
  IV U12466 ( .A(n12192), .Z(n12186) );
  NOR U12467 ( .A(n112), .B(n48), .Z(n12185) );
  IV U12468 ( .A(n12185), .Z(n12191) );
  NOR U12469 ( .A(n12186), .B(n12191), .Z(n12194) );
  XOR U12470 ( .A(n12188), .B(n12187), .Z(n12189) );
  XOR U12471 ( .A(n12190), .B(n12189), .Z(n12469) );
  XOR U12472 ( .A(n12192), .B(n12191), .Z(n12468) );
  NOR U12473 ( .A(n12469), .B(n12468), .Z(n12193) );
  NOR U12474 ( .A(n12194), .B(n12193), .Z(n12682) );
  IV U12475 ( .A(n12682), .Z(n12195) );
  NOR U12476 ( .A(n12196), .B(n12195), .Z(n12197) );
  NOR U12477 ( .A(n12198), .B(n12197), .Z(n12466) );
  IV U12478 ( .A(n12466), .Z(n12199) );
  NOR U12479 ( .A(n12465), .B(n12199), .Z(n12200) );
  NOR U12480 ( .A(n12201), .B(n12200), .Z(n12463) );
  IV U12481 ( .A(n12463), .Z(n12202) );
  NOR U12482 ( .A(n12203), .B(n12202), .Z(n12204) );
  NOR U12483 ( .A(n12205), .B(n12204), .Z(n12209) );
  IV U12484 ( .A(n12209), .Z(n12206) );
  NOR U12485 ( .A(n12210), .B(n12206), .Z(n12212) );
  XOR U12486 ( .A(n12208), .B(n12207), .Z(n12457) );
  XOR U12487 ( .A(n12210), .B(n12209), .Z(n12456) );
  NOR U12488 ( .A(n12457), .B(n12456), .Z(n12211) );
  NOR U12489 ( .A(n12212), .B(n12211), .Z(n12703) );
  XOR U12490 ( .A(n12214), .B(n12213), .Z(n12704) );
  IV U12491 ( .A(n12704), .Z(n12215) );
  NOR U12492 ( .A(n12703), .B(n12215), .Z(n12216) );
  NOR U12493 ( .A(n12217), .B(n12216), .Z(n12223) );
  XOR U12494 ( .A(n12219), .B(n12218), .Z(n12220) );
  XOR U12495 ( .A(n12221), .B(n12220), .Z(n12222) );
  NOR U12496 ( .A(n12223), .B(n12222), .Z(n12227) );
  XOR U12497 ( .A(n12223), .B(n12222), .Z(n12708) );
  IV U12498 ( .A(n12708), .Z(n12225) );
  NOR U12499 ( .A(n115), .B(n48), .Z(n12224) );
  IV U12500 ( .A(n12224), .Z(n12709) );
  NOR U12501 ( .A(n12225), .B(n12709), .Z(n12226) );
  NOR U12502 ( .A(n12227), .B(n12226), .Z(n12717) );
  NOR U12503 ( .A(n12228), .B(n12717), .Z(n12229) );
  NOR U12504 ( .A(n12230), .B(n12229), .Z(n12237) );
  NOR U12505 ( .A(n116), .B(n48), .Z(n12236) );
  IV U12506 ( .A(n12236), .Z(n12231) );
  NOR U12507 ( .A(n12237), .B(n12231), .Z(n12239) );
  XOR U12508 ( .A(n12233), .B(n12232), .Z(n12234) );
  XOR U12509 ( .A(n12235), .B(n12234), .Z(n12453) );
  XOR U12510 ( .A(n12237), .B(n12236), .Z(n12452) );
  NOR U12511 ( .A(n12453), .B(n12452), .Z(n12238) );
  NOR U12512 ( .A(n12239), .B(n12238), .Z(n12246) );
  XOR U12513 ( .A(n12241), .B(n12240), .Z(n12242) );
  XOR U12514 ( .A(n12243), .B(n12242), .Z(n12245) );
  IV U12515 ( .A(n12245), .Z(n12244) );
  NOR U12516 ( .A(n12246), .B(n12244), .Z(n12249) );
  XOR U12517 ( .A(n12246), .B(n12245), .Z(n12730) );
  NOR U12518 ( .A(n80), .B(n48), .Z(n12731) );
  IV U12519 ( .A(n12731), .Z(n12247) );
  NOR U12520 ( .A(n12730), .B(n12247), .Z(n12248) );
  NOR U12521 ( .A(n12249), .B(n12248), .Z(n12735) );
  XOR U12522 ( .A(n12251), .B(n12250), .Z(n12734) );
  NOR U12523 ( .A(n12735), .B(n12734), .Z(n12252) );
  NOR U12524 ( .A(n12253), .B(n12252), .Z(n12260) );
  NOR U12525 ( .A(n79), .B(n48), .Z(n12259) );
  IV U12526 ( .A(n12259), .Z(n12254) );
  NOR U12527 ( .A(n12260), .B(n12254), .Z(n12262) );
  XOR U12528 ( .A(n12256), .B(n12255), .Z(n12257) );
  XOR U12529 ( .A(n12258), .B(n12257), .Z(n12449) );
  XOR U12530 ( .A(n12260), .B(n12259), .Z(n12448) );
  NOR U12531 ( .A(n12449), .B(n12448), .Z(n12261) );
  NOR U12532 ( .A(n12262), .B(n12261), .Z(n12267) );
  XOR U12533 ( .A(n12264), .B(n12263), .Z(n12266) );
  IV U12534 ( .A(n12266), .Z(n12265) );
  NOR U12535 ( .A(n12267), .B(n12265), .Z(n12270) );
  XOR U12536 ( .A(n12267), .B(n12266), .Z(n12747) );
  NOR U12537 ( .A(n119), .B(n48), .Z(n12268) );
  IV U12538 ( .A(n12268), .Z(n12746) );
  NOR U12539 ( .A(n12747), .B(n12746), .Z(n12269) );
  NOR U12540 ( .A(n12270), .B(n12269), .Z(n12753) );
  XOR U12541 ( .A(n12272), .B(n12271), .Z(n12754) );
  NOR U12542 ( .A(n12753), .B(n12754), .Z(n12273) );
  NOR U12543 ( .A(n12274), .B(n12273), .Z(n12445) );
  XOR U12544 ( .A(n12276), .B(n12275), .Z(n12444) );
  NOR U12545 ( .A(n12445), .B(n12444), .Z(n12277) );
  NOR U12546 ( .A(n12278), .B(n12277), .Z(n12282) );
  XOR U12547 ( .A(n12280), .B(n12279), .Z(n12281) );
  NOR U12548 ( .A(n12282), .B(n12281), .Z(n12286) );
  XOR U12549 ( .A(n12282), .B(n12281), .Z(n12283) );
  IV U12550 ( .A(n12283), .Z(n12770) );
  NOR U12551 ( .A(n125), .B(n48), .Z(n12771) );
  IV U12552 ( .A(n12771), .Z(n12284) );
  NOR U12553 ( .A(n12770), .B(n12284), .Z(n12285) );
  NOR U12554 ( .A(n12286), .B(n12285), .Z(n12775) );
  XOR U12555 ( .A(n12288), .B(n12287), .Z(n12774) );
  NOR U12556 ( .A(n12775), .B(n12774), .Z(n12289) );
  NOR U12557 ( .A(n12290), .B(n12289), .Z(n12295) );
  NOR U12558 ( .A(n128), .B(n48), .Z(n12294) );
  IV U12559 ( .A(n12294), .Z(n12291) );
  NOR U12560 ( .A(n12295), .B(n12291), .Z(n12298) );
  XOR U12561 ( .A(n12293), .B(n12292), .Z(n12442) );
  IV U12562 ( .A(n12442), .Z(n12296) );
  XOR U12563 ( .A(n12295), .B(n12294), .Z(n12441) );
  NOR U12564 ( .A(n12296), .B(n12441), .Z(n12297) );
  NOR U12565 ( .A(n12298), .B(n12297), .Z(n12303) );
  XOR U12566 ( .A(n12300), .B(n12299), .Z(n12302) );
  IV U12567 ( .A(n12302), .Z(n12301) );
  NOR U12568 ( .A(n12303), .B(n12301), .Z(n12306) );
  XOR U12569 ( .A(n12303), .B(n12302), .Z(n12787) );
  NOR U12570 ( .A(n131), .B(n48), .Z(n12788) );
  IV U12571 ( .A(n12788), .Z(n12304) );
  NOR U12572 ( .A(n12787), .B(n12304), .Z(n12305) );
  NOR U12573 ( .A(n12306), .B(n12305), .Z(n12794) );
  XOR U12574 ( .A(n12308), .B(n12307), .Z(n12793) );
  NOR U12575 ( .A(n12794), .B(n12793), .Z(n12309) );
  NOR U12576 ( .A(n12310), .B(n12309), .Z(n12313) );
  NOR U12577 ( .A(n135), .B(n48), .Z(n12312) );
  IV U12578 ( .A(n12312), .Z(n12311) );
  NOR U12579 ( .A(n12313), .B(n12311), .Z(n12317) );
  XOR U12580 ( .A(n12313), .B(n12312), .Z(n12438) );
  XOR U12581 ( .A(n12315), .B(n12314), .Z(n12437) );
  NOR U12582 ( .A(n12438), .B(n12437), .Z(n12316) );
  NOR U12583 ( .A(n12317), .B(n12316), .Z(n12321) );
  XOR U12584 ( .A(n12319), .B(n12318), .Z(n12320) );
  NOR U12585 ( .A(n12321), .B(n12320), .Z(n12325) );
  XOR U12586 ( .A(n12321), .B(n12320), .Z(n12808) );
  IV U12587 ( .A(n12808), .Z(n12323) );
  NOR U12588 ( .A(n137), .B(n48), .Z(n12322) );
  IV U12589 ( .A(n12322), .Z(n12809) );
  NOR U12590 ( .A(n12323), .B(n12809), .Z(n12324) );
  NOR U12591 ( .A(n12325), .B(n12324), .Z(n12813) );
  XOR U12592 ( .A(n12327), .B(n12326), .Z(n12812) );
  NOR U12593 ( .A(n12813), .B(n12812), .Z(n12328) );
  NOR U12594 ( .A(n12329), .B(n12328), .Z(n12436) );
  XOR U12595 ( .A(n12331), .B(n12330), .Z(n12435) );
  NOR U12596 ( .A(n12436), .B(n12435), .Z(n12332) );
  NOR U12597 ( .A(n12333), .B(n12332), .Z(n12337) );
  XOR U12598 ( .A(n12335), .B(n12334), .Z(n12336) );
  NOR U12599 ( .A(n12337), .B(n12336), .Z(n12341) );
  XOR U12600 ( .A(n12337), .B(n12336), .Z(n12338) );
  IV U12601 ( .A(n12338), .Z(n12829) );
  NOR U12602 ( .A(n143), .B(n48), .Z(n12830) );
  IV U12603 ( .A(n12830), .Z(n12339) );
  NOR U12604 ( .A(n12829), .B(n12339), .Z(n12340) );
  NOR U12605 ( .A(n12341), .B(n12340), .Z(n12834) );
  XOR U12606 ( .A(n12343), .B(n12342), .Z(n12833) );
  NOR U12607 ( .A(n12834), .B(n12833), .Z(n12344) );
  NOR U12608 ( .A(n12345), .B(n12344), .Z(n12431) );
  XOR U12609 ( .A(n12347), .B(n12346), .Z(n12432) );
  NOR U12610 ( .A(n12431), .B(n12432), .Z(n12348) );
  NOR U12611 ( .A(n12349), .B(n12348), .Z(n12353) );
  XOR U12612 ( .A(n12351), .B(n12350), .Z(n12352) );
  NOR U12613 ( .A(n12353), .B(n12352), .Z(n12357) );
  XOR U12614 ( .A(n12353), .B(n12352), .Z(n12848) );
  IV U12615 ( .A(n12848), .Z(n12355) );
  NOR U12616 ( .A(n148), .B(n48), .Z(n12354) );
  IV U12617 ( .A(n12354), .Z(n12849) );
  NOR U12618 ( .A(n12355), .B(n12849), .Z(n12356) );
  NOR U12619 ( .A(n12357), .B(n12356), .Z(n12853) );
  XOR U12620 ( .A(n12359), .B(n12358), .Z(n12852) );
  NOR U12621 ( .A(n12853), .B(n12852), .Z(n12360) );
  NOR U12622 ( .A(n12361), .B(n12360), .Z(n12364) );
  NOR U12623 ( .A(n153), .B(n48), .Z(n12363) );
  IV U12624 ( .A(n12363), .Z(n12362) );
  NOR U12625 ( .A(n12364), .B(n12362), .Z(n12369) );
  XOR U12626 ( .A(n12364), .B(n12363), .Z(n12428) );
  XOR U12627 ( .A(n12366), .B(n12365), .Z(n12429) );
  IV U12628 ( .A(n12429), .Z(n12367) );
  NOR U12629 ( .A(n12428), .B(n12367), .Z(n12368) );
  NOR U12630 ( .A(n12369), .B(n12368), .Z(n12374) );
  XOR U12631 ( .A(n12371), .B(n12370), .Z(n12373) );
  IV U12632 ( .A(n12373), .Z(n12372) );
  NOR U12633 ( .A(n12374), .B(n12372), .Z(n12377) );
  XOR U12634 ( .A(n12374), .B(n12373), .Z(n12867) );
  NOR U12635 ( .A(n155), .B(n48), .Z(n12868) );
  IV U12636 ( .A(n12868), .Z(n12375) );
  NOR U12637 ( .A(n12867), .B(n12375), .Z(n12376) );
  NOR U12638 ( .A(n12377), .B(n12376), .Z(n12872) );
  XOR U12639 ( .A(n12379), .B(n12378), .Z(n12871) );
  NOR U12640 ( .A(n12872), .B(n12871), .Z(n12380) );
  NOR U12641 ( .A(n12381), .B(n12380), .Z(n12384) );
  NOR U12642 ( .A(n158), .B(n48), .Z(n12383) );
  IV U12643 ( .A(n12383), .Z(n12382) );
  NOR U12644 ( .A(n12384), .B(n12382), .Z(n12388) );
  XOR U12645 ( .A(n12384), .B(n12383), .Z(n12425) );
  XOR U12646 ( .A(n12386), .B(n12385), .Z(n12424) );
  NOR U12647 ( .A(n12425), .B(n12424), .Z(n12387) );
  NOR U12648 ( .A(n12388), .B(n12387), .Z(n12392) );
  XOR U12649 ( .A(n12390), .B(n12389), .Z(n12391) );
  NOR U12650 ( .A(n12392), .B(n12391), .Z(n12396) );
  XOR U12651 ( .A(n12392), .B(n12391), .Z(n12886) );
  IV U12652 ( .A(n12886), .Z(n12394) );
  NOR U12653 ( .A(n161), .B(n48), .Z(n12393) );
  IV U12654 ( .A(n12393), .Z(n12887) );
  NOR U12655 ( .A(n12394), .B(n12887), .Z(n12395) );
  NOR U12656 ( .A(n12396), .B(n12395), .Z(n12891) );
  XOR U12657 ( .A(n12398), .B(n12397), .Z(n12890) );
  NOR U12658 ( .A(n12891), .B(n12890), .Z(n12399) );
  NOR U12659 ( .A(n12400), .B(n12399), .Z(n12405) );
  XOR U12660 ( .A(n12402), .B(n12401), .Z(n12404) );
  IV U12661 ( .A(n12404), .Z(n12403) );
  NOR U12662 ( .A(n12405), .B(n12403), .Z(n12408) );
  XOR U12663 ( .A(n12405), .B(n12404), .Z(n12421) );
  NOR U12664 ( .A(n165), .B(n48), .Z(n12422) );
  IV U12665 ( .A(n12422), .Z(n12406) );
  NOR U12666 ( .A(n12421), .B(n12406), .Z(n12407) );
  NOR U12667 ( .A(n12408), .B(n12407), .Z(n12412) );
  XOR U12668 ( .A(n12410), .B(n12409), .Z(n12411) );
  NOR U12669 ( .A(n12412), .B(n12411), .Z(n12416) );
  XOR U12670 ( .A(n12412), .B(n12411), .Z(n12902) );
  IV U12671 ( .A(n12902), .Z(n12414) );
  NOR U12672 ( .A(n167), .B(n48), .Z(n12413) );
  IV U12673 ( .A(n12413), .Z(n12903) );
  NOR U12674 ( .A(n12414), .B(n12903), .Z(n12415) );
  NOR U12675 ( .A(n12416), .B(n12415), .Z(n12905) );
  XOR U12676 ( .A(n12418), .B(n12417), .Z(n12904) );
  NOR U12677 ( .A(n12905), .B(n12904), .Z(n28624) );
  XOR U12678 ( .A(n12420), .B(n12419), .Z(n28623) );
  NOR U12679 ( .A(n28624), .B(n28623), .Z(n28627) );
  XOR U12680 ( .A(n12422), .B(n12421), .Z(n12898) );
  NOR U12681 ( .A(n167), .B(n49), .Z(n12899) );
  IV U12682 ( .A(n12899), .Z(n12423) );
  NOR U12683 ( .A(n12898), .B(n12423), .Z(n12901) );
  IV U12684 ( .A(n12424), .Z(n12426) );
  XOR U12685 ( .A(n12426), .B(n12425), .Z(n12879) );
  NOR U12686 ( .A(n161), .B(n49), .Z(n12880) );
  IV U12687 ( .A(n12880), .Z(n12427) );
  NOR U12688 ( .A(n12879), .B(n12427), .Z(n12882) );
  XOR U12689 ( .A(n12429), .B(n12428), .Z(n12860) );
  NOR U12690 ( .A(n155), .B(n49), .Z(n12861) );
  IV U12691 ( .A(n12861), .Z(n12430) );
  NOR U12692 ( .A(n12860), .B(n12430), .Z(n12863) );
  IV U12693 ( .A(n12431), .Z(n12433) );
  XOR U12694 ( .A(n12433), .B(n12432), .Z(n12841) );
  NOR U12695 ( .A(n148), .B(n49), .Z(n12842) );
  IV U12696 ( .A(n12842), .Z(n12434) );
  NOR U12697 ( .A(n12841), .B(n12434), .Z(n12844) );
  XOR U12698 ( .A(n12436), .B(n12435), .Z(n12822) );
  IV U12699 ( .A(n12437), .Z(n12439) );
  XOR U12700 ( .A(n12439), .B(n12438), .Z(n12801) );
  NOR U12701 ( .A(n137), .B(n49), .Z(n12802) );
  IV U12702 ( .A(n12802), .Z(n12440) );
  NOR U12703 ( .A(n12801), .B(n12440), .Z(n12804) );
  XOR U12704 ( .A(n12442), .B(n12441), .Z(n12782) );
  NOR U12705 ( .A(n131), .B(n49), .Z(n12783) );
  IV U12706 ( .A(n12783), .Z(n12443) );
  NOR U12707 ( .A(n12782), .B(n12443), .Z(n12785) );
  NOR U12708 ( .A(n125), .B(n49), .Z(n12446) );
  XOR U12709 ( .A(n12445), .B(n12444), .Z(n12447) );
  NOR U12710 ( .A(n12446), .B(n12447), .Z(n12765) );
  IV U12711 ( .A(n12446), .Z(n13246) );
  IV U12712 ( .A(n12447), .Z(n13245) );
  NOR U12713 ( .A(n13246), .B(n13245), .Z(n12763) );
  NOR U12714 ( .A(n120), .B(n49), .Z(n12748) );
  NOR U12715 ( .A(n119), .B(n49), .Z(n12450) );
  XOR U12716 ( .A(n12449), .B(n12448), .Z(n12451) );
  NOR U12717 ( .A(n12450), .B(n12451), .Z(n12745) );
  IV U12718 ( .A(n12450), .Z(n13222) );
  IV U12719 ( .A(n12451), .Z(n13221) );
  NOR U12720 ( .A(n13222), .B(n13221), .Z(n12743) );
  XOR U12721 ( .A(n12453), .B(n12452), .Z(n12455) );
  IV U12722 ( .A(n12455), .Z(n13198) );
  NOR U12723 ( .A(n80), .B(n49), .Z(n13196) );
  IV U12724 ( .A(n13196), .Z(n12454) );
  NOR U12725 ( .A(n13198), .B(n12454), .Z(n12726) );
  NOR U12726 ( .A(n12455), .B(n13196), .Z(n12724) );
  XOR U12727 ( .A(n12457), .B(n12456), .Z(n12458) );
  IV U12728 ( .A(n12458), .Z(n12696) );
  NOR U12729 ( .A(n82), .B(n49), .Z(n12697) );
  IV U12730 ( .A(n12697), .Z(n12459) );
  NOR U12731 ( .A(n12696), .B(n12459), .Z(n12699) );
  XOR U12732 ( .A(n12461), .B(n12460), .Z(n12462) );
  XOR U12733 ( .A(n12463), .B(n12462), .Z(n12693) );
  NOR U12734 ( .A(n114), .B(n49), .Z(n12692) );
  IV U12735 ( .A(n12692), .Z(n12464) );
  NOR U12736 ( .A(n12693), .B(n12464), .Z(n12695) );
  NOR U12737 ( .A(n83), .B(n49), .Z(n12689) );
  IV U12738 ( .A(n12689), .Z(n12467) );
  XOR U12739 ( .A(n12466), .B(n12465), .Z(n12688) );
  NOR U12740 ( .A(n12467), .B(n12688), .Z(n12691) );
  XOR U12741 ( .A(n12469), .B(n12468), .Z(n12677) );
  IV U12742 ( .A(n12677), .Z(n12926) );
  NOR U12743 ( .A(n84), .B(n49), .Z(n12676) );
  IV U12744 ( .A(n12676), .Z(n12925) );
  NOR U12745 ( .A(n12926), .B(n12925), .Z(n12680) );
  XOR U12746 ( .A(n12471), .B(n12470), .Z(n12939) );
  IV U12747 ( .A(n12939), .Z(n12473) );
  NOR U12748 ( .A(n85), .B(n49), .Z(n12937) );
  IV U12749 ( .A(n12937), .Z(n12472) );
  NOR U12750 ( .A(n12473), .B(n12472), .Z(n12666) );
  XOR U12751 ( .A(n12475), .B(n12474), .Z(n12476) );
  XOR U12752 ( .A(n12477), .B(n12476), .Z(n12661) );
  NOR U12753 ( .A(n111), .B(n49), .Z(n12660) );
  IV U12754 ( .A(n12660), .Z(n12478) );
  NOR U12755 ( .A(n12661), .B(n12478), .Z(n12663) );
  XOR U12756 ( .A(n12480), .B(n12479), .Z(n12481) );
  IV U12757 ( .A(n12481), .Z(n12656) );
  NOR U12758 ( .A(n86), .B(n49), .Z(n12657) );
  IV U12759 ( .A(n12657), .Z(n12482) );
  NOR U12760 ( .A(n12656), .B(n12482), .Z(n12659) );
  XOR U12761 ( .A(n12484), .B(n12483), .Z(n12485) );
  IV U12762 ( .A(n12485), .Z(n12487) );
  NOR U12763 ( .A(n110), .B(n49), .Z(n12488) );
  IV U12764 ( .A(n12488), .Z(n12486) );
  NOR U12765 ( .A(n12487), .B(n12486), .Z(n12655) );
  XOR U12766 ( .A(n12488), .B(n12487), .Z(n12943) );
  XOR U12767 ( .A(n12490), .B(n12489), .Z(n12648) );
  NOR U12768 ( .A(n109), .B(n49), .Z(n12649) );
  NOR U12769 ( .A(n12648), .B(n12649), .Z(n12652) );
  XOR U12770 ( .A(n12492), .B(n12491), .Z(n12493) );
  XOR U12771 ( .A(n12494), .B(n12493), .Z(n12643) );
  XOR U12772 ( .A(n12496), .B(n12495), .Z(n12953) );
  IV U12773 ( .A(n12953), .Z(n12497) );
  NOR U12774 ( .A(n87), .B(n49), .Z(n12951) );
  NOR U12775 ( .A(n12497), .B(n12951), .Z(n12640) );
  IV U12776 ( .A(n12951), .Z(n12498) );
  NOR U12777 ( .A(n12953), .B(n12498), .Z(n12638) );
  NOR U12778 ( .A(n107), .B(n49), .Z(n12502) );
  XOR U12779 ( .A(n12500), .B(n12499), .Z(n12501) );
  NOR U12780 ( .A(n12502), .B(n12501), .Z(n12637) );
  IV U12781 ( .A(n12501), .Z(n12503) );
  XOR U12782 ( .A(n12503), .B(n12502), .Z(n12957) );
  NOR U12783 ( .A(n88), .B(n49), .Z(n12632) );
  IV U12784 ( .A(n12632), .Z(n12506) );
  XOR U12785 ( .A(n12505), .B(n12504), .Z(n12631) );
  NOR U12786 ( .A(n12506), .B(n12631), .Z(n12634) );
  XOR U12787 ( .A(n12508), .B(n12507), .Z(n12620) );
  IV U12788 ( .A(n12620), .Z(n13088) );
  NOR U12789 ( .A(n105), .B(n49), .Z(n12619) );
  IV U12790 ( .A(n12619), .Z(n13087) );
  NOR U12791 ( .A(n13088), .B(n13087), .Z(n12623) );
  XOR U12792 ( .A(n12510), .B(n12509), .Z(n12616) );
  NOR U12793 ( .A(n104), .B(n49), .Z(n12615) );
  IV U12794 ( .A(n12615), .Z(n12511) );
  NOR U12795 ( .A(n12616), .B(n12511), .Z(n12618) );
  XOR U12796 ( .A(n12513), .B(n12512), .Z(n12611) );
  NOR U12797 ( .A(n89), .B(n49), .Z(n12612) );
  IV U12798 ( .A(n12612), .Z(n12514) );
  NOR U12799 ( .A(n12611), .B(n12514), .Z(n12614) );
  XOR U12800 ( .A(n12516), .B(n12515), .Z(n12608) );
  NOR U12801 ( .A(n103), .B(n49), .Z(n12607) );
  IV U12802 ( .A(n12607), .Z(n12517) );
  NOR U12803 ( .A(n12608), .B(n12517), .Z(n12610) );
  XOR U12804 ( .A(n12519), .B(n12518), .Z(n12603) );
  NOR U12805 ( .A(n90), .B(n49), .Z(n12604) );
  IV U12806 ( .A(n12604), .Z(n12520) );
  NOR U12807 ( .A(n12603), .B(n12520), .Z(n12606) );
  XOR U12808 ( .A(n12522), .B(n12521), .Z(n12600) );
  NOR U12809 ( .A(n102), .B(n49), .Z(n12599) );
  IV U12810 ( .A(n12599), .Z(n12523) );
  NOR U12811 ( .A(n12600), .B(n12523), .Z(n12602) );
  IV U12812 ( .A(n12524), .Z(n12526) );
  XOR U12813 ( .A(n12526), .B(n12525), .Z(n12595) );
  NOR U12814 ( .A(n101), .B(n49), .Z(n12596) );
  IV U12815 ( .A(n12596), .Z(n12527) );
  NOR U12816 ( .A(n12595), .B(n12527), .Z(n12598) );
  IV U12817 ( .A(n12528), .Z(n12530) );
  XOR U12818 ( .A(n12530), .B(n12529), .Z(n12591) );
  NOR U12819 ( .A(n100), .B(n49), .Z(n12592) );
  IV U12820 ( .A(n12592), .Z(n12531) );
  NOR U12821 ( .A(n12591), .B(n12531), .Z(n12594) );
  IV U12822 ( .A(n12532), .Z(n12534) );
  XOR U12823 ( .A(n12534), .B(n12533), .Z(n12587) );
  NOR U12824 ( .A(n99), .B(n49), .Z(n12588) );
  IV U12825 ( .A(n12588), .Z(n12535) );
  NOR U12826 ( .A(n12587), .B(n12535), .Z(n12590) );
  IV U12827 ( .A(n12536), .Z(n12538) );
  XOR U12828 ( .A(n12538), .B(n12537), .Z(n12583) );
  NOR U12829 ( .A(n98), .B(n49), .Z(n12584) );
  IV U12830 ( .A(n12584), .Z(n12539) );
  NOR U12831 ( .A(n12583), .B(n12539), .Z(n12586) );
  IV U12832 ( .A(n12540), .Z(n12542) );
  XOR U12833 ( .A(n12542), .B(n12541), .Z(n12579) );
  NOR U12834 ( .A(n91), .B(n49), .Z(n12580) );
  IV U12835 ( .A(n12580), .Z(n12543) );
  NOR U12836 ( .A(n12579), .B(n12543), .Z(n12582) );
  XOR U12837 ( .A(n12545), .B(n12544), .Z(n12567) );
  IV U12838 ( .A(n12567), .Z(n12547) );
  NOR U12839 ( .A(n96), .B(n49), .Z(n12546) );
  IV U12840 ( .A(n12546), .Z(n12568) );
  NOR U12841 ( .A(n12547), .B(n12568), .Z(n12570) );
  NOR U12842 ( .A(n95), .B(n49), .Z(n12564) );
  IV U12843 ( .A(n12564), .Z(n12550) );
  XOR U12844 ( .A(n12549), .B(n12548), .Z(n12563) );
  NOR U12845 ( .A(n12550), .B(n12563), .Z(n12566) );
  NOR U12846 ( .A(n49), .B(n93), .Z(n13532) );
  IV U12847 ( .A(n13532), .Z(n12551) );
  NOR U12848 ( .A(n48), .B(n168), .Z(n12559) );
  IV U12849 ( .A(n12559), .Z(n12554) );
  NOR U12850 ( .A(n12551), .B(n12554), .Z(n12552) );
  IV U12851 ( .A(n12552), .Z(n12553) );
  NOR U12852 ( .A(n94), .B(n12553), .Z(n12562) );
  NOR U12853 ( .A(n12554), .B(n93), .Z(n12555) );
  XOR U12854 ( .A(n94), .B(n12555), .Z(n12556) );
  NOR U12855 ( .A(n49), .B(n12556), .Z(n12557) );
  IV U12856 ( .A(n12557), .Z(n13008) );
  XOR U12857 ( .A(n12559), .B(n12558), .Z(n13007) );
  IV U12858 ( .A(n13007), .Z(n12560) );
  NOR U12859 ( .A(n13008), .B(n12560), .Z(n12561) );
  NOR U12860 ( .A(n12562), .B(n12561), .Z(n13004) );
  XOR U12861 ( .A(n12564), .B(n12563), .Z(n13003) );
  NOR U12862 ( .A(n13004), .B(n13003), .Z(n12565) );
  NOR U12863 ( .A(n12566), .B(n12565), .Z(n13031) );
  XOR U12864 ( .A(n12568), .B(n12567), .Z(n13030) );
  NOR U12865 ( .A(n13031), .B(n13030), .Z(n12569) );
  NOR U12866 ( .A(n12570), .B(n12569), .Z(n12573) );
  NOR U12867 ( .A(n97), .B(n49), .Z(n12572) );
  IV U12868 ( .A(n12572), .Z(n12571) );
  NOR U12869 ( .A(n12573), .B(n12571), .Z(n12578) );
  XOR U12870 ( .A(n12573), .B(n12572), .Z(n13000) );
  XOR U12871 ( .A(n12575), .B(n12574), .Z(n13001) );
  IV U12872 ( .A(n13001), .Z(n12576) );
  NOR U12873 ( .A(n13000), .B(n12576), .Z(n12577) );
  NOR U12874 ( .A(n12578), .B(n12577), .Z(n12996) );
  XOR U12875 ( .A(n12580), .B(n12579), .Z(n12997) );
  NOR U12876 ( .A(n12996), .B(n12997), .Z(n12581) );
  NOR U12877 ( .A(n12582), .B(n12581), .Z(n12992) );
  XOR U12878 ( .A(n12584), .B(n12583), .Z(n12993) );
  NOR U12879 ( .A(n12992), .B(n12993), .Z(n12585) );
  NOR U12880 ( .A(n12586), .B(n12585), .Z(n12988) );
  XOR U12881 ( .A(n12588), .B(n12587), .Z(n12989) );
  NOR U12882 ( .A(n12988), .B(n12989), .Z(n12589) );
  NOR U12883 ( .A(n12590), .B(n12589), .Z(n12984) );
  XOR U12884 ( .A(n12592), .B(n12591), .Z(n12985) );
  NOR U12885 ( .A(n12984), .B(n12985), .Z(n12593) );
  NOR U12886 ( .A(n12594), .B(n12593), .Z(n12980) );
  XOR U12887 ( .A(n12596), .B(n12595), .Z(n12981) );
  NOR U12888 ( .A(n12980), .B(n12981), .Z(n12597) );
  NOR U12889 ( .A(n12598), .B(n12597), .Z(n12979) );
  XOR U12890 ( .A(n12600), .B(n12599), .Z(n12978) );
  NOR U12891 ( .A(n12979), .B(n12978), .Z(n12601) );
  NOR U12892 ( .A(n12602), .B(n12601), .Z(n12974) );
  XOR U12893 ( .A(n12604), .B(n12603), .Z(n12975) );
  NOR U12894 ( .A(n12974), .B(n12975), .Z(n12605) );
  NOR U12895 ( .A(n12606), .B(n12605), .Z(n12970) );
  XOR U12896 ( .A(n12608), .B(n12607), .Z(n12971) );
  NOR U12897 ( .A(n12970), .B(n12971), .Z(n12609) );
  NOR U12898 ( .A(n12610), .B(n12609), .Z(n12966) );
  XOR U12899 ( .A(n12612), .B(n12611), .Z(n12967) );
  NOR U12900 ( .A(n12966), .B(n12967), .Z(n12613) );
  NOR U12901 ( .A(n12614), .B(n12613), .Z(n12964) );
  XOR U12902 ( .A(n12616), .B(n12615), .Z(n12965) );
  NOR U12903 ( .A(n12964), .B(n12965), .Z(n12617) );
  NOR U12904 ( .A(n12618), .B(n12617), .Z(n13090) );
  NOR U12905 ( .A(n12620), .B(n12619), .Z(n12621) );
  NOR U12906 ( .A(n13090), .B(n12621), .Z(n12622) );
  NOR U12907 ( .A(n12623), .B(n12622), .Z(n12628) );
  NOR U12908 ( .A(n106), .B(n49), .Z(n12627) );
  IV U12909 ( .A(n12627), .Z(n12624) );
  NOR U12910 ( .A(n12628), .B(n12624), .Z(n12630) );
  XOR U12911 ( .A(n12626), .B(n12625), .Z(n12961) );
  XOR U12912 ( .A(n12628), .B(n12627), .Z(n12960) );
  NOR U12913 ( .A(n12961), .B(n12960), .Z(n12629) );
  NOR U12914 ( .A(n12630), .B(n12629), .Z(n13101) );
  XOR U12915 ( .A(n12632), .B(n12631), .Z(n13102) );
  NOR U12916 ( .A(n13101), .B(n13102), .Z(n12633) );
  NOR U12917 ( .A(n12634), .B(n12633), .Z(n12635) );
  IV U12918 ( .A(n12635), .Z(n12958) );
  NOR U12919 ( .A(n12957), .B(n12958), .Z(n12636) );
  NOR U12920 ( .A(n12637), .B(n12636), .Z(n12950) );
  NOR U12921 ( .A(n12638), .B(n12950), .Z(n12639) );
  NOR U12922 ( .A(n12640), .B(n12639), .Z(n12642) );
  IV U12923 ( .A(n12642), .Z(n12641) );
  NOR U12924 ( .A(n12643), .B(n12641), .Z(n12646) );
  XOR U12925 ( .A(n12643), .B(n12642), .Z(n12948) );
  NOR U12926 ( .A(n108), .B(n49), .Z(n12644) );
  IV U12927 ( .A(n12644), .Z(n12949) );
  NOR U12928 ( .A(n12948), .B(n12949), .Z(n12645) );
  NOR U12929 ( .A(n12646), .B(n12645), .Z(n12647) );
  IV U12930 ( .A(n12647), .Z(n12947) );
  XOR U12931 ( .A(n12649), .B(n12648), .Z(n12650) );
  IV U12932 ( .A(n12650), .Z(n12946) );
  NOR U12933 ( .A(n12947), .B(n12946), .Z(n12651) );
  NOR U12934 ( .A(n12652), .B(n12651), .Z(n12944) );
  IV U12935 ( .A(n12944), .Z(n12653) );
  NOR U12936 ( .A(n12943), .B(n12653), .Z(n12654) );
  NOR U12937 ( .A(n12655), .B(n12654), .Z(n13132) );
  XOR U12938 ( .A(n12657), .B(n12656), .Z(n13133) );
  NOR U12939 ( .A(n13132), .B(n13133), .Z(n12658) );
  NOR U12940 ( .A(n12659), .B(n12658), .Z(n12942) );
  XOR U12941 ( .A(n12661), .B(n12660), .Z(n12941) );
  NOR U12942 ( .A(n12942), .B(n12941), .Z(n12662) );
  NOR U12943 ( .A(n12663), .B(n12662), .Z(n12936) );
  NOR U12944 ( .A(n12939), .B(n12937), .Z(n12664) );
  NOR U12945 ( .A(n12936), .B(n12664), .Z(n12665) );
  NOR U12946 ( .A(n12666), .B(n12665), .Z(n12672) );
  NOR U12947 ( .A(n112), .B(n49), .Z(n12673) );
  IV U12948 ( .A(n12673), .Z(n12667) );
  NOR U12949 ( .A(n12672), .B(n12667), .Z(n12675) );
  XOR U12950 ( .A(n12669), .B(n12668), .Z(n12670) );
  XOR U12951 ( .A(n12671), .B(n12670), .Z(n12931) );
  XOR U12952 ( .A(n12673), .B(n12672), .Z(n12930) );
  NOR U12953 ( .A(n12931), .B(n12930), .Z(n12674) );
  NOR U12954 ( .A(n12675), .B(n12674), .Z(n12928) );
  NOR U12955 ( .A(n12677), .B(n12676), .Z(n12678) );
  NOR U12956 ( .A(n12928), .B(n12678), .Z(n12679) );
  NOR U12957 ( .A(n12680), .B(n12679), .Z(n12684) );
  NOR U12958 ( .A(n113), .B(n49), .Z(n12685) );
  IV U12959 ( .A(n12685), .Z(n12681) );
  NOR U12960 ( .A(n12684), .B(n12681), .Z(n12687) );
  XOR U12961 ( .A(n12683), .B(n12682), .Z(n12922) );
  XOR U12962 ( .A(n12685), .B(n12684), .Z(n12921) );
  NOR U12963 ( .A(n12922), .B(n12921), .Z(n12686) );
  NOR U12964 ( .A(n12687), .B(n12686), .Z(n12917) );
  XOR U12965 ( .A(n12689), .B(n12688), .Z(n12918) );
  NOR U12966 ( .A(n12917), .B(n12918), .Z(n12690) );
  NOR U12967 ( .A(n12691), .B(n12690), .Z(n12913) );
  XOR U12968 ( .A(n12693), .B(n12692), .Z(n12914) );
  NOR U12969 ( .A(n12913), .B(n12914), .Z(n12694) );
  NOR U12970 ( .A(n12695), .B(n12694), .Z(n12909) );
  XOR U12971 ( .A(n12697), .B(n12696), .Z(n12910) );
  NOR U12972 ( .A(n12909), .B(n12910), .Z(n12698) );
  NOR U12973 ( .A(n12699), .B(n12698), .Z(n12702) );
  NOR U12974 ( .A(n115), .B(n49), .Z(n12701) );
  IV U12975 ( .A(n12701), .Z(n12700) );
  NOR U12976 ( .A(n12702), .B(n12700), .Z(n12706) );
  XOR U12977 ( .A(n12702), .B(n12701), .Z(n13174) );
  XOR U12978 ( .A(n12704), .B(n12703), .Z(n13173) );
  NOR U12979 ( .A(n13174), .B(n13173), .Z(n12705) );
  NOR U12980 ( .A(n12706), .B(n12705), .Z(n12711) );
  NOR U12981 ( .A(n81), .B(n49), .Z(n12710) );
  IV U12982 ( .A(n12710), .Z(n12707) );
  NOR U12983 ( .A(n12711), .B(n12707), .Z(n12713) );
  XOR U12984 ( .A(n12709), .B(n12708), .Z(n13179) );
  XOR U12985 ( .A(n12711), .B(n12710), .Z(n13180) );
  NOR U12986 ( .A(n13179), .B(n13180), .Z(n12712) );
  NOR U12987 ( .A(n12713), .B(n12712), .Z(n12719) );
  XOR U12988 ( .A(n12715), .B(n12714), .Z(n12716) );
  XOR U12989 ( .A(n12717), .B(n12716), .Z(n12718) );
  NOR U12990 ( .A(n12719), .B(n12718), .Z(n12723) );
  XOR U12991 ( .A(n12719), .B(n12718), .Z(n12720) );
  IV U12992 ( .A(n12720), .Z(n13191) );
  NOR U12993 ( .A(n116), .B(n49), .Z(n12721) );
  IV U12994 ( .A(n12721), .Z(n13190) );
  NOR U12995 ( .A(n13191), .B(n13190), .Z(n12722) );
  NOR U12996 ( .A(n12723), .B(n12722), .Z(n13195) );
  NOR U12997 ( .A(n12724), .B(n13195), .Z(n12725) );
  NOR U12998 ( .A(n12726), .B(n12725), .Z(n12729) );
  NOR U12999 ( .A(n117), .B(n49), .Z(n12728) );
  IV U13000 ( .A(n12728), .Z(n12727) );
  NOR U13001 ( .A(n12729), .B(n12727), .Z(n12733) );
  XOR U13002 ( .A(n12729), .B(n12728), .Z(n13204) );
  XOR U13003 ( .A(n12731), .B(n12730), .Z(n13205) );
  NOR U13004 ( .A(n13204), .B(n13205), .Z(n12732) );
  NOR U13005 ( .A(n12733), .B(n12732), .Z(n12738) );
  XOR U13006 ( .A(n12735), .B(n12734), .Z(n12737) );
  IV U13007 ( .A(n12737), .Z(n12736) );
  NOR U13008 ( .A(n12738), .B(n12736), .Z(n12741) );
  XOR U13009 ( .A(n12738), .B(n12737), .Z(n13215) );
  NOR U13010 ( .A(n79), .B(n49), .Z(n12739) );
  IV U13011 ( .A(n12739), .Z(n13214) );
  NOR U13012 ( .A(n13215), .B(n13214), .Z(n12740) );
  NOR U13013 ( .A(n12741), .B(n12740), .Z(n13224) );
  IV U13014 ( .A(n13224), .Z(n12742) );
  NOR U13015 ( .A(n12743), .B(n12742), .Z(n12744) );
  NOR U13016 ( .A(n12745), .B(n12744), .Z(n12749) );
  NOR U13017 ( .A(n12748), .B(n12749), .Z(n12752) );
  XOR U13018 ( .A(n12747), .B(n12746), .Z(n13229) );
  IV U13019 ( .A(n12748), .Z(n12750) );
  XOR U13020 ( .A(n12750), .B(n12749), .Z(n13230) );
  NOR U13021 ( .A(n13229), .B(n13230), .Z(n12751) );
  NOR U13022 ( .A(n12752), .B(n12751), .Z(n12758) );
  IV U13023 ( .A(n12758), .Z(n12756) );
  IV U13024 ( .A(n12753), .Z(n12755) );
  XOR U13025 ( .A(n12755), .B(n12754), .Z(n12757) );
  NOR U13026 ( .A(n12756), .B(n12757), .Z(n12761) );
  XOR U13027 ( .A(n12758), .B(n12757), .Z(n13240) );
  NOR U13028 ( .A(n123), .B(n49), .Z(n13241) );
  IV U13029 ( .A(n13241), .Z(n12759) );
  NOR U13030 ( .A(n13240), .B(n12759), .Z(n12760) );
  NOR U13031 ( .A(n12761), .B(n12760), .Z(n13248) );
  IV U13032 ( .A(n13248), .Z(n12762) );
  NOR U13033 ( .A(n12763), .B(n12762), .Z(n12764) );
  NOR U13034 ( .A(n12765), .B(n12764), .Z(n12769) );
  IV U13035 ( .A(n12769), .Z(n12767) );
  NOR U13036 ( .A(n126), .B(n49), .Z(n12766) );
  IV U13037 ( .A(n12766), .Z(n12768) );
  NOR U13038 ( .A(n12767), .B(n12768), .Z(n12773) );
  XOR U13039 ( .A(n12769), .B(n12768), .Z(n13254) );
  XOR U13040 ( .A(n12771), .B(n12770), .Z(n13253) );
  NOR U13041 ( .A(n13254), .B(n13253), .Z(n12772) );
  NOR U13042 ( .A(n12773), .B(n12772), .Z(n12778) );
  XOR U13043 ( .A(n12775), .B(n12774), .Z(n12777) );
  IV U13044 ( .A(n12777), .Z(n12776) );
  NOR U13045 ( .A(n12778), .B(n12776), .Z(n12781) );
  XOR U13046 ( .A(n12778), .B(n12777), .Z(n13264) );
  NOR U13047 ( .A(n128), .B(n49), .Z(n13265) );
  IV U13048 ( .A(n13265), .Z(n12779) );
  NOR U13049 ( .A(n13264), .B(n12779), .Z(n12780) );
  NOR U13050 ( .A(n12781), .B(n12780), .Z(n13272) );
  XOR U13051 ( .A(n12783), .B(n12782), .Z(n13271) );
  NOR U13052 ( .A(n13272), .B(n13271), .Z(n12784) );
  NOR U13053 ( .A(n12785), .B(n12784), .Z(n12790) );
  NOR U13054 ( .A(n133), .B(n49), .Z(n12789) );
  IV U13055 ( .A(n12789), .Z(n12786) );
  NOR U13056 ( .A(n12790), .B(n12786), .Z(n12792) );
  XOR U13057 ( .A(n12788), .B(n12787), .Z(n13277) );
  XOR U13058 ( .A(n12790), .B(n12789), .Z(n13276) );
  NOR U13059 ( .A(n13277), .B(n13276), .Z(n12791) );
  NOR U13060 ( .A(n12792), .B(n12791), .Z(n12797) );
  XOR U13061 ( .A(n12794), .B(n12793), .Z(n12796) );
  IV U13062 ( .A(n12796), .Z(n12795) );
  NOR U13063 ( .A(n12797), .B(n12795), .Z(n12800) );
  XOR U13064 ( .A(n12797), .B(n12796), .Z(n12906) );
  NOR U13065 ( .A(n135), .B(n49), .Z(n12907) );
  IV U13066 ( .A(n12907), .Z(n12798) );
  NOR U13067 ( .A(n12906), .B(n12798), .Z(n12799) );
  NOR U13068 ( .A(n12800), .B(n12799), .Z(n13292) );
  XOR U13069 ( .A(n12802), .B(n12801), .Z(n13291) );
  NOR U13070 ( .A(n13292), .B(n13291), .Z(n12803) );
  NOR U13071 ( .A(n12804), .B(n12803), .Z(n12807) );
  NOR U13072 ( .A(n139), .B(n49), .Z(n12806) );
  IV U13073 ( .A(n12806), .Z(n12805) );
  NOR U13074 ( .A(n12807), .B(n12805), .Z(n12811) );
  XOR U13075 ( .A(n12807), .B(n12806), .Z(n13296) );
  XOR U13076 ( .A(n12809), .B(n12808), .Z(n13297) );
  NOR U13077 ( .A(n13296), .B(n13297), .Z(n12810) );
  NOR U13078 ( .A(n12811), .B(n12810), .Z(n12816) );
  XOR U13079 ( .A(n12813), .B(n12812), .Z(n12815) );
  IV U13080 ( .A(n12815), .Z(n12814) );
  NOR U13081 ( .A(n12816), .B(n12814), .Z(n12819) );
  XOR U13082 ( .A(n12816), .B(n12815), .Z(n13307) );
  NOR U13083 ( .A(n141), .B(n49), .Z(n13308) );
  IV U13084 ( .A(n13308), .Z(n12817) );
  NOR U13085 ( .A(n13307), .B(n12817), .Z(n12818) );
  NOR U13086 ( .A(n12819), .B(n12818), .Z(n12821) );
  IV U13087 ( .A(n12821), .Z(n12820) );
  NOR U13088 ( .A(n12822), .B(n12820), .Z(n12824) );
  NOR U13089 ( .A(n143), .B(n49), .Z(n13313) );
  XOR U13090 ( .A(n12822), .B(n12821), .Z(n13312) );
  NOR U13091 ( .A(n13313), .B(n13312), .Z(n12823) );
  NOR U13092 ( .A(n12824), .B(n12823), .Z(n12828) );
  IV U13093 ( .A(n12828), .Z(n12826) );
  NOR U13094 ( .A(n145), .B(n49), .Z(n12825) );
  IV U13095 ( .A(n12825), .Z(n12827) );
  NOR U13096 ( .A(n12826), .B(n12827), .Z(n12832) );
  XOR U13097 ( .A(n12828), .B(n12827), .Z(n13319) );
  XOR U13098 ( .A(n12830), .B(n12829), .Z(n13318) );
  NOR U13099 ( .A(n13319), .B(n13318), .Z(n12831) );
  NOR U13100 ( .A(n12832), .B(n12831), .Z(n12837) );
  XOR U13101 ( .A(n12834), .B(n12833), .Z(n12836) );
  IV U13102 ( .A(n12836), .Z(n12835) );
  NOR U13103 ( .A(n12837), .B(n12835), .Z(n12840) );
  XOR U13104 ( .A(n12837), .B(n12836), .Z(n13329) );
  NOR U13105 ( .A(n147), .B(n49), .Z(n13330) );
  IV U13106 ( .A(n13330), .Z(n12838) );
  NOR U13107 ( .A(n13329), .B(n12838), .Z(n12839) );
  NOR U13108 ( .A(n12840), .B(n12839), .Z(n13334) );
  XOR U13109 ( .A(n12842), .B(n12841), .Z(n13335) );
  NOR U13110 ( .A(n13334), .B(n13335), .Z(n12843) );
  NOR U13111 ( .A(n12844), .B(n12843), .Z(n12847) );
  NOR U13112 ( .A(n150), .B(n49), .Z(n12846) );
  IV U13113 ( .A(n12846), .Z(n12845) );
  NOR U13114 ( .A(n12847), .B(n12845), .Z(n12851) );
  XOR U13115 ( .A(n12847), .B(n12846), .Z(n13341) );
  XOR U13116 ( .A(n12849), .B(n12848), .Z(n13342) );
  NOR U13117 ( .A(n13341), .B(n13342), .Z(n12850) );
  NOR U13118 ( .A(n12851), .B(n12850), .Z(n12856) );
  XOR U13119 ( .A(n12853), .B(n12852), .Z(n12855) );
  IV U13120 ( .A(n12855), .Z(n12854) );
  NOR U13121 ( .A(n12856), .B(n12854), .Z(n12859) );
  XOR U13122 ( .A(n12856), .B(n12855), .Z(n13351) );
  NOR U13123 ( .A(n153), .B(n49), .Z(n12857) );
  IV U13124 ( .A(n12857), .Z(n13350) );
  NOR U13125 ( .A(n13351), .B(n13350), .Z(n12858) );
  NOR U13126 ( .A(n12859), .B(n12858), .Z(n13361) );
  XOR U13127 ( .A(n12861), .B(n12860), .Z(n13360) );
  NOR U13128 ( .A(n13361), .B(n13360), .Z(n12862) );
  NOR U13129 ( .A(n12863), .B(n12862), .Z(n12866) );
  NOR U13130 ( .A(n156), .B(n49), .Z(n12865) );
  IV U13131 ( .A(n12865), .Z(n12864) );
  NOR U13132 ( .A(n12866), .B(n12864), .Z(n12870) );
  XOR U13133 ( .A(n12866), .B(n12865), .Z(n13365) );
  XOR U13134 ( .A(n12868), .B(n12867), .Z(n13366) );
  NOR U13135 ( .A(n13365), .B(n13366), .Z(n12869) );
  NOR U13136 ( .A(n12870), .B(n12869), .Z(n12875) );
  XOR U13137 ( .A(n12872), .B(n12871), .Z(n12874) );
  IV U13138 ( .A(n12874), .Z(n12873) );
  NOR U13139 ( .A(n12875), .B(n12873), .Z(n12878) );
  XOR U13140 ( .A(n12875), .B(n12874), .Z(n13376) );
  NOR U13141 ( .A(n158), .B(n49), .Z(n13377) );
  IV U13142 ( .A(n13377), .Z(n12876) );
  NOR U13143 ( .A(n13376), .B(n12876), .Z(n12877) );
  NOR U13144 ( .A(n12878), .B(n12877), .Z(n13384) );
  XOR U13145 ( .A(n12880), .B(n12879), .Z(n13383) );
  NOR U13146 ( .A(n13384), .B(n13383), .Z(n12881) );
  NOR U13147 ( .A(n12882), .B(n12881), .Z(n12885) );
  NOR U13148 ( .A(n163), .B(n49), .Z(n12884) );
  IV U13149 ( .A(n12884), .Z(n12883) );
  NOR U13150 ( .A(n12885), .B(n12883), .Z(n12889) );
  XOR U13151 ( .A(n12885), .B(n12884), .Z(n13388) );
  XOR U13152 ( .A(n12887), .B(n12886), .Z(n13389) );
  NOR U13153 ( .A(n13388), .B(n13389), .Z(n12888) );
  NOR U13154 ( .A(n12889), .B(n12888), .Z(n12894) );
  XOR U13155 ( .A(n12891), .B(n12890), .Z(n12893) );
  IV U13156 ( .A(n12893), .Z(n12892) );
  NOR U13157 ( .A(n12894), .B(n12892), .Z(n12897) );
  XOR U13158 ( .A(n12894), .B(n12893), .Z(n13399) );
  NOR U13159 ( .A(n165), .B(n49), .Z(n12895) );
  IV U13160 ( .A(n12895), .Z(n13400) );
  NOR U13161 ( .A(n13399), .B(n13400), .Z(n12896) );
  NOR U13162 ( .A(n12897), .B(n12896), .Z(n13404) );
  XOR U13163 ( .A(n12899), .B(n12898), .Z(n13405) );
  NOR U13164 ( .A(n13404), .B(n13405), .Z(n12900) );
  NOR U13165 ( .A(n12901), .B(n12900), .Z(n13407) );
  XOR U13166 ( .A(n12903), .B(n12902), .Z(n13408) );
  NOR U13167 ( .A(n13407), .B(n13408), .Z(n28619) );
  XOR U13168 ( .A(n12905), .B(n12904), .Z(n28618) );
  NOR U13169 ( .A(n28619), .B(n28618), .Z(n28622) );
  NOR U13170 ( .A(n155), .B(n50), .Z(n13353) );
  XOR U13171 ( .A(n12907), .B(n12906), .Z(n13284) );
  NOR U13172 ( .A(n137), .B(n50), .Z(n13285) );
  IV U13173 ( .A(n13285), .Z(n12908) );
  NOR U13174 ( .A(n13284), .B(n12908), .Z(n13287) );
  NOR U13175 ( .A(n119), .B(n50), .Z(n13212) );
  NOR U13176 ( .A(n117), .B(n50), .Z(n13200) );
  NOR U13177 ( .A(n80), .B(n50), .Z(n13188) );
  NOR U13178 ( .A(n81), .B(n50), .Z(n13175) );
  XOR U13179 ( .A(n12910), .B(n12909), .Z(n12911) );
  IV U13180 ( .A(n12911), .Z(n13168) );
  NOR U13181 ( .A(n115), .B(n50), .Z(n13169) );
  IV U13182 ( .A(n13169), .Z(n12912) );
  NOR U13183 ( .A(n13168), .B(n12912), .Z(n13171) );
  NOR U13184 ( .A(n82), .B(n50), .Z(n13165) );
  IV U13185 ( .A(n13165), .Z(n12916) );
  XOR U13186 ( .A(n12914), .B(n12913), .Z(n12915) );
  IV U13187 ( .A(n12915), .Z(n13164) );
  NOR U13188 ( .A(n12916), .B(n13164), .Z(n13167) );
  XOR U13189 ( .A(n12918), .B(n12917), .Z(n12919) );
  IV U13190 ( .A(n12919), .Z(n13160) );
  NOR U13191 ( .A(n114), .B(n50), .Z(n13161) );
  IV U13192 ( .A(n13161), .Z(n12920) );
  NOR U13193 ( .A(n13160), .B(n12920), .Z(n13163) );
  NOR U13194 ( .A(n83), .B(n50), .Z(n13157) );
  IV U13195 ( .A(n13157), .Z(n12924) );
  XOR U13196 ( .A(n12922), .B(n12921), .Z(n12923) );
  IV U13197 ( .A(n12923), .Z(n13156) );
  NOR U13198 ( .A(n12924), .B(n13156), .Z(n13159) );
  XOR U13199 ( .A(n12926), .B(n12925), .Z(n12927) );
  XOR U13200 ( .A(n12928), .B(n12927), .Z(n13152) );
  NOR U13201 ( .A(n113), .B(n50), .Z(n13153) );
  IV U13202 ( .A(n13153), .Z(n12929) );
  NOR U13203 ( .A(n13152), .B(n12929), .Z(n13155) );
  XOR U13204 ( .A(n12931), .B(n12930), .Z(n12932) );
  IV U13205 ( .A(n12932), .Z(n12934) );
  NOR U13206 ( .A(n84), .B(n50), .Z(n12935) );
  IV U13207 ( .A(n12935), .Z(n12933) );
  NOR U13208 ( .A(n12934), .B(n12933), .Z(n13151) );
  XOR U13209 ( .A(n12935), .B(n12934), .Z(n13434) );
  NOR U13210 ( .A(n112), .B(n50), .Z(n13145) );
  XOR U13211 ( .A(n12937), .B(n12936), .Z(n12938) );
  XOR U13212 ( .A(n12939), .B(n12938), .Z(n13146) );
  IV U13213 ( .A(n13146), .Z(n12940) );
  NOR U13214 ( .A(n13145), .B(n12940), .Z(n13148) );
  XOR U13215 ( .A(n12942), .B(n12941), .Z(n13140) );
  NOR U13216 ( .A(n85), .B(n50), .Z(n13141) );
  NOR U13217 ( .A(n13140), .B(n13141), .Z(n13144) );
  XOR U13218 ( .A(n12944), .B(n12943), .Z(n13127) );
  NOR U13219 ( .A(n86), .B(n50), .Z(n13128) );
  IV U13220 ( .A(n13128), .Z(n12945) );
  NOR U13221 ( .A(n13127), .B(n12945), .Z(n13130) );
  XOR U13222 ( .A(n12947), .B(n12946), .Z(n13121) );
  XOR U13223 ( .A(n12949), .B(n12948), .Z(n13117) );
  IV U13224 ( .A(n13117), .Z(n13454) );
  NOR U13225 ( .A(n109), .B(n50), .Z(n13116) );
  IV U13226 ( .A(n13116), .Z(n13453) );
  NOR U13227 ( .A(n13454), .B(n13453), .Z(n13120) );
  XOR U13228 ( .A(n12951), .B(n12950), .Z(n12952) );
  XOR U13229 ( .A(n12953), .B(n12952), .Z(n12955) );
  NOR U13230 ( .A(n108), .B(n50), .Z(n12956) );
  IV U13231 ( .A(n12956), .Z(n12954) );
  NOR U13232 ( .A(n12955), .B(n12954), .Z(n13115) );
  XOR U13233 ( .A(n12956), .B(n12955), .Z(n13458) );
  NOR U13234 ( .A(n87), .B(n50), .Z(n13109) );
  XOR U13235 ( .A(n12958), .B(n12957), .Z(n13110) );
  IV U13236 ( .A(n13110), .Z(n12959) );
  NOR U13237 ( .A(n13109), .B(n12959), .Z(n13112) );
  XOR U13238 ( .A(n12961), .B(n12960), .Z(n12962) );
  NOR U13239 ( .A(n88), .B(n50), .Z(n12963) );
  NOR U13240 ( .A(n12962), .B(n12963), .Z(n13098) );
  IV U13241 ( .A(n12962), .Z(n13464) );
  IV U13242 ( .A(n12963), .Z(n13463) );
  NOR U13243 ( .A(n13464), .B(n13463), .Z(n13096) );
  XOR U13244 ( .A(n12965), .B(n12964), .Z(n13082) );
  IV U13245 ( .A(n13082), .Z(n13473) );
  NOR U13246 ( .A(n105), .B(n50), .Z(n13081) );
  IV U13247 ( .A(n13081), .Z(n13472) );
  NOR U13248 ( .A(n13473), .B(n13472), .Z(n13085) );
  IV U13249 ( .A(n12966), .Z(n12968) );
  XOR U13250 ( .A(n12968), .B(n12967), .Z(n13077) );
  NOR U13251 ( .A(n104), .B(n50), .Z(n13078) );
  IV U13252 ( .A(n13078), .Z(n12969) );
  NOR U13253 ( .A(n13077), .B(n12969), .Z(n13080) );
  IV U13254 ( .A(n12970), .Z(n12972) );
  XOR U13255 ( .A(n12972), .B(n12971), .Z(n13073) );
  NOR U13256 ( .A(n89), .B(n50), .Z(n13074) );
  IV U13257 ( .A(n13074), .Z(n12973) );
  NOR U13258 ( .A(n13073), .B(n12973), .Z(n13076) );
  IV U13259 ( .A(n12974), .Z(n12976) );
  XOR U13260 ( .A(n12976), .B(n12975), .Z(n13068) );
  NOR U13261 ( .A(n103), .B(n50), .Z(n13069) );
  IV U13262 ( .A(n13069), .Z(n12977) );
  NOR U13263 ( .A(n13068), .B(n12977), .Z(n13072) );
  NOR U13264 ( .A(n90), .B(n50), .Z(n13064) );
  XOR U13265 ( .A(n12979), .B(n12978), .Z(n13063) );
  NOR U13266 ( .A(n13064), .B(n13063), .Z(n13067) );
  IV U13267 ( .A(n12980), .Z(n12982) );
  XOR U13268 ( .A(n12982), .B(n12981), .Z(n13058) );
  NOR U13269 ( .A(n102), .B(n50), .Z(n13059) );
  IV U13270 ( .A(n13059), .Z(n12983) );
  NOR U13271 ( .A(n13058), .B(n12983), .Z(n13061) );
  IV U13272 ( .A(n12984), .Z(n12986) );
  XOR U13273 ( .A(n12986), .B(n12985), .Z(n13054) );
  NOR U13274 ( .A(n101), .B(n50), .Z(n13055) );
  IV U13275 ( .A(n13055), .Z(n12987) );
  NOR U13276 ( .A(n13054), .B(n12987), .Z(n13057) );
  IV U13277 ( .A(n12988), .Z(n12990) );
  XOR U13278 ( .A(n12990), .B(n12989), .Z(n13050) );
  NOR U13279 ( .A(n100), .B(n50), .Z(n13051) );
  IV U13280 ( .A(n13051), .Z(n12991) );
  NOR U13281 ( .A(n13050), .B(n12991), .Z(n13053) );
  IV U13282 ( .A(n12992), .Z(n12994) );
  XOR U13283 ( .A(n12994), .B(n12993), .Z(n13046) );
  NOR U13284 ( .A(n99), .B(n50), .Z(n13047) );
  IV U13285 ( .A(n13047), .Z(n12995) );
  NOR U13286 ( .A(n13046), .B(n12995), .Z(n13049) );
  IV U13287 ( .A(n12996), .Z(n12998) );
  XOR U13288 ( .A(n12998), .B(n12997), .Z(n13042) );
  NOR U13289 ( .A(n98), .B(n50), .Z(n13043) );
  IV U13290 ( .A(n13043), .Z(n12999) );
  NOR U13291 ( .A(n13042), .B(n12999), .Z(n13045) );
  XOR U13292 ( .A(n13001), .B(n13000), .Z(n13038) );
  NOR U13293 ( .A(n91), .B(n50), .Z(n13039) );
  IV U13294 ( .A(n13039), .Z(n13002) );
  NOR U13295 ( .A(n13038), .B(n13002), .Z(n13041) );
  XOR U13296 ( .A(n13004), .B(n13003), .Z(n13026) );
  IV U13297 ( .A(n13026), .Z(n13006) );
  NOR U13298 ( .A(n96), .B(n50), .Z(n13005) );
  IV U13299 ( .A(n13005), .Z(n13027) );
  NOR U13300 ( .A(n13006), .B(n13027), .Z(n13029) );
  NOR U13301 ( .A(n95), .B(n50), .Z(n13023) );
  IV U13302 ( .A(n13023), .Z(n13009) );
  XOR U13303 ( .A(n13008), .B(n13007), .Z(n13022) );
  NOR U13304 ( .A(n13009), .B(n13022), .Z(n13025) );
  NOR U13305 ( .A(n50), .B(n93), .Z(n14041) );
  IV U13306 ( .A(n14041), .Z(n13010) );
  NOR U13307 ( .A(n49), .B(n168), .Z(n13018) );
  IV U13308 ( .A(n13018), .Z(n13013) );
  NOR U13309 ( .A(n13010), .B(n13013), .Z(n13011) );
  IV U13310 ( .A(n13011), .Z(n13012) );
  NOR U13311 ( .A(n94), .B(n13012), .Z(n13021) );
  NOR U13312 ( .A(n13013), .B(n93), .Z(n13014) );
  XOR U13313 ( .A(n94), .B(n13014), .Z(n13015) );
  NOR U13314 ( .A(n50), .B(n13015), .Z(n13016) );
  IV U13315 ( .A(n13016), .Z(n13523) );
  XOR U13316 ( .A(n13018), .B(n13017), .Z(n13522) );
  IV U13317 ( .A(n13522), .Z(n13019) );
  NOR U13318 ( .A(n13523), .B(n13019), .Z(n13020) );
  NOR U13319 ( .A(n13021), .B(n13020), .Z(n13519) );
  XOR U13320 ( .A(n13023), .B(n13022), .Z(n13518) );
  NOR U13321 ( .A(n13519), .B(n13518), .Z(n13024) );
  NOR U13322 ( .A(n13025), .B(n13024), .Z(n13549) );
  XOR U13323 ( .A(n13027), .B(n13026), .Z(n13548) );
  NOR U13324 ( .A(n13549), .B(n13548), .Z(n13028) );
  NOR U13325 ( .A(n13029), .B(n13028), .Z(n13034) );
  XOR U13326 ( .A(n13031), .B(n13030), .Z(n13033) );
  IV U13327 ( .A(n13033), .Z(n13032) );
  NOR U13328 ( .A(n13034), .B(n13032), .Z(n13037) );
  XOR U13329 ( .A(n13034), .B(n13033), .Z(n13515) );
  NOR U13330 ( .A(n97), .B(n50), .Z(n13516) );
  IV U13331 ( .A(n13516), .Z(n13035) );
  NOR U13332 ( .A(n13515), .B(n13035), .Z(n13036) );
  NOR U13333 ( .A(n13037), .B(n13036), .Z(n13511) );
  XOR U13334 ( .A(n13039), .B(n13038), .Z(n13512) );
  NOR U13335 ( .A(n13511), .B(n13512), .Z(n13040) );
  NOR U13336 ( .A(n13041), .B(n13040), .Z(n13507) );
  XOR U13337 ( .A(n13043), .B(n13042), .Z(n13508) );
  NOR U13338 ( .A(n13507), .B(n13508), .Z(n13044) );
  NOR U13339 ( .A(n13045), .B(n13044), .Z(n13503) );
  XOR U13340 ( .A(n13047), .B(n13046), .Z(n13504) );
  NOR U13341 ( .A(n13503), .B(n13504), .Z(n13048) );
  NOR U13342 ( .A(n13049), .B(n13048), .Z(n13499) );
  XOR U13343 ( .A(n13051), .B(n13050), .Z(n13500) );
  NOR U13344 ( .A(n13499), .B(n13500), .Z(n13052) );
  NOR U13345 ( .A(n13053), .B(n13052), .Z(n13495) );
  XOR U13346 ( .A(n13055), .B(n13054), .Z(n13496) );
  NOR U13347 ( .A(n13495), .B(n13496), .Z(n13056) );
  NOR U13348 ( .A(n13057), .B(n13056), .Z(n13491) );
  XOR U13349 ( .A(n13059), .B(n13058), .Z(n13492) );
  NOR U13350 ( .A(n13491), .B(n13492), .Z(n13060) );
  NOR U13351 ( .A(n13061), .B(n13060), .Z(n13062) );
  IV U13352 ( .A(n13062), .Z(n13489) );
  XOR U13353 ( .A(n13064), .B(n13063), .Z(n13065) );
  IV U13354 ( .A(n13065), .Z(n13488) );
  NOR U13355 ( .A(n13489), .B(n13488), .Z(n13066) );
  NOR U13356 ( .A(n13067), .B(n13066), .Z(n13486) );
  IV U13357 ( .A(n13486), .Z(n13070) );
  XOR U13358 ( .A(n13069), .B(n13068), .Z(n13485) );
  NOR U13359 ( .A(n13070), .B(n13485), .Z(n13071) );
  NOR U13360 ( .A(n13072), .B(n13071), .Z(n13481) );
  XOR U13361 ( .A(n13074), .B(n13073), .Z(n13482) );
  NOR U13362 ( .A(n13481), .B(n13482), .Z(n13075) );
  NOR U13363 ( .A(n13076), .B(n13075), .Z(n13477) );
  XOR U13364 ( .A(n13078), .B(n13077), .Z(n13478) );
  NOR U13365 ( .A(n13477), .B(n13478), .Z(n13079) );
  NOR U13366 ( .A(n13080), .B(n13079), .Z(n13475) );
  NOR U13367 ( .A(n13082), .B(n13081), .Z(n13083) );
  NOR U13368 ( .A(n13475), .B(n13083), .Z(n13084) );
  NOR U13369 ( .A(n13085), .B(n13084), .Z(n13092) );
  NOR U13370 ( .A(n106), .B(n50), .Z(n13091) );
  IV U13371 ( .A(n13091), .Z(n13086) );
  NOR U13372 ( .A(n13092), .B(n13086), .Z(n13094) );
  XOR U13373 ( .A(n13088), .B(n13087), .Z(n13089) );
  XOR U13374 ( .A(n13090), .B(n13089), .Z(n13471) );
  XOR U13375 ( .A(n13092), .B(n13091), .Z(n13470) );
  NOR U13376 ( .A(n13471), .B(n13470), .Z(n13093) );
  NOR U13377 ( .A(n13094), .B(n13093), .Z(n13466) );
  IV U13378 ( .A(n13466), .Z(n13095) );
  NOR U13379 ( .A(n13096), .B(n13095), .Z(n13097) );
  NOR U13380 ( .A(n13098), .B(n13097), .Z(n13105) );
  IV U13381 ( .A(n13105), .Z(n13100) );
  NOR U13382 ( .A(n107), .B(n50), .Z(n13099) );
  IV U13383 ( .A(n13099), .Z(n13104) );
  NOR U13384 ( .A(n13100), .B(n13104), .Z(n13107) );
  XOR U13385 ( .A(n13102), .B(n13101), .Z(n13103) );
  IV U13386 ( .A(n13103), .Z(n13461) );
  XOR U13387 ( .A(n13105), .B(n13104), .Z(n13462) );
  NOR U13388 ( .A(n13461), .B(n13462), .Z(n13106) );
  NOR U13389 ( .A(n13107), .B(n13106), .Z(n13108) );
  IV U13390 ( .A(n13108), .Z(n13617) );
  XOR U13391 ( .A(n13110), .B(n13109), .Z(n13616) );
  NOR U13392 ( .A(n13617), .B(n13616), .Z(n13111) );
  NOR U13393 ( .A(n13112), .B(n13111), .Z(n13459) );
  IV U13394 ( .A(n13459), .Z(n13113) );
  NOR U13395 ( .A(n13458), .B(n13113), .Z(n13114) );
  NOR U13396 ( .A(n13115), .B(n13114), .Z(n13456) );
  NOR U13397 ( .A(n13117), .B(n13116), .Z(n13118) );
  NOR U13398 ( .A(n13456), .B(n13118), .Z(n13119) );
  NOR U13399 ( .A(n13120), .B(n13119), .Z(n13122) );
  NOR U13400 ( .A(n13121), .B(n13122), .Z(n13126) );
  XOR U13401 ( .A(n13122), .B(n13121), .Z(n13449) );
  IV U13402 ( .A(n13449), .Z(n13124) );
  NOR U13403 ( .A(n110), .B(n50), .Z(n13448) );
  IV U13404 ( .A(n13448), .Z(n13123) );
  NOR U13405 ( .A(n13124), .B(n13123), .Z(n13125) );
  NOR U13406 ( .A(n13126), .B(n13125), .Z(n13444) );
  XOR U13407 ( .A(n13128), .B(n13127), .Z(n13445) );
  NOR U13408 ( .A(n13444), .B(n13445), .Z(n13129) );
  NOR U13409 ( .A(n13130), .B(n13129), .Z(n13136) );
  NOR U13410 ( .A(n111), .B(n50), .Z(n13135) );
  IV U13411 ( .A(n13135), .Z(n13131) );
  NOR U13412 ( .A(n13136), .B(n13131), .Z(n13138) );
  XOR U13413 ( .A(n13133), .B(n13132), .Z(n13134) );
  IV U13414 ( .A(n13134), .Z(n13441) );
  XOR U13415 ( .A(n13136), .B(n13135), .Z(n13440) );
  NOR U13416 ( .A(n13441), .B(n13440), .Z(n13137) );
  NOR U13417 ( .A(n13138), .B(n13137), .Z(n13139) );
  IV U13418 ( .A(n13139), .Z(n13645) );
  XOR U13419 ( .A(n13141), .B(n13140), .Z(n13142) );
  IV U13420 ( .A(n13142), .Z(n13644) );
  NOR U13421 ( .A(n13645), .B(n13644), .Z(n13143) );
  NOR U13422 ( .A(n13144), .B(n13143), .Z(n13438) );
  XOR U13423 ( .A(n13146), .B(n13145), .Z(n13437) );
  NOR U13424 ( .A(n13438), .B(n13437), .Z(n13147) );
  NOR U13425 ( .A(n13148), .B(n13147), .Z(n13435) );
  IV U13426 ( .A(n13435), .Z(n13149) );
  NOR U13427 ( .A(n13434), .B(n13149), .Z(n13150) );
  NOR U13428 ( .A(n13151), .B(n13150), .Z(n13431) );
  XOR U13429 ( .A(n13153), .B(n13152), .Z(n13430) );
  NOR U13430 ( .A(n13431), .B(n13430), .Z(n13154) );
  NOR U13431 ( .A(n13155), .B(n13154), .Z(n13427) );
  XOR U13432 ( .A(n13157), .B(n13156), .Z(n13428) );
  NOR U13433 ( .A(n13427), .B(n13428), .Z(n13158) );
  NOR U13434 ( .A(n13159), .B(n13158), .Z(n13424) );
  XOR U13435 ( .A(n13161), .B(n13160), .Z(n13423) );
  NOR U13436 ( .A(n13424), .B(n13423), .Z(n13162) );
  NOR U13437 ( .A(n13163), .B(n13162), .Z(n13419) );
  XOR U13438 ( .A(n13165), .B(n13164), .Z(n13420) );
  NOR U13439 ( .A(n13419), .B(n13420), .Z(n13166) );
  NOR U13440 ( .A(n13167), .B(n13166), .Z(n13416) );
  XOR U13441 ( .A(n13169), .B(n13168), .Z(n13415) );
  NOR U13442 ( .A(n13416), .B(n13415), .Z(n13170) );
  NOR U13443 ( .A(n13171), .B(n13170), .Z(n13176) );
  IV U13444 ( .A(n13176), .Z(n13172) );
  NOR U13445 ( .A(n13175), .B(n13172), .Z(n13178) );
  XOR U13446 ( .A(n13174), .B(n13173), .Z(n13684) );
  XOR U13447 ( .A(n13176), .B(n13175), .Z(n13683) );
  NOR U13448 ( .A(n13684), .B(n13683), .Z(n13177) );
  NOR U13449 ( .A(n13178), .B(n13177), .Z(n13184) );
  IV U13450 ( .A(n13184), .Z(n13182) );
  IV U13451 ( .A(n13179), .Z(n13181) );
  XOR U13452 ( .A(n13181), .B(n13180), .Z(n13183) );
  NOR U13453 ( .A(n13182), .B(n13183), .Z(n13187) );
  XOR U13454 ( .A(n13184), .B(n13183), .Z(n13692) );
  NOR U13455 ( .A(n116), .B(n50), .Z(n13185) );
  IV U13456 ( .A(n13185), .Z(n13691) );
  NOR U13457 ( .A(n13692), .B(n13691), .Z(n13186) );
  NOR U13458 ( .A(n13187), .B(n13186), .Z(n13189) );
  IV U13459 ( .A(n13189), .Z(n13698) );
  NOR U13460 ( .A(n13188), .B(n13698), .Z(n13194) );
  IV U13461 ( .A(n13188), .Z(n13699) );
  NOR U13462 ( .A(n13189), .B(n13699), .Z(n13192) );
  XOR U13463 ( .A(n13191), .B(n13190), .Z(n13701) );
  NOR U13464 ( .A(n13192), .B(n13701), .Z(n13193) );
  NOR U13465 ( .A(n13194), .B(n13193), .Z(n13199) );
  NOR U13466 ( .A(n13200), .B(n13199), .Z(n13203) );
  XOR U13467 ( .A(n13196), .B(n13195), .Z(n13197) );
  XOR U13468 ( .A(n13198), .B(n13197), .Z(n13707) );
  XOR U13469 ( .A(n13200), .B(n13199), .Z(n13201) );
  IV U13470 ( .A(n13201), .Z(n13706) );
  NOR U13471 ( .A(n13707), .B(n13706), .Z(n13202) );
  NOR U13472 ( .A(n13203), .B(n13202), .Z(n13207) );
  IV U13473 ( .A(n13207), .Z(n13717) );
  XOR U13474 ( .A(n13205), .B(n13204), .Z(n13206) );
  IV U13475 ( .A(n13206), .Z(n13716) );
  NOR U13476 ( .A(n13717), .B(n13716), .Z(n13211) );
  NOR U13477 ( .A(n13207), .B(n13206), .Z(n13209) );
  NOR U13478 ( .A(n79), .B(n50), .Z(n13719) );
  IV U13479 ( .A(n13719), .Z(n13208) );
  NOR U13480 ( .A(n13209), .B(n13208), .Z(n13210) );
  NOR U13481 ( .A(n13211), .B(n13210), .Z(n13213) );
  IV U13482 ( .A(n13213), .Z(n13725) );
  NOR U13483 ( .A(n13212), .B(n13725), .Z(n13218) );
  IV U13484 ( .A(n13212), .Z(n13726) );
  NOR U13485 ( .A(n13213), .B(n13726), .Z(n13216) );
  XOR U13486 ( .A(n13215), .B(n13214), .Z(n13728) );
  NOR U13487 ( .A(n13216), .B(n13728), .Z(n13217) );
  NOR U13488 ( .A(n13218), .B(n13217), .Z(n13226) );
  IV U13489 ( .A(n13226), .Z(n13220) );
  NOR U13490 ( .A(n120), .B(n50), .Z(n13219) );
  IV U13491 ( .A(n13219), .Z(n13225) );
  NOR U13492 ( .A(n13220), .B(n13225), .Z(n13228) );
  XOR U13493 ( .A(n13222), .B(n13221), .Z(n13223) );
  XOR U13494 ( .A(n13224), .B(n13223), .Z(n13734) );
  XOR U13495 ( .A(n13226), .B(n13225), .Z(n13733) );
  NOR U13496 ( .A(n13734), .B(n13733), .Z(n13227) );
  NOR U13497 ( .A(n13228), .B(n13227), .Z(n13231) );
  XOR U13498 ( .A(n13230), .B(n13229), .Z(n13232) );
  NOR U13499 ( .A(n13231), .B(n13232), .Z(n13236) );
  IV U13500 ( .A(n13231), .Z(n13233) );
  XOR U13501 ( .A(n13233), .B(n13232), .Z(n13741) );
  NOR U13502 ( .A(n123), .B(n50), .Z(n13234) );
  IV U13503 ( .A(n13234), .Z(n13742) );
  NOR U13504 ( .A(n13741), .B(n13742), .Z(n13235) );
  NOR U13505 ( .A(n13236), .B(n13235), .Z(n13239) );
  NOR U13506 ( .A(n125), .B(n50), .Z(n13238) );
  IV U13507 ( .A(n13238), .Z(n13237) );
  NOR U13508 ( .A(n13239), .B(n13237), .Z(n13243) );
  XOR U13509 ( .A(n13239), .B(n13238), .Z(n13750) );
  XOR U13510 ( .A(n13241), .B(n13240), .Z(n13751) );
  NOR U13511 ( .A(n13750), .B(n13751), .Z(n13242) );
  NOR U13512 ( .A(n13243), .B(n13242), .Z(n13250) );
  NOR U13513 ( .A(n126), .B(n50), .Z(n13249) );
  IV U13514 ( .A(n13249), .Z(n13244) );
  NOR U13515 ( .A(n13250), .B(n13244), .Z(n13252) );
  XOR U13516 ( .A(n13246), .B(n13245), .Z(n13247) );
  XOR U13517 ( .A(n13248), .B(n13247), .Z(n13758) );
  XOR U13518 ( .A(n13250), .B(n13249), .Z(n13757) );
  NOR U13519 ( .A(n13758), .B(n13757), .Z(n13251) );
  NOR U13520 ( .A(n13252), .B(n13251), .Z(n13257) );
  XOR U13521 ( .A(n13254), .B(n13253), .Z(n13256) );
  IV U13522 ( .A(n13256), .Z(n13255) );
  NOR U13523 ( .A(n13257), .B(n13255), .Z(n13260) );
  XOR U13524 ( .A(n13257), .B(n13256), .Z(n13412) );
  NOR U13525 ( .A(n128), .B(n50), .Z(n13413) );
  IV U13526 ( .A(n13413), .Z(n13258) );
  NOR U13527 ( .A(n13412), .B(n13258), .Z(n13259) );
  NOR U13528 ( .A(n13260), .B(n13259), .Z(n13263) );
  NOR U13529 ( .A(n131), .B(n50), .Z(n13262) );
  IV U13530 ( .A(n13262), .Z(n13261) );
  NOR U13531 ( .A(n13263), .B(n13261), .Z(n13267) );
  XOR U13532 ( .A(n13263), .B(n13262), .Z(n13772) );
  XOR U13533 ( .A(n13265), .B(n13264), .Z(n13773) );
  NOR U13534 ( .A(n13772), .B(n13773), .Z(n13266) );
  NOR U13535 ( .A(n13267), .B(n13266), .Z(n13270) );
  NOR U13536 ( .A(n133), .B(n50), .Z(n13269) );
  IV U13537 ( .A(n13269), .Z(n13268) );
  NOR U13538 ( .A(n13270), .B(n13268), .Z(n13275) );
  XOR U13539 ( .A(n13270), .B(n13269), .Z(n13777) );
  XOR U13540 ( .A(n13272), .B(n13271), .Z(n13778) );
  IV U13541 ( .A(n13778), .Z(n13273) );
  NOR U13542 ( .A(n13777), .B(n13273), .Z(n13274) );
  NOR U13543 ( .A(n13275), .B(n13274), .Z(n13280) );
  XOR U13544 ( .A(n13277), .B(n13276), .Z(n13279) );
  IV U13545 ( .A(n13279), .Z(n13278) );
  NOR U13546 ( .A(n13280), .B(n13278), .Z(n13283) );
  XOR U13547 ( .A(n13280), .B(n13279), .Z(n13788) );
  NOR U13548 ( .A(n135), .B(n50), .Z(n13789) );
  IV U13549 ( .A(n13789), .Z(n13281) );
  NOR U13550 ( .A(n13788), .B(n13281), .Z(n13282) );
  NOR U13551 ( .A(n13283), .B(n13282), .Z(n13796) );
  XOR U13552 ( .A(n13285), .B(n13284), .Z(n13795) );
  NOR U13553 ( .A(n13796), .B(n13795), .Z(n13286) );
  NOR U13554 ( .A(n13287), .B(n13286), .Z(n13290) );
  NOR U13555 ( .A(n139), .B(n50), .Z(n13289) );
  IV U13556 ( .A(n13289), .Z(n13288) );
  NOR U13557 ( .A(n13290), .B(n13288), .Z(n13295) );
  XOR U13558 ( .A(n13290), .B(n13289), .Z(n13800) );
  XOR U13559 ( .A(n13292), .B(n13291), .Z(n13801) );
  IV U13560 ( .A(n13801), .Z(n13293) );
  NOR U13561 ( .A(n13800), .B(n13293), .Z(n13294) );
  NOR U13562 ( .A(n13295), .B(n13294), .Z(n13300) );
  XOR U13563 ( .A(n13297), .B(n13296), .Z(n13299) );
  IV U13564 ( .A(n13299), .Z(n13298) );
  NOR U13565 ( .A(n13300), .B(n13298), .Z(n13303) );
  XOR U13566 ( .A(n13300), .B(n13299), .Z(n13811) );
  NOR U13567 ( .A(n141), .B(n50), .Z(n13812) );
  IV U13568 ( .A(n13812), .Z(n13301) );
  NOR U13569 ( .A(n13811), .B(n13301), .Z(n13302) );
  NOR U13570 ( .A(n13303), .B(n13302), .Z(n13306) );
  NOR U13571 ( .A(n143), .B(n50), .Z(n13305) );
  IV U13572 ( .A(n13305), .Z(n13304) );
  NOR U13573 ( .A(n13306), .B(n13304), .Z(n13310) );
  XOR U13574 ( .A(n13306), .B(n13305), .Z(n13816) );
  XOR U13575 ( .A(n13308), .B(n13307), .Z(n13817) );
  NOR U13576 ( .A(n13816), .B(n13817), .Z(n13309) );
  NOR U13577 ( .A(n13310), .B(n13309), .Z(n13315) );
  NOR U13578 ( .A(n145), .B(n50), .Z(n13314) );
  IV U13579 ( .A(n13314), .Z(n13311) );
  NOR U13580 ( .A(n13315), .B(n13311), .Z(n13317) );
  XOR U13581 ( .A(n13313), .B(n13312), .Z(n13824) );
  XOR U13582 ( .A(n13315), .B(n13314), .Z(n13823) );
  NOR U13583 ( .A(n13824), .B(n13823), .Z(n13316) );
  NOR U13584 ( .A(n13317), .B(n13316), .Z(n13322) );
  XOR U13585 ( .A(n13319), .B(n13318), .Z(n13321) );
  IV U13586 ( .A(n13321), .Z(n13320) );
  NOR U13587 ( .A(n13322), .B(n13320), .Z(n13325) );
  XOR U13588 ( .A(n13322), .B(n13321), .Z(n13831) );
  NOR U13589 ( .A(n147), .B(n50), .Z(n13832) );
  IV U13590 ( .A(n13832), .Z(n13323) );
  NOR U13591 ( .A(n13831), .B(n13323), .Z(n13324) );
  NOR U13592 ( .A(n13325), .B(n13324), .Z(n13328) );
  NOR U13593 ( .A(n148), .B(n50), .Z(n13327) );
  IV U13594 ( .A(n13327), .Z(n13326) );
  NOR U13595 ( .A(n13328), .B(n13326), .Z(n13332) );
  XOR U13596 ( .A(n13328), .B(n13327), .Z(n13842) );
  XOR U13597 ( .A(n13330), .B(n13329), .Z(n13843) );
  NOR U13598 ( .A(n13842), .B(n13843), .Z(n13331) );
  NOR U13599 ( .A(n13332), .B(n13331), .Z(n13338) );
  NOR U13600 ( .A(n150), .B(n50), .Z(n13337) );
  IV U13601 ( .A(n13337), .Z(n13333) );
  NOR U13602 ( .A(n13338), .B(n13333), .Z(n13340) );
  IV U13603 ( .A(n13334), .Z(n13336) );
  XOR U13604 ( .A(n13336), .B(n13335), .Z(n13411) );
  XOR U13605 ( .A(n13338), .B(n13337), .Z(n13410) );
  NOR U13606 ( .A(n13411), .B(n13410), .Z(n13339) );
  NOR U13607 ( .A(n13340), .B(n13339), .Z(n13345) );
  XOR U13608 ( .A(n13342), .B(n13341), .Z(n13344) );
  IV U13609 ( .A(n13344), .Z(n13343) );
  NOR U13610 ( .A(n13345), .B(n13343), .Z(n13348) );
  XOR U13611 ( .A(n13345), .B(n13344), .Z(n13853) );
  NOR U13612 ( .A(n153), .B(n50), .Z(n13346) );
  IV U13613 ( .A(n13346), .Z(n13852) );
  NOR U13614 ( .A(n13853), .B(n13852), .Z(n13347) );
  NOR U13615 ( .A(n13348), .B(n13347), .Z(n13352) );
  IV U13616 ( .A(n13352), .Z(n13349) );
  NOR U13617 ( .A(n13353), .B(n13349), .Z(n13355) );
  XOR U13618 ( .A(n13351), .B(n13350), .Z(n13862) );
  XOR U13619 ( .A(n13353), .B(n13352), .Z(n13861) );
  NOR U13620 ( .A(n13862), .B(n13861), .Z(n13354) );
  NOR U13621 ( .A(n13355), .B(n13354), .Z(n13359) );
  IV U13622 ( .A(n13359), .Z(n13357) );
  NOR U13623 ( .A(n156), .B(n50), .Z(n13356) );
  IV U13624 ( .A(n13356), .Z(n13358) );
  NOR U13625 ( .A(n13357), .B(n13358), .Z(n13364) );
  XOR U13626 ( .A(n13359), .B(n13358), .Z(n13868) );
  XOR U13627 ( .A(n13361), .B(n13360), .Z(n13867) );
  IV U13628 ( .A(n13867), .Z(n13362) );
  NOR U13629 ( .A(n13868), .B(n13362), .Z(n13363) );
  NOR U13630 ( .A(n13364), .B(n13363), .Z(n13369) );
  XOR U13631 ( .A(n13366), .B(n13365), .Z(n13368) );
  IV U13632 ( .A(n13368), .Z(n13367) );
  NOR U13633 ( .A(n13369), .B(n13367), .Z(n13372) );
  XOR U13634 ( .A(n13369), .B(n13368), .Z(n13878) );
  NOR U13635 ( .A(n158), .B(n50), .Z(n13879) );
  IV U13636 ( .A(n13879), .Z(n13370) );
  NOR U13637 ( .A(n13878), .B(n13370), .Z(n13371) );
  NOR U13638 ( .A(n13372), .B(n13371), .Z(n13375) );
  NOR U13639 ( .A(n161), .B(n50), .Z(n13374) );
  IV U13640 ( .A(n13374), .Z(n13373) );
  NOR U13641 ( .A(n13375), .B(n13373), .Z(n13379) );
  XOR U13642 ( .A(n13375), .B(n13374), .Z(n13883) );
  XOR U13643 ( .A(n13377), .B(n13376), .Z(n13884) );
  NOR U13644 ( .A(n13883), .B(n13884), .Z(n13378) );
  NOR U13645 ( .A(n13379), .B(n13378), .Z(n13382) );
  NOR U13646 ( .A(n163), .B(n50), .Z(n13381) );
  IV U13647 ( .A(n13381), .Z(n13380) );
  NOR U13648 ( .A(n13382), .B(n13380), .Z(n13387) );
  XOR U13649 ( .A(n13382), .B(n13381), .Z(n13890) );
  XOR U13650 ( .A(n13384), .B(n13383), .Z(n13891) );
  IV U13651 ( .A(n13891), .Z(n13385) );
  NOR U13652 ( .A(n13890), .B(n13385), .Z(n13386) );
  NOR U13653 ( .A(n13387), .B(n13386), .Z(n13392) );
  XOR U13654 ( .A(n13389), .B(n13388), .Z(n13391) );
  IV U13655 ( .A(n13391), .Z(n13390) );
  NOR U13656 ( .A(n13392), .B(n13390), .Z(n13395) );
  XOR U13657 ( .A(n13392), .B(n13391), .Z(n13901) );
  NOR U13658 ( .A(n165), .B(n50), .Z(n13393) );
  IV U13659 ( .A(n13393), .Z(n13902) );
  NOR U13660 ( .A(n13901), .B(n13902), .Z(n13394) );
  NOR U13661 ( .A(n13395), .B(n13394), .Z(n13398) );
  NOR U13662 ( .A(n167), .B(n50), .Z(n13397) );
  IV U13663 ( .A(n13397), .Z(n13396) );
  NOR U13664 ( .A(n13398), .B(n13396), .Z(n13403) );
  XOR U13665 ( .A(n13398), .B(n13397), .Z(n13906) );
  XOR U13666 ( .A(n13400), .B(n13399), .Z(n13907) );
  IV U13667 ( .A(n13907), .Z(n13401) );
  NOR U13668 ( .A(n13906), .B(n13401), .Z(n13402) );
  NOR U13669 ( .A(n13403), .B(n13402), .Z(n13909) );
  IV U13670 ( .A(n13404), .Z(n13406) );
  XOR U13671 ( .A(n13406), .B(n13405), .Z(n13908) );
  NOR U13672 ( .A(n13909), .B(n13908), .Z(n31648) );
  IV U13673 ( .A(n13407), .Z(n13409) );
  XOR U13674 ( .A(n13409), .B(n13408), .Z(n31655) );
  XOR U13675 ( .A(n31648), .B(n31655), .Z(n28614) );
  XOR U13676 ( .A(n13411), .B(n13410), .Z(n13849) );
  XOR U13677 ( .A(n13413), .B(n13412), .Z(n13765) );
  NOR U13678 ( .A(n131), .B(n51), .Z(n13766) );
  IV U13679 ( .A(n13766), .Z(n13414) );
  NOR U13680 ( .A(n13765), .B(n13414), .Z(n13768) );
  NOR U13681 ( .A(n119), .B(n51), .Z(n13714) );
  NOR U13682 ( .A(n80), .B(n51), .Z(n13689) );
  XOR U13683 ( .A(n13416), .B(n13415), .Z(n13930) );
  NOR U13684 ( .A(n81), .B(n51), .Z(n13417) );
  NOR U13685 ( .A(n13930), .B(n13417), .Z(n13680) );
  IV U13686 ( .A(n13930), .Z(n13418) );
  IV U13687 ( .A(n13417), .Z(n13928) );
  NOR U13688 ( .A(n13418), .B(n13928), .Z(n13678) );
  XOR U13689 ( .A(n13420), .B(n13419), .Z(n13421) );
  IV U13690 ( .A(n13421), .Z(n13673) );
  NOR U13691 ( .A(n115), .B(n51), .Z(n13674) );
  IV U13692 ( .A(n13674), .Z(n13422) );
  NOR U13693 ( .A(n13673), .B(n13422), .Z(n13676) );
  NOR U13694 ( .A(n82), .B(n51), .Z(n13669) );
  IV U13695 ( .A(n13669), .Z(n13426) );
  XOR U13696 ( .A(n13424), .B(n13423), .Z(n13668) );
  IV U13697 ( .A(n13668), .Z(n13425) );
  NOR U13698 ( .A(n13426), .B(n13425), .Z(n13672) );
  XOR U13699 ( .A(n13428), .B(n13427), .Z(n13429) );
  IV U13700 ( .A(n13429), .Z(n13663) );
  XOR U13701 ( .A(n13431), .B(n13430), .Z(n13432) );
  NOR U13702 ( .A(n83), .B(n51), .Z(n13433) );
  NOR U13703 ( .A(n13432), .B(n13433), .Z(n13661) );
  IV U13704 ( .A(n13432), .Z(n14179) );
  IV U13705 ( .A(n13433), .Z(n14178) );
  NOR U13706 ( .A(n14179), .B(n14178), .Z(n13659) );
  XOR U13707 ( .A(n13435), .B(n13434), .Z(n13654) );
  NOR U13708 ( .A(n113), .B(n51), .Z(n13655) );
  IV U13709 ( .A(n13655), .Z(n13436) );
  NOR U13710 ( .A(n13654), .B(n13436), .Z(n13657) );
  XOR U13711 ( .A(n13438), .B(n13437), .Z(n13651) );
  NOR U13712 ( .A(n84), .B(n51), .Z(n13650) );
  IV U13713 ( .A(n13650), .Z(n13439) );
  NOR U13714 ( .A(n13651), .B(n13439), .Z(n13653) );
  XOR U13715 ( .A(n13441), .B(n13440), .Z(n13442) );
  NOR U13716 ( .A(n85), .B(n51), .Z(n13443) );
  NOR U13717 ( .A(n13442), .B(n13443), .Z(n13641) );
  IV U13718 ( .A(n13442), .Z(n14159) );
  IV U13719 ( .A(n13443), .Z(n14158) );
  NOR U13720 ( .A(n14159), .B(n14158), .Z(n13639) );
  IV U13721 ( .A(n13444), .Z(n13446) );
  XOR U13722 ( .A(n13446), .B(n13445), .Z(n13633) );
  NOR U13723 ( .A(n111), .B(n51), .Z(n13634) );
  IV U13724 ( .A(n13634), .Z(n13447) );
  NOR U13725 ( .A(n13633), .B(n13447), .Z(n13637) );
  NOR U13726 ( .A(n86), .B(n51), .Z(n13451) );
  XOR U13727 ( .A(n13449), .B(n13448), .Z(n13450) );
  NOR U13728 ( .A(n13451), .B(n13450), .Z(n13632) );
  XOR U13729 ( .A(n13451), .B(n13450), .Z(n13452) );
  IV U13730 ( .A(n13452), .Z(n13956) );
  XOR U13731 ( .A(n13454), .B(n13453), .Z(n13455) );
  XOR U13732 ( .A(n13456), .B(n13455), .Z(n13627) );
  NOR U13733 ( .A(n110), .B(n51), .Z(n13626) );
  IV U13734 ( .A(n13626), .Z(n13457) );
  NOR U13735 ( .A(n13627), .B(n13457), .Z(n13629) );
  NOR U13736 ( .A(n109), .B(n51), .Z(n13623) );
  IV U13737 ( .A(n13623), .Z(n13460) );
  XOR U13738 ( .A(n13459), .B(n13458), .Z(n13622) );
  NOR U13739 ( .A(n13460), .B(n13622), .Z(n13625) );
  XOR U13740 ( .A(n13462), .B(n13461), .Z(n13611) );
  IV U13741 ( .A(n13611), .Z(n13969) );
  NOR U13742 ( .A(n87), .B(n51), .Z(n13610) );
  IV U13743 ( .A(n13610), .Z(n13968) );
  NOR U13744 ( .A(n13969), .B(n13968), .Z(n13614) );
  XOR U13745 ( .A(n13464), .B(n13463), .Z(n13465) );
  XOR U13746 ( .A(n13466), .B(n13465), .Z(n13469) );
  NOR U13747 ( .A(n107), .B(n51), .Z(n13468) );
  IV U13748 ( .A(n13468), .Z(n13467) );
  NOR U13749 ( .A(n13469), .B(n13467), .Z(n13609) );
  XOR U13750 ( .A(n13469), .B(n13468), .Z(n13974) );
  NOR U13751 ( .A(n88), .B(n51), .Z(n13603) );
  XOR U13752 ( .A(n13471), .B(n13470), .Z(n13602) );
  NOR U13753 ( .A(n13603), .B(n13602), .Z(n13606) );
  XOR U13754 ( .A(n13473), .B(n13472), .Z(n13474) );
  XOR U13755 ( .A(n13475), .B(n13474), .Z(n13598) );
  NOR U13756 ( .A(n106), .B(n51), .Z(n13597) );
  IV U13757 ( .A(n13597), .Z(n13476) );
  NOR U13758 ( .A(n13598), .B(n13476), .Z(n13600) );
  IV U13759 ( .A(n13477), .Z(n13479) );
  XOR U13760 ( .A(n13479), .B(n13478), .Z(n13593) );
  NOR U13761 ( .A(n105), .B(n51), .Z(n13594) );
  IV U13762 ( .A(n13594), .Z(n13480) );
  NOR U13763 ( .A(n13593), .B(n13480), .Z(n13596) );
  IV U13764 ( .A(n13481), .Z(n13483) );
  XOR U13765 ( .A(n13483), .B(n13482), .Z(n13589) );
  NOR U13766 ( .A(n104), .B(n51), .Z(n13590) );
  IV U13767 ( .A(n13590), .Z(n13484) );
  NOR U13768 ( .A(n13589), .B(n13484), .Z(n13592) );
  XOR U13769 ( .A(n13486), .B(n13485), .Z(n13585) );
  NOR U13770 ( .A(n89), .B(n51), .Z(n13586) );
  IV U13771 ( .A(n13586), .Z(n13487) );
  NOR U13772 ( .A(n13585), .B(n13487), .Z(n13588) );
  XOR U13773 ( .A(n13489), .B(n13488), .Z(n13582) );
  NOR U13774 ( .A(n103), .B(n51), .Z(n13581) );
  IV U13775 ( .A(n13581), .Z(n13490) );
  NOR U13776 ( .A(n13582), .B(n13490), .Z(n13584) );
  IV U13777 ( .A(n13491), .Z(n13493) );
  XOR U13778 ( .A(n13493), .B(n13492), .Z(n13577) );
  NOR U13779 ( .A(n90), .B(n51), .Z(n13578) );
  IV U13780 ( .A(n13578), .Z(n13494) );
  NOR U13781 ( .A(n13577), .B(n13494), .Z(n13580) );
  IV U13782 ( .A(n13495), .Z(n13497) );
  XOR U13783 ( .A(n13497), .B(n13496), .Z(n13573) );
  NOR U13784 ( .A(n102), .B(n51), .Z(n13574) );
  IV U13785 ( .A(n13574), .Z(n13498) );
  NOR U13786 ( .A(n13573), .B(n13498), .Z(n13576) );
  IV U13787 ( .A(n13499), .Z(n13501) );
  XOR U13788 ( .A(n13501), .B(n13500), .Z(n13569) );
  NOR U13789 ( .A(n101), .B(n51), .Z(n13570) );
  IV U13790 ( .A(n13570), .Z(n13502) );
  NOR U13791 ( .A(n13569), .B(n13502), .Z(n13572) );
  IV U13792 ( .A(n13503), .Z(n13505) );
  XOR U13793 ( .A(n13505), .B(n13504), .Z(n13565) );
  NOR U13794 ( .A(n100), .B(n51), .Z(n13566) );
  IV U13795 ( .A(n13566), .Z(n13506) );
  NOR U13796 ( .A(n13565), .B(n13506), .Z(n13568) );
  IV U13797 ( .A(n13507), .Z(n13509) );
  XOR U13798 ( .A(n13509), .B(n13508), .Z(n13561) );
  NOR U13799 ( .A(n99), .B(n51), .Z(n13562) );
  IV U13800 ( .A(n13562), .Z(n13510) );
  NOR U13801 ( .A(n13561), .B(n13510), .Z(n13564) );
  IV U13802 ( .A(n13511), .Z(n13513) );
  XOR U13803 ( .A(n13513), .B(n13512), .Z(n13557) );
  NOR U13804 ( .A(n98), .B(n51), .Z(n13558) );
  IV U13805 ( .A(n13558), .Z(n13514) );
  NOR U13806 ( .A(n13557), .B(n13514), .Z(n13560) );
  XOR U13807 ( .A(n13516), .B(n13515), .Z(n13553) );
  NOR U13808 ( .A(n91), .B(n51), .Z(n13554) );
  IV U13809 ( .A(n13554), .Z(n13517) );
  NOR U13810 ( .A(n13553), .B(n13517), .Z(n13556) );
  XOR U13811 ( .A(n13519), .B(n13518), .Z(n13541) );
  IV U13812 ( .A(n13541), .Z(n13521) );
  NOR U13813 ( .A(n96), .B(n51), .Z(n13520) );
  IV U13814 ( .A(n13520), .Z(n13542) );
  NOR U13815 ( .A(n13521), .B(n13542), .Z(n13544) );
  NOR U13816 ( .A(n95), .B(n51), .Z(n13538) );
  IV U13817 ( .A(n13538), .Z(n13524) );
  XOR U13818 ( .A(n13523), .B(n13522), .Z(n13537) );
  NOR U13819 ( .A(n13524), .B(n13537), .Z(n13540) );
  NOR U13820 ( .A(n51), .B(n93), .Z(n14552) );
  IV U13821 ( .A(n14552), .Z(n13525) );
  NOR U13822 ( .A(n50), .B(n168), .Z(n13533) );
  IV U13823 ( .A(n13533), .Z(n13528) );
  NOR U13824 ( .A(n13525), .B(n13528), .Z(n13526) );
  IV U13825 ( .A(n13526), .Z(n13527) );
  NOR U13826 ( .A(n94), .B(n13527), .Z(n13536) );
  NOR U13827 ( .A(n13528), .B(n93), .Z(n13529) );
  XOR U13828 ( .A(n94), .B(n13529), .Z(n13530) );
  NOR U13829 ( .A(n51), .B(n13530), .Z(n13531) );
  IV U13830 ( .A(n13531), .Z(n14032) );
  XOR U13831 ( .A(n13533), .B(n13532), .Z(n14031) );
  IV U13832 ( .A(n14031), .Z(n13534) );
  NOR U13833 ( .A(n14032), .B(n13534), .Z(n13535) );
  NOR U13834 ( .A(n13536), .B(n13535), .Z(n14028) );
  XOR U13835 ( .A(n13538), .B(n13537), .Z(n14027) );
  NOR U13836 ( .A(n14028), .B(n14027), .Z(n13539) );
  NOR U13837 ( .A(n13540), .B(n13539), .Z(n14055) );
  XOR U13838 ( .A(n13542), .B(n13541), .Z(n14054) );
  NOR U13839 ( .A(n14055), .B(n14054), .Z(n13543) );
  NOR U13840 ( .A(n13544), .B(n13543), .Z(n13547) );
  NOR U13841 ( .A(n97), .B(n51), .Z(n13546) );
  IV U13842 ( .A(n13546), .Z(n13545) );
  NOR U13843 ( .A(n13547), .B(n13545), .Z(n13552) );
  XOR U13844 ( .A(n13547), .B(n13546), .Z(n14024) );
  XOR U13845 ( .A(n13549), .B(n13548), .Z(n14025) );
  IV U13846 ( .A(n14025), .Z(n13550) );
  NOR U13847 ( .A(n14024), .B(n13550), .Z(n13551) );
  NOR U13848 ( .A(n13552), .B(n13551), .Z(n14020) );
  XOR U13849 ( .A(n13554), .B(n13553), .Z(n14021) );
  NOR U13850 ( .A(n14020), .B(n14021), .Z(n13555) );
  NOR U13851 ( .A(n13556), .B(n13555), .Z(n14016) );
  XOR U13852 ( .A(n13558), .B(n13557), .Z(n14017) );
  NOR U13853 ( .A(n14016), .B(n14017), .Z(n13559) );
  NOR U13854 ( .A(n13560), .B(n13559), .Z(n14012) );
  XOR U13855 ( .A(n13562), .B(n13561), .Z(n14013) );
  NOR U13856 ( .A(n14012), .B(n14013), .Z(n13563) );
  NOR U13857 ( .A(n13564), .B(n13563), .Z(n14008) );
  XOR U13858 ( .A(n13566), .B(n13565), .Z(n14009) );
  NOR U13859 ( .A(n14008), .B(n14009), .Z(n13567) );
  NOR U13860 ( .A(n13568), .B(n13567), .Z(n14004) );
  XOR U13861 ( .A(n13570), .B(n13569), .Z(n14005) );
  NOR U13862 ( .A(n14004), .B(n14005), .Z(n13571) );
  NOR U13863 ( .A(n13572), .B(n13571), .Z(n14000) );
  XOR U13864 ( .A(n13574), .B(n13573), .Z(n14001) );
  NOR U13865 ( .A(n14000), .B(n14001), .Z(n13575) );
  NOR U13866 ( .A(n13576), .B(n13575), .Z(n13996) );
  XOR U13867 ( .A(n13578), .B(n13577), .Z(n13997) );
  NOR U13868 ( .A(n13996), .B(n13997), .Z(n13579) );
  NOR U13869 ( .A(n13580), .B(n13579), .Z(n13995) );
  XOR U13870 ( .A(n13582), .B(n13581), .Z(n13994) );
  NOR U13871 ( .A(n13995), .B(n13994), .Z(n13583) );
  NOR U13872 ( .A(n13584), .B(n13583), .Z(n13990) );
  XOR U13873 ( .A(n13586), .B(n13585), .Z(n13991) );
  NOR U13874 ( .A(n13990), .B(n13991), .Z(n13587) );
  NOR U13875 ( .A(n13588), .B(n13587), .Z(n13989) );
  XOR U13876 ( .A(n13590), .B(n13589), .Z(n13988) );
  NOR U13877 ( .A(n13989), .B(n13988), .Z(n13591) );
  NOR U13878 ( .A(n13592), .B(n13591), .Z(n13982) );
  XOR U13879 ( .A(n13594), .B(n13593), .Z(n13983) );
  NOR U13880 ( .A(n13982), .B(n13983), .Z(n13595) );
  NOR U13881 ( .A(n13596), .B(n13595), .Z(n13978) );
  XOR U13882 ( .A(n13598), .B(n13597), .Z(n13979) );
  NOR U13883 ( .A(n13978), .B(n13979), .Z(n13599) );
  NOR U13884 ( .A(n13600), .B(n13599), .Z(n13601) );
  IV U13885 ( .A(n13601), .Z(n13976) );
  XOR U13886 ( .A(n13603), .B(n13602), .Z(n13604) );
  IV U13887 ( .A(n13604), .Z(n13975) );
  NOR U13888 ( .A(n13976), .B(n13975), .Z(n13605) );
  NOR U13889 ( .A(n13606), .B(n13605), .Z(n13607) );
  IV U13890 ( .A(n13607), .Z(n13973) );
  NOR U13891 ( .A(n13974), .B(n13973), .Z(n13608) );
  NOR U13892 ( .A(n13609), .B(n13608), .Z(n13971) );
  NOR U13893 ( .A(n13611), .B(n13610), .Z(n13612) );
  NOR U13894 ( .A(n13971), .B(n13612), .Z(n13613) );
  NOR U13895 ( .A(n13614), .B(n13613), .Z(n13619) );
  NOR U13896 ( .A(n108), .B(n51), .Z(n13618) );
  IV U13897 ( .A(n13618), .Z(n13615) );
  NOR U13898 ( .A(n13619), .B(n13615), .Z(n13621) );
  XOR U13899 ( .A(n13617), .B(n13616), .Z(n13965) );
  XOR U13900 ( .A(n13619), .B(n13618), .Z(n13964) );
  NOR U13901 ( .A(n13965), .B(n13964), .Z(n13620) );
  NOR U13902 ( .A(n13621), .B(n13620), .Z(n14139) );
  XOR U13903 ( .A(n13623), .B(n13622), .Z(n14138) );
  NOR U13904 ( .A(n14139), .B(n14138), .Z(n13624) );
  NOR U13905 ( .A(n13625), .B(n13624), .Z(n13959) );
  XOR U13906 ( .A(n13627), .B(n13626), .Z(n13958) );
  NOR U13907 ( .A(n13959), .B(n13958), .Z(n13628) );
  NOR U13908 ( .A(n13629), .B(n13628), .Z(n13630) );
  IV U13909 ( .A(n13630), .Z(n13955) );
  NOR U13910 ( .A(n13956), .B(n13955), .Z(n13631) );
  NOR U13911 ( .A(n13632), .B(n13631), .Z(n13953) );
  IV U13912 ( .A(n13953), .Z(n13635) );
  XOR U13913 ( .A(n13634), .B(n13633), .Z(n13952) );
  NOR U13914 ( .A(n13635), .B(n13952), .Z(n13636) );
  NOR U13915 ( .A(n13637), .B(n13636), .Z(n14161) );
  IV U13916 ( .A(n14161), .Z(n13638) );
  NOR U13917 ( .A(n13639), .B(n13638), .Z(n13640) );
  NOR U13918 ( .A(n13641), .B(n13640), .Z(n13642) );
  IV U13919 ( .A(n13642), .Z(n13647) );
  NOR U13920 ( .A(n112), .B(n51), .Z(n13646) );
  IV U13921 ( .A(n13646), .Z(n13643) );
  NOR U13922 ( .A(n13647), .B(n13643), .Z(n13649) );
  XOR U13923 ( .A(n13645), .B(n13644), .Z(n13949) );
  XOR U13924 ( .A(n13647), .B(n13646), .Z(n13948) );
  NOR U13925 ( .A(n13949), .B(n13948), .Z(n13648) );
  NOR U13926 ( .A(n13649), .B(n13648), .Z(n13944) );
  XOR U13927 ( .A(n13651), .B(n13650), .Z(n13943) );
  NOR U13928 ( .A(n13944), .B(n13943), .Z(n13652) );
  NOR U13929 ( .A(n13653), .B(n13652), .Z(n13940) );
  XOR U13930 ( .A(n13655), .B(n13654), .Z(n13939) );
  NOR U13931 ( .A(n13940), .B(n13939), .Z(n13656) );
  NOR U13932 ( .A(n13657), .B(n13656), .Z(n14181) );
  IV U13933 ( .A(n14181), .Z(n13658) );
  NOR U13934 ( .A(n13659), .B(n13658), .Z(n13660) );
  NOR U13935 ( .A(n13661), .B(n13660), .Z(n13664) );
  IV U13936 ( .A(n13664), .Z(n13662) );
  NOR U13937 ( .A(n13663), .B(n13662), .Z(n13667) );
  XOR U13938 ( .A(n13664), .B(n13663), .Z(n13935) );
  NOR U13939 ( .A(n114), .B(n51), .Z(n13665) );
  IV U13940 ( .A(n13665), .Z(n13934) );
  NOR U13941 ( .A(n13935), .B(n13934), .Z(n13666) );
  NOR U13942 ( .A(n13667), .B(n13666), .Z(n14193) );
  XOR U13943 ( .A(n13669), .B(n13668), .Z(n14194) );
  IV U13944 ( .A(n14194), .Z(n13670) );
  NOR U13945 ( .A(n14193), .B(n13670), .Z(n13671) );
  NOR U13946 ( .A(n13672), .B(n13671), .Z(n13933) );
  XOR U13947 ( .A(n13674), .B(n13673), .Z(n13932) );
  NOR U13948 ( .A(n13933), .B(n13932), .Z(n13675) );
  NOR U13949 ( .A(n13676), .B(n13675), .Z(n13677) );
  IV U13950 ( .A(n13677), .Z(n13927) );
  NOR U13951 ( .A(n13678), .B(n13927), .Z(n13679) );
  NOR U13952 ( .A(n13680), .B(n13679), .Z(n13681) );
  IV U13953 ( .A(n13681), .Z(n13686) );
  NOR U13954 ( .A(n116), .B(n51), .Z(n13685) );
  IV U13955 ( .A(n13685), .Z(n13682) );
  NOR U13956 ( .A(n13686), .B(n13682), .Z(n13688) );
  XOR U13957 ( .A(n13684), .B(n13683), .Z(n14210) );
  XOR U13958 ( .A(n13686), .B(n13685), .Z(n14209) );
  NOR U13959 ( .A(n14210), .B(n14209), .Z(n13687) );
  NOR U13960 ( .A(n13688), .B(n13687), .Z(n13690) );
  IV U13961 ( .A(n13690), .Z(n14216) );
  NOR U13962 ( .A(n13689), .B(n14216), .Z(n13695) );
  IV U13963 ( .A(n13689), .Z(n14217) );
  NOR U13964 ( .A(n13690), .B(n14217), .Z(n13693) );
  XOR U13965 ( .A(n13692), .B(n13691), .Z(n14219) );
  NOR U13966 ( .A(n13693), .B(n14219), .Z(n13694) );
  NOR U13967 ( .A(n13695), .B(n13694), .Z(n13696) );
  IV U13968 ( .A(n13696), .Z(n13703) );
  NOR U13969 ( .A(n117), .B(n51), .Z(n13702) );
  IV U13970 ( .A(n13702), .Z(n13697) );
  NOR U13971 ( .A(n13703), .B(n13697), .Z(n13705) );
  XOR U13972 ( .A(n13699), .B(n13698), .Z(n13700) );
  XOR U13973 ( .A(n13701), .B(n13700), .Z(n13923) );
  XOR U13974 ( .A(n13703), .B(n13702), .Z(n13924) );
  NOR U13975 ( .A(n13923), .B(n13924), .Z(n13704) );
  NOR U13976 ( .A(n13705), .B(n13704), .Z(n13708) );
  XOR U13977 ( .A(n13707), .B(n13706), .Z(n13709) );
  NOR U13978 ( .A(n13708), .B(n13709), .Z(n13713) );
  IV U13979 ( .A(n13708), .Z(n14233) );
  IV U13980 ( .A(n13709), .Z(n14232) );
  NOR U13981 ( .A(n14233), .B(n14232), .Z(n13711) );
  NOR U13982 ( .A(n79), .B(n51), .Z(n14235) );
  IV U13983 ( .A(n14235), .Z(n13710) );
  NOR U13984 ( .A(n13711), .B(n13710), .Z(n13712) );
  NOR U13985 ( .A(n13713), .B(n13712), .Z(n13715) );
  IV U13986 ( .A(n13715), .Z(n14241) );
  NOR U13987 ( .A(n13714), .B(n14241), .Z(n13722) );
  IV U13988 ( .A(n13714), .Z(n14242) );
  NOR U13989 ( .A(n13715), .B(n14242), .Z(n13720) );
  XOR U13990 ( .A(n13717), .B(n13716), .Z(n13718) );
  XOR U13991 ( .A(n13719), .B(n13718), .Z(n14244) );
  NOR U13992 ( .A(n13720), .B(n14244), .Z(n13721) );
  NOR U13993 ( .A(n13722), .B(n13721), .Z(n13730) );
  IV U13994 ( .A(n13730), .Z(n13724) );
  NOR U13995 ( .A(n120), .B(n51), .Z(n13723) );
  IV U13996 ( .A(n13723), .Z(n13729) );
  NOR U13997 ( .A(n13724), .B(n13729), .Z(n13732) );
  XOR U13998 ( .A(n13726), .B(n13725), .Z(n13727) );
  XOR U13999 ( .A(n13728), .B(n13727), .Z(n14249) );
  XOR U14000 ( .A(n13730), .B(n13729), .Z(n14250) );
  NOR U14001 ( .A(n14249), .B(n14250), .Z(n13731) );
  NOR U14002 ( .A(n13732), .B(n13731), .Z(n13737) );
  XOR U14003 ( .A(n13734), .B(n13733), .Z(n13736) );
  IV U14004 ( .A(n13736), .Z(n13735) );
  NOR U14005 ( .A(n13737), .B(n13735), .Z(n13740) );
  XOR U14006 ( .A(n13737), .B(n13736), .Z(n13920) );
  NOR U14007 ( .A(n123), .B(n51), .Z(n13921) );
  IV U14008 ( .A(n13921), .Z(n13738) );
  NOR U14009 ( .A(n13920), .B(n13738), .Z(n13739) );
  NOR U14010 ( .A(n13740), .B(n13739), .Z(n13743) );
  XOR U14011 ( .A(n13742), .B(n13741), .Z(n13744) );
  IV U14012 ( .A(n13744), .Z(n14262) );
  NOR U14013 ( .A(n13743), .B(n14262), .Z(n13748) );
  IV U14014 ( .A(n13743), .Z(n14263) );
  NOR U14015 ( .A(n13744), .B(n14263), .Z(n13746) );
  NOR U14016 ( .A(n125), .B(n51), .Z(n14265) );
  IV U14017 ( .A(n14265), .Z(n13745) );
  NOR U14018 ( .A(n13746), .B(n13745), .Z(n13747) );
  NOR U14019 ( .A(n13748), .B(n13747), .Z(n13753) );
  NOR U14020 ( .A(n126), .B(n51), .Z(n13752) );
  IV U14021 ( .A(n13752), .Z(n13749) );
  NOR U14022 ( .A(n13753), .B(n13749), .Z(n13756) );
  XOR U14023 ( .A(n13751), .B(n13750), .Z(n14271) );
  IV U14024 ( .A(n14271), .Z(n13754) );
  XOR U14025 ( .A(n13753), .B(n13752), .Z(n14270) );
  NOR U14026 ( .A(n13754), .B(n14270), .Z(n13755) );
  NOR U14027 ( .A(n13756), .B(n13755), .Z(n13761) );
  XOR U14028 ( .A(n13758), .B(n13757), .Z(n13760) );
  IV U14029 ( .A(n13760), .Z(n13759) );
  NOR U14030 ( .A(n13761), .B(n13759), .Z(n13764) );
  XOR U14031 ( .A(n13761), .B(n13760), .Z(n14281) );
  NOR U14032 ( .A(n128), .B(n51), .Z(n14282) );
  IV U14033 ( .A(n14282), .Z(n13762) );
  NOR U14034 ( .A(n14281), .B(n13762), .Z(n13763) );
  NOR U14035 ( .A(n13764), .B(n13763), .Z(n14289) );
  XOR U14036 ( .A(n13766), .B(n13765), .Z(n14288) );
  NOR U14037 ( .A(n14289), .B(n14288), .Z(n13767) );
  NOR U14038 ( .A(n13768), .B(n13767), .Z(n13771) );
  NOR U14039 ( .A(n133), .B(n51), .Z(n13770) );
  IV U14040 ( .A(n13770), .Z(n13769) );
  NOR U14041 ( .A(n13771), .B(n13769), .Z(n13776) );
  XOR U14042 ( .A(n13771), .B(n13770), .Z(n14293) );
  XOR U14043 ( .A(n13773), .B(n13772), .Z(n14294) );
  IV U14044 ( .A(n14294), .Z(n13774) );
  NOR U14045 ( .A(n14293), .B(n13774), .Z(n13775) );
  NOR U14046 ( .A(n13776), .B(n13775), .Z(n13780) );
  XOR U14047 ( .A(n13778), .B(n13777), .Z(n13779) );
  NOR U14048 ( .A(n13780), .B(n13779), .Z(n13784) );
  XOR U14049 ( .A(n13780), .B(n13779), .Z(n13781) );
  IV U14050 ( .A(n13781), .Z(n14304) );
  NOR U14051 ( .A(n135), .B(n51), .Z(n14305) );
  IV U14052 ( .A(n14305), .Z(n13782) );
  NOR U14053 ( .A(n14304), .B(n13782), .Z(n13783) );
  NOR U14054 ( .A(n13784), .B(n13783), .Z(n13787) );
  NOR U14055 ( .A(n137), .B(n51), .Z(n13786) );
  IV U14056 ( .A(n13786), .Z(n13785) );
  NOR U14057 ( .A(n13787), .B(n13785), .Z(n13791) );
  XOR U14058 ( .A(n13787), .B(n13786), .Z(n14311) );
  XOR U14059 ( .A(n13789), .B(n13788), .Z(n14312) );
  NOR U14060 ( .A(n14311), .B(n14312), .Z(n13790) );
  NOR U14061 ( .A(n13791), .B(n13790), .Z(n13794) );
  NOR U14062 ( .A(n139), .B(n51), .Z(n13793) );
  IV U14063 ( .A(n13793), .Z(n13792) );
  NOR U14064 ( .A(n13794), .B(n13792), .Z(n13799) );
  XOR U14065 ( .A(n13794), .B(n13793), .Z(n14316) );
  XOR U14066 ( .A(n13796), .B(n13795), .Z(n14317) );
  IV U14067 ( .A(n14317), .Z(n13797) );
  NOR U14068 ( .A(n14316), .B(n13797), .Z(n13798) );
  NOR U14069 ( .A(n13799), .B(n13798), .Z(n13803) );
  XOR U14070 ( .A(n13801), .B(n13800), .Z(n13802) );
  NOR U14071 ( .A(n13803), .B(n13802), .Z(n13807) );
  XOR U14072 ( .A(n13803), .B(n13802), .Z(n13804) );
  IV U14073 ( .A(n13804), .Z(n14327) );
  NOR U14074 ( .A(n141), .B(n51), .Z(n14328) );
  IV U14075 ( .A(n14328), .Z(n13805) );
  NOR U14076 ( .A(n14327), .B(n13805), .Z(n13806) );
  NOR U14077 ( .A(n13807), .B(n13806), .Z(n13810) );
  NOR U14078 ( .A(n143), .B(n51), .Z(n13809) );
  IV U14079 ( .A(n13809), .Z(n13808) );
  NOR U14080 ( .A(n13810), .B(n13808), .Z(n13814) );
  XOR U14081 ( .A(n13810), .B(n13809), .Z(n14334) );
  XOR U14082 ( .A(n13812), .B(n13811), .Z(n14335) );
  NOR U14083 ( .A(n14334), .B(n14335), .Z(n13813) );
  NOR U14084 ( .A(n13814), .B(n13813), .Z(n13819) );
  NOR U14085 ( .A(n145), .B(n51), .Z(n13818) );
  IV U14086 ( .A(n13818), .Z(n13815) );
  NOR U14087 ( .A(n13819), .B(n13815), .Z(n13822) );
  XOR U14088 ( .A(n13817), .B(n13816), .Z(n14340) );
  IV U14089 ( .A(n14340), .Z(n13820) );
  XOR U14090 ( .A(n13819), .B(n13818), .Z(n14339) );
  NOR U14091 ( .A(n13820), .B(n14339), .Z(n13821) );
  NOR U14092 ( .A(n13822), .B(n13821), .Z(n13827) );
  XOR U14093 ( .A(n13824), .B(n13823), .Z(n13826) );
  IV U14094 ( .A(n13826), .Z(n13825) );
  NOR U14095 ( .A(n13827), .B(n13825), .Z(n13830) );
  XOR U14096 ( .A(n13827), .B(n13826), .Z(n14349) );
  NOR U14097 ( .A(n147), .B(n51), .Z(n13828) );
  IV U14098 ( .A(n13828), .Z(n14348) );
  NOR U14099 ( .A(n14349), .B(n14348), .Z(n13829) );
  NOR U14100 ( .A(n13830), .B(n13829), .Z(n13833) );
  XOR U14101 ( .A(n13832), .B(n13831), .Z(n13834) );
  NOR U14102 ( .A(n13833), .B(n13834), .Z(n13838) );
  IV U14103 ( .A(n13833), .Z(n13835) );
  XOR U14104 ( .A(n13835), .B(n13834), .Z(n14358) );
  NOR U14105 ( .A(n148), .B(n51), .Z(n14359) );
  IV U14106 ( .A(n14359), .Z(n13836) );
  NOR U14107 ( .A(n14358), .B(n13836), .Z(n13837) );
  NOR U14108 ( .A(n13838), .B(n13837), .Z(n13841) );
  NOR U14109 ( .A(n150), .B(n51), .Z(n13840) );
  IV U14110 ( .A(n13840), .Z(n13839) );
  NOR U14111 ( .A(n13841), .B(n13839), .Z(n13846) );
  XOR U14112 ( .A(n13841), .B(n13840), .Z(n14362) );
  XOR U14113 ( .A(n13843), .B(n13842), .Z(n14363) );
  IV U14114 ( .A(n14363), .Z(n13844) );
  NOR U14115 ( .A(n14362), .B(n13844), .Z(n13845) );
  NOR U14116 ( .A(n13846), .B(n13845), .Z(n13848) );
  IV U14117 ( .A(n13848), .Z(n13847) );
  NOR U14118 ( .A(n13849), .B(n13847), .Z(n13851) );
  NOR U14119 ( .A(n153), .B(n51), .Z(n13918) );
  XOR U14120 ( .A(n13849), .B(n13848), .Z(n13917) );
  NOR U14121 ( .A(n13918), .B(n13917), .Z(n13850) );
  NOR U14122 ( .A(n13851), .B(n13850), .Z(n13854) );
  XOR U14123 ( .A(n13853), .B(n13852), .Z(n13855) );
  NOR U14124 ( .A(n13854), .B(n13855), .Z(n13858) );
  NOR U14125 ( .A(n155), .B(n51), .Z(n14376) );
  IV U14126 ( .A(n13854), .Z(n13856) );
  XOR U14127 ( .A(n13856), .B(n13855), .Z(n14375) );
  NOR U14128 ( .A(n14376), .B(n14375), .Z(n13857) );
  NOR U14129 ( .A(n13858), .B(n13857), .Z(n13864) );
  IV U14130 ( .A(n13864), .Z(n13860) );
  NOR U14131 ( .A(n156), .B(n51), .Z(n13859) );
  IV U14132 ( .A(n13859), .Z(n13863) );
  NOR U14133 ( .A(n13860), .B(n13863), .Z(n13866) );
  XOR U14134 ( .A(n13862), .B(n13861), .Z(n14382) );
  XOR U14135 ( .A(n13864), .B(n13863), .Z(n14381) );
  NOR U14136 ( .A(n14382), .B(n14381), .Z(n13865) );
  NOR U14137 ( .A(n13866), .B(n13865), .Z(n13869) );
  XOR U14138 ( .A(n13868), .B(n13867), .Z(n13870) );
  NOR U14139 ( .A(n13869), .B(n13870), .Z(n13874) );
  IV U14140 ( .A(n13869), .Z(n13871) );
  XOR U14141 ( .A(n13871), .B(n13870), .Z(n13914) );
  NOR U14142 ( .A(n158), .B(n51), .Z(n13915) );
  IV U14143 ( .A(n13915), .Z(n13872) );
  NOR U14144 ( .A(n13914), .B(n13872), .Z(n13873) );
  NOR U14145 ( .A(n13874), .B(n13873), .Z(n13877) );
  NOR U14146 ( .A(n161), .B(n51), .Z(n13876) );
  IV U14147 ( .A(n13876), .Z(n13875) );
  NOR U14148 ( .A(n13877), .B(n13875), .Z(n13881) );
  XOR U14149 ( .A(n13877), .B(n13876), .Z(n14394) );
  XOR U14150 ( .A(n13879), .B(n13878), .Z(n14395) );
  NOR U14151 ( .A(n14394), .B(n14395), .Z(n13880) );
  NOR U14152 ( .A(n13881), .B(n13880), .Z(n13886) );
  NOR U14153 ( .A(n163), .B(n51), .Z(n13885) );
  IV U14154 ( .A(n13885), .Z(n13882) );
  NOR U14155 ( .A(n13886), .B(n13882), .Z(n13889) );
  XOR U14156 ( .A(n13884), .B(n13883), .Z(n14402) );
  IV U14157 ( .A(n14402), .Z(n13887) );
  XOR U14158 ( .A(n13886), .B(n13885), .Z(n14401) );
  NOR U14159 ( .A(n13887), .B(n14401), .Z(n13888) );
  NOR U14160 ( .A(n13889), .B(n13888), .Z(n13893) );
  XOR U14161 ( .A(n13891), .B(n13890), .Z(n13892) );
  NOR U14162 ( .A(n13893), .B(n13892), .Z(n13897) );
  XOR U14163 ( .A(n13893), .B(n13892), .Z(n13894) );
  IV U14164 ( .A(n13894), .Z(n14412) );
  NOR U14165 ( .A(n165), .B(n51), .Z(n13895) );
  IV U14166 ( .A(n13895), .Z(n14413) );
  NOR U14167 ( .A(n14412), .B(n14413), .Z(n13896) );
  NOR U14168 ( .A(n13897), .B(n13896), .Z(n13900) );
  NOR U14169 ( .A(n167), .B(n51), .Z(n13899) );
  IV U14170 ( .A(n13899), .Z(n13898) );
  NOR U14171 ( .A(n13900), .B(n13898), .Z(n13905) );
  XOR U14172 ( .A(n13900), .B(n13899), .Z(n14417) );
  XOR U14173 ( .A(n13902), .B(n13901), .Z(n14418) );
  IV U14174 ( .A(n14418), .Z(n13903) );
  NOR U14175 ( .A(n14417), .B(n13903), .Z(n13904) );
  NOR U14176 ( .A(n13905), .B(n13904), .Z(n13913) );
  XOR U14177 ( .A(n13907), .B(n13906), .Z(n13912) );
  NOR U14178 ( .A(n13913), .B(n13912), .Z(n13910) );
  XOR U14179 ( .A(n13909), .B(n13908), .Z(n13911) );
  NOR U14180 ( .A(n13910), .B(n13911), .Z(n28612) );
  IV U14181 ( .A(n13910), .Z(n31649) );
  XOR U14182 ( .A(n31649), .B(n13911), .Z(n31646) );
  XOR U14183 ( .A(n13913), .B(n13912), .Z(n28601) );
  IV U14184 ( .A(n28601), .Z(n31645) );
  XOR U14185 ( .A(n13915), .B(n13914), .Z(n14389) );
  NOR U14186 ( .A(n161), .B(n52), .Z(n14390) );
  IV U14187 ( .A(n14390), .Z(n13916) );
  NOR U14188 ( .A(n14389), .B(n13916), .Z(n14392) );
  XOR U14189 ( .A(n13918), .B(n13917), .Z(n14371) );
  NOR U14190 ( .A(n155), .B(n52), .Z(n14370) );
  IV U14191 ( .A(n14370), .Z(n13919) );
  NOR U14192 ( .A(n14371), .B(n13919), .Z(n14373) );
  NOR U14193 ( .A(n148), .B(n52), .Z(n14846) );
  XOR U14194 ( .A(n13921), .B(n13920), .Z(n14257) );
  NOR U14195 ( .A(n125), .B(n52), .Z(n14258) );
  IV U14196 ( .A(n14258), .Z(n13922) );
  NOR U14197 ( .A(n14257), .B(n13922), .Z(n14260) );
  NOR U14198 ( .A(n119), .B(n52), .Z(n14230) );
  XOR U14199 ( .A(n13924), .B(n13923), .Z(n13925) );
  IV U14200 ( .A(n13925), .Z(n14226) );
  NOR U14201 ( .A(n79), .B(n52), .Z(n14227) );
  IV U14202 ( .A(n14227), .Z(n13926) );
  NOR U14203 ( .A(n14226), .B(n13926), .Z(n14229) );
  NOR U14204 ( .A(n80), .B(n52), .Z(n14212) );
  IV U14205 ( .A(n14212), .Z(n14208) );
  NOR U14206 ( .A(n116), .B(n52), .Z(n14203) );
  XOR U14207 ( .A(n13928), .B(n13927), .Z(n13929) );
  XOR U14208 ( .A(n13930), .B(n13929), .Z(n14204) );
  IV U14209 ( .A(n14204), .Z(n13931) );
  NOR U14210 ( .A(n14203), .B(n13931), .Z(n14206) );
  NOR U14211 ( .A(n81), .B(n52), .Z(n14199) );
  XOR U14212 ( .A(n13933), .B(n13932), .Z(n14198) );
  NOR U14213 ( .A(n14199), .B(n14198), .Z(n14202) );
  XOR U14214 ( .A(n13935), .B(n13934), .Z(n13936) );
  NOR U14215 ( .A(n82), .B(n52), .Z(n13937) );
  NOR U14216 ( .A(n13936), .B(n13937), .Z(n14188) );
  XOR U14217 ( .A(n13937), .B(n13936), .Z(n13938) );
  IV U14218 ( .A(n13938), .Z(n14698) );
  XOR U14219 ( .A(n13940), .B(n13939), .Z(n13941) );
  NOR U14220 ( .A(n83), .B(n52), .Z(n14452) );
  NOR U14221 ( .A(n13941), .B(n14452), .Z(n14175) );
  IV U14222 ( .A(n13941), .Z(n14454) );
  IV U14223 ( .A(n14452), .Z(n13942) );
  NOR U14224 ( .A(n14454), .B(n13942), .Z(n14173) );
  XOR U14225 ( .A(n13944), .B(n13943), .Z(n13945) );
  NOR U14226 ( .A(n113), .B(n52), .Z(n13946) );
  NOR U14227 ( .A(n13945), .B(n13946), .Z(n14172) );
  XOR U14228 ( .A(n13946), .B(n13945), .Z(n13947) );
  IV U14229 ( .A(n13947), .Z(n14457) );
  XOR U14230 ( .A(n13949), .B(n13948), .Z(n13950) );
  IV U14231 ( .A(n13950), .Z(n14166) );
  NOR U14232 ( .A(n84), .B(n52), .Z(n14167) );
  IV U14233 ( .A(n14167), .Z(n13951) );
  NOR U14234 ( .A(n14166), .B(n13951), .Z(n14169) );
  NOR U14235 ( .A(n85), .B(n52), .Z(n14154) );
  IV U14236 ( .A(n14154), .Z(n13954) );
  XOR U14237 ( .A(n13953), .B(n13952), .Z(n14153) );
  NOR U14238 ( .A(n13954), .B(n14153), .Z(n14156) );
  XOR U14239 ( .A(n13956), .B(n13955), .Z(n14150) );
  NOR U14240 ( .A(n111), .B(n52), .Z(n14149) );
  IV U14241 ( .A(n14149), .Z(n13957) );
  NOR U14242 ( .A(n14150), .B(n13957), .Z(n14152) );
  NOR U14243 ( .A(n86), .B(n52), .Z(n13961) );
  XOR U14244 ( .A(n13959), .B(n13958), .Z(n13960) );
  NOR U14245 ( .A(n13961), .B(n13960), .Z(n14147) );
  XOR U14246 ( .A(n13961), .B(n13960), .Z(n13962) );
  IV U14247 ( .A(n13962), .Z(n14471) );
  NOR U14248 ( .A(n110), .B(n52), .Z(n13963) );
  IV U14249 ( .A(n13963), .Z(n14141) );
  XOR U14250 ( .A(n13965), .B(n13964), .Z(n13966) );
  NOR U14251 ( .A(n109), .B(n52), .Z(n13967) );
  NOR U14252 ( .A(n13966), .B(n13967), .Z(n14136) );
  IV U14253 ( .A(n13966), .Z(n14477) );
  IV U14254 ( .A(n13967), .Z(n14476) );
  NOR U14255 ( .A(n14477), .B(n14476), .Z(n14134) );
  XOR U14256 ( .A(n13969), .B(n13968), .Z(n13970) );
  XOR U14257 ( .A(n13971), .B(n13970), .Z(n14129) );
  NOR U14258 ( .A(n108), .B(n52), .Z(n14128) );
  IV U14259 ( .A(n14128), .Z(n13972) );
  NOR U14260 ( .A(n14129), .B(n13972), .Z(n14132) );
  NOR U14261 ( .A(n87), .B(n52), .Z(n14124) );
  XOR U14262 ( .A(n13974), .B(n13973), .Z(n14123) );
  NOR U14263 ( .A(n14124), .B(n14123), .Z(n14127) );
  XOR U14264 ( .A(n13976), .B(n13975), .Z(n14119) );
  NOR U14265 ( .A(n107), .B(n52), .Z(n14118) );
  IV U14266 ( .A(n14118), .Z(n13977) );
  NOR U14267 ( .A(n14119), .B(n13977), .Z(n14121) );
  IV U14268 ( .A(n13978), .Z(n13980) );
  XOR U14269 ( .A(n13980), .B(n13979), .Z(n14114) );
  NOR U14270 ( .A(n88), .B(n52), .Z(n14115) );
  IV U14271 ( .A(n14115), .Z(n13981) );
  NOR U14272 ( .A(n14114), .B(n13981), .Z(n14117) );
  IV U14273 ( .A(n13982), .Z(n13984) );
  XOR U14274 ( .A(n13984), .B(n13983), .Z(n13986) );
  NOR U14275 ( .A(n106), .B(n52), .Z(n13987) );
  IV U14276 ( .A(n13987), .Z(n13985) );
  NOR U14277 ( .A(n13986), .B(n13985), .Z(n14113) );
  XOR U14278 ( .A(n13987), .B(n13986), .Z(n14493) );
  NOR U14279 ( .A(n105), .B(n52), .Z(n14107) );
  XOR U14280 ( .A(n13989), .B(n13988), .Z(n14106) );
  NOR U14281 ( .A(n14107), .B(n14106), .Z(n14110) );
  IV U14282 ( .A(n13990), .Z(n13992) );
  XOR U14283 ( .A(n13992), .B(n13991), .Z(n14100) );
  NOR U14284 ( .A(n104), .B(n52), .Z(n14101) );
  IV U14285 ( .A(n14101), .Z(n13993) );
  NOR U14286 ( .A(n14100), .B(n13993), .Z(n14104) );
  NOR U14287 ( .A(n89), .B(n52), .Z(n14096) );
  XOR U14288 ( .A(n13995), .B(n13994), .Z(n14095) );
  NOR U14289 ( .A(n14096), .B(n14095), .Z(n14099) );
  IV U14290 ( .A(n13996), .Z(n13998) );
  XOR U14291 ( .A(n13998), .B(n13997), .Z(n14090) );
  NOR U14292 ( .A(n103), .B(n52), .Z(n14091) );
  IV U14293 ( .A(n14091), .Z(n13999) );
  NOR U14294 ( .A(n14090), .B(n13999), .Z(n14093) );
  IV U14295 ( .A(n14000), .Z(n14002) );
  XOR U14296 ( .A(n14002), .B(n14001), .Z(n14086) );
  NOR U14297 ( .A(n90), .B(n52), .Z(n14087) );
  IV U14298 ( .A(n14087), .Z(n14003) );
  NOR U14299 ( .A(n14086), .B(n14003), .Z(n14089) );
  IV U14300 ( .A(n14004), .Z(n14006) );
  XOR U14301 ( .A(n14006), .B(n14005), .Z(n14082) );
  NOR U14302 ( .A(n102), .B(n52), .Z(n14083) );
  IV U14303 ( .A(n14083), .Z(n14007) );
  NOR U14304 ( .A(n14082), .B(n14007), .Z(n14085) );
  IV U14305 ( .A(n14008), .Z(n14010) );
  XOR U14306 ( .A(n14010), .B(n14009), .Z(n14078) );
  NOR U14307 ( .A(n101), .B(n52), .Z(n14079) );
  IV U14308 ( .A(n14079), .Z(n14011) );
  NOR U14309 ( .A(n14078), .B(n14011), .Z(n14081) );
  IV U14310 ( .A(n14012), .Z(n14014) );
  XOR U14311 ( .A(n14014), .B(n14013), .Z(n14074) );
  NOR U14312 ( .A(n100), .B(n52), .Z(n14075) );
  IV U14313 ( .A(n14075), .Z(n14015) );
  NOR U14314 ( .A(n14074), .B(n14015), .Z(n14077) );
  IV U14315 ( .A(n14016), .Z(n14018) );
  XOR U14316 ( .A(n14018), .B(n14017), .Z(n14070) );
  NOR U14317 ( .A(n99), .B(n52), .Z(n14071) );
  IV U14318 ( .A(n14071), .Z(n14019) );
  NOR U14319 ( .A(n14070), .B(n14019), .Z(n14073) );
  IV U14320 ( .A(n14020), .Z(n14022) );
  XOR U14321 ( .A(n14022), .B(n14021), .Z(n14066) );
  NOR U14322 ( .A(n98), .B(n52), .Z(n14067) );
  IV U14323 ( .A(n14067), .Z(n14023) );
  NOR U14324 ( .A(n14066), .B(n14023), .Z(n14069) );
  XOR U14325 ( .A(n14025), .B(n14024), .Z(n14062) );
  NOR U14326 ( .A(n91), .B(n52), .Z(n14063) );
  IV U14327 ( .A(n14063), .Z(n14026) );
  NOR U14328 ( .A(n14062), .B(n14026), .Z(n14065) );
  XOR U14329 ( .A(n14028), .B(n14027), .Z(n14050) );
  IV U14330 ( .A(n14050), .Z(n14030) );
  NOR U14331 ( .A(n96), .B(n52), .Z(n14029) );
  IV U14332 ( .A(n14029), .Z(n14051) );
  NOR U14333 ( .A(n14030), .B(n14051), .Z(n14053) );
  NOR U14334 ( .A(n95), .B(n52), .Z(n14047) );
  IV U14335 ( .A(n14047), .Z(n14033) );
  XOR U14336 ( .A(n14032), .B(n14031), .Z(n14046) );
  NOR U14337 ( .A(n14033), .B(n14046), .Z(n14049) );
  NOR U14338 ( .A(n93), .B(n52), .Z(n15033) );
  IV U14339 ( .A(n15033), .Z(n14034) );
  NOR U14340 ( .A(n51), .B(n168), .Z(n14042) );
  IV U14341 ( .A(n14042), .Z(n14037) );
  NOR U14342 ( .A(n14034), .B(n14037), .Z(n14035) );
  IV U14343 ( .A(n14035), .Z(n14036) );
  NOR U14344 ( .A(n94), .B(n14036), .Z(n14045) );
  NOR U14345 ( .A(n14037), .B(n93), .Z(n14038) );
  XOR U14346 ( .A(n94), .B(n14038), .Z(n14039) );
  NOR U14347 ( .A(n52), .B(n14039), .Z(n14040) );
  IV U14348 ( .A(n14040), .Z(n14543) );
  XOR U14349 ( .A(n14042), .B(n14041), .Z(n14542) );
  IV U14350 ( .A(n14542), .Z(n14043) );
  NOR U14351 ( .A(n14543), .B(n14043), .Z(n14044) );
  NOR U14352 ( .A(n14045), .B(n14044), .Z(n14539) );
  XOR U14353 ( .A(n14047), .B(n14046), .Z(n14538) );
  NOR U14354 ( .A(n14539), .B(n14538), .Z(n14048) );
  NOR U14355 ( .A(n14049), .B(n14048), .Z(n14566) );
  XOR U14356 ( .A(n14051), .B(n14050), .Z(n14565) );
  NOR U14357 ( .A(n14566), .B(n14565), .Z(n14052) );
  NOR U14358 ( .A(n14053), .B(n14052), .Z(n14058) );
  XOR U14359 ( .A(n14055), .B(n14054), .Z(n14057) );
  IV U14360 ( .A(n14057), .Z(n14056) );
  NOR U14361 ( .A(n14058), .B(n14056), .Z(n14061) );
  XOR U14362 ( .A(n14058), .B(n14057), .Z(n14535) );
  NOR U14363 ( .A(n97), .B(n52), .Z(n14536) );
  IV U14364 ( .A(n14536), .Z(n14059) );
  NOR U14365 ( .A(n14535), .B(n14059), .Z(n14060) );
  NOR U14366 ( .A(n14061), .B(n14060), .Z(n14531) );
  XOR U14367 ( .A(n14063), .B(n14062), .Z(n14532) );
  NOR U14368 ( .A(n14531), .B(n14532), .Z(n14064) );
  NOR U14369 ( .A(n14065), .B(n14064), .Z(n14527) );
  XOR U14370 ( .A(n14067), .B(n14066), .Z(n14528) );
  NOR U14371 ( .A(n14527), .B(n14528), .Z(n14068) );
  NOR U14372 ( .A(n14069), .B(n14068), .Z(n14523) );
  XOR U14373 ( .A(n14071), .B(n14070), .Z(n14524) );
  NOR U14374 ( .A(n14523), .B(n14524), .Z(n14072) );
  NOR U14375 ( .A(n14073), .B(n14072), .Z(n14519) );
  XOR U14376 ( .A(n14075), .B(n14074), .Z(n14520) );
  NOR U14377 ( .A(n14519), .B(n14520), .Z(n14076) );
  NOR U14378 ( .A(n14077), .B(n14076), .Z(n14515) );
  XOR U14379 ( .A(n14079), .B(n14078), .Z(n14516) );
  NOR U14380 ( .A(n14515), .B(n14516), .Z(n14080) );
  NOR U14381 ( .A(n14081), .B(n14080), .Z(n14511) );
  XOR U14382 ( .A(n14083), .B(n14082), .Z(n14512) );
  NOR U14383 ( .A(n14511), .B(n14512), .Z(n14084) );
  NOR U14384 ( .A(n14085), .B(n14084), .Z(n14507) );
  XOR U14385 ( .A(n14087), .B(n14086), .Z(n14508) );
  NOR U14386 ( .A(n14507), .B(n14508), .Z(n14088) );
  NOR U14387 ( .A(n14089), .B(n14088), .Z(n14503) );
  XOR U14388 ( .A(n14091), .B(n14090), .Z(n14504) );
  NOR U14389 ( .A(n14503), .B(n14504), .Z(n14092) );
  NOR U14390 ( .A(n14093), .B(n14092), .Z(n14094) );
  IV U14391 ( .A(n14094), .Z(n14501) );
  XOR U14392 ( .A(n14096), .B(n14095), .Z(n14097) );
  IV U14393 ( .A(n14097), .Z(n14500) );
  NOR U14394 ( .A(n14501), .B(n14500), .Z(n14098) );
  NOR U14395 ( .A(n14099), .B(n14098), .Z(n14498) );
  IV U14396 ( .A(n14498), .Z(n14102) );
  XOR U14397 ( .A(n14101), .B(n14100), .Z(n14497) );
  NOR U14398 ( .A(n14102), .B(n14497), .Z(n14103) );
  NOR U14399 ( .A(n14104), .B(n14103), .Z(n14105) );
  IV U14400 ( .A(n14105), .Z(n14495) );
  XOR U14401 ( .A(n14107), .B(n14106), .Z(n14108) );
  IV U14402 ( .A(n14108), .Z(n14494) );
  NOR U14403 ( .A(n14495), .B(n14494), .Z(n14109) );
  NOR U14404 ( .A(n14110), .B(n14109), .Z(n14111) );
  IV U14405 ( .A(n14111), .Z(n14492) );
  NOR U14406 ( .A(n14493), .B(n14492), .Z(n14112) );
  NOR U14407 ( .A(n14113), .B(n14112), .Z(n14489) );
  XOR U14408 ( .A(n14115), .B(n14114), .Z(n14488) );
  NOR U14409 ( .A(n14489), .B(n14488), .Z(n14116) );
  NOR U14410 ( .A(n14117), .B(n14116), .Z(n14485) );
  XOR U14411 ( .A(n14119), .B(n14118), .Z(n14484) );
  NOR U14412 ( .A(n14485), .B(n14484), .Z(n14120) );
  NOR U14413 ( .A(n14121), .B(n14120), .Z(n14122) );
  IV U14414 ( .A(n14122), .Z(n14639) );
  XOR U14415 ( .A(n14124), .B(n14123), .Z(n14125) );
  IV U14416 ( .A(n14125), .Z(n14638) );
  NOR U14417 ( .A(n14639), .B(n14638), .Z(n14126) );
  NOR U14418 ( .A(n14127), .B(n14126), .Z(n14482) );
  IV U14419 ( .A(n14482), .Z(n14130) );
  XOR U14420 ( .A(n14129), .B(n14128), .Z(n14481) );
  NOR U14421 ( .A(n14130), .B(n14481), .Z(n14131) );
  NOR U14422 ( .A(n14132), .B(n14131), .Z(n14479) );
  IV U14423 ( .A(n14479), .Z(n14133) );
  NOR U14424 ( .A(n14134), .B(n14133), .Z(n14135) );
  NOR U14425 ( .A(n14136), .B(n14135), .Z(n14140) );
  IV U14426 ( .A(n14140), .Z(n14137) );
  NOR U14427 ( .A(n14141), .B(n14137), .Z(n14144) );
  XOR U14428 ( .A(n14139), .B(n14138), .Z(n14473) );
  IV U14429 ( .A(n14473), .Z(n14142) );
  XOR U14430 ( .A(n14141), .B(n14140), .Z(n14474) );
  NOR U14431 ( .A(n14142), .B(n14474), .Z(n14143) );
  NOR U14432 ( .A(n14144), .B(n14143), .Z(n14145) );
  IV U14433 ( .A(n14145), .Z(n14470) );
  NOR U14434 ( .A(n14471), .B(n14470), .Z(n14146) );
  NOR U14435 ( .A(n14147), .B(n14146), .Z(n14148) );
  IV U14436 ( .A(n14148), .Z(n14469) );
  XOR U14437 ( .A(n14150), .B(n14149), .Z(n14468) );
  NOR U14438 ( .A(n14469), .B(n14468), .Z(n14151) );
  NOR U14439 ( .A(n14152), .B(n14151), .Z(n14669) );
  XOR U14440 ( .A(n14154), .B(n14153), .Z(n14670) );
  NOR U14441 ( .A(n14669), .B(n14670), .Z(n14155) );
  NOR U14442 ( .A(n14156), .B(n14155), .Z(n14163) );
  NOR U14443 ( .A(n112), .B(n52), .Z(n14162) );
  IV U14444 ( .A(n14162), .Z(n14157) );
  NOR U14445 ( .A(n14163), .B(n14157), .Z(n14165) );
  XOR U14446 ( .A(n14159), .B(n14158), .Z(n14160) );
  XOR U14447 ( .A(n14161), .B(n14160), .Z(n14464) );
  XOR U14448 ( .A(n14163), .B(n14162), .Z(n14465) );
  NOR U14449 ( .A(n14464), .B(n14465), .Z(n14164) );
  NOR U14450 ( .A(n14165), .B(n14164), .Z(n14460) );
  XOR U14451 ( .A(n14167), .B(n14166), .Z(n14459) );
  NOR U14452 ( .A(n14460), .B(n14459), .Z(n14168) );
  NOR U14453 ( .A(n14169), .B(n14168), .Z(n14170) );
  IV U14454 ( .A(n14170), .Z(n14456) );
  NOR U14455 ( .A(n14457), .B(n14456), .Z(n14171) );
  NOR U14456 ( .A(n14172), .B(n14171), .Z(n14451) );
  NOR U14457 ( .A(n14173), .B(n14451), .Z(n14174) );
  NOR U14458 ( .A(n14175), .B(n14174), .Z(n14176) );
  IV U14459 ( .A(n14176), .Z(n14183) );
  NOR U14460 ( .A(n114), .B(n52), .Z(n14182) );
  IV U14461 ( .A(n14182), .Z(n14177) );
  NOR U14462 ( .A(n14183), .B(n14177), .Z(n14185) );
  XOR U14463 ( .A(n14179), .B(n14178), .Z(n14180) );
  XOR U14464 ( .A(n14181), .B(n14180), .Z(n14447) );
  XOR U14465 ( .A(n14183), .B(n14182), .Z(n14448) );
  NOR U14466 ( .A(n14447), .B(n14448), .Z(n14184) );
  NOR U14467 ( .A(n14185), .B(n14184), .Z(n14186) );
  IV U14468 ( .A(n14186), .Z(n14697) );
  NOR U14469 ( .A(n14698), .B(n14697), .Z(n14187) );
  NOR U14470 ( .A(n14188), .B(n14187), .Z(n14189) );
  IV U14471 ( .A(n14189), .Z(n14192) );
  NOR U14472 ( .A(n115), .B(n52), .Z(n14191) );
  IV U14473 ( .A(n14191), .Z(n14190) );
  NOR U14474 ( .A(n14192), .B(n14190), .Z(n14196) );
  XOR U14475 ( .A(n14192), .B(n14191), .Z(n14443) );
  XOR U14476 ( .A(n14194), .B(n14193), .Z(n14442) );
  NOR U14477 ( .A(n14443), .B(n14442), .Z(n14195) );
  NOR U14478 ( .A(n14196), .B(n14195), .Z(n14197) );
  IV U14479 ( .A(n14197), .Z(n14710) );
  XOR U14480 ( .A(n14199), .B(n14198), .Z(n14200) );
  IV U14481 ( .A(n14200), .Z(n14709) );
  NOR U14482 ( .A(n14710), .B(n14709), .Z(n14201) );
  NOR U14483 ( .A(n14202), .B(n14201), .Z(n14438) );
  XOR U14484 ( .A(n14204), .B(n14203), .Z(n14439) );
  NOR U14485 ( .A(n14438), .B(n14439), .Z(n14205) );
  NOR U14486 ( .A(n14206), .B(n14205), .Z(n14207) );
  IV U14487 ( .A(n14207), .Z(n14211) );
  NOR U14488 ( .A(n14208), .B(n14211), .Z(n14215) );
  XOR U14489 ( .A(n14210), .B(n14209), .Z(n14721) );
  IV U14490 ( .A(n14721), .Z(n14213) );
  XOR U14491 ( .A(n14212), .B(n14211), .Z(n14722) );
  NOR U14492 ( .A(n14213), .B(n14722), .Z(n14214) );
  NOR U14493 ( .A(n14215), .B(n14214), .Z(n14220) );
  XOR U14494 ( .A(n14217), .B(n14216), .Z(n14218) );
  XOR U14495 ( .A(n14219), .B(n14218), .Z(n14221) );
  NOR U14496 ( .A(n14220), .B(n14221), .Z(n14225) );
  XOR U14497 ( .A(n14221), .B(n14220), .Z(n14729) );
  IV U14498 ( .A(n14729), .Z(n14223) );
  NOR U14499 ( .A(n117), .B(n52), .Z(n14222) );
  IV U14500 ( .A(n14222), .Z(n14730) );
  NOR U14501 ( .A(n14223), .B(n14730), .Z(n14224) );
  NOR U14502 ( .A(n14225), .B(n14224), .Z(n14437) );
  XOR U14503 ( .A(n14227), .B(n14226), .Z(n14436) );
  NOR U14504 ( .A(n14437), .B(n14436), .Z(n14228) );
  NOR U14505 ( .A(n14229), .B(n14228), .Z(n14231) );
  IV U14506 ( .A(n14231), .Z(n14430) );
  NOR U14507 ( .A(n14230), .B(n14430), .Z(n14238) );
  IV U14508 ( .A(n14230), .Z(n14431) );
  NOR U14509 ( .A(n14231), .B(n14431), .Z(n14236) );
  XOR U14510 ( .A(n14233), .B(n14232), .Z(n14234) );
  XOR U14511 ( .A(n14235), .B(n14234), .Z(n14433) );
  NOR U14512 ( .A(n14236), .B(n14433), .Z(n14237) );
  NOR U14513 ( .A(n14238), .B(n14237), .Z(n14239) );
  IV U14514 ( .A(n14239), .Z(n14246) );
  NOR U14515 ( .A(n120), .B(n52), .Z(n14245) );
  IV U14516 ( .A(n14245), .Z(n14240) );
  NOR U14517 ( .A(n14246), .B(n14240), .Z(n14248) );
  XOR U14518 ( .A(n14242), .B(n14241), .Z(n14243) );
  XOR U14519 ( .A(n14244), .B(n14243), .Z(n14429) );
  XOR U14520 ( .A(n14246), .B(n14245), .Z(n14428) );
  NOR U14521 ( .A(n14429), .B(n14428), .Z(n14247) );
  NOR U14522 ( .A(n14248), .B(n14247), .Z(n14253) );
  XOR U14523 ( .A(n14250), .B(n14249), .Z(n14252) );
  IV U14524 ( .A(n14252), .Z(n14251) );
  NOR U14525 ( .A(n14253), .B(n14251), .Z(n14256) );
  XOR U14526 ( .A(n14253), .B(n14252), .Z(n14748) );
  NOR U14527 ( .A(n123), .B(n52), .Z(n14254) );
  IV U14528 ( .A(n14254), .Z(n14747) );
  NOR U14529 ( .A(n14748), .B(n14747), .Z(n14255) );
  NOR U14530 ( .A(n14256), .B(n14255), .Z(n14759) );
  XOR U14531 ( .A(n14258), .B(n14257), .Z(n14758) );
  NOR U14532 ( .A(n14759), .B(n14758), .Z(n14259) );
  NOR U14533 ( .A(n14260), .B(n14259), .Z(n14267) );
  NOR U14534 ( .A(n126), .B(n52), .Z(n14266) );
  IV U14535 ( .A(n14266), .Z(n14261) );
  NOR U14536 ( .A(n14267), .B(n14261), .Z(n14269) );
  XOR U14537 ( .A(n14263), .B(n14262), .Z(n14264) );
  XOR U14538 ( .A(n14265), .B(n14264), .Z(n14764) );
  XOR U14539 ( .A(n14267), .B(n14266), .Z(n14763) );
  NOR U14540 ( .A(n14764), .B(n14763), .Z(n14268) );
  NOR U14541 ( .A(n14269), .B(n14268), .Z(n14273) );
  XOR U14542 ( .A(n14271), .B(n14270), .Z(n14272) );
  NOR U14543 ( .A(n14273), .B(n14272), .Z(n14277) );
  XOR U14544 ( .A(n14273), .B(n14272), .Z(n14274) );
  IV U14545 ( .A(n14274), .Z(n14773) );
  NOR U14546 ( .A(n128), .B(n52), .Z(n14275) );
  IV U14547 ( .A(n14275), .Z(n14772) );
  NOR U14548 ( .A(n14773), .B(n14772), .Z(n14276) );
  NOR U14549 ( .A(n14277), .B(n14276), .Z(n14280) );
  NOR U14550 ( .A(n131), .B(n52), .Z(n14279) );
  IV U14551 ( .A(n14279), .Z(n14278) );
  NOR U14552 ( .A(n14280), .B(n14278), .Z(n14284) );
  XOR U14553 ( .A(n14280), .B(n14279), .Z(n14782) );
  XOR U14554 ( .A(n14282), .B(n14281), .Z(n14783) );
  NOR U14555 ( .A(n14782), .B(n14783), .Z(n14283) );
  NOR U14556 ( .A(n14284), .B(n14283), .Z(n14287) );
  NOR U14557 ( .A(n133), .B(n52), .Z(n14286) );
  IV U14558 ( .A(n14286), .Z(n14285) );
  NOR U14559 ( .A(n14287), .B(n14285), .Z(n14292) );
  XOR U14560 ( .A(n14287), .B(n14286), .Z(n14787) );
  XOR U14561 ( .A(n14289), .B(n14288), .Z(n14788) );
  IV U14562 ( .A(n14788), .Z(n14290) );
  NOR U14563 ( .A(n14787), .B(n14290), .Z(n14291) );
  NOR U14564 ( .A(n14292), .B(n14291), .Z(n14296) );
  XOR U14565 ( .A(n14294), .B(n14293), .Z(n14295) );
  NOR U14566 ( .A(n14296), .B(n14295), .Z(n14300) );
  XOR U14567 ( .A(n14296), .B(n14295), .Z(n14798) );
  IV U14568 ( .A(n14798), .Z(n14298) );
  NOR U14569 ( .A(n135), .B(n52), .Z(n14297) );
  IV U14570 ( .A(n14297), .Z(n14799) );
  NOR U14571 ( .A(n14298), .B(n14799), .Z(n14299) );
  NOR U14572 ( .A(n14300), .B(n14299), .Z(n14303) );
  NOR U14573 ( .A(n137), .B(n52), .Z(n14302) );
  IV U14574 ( .A(n14302), .Z(n14301) );
  NOR U14575 ( .A(n14303), .B(n14301), .Z(n14307) );
  XOR U14576 ( .A(n14303), .B(n14302), .Z(n14803) );
  XOR U14577 ( .A(n14305), .B(n14304), .Z(n14804) );
  NOR U14578 ( .A(n14803), .B(n14804), .Z(n14306) );
  NOR U14579 ( .A(n14307), .B(n14306), .Z(n14310) );
  NOR U14580 ( .A(n139), .B(n52), .Z(n14309) );
  IV U14581 ( .A(n14309), .Z(n14308) );
  NOR U14582 ( .A(n14310), .B(n14308), .Z(n14315) );
  XOR U14583 ( .A(n14310), .B(n14309), .Z(n14810) );
  XOR U14584 ( .A(n14312), .B(n14311), .Z(n14811) );
  IV U14585 ( .A(n14811), .Z(n14313) );
  NOR U14586 ( .A(n14810), .B(n14313), .Z(n14314) );
  NOR U14587 ( .A(n14315), .B(n14314), .Z(n14319) );
  XOR U14588 ( .A(n14317), .B(n14316), .Z(n14318) );
  NOR U14589 ( .A(n14319), .B(n14318), .Z(n14323) );
  XOR U14590 ( .A(n14319), .B(n14318), .Z(n14320) );
  IV U14591 ( .A(n14320), .Z(n14425) );
  NOR U14592 ( .A(n141), .B(n52), .Z(n14426) );
  IV U14593 ( .A(n14426), .Z(n14321) );
  NOR U14594 ( .A(n14425), .B(n14321), .Z(n14322) );
  NOR U14595 ( .A(n14323), .B(n14322), .Z(n14326) );
  NOR U14596 ( .A(n143), .B(n52), .Z(n14325) );
  IV U14597 ( .A(n14325), .Z(n14324) );
  NOR U14598 ( .A(n14326), .B(n14324), .Z(n14330) );
  XOR U14599 ( .A(n14326), .B(n14325), .Z(n14825) );
  XOR U14600 ( .A(n14328), .B(n14327), .Z(n14826) );
  NOR U14601 ( .A(n14825), .B(n14826), .Z(n14329) );
  NOR U14602 ( .A(n14330), .B(n14329), .Z(n14333) );
  NOR U14603 ( .A(n145), .B(n52), .Z(n14332) );
  IV U14604 ( .A(n14332), .Z(n14331) );
  NOR U14605 ( .A(n14333), .B(n14331), .Z(n14338) );
  XOR U14606 ( .A(n14333), .B(n14332), .Z(n14830) );
  XOR U14607 ( .A(n14335), .B(n14334), .Z(n14831) );
  IV U14608 ( .A(n14831), .Z(n14336) );
  NOR U14609 ( .A(n14830), .B(n14336), .Z(n14337) );
  NOR U14610 ( .A(n14338), .B(n14337), .Z(n14342) );
  XOR U14611 ( .A(n14340), .B(n14339), .Z(n14341) );
  NOR U14612 ( .A(n14342), .B(n14341), .Z(n14346) );
  XOR U14613 ( .A(n14342), .B(n14341), .Z(n14841) );
  IV U14614 ( .A(n14841), .Z(n14344) );
  NOR U14615 ( .A(n147), .B(n52), .Z(n14343) );
  IV U14616 ( .A(n14343), .Z(n14842) );
  NOR U14617 ( .A(n14344), .B(n14842), .Z(n14345) );
  NOR U14618 ( .A(n14346), .B(n14345), .Z(n14849) );
  IV U14619 ( .A(n14849), .Z(n14347) );
  NOR U14620 ( .A(n14846), .B(n14347), .Z(n14353) );
  XOR U14621 ( .A(n14349), .B(n14348), .Z(n14847) );
  IV U14622 ( .A(n14846), .Z(n14350) );
  NOR U14623 ( .A(n14849), .B(n14350), .Z(n14351) );
  NOR U14624 ( .A(n14847), .B(n14351), .Z(n14352) );
  NOR U14625 ( .A(n14353), .B(n14352), .Z(n14357) );
  IV U14626 ( .A(n14357), .Z(n14355) );
  NOR U14627 ( .A(n150), .B(n52), .Z(n14354) );
  IV U14628 ( .A(n14354), .Z(n14356) );
  NOR U14629 ( .A(n14355), .B(n14356), .Z(n14361) );
  XOR U14630 ( .A(n14357), .B(n14356), .Z(n14855) );
  XOR U14631 ( .A(n14359), .B(n14358), .Z(n14854) );
  NOR U14632 ( .A(n14855), .B(n14854), .Z(n14360) );
  NOR U14633 ( .A(n14361), .B(n14360), .Z(n14365) );
  XOR U14634 ( .A(n14363), .B(n14362), .Z(n14364) );
  NOR U14635 ( .A(n14365), .B(n14364), .Z(n14369) );
  XOR U14636 ( .A(n14365), .B(n14364), .Z(n14366) );
  IV U14637 ( .A(n14366), .Z(n14865) );
  NOR U14638 ( .A(n153), .B(n52), .Z(n14866) );
  IV U14639 ( .A(n14866), .Z(n14367) );
  NOR U14640 ( .A(n14865), .B(n14367), .Z(n14368) );
  NOR U14641 ( .A(n14369), .B(n14368), .Z(n14871) );
  XOR U14642 ( .A(n14371), .B(n14370), .Z(n14870) );
  NOR U14643 ( .A(n14871), .B(n14870), .Z(n14372) );
  NOR U14644 ( .A(n14373), .B(n14372), .Z(n14378) );
  NOR U14645 ( .A(n156), .B(n52), .Z(n14377) );
  IV U14646 ( .A(n14377), .Z(n14374) );
  NOR U14647 ( .A(n14378), .B(n14374), .Z(n14380) );
  XOR U14648 ( .A(n14376), .B(n14375), .Z(n14878) );
  XOR U14649 ( .A(n14378), .B(n14377), .Z(n14877) );
  NOR U14650 ( .A(n14878), .B(n14877), .Z(n14379) );
  NOR U14651 ( .A(n14380), .B(n14379), .Z(n14385) );
  XOR U14652 ( .A(n14382), .B(n14381), .Z(n14384) );
  IV U14653 ( .A(n14384), .Z(n14383) );
  NOR U14654 ( .A(n14385), .B(n14383), .Z(n14388) );
  XOR U14655 ( .A(n14385), .B(n14384), .Z(n14422) );
  NOR U14656 ( .A(n158), .B(n52), .Z(n14423) );
  IV U14657 ( .A(n14423), .Z(n14386) );
  NOR U14658 ( .A(n14422), .B(n14386), .Z(n14387) );
  NOR U14659 ( .A(n14388), .B(n14387), .Z(n14893) );
  XOR U14660 ( .A(n14390), .B(n14389), .Z(n14892) );
  NOR U14661 ( .A(n14893), .B(n14892), .Z(n14391) );
  NOR U14662 ( .A(n14392), .B(n14391), .Z(n14397) );
  NOR U14663 ( .A(n163), .B(n52), .Z(n14396) );
  IV U14664 ( .A(n14396), .Z(n14393) );
  NOR U14665 ( .A(n14397), .B(n14393), .Z(n14400) );
  XOR U14666 ( .A(n14395), .B(n14394), .Z(n14898) );
  IV U14667 ( .A(n14898), .Z(n14398) );
  XOR U14668 ( .A(n14397), .B(n14396), .Z(n14897) );
  NOR U14669 ( .A(n14398), .B(n14897), .Z(n14399) );
  NOR U14670 ( .A(n14400), .B(n14399), .Z(n14404) );
  XOR U14671 ( .A(n14402), .B(n14401), .Z(n14403) );
  NOR U14672 ( .A(n14404), .B(n14403), .Z(n14408) );
  XOR U14673 ( .A(n14404), .B(n14403), .Z(n14419) );
  IV U14674 ( .A(n14419), .Z(n14406) );
  NOR U14675 ( .A(n165), .B(n52), .Z(n14405) );
  IV U14676 ( .A(n14405), .Z(n14420) );
  NOR U14677 ( .A(n14406), .B(n14420), .Z(n14407) );
  NOR U14678 ( .A(n14408), .B(n14407), .Z(n14411) );
  NOR U14679 ( .A(n167), .B(n52), .Z(n14410) );
  IV U14680 ( .A(n14410), .Z(n14409) );
  NOR U14681 ( .A(n14411), .B(n14409), .Z(n14416) );
  XOR U14682 ( .A(n14411), .B(n14410), .Z(n14909) );
  XOR U14683 ( .A(n14413), .B(n14412), .Z(n14910) );
  IV U14684 ( .A(n14910), .Z(n14414) );
  NOR U14685 ( .A(n14909), .B(n14414), .Z(n14415) );
  NOR U14686 ( .A(n14416), .B(n14415), .Z(n14912) );
  XOR U14687 ( .A(n14418), .B(n14417), .Z(n14911) );
  NOR U14688 ( .A(n14912), .B(n14911), .Z(n31643) );
  XOR U14689 ( .A(n14420), .B(n14419), .Z(n14905) );
  NOR U14690 ( .A(n167), .B(n53), .Z(n14906) );
  IV U14691 ( .A(n14906), .Z(n14421) );
  NOR U14692 ( .A(n14905), .B(n14421), .Z(n14908) );
  XOR U14693 ( .A(n14423), .B(n14422), .Z(n14885) );
  NOR U14694 ( .A(n161), .B(n53), .Z(n14886) );
  IV U14695 ( .A(n14886), .Z(n14424) );
  NOR U14696 ( .A(n14885), .B(n14424), .Z(n14888) );
  XOR U14697 ( .A(n14426), .B(n14425), .Z(n14818) );
  NOR U14698 ( .A(n143), .B(n53), .Z(n14819) );
  IV U14699 ( .A(n14819), .Z(n14427) );
  NOR U14700 ( .A(n14818), .B(n14427), .Z(n14821) );
  NOR U14701 ( .A(n131), .B(n53), .Z(n15284) );
  NOR U14702 ( .A(n125), .B(n53), .Z(n14749) );
  XOR U14703 ( .A(n14429), .B(n14428), .Z(n14743) );
  XOR U14704 ( .A(n14431), .B(n14430), .Z(n14432) );
  XOR U14705 ( .A(n14433), .B(n14432), .Z(n15240) );
  NOR U14706 ( .A(n120), .B(n53), .Z(n14434) );
  IV U14707 ( .A(n14434), .Z(n15237) );
  NOR U14708 ( .A(n15240), .B(n15237), .Z(n14741) );
  IV U14709 ( .A(n15240), .Z(n14435) );
  NOR U14710 ( .A(n14435), .B(n14434), .Z(n14739) );
  XOR U14711 ( .A(n14437), .B(n14436), .Z(n14735) );
  NOR U14712 ( .A(n80), .B(n53), .Z(n14440) );
  XOR U14713 ( .A(n14439), .B(n14438), .Z(n14441) );
  IV U14714 ( .A(n14441), .Z(n15215) );
  NOR U14715 ( .A(n14440), .B(n15215), .Z(n14718) );
  IV U14716 ( .A(n14440), .Z(n15213) );
  NOR U14717 ( .A(n14441), .B(n15213), .Z(n14716) );
  XOR U14718 ( .A(n14443), .B(n14442), .Z(n14444) );
  NOR U14719 ( .A(n81), .B(n53), .Z(n14445) );
  NOR U14720 ( .A(n14444), .B(n14445), .Z(n14706) );
  IV U14721 ( .A(n14444), .Z(n15199) );
  IV U14722 ( .A(n14445), .Z(n15198) );
  NOR U14723 ( .A(n15199), .B(n15198), .Z(n14704) );
  NOR U14724 ( .A(n115), .B(n53), .Z(n14446) );
  IV U14725 ( .A(n14446), .Z(n14700) );
  XOR U14726 ( .A(n14448), .B(n14447), .Z(n14449) );
  NOR U14727 ( .A(n82), .B(n53), .Z(n14450) );
  NOR U14728 ( .A(n14449), .B(n14450), .Z(n14695) );
  IV U14729 ( .A(n14449), .Z(n14934) );
  IV U14730 ( .A(n14450), .Z(n14932) );
  NOR U14731 ( .A(n14934), .B(n14932), .Z(n14693) );
  XOR U14732 ( .A(n14452), .B(n14451), .Z(n14453) );
  XOR U14733 ( .A(n14454), .B(n14453), .Z(n14688) );
  NOR U14734 ( .A(n114), .B(n53), .Z(n14689) );
  IV U14735 ( .A(n14689), .Z(n14455) );
  NOR U14736 ( .A(n14688), .B(n14455), .Z(n14691) );
  XOR U14737 ( .A(n14457), .B(n14456), .Z(n14684) );
  NOR U14738 ( .A(n83), .B(n53), .Z(n14458) );
  IV U14739 ( .A(n14458), .Z(n14683) );
  NOR U14740 ( .A(n14684), .B(n14683), .Z(n14687) );
  XOR U14741 ( .A(n14460), .B(n14459), .Z(n14679) );
  IV U14742 ( .A(n14679), .Z(n14462) );
  NOR U14743 ( .A(n113), .B(n53), .Z(n14461) );
  IV U14744 ( .A(n14461), .Z(n14680) );
  NOR U14745 ( .A(n14462), .B(n14680), .Z(n14682) );
  NOR U14746 ( .A(n84), .B(n53), .Z(n14463) );
  IV U14747 ( .A(n14463), .Z(n14675) );
  IV U14748 ( .A(n14464), .Z(n14466) );
  XOR U14749 ( .A(n14466), .B(n14465), .Z(n14674) );
  NOR U14750 ( .A(n14675), .B(n14674), .Z(n14678) );
  NOR U14751 ( .A(n112), .B(n53), .Z(n14467) );
  IV U14752 ( .A(n14467), .Z(n14668) );
  NOR U14753 ( .A(n85), .B(n53), .Z(n14662) );
  XOR U14754 ( .A(n14469), .B(n14468), .Z(n14661) );
  NOR U14755 ( .A(n14662), .B(n14661), .Z(n14665) );
  XOR U14756 ( .A(n14471), .B(n14470), .Z(n14657) );
  NOR U14757 ( .A(n111), .B(n53), .Z(n14656) );
  IV U14758 ( .A(n14656), .Z(n14472) );
  NOR U14759 ( .A(n14657), .B(n14472), .Z(n14659) );
  XOR U14760 ( .A(n14474), .B(n14473), .Z(n14652) );
  NOR U14761 ( .A(n86), .B(n53), .Z(n14653) );
  IV U14762 ( .A(n14653), .Z(n14475) );
  NOR U14763 ( .A(n14652), .B(n14475), .Z(n14655) );
  XOR U14764 ( .A(n14477), .B(n14476), .Z(n14478) );
  XOR U14765 ( .A(n14479), .B(n14478), .Z(n14649) );
  NOR U14766 ( .A(n110), .B(n53), .Z(n14648) );
  IV U14767 ( .A(n14648), .Z(n14480) );
  NOR U14768 ( .A(n14649), .B(n14480), .Z(n14651) );
  XOR U14769 ( .A(n14482), .B(n14481), .Z(n14644) );
  NOR U14770 ( .A(n109), .B(n53), .Z(n14645) );
  IV U14771 ( .A(n14645), .Z(n14483) );
  NOR U14772 ( .A(n14644), .B(n14483), .Z(n14647) );
  NOR U14773 ( .A(n87), .B(n53), .Z(n14486) );
  XOR U14774 ( .A(n14485), .B(n14484), .Z(n14487) );
  NOR U14775 ( .A(n14486), .B(n14487), .Z(n14635) );
  IV U14776 ( .A(n14486), .Z(n14960) );
  IV U14777 ( .A(n14487), .Z(n14959) );
  NOR U14778 ( .A(n14960), .B(n14959), .Z(n14633) );
  XOR U14779 ( .A(n14489), .B(n14488), .Z(n14628) );
  IV U14780 ( .A(n14628), .Z(n14491) );
  NOR U14781 ( .A(n107), .B(n53), .Z(n14490) );
  IV U14782 ( .A(n14490), .Z(n14629) );
  NOR U14783 ( .A(n14491), .B(n14629), .Z(n14631) );
  NOR U14784 ( .A(n88), .B(n53), .Z(n14623) );
  XOR U14785 ( .A(n14493), .B(n14492), .Z(n14622) );
  NOR U14786 ( .A(n14623), .B(n14622), .Z(n14626) );
  XOR U14787 ( .A(n14495), .B(n14494), .Z(n14618) );
  NOR U14788 ( .A(n106), .B(n53), .Z(n14617) );
  IV U14789 ( .A(n14617), .Z(n14496) );
  NOR U14790 ( .A(n14618), .B(n14496), .Z(n14620) );
  XOR U14791 ( .A(n14498), .B(n14497), .Z(n14613) );
  NOR U14792 ( .A(n105), .B(n53), .Z(n14614) );
  IV U14793 ( .A(n14614), .Z(n14499) );
  NOR U14794 ( .A(n14613), .B(n14499), .Z(n14616) );
  XOR U14795 ( .A(n14501), .B(n14500), .Z(n14610) );
  NOR U14796 ( .A(n104), .B(n53), .Z(n14609) );
  IV U14797 ( .A(n14609), .Z(n14502) );
  NOR U14798 ( .A(n14610), .B(n14502), .Z(n14612) );
  IV U14799 ( .A(n14503), .Z(n14505) );
  XOR U14800 ( .A(n14505), .B(n14504), .Z(n14605) );
  NOR U14801 ( .A(n89), .B(n53), .Z(n14606) );
  IV U14802 ( .A(n14606), .Z(n14506) );
  NOR U14803 ( .A(n14605), .B(n14506), .Z(n14608) );
  IV U14804 ( .A(n14507), .Z(n14509) );
  XOR U14805 ( .A(n14509), .B(n14508), .Z(n14601) );
  NOR U14806 ( .A(n103), .B(n53), .Z(n14602) );
  IV U14807 ( .A(n14602), .Z(n14510) );
  NOR U14808 ( .A(n14601), .B(n14510), .Z(n14604) );
  IV U14809 ( .A(n14511), .Z(n14513) );
  XOR U14810 ( .A(n14513), .B(n14512), .Z(n14597) );
  NOR U14811 ( .A(n90), .B(n53), .Z(n14598) );
  IV U14812 ( .A(n14598), .Z(n14514) );
  NOR U14813 ( .A(n14597), .B(n14514), .Z(n14600) );
  IV U14814 ( .A(n14515), .Z(n14517) );
  XOR U14815 ( .A(n14517), .B(n14516), .Z(n14593) );
  NOR U14816 ( .A(n102), .B(n53), .Z(n14594) );
  IV U14817 ( .A(n14594), .Z(n14518) );
  NOR U14818 ( .A(n14593), .B(n14518), .Z(n14596) );
  IV U14819 ( .A(n14519), .Z(n14521) );
  XOR U14820 ( .A(n14521), .B(n14520), .Z(n14589) );
  NOR U14821 ( .A(n101), .B(n53), .Z(n14590) );
  IV U14822 ( .A(n14590), .Z(n14522) );
  NOR U14823 ( .A(n14589), .B(n14522), .Z(n14592) );
  IV U14824 ( .A(n14523), .Z(n14525) );
  XOR U14825 ( .A(n14525), .B(n14524), .Z(n14585) );
  NOR U14826 ( .A(n100), .B(n53), .Z(n14586) );
  IV U14827 ( .A(n14586), .Z(n14526) );
  NOR U14828 ( .A(n14585), .B(n14526), .Z(n14588) );
  IV U14829 ( .A(n14527), .Z(n14529) );
  XOR U14830 ( .A(n14529), .B(n14528), .Z(n14581) );
  NOR U14831 ( .A(n99), .B(n53), .Z(n14582) );
  IV U14832 ( .A(n14582), .Z(n14530) );
  NOR U14833 ( .A(n14581), .B(n14530), .Z(n14584) );
  IV U14834 ( .A(n14531), .Z(n14533) );
  XOR U14835 ( .A(n14533), .B(n14532), .Z(n14577) );
  NOR U14836 ( .A(n98), .B(n53), .Z(n14578) );
  IV U14837 ( .A(n14578), .Z(n14534) );
  NOR U14838 ( .A(n14577), .B(n14534), .Z(n14580) );
  XOR U14839 ( .A(n14536), .B(n14535), .Z(n14573) );
  NOR U14840 ( .A(n91), .B(n53), .Z(n14574) );
  IV U14841 ( .A(n14574), .Z(n14537) );
  NOR U14842 ( .A(n14573), .B(n14537), .Z(n14576) );
  XOR U14843 ( .A(n14539), .B(n14538), .Z(n14561) );
  IV U14844 ( .A(n14561), .Z(n14541) );
  NOR U14845 ( .A(n96), .B(n53), .Z(n14540) );
  IV U14846 ( .A(n14540), .Z(n14562) );
  NOR U14847 ( .A(n14541), .B(n14562), .Z(n14564) );
  NOR U14848 ( .A(n95), .B(n53), .Z(n14558) );
  IV U14849 ( .A(n14558), .Z(n14544) );
  XOR U14850 ( .A(n14543), .B(n14542), .Z(n14557) );
  NOR U14851 ( .A(n14544), .B(n14557), .Z(n14560) );
  NOR U14852 ( .A(n93), .B(n53), .Z(n15547) );
  IV U14853 ( .A(n15547), .Z(n14545) );
  NOR U14854 ( .A(n52), .B(n168), .Z(n14553) );
  IV U14855 ( .A(n14553), .Z(n14548) );
  NOR U14856 ( .A(n14545), .B(n14548), .Z(n14546) );
  IV U14857 ( .A(n14546), .Z(n14547) );
  NOR U14858 ( .A(n94), .B(n14547), .Z(n14556) );
  NOR U14859 ( .A(n14548), .B(n93), .Z(n14549) );
  XOR U14860 ( .A(n94), .B(n14549), .Z(n14550) );
  NOR U14861 ( .A(n53), .B(n14550), .Z(n14551) );
  IV U14862 ( .A(n14551), .Z(n15024) );
  XOR U14863 ( .A(n14553), .B(n14552), .Z(n15023) );
  IV U14864 ( .A(n15023), .Z(n14554) );
  NOR U14865 ( .A(n15024), .B(n14554), .Z(n14555) );
  NOR U14866 ( .A(n14556), .B(n14555), .Z(n15020) );
  XOR U14867 ( .A(n14558), .B(n14557), .Z(n15019) );
  NOR U14868 ( .A(n15020), .B(n15019), .Z(n14559) );
  NOR U14869 ( .A(n14560), .B(n14559), .Z(n15047) );
  XOR U14870 ( .A(n14562), .B(n14561), .Z(n15046) );
  NOR U14871 ( .A(n15047), .B(n15046), .Z(n14563) );
  NOR U14872 ( .A(n14564), .B(n14563), .Z(n14569) );
  XOR U14873 ( .A(n14566), .B(n14565), .Z(n14568) );
  IV U14874 ( .A(n14568), .Z(n14567) );
  NOR U14875 ( .A(n14569), .B(n14567), .Z(n14572) );
  XOR U14876 ( .A(n14569), .B(n14568), .Z(n15016) );
  NOR U14877 ( .A(n97), .B(n53), .Z(n15017) );
  IV U14878 ( .A(n15017), .Z(n14570) );
  NOR U14879 ( .A(n15016), .B(n14570), .Z(n14571) );
  NOR U14880 ( .A(n14572), .B(n14571), .Z(n15012) );
  XOR U14881 ( .A(n14574), .B(n14573), .Z(n15013) );
  NOR U14882 ( .A(n15012), .B(n15013), .Z(n14575) );
  NOR U14883 ( .A(n14576), .B(n14575), .Z(n15008) );
  XOR U14884 ( .A(n14578), .B(n14577), .Z(n15009) );
  NOR U14885 ( .A(n15008), .B(n15009), .Z(n14579) );
  NOR U14886 ( .A(n14580), .B(n14579), .Z(n15004) );
  XOR U14887 ( .A(n14582), .B(n14581), .Z(n15005) );
  NOR U14888 ( .A(n15004), .B(n15005), .Z(n14583) );
  NOR U14889 ( .A(n14584), .B(n14583), .Z(n15000) );
  XOR U14890 ( .A(n14586), .B(n14585), .Z(n15001) );
  NOR U14891 ( .A(n15000), .B(n15001), .Z(n14587) );
  NOR U14892 ( .A(n14588), .B(n14587), .Z(n14996) );
  XOR U14893 ( .A(n14590), .B(n14589), .Z(n14997) );
  NOR U14894 ( .A(n14996), .B(n14997), .Z(n14591) );
  NOR U14895 ( .A(n14592), .B(n14591), .Z(n14993) );
  XOR U14896 ( .A(n14594), .B(n14593), .Z(n14992) );
  NOR U14897 ( .A(n14993), .B(n14992), .Z(n14595) );
  NOR U14898 ( .A(n14596), .B(n14595), .Z(n14988) );
  XOR U14899 ( .A(n14598), .B(n14597), .Z(n14989) );
  NOR U14900 ( .A(n14988), .B(n14989), .Z(n14599) );
  NOR U14901 ( .A(n14600), .B(n14599), .Z(n14984) );
  XOR U14902 ( .A(n14602), .B(n14601), .Z(n14985) );
  NOR U14903 ( .A(n14984), .B(n14985), .Z(n14603) );
  NOR U14904 ( .A(n14604), .B(n14603), .Z(n14980) );
  XOR U14905 ( .A(n14606), .B(n14605), .Z(n14981) );
  NOR U14906 ( .A(n14980), .B(n14981), .Z(n14607) );
  NOR U14907 ( .A(n14608), .B(n14607), .Z(n14979) );
  XOR U14908 ( .A(n14610), .B(n14609), .Z(n14978) );
  NOR U14909 ( .A(n14979), .B(n14978), .Z(n14611) );
  NOR U14910 ( .A(n14612), .B(n14611), .Z(n14974) );
  XOR U14911 ( .A(n14614), .B(n14613), .Z(n14975) );
  NOR U14912 ( .A(n14974), .B(n14975), .Z(n14615) );
  NOR U14913 ( .A(n14616), .B(n14615), .Z(n14973) );
  XOR U14914 ( .A(n14618), .B(n14617), .Z(n14972) );
  NOR U14915 ( .A(n14973), .B(n14972), .Z(n14619) );
  NOR U14916 ( .A(n14620), .B(n14619), .Z(n14621) );
  IV U14917 ( .A(n14621), .Z(n14970) );
  XOR U14918 ( .A(n14623), .B(n14622), .Z(n14624) );
  IV U14919 ( .A(n14624), .Z(n14969) );
  NOR U14920 ( .A(n14970), .B(n14969), .Z(n14625) );
  NOR U14921 ( .A(n14626), .B(n14625), .Z(n14627) );
  IV U14922 ( .A(n14627), .Z(n14965) );
  XOR U14923 ( .A(n14629), .B(n14628), .Z(n14964) );
  NOR U14924 ( .A(n14965), .B(n14964), .Z(n14630) );
  NOR U14925 ( .A(n14631), .B(n14630), .Z(n14962) );
  IV U14926 ( .A(n14962), .Z(n14632) );
  NOR U14927 ( .A(n14633), .B(n14632), .Z(n14634) );
  NOR U14928 ( .A(n14635), .B(n14634), .Z(n14636) );
  IV U14929 ( .A(n14636), .Z(n14641) );
  NOR U14930 ( .A(n108), .B(n53), .Z(n14640) );
  IV U14931 ( .A(n14640), .Z(n14637) );
  NOR U14932 ( .A(n14641), .B(n14637), .Z(n14643) );
  XOR U14933 ( .A(n14639), .B(n14638), .Z(n14957) );
  XOR U14934 ( .A(n14641), .B(n14640), .Z(n14958) );
  NOR U14935 ( .A(n14957), .B(n14958), .Z(n14642) );
  NOR U14936 ( .A(n14643), .B(n14642), .Z(n14954) );
  XOR U14937 ( .A(n14645), .B(n14644), .Z(n14953) );
  NOR U14938 ( .A(n14954), .B(n14953), .Z(n14646) );
  NOR U14939 ( .A(n14647), .B(n14646), .Z(n14952) );
  XOR U14940 ( .A(n14649), .B(n14648), .Z(n14951) );
  NOR U14941 ( .A(n14952), .B(n14951), .Z(n14650) );
  NOR U14942 ( .A(n14651), .B(n14650), .Z(n15141) );
  XOR U14943 ( .A(n14653), .B(n14652), .Z(n15142) );
  NOR U14944 ( .A(n15141), .B(n15142), .Z(n14654) );
  NOR U14945 ( .A(n14655), .B(n14654), .Z(n14947) );
  XOR U14946 ( .A(n14657), .B(n14656), .Z(n14948) );
  NOR U14947 ( .A(n14947), .B(n14948), .Z(n14658) );
  NOR U14948 ( .A(n14659), .B(n14658), .Z(n14660) );
  IV U14949 ( .A(n14660), .Z(n14945) );
  XOR U14950 ( .A(n14662), .B(n14661), .Z(n14663) );
  IV U14951 ( .A(n14663), .Z(n14944) );
  NOR U14952 ( .A(n14945), .B(n14944), .Z(n14664) );
  NOR U14953 ( .A(n14665), .B(n14664), .Z(n14667) );
  IV U14954 ( .A(n14667), .Z(n14666) );
  NOR U14955 ( .A(n14668), .B(n14666), .Z(n14673) );
  XOR U14956 ( .A(n14668), .B(n14667), .Z(n14943) );
  XOR U14957 ( .A(n14670), .B(n14669), .Z(n14671) );
  IV U14958 ( .A(n14671), .Z(n14942) );
  NOR U14959 ( .A(n14943), .B(n14942), .Z(n14672) );
  NOR U14960 ( .A(n14673), .B(n14672), .Z(n15167) );
  XOR U14961 ( .A(n14675), .B(n14674), .Z(n15168) );
  IV U14962 ( .A(n15168), .Z(n14676) );
  NOR U14963 ( .A(n15167), .B(n14676), .Z(n14677) );
  NOR U14964 ( .A(n14678), .B(n14677), .Z(n14938) );
  XOR U14965 ( .A(n14680), .B(n14679), .Z(n14937) );
  NOR U14966 ( .A(n14938), .B(n14937), .Z(n14681) );
  NOR U14967 ( .A(n14682), .B(n14681), .Z(n15175) );
  XOR U14968 ( .A(n14684), .B(n14683), .Z(n15176) );
  IV U14969 ( .A(n15176), .Z(n14685) );
  NOR U14970 ( .A(n15175), .B(n14685), .Z(n14686) );
  NOR U14971 ( .A(n14687), .B(n14686), .Z(n14936) );
  XOR U14972 ( .A(n14689), .B(n14688), .Z(n14935) );
  NOR U14973 ( .A(n14936), .B(n14935), .Z(n14690) );
  NOR U14974 ( .A(n14691), .B(n14690), .Z(n14692) );
  IV U14975 ( .A(n14692), .Z(n14931) );
  NOR U14976 ( .A(n14693), .B(n14931), .Z(n14694) );
  NOR U14977 ( .A(n14695), .B(n14694), .Z(n14699) );
  IV U14978 ( .A(n14699), .Z(n14696) );
  NOR U14979 ( .A(n14700), .B(n14696), .Z(n14702) );
  XOR U14980 ( .A(n14698), .B(n14697), .Z(n14927) );
  XOR U14981 ( .A(n14700), .B(n14699), .Z(n14928) );
  NOR U14982 ( .A(n14927), .B(n14928), .Z(n14701) );
  NOR U14983 ( .A(n14702), .B(n14701), .Z(n15201) );
  IV U14984 ( .A(n15201), .Z(n14703) );
  NOR U14985 ( .A(n14704), .B(n14703), .Z(n14705) );
  NOR U14986 ( .A(n14706), .B(n14705), .Z(n14707) );
  IV U14987 ( .A(n14707), .Z(n14712) );
  NOR U14988 ( .A(n116), .B(n53), .Z(n14711) );
  IV U14989 ( .A(n14711), .Z(n14708) );
  NOR U14990 ( .A(n14712), .B(n14708), .Z(n14714) );
  XOR U14991 ( .A(n14710), .B(n14709), .Z(n14923) );
  XOR U14992 ( .A(n14712), .B(n14711), .Z(n14924) );
  NOR U14993 ( .A(n14923), .B(n14924), .Z(n14713) );
  NOR U14994 ( .A(n14714), .B(n14713), .Z(n14715) );
  IV U14995 ( .A(n14715), .Z(n15212) );
  NOR U14996 ( .A(n14716), .B(n15212), .Z(n14717) );
  NOR U14997 ( .A(n14718), .B(n14717), .Z(n14720) );
  IV U14998 ( .A(n14720), .Z(n14918) );
  NOR U14999 ( .A(n117), .B(n53), .Z(n14719) );
  IV U15000 ( .A(n14719), .Z(n14917) );
  NOR U15001 ( .A(n14918), .B(n14917), .Z(n14725) );
  NOR U15002 ( .A(n14720), .B(n14719), .Z(n14723) );
  XOR U15003 ( .A(n14722), .B(n14721), .Z(n14920) );
  NOR U15004 ( .A(n14723), .B(n14920), .Z(n14724) );
  NOR U15005 ( .A(n14725), .B(n14724), .Z(n14728) );
  NOR U15006 ( .A(n79), .B(n53), .Z(n14727) );
  IV U15007 ( .A(n14727), .Z(n14726) );
  NOR U15008 ( .A(n14728), .B(n14726), .Z(n14732) );
  XOR U15009 ( .A(n14728), .B(n14727), .Z(n14916) );
  XOR U15010 ( .A(n14730), .B(n14729), .Z(n14915) );
  NOR U15011 ( .A(n14916), .B(n14915), .Z(n14731) );
  NOR U15012 ( .A(n14732), .B(n14731), .Z(n14734) );
  IV U15013 ( .A(n14734), .Z(n14733) );
  NOR U15014 ( .A(n14735), .B(n14733), .Z(n14737) );
  NOR U15015 ( .A(n119), .B(n53), .Z(n15232) );
  XOR U15016 ( .A(n14735), .B(n14734), .Z(n15231) );
  NOR U15017 ( .A(n15232), .B(n15231), .Z(n14736) );
  NOR U15018 ( .A(n14737), .B(n14736), .Z(n14738) );
  IV U15019 ( .A(n14738), .Z(n15238) );
  NOR U15020 ( .A(n14739), .B(n15238), .Z(n14740) );
  NOR U15021 ( .A(n14741), .B(n14740), .Z(n15247) );
  IV U15022 ( .A(n15247), .Z(n14742) );
  NOR U15023 ( .A(n14743), .B(n14742), .Z(n14746) );
  NOR U15024 ( .A(n123), .B(n53), .Z(n15248) );
  IV U15025 ( .A(n14743), .Z(n15250) );
  NOR U15026 ( .A(n15247), .B(n15250), .Z(n14744) );
  NOR U15027 ( .A(n15248), .B(n14744), .Z(n14745) );
  NOR U15028 ( .A(n14746), .B(n14745), .Z(n14750) );
  NOR U15029 ( .A(n14749), .B(n14750), .Z(n14753) );
  XOR U15030 ( .A(n14748), .B(n14747), .Z(n15259) );
  IV U15031 ( .A(n14749), .Z(n15257) );
  IV U15032 ( .A(n14750), .Z(n15256) );
  NOR U15033 ( .A(n15257), .B(n15256), .Z(n14751) );
  NOR U15034 ( .A(n15259), .B(n14751), .Z(n14752) );
  NOR U15035 ( .A(n14753), .B(n14752), .Z(n14757) );
  IV U15036 ( .A(n14757), .Z(n14755) );
  NOR U15037 ( .A(n126), .B(n53), .Z(n14754) );
  IV U15038 ( .A(n14754), .Z(n14756) );
  NOR U15039 ( .A(n14755), .B(n14756), .Z(n14762) );
  XOR U15040 ( .A(n14757), .B(n14756), .Z(n15266) );
  XOR U15041 ( .A(n14759), .B(n14758), .Z(n15265) );
  IV U15042 ( .A(n15265), .Z(n14760) );
  NOR U15043 ( .A(n15266), .B(n14760), .Z(n14761) );
  NOR U15044 ( .A(n14762), .B(n14761), .Z(n14765) );
  XOR U15045 ( .A(n14764), .B(n14763), .Z(n14766) );
  IV U15046 ( .A(n14766), .Z(n15277) );
  NOR U15047 ( .A(n14765), .B(n15277), .Z(n14770) );
  IV U15048 ( .A(n14765), .Z(n15274) );
  NOR U15049 ( .A(n14766), .B(n15274), .Z(n14768) );
  NOR U15050 ( .A(n128), .B(n53), .Z(n14767) );
  IV U15051 ( .A(n14767), .Z(n15275) );
  NOR U15052 ( .A(n14768), .B(n15275), .Z(n14769) );
  NOR U15053 ( .A(n14770), .B(n14769), .Z(n15287) );
  IV U15054 ( .A(n15287), .Z(n14771) );
  NOR U15055 ( .A(n15284), .B(n14771), .Z(n14777) );
  XOR U15056 ( .A(n14773), .B(n14772), .Z(n15285) );
  IV U15057 ( .A(n15284), .Z(n14774) );
  NOR U15058 ( .A(n15287), .B(n14774), .Z(n14775) );
  NOR U15059 ( .A(n15285), .B(n14775), .Z(n14776) );
  NOR U15060 ( .A(n14777), .B(n14776), .Z(n14781) );
  IV U15061 ( .A(n14781), .Z(n14779) );
  NOR U15062 ( .A(n133), .B(n53), .Z(n14778) );
  IV U15063 ( .A(n14778), .Z(n14780) );
  NOR U15064 ( .A(n14779), .B(n14780), .Z(n14786) );
  XOR U15065 ( .A(n14781), .B(n14780), .Z(n15293) );
  XOR U15066 ( .A(n14783), .B(n14782), .Z(n15292) );
  IV U15067 ( .A(n15292), .Z(n14784) );
  NOR U15068 ( .A(n15293), .B(n14784), .Z(n14785) );
  NOR U15069 ( .A(n14786), .B(n14785), .Z(n14790) );
  XOR U15070 ( .A(n14788), .B(n14787), .Z(n14789) );
  NOR U15071 ( .A(n14790), .B(n14789), .Z(n14794) );
  XOR U15072 ( .A(n14790), .B(n14789), .Z(n15303) );
  IV U15073 ( .A(n15303), .Z(n14792) );
  NOR U15074 ( .A(n135), .B(n53), .Z(n14791) );
  IV U15075 ( .A(n14791), .Z(n15304) );
  NOR U15076 ( .A(n14792), .B(n15304), .Z(n14793) );
  NOR U15077 ( .A(n14794), .B(n14793), .Z(n14797) );
  NOR U15078 ( .A(n137), .B(n53), .Z(n14796) );
  IV U15079 ( .A(n14796), .Z(n14795) );
  NOR U15080 ( .A(n14797), .B(n14795), .Z(n14801) );
  XOR U15081 ( .A(n14797), .B(n14796), .Z(n15310) );
  XOR U15082 ( .A(n14799), .B(n14798), .Z(n15311) );
  NOR U15083 ( .A(n15310), .B(n15311), .Z(n14800) );
  NOR U15084 ( .A(n14801), .B(n14800), .Z(n14806) );
  NOR U15085 ( .A(n139), .B(n53), .Z(n14805) );
  IV U15086 ( .A(n14805), .Z(n14802) );
  NOR U15087 ( .A(n14806), .B(n14802), .Z(n14809) );
  XOR U15088 ( .A(n14804), .B(n14803), .Z(n15316) );
  IV U15089 ( .A(n15316), .Z(n14807) );
  XOR U15090 ( .A(n14806), .B(n14805), .Z(n15315) );
  NOR U15091 ( .A(n14807), .B(n15315), .Z(n14808) );
  NOR U15092 ( .A(n14809), .B(n14808), .Z(n14813) );
  XOR U15093 ( .A(n14811), .B(n14810), .Z(n14812) );
  NOR U15094 ( .A(n14813), .B(n14812), .Z(n14817) );
  XOR U15095 ( .A(n14813), .B(n14812), .Z(n14814) );
  IV U15096 ( .A(n14814), .Z(n15326) );
  NOR U15097 ( .A(n141), .B(n53), .Z(n15327) );
  IV U15098 ( .A(n15327), .Z(n14815) );
  NOR U15099 ( .A(n15326), .B(n14815), .Z(n14816) );
  NOR U15100 ( .A(n14817), .B(n14816), .Z(n15332) );
  XOR U15101 ( .A(n14819), .B(n14818), .Z(n15331) );
  NOR U15102 ( .A(n15332), .B(n15331), .Z(n14820) );
  NOR U15103 ( .A(n14821), .B(n14820), .Z(n14824) );
  NOR U15104 ( .A(n145), .B(n53), .Z(n14823) );
  IV U15105 ( .A(n14823), .Z(n14822) );
  NOR U15106 ( .A(n14824), .B(n14822), .Z(n14829) );
  XOR U15107 ( .A(n14824), .B(n14823), .Z(n15338) );
  XOR U15108 ( .A(n14826), .B(n14825), .Z(n15339) );
  IV U15109 ( .A(n15339), .Z(n14827) );
  NOR U15110 ( .A(n15338), .B(n14827), .Z(n14828) );
  NOR U15111 ( .A(n14829), .B(n14828), .Z(n14833) );
  XOR U15112 ( .A(n14831), .B(n14830), .Z(n14832) );
  NOR U15113 ( .A(n14833), .B(n14832), .Z(n14837) );
  XOR U15114 ( .A(n14833), .B(n14832), .Z(n14834) );
  IV U15115 ( .A(n14834), .Z(n15349) );
  NOR U15116 ( .A(n147), .B(n53), .Z(n15350) );
  IV U15117 ( .A(n15350), .Z(n14835) );
  NOR U15118 ( .A(n15349), .B(n14835), .Z(n14836) );
  NOR U15119 ( .A(n14837), .B(n14836), .Z(n14840) );
  NOR U15120 ( .A(n148), .B(n53), .Z(n14839) );
  IV U15121 ( .A(n14839), .Z(n14838) );
  NOR U15122 ( .A(n14840), .B(n14838), .Z(n14844) );
  XOR U15123 ( .A(n14840), .B(n14839), .Z(n15354) );
  XOR U15124 ( .A(n14842), .B(n14841), .Z(n15355) );
  NOR U15125 ( .A(n15354), .B(n15355), .Z(n14843) );
  NOR U15126 ( .A(n14844), .B(n14843), .Z(n14851) );
  NOR U15127 ( .A(n150), .B(n53), .Z(n14850) );
  IV U15128 ( .A(n14850), .Z(n14845) );
  NOR U15129 ( .A(n14851), .B(n14845), .Z(n14853) );
  XOR U15130 ( .A(n14847), .B(n14846), .Z(n14848) );
  XOR U15131 ( .A(n14849), .B(n14848), .Z(n15362) );
  XOR U15132 ( .A(n14851), .B(n14850), .Z(n15361) );
  NOR U15133 ( .A(n15362), .B(n15361), .Z(n14852) );
  NOR U15134 ( .A(n14853), .B(n14852), .Z(n14858) );
  XOR U15135 ( .A(n14855), .B(n14854), .Z(n14857) );
  IV U15136 ( .A(n14857), .Z(n14856) );
  NOR U15137 ( .A(n14858), .B(n14856), .Z(n14861) );
  XOR U15138 ( .A(n14858), .B(n14857), .Z(n15372) );
  NOR U15139 ( .A(n153), .B(n53), .Z(n15373) );
  IV U15140 ( .A(n15373), .Z(n14859) );
  NOR U15141 ( .A(n15372), .B(n14859), .Z(n14860) );
  NOR U15142 ( .A(n14861), .B(n14860), .Z(n14864) );
  NOR U15143 ( .A(n155), .B(n53), .Z(n14863) );
  IV U15144 ( .A(n14863), .Z(n14862) );
  NOR U15145 ( .A(n14864), .B(n14862), .Z(n14868) );
  XOR U15146 ( .A(n14864), .B(n14863), .Z(n15379) );
  XOR U15147 ( .A(n14866), .B(n14865), .Z(n15380) );
  NOR U15148 ( .A(n15379), .B(n15380), .Z(n14867) );
  NOR U15149 ( .A(n14868), .B(n14867), .Z(n14873) );
  NOR U15150 ( .A(n156), .B(n53), .Z(n14872) );
  IV U15151 ( .A(n14872), .Z(n14869) );
  NOR U15152 ( .A(n14873), .B(n14869), .Z(n14876) );
  XOR U15153 ( .A(n14871), .B(n14870), .Z(n15385) );
  IV U15154 ( .A(n15385), .Z(n14874) );
  XOR U15155 ( .A(n14873), .B(n14872), .Z(n15384) );
  NOR U15156 ( .A(n14874), .B(n15384), .Z(n14875) );
  NOR U15157 ( .A(n14876), .B(n14875), .Z(n14881) );
  XOR U15158 ( .A(n14878), .B(n14877), .Z(n14880) );
  IV U15159 ( .A(n14880), .Z(n14879) );
  NOR U15160 ( .A(n14881), .B(n14879), .Z(n14884) );
  XOR U15161 ( .A(n14881), .B(n14880), .Z(n15395) );
  NOR U15162 ( .A(n158), .B(n53), .Z(n15396) );
  IV U15163 ( .A(n15396), .Z(n14882) );
  NOR U15164 ( .A(n15395), .B(n14882), .Z(n14883) );
  NOR U15165 ( .A(n14884), .B(n14883), .Z(n15401) );
  XOR U15166 ( .A(n14886), .B(n14885), .Z(n15400) );
  NOR U15167 ( .A(n15401), .B(n15400), .Z(n14887) );
  NOR U15168 ( .A(n14888), .B(n14887), .Z(n14891) );
  NOR U15169 ( .A(n163), .B(n53), .Z(n14890) );
  IV U15170 ( .A(n14890), .Z(n14889) );
  NOR U15171 ( .A(n14891), .B(n14889), .Z(n14896) );
  XOR U15172 ( .A(n14891), .B(n14890), .Z(n15407) );
  XOR U15173 ( .A(n14893), .B(n14892), .Z(n15408) );
  IV U15174 ( .A(n15408), .Z(n14894) );
  NOR U15175 ( .A(n15407), .B(n14894), .Z(n14895) );
  NOR U15176 ( .A(n14896), .B(n14895), .Z(n14900) );
  XOR U15177 ( .A(n14898), .B(n14897), .Z(n14899) );
  NOR U15178 ( .A(n14900), .B(n14899), .Z(n14904) );
  XOR U15179 ( .A(n14900), .B(n14899), .Z(n15418) );
  IV U15180 ( .A(n15418), .Z(n14902) );
  NOR U15181 ( .A(n165), .B(n53), .Z(n14901) );
  IV U15182 ( .A(n14901), .Z(n15419) );
  NOR U15183 ( .A(n14902), .B(n15419), .Z(n14903) );
  NOR U15184 ( .A(n14904), .B(n14903), .Z(n15423) );
  XOR U15185 ( .A(n14906), .B(n14905), .Z(n15422) );
  NOR U15186 ( .A(n15423), .B(n15422), .Z(n14907) );
  NOR U15187 ( .A(n14908), .B(n14907), .Z(n15426) );
  XOR U15188 ( .A(n14910), .B(n14909), .Z(n15425) );
  NOR U15189 ( .A(n15426), .B(n15425), .Z(n28602) );
  IV U15190 ( .A(n28602), .Z(n31637) );
  XOR U15191 ( .A(n14912), .B(n14911), .Z(n31636) );
  IV U15192 ( .A(n31636), .Z(n14913) );
  NOR U15193 ( .A(n31637), .B(n14913), .Z(n31641) );
  NOR U15194 ( .A(n31643), .B(n31641), .Z(n14914) );
  NOR U15195 ( .A(n31645), .B(n14914), .Z(n28609) );
  NOR U15196 ( .A(n125), .B(n54), .Z(n15245) );
  XOR U15197 ( .A(n14916), .B(n14915), .Z(n15224) );
  XOR U15198 ( .A(n14918), .B(n14917), .Z(n14919) );
  XOR U15199 ( .A(n14920), .B(n14919), .Z(n15735) );
  IV U15200 ( .A(n15735), .Z(n14921) );
  NOR U15201 ( .A(n79), .B(n54), .Z(n14922) );
  NOR U15202 ( .A(n14921), .B(n14922), .Z(n15223) );
  IV U15203 ( .A(n14922), .Z(n15734) );
  NOR U15204 ( .A(n15735), .B(n15734), .Z(n15221) );
  NOR U15205 ( .A(n80), .B(n54), .Z(n14925) );
  XOR U15206 ( .A(n14924), .B(n14923), .Z(n14926) );
  NOR U15207 ( .A(n14925), .B(n14926), .Z(n15209) );
  IV U15208 ( .A(n14925), .Z(n15721) );
  IV U15209 ( .A(n14926), .Z(n15720) );
  NOR U15210 ( .A(n15721), .B(n15720), .Z(n15207) );
  XOR U15211 ( .A(n14928), .B(n14927), .Z(n14929) );
  IV U15212 ( .A(n14929), .Z(n15192) );
  NOR U15213 ( .A(n81), .B(n54), .Z(n15193) );
  IV U15214 ( .A(n15193), .Z(n14930) );
  NOR U15215 ( .A(n15192), .B(n14930), .Z(n15196) );
  NOR U15216 ( .A(n115), .B(n54), .Z(n15187) );
  XOR U15217 ( .A(n14932), .B(n14931), .Z(n14933) );
  XOR U15218 ( .A(n14934), .B(n14933), .Z(n15188) );
  NOR U15219 ( .A(n15187), .B(n15188), .Z(n15191) );
  NOR U15220 ( .A(n82), .B(n54), .Z(n15183) );
  XOR U15221 ( .A(n14936), .B(n14935), .Z(n15182) );
  NOR U15222 ( .A(n15183), .B(n15182), .Z(n15186) );
  NOR U15223 ( .A(n83), .B(n54), .Z(n14940) );
  IV U15224 ( .A(n14940), .Z(n15688) );
  XOR U15225 ( .A(n14938), .B(n14937), .Z(n14939) );
  IV U15226 ( .A(n14939), .Z(n15687) );
  NOR U15227 ( .A(n15688), .B(n15687), .Z(n15173) );
  NOR U15228 ( .A(n14940), .B(n14939), .Z(n15171) );
  NOR U15229 ( .A(n113), .B(n54), .Z(n14941) );
  IV U15230 ( .A(n14941), .Z(n15166) );
  NOR U15231 ( .A(n84), .B(n54), .Z(n15160) );
  XOR U15232 ( .A(n14943), .B(n14942), .Z(n15159) );
  NOR U15233 ( .A(n15160), .B(n15159), .Z(n15163) );
  XOR U15234 ( .A(n14945), .B(n14944), .Z(n15155) );
  NOR U15235 ( .A(n112), .B(n54), .Z(n15154) );
  IV U15236 ( .A(n15154), .Z(n14946) );
  NOR U15237 ( .A(n15155), .B(n14946), .Z(n15157) );
  IV U15238 ( .A(n14947), .Z(n14949) );
  XOR U15239 ( .A(n14949), .B(n14948), .Z(n15150) );
  NOR U15240 ( .A(n85), .B(n54), .Z(n15151) );
  IV U15241 ( .A(n15151), .Z(n14950) );
  NOR U15242 ( .A(n15150), .B(n14950), .Z(n15153) );
  XOR U15243 ( .A(n14952), .B(n14951), .Z(n15135) );
  NOR U15244 ( .A(n86), .B(n54), .Z(n15136) );
  NOR U15245 ( .A(n15135), .B(n15136), .Z(n15140) );
  XOR U15246 ( .A(n14954), .B(n14953), .Z(n15131) );
  IV U15247 ( .A(n15131), .Z(n14956) );
  NOR U15248 ( .A(n110), .B(n54), .Z(n14955) );
  IV U15249 ( .A(n14955), .Z(n15132) );
  NOR U15250 ( .A(n14956), .B(n15132), .Z(n15134) );
  NOR U15251 ( .A(n109), .B(n54), .Z(n15126) );
  XOR U15252 ( .A(n14958), .B(n14957), .Z(n15125) );
  NOR U15253 ( .A(n15126), .B(n15125), .Z(n15129) );
  XOR U15254 ( .A(n14960), .B(n14959), .Z(n14961) );
  XOR U15255 ( .A(n14962), .B(n14961), .Z(n15120) );
  NOR U15256 ( .A(n108), .B(n54), .Z(n15119) );
  IV U15257 ( .A(n15119), .Z(n14963) );
  NOR U15258 ( .A(n15120), .B(n14963), .Z(n15123) );
  NOR U15259 ( .A(n87), .B(n54), .Z(n14967) );
  XOR U15260 ( .A(n14965), .B(n14964), .Z(n14966) );
  NOR U15261 ( .A(n14967), .B(n14966), .Z(n15118) );
  XOR U15262 ( .A(n14967), .B(n14966), .Z(n14968) );
  IV U15263 ( .A(n14968), .Z(n15481) );
  XOR U15264 ( .A(n14970), .B(n14969), .Z(n15113) );
  NOR U15265 ( .A(n107), .B(n54), .Z(n15112) );
  IV U15266 ( .A(n15112), .Z(n14971) );
  NOR U15267 ( .A(n15113), .B(n14971), .Z(n15115) );
  NOR U15268 ( .A(n88), .B(n54), .Z(n15107) );
  XOR U15269 ( .A(n14973), .B(n14972), .Z(n15106) );
  NOR U15270 ( .A(n15107), .B(n15106), .Z(n15110) );
  IV U15271 ( .A(n14974), .Z(n14976) );
  XOR U15272 ( .A(n14976), .B(n14975), .Z(n15100) );
  NOR U15273 ( .A(n106), .B(n54), .Z(n15101) );
  IV U15274 ( .A(n15101), .Z(n14977) );
  NOR U15275 ( .A(n15100), .B(n14977), .Z(n15104) );
  NOR U15276 ( .A(n105), .B(n54), .Z(n15096) );
  XOR U15277 ( .A(n14979), .B(n14978), .Z(n15095) );
  NOR U15278 ( .A(n15096), .B(n15095), .Z(n15099) );
  IV U15279 ( .A(n14980), .Z(n14982) );
  XOR U15280 ( .A(n14982), .B(n14981), .Z(n15090) );
  NOR U15281 ( .A(n104), .B(n54), .Z(n15091) );
  IV U15282 ( .A(n15091), .Z(n14983) );
  NOR U15283 ( .A(n15090), .B(n14983), .Z(n15093) );
  IV U15284 ( .A(n14984), .Z(n14986) );
  XOR U15285 ( .A(n14986), .B(n14985), .Z(n15086) );
  NOR U15286 ( .A(n89), .B(n54), .Z(n15087) );
  IV U15287 ( .A(n15087), .Z(n14987) );
  NOR U15288 ( .A(n15086), .B(n14987), .Z(n15089) );
  IV U15289 ( .A(n14988), .Z(n14990) );
  XOR U15290 ( .A(n14990), .B(n14989), .Z(n15082) );
  NOR U15291 ( .A(n103), .B(n54), .Z(n15083) );
  IV U15292 ( .A(n15083), .Z(n14991) );
  NOR U15293 ( .A(n15082), .B(n14991), .Z(n15085) );
  XOR U15294 ( .A(n14993), .B(n14992), .Z(n15078) );
  IV U15295 ( .A(n15078), .Z(n14995) );
  NOR U15296 ( .A(n90), .B(n54), .Z(n14994) );
  IV U15297 ( .A(n14994), .Z(n15079) );
  NOR U15298 ( .A(n14995), .B(n15079), .Z(n15081) );
  IV U15299 ( .A(n14996), .Z(n14998) );
  XOR U15300 ( .A(n14998), .B(n14997), .Z(n15074) );
  NOR U15301 ( .A(n102), .B(n54), .Z(n15075) );
  IV U15302 ( .A(n15075), .Z(n14999) );
  NOR U15303 ( .A(n15074), .B(n14999), .Z(n15077) );
  IV U15304 ( .A(n15000), .Z(n15002) );
  XOR U15305 ( .A(n15002), .B(n15001), .Z(n15070) );
  NOR U15306 ( .A(n101), .B(n54), .Z(n15071) );
  IV U15307 ( .A(n15071), .Z(n15003) );
  NOR U15308 ( .A(n15070), .B(n15003), .Z(n15073) );
  IV U15309 ( .A(n15004), .Z(n15006) );
  XOR U15310 ( .A(n15006), .B(n15005), .Z(n15066) );
  NOR U15311 ( .A(n100), .B(n54), .Z(n15067) );
  IV U15312 ( .A(n15067), .Z(n15007) );
  NOR U15313 ( .A(n15066), .B(n15007), .Z(n15069) );
  IV U15314 ( .A(n15008), .Z(n15010) );
  XOR U15315 ( .A(n15010), .B(n15009), .Z(n15062) );
  NOR U15316 ( .A(n99), .B(n54), .Z(n15063) );
  IV U15317 ( .A(n15063), .Z(n15011) );
  NOR U15318 ( .A(n15062), .B(n15011), .Z(n15065) );
  IV U15319 ( .A(n15012), .Z(n15014) );
  XOR U15320 ( .A(n15014), .B(n15013), .Z(n15058) );
  NOR U15321 ( .A(n98), .B(n54), .Z(n15059) );
  IV U15322 ( .A(n15059), .Z(n15015) );
  NOR U15323 ( .A(n15058), .B(n15015), .Z(n15061) );
  XOR U15324 ( .A(n15017), .B(n15016), .Z(n15054) );
  NOR U15325 ( .A(n91), .B(n54), .Z(n15055) );
  IV U15326 ( .A(n15055), .Z(n15018) );
  NOR U15327 ( .A(n15054), .B(n15018), .Z(n15057) );
  XOR U15328 ( .A(n15020), .B(n15019), .Z(n15042) );
  IV U15329 ( .A(n15042), .Z(n15022) );
  NOR U15330 ( .A(n96), .B(n54), .Z(n15021) );
  IV U15331 ( .A(n15021), .Z(n15043) );
  NOR U15332 ( .A(n15022), .B(n15043), .Z(n15045) );
  NOR U15333 ( .A(n95), .B(n54), .Z(n15039) );
  IV U15334 ( .A(n15039), .Z(n15025) );
  XOR U15335 ( .A(n15024), .B(n15023), .Z(n15038) );
  NOR U15336 ( .A(n15025), .B(n15038), .Z(n15041) );
  NOR U15337 ( .A(n93), .B(n54), .Z(n16050) );
  IV U15338 ( .A(n16050), .Z(n15026) );
  NOR U15339 ( .A(n53), .B(n168), .Z(n15034) );
  IV U15340 ( .A(n15034), .Z(n15029) );
  NOR U15341 ( .A(n15026), .B(n15029), .Z(n15027) );
  IV U15342 ( .A(n15027), .Z(n15028) );
  NOR U15343 ( .A(n94), .B(n15028), .Z(n15037) );
  NOR U15344 ( .A(n15029), .B(n93), .Z(n15030) );
  XOR U15345 ( .A(n94), .B(n15030), .Z(n15031) );
  NOR U15346 ( .A(n54), .B(n15031), .Z(n15032) );
  IV U15347 ( .A(n15032), .Z(n15538) );
  XOR U15348 ( .A(n15034), .B(n15033), .Z(n15537) );
  IV U15349 ( .A(n15537), .Z(n15035) );
  NOR U15350 ( .A(n15538), .B(n15035), .Z(n15036) );
  NOR U15351 ( .A(n15037), .B(n15036), .Z(n15533) );
  XOR U15352 ( .A(n15039), .B(n15038), .Z(n15534) );
  NOR U15353 ( .A(n15533), .B(n15534), .Z(n15040) );
  NOR U15354 ( .A(n15041), .B(n15040), .Z(n15561) );
  XOR U15355 ( .A(n15043), .B(n15042), .Z(n15560) );
  NOR U15356 ( .A(n15561), .B(n15560), .Z(n15044) );
  NOR U15357 ( .A(n15045), .B(n15044), .Z(n15050) );
  XOR U15358 ( .A(n15047), .B(n15046), .Z(n15049) );
  IV U15359 ( .A(n15049), .Z(n15048) );
  NOR U15360 ( .A(n15050), .B(n15048), .Z(n15053) );
  XOR U15361 ( .A(n15050), .B(n15049), .Z(n15530) );
  NOR U15362 ( .A(n97), .B(n54), .Z(n15531) );
  IV U15363 ( .A(n15531), .Z(n15051) );
  NOR U15364 ( .A(n15530), .B(n15051), .Z(n15052) );
  NOR U15365 ( .A(n15053), .B(n15052), .Z(n15526) );
  XOR U15366 ( .A(n15055), .B(n15054), .Z(n15527) );
  NOR U15367 ( .A(n15526), .B(n15527), .Z(n15056) );
  NOR U15368 ( .A(n15057), .B(n15056), .Z(n15522) );
  XOR U15369 ( .A(n15059), .B(n15058), .Z(n15523) );
  NOR U15370 ( .A(n15522), .B(n15523), .Z(n15060) );
  NOR U15371 ( .A(n15061), .B(n15060), .Z(n15518) );
  XOR U15372 ( .A(n15063), .B(n15062), .Z(n15519) );
  NOR U15373 ( .A(n15518), .B(n15519), .Z(n15064) );
  NOR U15374 ( .A(n15065), .B(n15064), .Z(n15514) );
  XOR U15375 ( .A(n15067), .B(n15066), .Z(n15515) );
  NOR U15376 ( .A(n15514), .B(n15515), .Z(n15068) );
  NOR U15377 ( .A(n15069), .B(n15068), .Z(n15510) );
  XOR U15378 ( .A(n15071), .B(n15070), .Z(n15511) );
  NOR U15379 ( .A(n15510), .B(n15511), .Z(n15072) );
  NOR U15380 ( .A(n15073), .B(n15072), .Z(n15506) );
  XOR U15381 ( .A(n15075), .B(n15074), .Z(n15507) );
  NOR U15382 ( .A(n15506), .B(n15507), .Z(n15076) );
  NOR U15383 ( .A(n15077), .B(n15076), .Z(n15597) );
  XOR U15384 ( .A(n15079), .B(n15078), .Z(n15596) );
  NOR U15385 ( .A(n15597), .B(n15596), .Z(n15080) );
  NOR U15386 ( .A(n15081), .B(n15080), .Z(n15502) );
  XOR U15387 ( .A(n15083), .B(n15082), .Z(n15503) );
  NOR U15388 ( .A(n15502), .B(n15503), .Z(n15084) );
  NOR U15389 ( .A(n15085), .B(n15084), .Z(n15498) );
  XOR U15390 ( .A(n15087), .B(n15086), .Z(n15499) );
  NOR U15391 ( .A(n15498), .B(n15499), .Z(n15088) );
  NOR U15392 ( .A(n15089), .B(n15088), .Z(n15494) );
  XOR U15393 ( .A(n15091), .B(n15090), .Z(n15495) );
  NOR U15394 ( .A(n15494), .B(n15495), .Z(n15092) );
  NOR U15395 ( .A(n15093), .B(n15092), .Z(n15094) );
  IV U15396 ( .A(n15094), .Z(n15492) );
  XOR U15397 ( .A(n15096), .B(n15095), .Z(n15097) );
  IV U15398 ( .A(n15097), .Z(n15491) );
  NOR U15399 ( .A(n15492), .B(n15491), .Z(n15098) );
  NOR U15400 ( .A(n15099), .B(n15098), .Z(n15489) );
  IV U15401 ( .A(n15489), .Z(n15102) );
  XOR U15402 ( .A(n15101), .B(n15100), .Z(n15488) );
  NOR U15403 ( .A(n15102), .B(n15488), .Z(n15103) );
  NOR U15404 ( .A(n15104), .B(n15103), .Z(n15105) );
  IV U15405 ( .A(n15105), .Z(n15486) );
  XOR U15406 ( .A(n15107), .B(n15106), .Z(n15108) );
  IV U15407 ( .A(n15108), .Z(n15485) );
  NOR U15408 ( .A(n15486), .B(n15485), .Z(n15109) );
  NOR U15409 ( .A(n15110), .B(n15109), .Z(n15111) );
  IV U15410 ( .A(n15111), .Z(n15484) );
  XOR U15411 ( .A(n15113), .B(n15112), .Z(n15483) );
  NOR U15412 ( .A(n15484), .B(n15483), .Z(n15114) );
  NOR U15413 ( .A(n15115), .B(n15114), .Z(n15116) );
  IV U15414 ( .A(n15116), .Z(n15480) );
  NOR U15415 ( .A(n15481), .B(n15480), .Z(n15117) );
  NOR U15416 ( .A(n15118), .B(n15117), .Z(n15478) );
  IV U15417 ( .A(n15478), .Z(n15121) );
  XOR U15418 ( .A(n15120), .B(n15119), .Z(n15477) );
  NOR U15419 ( .A(n15121), .B(n15477), .Z(n15122) );
  NOR U15420 ( .A(n15123), .B(n15122), .Z(n15124) );
  IV U15421 ( .A(n15124), .Z(n15475) );
  XOR U15422 ( .A(n15126), .B(n15125), .Z(n15127) );
  IV U15423 ( .A(n15127), .Z(n15474) );
  NOR U15424 ( .A(n15475), .B(n15474), .Z(n15128) );
  NOR U15425 ( .A(n15129), .B(n15128), .Z(n15130) );
  IV U15426 ( .A(n15130), .Z(n15473) );
  XOR U15427 ( .A(n15132), .B(n15131), .Z(n15472) );
  NOR U15428 ( .A(n15473), .B(n15472), .Z(n15133) );
  NOR U15429 ( .A(n15134), .B(n15133), .Z(n15468) );
  IV U15430 ( .A(n15468), .Z(n15138) );
  IV U15431 ( .A(n15135), .Z(n15466) );
  IV U15432 ( .A(n15136), .Z(n15465) );
  NOR U15433 ( .A(n15466), .B(n15465), .Z(n15137) );
  NOR U15434 ( .A(n15138), .B(n15137), .Z(n15139) );
  NOR U15435 ( .A(n15140), .B(n15139), .Z(n15146) );
  IV U15436 ( .A(n15146), .Z(n15144) );
  IV U15437 ( .A(n15141), .Z(n15143) );
  XOR U15438 ( .A(n15143), .B(n15142), .Z(n15145) );
  NOR U15439 ( .A(n15144), .B(n15145), .Z(n15149) );
  XOR U15440 ( .A(n15146), .B(n15145), .Z(n15463) );
  NOR U15441 ( .A(n111), .B(n54), .Z(n15147) );
  IV U15442 ( .A(n15147), .Z(n15464) );
  NOR U15443 ( .A(n15463), .B(n15464), .Z(n15148) );
  NOR U15444 ( .A(n15149), .B(n15148), .Z(n15662) );
  XOR U15445 ( .A(n15151), .B(n15150), .Z(n15663) );
  NOR U15446 ( .A(n15662), .B(n15663), .Z(n15152) );
  NOR U15447 ( .A(n15153), .B(n15152), .Z(n15460) );
  XOR U15448 ( .A(n15155), .B(n15154), .Z(n15459) );
  NOR U15449 ( .A(n15460), .B(n15459), .Z(n15156) );
  NOR U15450 ( .A(n15157), .B(n15156), .Z(n15158) );
  IV U15451 ( .A(n15158), .Z(n15676) );
  XOR U15452 ( .A(n15160), .B(n15159), .Z(n15161) );
  IV U15453 ( .A(n15161), .Z(n15675) );
  NOR U15454 ( .A(n15676), .B(n15675), .Z(n15162) );
  NOR U15455 ( .A(n15163), .B(n15162), .Z(n15165) );
  IV U15456 ( .A(n15165), .Z(n15164) );
  NOR U15457 ( .A(n15166), .B(n15164), .Z(n15170) );
  XOR U15458 ( .A(n15166), .B(n15165), .Z(n15456) );
  XOR U15459 ( .A(n15168), .B(n15167), .Z(n15455) );
  NOR U15460 ( .A(n15456), .B(n15455), .Z(n15169) );
  NOR U15461 ( .A(n15170), .B(n15169), .Z(n15690) );
  NOR U15462 ( .A(n15171), .B(n15690), .Z(n15172) );
  NOR U15463 ( .A(n15173), .B(n15172), .Z(n15177) );
  NOR U15464 ( .A(n114), .B(n54), .Z(n15178) );
  IV U15465 ( .A(n15178), .Z(n15174) );
  NOR U15466 ( .A(n15177), .B(n15174), .Z(n15180) );
  XOR U15467 ( .A(n15176), .B(n15175), .Z(n15452) );
  XOR U15468 ( .A(n15178), .B(n15177), .Z(n15451) );
  NOR U15469 ( .A(n15452), .B(n15451), .Z(n15179) );
  NOR U15470 ( .A(n15180), .B(n15179), .Z(n15181) );
  IV U15471 ( .A(n15181), .Z(n15700) );
  XOR U15472 ( .A(n15183), .B(n15182), .Z(n15184) );
  IV U15473 ( .A(n15184), .Z(n15699) );
  NOR U15474 ( .A(n15700), .B(n15699), .Z(n15185) );
  NOR U15475 ( .A(n15186), .B(n15185), .Z(n15449) );
  XOR U15476 ( .A(n15188), .B(n15187), .Z(n15450) );
  IV U15477 ( .A(n15450), .Z(n15189) );
  NOR U15478 ( .A(n15449), .B(n15189), .Z(n15190) );
  NOR U15479 ( .A(n15191), .B(n15190), .Z(n15447) );
  IV U15480 ( .A(n15447), .Z(n15194) );
  XOR U15481 ( .A(n15193), .B(n15192), .Z(n15446) );
  NOR U15482 ( .A(n15194), .B(n15446), .Z(n15195) );
  NOR U15483 ( .A(n15196), .B(n15195), .Z(n15202) );
  NOR U15484 ( .A(n116), .B(n54), .Z(n15203) );
  IV U15485 ( .A(n15203), .Z(n15197) );
  NOR U15486 ( .A(n15202), .B(n15197), .Z(n15205) );
  XOR U15487 ( .A(n15199), .B(n15198), .Z(n15200) );
  XOR U15488 ( .A(n15201), .B(n15200), .Z(n15443) );
  XOR U15489 ( .A(n15203), .B(n15202), .Z(n15442) );
  NOR U15490 ( .A(n15443), .B(n15442), .Z(n15204) );
  NOR U15491 ( .A(n15205), .B(n15204), .Z(n15723) );
  IV U15492 ( .A(n15723), .Z(n15206) );
  NOR U15493 ( .A(n15207), .B(n15206), .Z(n15208) );
  NOR U15494 ( .A(n15209), .B(n15208), .Z(n15210) );
  IV U15495 ( .A(n15210), .Z(n15217) );
  NOR U15496 ( .A(n117), .B(n54), .Z(n15216) );
  IV U15497 ( .A(n15216), .Z(n15211) );
  NOR U15498 ( .A(n15217), .B(n15211), .Z(n15219) );
  XOR U15499 ( .A(n15213), .B(n15212), .Z(n15214) );
  XOR U15500 ( .A(n15215), .B(n15214), .Z(n15438) );
  XOR U15501 ( .A(n15217), .B(n15216), .Z(n15439) );
  NOR U15502 ( .A(n15438), .B(n15439), .Z(n15218) );
  NOR U15503 ( .A(n15219), .B(n15218), .Z(n15737) );
  IV U15504 ( .A(n15737), .Z(n15220) );
  NOR U15505 ( .A(n15221), .B(n15220), .Z(n15222) );
  NOR U15506 ( .A(n15223), .B(n15222), .Z(n15745) );
  NOR U15507 ( .A(n15224), .B(n15745), .Z(n15228) );
  IV U15508 ( .A(n15224), .Z(n15747) );
  IV U15509 ( .A(n15745), .Z(n15225) );
  NOR U15510 ( .A(n15747), .B(n15225), .Z(n15226) );
  NOR U15511 ( .A(n119), .B(n54), .Z(n15744) );
  NOR U15512 ( .A(n15226), .B(n15744), .Z(n15227) );
  NOR U15513 ( .A(n15228), .B(n15227), .Z(n15230) );
  IV U15514 ( .A(n15230), .Z(n15753) );
  NOR U15515 ( .A(n120), .B(n54), .Z(n15229) );
  IV U15516 ( .A(n15229), .Z(n15752) );
  NOR U15517 ( .A(n15753), .B(n15752), .Z(n15235) );
  NOR U15518 ( .A(n15230), .B(n15229), .Z(n15233) );
  XOR U15519 ( .A(n15232), .B(n15231), .Z(n15755) );
  NOR U15520 ( .A(n15233), .B(n15755), .Z(n15234) );
  NOR U15521 ( .A(n15235), .B(n15234), .Z(n15242) );
  NOR U15522 ( .A(n123), .B(n54), .Z(n15241) );
  IV U15523 ( .A(n15241), .Z(n15236) );
  NOR U15524 ( .A(n15242), .B(n15236), .Z(n15244) );
  XOR U15525 ( .A(n15238), .B(n15237), .Z(n15239) );
  XOR U15526 ( .A(n15240), .B(n15239), .Z(n15437) );
  XOR U15527 ( .A(n15242), .B(n15241), .Z(n15436) );
  NOR U15528 ( .A(n15437), .B(n15436), .Z(n15243) );
  NOR U15529 ( .A(n15244), .B(n15243), .Z(n15246) );
  IV U15530 ( .A(n15246), .Z(n15765) );
  NOR U15531 ( .A(n15245), .B(n15765), .Z(n15253) );
  IV U15532 ( .A(n15245), .Z(n15766) );
  NOR U15533 ( .A(n15246), .B(n15766), .Z(n15251) );
  XOR U15534 ( .A(n15248), .B(n15247), .Z(n15249) );
  XOR U15535 ( .A(n15250), .B(n15249), .Z(n15768) );
  NOR U15536 ( .A(n15251), .B(n15768), .Z(n15252) );
  NOR U15537 ( .A(n15253), .B(n15252), .Z(n15254) );
  IV U15538 ( .A(n15254), .Z(n15261) );
  NOR U15539 ( .A(n126), .B(n54), .Z(n15260) );
  IV U15540 ( .A(n15260), .Z(n15255) );
  NOR U15541 ( .A(n15261), .B(n15255), .Z(n15264) );
  XOR U15542 ( .A(n15257), .B(n15256), .Z(n15258) );
  XOR U15543 ( .A(n15259), .B(n15258), .Z(n15779) );
  IV U15544 ( .A(n15779), .Z(n15262) );
  XOR U15545 ( .A(n15261), .B(n15260), .Z(n15780) );
  NOR U15546 ( .A(n15262), .B(n15780), .Z(n15263) );
  NOR U15547 ( .A(n15264), .B(n15263), .Z(n15268) );
  XOR U15548 ( .A(n15266), .B(n15265), .Z(n15267) );
  NOR U15549 ( .A(n15268), .B(n15267), .Z(n15272) );
  XOR U15550 ( .A(n15268), .B(n15267), .Z(n15434) );
  IV U15551 ( .A(n15434), .Z(n15270) );
  NOR U15552 ( .A(n128), .B(n54), .Z(n15269) );
  IV U15553 ( .A(n15269), .Z(n15433) );
  NOR U15554 ( .A(n15270), .B(n15433), .Z(n15271) );
  NOR U15555 ( .A(n15272), .B(n15271), .Z(n15279) );
  NOR U15556 ( .A(n131), .B(n54), .Z(n15278) );
  IV U15557 ( .A(n15278), .Z(n15273) );
  NOR U15558 ( .A(n15279), .B(n15273), .Z(n15282) );
  XOR U15559 ( .A(n15275), .B(n15274), .Z(n15276) );
  XOR U15560 ( .A(n15277), .B(n15276), .Z(n15787) );
  IV U15561 ( .A(n15787), .Z(n15280) );
  XOR U15562 ( .A(n15279), .B(n15278), .Z(n15786) );
  NOR U15563 ( .A(n15280), .B(n15786), .Z(n15281) );
  NOR U15564 ( .A(n15282), .B(n15281), .Z(n15289) );
  NOR U15565 ( .A(n133), .B(n54), .Z(n15288) );
  IV U15566 ( .A(n15288), .Z(n15283) );
  NOR U15567 ( .A(n15289), .B(n15283), .Z(n15291) );
  XOR U15568 ( .A(n15285), .B(n15284), .Z(n15286) );
  XOR U15569 ( .A(n15287), .B(n15286), .Z(n15791) );
  XOR U15570 ( .A(n15289), .B(n15288), .Z(n15790) );
  NOR U15571 ( .A(n15791), .B(n15790), .Z(n15290) );
  NOR U15572 ( .A(n15291), .B(n15290), .Z(n15294) );
  XOR U15573 ( .A(n15293), .B(n15292), .Z(n15295) );
  NOR U15574 ( .A(n15294), .B(n15295), .Z(n15299) );
  IV U15575 ( .A(n15294), .Z(n15296) );
  XOR U15576 ( .A(n15296), .B(n15295), .Z(n15430) );
  NOR U15577 ( .A(n135), .B(n54), .Z(n15431) );
  IV U15578 ( .A(n15431), .Z(n15297) );
  NOR U15579 ( .A(n15430), .B(n15297), .Z(n15298) );
  NOR U15580 ( .A(n15299), .B(n15298), .Z(n15302) );
  NOR U15581 ( .A(n137), .B(n54), .Z(n15301) );
  IV U15582 ( .A(n15301), .Z(n15300) );
  NOR U15583 ( .A(n15302), .B(n15300), .Z(n15306) );
  XOR U15584 ( .A(n15302), .B(n15301), .Z(n15805) );
  XOR U15585 ( .A(n15304), .B(n15303), .Z(n15806) );
  NOR U15586 ( .A(n15805), .B(n15806), .Z(n15305) );
  NOR U15587 ( .A(n15306), .B(n15305), .Z(n15309) );
  NOR U15588 ( .A(n139), .B(n54), .Z(n15308) );
  IV U15589 ( .A(n15308), .Z(n15307) );
  NOR U15590 ( .A(n15309), .B(n15307), .Z(n15314) );
  XOR U15591 ( .A(n15309), .B(n15308), .Z(n15810) );
  XOR U15592 ( .A(n15311), .B(n15310), .Z(n15811) );
  IV U15593 ( .A(n15811), .Z(n15312) );
  NOR U15594 ( .A(n15810), .B(n15312), .Z(n15313) );
  NOR U15595 ( .A(n15314), .B(n15313), .Z(n15318) );
  XOR U15596 ( .A(n15316), .B(n15315), .Z(n15317) );
  NOR U15597 ( .A(n15318), .B(n15317), .Z(n15322) );
  XOR U15598 ( .A(n15318), .B(n15317), .Z(n15427) );
  IV U15599 ( .A(n15427), .Z(n15320) );
  NOR U15600 ( .A(n141), .B(n54), .Z(n15319) );
  IV U15601 ( .A(n15319), .Z(n15428) );
  NOR U15602 ( .A(n15320), .B(n15428), .Z(n15321) );
  NOR U15603 ( .A(n15322), .B(n15321), .Z(n15325) );
  NOR U15604 ( .A(n143), .B(n54), .Z(n15324) );
  IV U15605 ( .A(n15324), .Z(n15323) );
  NOR U15606 ( .A(n15325), .B(n15323), .Z(n15329) );
  XOR U15607 ( .A(n15325), .B(n15324), .Z(n15823) );
  XOR U15608 ( .A(n15327), .B(n15326), .Z(n15824) );
  NOR U15609 ( .A(n15823), .B(n15824), .Z(n15328) );
  NOR U15610 ( .A(n15329), .B(n15328), .Z(n15334) );
  NOR U15611 ( .A(n145), .B(n54), .Z(n15333) );
  IV U15612 ( .A(n15333), .Z(n15330) );
  NOR U15613 ( .A(n15334), .B(n15330), .Z(n15337) );
  XOR U15614 ( .A(n15332), .B(n15331), .Z(n15831) );
  IV U15615 ( .A(n15831), .Z(n15335) );
  XOR U15616 ( .A(n15334), .B(n15333), .Z(n15830) );
  NOR U15617 ( .A(n15335), .B(n15830), .Z(n15336) );
  NOR U15618 ( .A(n15337), .B(n15336), .Z(n15341) );
  XOR U15619 ( .A(n15339), .B(n15338), .Z(n15340) );
  NOR U15620 ( .A(n15341), .B(n15340), .Z(n15345) );
  XOR U15621 ( .A(n15341), .B(n15340), .Z(n15841) );
  IV U15622 ( .A(n15841), .Z(n15343) );
  NOR U15623 ( .A(n147), .B(n54), .Z(n15342) );
  IV U15624 ( .A(n15342), .Z(n15842) );
  NOR U15625 ( .A(n15343), .B(n15842), .Z(n15344) );
  NOR U15626 ( .A(n15345), .B(n15344), .Z(n15348) );
  NOR U15627 ( .A(n148), .B(n54), .Z(n15347) );
  IV U15628 ( .A(n15347), .Z(n15346) );
  NOR U15629 ( .A(n15348), .B(n15346), .Z(n15352) );
  XOR U15630 ( .A(n15348), .B(n15347), .Z(n15846) );
  XOR U15631 ( .A(n15350), .B(n15349), .Z(n15847) );
  NOR U15632 ( .A(n15846), .B(n15847), .Z(n15351) );
  NOR U15633 ( .A(n15352), .B(n15351), .Z(n15357) );
  NOR U15634 ( .A(n150), .B(n54), .Z(n15356) );
  IV U15635 ( .A(n15356), .Z(n15353) );
  NOR U15636 ( .A(n15357), .B(n15353), .Z(n15360) );
  XOR U15637 ( .A(n15355), .B(n15354), .Z(n15854) );
  IV U15638 ( .A(n15854), .Z(n15358) );
  XOR U15639 ( .A(n15357), .B(n15356), .Z(n15853) );
  NOR U15640 ( .A(n15358), .B(n15853), .Z(n15359) );
  NOR U15641 ( .A(n15360), .B(n15359), .Z(n15365) );
  XOR U15642 ( .A(n15362), .B(n15361), .Z(n15364) );
  IV U15643 ( .A(n15364), .Z(n15363) );
  NOR U15644 ( .A(n15365), .B(n15363), .Z(n15368) );
  XOR U15645 ( .A(n15365), .B(n15364), .Z(n15861) );
  NOR U15646 ( .A(n153), .B(n54), .Z(n15862) );
  IV U15647 ( .A(n15862), .Z(n15366) );
  NOR U15648 ( .A(n15861), .B(n15366), .Z(n15367) );
  NOR U15649 ( .A(n15368), .B(n15367), .Z(n15371) );
  NOR U15650 ( .A(n155), .B(n54), .Z(n15370) );
  IV U15651 ( .A(n15370), .Z(n15369) );
  NOR U15652 ( .A(n15371), .B(n15369), .Z(n15375) );
  XOR U15653 ( .A(n15371), .B(n15370), .Z(n15870) );
  XOR U15654 ( .A(n15373), .B(n15372), .Z(n15871) );
  NOR U15655 ( .A(n15870), .B(n15871), .Z(n15374) );
  NOR U15656 ( .A(n15375), .B(n15374), .Z(n15378) );
  NOR U15657 ( .A(n156), .B(n54), .Z(n15377) );
  IV U15658 ( .A(n15377), .Z(n15376) );
  NOR U15659 ( .A(n15378), .B(n15376), .Z(n15383) );
  XOR U15660 ( .A(n15378), .B(n15377), .Z(n15877) );
  XOR U15661 ( .A(n15380), .B(n15379), .Z(n15878) );
  IV U15662 ( .A(n15878), .Z(n15381) );
  NOR U15663 ( .A(n15877), .B(n15381), .Z(n15382) );
  NOR U15664 ( .A(n15383), .B(n15382), .Z(n15387) );
  XOR U15665 ( .A(n15385), .B(n15384), .Z(n15386) );
  NOR U15666 ( .A(n15387), .B(n15386), .Z(n15391) );
  XOR U15667 ( .A(n15387), .B(n15386), .Z(n15388) );
  IV U15668 ( .A(n15388), .Z(n15887) );
  NOR U15669 ( .A(n158), .B(n54), .Z(n15389) );
  IV U15670 ( .A(n15389), .Z(n15886) );
  NOR U15671 ( .A(n15887), .B(n15886), .Z(n15390) );
  NOR U15672 ( .A(n15391), .B(n15390), .Z(n15394) );
  NOR U15673 ( .A(n161), .B(n54), .Z(n15393) );
  IV U15674 ( .A(n15393), .Z(n15392) );
  NOR U15675 ( .A(n15394), .B(n15392), .Z(n15398) );
  XOR U15676 ( .A(n15394), .B(n15393), .Z(n15896) );
  XOR U15677 ( .A(n15396), .B(n15395), .Z(n15897) );
  NOR U15678 ( .A(n15896), .B(n15897), .Z(n15397) );
  NOR U15679 ( .A(n15398), .B(n15397), .Z(n15403) );
  NOR U15680 ( .A(n163), .B(n54), .Z(n15402) );
  IV U15681 ( .A(n15402), .Z(n15399) );
  NOR U15682 ( .A(n15403), .B(n15399), .Z(n15406) );
  XOR U15683 ( .A(n15401), .B(n15400), .Z(n15902) );
  IV U15684 ( .A(n15902), .Z(n15404) );
  XOR U15685 ( .A(n15403), .B(n15402), .Z(n15901) );
  NOR U15686 ( .A(n15404), .B(n15901), .Z(n15405) );
  NOR U15687 ( .A(n15406), .B(n15405), .Z(n15410) );
  XOR U15688 ( .A(n15408), .B(n15407), .Z(n15409) );
  NOR U15689 ( .A(n15410), .B(n15409), .Z(n15414) );
  XOR U15690 ( .A(n15410), .B(n15409), .Z(n15411) );
  IV U15691 ( .A(n15411), .Z(n15912) );
  NOR U15692 ( .A(n165), .B(n54), .Z(n15913) );
  IV U15693 ( .A(n15913), .Z(n15412) );
  NOR U15694 ( .A(n15912), .B(n15412), .Z(n15413) );
  NOR U15695 ( .A(n15414), .B(n15413), .Z(n15417) );
  NOR U15696 ( .A(n167), .B(n54), .Z(n15416) );
  IV U15697 ( .A(n15416), .Z(n15415) );
  NOR U15698 ( .A(n15417), .B(n15415), .Z(n15421) );
  XOR U15699 ( .A(n15417), .B(n15416), .Z(n15916) );
  XOR U15700 ( .A(n15419), .B(n15418), .Z(n15917) );
  NOR U15701 ( .A(n15916), .B(n15917), .Z(n15420) );
  NOR U15702 ( .A(n15421), .B(n15420), .Z(n28590) );
  XOR U15703 ( .A(n15423), .B(n15422), .Z(n15424) );
  IV U15704 ( .A(n15424), .Z(n28589) );
  NOR U15705 ( .A(n28590), .B(n28589), .Z(n31626) );
  XOR U15706 ( .A(n15426), .B(n15425), .Z(n28597) );
  NOR U15707 ( .A(n31626), .B(n28597), .Z(n28594) );
  NOR U15708 ( .A(n161), .B(n55), .Z(n16396) );
  XOR U15709 ( .A(n15428), .B(n15427), .Z(n15818) );
  NOR U15710 ( .A(n143), .B(n55), .Z(n15819) );
  IV U15711 ( .A(n15819), .Z(n15429) );
  NOR U15712 ( .A(n15818), .B(n15429), .Z(n15821) );
  XOR U15713 ( .A(n15431), .B(n15430), .Z(n15798) );
  NOR U15714 ( .A(n137), .B(n55), .Z(n15799) );
  IV U15715 ( .A(n15799), .Z(n15432) );
  NOR U15716 ( .A(n15798), .B(n15432), .Z(n15801) );
  NOR U15717 ( .A(n131), .B(n55), .Z(n15435) );
  XOR U15718 ( .A(n15434), .B(n15433), .Z(n16282) );
  IV U15719 ( .A(n15435), .Z(n16283) );
  NOR U15720 ( .A(n126), .B(n55), .Z(n15769) );
  XOR U15721 ( .A(n15437), .B(n15436), .Z(n15760) );
  NOR U15722 ( .A(n79), .B(n55), .Z(n15440) );
  XOR U15723 ( .A(n15439), .B(n15438), .Z(n15441) );
  NOR U15724 ( .A(n15440), .B(n15441), .Z(n15731) );
  IV U15725 ( .A(n15440), .Z(n16232) );
  IV U15726 ( .A(n15441), .Z(n16231) );
  NOR U15727 ( .A(n16232), .B(n16231), .Z(n15729) );
  XOR U15728 ( .A(n15443), .B(n15442), .Z(n15445) );
  IV U15729 ( .A(n15445), .Z(n16218) );
  NOR U15730 ( .A(n80), .B(n55), .Z(n15444) );
  IV U15731 ( .A(n15444), .Z(n16217) );
  NOR U15732 ( .A(n16218), .B(n16217), .Z(n15718) );
  NOR U15733 ( .A(n15445), .B(n15444), .Z(n15716) );
  XOR U15734 ( .A(n15447), .B(n15446), .Z(n15711) );
  NOR U15735 ( .A(n116), .B(n55), .Z(n15712) );
  IV U15736 ( .A(n15712), .Z(n15448) );
  NOR U15737 ( .A(n15711), .B(n15448), .Z(n15715) );
  NOR U15738 ( .A(n81), .B(n55), .Z(n15706) );
  XOR U15739 ( .A(n15450), .B(n15449), .Z(n15707) );
  NOR U15740 ( .A(n15706), .B(n15707), .Z(n15710) );
  NOR U15741 ( .A(n82), .B(n55), .Z(n15454) );
  IV U15742 ( .A(n15454), .Z(n16195) );
  XOR U15743 ( .A(n15452), .B(n15451), .Z(n15453) );
  IV U15744 ( .A(n15453), .Z(n16194) );
  NOR U15745 ( .A(n16195), .B(n16194), .Z(n15697) );
  NOR U15746 ( .A(n15454), .B(n15453), .Z(n15695) );
  XOR U15747 ( .A(n15456), .B(n15455), .Z(n15457) );
  NOR U15748 ( .A(n83), .B(n55), .Z(n15458) );
  NOR U15749 ( .A(n15457), .B(n15458), .Z(n15684) );
  IV U15750 ( .A(n15457), .Z(n16183) );
  IV U15751 ( .A(n15458), .Z(n16182) );
  NOR U15752 ( .A(n16183), .B(n16182), .Z(n15682) );
  XOR U15753 ( .A(n15460), .B(n15459), .Z(n15461) );
  NOR U15754 ( .A(n84), .B(n55), .Z(n15462) );
  NOR U15755 ( .A(n15461), .B(n15462), .Z(n15672) );
  IV U15756 ( .A(n15461), .Z(n16169) );
  IV U15757 ( .A(n15462), .Z(n16168) );
  NOR U15758 ( .A(n16169), .B(n16168), .Z(n15670) );
  XOR U15759 ( .A(n15464), .B(n15463), .Z(n15657) );
  IV U15760 ( .A(n15657), .Z(n15955) );
  NOR U15761 ( .A(n85), .B(n55), .Z(n15656) );
  IV U15762 ( .A(n15656), .Z(n15954) );
  NOR U15763 ( .A(n15955), .B(n15954), .Z(n15660) );
  XOR U15764 ( .A(n15466), .B(n15465), .Z(n15467) );
  XOR U15765 ( .A(n15468), .B(n15467), .Z(n15471) );
  NOR U15766 ( .A(n111), .B(n55), .Z(n15470) );
  IV U15767 ( .A(n15470), .Z(n15469) );
  NOR U15768 ( .A(n15471), .B(n15469), .Z(n15655) );
  XOR U15769 ( .A(n15471), .B(n15470), .Z(n15959) );
  NOR U15770 ( .A(n86), .B(n55), .Z(n15649) );
  XOR U15771 ( .A(n15473), .B(n15472), .Z(n15648) );
  NOR U15772 ( .A(n15649), .B(n15648), .Z(n15652) );
  XOR U15773 ( .A(n15475), .B(n15474), .Z(n15644) );
  NOR U15774 ( .A(n110), .B(n55), .Z(n15643) );
  IV U15775 ( .A(n15643), .Z(n15476) );
  NOR U15776 ( .A(n15644), .B(n15476), .Z(n15646) );
  XOR U15777 ( .A(n15478), .B(n15477), .Z(n15639) );
  NOR U15778 ( .A(n109), .B(n55), .Z(n15640) );
  IV U15779 ( .A(n15640), .Z(n15479) );
  NOR U15780 ( .A(n15639), .B(n15479), .Z(n15642) );
  XOR U15781 ( .A(n15481), .B(n15480), .Z(n15636) );
  NOR U15782 ( .A(n108), .B(n55), .Z(n15635) );
  IV U15783 ( .A(n15635), .Z(n15482) );
  NOR U15784 ( .A(n15636), .B(n15482), .Z(n15638) );
  NOR U15785 ( .A(n87), .B(n55), .Z(n15630) );
  XOR U15786 ( .A(n15484), .B(n15483), .Z(n15629) );
  NOR U15787 ( .A(n15630), .B(n15629), .Z(n15633) );
  XOR U15788 ( .A(n15486), .B(n15485), .Z(n15625) );
  NOR U15789 ( .A(n107), .B(n55), .Z(n15624) );
  IV U15790 ( .A(n15624), .Z(n15487) );
  NOR U15791 ( .A(n15625), .B(n15487), .Z(n15627) );
  XOR U15792 ( .A(n15489), .B(n15488), .Z(n15620) );
  NOR U15793 ( .A(n88), .B(n55), .Z(n15621) );
  IV U15794 ( .A(n15621), .Z(n15490) );
  NOR U15795 ( .A(n15620), .B(n15490), .Z(n15623) );
  XOR U15796 ( .A(n15492), .B(n15491), .Z(n15617) );
  NOR U15797 ( .A(n106), .B(n55), .Z(n15616) );
  IV U15798 ( .A(n15616), .Z(n15493) );
  NOR U15799 ( .A(n15617), .B(n15493), .Z(n15619) );
  IV U15800 ( .A(n15494), .Z(n15496) );
  XOR U15801 ( .A(n15496), .B(n15495), .Z(n15612) );
  NOR U15802 ( .A(n105), .B(n55), .Z(n15613) );
  IV U15803 ( .A(n15613), .Z(n15497) );
  NOR U15804 ( .A(n15612), .B(n15497), .Z(n15615) );
  IV U15805 ( .A(n15498), .Z(n15500) );
  XOR U15806 ( .A(n15500), .B(n15499), .Z(n15608) );
  NOR U15807 ( .A(n104), .B(n55), .Z(n15609) );
  IV U15808 ( .A(n15609), .Z(n15501) );
  NOR U15809 ( .A(n15608), .B(n15501), .Z(n15611) );
  IV U15810 ( .A(n15502), .Z(n15504) );
  XOR U15811 ( .A(n15504), .B(n15503), .Z(n15604) );
  NOR U15812 ( .A(n89), .B(n55), .Z(n15605) );
  IV U15813 ( .A(n15605), .Z(n15505) );
  NOR U15814 ( .A(n15604), .B(n15505), .Z(n15607) );
  IV U15815 ( .A(n15506), .Z(n15508) );
  XOR U15816 ( .A(n15508), .B(n15507), .Z(n15592) );
  NOR U15817 ( .A(n90), .B(n55), .Z(n15593) );
  IV U15818 ( .A(n15593), .Z(n15509) );
  NOR U15819 ( .A(n15592), .B(n15509), .Z(n15595) );
  IV U15820 ( .A(n15510), .Z(n15512) );
  XOR U15821 ( .A(n15512), .B(n15511), .Z(n15588) );
  NOR U15822 ( .A(n102), .B(n55), .Z(n15589) );
  IV U15823 ( .A(n15589), .Z(n15513) );
  NOR U15824 ( .A(n15588), .B(n15513), .Z(n15591) );
  IV U15825 ( .A(n15514), .Z(n15516) );
  XOR U15826 ( .A(n15516), .B(n15515), .Z(n15584) );
  NOR U15827 ( .A(n101), .B(n55), .Z(n15585) );
  IV U15828 ( .A(n15585), .Z(n15517) );
  NOR U15829 ( .A(n15584), .B(n15517), .Z(n15587) );
  IV U15830 ( .A(n15518), .Z(n15520) );
  XOR U15831 ( .A(n15520), .B(n15519), .Z(n15580) );
  NOR U15832 ( .A(n100), .B(n55), .Z(n15581) );
  IV U15833 ( .A(n15581), .Z(n15521) );
  NOR U15834 ( .A(n15580), .B(n15521), .Z(n15583) );
  IV U15835 ( .A(n15522), .Z(n15524) );
  XOR U15836 ( .A(n15524), .B(n15523), .Z(n15576) );
  NOR U15837 ( .A(n99), .B(n55), .Z(n15577) );
  IV U15838 ( .A(n15577), .Z(n15525) );
  NOR U15839 ( .A(n15576), .B(n15525), .Z(n15579) );
  IV U15840 ( .A(n15526), .Z(n15528) );
  XOR U15841 ( .A(n15528), .B(n15527), .Z(n15572) );
  NOR U15842 ( .A(n98), .B(n55), .Z(n15573) );
  IV U15843 ( .A(n15573), .Z(n15529) );
  NOR U15844 ( .A(n15572), .B(n15529), .Z(n15575) );
  XOR U15845 ( .A(n15531), .B(n15530), .Z(n15568) );
  NOR U15846 ( .A(n91), .B(n55), .Z(n15569) );
  IV U15847 ( .A(n15569), .Z(n15532) );
  NOR U15848 ( .A(n15568), .B(n15532), .Z(n15571) );
  IV U15849 ( .A(n15533), .Z(n15535) );
  XOR U15850 ( .A(n15535), .B(n15534), .Z(n15556) );
  NOR U15851 ( .A(n96), .B(n55), .Z(n15557) );
  IV U15852 ( .A(n15557), .Z(n15536) );
  NOR U15853 ( .A(n15556), .B(n15536), .Z(n15559) );
  NOR U15854 ( .A(n95), .B(n55), .Z(n15553) );
  IV U15855 ( .A(n15553), .Z(n15539) );
  XOR U15856 ( .A(n15538), .B(n15537), .Z(n15552) );
  NOR U15857 ( .A(n15539), .B(n15552), .Z(n15555) );
  NOR U15858 ( .A(n93), .B(n55), .Z(n16530) );
  IV U15859 ( .A(n16530), .Z(n15540) );
  NOR U15860 ( .A(n54), .B(n168), .Z(n15548) );
  IV U15861 ( .A(n15548), .Z(n15543) );
  NOR U15862 ( .A(n15540), .B(n15543), .Z(n15541) );
  IV U15863 ( .A(n15541), .Z(n15542) );
  NOR U15864 ( .A(n94), .B(n15542), .Z(n15551) );
  NOR U15865 ( .A(n15543), .B(n93), .Z(n15544) );
  XOR U15866 ( .A(n94), .B(n15544), .Z(n15545) );
  NOR U15867 ( .A(n55), .B(n15545), .Z(n15546) );
  IV U15868 ( .A(n15546), .Z(n16041) );
  XOR U15869 ( .A(n15548), .B(n15547), .Z(n16040) );
  IV U15870 ( .A(n16040), .Z(n15549) );
  NOR U15871 ( .A(n16041), .B(n15549), .Z(n15550) );
  NOR U15872 ( .A(n15551), .B(n15550), .Z(n16037) );
  XOR U15873 ( .A(n15553), .B(n15552), .Z(n16036) );
  NOR U15874 ( .A(n16037), .B(n16036), .Z(n15554) );
  NOR U15875 ( .A(n15555), .B(n15554), .Z(n16032) );
  XOR U15876 ( .A(n15557), .B(n15556), .Z(n16033) );
  NOR U15877 ( .A(n16032), .B(n16033), .Z(n15558) );
  NOR U15878 ( .A(n15559), .B(n15558), .Z(n15564) );
  XOR U15879 ( .A(n15561), .B(n15560), .Z(n15563) );
  IV U15880 ( .A(n15563), .Z(n15562) );
  NOR U15881 ( .A(n15564), .B(n15562), .Z(n15567) );
  XOR U15882 ( .A(n15564), .B(n15563), .Z(n16029) );
  NOR U15883 ( .A(n97), .B(n55), .Z(n16030) );
  IV U15884 ( .A(n16030), .Z(n15565) );
  NOR U15885 ( .A(n16029), .B(n15565), .Z(n15566) );
  NOR U15886 ( .A(n15567), .B(n15566), .Z(n16025) );
  XOR U15887 ( .A(n15569), .B(n15568), .Z(n16026) );
  NOR U15888 ( .A(n16025), .B(n16026), .Z(n15570) );
  NOR U15889 ( .A(n15571), .B(n15570), .Z(n16021) );
  XOR U15890 ( .A(n15573), .B(n15572), .Z(n16022) );
  NOR U15891 ( .A(n16021), .B(n16022), .Z(n15574) );
  NOR U15892 ( .A(n15575), .B(n15574), .Z(n16017) );
  XOR U15893 ( .A(n15577), .B(n15576), .Z(n16018) );
  NOR U15894 ( .A(n16017), .B(n16018), .Z(n15578) );
  NOR U15895 ( .A(n15579), .B(n15578), .Z(n16013) );
  XOR U15896 ( .A(n15581), .B(n15580), .Z(n16014) );
  NOR U15897 ( .A(n16013), .B(n16014), .Z(n15582) );
  NOR U15898 ( .A(n15583), .B(n15582), .Z(n16009) );
  XOR U15899 ( .A(n15585), .B(n15584), .Z(n16010) );
  NOR U15900 ( .A(n16009), .B(n16010), .Z(n15586) );
  NOR U15901 ( .A(n15587), .B(n15586), .Z(n16005) );
  XOR U15902 ( .A(n15589), .B(n15588), .Z(n16006) );
  NOR U15903 ( .A(n16005), .B(n16006), .Z(n15590) );
  NOR U15904 ( .A(n15591), .B(n15590), .Z(n16001) );
  XOR U15905 ( .A(n15593), .B(n15592), .Z(n16002) );
  NOR U15906 ( .A(n16001), .B(n16002), .Z(n15594) );
  NOR U15907 ( .A(n15595), .B(n15594), .Z(n15600) );
  XOR U15908 ( .A(n15597), .B(n15596), .Z(n15599) );
  IV U15909 ( .A(n15599), .Z(n15598) );
  NOR U15910 ( .A(n15600), .B(n15598), .Z(n15603) );
  XOR U15911 ( .A(n15600), .B(n15599), .Z(n15998) );
  NOR U15912 ( .A(n103), .B(n55), .Z(n15999) );
  IV U15913 ( .A(n15999), .Z(n15601) );
  NOR U15914 ( .A(n15998), .B(n15601), .Z(n15602) );
  NOR U15915 ( .A(n15603), .B(n15602), .Z(n15994) );
  XOR U15916 ( .A(n15605), .B(n15604), .Z(n15995) );
  NOR U15917 ( .A(n15994), .B(n15995), .Z(n15606) );
  NOR U15918 ( .A(n15607), .B(n15606), .Z(n15991) );
  XOR U15919 ( .A(n15609), .B(n15608), .Z(n15990) );
  NOR U15920 ( .A(n15991), .B(n15990), .Z(n15610) );
  NOR U15921 ( .A(n15611), .B(n15610), .Z(n15986) );
  XOR U15922 ( .A(n15613), .B(n15612), .Z(n15987) );
  NOR U15923 ( .A(n15986), .B(n15987), .Z(n15614) );
  NOR U15924 ( .A(n15615), .B(n15614), .Z(n15983) );
  XOR U15925 ( .A(n15617), .B(n15616), .Z(n15982) );
  NOR U15926 ( .A(n15983), .B(n15982), .Z(n15618) );
  NOR U15927 ( .A(n15619), .B(n15618), .Z(n15978) );
  XOR U15928 ( .A(n15621), .B(n15620), .Z(n15979) );
  NOR U15929 ( .A(n15978), .B(n15979), .Z(n15622) );
  NOR U15930 ( .A(n15623), .B(n15622), .Z(n15977) );
  XOR U15931 ( .A(n15625), .B(n15624), .Z(n15976) );
  NOR U15932 ( .A(n15977), .B(n15976), .Z(n15626) );
  NOR U15933 ( .A(n15627), .B(n15626), .Z(n15628) );
  IV U15934 ( .A(n15628), .Z(n15974) );
  XOR U15935 ( .A(n15630), .B(n15629), .Z(n15631) );
  IV U15936 ( .A(n15631), .Z(n15973) );
  NOR U15937 ( .A(n15974), .B(n15973), .Z(n15632) );
  NOR U15938 ( .A(n15633), .B(n15632), .Z(n15634) );
  IV U15939 ( .A(n15634), .Z(n15969) );
  XOR U15940 ( .A(n15636), .B(n15635), .Z(n15968) );
  NOR U15941 ( .A(n15969), .B(n15968), .Z(n15637) );
  NOR U15942 ( .A(n15638), .B(n15637), .Z(n15965) );
  XOR U15943 ( .A(n15640), .B(n15639), .Z(n15964) );
  NOR U15944 ( .A(n15965), .B(n15964), .Z(n15641) );
  NOR U15945 ( .A(n15642), .B(n15641), .Z(n15963) );
  XOR U15946 ( .A(n15644), .B(n15643), .Z(n15962) );
  NOR U15947 ( .A(n15963), .B(n15962), .Z(n15645) );
  NOR U15948 ( .A(n15646), .B(n15645), .Z(n15647) );
  IV U15949 ( .A(n15647), .Z(n16149) );
  XOR U15950 ( .A(n15649), .B(n15648), .Z(n15650) );
  IV U15951 ( .A(n15650), .Z(n16148) );
  NOR U15952 ( .A(n16149), .B(n16148), .Z(n15651) );
  NOR U15953 ( .A(n15652), .B(n15651), .Z(n15960) );
  IV U15954 ( .A(n15960), .Z(n15653) );
  NOR U15955 ( .A(n15959), .B(n15653), .Z(n15654) );
  NOR U15956 ( .A(n15655), .B(n15654), .Z(n15957) );
  NOR U15957 ( .A(n15657), .B(n15656), .Z(n15658) );
  NOR U15958 ( .A(n15957), .B(n15658), .Z(n15659) );
  NOR U15959 ( .A(n15660), .B(n15659), .Z(n15666) );
  NOR U15960 ( .A(n112), .B(n55), .Z(n15665) );
  IV U15961 ( .A(n15665), .Z(n15661) );
  NOR U15962 ( .A(n15666), .B(n15661), .Z(n15668) );
  XOR U15963 ( .A(n15663), .B(n15662), .Z(n15664) );
  IV U15964 ( .A(n15664), .Z(n15951) );
  XOR U15965 ( .A(n15666), .B(n15665), .Z(n15950) );
  NOR U15966 ( .A(n15951), .B(n15950), .Z(n15667) );
  NOR U15967 ( .A(n15668), .B(n15667), .Z(n16171) );
  IV U15968 ( .A(n16171), .Z(n15669) );
  NOR U15969 ( .A(n15670), .B(n15669), .Z(n15671) );
  NOR U15970 ( .A(n15672), .B(n15671), .Z(n15678) );
  IV U15971 ( .A(n15678), .Z(n15674) );
  NOR U15972 ( .A(n113), .B(n55), .Z(n15673) );
  IV U15973 ( .A(n15673), .Z(n15677) );
  NOR U15974 ( .A(n15674), .B(n15677), .Z(n15680) );
  XOR U15975 ( .A(n15676), .B(n15675), .Z(n15949) );
  XOR U15976 ( .A(n15678), .B(n15677), .Z(n15948) );
  NOR U15977 ( .A(n15949), .B(n15948), .Z(n15679) );
  NOR U15978 ( .A(n15680), .B(n15679), .Z(n16185) );
  IV U15979 ( .A(n16185), .Z(n15681) );
  NOR U15980 ( .A(n15682), .B(n15681), .Z(n15683) );
  NOR U15981 ( .A(n15684), .B(n15683), .Z(n15692) );
  IV U15982 ( .A(n15692), .Z(n15686) );
  NOR U15983 ( .A(n114), .B(n55), .Z(n15685) );
  IV U15984 ( .A(n15685), .Z(n15691) );
  NOR U15985 ( .A(n15686), .B(n15691), .Z(n15694) );
  XOR U15986 ( .A(n15688), .B(n15687), .Z(n15689) );
  XOR U15987 ( .A(n15690), .B(n15689), .Z(n15945) );
  XOR U15988 ( .A(n15692), .B(n15691), .Z(n15944) );
  NOR U15989 ( .A(n15945), .B(n15944), .Z(n15693) );
  NOR U15990 ( .A(n15694), .B(n15693), .Z(n16197) );
  NOR U15991 ( .A(n15695), .B(n16197), .Z(n15696) );
  NOR U15992 ( .A(n15697), .B(n15696), .Z(n15702) );
  NOR U15993 ( .A(n115), .B(n55), .Z(n15701) );
  IV U15994 ( .A(n15701), .Z(n15698) );
  NOR U15995 ( .A(n15702), .B(n15698), .Z(n15704) );
  XOR U15996 ( .A(n15700), .B(n15699), .Z(n15940) );
  XOR U15997 ( .A(n15702), .B(n15701), .Z(n15941) );
  NOR U15998 ( .A(n15940), .B(n15941), .Z(n15703) );
  NOR U15999 ( .A(n15704), .B(n15703), .Z(n15705) );
  IV U16000 ( .A(n15705), .Z(n16207) );
  XOR U16001 ( .A(n15707), .B(n15706), .Z(n15708) );
  IV U16002 ( .A(n15708), .Z(n16206) );
  NOR U16003 ( .A(n16207), .B(n16206), .Z(n15709) );
  NOR U16004 ( .A(n15710), .B(n15709), .Z(n15937) );
  IV U16005 ( .A(n15937), .Z(n15713) );
  XOR U16006 ( .A(n15712), .B(n15711), .Z(n15936) );
  NOR U16007 ( .A(n15713), .B(n15936), .Z(n15714) );
  NOR U16008 ( .A(n15715), .B(n15714), .Z(n16220) );
  NOR U16009 ( .A(n15716), .B(n16220), .Z(n15717) );
  NOR U16010 ( .A(n15718), .B(n15717), .Z(n15725) );
  NOR U16011 ( .A(n117), .B(n55), .Z(n15724) );
  IV U16012 ( .A(n15724), .Z(n15719) );
  NOR U16013 ( .A(n15725), .B(n15719), .Z(n15727) );
  XOR U16014 ( .A(n15721), .B(n15720), .Z(n15722) );
  XOR U16015 ( .A(n15723), .B(n15722), .Z(n15934) );
  XOR U16016 ( .A(n15725), .B(n15724), .Z(n15933) );
  NOR U16017 ( .A(n15934), .B(n15933), .Z(n15726) );
  NOR U16018 ( .A(n15727), .B(n15726), .Z(n16234) );
  IV U16019 ( .A(n16234), .Z(n15728) );
  NOR U16020 ( .A(n15729), .B(n15728), .Z(n15730) );
  NOR U16021 ( .A(n15731), .B(n15730), .Z(n15732) );
  IV U16022 ( .A(n15732), .Z(n15739) );
  NOR U16023 ( .A(n119), .B(n55), .Z(n15738) );
  IV U16024 ( .A(n15738), .Z(n15733) );
  NOR U16025 ( .A(n15739), .B(n15733), .Z(n15741) );
  XOR U16026 ( .A(n15735), .B(n15734), .Z(n15736) );
  XOR U16027 ( .A(n15737), .B(n15736), .Z(n15930) );
  XOR U16028 ( .A(n15739), .B(n15738), .Z(n15929) );
  NOR U16029 ( .A(n15930), .B(n15929), .Z(n15740) );
  NOR U16030 ( .A(n15741), .B(n15740), .Z(n15742) );
  NOR U16031 ( .A(n120), .B(n55), .Z(n15743) );
  IV U16032 ( .A(n15743), .Z(n16243) );
  NOR U16033 ( .A(n15742), .B(n16243), .Z(n15750) );
  IV U16034 ( .A(n15742), .Z(n16244) );
  NOR U16035 ( .A(n15743), .B(n16244), .Z(n15748) );
  XOR U16036 ( .A(n15745), .B(n15744), .Z(n15746) );
  XOR U16037 ( .A(n15747), .B(n15746), .Z(n16246) );
  NOR U16038 ( .A(n15748), .B(n16246), .Z(n15749) );
  NOR U16039 ( .A(n15750), .B(n15749), .Z(n15757) );
  NOR U16040 ( .A(n123), .B(n55), .Z(n15756) );
  IV U16041 ( .A(n15756), .Z(n15751) );
  NOR U16042 ( .A(n15757), .B(n15751), .Z(n15759) );
  XOR U16043 ( .A(n15753), .B(n15752), .Z(n15754) );
  XOR U16044 ( .A(n15755), .B(n15754), .Z(n15926) );
  XOR U16045 ( .A(n15757), .B(n15756), .Z(n15925) );
  NOR U16046 ( .A(n15926), .B(n15925), .Z(n15758) );
  NOR U16047 ( .A(n15759), .B(n15758), .Z(n15761) );
  IV U16048 ( .A(n15761), .Z(n16259) );
  NOR U16049 ( .A(n15760), .B(n16259), .Z(n15764) );
  IV U16050 ( .A(n15760), .Z(n16260) );
  NOR U16051 ( .A(n15761), .B(n16260), .Z(n15762) );
  NOR U16052 ( .A(n125), .B(n55), .Z(n16262) );
  NOR U16053 ( .A(n15762), .B(n16262), .Z(n15763) );
  NOR U16054 ( .A(n15764), .B(n15763), .Z(n15770) );
  NOR U16055 ( .A(n15769), .B(n15770), .Z(n15774) );
  XOR U16056 ( .A(n15766), .B(n15765), .Z(n15767) );
  XOR U16057 ( .A(n15768), .B(n15767), .Z(n16270) );
  IV U16058 ( .A(n16270), .Z(n15772) );
  IV U16059 ( .A(n15769), .Z(n16268) );
  IV U16060 ( .A(n15770), .Z(n16267) );
  NOR U16061 ( .A(n16268), .B(n16267), .Z(n15771) );
  NOR U16062 ( .A(n15772), .B(n15771), .Z(n15773) );
  NOR U16063 ( .A(n15774), .B(n15773), .Z(n15775) );
  IV U16064 ( .A(n15775), .Z(n15778) );
  NOR U16065 ( .A(n128), .B(n55), .Z(n15777) );
  IV U16066 ( .A(n15777), .Z(n15776) );
  NOR U16067 ( .A(n15778), .B(n15776), .Z(n15782) );
  XOR U16068 ( .A(n15778), .B(n15777), .Z(n15922) );
  XOR U16069 ( .A(n15780), .B(n15779), .Z(n15921) );
  NOR U16070 ( .A(n15922), .B(n15921), .Z(n15781) );
  NOR U16071 ( .A(n15782), .B(n15781), .Z(n16285) );
  NOR U16072 ( .A(n133), .B(n55), .Z(n15784) );
  IV U16073 ( .A(n15784), .Z(n15783) );
  NOR U16074 ( .A(n15785), .B(n15783), .Z(n15789) );
  XOR U16075 ( .A(n15785), .B(n15784), .Z(n15920) );
  XOR U16076 ( .A(n15787), .B(n15786), .Z(n15919) );
  NOR U16077 ( .A(n15920), .B(n15919), .Z(n15788) );
  NOR U16078 ( .A(n15789), .B(n15788), .Z(n15794) );
  XOR U16079 ( .A(n15791), .B(n15790), .Z(n15793) );
  IV U16080 ( .A(n15793), .Z(n15792) );
  NOR U16081 ( .A(n15794), .B(n15792), .Z(n15797) );
  XOR U16082 ( .A(n15794), .B(n15793), .Z(n16299) );
  NOR U16083 ( .A(n135), .B(n55), .Z(n16300) );
  IV U16084 ( .A(n16300), .Z(n15795) );
  NOR U16085 ( .A(n16299), .B(n15795), .Z(n15796) );
  NOR U16086 ( .A(n15797), .B(n15796), .Z(n16305) );
  XOR U16087 ( .A(n15799), .B(n15798), .Z(n16304) );
  NOR U16088 ( .A(n16305), .B(n16304), .Z(n15800) );
  NOR U16089 ( .A(n15801), .B(n15800), .Z(n15804) );
  NOR U16090 ( .A(n139), .B(n55), .Z(n15803) );
  IV U16091 ( .A(n15803), .Z(n15802) );
  NOR U16092 ( .A(n15804), .B(n15802), .Z(n15809) );
  XOR U16093 ( .A(n15804), .B(n15803), .Z(n16311) );
  XOR U16094 ( .A(n15806), .B(n15805), .Z(n16312) );
  IV U16095 ( .A(n16312), .Z(n15807) );
  NOR U16096 ( .A(n16311), .B(n15807), .Z(n15808) );
  NOR U16097 ( .A(n15809), .B(n15808), .Z(n15813) );
  XOR U16098 ( .A(n15811), .B(n15810), .Z(n15812) );
  NOR U16099 ( .A(n15813), .B(n15812), .Z(n15817) );
  XOR U16100 ( .A(n15813), .B(n15812), .Z(n16322) );
  IV U16101 ( .A(n16322), .Z(n15815) );
  NOR U16102 ( .A(n141), .B(n55), .Z(n15814) );
  IV U16103 ( .A(n15814), .Z(n16323) );
  NOR U16104 ( .A(n15815), .B(n16323), .Z(n15816) );
  NOR U16105 ( .A(n15817), .B(n15816), .Z(n16328) );
  XOR U16106 ( .A(n15819), .B(n15818), .Z(n16327) );
  NOR U16107 ( .A(n16328), .B(n16327), .Z(n15820) );
  NOR U16108 ( .A(n15821), .B(n15820), .Z(n15826) );
  NOR U16109 ( .A(n145), .B(n55), .Z(n15825) );
  IV U16110 ( .A(n15825), .Z(n15822) );
  NOR U16111 ( .A(n15826), .B(n15822), .Z(n15829) );
  XOR U16112 ( .A(n15824), .B(n15823), .Z(n16335) );
  IV U16113 ( .A(n16335), .Z(n15827) );
  XOR U16114 ( .A(n15826), .B(n15825), .Z(n16334) );
  NOR U16115 ( .A(n15827), .B(n16334), .Z(n15828) );
  NOR U16116 ( .A(n15829), .B(n15828), .Z(n15833) );
  XOR U16117 ( .A(n15831), .B(n15830), .Z(n15832) );
  NOR U16118 ( .A(n15833), .B(n15832), .Z(n15837) );
  XOR U16119 ( .A(n15833), .B(n15832), .Z(n15834) );
  IV U16120 ( .A(n15834), .Z(n16345) );
  NOR U16121 ( .A(n147), .B(n55), .Z(n16346) );
  IV U16122 ( .A(n16346), .Z(n15835) );
  NOR U16123 ( .A(n16345), .B(n15835), .Z(n15836) );
  NOR U16124 ( .A(n15837), .B(n15836), .Z(n15840) );
  NOR U16125 ( .A(n148), .B(n55), .Z(n15839) );
  IV U16126 ( .A(n15839), .Z(n15838) );
  NOR U16127 ( .A(n15840), .B(n15838), .Z(n15844) );
  XOR U16128 ( .A(n15840), .B(n15839), .Z(n16352) );
  XOR U16129 ( .A(n15842), .B(n15841), .Z(n16353) );
  NOR U16130 ( .A(n16352), .B(n16353), .Z(n15843) );
  NOR U16131 ( .A(n15844), .B(n15843), .Z(n15849) );
  NOR U16132 ( .A(n150), .B(n55), .Z(n15848) );
  IV U16133 ( .A(n15848), .Z(n15845) );
  NOR U16134 ( .A(n15849), .B(n15845), .Z(n15852) );
  XOR U16135 ( .A(n15847), .B(n15846), .Z(n16358) );
  IV U16136 ( .A(n16358), .Z(n15850) );
  XOR U16137 ( .A(n15849), .B(n15848), .Z(n16357) );
  NOR U16138 ( .A(n15850), .B(n16357), .Z(n15851) );
  NOR U16139 ( .A(n15852), .B(n15851), .Z(n15856) );
  XOR U16140 ( .A(n15854), .B(n15853), .Z(n15855) );
  NOR U16141 ( .A(n15856), .B(n15855), .Z(n15860) );
  XOR U16142 ( .A(n15856), .B(n15855), .Z(n16368) );
  IV U16143 ( .A(n16368), .Z(n15858) );
  NOR U16144 ( .A(n153), .B(n55), .Z(n15857) );
  IV U16145 ( .A(n15857), .Z(n16369) );
  NOR U16146 ( .A(n15858), .B(n16369), .Z(n15859) );
  NOR U16147 ( .A(n15860), .B(n15859), .Z(n15863) );
  XOR U16148 ( .A(n15862), .B(n15861), .Z(n15864) );
  NOR U16149 ( .A(n15863), .B(n15864), .Z(n15868) );
  IV U16150 ( .A(n15863), .Z(n15865) );
  XOR U16151 ( .A(n15865), .B(n15864), .Z(n16373) );
  NOR U16152 ( .A(n155), .B(n55), .Z(n16374) );
  IV U16153 ( .A(n16374), .Z(n15866) );
  NOR U16154 ( .A(n16373), .B(n15866), .Z(n15867) );
  NOR U16155 ( .A(n15868), .B(n15867), .Z(n15873) );
  NOR U16156 ( .A(n156), .B(n55), .Z(n15872) );
  IV U16157 ( .A(n15872), .Z(n15869) );
  NOR U16158 ( .A(n15873), .B(n15869), .Z(n15876) );
  XOR U16159 ( .A(n15871), .B(n15870), .Z(n16380) );
  IV U16160 ( .A(n16380), .Z(n15874) );
  XOR U16161 ( .A(n15873), .B(n15872), .Z(n16379) );
  NOR U16162 ( .A(n15874), .B(n16379), .Z(n15875) );
  NOR U16163 ( .A(n15876), .B(n15875), .Z(n15880) );
  XOR U16164 ( .A(n15878), .B(n15877), .Z(n15879) );
  NOR U16165 ( .A(n15880), .B(n15879), .Z(n15884) );
  XOR U16166 ( .A(n15880), .B(n15879), .Z(n16390) );
  IV U16167 ( .A(n16390), .Z(n15882) );
  NOR U16168 ( .A(n158), .B(n55), .Z(n16389) );
  IV U16169 ( .A(n16389), .Z(n15881) );
  NOR U16170 ( .A(n15882), .B(n15881), .Z(n15883) );
  NOR U16171 ( .A(n15884), .B(n15883), .Z(n16399) );
  IV U16172 ( .A(n16399), .Z(n15885) );
  NOR U16173 ( .A(n16396), .B(n15885), .Z(n15891) );
  XOR U16174 ( .A(n15887), .B(n15886), .Z(n16397) );
  IV U16175 ( .A(n16396), .Z(n15888) );
  NOR U16176 ( .A(n16399), .B(n15888), .Z(n15889) );
  NOR U16177 ( .A(n16397), .B(n15889), .Z(n15890) );
  NOR U16178 ( .A(n15891), .B(n15890), .Z(n15895) );
  IV U16179 ( .A(n15895), .Z(n15893) );
  NOR U16180 ( .A(n163), .B(n55), .Z(n15892) );
  IV U16181 ( .A(n15892), .Z(n15894) );
  NOR U16182 ( .A(n15893), .B(n15894), .Z(n15900) );
  XOR U16183 ( .A(n15895), .B(n15894), .Z(n16405) );
  XOR U16184 ( .A(n15897), .B(n15896), .Z(n16404) );
  IV U16185 ( .A(n16404), .Z(n15898) );
  NOR U16186 ( .A(n16405), .B(n15898), .Z(n15899) );
  NOR U16187 ( .A(n15900), .B(n15899), .Z(n15904) );
  XOR U16188 ( .A(n15902), .B(n15901), .Z(n15903) );
  NOR U16189 ( .A(n15904), .B(n15903), .Z(n15908) );
  XOR U16190 ( .A(n15904), .B(n15903), .Z(n15905) );
  IV U16191 ( .A(n15905), .Z(n16908) );
  NOR U16192 ( .A(n165), .B(n55), .Z(n16909) );
  IV U16193 ( .A(n16909), .Z(n15906) );
  NOR U16194 ( .A(n16908), .B(n15906), .Z(n15907) );
  NOR U16195 ( .A(n15908), .B(n15907), .Z(n15911) );
  NOR U16196 ( .A(n167), .B(n55), .Z(n15910) );
  IV U16197 ( .A(n15910), .Z(n15909) );
  NOR U16198 ( .A(n15911), .B(n15909), .Z(n15915) );
  XOR U16199 ( .A(n15911), .B(n15910), .Z(n16925) );
  XOR U16200 ( .A(n15913), .B(n15912), .Z(n16926) );
  NOR U16201 ( .A(n16925), .B(n16926), .Z(n15914) );
  NOR U16202 ( .A(n15915), .B(n15914), .Z(n28588) );
  XOR U16203 ( .A(n15917), .B(n15916), .Z(n15918) );
  IV U16204 ( .A(n15918), .Z(n28587) );
  XOR U16205 ( .A(n28588), .B(n28587), .Z(n31617) );
  NOR U16206 ( .A(n165), .B(n56), .Z(n16912) );
  NOR U16207 ( .A(n161), .B(n56), .Z(n16387) );
  XOR U16208 ( .A(n15920), .B(n15919), .Z(n16290) );
  XOR U16209 ( .A(n15922), .B(n15921), .Z(n15923) );
  IV U16210 ( .A(n15923), .Z(n16277) );
  NOR U16211 ( .A(n131), .B(n56), .Z(n16278) );
  IV U16212 ( .A(n16278), .Z(n15924) );
  NOR U16213 ( .A(n16277), .B(n15924), .Z(n16280) );
  NOR U16214 ( .A(n125), .B(n56), .Z(n15927) );
  XOR U16215 ( .A(n15926), .B(n15925), .Z(n16757) );
  NOR U16216 ( .A(n15927), .B(n16757), .Z(n16256) );
  IV U16217 ( .A(n15927), .Z(n16755) );
  IV U16218 ( .A(n16757), .Z(n15928) );
  NOR U16219 ( .A(n16755), .B(n15928), .Z(n16254) );
  NOR U16220 ( .A(n120), .B(n56), .Z(n16240) );
  IV U16221 ( .A(n16240), .Z(n15932) );
  XOR U16222 ( .A(n15930), .B(n15929), .Z(n15931) );
  IV U16223 ( .A(n15931), .Z(n16239) );
  NOR U16224 ( .A(n15932), .B(n16239), .Z(n16242) );
  XOR U16225 ( .A(n15934), .B(n15933), .Z(n16226) );
  IV U16226 ( .A(n16226), .Z(n16727) );
  NOR U16227 ( .A(n79), .B(n56), .Z(n16225) );
  IV U16228 ( .A(n16225), .Z(n16726) );
  NOR U16229 ( .A(n16727), .B(n16726), .Z(n16229) );
  NOR U16230 ( .A(n117), .B(n56), .Z(n15935) );
  IV U16231 ( .A(n15935), .Z(n16222) );
  XOR U16232 ( .A(n15937), .B(n15936), .Z(n16713) );
  IV U16233 ( .A(n16713), .Z(n15938) );
  NOR U16234 ( .A(n80), .B(n56), .Z(n15939) );
  NOR U16235 ( .A(n15938), .B(n15939), .Z(n16215) );
  IV U16236 ( .A(n15939), .Z(n16712) );
  NOR U16237 ( .A(n16713), .B(n16712), .Z(n16213) );
  XOR U16238 ( .A(n15941), .B(n15940), .Z(n15943) );
  IV U16239 ( .A(n15943), .Z(n16700) );
  NOR U16240 ( .A(n81), .B(n56), .Z(n15942) );
  IV U16241 ( .A(n15942), .Z(n16699) );
  NOR U16242 ( .A(n16700), .B(n16699), .Z(n16204) );
  NOR U16243 ( .A(n15943), .B(n15942), .Z(n16202) );
  NOR U16244 ( .A(n82), .B(n56), .Z(n15947) );
  IV U16245 ( .A(n15947), .Z(n16686) );
  XOR U16246 ( .A(n15945), .B(n15944), .Z(n15946) );
  IV U16247 ( .A(n15946), .Z(n16685) );
  NOR U16248 ( .A(n16686), .B(n16685), .Z(n16192) );
  NOR U16249 ( .A(n15947), .B(n15946), .Z(n16190) );
  XOR U16250 ( .A(n15949), .B(n15948), .Z(n16177) );
  IV U16251 ( .A(n16177), .Z(n16672) );
  NOR U16252 ( .A(n83), .B(n56), .Z(n16176) );
  IV U16253 ( .A(n16176), .Z(n16671) );
  NOR U16254 ( .A(n16672), .B(n16671), .Z(n16180) );
  XOR U16255 ( .A(n15951), .B(n15950), .Z(n15952) );
  NOR U16256 ( .A(n84), .B(n56), .Z(n15953) );
  NOR U16257 ( .A(n15952), .B(n15953), .Z(n16165) );
  IV U16258 ( .A(n15952), .Z(n16439) );
  IV U16259 ( .A(n15953), .Z(n16438) );
  NOR U16260 ( .A(n16439), .B(n16438), .Z(n16163) );
  XOR U16261 ( .A(n15955), .B(n15954), .Z(n15956) );
  XOR U16262 ( .A(n15957), .B(n15956), .Z(n16159) );
  NOR U16263 ( .A(n112), .B(n56), .Z(n16158) );
  IV U16264 ( .A(n16158), .Z(n15958) );
  NOR U16265 ( .A(n16159), .B(n15958), .Z(n16161) );
  NOR U16266 ( .A(n85), .B(n56), .Z(n16155) );
  IV U16267 ( .A(n16155), .Z(n15961) );
  XOR U16268 ( .A(n15960), .B(n15959), .Z(n16154) );
  NOR U16269 ( .A(n15961), .B(n16154), .Z(n16157) );
  XOR U16270 ( .A(n15963), .B(n15962), .Z(n16143) );
  IV U16271 ( .A(n16143), .Z(n16450) );
  NOR U16272 ( .A(n86), .B(n56), .Z(n16142) );
  IV U16273 ( .A(n16142), .Z(n16449) );
  NOR U16274 ( .A(n16450), .B(n16449), .Z(n16146) );
  XOR U16275 ( .A(n15965), .B(n15964), .Z(n16138) );
  IV U16276 ( .A(n16138), .Z(n15967) );
  NOR U16277 ( .A(n110), .B(n56), .Z(n15966) );
  IV U16278 ( .A(n15966), .Z(n16139) );
  NOR U16279 ( .A(n15967), .B(n16139), .Z(n16141) );
  NOR U16280 ( .A(n109), .B(n56), .Z(n15971) );
  XOR U16281 ( .A(n15969), .B(n15968), .Z(n15970) );
  NOR U16282 ( .A(n15971), .B(n15970), .Z(n16136) );
  XOR U16283 ( .A(n15971), .B(n15970), .Z(n15972) );
  IV U16284 ( .A(n15972), .Z(n16457) );
  XOR U16285 ( .A(n15974), .B(n15973), .Z(n16130) );
  NOR U16286 ( .A(n108), .B(n56), .Z(n16129) );
  IV U16287 ( .A(n16129), .Z(n15975) );
  NOR U16288 ( .A(n16130), .B(n15975), .Z(n16133) );
  NOR U16289 ( .A(n87), .B(n56), .Z(n16125) );
  XOR U16290 ( .A(n15977), .B(n15976), .Z(n16124) );
  NOR U16291 ( .A(n16125), .B(n16124), .Z(n16128) );
  IV U16292 ( .A(n15978), .Z(n15980) );
  XOR U16293 ( .A(n15980), .B(n15979), .Z(n16119) );
  NOR U16294 ( .A(n107), .B(n56), .Z(n16120) );
  IV U16295 ( .A(n16120), .Z(n15981) );
  NOR U16296 ( .A(n16119), .B(n15981), .Z(n16122) );
  XOR U16297 ( .A(n15983), .B(n15982), .Z(n16115) );
  IV U16298 ( .A(n16115), .Z(n15985) );
  NOR U16299 ( .A(n88), .B(n56), .Z(n15984) );
  IV U16300 ( .A(n15984), .Z(n16116) );
  NOR U16301 ( .A(n15985), .B(n16116), .Z(n16118) );
  IV U16302 ( .A(n15986), .Z(n15988) );
  XOR U16303 ( .A(n15988), .B(n15987), .Z(n16111) );
  NOR U16304 ( .A(n106), .B(n56), .Z(n16112) );
  IV U16305 ( .A(n16112), .Z(n15989) );
  NOR U16306 ( .A(n16111), .B(n15989), .Z(n16114) );
  XOR U16307 ( .A(n15991), .B(n15990), .Z(n16107) );
  IV U16308 ( .A(n16107), .Z(n15993) );
  NOR U16309 ( .A(n105), .B(n56), .Z(n15992) );
  IV U16310 ( .A(n15992), .Z(n16108) );
  NOR U16311 ( .A(n15993), .B(n16108), .Z(n16110) );
  IV U16312 ( .A(n15994), .Z(n15996) );
  XOR U16313 ( .A(n15996), .B(n15995), .Z(n16103) );
  NOR U16314 ( .A(n104), .B(n56), .Z(n16104) );
  IV U16315 ( .A(n16104), .Z(n15997) );
  NOR U16316 ( .A(n16103), .B(n15997), .Z(n16106) );
  XOR U16317 ( .A(n15999), .B(n15998), .Z(n16099) );
  NOR U16318 ( .A(n89), .B(n56), .Z(n16100) );
  IV U16319 ( .A(n16100), .Z(n16000) );
  NOR U16320 ( .A(n16099), .B(n16000), .Z(n16102) );
  IV U16321 ( .A(n16001), .Z(n16003) );
  XOR U16322 ( .A(n16003), .B(n16002), .Z(n16095) );
  NOR U16323 ( .A(n103), .B(n56), .Z(n16096) );
  IV U16324 ( .A(n16096), .Z(n16004) );
  NOR U16325 ( .A(n16095), .B(n16004), .Z(n16098) );
  IV U16326 ( .A(n16005), .Z(n16007) );
  XOR U16327 ( .A(n16007), .B(n16006), .Z(n16091) );
  NOR U16328 ( .A(n90), .B(n56), .Z(n16092) );
  IV U16329 ( .A(n16092), .Z(n16008) );
  NOR U16330 ( .A(n16091), .B(n16008), .Z(n16094) );
  IV U16331 ( .A(n16009), .Z(n16011) );
  XOR U16332 ( .A(n16011), .B(n16010), .Z(n16087) );
  NOR U16333 ( .A(n102), .B(n56), .Z(n16088) );
  IV U16334 ( .A(n16088), .Z(n16012) );
  NOR U16335 ( .A(n16087), .B(n16012), .Z(n16090) );
  IV U16336 ( .A(n16013), .Z(n16015) );
  XOR U16337 ( .A(n16015), .B(n16014), .Z(n16083) );
  NOR U16338 ( .A(n101), .B(n56), .Z(n16084) );
  IV U16339 ( .A(n16084), .Z(n16016) );
  NOR U16340 ( .A(n16083), .B(n16016), .Z(n16086) );
  IV U16341 ( .A(n16017), .Z(n16019) );
  XOR U16342 ( .A(n16019), .B(n16018), .Z(n16079) );
  NOR U16343 ( .A(n100), .B(n56), .Z(n16080) );
  IV U16344 ( .A(n16080), .Z(n16020) );
  NOR U16345 ( .A(n16079), .B(n16020), .Z(n16082) );
  IV U16346 ( .A(n16021), .Z(n16023) );
  XOR U16347 ( .A(n16023), .B(n16022), .Z(n16075) );
  NOR U16348 ( .A(n99), .B(n56), .Z(n16076) );
  IV U16349 ( .A(n16076), .Z(n16024) );
  NOR U16350 ( .A(n16075), .B(n16024), .Z(n16078) );
  IV U16351 ( .A(n16025), .Z(n16027) );
  XOR U16352 ( .A(n16027), .B(n16026), .Z(n16071) );
  NOR U16353 ( .A(n98), .B(n56), .Z(n16072) );
  IV U16354 ( .A(n16072), .Z(n16028) );
  NOR U16355 ( .A(n16071), .B(n16028), .Z(n16074) );
  XOR U16356 ( .A(n16030), .B(n16029), .Z(n16067) );
  NOR U16357 ( .A(n91), .B(n56), .Z(n16068) );
  IV U16358 ( .A(n16068), .Z(n16031) );
  NOR U16359 ( .A(n16067), .B(n16031), .Z(n16070) );
  IV U16360 ( .A(n16032), .Z(n16034) );
  XOR U16361 ( .A(n16034), .B(n16033), .Z(n16063) );
  NOR U16362 ( .A(n97), .B(n56), .Z(n16064) );
  IV U16363 ( .A(n16064), .Z(n16035) );
  NOR U16364 ( .A(n16063), .B(n16035), .Z(n16066) );
  XOR U16365 ( .A(n16037), .B(n16036), .Z(n16059) );
  IV U16366 ( .A(n16059), .Z(n16039) );
  NOR U16367 ( .A(n96), .B(n56), .Z(n16038) );
  IV U16368 ( .A(n16038), .Z(n16060) );
  NOR U16369 ( .A(n16039), .B(n16060), .Z(n16062) );
  NOR U16370 ( .A(n95), .B(n56), .Z(n16056) );
  IV U16371 ( .A(n16056), .Z(n16042) );
  XOR U16372 ( .A(n16041), .B(n16040), .Z(n16055) );
  NOR U16373 ( .A(n16042), .B(n16055), .Z(n16058) );
  NOR U16374 ( .A(n56), .B(n93), .Z(n17068) );
  IV U16375 ( .A(n17068), .Z(n16043) );
  NOR U16376 ( .A(n55), .B(n168), .Z(n16051) );
  IV U16377 ( .A(n16051), .Z(n16046) );
  NOR U16378 ( .A(n16043), .B(n16046), .Z(n16044) );
  IV U16379 ( .A(n16044), .Z(n16045) );
  NOR U16380 ( .A(n94), .B(n16045), .Z(n16054) );
  NOR U16381 ( .A(n16046), .B(n93), .Z(n16047) );
  XOR U16382 ( .A(n94), .B(n16047), .Z(n16048) );
  NOR U16383 ( .A(n56), .B(n16048), .Z(n16049) );
  IV U16384 ( .A(n16049), .Z(n16521) );
  XOR U16385 ( .A(n16051), .B(n16050), .Z(n16520) );
  IV U16386 ( .A(n16520), .Z(n16052) );
  NOR U16387 ( .A(n16521), .B(n16052), .Z(n16053) );
  NOR U16388 ( .A(n16054), .B(n16053), .Z(n16517) );
  XOR U16389 ( .A(n16056), .B(n16055), .Z(n16516) );
  NOR U16390 ( .A(n16517), .B(n16516), .Z(n16057) );
  NOR U16391 ( .A(n16058), .B(n16057), .Z(n16544) );
  XOR U16392 ( .A(n16060), .B(n16059), .Z(n16543) );
  NOR U16393 ( .A(n16544), .B(n16543), .Z(n16061) );
  NOR U16394 ( .A(n16062), .B(n16061), .Z(n16512) );
  XOR U16395 ( .A(n16064), .B(n16063), .Z(n16513) );
  NOR U16396 ( .A(n16512), .B(n16513), .Z(n16065) );
  NOR U16397 ( .A(n16066), .B(n16065), .Z(n16508) );
  XOR U16398 ( .A(n16068), .B(n16067), .Z(n16509) );
  NOR U16399 ( .A(n16508), .B(n16509), .Z(n16069) );
  NOR U16400 ( .A(n16070), .B(n16069), .Z(n16504) );
  XOR U16401 ( .A(n16072), .B(n16071), .Z(n16505) );
  NOR U16402 ( .A(n16504), .B(n16505), .Z(n16073) );
  NOR U16403 ( .A(n16074), .B(n16073), .Z(n16500) );
  XOR U16404 ( .A(n16076), .B(n16075), .Z(n16501) );
  NOR U16405 ( .A(n16500), .B(n16501), .Z(n16077) );
  NOR U16406 ( .A(n16078), .B(n16077), .Z(n16496) );
  XOR U16407 ( .A(n16080), .B(n16079), .Z(n16497) );
  NOR U16408 ( .A(n16496), .B(n16497), .Z(n16081) );
  NOR U16409 ( .A(n16082), .B(n16081), .Z(n16492) );
  XOR U16410 ( .A(n16084), .B(n16083), .Z(n16493) );
  NOR U16411 ( .A(n16492), .B(n16493), .Z(n16085) );
  NOR U16412 ( .A(n16086), .B(n16085), .Z(n16488) );
  XOR U16413 ( .A(n16088), .B(n16087), .Z(n16489) );
  NOR U16414 ( .A(n16488), .B(n16489), .Z(n16089) );
  NOR U16415 ( .A(n16090), .B(n16089), .Z(n16484) );
  XOR U16416 ( .A(n16092), .B(n16091), .Z(n16485) );
  NOR U16417 ( .A(n16484), .B(n16485), .Z(n16093) );
  NOR U16418 ( .A(n16094), .B(n16093), .Z(n16481) );
  XOR U16419 ( .A(n16096), .B(n16095), .Z(n16480) );
  NOR U16420 ( .A(n16481), .B(n16480), .Z(n16097) );
  NOR U16421 ( .A(n16098), .B(n16097), .Z(n16476) );
  XOR U16422 ( .A(n16100), .B(n16099), .Z(n16477) );
  NOR U16423 ( .A(n16476), .B(n16477), .Z(n16101) );
  NOR U16424 ( .A(n16102), .B(n16101), .Z(n16472) );
  XOR U16425 ( .A(n16104), .B(n16103), .Z(n16473) );
  NOR U16426 ( .A(n16472), .B(n16473), .Z(n16105) );
  NOR U16427 ( .A(n16106), .B(n16105), .Z(n16596) );
  XOR U16428 ( .A(n16108), .B(n16107), .Z(n16595) );
  NOR U16429 ( .A(n16596), .B(n16595), .Z(n16109) );
  NOR U16430 ( .A(n16110), .B(n16109), .Z(n16468) );
  XOR U16431 ( .A(n16112), .B(n16111), .Z(n16469) );
  NOR U16432 ( .A(n16468), .B(n16469), .Z(n16113) );
  NOR U16433 ( .A(n16114), .B(n16113), .Z(n16609) );
  XOR U16434 ( .A(n16116), .B(n16115), .Z(n16608) );
  NOR U16435 ( .A(n16609), .B(n16608), .Z(n16117) );
  NOR U16436 ( .A(n16118), .B(n16117), .Z(n16464) );
  XOR U16437 ( .A(n16120), .B(n16119), .Z(n16465) );
  NOR U16438 ( .A(n16464), .B(n16465), .Z(n16121) );
  NOR U16439 ( .A(n16122), .B(n16121), .Z(n16123) );
  IV U16440 ( .A(n16123), .Z(n16463) );
  XOR U16441 ( .A(n16125), .B(n16124), .Z(n16126) );
  IV U16442 ( .A(n16126), .Z(n16462) );
  NOR U16443 ( .A(n16463), .B(n16462), .Z(n16127) );
  NOR U16444 ( .A(n16128), .B(n16127), .Z(n16460) );
  IV U16445 ( .A(n16460), .Z(n16131) );
  XOR U16446 ( .A(n16130), .B(n16129), .Z(n16459) );
  NOR U16447 ( .A(n16131), .B(n16459), .Z(n16132) );
  NOR U16448 ( .A(n16133), .B(n16132), .Z(n16134) );
  IV U16449 ( .A(n16134), .Z(n16456) );
  NOR U16450 ( .A(n16457), .B(n16456), .Z(n16135) );
  NOR U16451 ( .A(n16136), .B(n16135), .Z(n16137) );
  IV U16452 ( .A(n16137), .Z(n16455) );
  XOR U16453 ( .A(n16139), .B(n16138), .Z(n16454) );
  NOR U16454 ( .A(n16455), .B(n16454), .Z(n16140) );
  NOR U16455 ( .A(n16141), .B(n16140), .Z(n16452) );
  NOR U16456 ( .A(n16143), .B(n16142), .Z(n16144) );
  NOR U16457 ( .A(n16452), .B(n16144), .Z(n16145) );
  NOR U16458 ( .A(n16146), .B(n16145), .Z(n16151) );
  NOR U16459 ( .A(n111), .B(n56), .Z(n16150) );
  IV U16460 ( .A(n16150), .Z(n16147) );
  NOR U16461 ( .A(n16151), .B(n16147), .Z(n16153) );
  XOR U16462 ( .A(n16149), .B(n16148), .Z(n16447) );
  XOR U16463 ( .A(n16151), .B(n16150), .Z(n16448) );
  NOR U16464 ( .A(n16447), .B(n16448), .Z(n16152) );
  NOR U16465 ( .A(n16153), .B(n16152), .Z(n16652) );
  XOR U16466 ( .A(n16155), .B(n16154), .Z(n16653) );
  NOR U16467 ( .A(n16652), .B(n16653), .Z(n16156) );
  NOR U16468 ( .A(n16157), .B(n16156), .Z(n16443) );
  XOR U16469 ( .A(n16159), .B(n16158), .Z(n16444) );
  NOR U16470 ( .A(n16443), .B(n16444), .Z(n16160) );
  NOR U16471 ( .A(n16161), .B(n16160), .Z(n16441) );
  IV U16472 ( .A(n16441), .Z(n16162) );
  NOR U16473 ( .A(n16163), .B(n16162), .Z(n16164) );
  NOR U16474 ( .A(n16165), .B(n16164), .Z(n16166) );
  IV U16475 ( .A(n16166), .Z(n16173) );
  NOR U16476 ( .A(n113), .B(n56), .Z(n16172) );
  IV U16477 ( .A(n16172), .Z(n16167) );
  NOR U16478 ( .A(n16173), .B(n16167), .Z(n16175) );
  XOR U16479 ( .A(n16169), .B(n16168), .Z(n16170) );
  XOR U16480 ( .A(n16171), .B(n16170), .Z(n16434) );
  XOR U16481 ( .A(n16173), .B(n16172), .Z(n16435) );
  NOR U16482 ( .A(n16434), .B(n16435), .Z(n16174) );
  NOR U16483 ( .A(n16175), .B(n16174), .Z(n16674) );
  NOR U16484 ( .A(n16177), .B(n16176), .Z(n16178) );
  NOR U16485 ( .A(n16674), .B(n16178), .Z(n16179) );
  NOR U16486 ( .A(n16180), .B(n16179), .Z(n16187) );
  NOR U16487 ( .A(n114), .B(n56), .Z(n16186) );
  IV U16488 ( .A(n16186), .Z(n16181) );
  NOR U16489 ( .A(n16187), .B(n16181), .Z(n16189) );
  XOR U16490 ( .A(n16183), .B(n16182), .Z(n16184) );
  XOR U16491 ( .A(n16185), .B(n16184), .Z(n16433) );
  XOR U16492 ( .A(n16187), .B(n16186), .Z(n16432) );
  NOR U16493 ( .A(n16433), .B(n16432), .Z(n16188) );
  NOR U16494 ( .A(n16189), .B(n16188), .Z(n16688) );
  NOR U16495 ( .A(n16190), .B(n16688), .Z(n16191) );
  NOR U16496 ( .A(n16192), .B(n16191), .Z(n16199) );
  NOR U16497 ( .A(n115), .B(n56), .Z(n16198) );
  IV U16498 ( .A(n16198), .Z(n16193) );
  NOR U16499 ( .A(n16199), .B(n16193), .Z(n16201) );
  XOR U16500 ( .A(n16195), .B(n16194), .Z(n16196) );
  XOR U16501 ( .A(n16197), .B(n16196), .Z(n16429) );
  XOR U16502 ( .A(n16199), .B(n16198), .Z(n16428) );
  NOR U16503 ( .A(n16429), .B(n16428), .Z(n16200) );
  NOR U16504 ( .A(n16201), .B(n16200), .Z(n16702) );
  NOR U16505 ( .A(n16202), .B(n16702), .Z(n16203) );
  NOR U16506 ( .A(n16204), .B(n16203), .Z(n16208) );
  NOR U16507 ( .A(n116), .B(n56), .Z(n16209) );
  IV U16508 ( .A(n16209), .Z(n16205) );
  NOR U16509 ( .A(n16208), .B(n16205), .Z(n16211) );
  XOR U16510 ( .A(n16207), .B(n16206), .Z(n16425) );
  XOR U16511 ( .A(n16209), .B(n16208), .Z(n16424) );
  NOR U16512 ( .A(n16425), .B(n16424), .Z(n16210) );
  NOR U16513 ( .A(n16211), .B(n16210), .Z(n16715) );
  IV U16514 ( .A(n16715), .Z(n16212) );
  NOR U16515 ( .A(n16213), .B(n16212), .Z(n16214) );
  NOR U16516 ( .A(n16215), .B(n16214), .Z(n16221) );
  IV U16517 ( .A(n16221), .Z(n16216) );
  NOR U16518 ( .A(n16222), .B(n16216), .Z(n16224) );
  XOR U16519 ( .A(n16218), .B(n16217), .Z(n16219) );
  XOR U16520 ( .A(n16220), .B(n16219), .Z(n16420) );
  XOR U16521 ( .A(n16222), .B(n16221), .Z(n16419) );
  NOR U16522 ( .A(n16420), .B(n16419), .Z(n16223) );
  NOR U16523 ( .A(n16224), .B(n16223), .Z(n16729) );
  NOR U16524 ( .A(n16226), .B(n16225), .Z(n16227) );
  NOR U16525 ( .A(n16729), .B(n16227), .Z(n16228) );
  NOR U16526 ( .A(n16229), .B(n16228), .Z(n16236) );
  NOR U16527 ( .A(n119), .B(n56), .Z(n16235) );
  IV U16528 ( .A(n16235), .Z(n16230) );
  NOR U16529 ( .A(n16236), .B(n16230), .Z(n16238) );
  XOR U16530 ( .A(n16232), .B(n16231), .Z(n16233) );
  XOR U16531 ( .A(n16234), .B(n16233), .Z(n16418) );
  XOR U16532 ( .A(n16236), .B(n16235), .Z(n16417) );
  NOR U16533 ( .A(n16418), .B(n16417), .Z(n16237) );
  NOR U16534 ( .A(n16238), .B(n16237), .Z(n16743) );
  XOR U16535 ( .A(n16240), .B(n16239), .Z(n16742) );
  NOR U16536 ( .A(n16743), .B(n16742), .Z(n16241) );
  NOR U16537 ( .A(n16242), .B(n16241), .Z(n16249) );
  XOR U16538 ( .A(n16244), .B(n16243), .Z(n16245) );
  XOR U16539 ( .A(n16246), .B(n16245), .Z(n16248) );
  IV U16540 ( .A(n16248), .Z(n16247) );
  NOR U16541 ( .A(n16249), .B(n16247), .Z(n16252) );
  XOR U16542 ( .A(n16249), .B(n16248), .Z(n16749) );
  NOR U16543 ( .A(n123), .B(n56), .Z(n16748) );
  IV U16544 ( .A(n16748), .Z(n16250) );
  NOR U16545 ( .A(n16749), .B(n16250), .Z(n16251) );
  NOR U16546 ( .A(n16252), .B(n16251), .Z(n16253) );
  IV U16547 ( .A(n16253), .Z(n16754) );
  NOR U16548 ( .A(n16254), .B(n16754), .Z(n16255) );
  NOR U16549 ( .A(n16256), .B(n16255), .Z(n16257) );
  IV U16550 ( .A(n16257), .Z(n16264) );
  NOR U16551 ( .A(n126), .B(n56), .Z(n16263) );
  IV U16552 ( .A(n16263), .Z(n16258) );
  NOR U16553 ( .A(n16264), .B(n16258), .Z(n16266) );
  XOR U16554 ( .A(n16260), .B(n16259), .Z(n16261) );
  XOR U16555 ( .A(n16262), .B(n16261), .Z(n16414) );
  XOR U16556 ( .A(n16264), .B(n16263), .Z(n16413) );
  NOR U16557 ( .A(n16414), .B(n16413), .Z(n16265) );
  NOR U16558 ( .A(n16266), .B(n16265), .Z(n16272) );
  XOR U16559 ( .A(n16268), .B(n16267), .Z(n16269) );
  XOR U16560 ( .A(n16270), .B(n16269), .Z(n16271) );
  NOR U16561 ( .A(n16272), .B(n16271), .Z(n16276) );
  XOR U16562 ( .A(n16272), .B(n16271), .Z(n16773) );
  IV U16563 ( .A(n16773), .Z(n16274) );
  NOR U16564 ( .A(n128), .B(n56), .Z(n16273) );
  IV U16565 ( .A(n16273), .Z(n16772) );
  NOR U16566 ( .A(n16274), .B(n16772), .Z(n16275) );
  NOR U16567 ( .A(n16276), .B(n16275), .Z(n16412) );
  XOR U16568 ( .A(n16278), .B(n16277), .Z(n16411) );
  NOR U16569 ( .A(n16412), .B(n16411), .Z(n16279) );
  NOR U16570 ( .A(n16280), .B(n16279), .Z(n16287) );
  NOR U16571 ( .A(n133), .B(n56), .Z(n16286) );
  IV U16572 ( .A(n16286), .Z(n16281) );
  NOR U16573 ( .A(n16287), .B(n16281), .Z(n16289) );
  XOR U16574 ( .A(n16283), .B(n16282), .Z(n16284) );
  XOR U16575 ( .A(n16285), .B(n16284), .Z(n16784) );
  XOR U16576 ( .A(n16287), .B(n16286), .Z(n16783) );
  NOR U16577 ( .A(n16784), .B(n16783), .Z(n16288) );
  NOR U16578 ( .A(n16289), .B(n16288), .Z(n16291) );
  IV U16579 ( .A(n16291), .Z(n16790) );
  NOR U16580 ( .A(n16290), .B(n16790), .Z(n16294) );
  IV U16581 ( .A(n16290), .Z(n16791) );
  NOR U16582 ( .A(n16291), .B(n16791), .Z(n16292) );
  NOR U16583 ( .A(n135), .B(n56), .Z(n16793) );
  NOR U16584 ( .A(n16292), .B(n16793), .Z(n16293) );
  NOR U16585 ( .A(n16294), .B(n16293), .Z(n16295) );
  IV U16586 ( .A(n16295), .Z(n16298) );
  NOR U16587 ( .A(n137), .B(n56), .Z(n16297) );
  IV U16588 ( .A(n16297), .Z(n16296) );
  NOR U16589 ( .A(n16298), .B(n16296), .Z(n16302) );
  XOR U16590 ( .A(n16298), .B(n16297), .Z(n16800) );
  XOR U16591 ( .A(n16300), .B(n16299), .Z(n16799) );
  NOR U16592 ( .A(n16800), .B(n16799), .Z(n16301) );
  NOR U16593 ( .A(n16302), .B(n16301), .Z(n16307) );
  NOR U16594 ( .A(n139), .B(n56), .Z(n16306) );
  IV U16595 ( .A(n16306), .Z(n16303) );
  NOR U16596 ( .A(n16307), .B(n16303), .Z(n16310) );
  XOR U16597 ( .A(n16305), .B(n16304), .Z(n16807) );
  IV U16598 ( .A(n16807), .Z(n16308) );
  XOR U16599 ( .A(n16307), .B(n16306), .Z(n16806) );
  NOR U16600 ( .A(n16308), .B(n16806), .Z(n16309) );
  NOR U16601 ( .A(n16310), .B(n16309), .Z(n16314) );
  XOR U16602 ( .A(n16312), .B(n16311), .Z(n16313) );
  NOR U16603 ( .A(n16314), .B(n16313), .Z(n16318) );
  XOR U16604 ( .A(n16314), .B(n16313), .Z(n16818) );
  IV U16605 ( .A(n16818), .Z(n16316) );
  NOR U16606 ( .A(n141), .B(n56), .Z(n16315) );
  IV U16607 ( .A(n16315), .Z(n16817) );
  NOR U16608 ( .A(n16316), .B(n16817), .Z(n16317) );
  NOR U16609 ( .A(n16318), .B(n16317), .Z(n16321) );
  NOR U16610 ( .A(n143), .B(n56), .Z(n16320) );
  IV U16611 ( .A(n16320), .Z(n16319) );
  NOR U16612 ( .A(n16321), .B(n16319), .Z(n16325) );
  XOR U16613 ( .A(n16321), .B(n16320), .Z(n16825) );
  XOR U16614 ( .A(n16323), .B(n16322), .Z(n16824) );
  NOR U16615 ( .A(n16825), .B(n16824), .Z(n16324) );
  NOR U16616 ( .A(n16325), .B(n16324), .Z(n16330) );
  NOR U16617 ( .A(n145), .B(n56), .Z(n16329) );
  IV U16618 ( .A(n16329), .Z(n16326) );
  NOR U16619 ( .A(n16330), .B(n16326), .Z(n16333) );
  XOR U16620 ( .A(n16328), .B(n16327), .Z(n16830) );
  IV U16621 ( .A(n16830), .Z(n16331) );
  XOR U16622 ( .A(n16330), .B(n16329), .Z(n16829) );
  NOR U16623 ( .A(n16331), .B(n16829), .Z(n16332) );
  NOR U16624 ( .A(n16333), .B(n16332), .Z(n16337) );
  XOR U16625 ( .A(n16335), .B(n16334), .Z(n16336) );
  NOR U16626 ( .A(n16337), .B(n16336), .Z(n16341) );
  XOR U16627 ( .A(n16337), .B(n16336), .Z(n16841) );
  IV U16628 ( .A(n16841), .Z(n16339) );
  NOR U16629 ( .A(n147), .B(n56), .Z(n16338) );
  IV U16630 ( .A(n16338), .Z(n16840) );
  NOR U16631 ( .A(n16339), .B(n16840), .Z(n16340) );
  NOR U16632 ( .A(n16341), .B(n16340), .Z(n16344) );
  NOR U16633 ( .A(n148), .B(n56), .Z(n16343) );
  IV U16634 ( .A(n16343), .Z(n16342) );
  NOR U16635 ( .A(n16344), .B(n16342), .Z(n16348) );
  XOR U16636 ( .A(n16344), .B(n16343), .Z(n16846) );
  XOR U16637 ( .A(n16346), .B(n16345), .Z(n16845) );
  NOR U16638 ( .A(n16846), .B(n16845), .Z(n16347) );
  NOR U16639 ( .A(n16348), .B(n16347), .Z(n16351) );
  NOR U16640 ( .A(n150), .B(n56), .Z(n16350) );
  IV U16641 ( .A(n16350), .Z(n16349) );
  NOR U16642 ( .A(n16351), .B(n16349), .Z(n16356) );
  XOR U16643 ( .A(n16351), .B(n16350), .Z(n16853) );
  XOR U16644 ( .A(n16353), .B(n16352), .Z(n16852) );
  IV U16645 ( .A(n16852), .Z(n16354) );
  NOR U16646 ( .A(n16853), .B(n16354), .Z(n16355) );
  NOR U16647 ( .A(n16356), .B(n16355), .Z(n16360) );
  XOR U16648 ( .A(n16358), .B(n16357), .Z(n16359) );
  NOR U16649 ( .A(n16360), .B(n16359), .Z(n16364) );
  XOR U16650 ( .A(n16360), .B(n16359), .Z(n16409) );
  IV U16651 ( .A(n16409), .Z(n16362) );
  NOR U16652 ( .A(n153), .B(n56), .Z(n16361) );
  IV U16653 ( .A(n16361), .Z(n16408) );
  NOR U16654 ( .A(n16362), .B(n16408), .Z(n16363) );
  NOR U16655 ( .A(n16364), .B(n16363), .Z(n16367) );
  NOR U16656 ( .A(n155), .B(n56), .Z(n16366) );
  IV U16657 ( .A(n16366), .Z(n16365) );
  NOR U16658 ( .A(n16367), .B(n16365), .Z(n16371) );
  XOR U16659 ( .A(n16367), .B(n16366), .Z(n16866) );
  XOR U16660 ( .A(n16369), .B(n16368), .Z(n16865) );
  NOR U16661 ( .A(n16866), .B(n16865), .Z(n16370) );
  NOR U16662 ( .A(n16371), .B(n16370), .Z(n16376) );
  NOR U16663 ( .A(n156), .B(n56), .Z(n16375) );
  IV U16664 ( .A(n16375), .Z(n16372) );
  NOR U16665 ( .A(n16376), .B(n16372), .Z(n16378) );
  XOR U16666 ( .A(n16374), .B(n16373), .Z(n16873) );
  XOR U16667 ( .A(n16376), .B(n16375), .Z(n16872) );
  NOR U16668 ( .A(n16873), .B(n16872), .Z(n16377) );
  NOR U16669 ( .A(n16378), .B(n16377), .Z(n16382) );
  XOR U16670 ( .A(n16380), .B(n16379), .Z(n16381) );
  NOR U16671 ( .A(n16382), .B(n16381), .Z(n16386) );
  XOR U16672 ( .A(n16382), .B(n16381), .Z(n16884) );
  IV U16673 ( .A(n16884), .Z(n16384) );
  NOR U16674 ( .A(n158), .B(n56), .Z(n16383) );
  IV U16675 ( .A(n16383), .Z(n16883) );
  NOR U16676 ( .A(n16384), .B(n16883), .Z(n16385) );
  NOR U16677 ( .A(n16386), .B(n16385), .Z(n16388) );
  IV U16678 ( .A(n16388), .Z(n16888) );
  NOR U16679 ( .A(n16387), .B(n16888), .Z(n16393) );
  IV U16680 ( .A(n16387), .Z(n16889) );
  NOR U16681 ( .A(n16388), .B(n16889), .Z(n16391) );
  XOR U16682 ( .A(n16390), .B(n16389), .Z(n16891) );
  NOR U16683 ( .A(n16391), .B(n16891), .Z(n16392) );
  NOR U16684 ( .A(n16393), .B(n16392), .Z(n16401) );
  IV U16685 ( .A(n16401), .Z(n16395) );
  NOR U16686 ( .A(n163), .B(n56), .Z(n16394) );
  IV U16687 ( .A(n16394), .Z(n16400) );
  NOR U16688 ( .A(n16395), .B(n16400), .Z(n16403) );
  XOR U16689 ( .A(n16397), .B(n16396), .Z(n16398) );
  XOR U16690 ( .A(n16399), .B(n16398), .Z(n16897) );
  XOR U16691 ( .A(n16401), .B(n16400), .Z(n16896) );
  NOR U16692 ( .A(n16897), .B(n16896), .Z(n16402) );
  NOR U16693 ( .A(n16403), .B(n16402), .Z(n16911) );
  IV U16694 ( .A(n16911), .Z(n16406) );
  XOR U16695 ( .A(n16405), .B(n16404), .Z(n16910) );
  XOR U16696 ( .A(n16406), .B(n16910), .Z(n16914) );
  XOR U16697 ( .A(n16912), .B(n16914), .Z(n16904) );
  NOR U16698 ( .A(n167), .B(n57), .Z(n16905) );
  IV U16699 ( .A(n16905), .Z(n16407) );
  NOR U16700 ( .A(n16904), .B(n16407), .Z(n16907) );
  XOR U16701 ( .A(n16409), .B(n16408), .Z(n16861) );
  NOR U16702 ( .A(n155), .B(n57), .Z(n16860) );
  IV U16703 ( .A(n16860), .Z(n16410) );
  NOR U16704 ( .A(n16861), .B(n16410), .Z(n16863) );
  NOR U16705 ( .A(n135), .B(n57), .Z(n16781) );
  XOR U16706 ( .A(n16412), .B(n16411), .Z(n16776) );
  NOR U16707 ( .A(n128), .B(n57), .Z(n16415) );
  XOR U16708 ( .A(n16414), .B(n16413), .Z(n16416) );
  NOR U16709 ( .A(n16415), .B(n16416), .Z(n16767) );
  IV U16710 ( .A(n16415), .Z(n17298) );
  IV U16711 ( .A(n16416), .Z(n17297) );
  NOR U16712 ( .A(n17298), .B(n17297), .Z(n16765) );
  XOR U16713 ( .A(n16418), .B(n16417), .Z(n16735) );
  IV U16714 ( .A(n16735), .Z(n17271) );
  NOR U16715 ( .A(n120), .B(n57), .Z(n16734) );
  IV U16716 ( .A(n16734), .Z(n17270) );
  NOR U16717 ( .A(n17271), .B(n17270), .Z(n16738) );
  NOR U16718 ( .A(n119), .B(n57), .Z(n16731) );
  IV U16719 ( .A(n16731), .Z(n16725) );
  NOR U16720 ( .A(n79), .B(n57), .Z(n16421) );
  XOR U16721 ( .A(n16420), .B(n16419), .Z(n16422) );
  NOR U16722 ( .A(n16421), .B(n16422), .Z(n16723) );
  IV U16723 ( .A(n16421), .Z(n17257) );
  IV U16724 ( .A(n16422), .Z(n17256) );
  NOR U16725 ( .A(n17257), .B(n17256), .Z(n16721) );
  NOR U16726 ( .A(n117), .B(n57), .Z(n16423) );
  IV U16727 ( .A(n16423), .Z(n16717) );
  NOR U16728 ( .A(n80), .B(n57), .Z(n16426) );
  XOR U16729 ( .A(n16425), .B(n16424), .Z(n16427) );
  NOR U16730 ( .A(n16426), .B(n16427), .Z(n16710) );
  IV U16731 ( .A(n16426), .Z(n17243) );
  IV U16732 ( .A(n16427), .Z(n17242) );
  NOR U16733 ( .A(n17243), .B(n17242), .Z(n16708) );
  NOR U16734 ( .A(n81), .B(n57), .Z(n16430) );
  XOR U16735 ( .A(n16429), .B(n16428), .Z(n16431) );
  NOR U16736 ( .A(n16430), .B(n16431), .Z(n16696) );
  IV U16737 ( .A(n16430), .Z(n17229) );
  IV U16738 ( .A(n16431), .Z(n17228) );
  NOR U16739 ( .A(n17229), .B(n17228), .Z(n16694) );
  XOR U16740 ( .A(n16433), .B(n16432), .Z(n16680) );
  IV U16741 ( .A(n16680), .Z(n17215) );
  NOR U16742 ( .A(n82), .B(n57), .Z(n16679) );
  IV U16743 ( .A(n16679), .Z(n17214) );
  NOR U16744 ( .A(n17215), .B(n17214), .Z(n16683) );
  XOR U16745 ( .A(n16435), .B(n16434), .Z(n16436) );
  NOR U16746 ( .A(n83), .B(n57), .Z(n16437) );
  NOR U16747 ( .A(n16436), .B(n16437), .Z(n16668) );
  IV U16748 ( .A(n16436), .Z(n16966) );
  IV U16749 ( .A(n16437), .Z(n16965) );
  NOR U16750 ( .A(n16966), .B(n16965), .Z(n16666) );
  XOR U16751 ( .A(n16439), .B(n16438), .Z(n16440) );
  XOR U16752 ( .A(n16441), .B(n16440), .Z(n16662) );
  NOR U16753 ( .A(n113), .B(n57), .Z(n16661) );
  IV U16754 ( .A(n16661), .Z(n16442) );
  NOR U16755 ( .A(n16662), .B(n16442), .Z(n16664) );
  NOR U16756 ( .A(n84), .B(n57), .Z(n16658) );
  IV U16757 ( .A(n16658), .Z(n16446) );
  IV U16758 ( .A(n16443), .Z(n16445) );
  XOR U16759 ( .A(n16445), .B(n16444), .Z(n16657) );
  NOR U16760 ( .A(n16446), .B(n16657), .Z(n16660) );
  XOR U16761 ( .A(n16448), .B(n16447), .Z(n16645) );
  IV U16762 ( .A(n16645), .Z(n16977) );
  NOR U16763 ( .A(n85), .B(n57), .Z(n16644) );
  IV U16764 ( .A(n16644), .Z(n16976) );
  NOR U16765 ( .A(n16977), .B(n16976), .Z(n16648) );
  XOR U16766 ( .A(n16450), .B(n16449), .Z(n16451) );
  XOR U16767 ( .A(n16452), .B(n16451), .Z(n16641) );
  NOR U16768 ( .A(n111), .B(n57), .Z(n16640) );
  IV U16769 ( .A(n16640), .Z(n16453) );
  NOR U16770 ( .A(n16641), .B(n16453), .Z(n16643) );
  NOR U16771 ( .A(n86), .B(n57), .Z(n16635) );
  XOR U16772 ( .A(n16455), .B(n16454), .Z(n16634) );
  NOR U16773 ( .A(n16635), .B(n16634), .Z(n16638) );
  XOR U16774 ( .A(n16457), .B(n16456), .Z(n16630) );
  NOR U16775 ( .A(n110), .B(n57), .Z(n16629) );
  IV U16776 ( .A(n16629), .Z(n16458) );
  NOR U16777 ( .A(n16630), .B(n16458), .Z(n16632) );
  XOR U16778 ( .A(n16460), .B(n16459), .Z(n16625) );
  NOR U16779 ( .A(n109), .B(n57), .Z(n16626) );
  IV U16780 ( .A(n16626), .Z(n16461) );
  NOR U16781 ( .A(n16625), .B(n16461), .Z(n16628) );
  XOR U16782 ( .A(n16463), .B(n16462), .Z(n16620) );
  IV U16783 ( .A(n16464), .Z(n16466) );
  XOR U16784 ( .A(n16466), .B(n16465), .Z(n16615) );
  NOR U16785 ( .A(n87), .B(n57), .Z(n16616) );
  IV U16786 ( .A(n16616), .Z(n16467) );
  NOR U16787 ( .A(n16615), .B(n16467), .Z(n16618) );
  IV U16788 ( .A(n16468), .Z(n16470) );
  XOR U16789 ( .A(n16470), .B(n16469), .Z(n16603) );
  NOR U16790 ( .A(n88), .B(n57), .Z(n16604) );
  IV U16791 ( .A(n16604), .Z(n16471) );
  NOR U16792 ( .A(n16603), .B(n16471), .Z(n16606) );
  IV U16793 ( .A(n16472), .Z(n16474) );
  XOR U16794 ( .A(n16474), .B(n16473), .Z(n16591) );
  NOR U16795 ( .A(n105), .B(n57), .Z(n16592) );
  IV U16796 ( .A(n16592), .Z(n16475) );
  NOR U16797 ( .A(n16591), .B(n16475), .Z(n16594) );
  IV U16798 ( .A(n16476), .Z(n16478) );
  XOR U16799 ( .A(n16478), .B(n16477), .Z(n16587) );
  NOR U16800 ( .A(n104), .B(n57), .Z(n16588) );
  IV U16801 ( .A(n16588), .Z(n16479) );
  NOR U16802 ( .A(n16587), .B(n16479), .Z(n16590) );
  XOR U16803 ( .A(n16481), .B(n16480), .Z(n16583) );
  IV U16804 ( .A(n16583), .Z(n16483) );
  NOR U16805 ( .A(n89), .B(n57), .Z(n16482) );
  IV U16806 ( .A(n16482), .Z(n16584) );
  NOR U16807 ( .A(n16483), .B(n16584), .Z(n16586) );
  IV U16808 ( .A(n16484), .Z(n16486) );
  XOR U16809 ( .A(n16486), .B(n16485), .Z(n16579) );
  NOR U16810 ( .A(n103), .B(n57), .Z(n16580) );
  IV U16811 ( .A(n16580), .Z(n16487) );
  NOR U16812 ( .A(n16579), .B(n16487), .Z(n16582) );
  IV U16813 ( .A(n16488), .Z(n16490) );
  XOR U16814 ( .A(n16490), .B(n16489), .Z(n16575) );
  NOR U16815 ( .A(n90), .B(n57), .Z(n16576) );
  IV U16816 ( .A(n16576), .Z(n16491) );
  NOR U16817 ( .A(n16575), .B(n16491), .Z(n16578) );
  IV U16818 ( .A(n16492), .Z(n16494) );
  XOR U16819 ( .A(n16494), .B(n16493), .Z(n16571) );
  NOR U16820 ( .A(n102), .B(n57), .Z(n16572) );
  IV U16821 ( .A(n16572), .Z(n16495) );
  NOR U16822 ( .A(n16571), .B(n16495), .Z(n16574) );
  IV U16823 ( .A(n16496), .Z(n16498) );
  XOR U16824 ( .A(n16498), .B(n16497), .Z(n16567) );
  NOR U16825 ( .A(n101), .B(n57), .Z(n16568) );
  IV U16826 ( .A(n16568), .Z(n16499) );
  NOR U16827 ( .A(n16567), .B(n16499), .Z(n16570) );
  IV U16828 ( .A(n16500), .Z(n16502) );
  XOR U16829 ( .A(n16502), .B(n16501), .Z(n16563) );
  NOR U16830 ( .A(n100), .B(n57), .Z(n16564) );
  IV U16831 ( .A(n16564), .Z(n16503) );
  NOR U16832 ( .A(n16563), .B(n16503), .Z(n16566) );
  IV U16833 ( .A(n16504), .Z(n16506) );
  XOR U16834 ( .A(n16506), .B(n16505), .Z(n16559) );
  NOR U16835 ( .A(n99), .B(n57), .Z(n16560) );
  IV U16836 ( .A(n16560), .Z(n16507) );
  NOR U16837 ( .A(n16559), .B(n16507), .Z(n16562) );
  IV U16838 ( .A(n16508), .Z(n16510) );
  XOR U16839 ( .A(n16510), .B(n16509), .Z(n16555) );
  NOR U16840 ( .A(n98), .B(n57), .Z(n16556) );
  IV U16841 ( .A(n16556), .Z(n16511) );
  NOR U16842 ( .A(n16555), .B(n16511), .Z(n16558) );
  IV U16843 ( .A(n16512), .Z(n16514) );
  XOR U16844 ( .A(n16514), .B(n16513), .Z(n16551) );
  NOR U16845 ( .A(n91), .B(n57), .Z(n16552) );
  IV U16846 ( .A(n16552), .Z(n16515) );
  NOR U16847 ( .A(n16551), .B(n16515), .Z(n16554) );
  XOR U16848 ( .A(n16517), .B(n16516), .Z(n16539) );
  IV U16849 ( .A(n16539), .Z(n16519) );
  NOR U16850 ( .A(n96), .B(n57), .Z(n16518) );
  IV U16851 ( .A(n16518), .Z(n16540) );
  NOR U16852 ( .A(n16519), .B(n16540), .Z(n16542) );
  NOR U16853 ( .A(n95), .B(n57), .Z(n16536) );
  IV U16854 ( .A(n16536), .Z(n16522) );
  XOR U16855 ( .A(n16521), .B(n16520), .Z(n16535) );
  NOR U16856 ( .A(n16522), .B(n16535), .Z(n16538) );
  NOR U16857 ( .A(n57), .B(n93), .Z(n17571) );
  IV U16858 ( .A(n17571), .Z(n16523) );
  NOR U16859 ( .A(n56), .B(n168), .Z(n16531) );
  IV U16860 ( .A(n16531), .Z(n16526) );
  NOR U16861 ( .A(n16523), .B(n16526), .Z(n16524) );
  IV U16862 ( .A(n16524), .Z(n16525) );
  NOR U16863 ( .A(n94), .B(n16525), .Z(n16534) );
  NOR U16864 ( .A(n16526), .B(n93), .Z(n16527) );
  XOR U16865 ( .A(n94), .B(n16527), .Z(n16528) );
  NOR U16866 ( .A(n57), .B(n16528), .Z(n16529) );
  IV U16867 ( .A(n16529), .Z(n17059) );
  XOR U16868 ( .A(n16531), .B(n16530), .Z(n17058) );
  IV U16869 ( .A(n17058), .Z(n16532) );
  NOR U16870 ( .A(n17059), .B(n16532), .Z(n16533) );
  NOR U16871 ( .A(n16534), .B(n16533), .Z(n17055) );
  XOR U16872 ( .A(n16536), .B(n16535), .Z(n17054) );
  NOR U16873 ( .A(n17055), .B(n17054), .Z(n16537) );
  NOR U16874 ( .A(n16538), .B(n16537), .Z(n17082) );
  XOR U16875 ( .A(n16540), .B(n16539), .Z(n17081) );
  NOR U16876 ( .A(n17082), .B(n17081), .Z(n16541) );
  NOR U16877 ( .A(n16542), .B(n16541), .Z(n16547) );
  XOR U16878 ( .A(n16544), .B(n16543), .Z(n16546) );
  IV U16879 ( .A(n16546), .Z(n16545) );
  NOR U16880 ( .A(n16547), .B(n16545), .Z(n16550) );
  XOR U16881 ( .A(n16547), .B(n16546), .Z(n17051) );
  NOR U16882 ( .A(n97), .B(n57), .Z(n17052) );
  IV U16883 ( .A(n17052), .Z(n16548) );
  NOR U16884 ( .A(n17051), .B(n16548), .Z(n16549) );
  NOR U16885 ( .A(n16550), .B(n16549), .Z(n17047) );
  XOR U16886 ( .A(n16552), .B(n16551), .Z(n17048) );
  NOR U16887 ( .A(n17047), .B(n17048), .Z(n16553) );
  NOR U16888 ( .A(n16554), .B(n16553), .Z(n17043) );
  XOR U16889 ( .A(n16556), .B(n16555), .Z(n17044) );
  NOR U16890 ( .A(n17043), .B(n17044), .Z(n16557) );
  NOR U16891 ( .A(n16558), .B(n16557), .Z(n17039) );
  XOR U16892 ( .A(n16560), .B(n16559), .Z(n17040) );
  NOR U16893 ( .A(n17039), .B(n17040), .Z(n16561) );
  NOR U16894 ( .A(n16562), .B(n16561), .Z(n17035) );
  XOR U16895 ( .A(n16564), .B(n16563), .Z(n17036) );
  NOR U16896 ( .A(n17035), .B(n17036), .Z(n16565) );
  NOR U16897 ( .A(n16566), .B(n16565), .Z(n17031) );
  XOR U16898 ( .A(n16568), .B(n16567), .Z(n17032) );
  NOR U16899 ( .A(n17031), .B(n17032), .Z(n16569) );
  NOR U16900 ( .A(n16570), .B(n16569), .Z(n17027) );
  XOR U16901 ( .A(n16572), .B(n16571), .Z(n17028) );
  NOR U16902 ( .A(n17027), .B(n17028), .Z(n16573) );
  NOR U16903 ( .A(n16574), .B(n16573), .Z(n17023) );
  XOR U16904 ( .A(n16576), .B(n16575), .Z(n17024) );
  NOR U16905 ( .A(n17023), .B(n17024), .Z(n16577) );
  NOR U16906 ( .A(n16578), .B(n16577), .Z(n17019) );
  XOR U16907 ( .A(n16580), .B(n16579), .Z(n17020) );
  NOR U16908 ( .A(n17019), .B(n17020), .Z(n16581) );
  NOR U16909 ( .A(n16582), .B(n16581), .Z(n17126) );
  XOR U16910 ( .A(n16584), .B(n16583), .Z(n17125) );
  NOR U16911 ( .A(n17126), .B(n17125), .Z(n16585) );
  NOR U16912 ( .A(n16586), .B(n16585), .Z(n17016) );
  XOR U16913 ( .A(n16588), .B(n16587), .Z(n17015) );
  NOR U16914 ( .A(n17016), .B(n17015), .Z(n16589) );
  NOR U16915 ( .A(n16590), .B(n16589), .Z(n17011) );
  XOR U16916 ( .A(n16592), .B(n16591), .Z(n17012) );
  NOR U16917 ( .A(n17011), .B(n17012), .Z(n16593) );
  NOR U16918 ( .A(n16594), .B(n16593), .Z(n16599) );
  XOR U16919 ( .A(n16596), .B(n16595), .Z(n16598) );
  IV U16920 ( .A(n16598), .Z(n16597) );
  NOR U16921 ( .A(n16599), .B(n16597), .Z(n16602) );
  XOR U16922 ( .A(n16599), .B(n16598), .Z(n17008) );
  NOR U16923 ( .A(n106), .B(n57), .Z(n17009) );
  IV U16924 ( .A(n17009), .Z(n16600) );
  NOR U16925 ( .A(n17008), .B(n16600), .Z(n16601) );
  NOR U16926 ( .A(n16602), .B(n16601), .Z(n17004) );
  XOR U16927 ( .A(n16604), .B(n16603), .Z(n17005) );
  NOR U16928 ( .A(n17004), .B(n17005), .Z(n16605) );
  NOR U16929 ( .A(n16606), .B(n16605), .Z(n16611) );
  NOR U16930 ( .A(n107), .B(n57), .Z(n16610) );
  IV U16931 ( .A(n16610), .Z(n16607) );
  NOR U16932 ( .A(n16611), .B(n16607), .Z(n16614) );
  XOR U16933 ( .A(n16609), .B(n16608), .Z(n17002) );
  IV U16934 ( .A(n17002), .Z(n16612) );
  XOR U16935 ( .A(n16611), .B(n16610), .Z(n17001) );
  NOR U16936 ( .A(n16612), .B(n17001), .Z(n16613) );
  NOR U16937 ( .A(n16614), .B(n16613), .Z(n16997) );
  XOR U16938 ( .A(n16616), .B(n16615), .Z(n16998) );
  NOR U16939 ( .A(n16997), .B(n16998), .Z(n16617) );
  NOR U16940 ( .A(n16618), .B(n16617), .Z(n16619) );
  NOR U16941 ( .A(n16620), .B(n16619), .Z(n16624) );
  IV U16942 ( .A(n16619), .Z(n16621) );
  XOR U16943 ( .A(n16621), .B(n16620), .Z(n16994) );
  NOR U16944 ( .A(n108), .B(n57), .Z(n16995) );
  IV U16945 ( .A(n16995), .Z(n16622) );
  NOR U16946 ( .A(n16994), .B(n16622), .Z(n16623) );
  NOR U16947 ( .A(n16624), .B(n16623), .Z(n16990) );
  XOR U16948 ( .A(n16626), .B(n16625), .Z(n16991) );
  NOR U16949 ( .A(n16990), .B(n16991), .Z(n16627) );
  NOR U16950 ( .A(n16628), .B(n16627), .Z(n16986) );
  XOR U16951 ( .A(n16630), .B(n16629), .Z(n16987) );
  NOR U16952 ( .A(n16986), .B(n16987), .Z(n16631) );
  NOR U16953 ( .A(n16632), .B(n16631), .Z(n16633) );
  IV U16954 ( .A(n16633), .Z(n16984) );
  XOR U16955 ( .A(n16635), .B(n16634), .Z(n16636) );
  IV U16956 ( .A(n16636), .Z(n16983) );
  NOR U16957 ( .A(n16984), .B(n16983), .Z(n16637) );
  NOR U16958 ( .A(n16638), .B(n16637), .Z(n16639) );
  IV U16959 ( .A(n16639), .Z(n16982) );
  XOR U16960 ( .A(n16641), .B(n16640), .Z(n16981) );
  NOR U16961 ( .A(n16982), .B(n16981), .Z(n16642) );
  NOR U16962 ( .A(n16643), .B(n16642), .Z(n16979) );
  NOR U16963 ( .A(n16645), .B(n16644), .Z(n16646) );
  NOR U16964 ( .A(n16979), .B(n16646), .Z(n16647) );
  NOR U16965 ( .A(n16648), .B(n16647), .Z(n16650) );
  NOR U16966 ( .A(n112), .B(n57), .Z(n16651) );
  IV U16967 ( .A(n16651), .Z(n16649) );
  NOR U16968 ( .A(n16650), .B(n16649), .Z(n16656) );
  XOR U16969 ( .A(n16651), .B(n16650), .Z(n16973) );
  IV U16970 ( .A(n16652), .Z(n16654) );
  XOR U16971 ( .A(n16654), .B(n16653), .Z(n16972) );
  NOR U16972 ( .A(n16973), .B(n16972), .Z(n16655) );
  NOR U16973 ( .A(n16656), .B(n16655), .Z(n17190) );
  XOR U16974 ( .A(n16658), .B(n16657), .Z(n17191) );
  NOR U16975 ( .A(n17190), .B(n17191), .Z(n16659) );
  NOR U16976 ( .A(n16660), .B(n16659), .Z(n16971) );
  XOR U16977 ( .A(n16662), .B(n16661), .Z(n16970) );
  NOR U16978 ( .A(n16971), .B(n16970), .Z(n16663) );
  NOR U16979 ( .A(n16664), .B(n16663), .Z(n16968) );
  IV U16980 ( .A(n16968), .Z(n16665) );
  NOR U16981 ( .A(n16666), .B(n16665), .Z(n16667) );
  NOR U16982 ( .A(n16668), .B(n16667), .Z(n16669) );
  IV U16983 ( .A(n16669), .Z(n16676) );
  NOR U16984 ( .A(n114), .B(n57), .Z(n16675) );
  IV U16985 ( .A(n16675), .Z(n16670) );
  NOR U16986 ( .A(n16676), .B(n16670), .Z(n16678) );
  XOR U16987 ( .A(n16672), .B(n16671), .Z(n16673) );
  XOR U16988 ( .A(n16674), .B(n16673), .Z(n16961) );
  XOR U16989 ( .A(n16676), .B(n16675), .Z(n16962) );
  NOR U16990 ( .A(n16961), .B(n16962), .Z(n16677) );
  NOR U16991 ( .A(n16678), .B(n16677), .Z(n17217) );
  NOR U16992 ( .A(n16680), .B(n16679), .Z(n16681) );
  NOR U16993 ( .A(n17217), .B(n16681), .Z(n16682) );
  NOR U16994 ( .A(n16683), .B(n16682), .Z(n16690) );
  NOR U16995 ( .A(n115), .B(n57), .Z(n16689) );
  IV U16996 ( .A(n16689), .Z(n16684) );
  NOR U16997 ( .A(n16690), .B(n16684), .Z(n16692) );
  XOR U16998 ( .A(n16686), .B(n16685), .Z(n16687) );
  XOR U16999 ( .A(n16688), .B(n16687), .Z(n16958) );
  XOR U17000 ( .A(n16690), .B(n16689), .Z(n16957) );
  NOR U17001 ( .A(n16958), .B(n16957), .Z(n16691) );
  NOR U17002 ( .A(n16692), .B(n16691), .Z(n17231) );
  IV U17003 ( .A(n17231), .Z(n16693) );
  NOR U17004 ( .A(n16694), .B(n16693), .Z(n16695) );
  NOR U17005 ( .A(n16696), .B(n16695), .Z(n16704) );
  IV U17006 ( .A(n16704), .Z(n16698) );
  NOR U17007 ( .A(n116), .B(n57), .Z(n16697) );
  IV U17008 ( .A(n16697), .Z(n16703) );
  NOR U17009 ( .A(n16698), .B(n16703), .Z(n16706) );
  XOR U17010 ( .A(n16700), .B(n16699), .Z(n16701) );
  XOR U17011 ( .A(n16702), .B(n16701), .Z(n16956) );
  XOR U17012 ( .A(n16704), .B(n16703), .Z(n16955) );
  NOR U17013 ( .A(n16956), .B(n16955), .Z(n16705) );
  NOR U17014 ( .A(n16706), .B(n16705), .Z(n17245) );
  IV U17015 ( .A(n17245), .Z(n16707) );
  NOR U17016 ( .A(n16708), .B(n16707), .Z(n16709) );
  NOR U17017 ( .A(n16710), .B(n16709), .Z(n16716) );
  IV U17018 ( .A(n16716), .Z(n16711) );
  NOR U17019 ( .A(n16717), .B(n16711), .Z(n16719) );
  XOR U17020 ( .A(n16713), .B(n16712), .Z(n16714) );
  XOR U17021 ( .A(n16715), .B(n16714), .Z(n16951) );
  XOR U17022 ( .A(n16717), .B(n16716), .Z(n16952) );
  NOR U17023 ( .A(n16951), .B(n16952), .Z(n16718) );
  NOR U17024 ( .A(n16719), .B(n16718), .Z(n17259) );
  IV U17025 ( .A(n17259), .Z(n16720) );
  NOR U17026 ( .A(n16721), .B(n16720), .Z(n16722) );
  NOR U17027 ( .A(n16723), .B(n16722), .Z(n16724) );
  IV U17028 ( .A(n16724), .Z(n16730) );
  NOR U17029 ( .A(n16725), .B(n16730), .Z(n16733) );
  XOR U17030 ( .A(n16727), .B(n16726), .Z(n16728) );
  XOR U17031 ( .A(n16729), .B(n16728), .Z(n16950) );
  XOR U17032 ( .A(n16731), .B(n16730), .Z(n16949) );
  NOR U17033 ( .A(n16950), .B(n16949), .Z(n16732) );
  NOR U17034 ( .A(n16733), .B(n16732), .Z(n17273) );
  NOR U17035 ( .A(n16735), .B(n16734), .Z(n16736) );
  NOR U17036 ( .A(n17273), .B(n16736), .Z(n16737) );
  NOR U17037 ( .A(n16738), .B(n16737), .Z(n16741) );
  NOR U17038 ( .A(n123), .B(n57), .Z(n16740) );
  IV U17039 ( .A(n16740), .Z(n16739) );
  NOR U17040 ( .A(n16741), .B(n16739), .Z(n16746) );
  XOR U17041 ( .A(n16741), .B(n16740), .Z(n16946) );
  XOR U17042 ( .A(n16743), .B(n16742), .Z(n16947) );
  IV U17043 ( .A(n16947), .Z(n16744) );
  NOR U17044 ( .A(n16946), .B(n16744), .Z(n16745) );
  NOR U17045 ( .A(n16746), .B(n16745), .Z(n16751) );
  NOR U17046 ( .A(n125), .B(n57), .Z(n16750) );
  IV U17047 ( .A(n16750), .Z(n16747) );
  NOR U17048 ( .A(n16751), .B(n16747), .Z(n16753) );
  XOR U17049 ( .A(n16749), .B(n16748), .Z(n17283) );
  XOR U17050 ( .A(n16751), .B(n16750), .Z(n17282) );
  NOR U17051 ( .A(n17283), .B(n17282), .Z(n16752) );
  NOR U17052 ( .A(n16753), .B(n16752), .Z(n16759) );
  XOR U17053 ( .A(n16755), .B(n16754), .Z(n16756) );
  XOR U17054 ( .A(n16757), .B(n16756), .Z(n16758) );
  NOR U17055 ( .A(n16759), .B(n16758), .Z(n16763) );
  XOR U17056 ( .A(n16759), .B(n16758), .Z(n17292) );
  IV U17057 ( .A(n17292), .Z(n16761) );
  NOR U17058 ( .A(n126), .B(n57), .Z(n17293) );
  IV U17059 ( .A(n17293), .Z(n16760) );
  NOR U17060 ( .A(n16761), .B(n16760), .Z(n16762) );
  NOR U17061 ( .A(n16763), .B(n16762), .Z(n16764) );
  IV U17062 ( .A(n16764), .Z(n17300) );
  NOR U17063 ( .A(n16765), .B(n17300), .Z(n16766) );
  NOR U17064 ( .A(n16767), .B(n16766), .Z(n16771) );
  IV U17065 ( .A(n16771), .Z(n16769) );
  NOR U17066 ( .A(n131), .B(n57), .Z(n16768) );
  IV U17067 ( .A(n16768), .Z(n16770) );
  NOR U17068 ( .A(n16769), .B(n16770), .Z(n16775) );
  XOR U17069 ( .A(n16771), .B(n16770), .Z(n16945) );
  XOR U17070 ( .A(n16773), .B(n16772), .Z(n16944) );
  NOR U17071 ( .A(n16945), .B(n16944), .Z(n16774) );
  NOR U17072 ( .A(n16775), .B(n16774), .Z(n16777) );
  IV U17073 ( .A(n16777), .Z(n17313) );
  NOR U17074 ( .A(n16776), .B(n17313), .Z(n16780) );
  IV U17075 ( .A(n16776), .Z(n17314) );
  NOR U17076 ( .A(n16777), .B(n17314), .Z(n16778) );
  NOR U17077 ( .A(n133), .B(n57), .Z(n17316) );
  NOR U17078 ( .A(n16778), .B(n17316), .Z(n16779) );
  NOR U17079 ( .A(n16780), .B(n16779), .Z(n16782) );
  NOR U17080 ( .A(n16781), .B(n16782), .Z(n16787) );
  IV U17081 ( .A(n16781), .Z(n17324) );
  IV U17082 ( .A(n16782), .Z(n17323) );
  NOR U17083 ( .A(n17324), .B(n17323), .Z(n16785) );
  XOR U17084 ( .A(n16784), .B(n16783), .Z(n17326) );
  NOR U17085 ( .A(n16785), .B(n17326), .Z(n16786) );
  NOR U17086 ( .A(n16787), .B(n16786), .Z(n16795) );
  IV U17087 ( .A(n16795), .Z(n16789) );
  NOR U17088 ( .A(n137), .B(n57), .Z(n16788) );
  IV U17089 ( .A(n16788), .Z(n16794) );
  NOR U17090 ( .A(n16789), .B(n16794), .Z(n16797) );
  XOR U17091 ( .A(n16791), .B(n16790), .Z(n16792) );
  XOR U17092 ( .A(n16793), .B(n16792), .Z(n17332) );
  XOR U17093 ( .A(n16795), .B(n16794), .Z(n17333) );
  NOR U17094 ( .A(n17332), .B(n17333), .Z(n16796) );
  NOR U17095 ( .A(n16797), .B(n16796), .Z(n16802) );
  NOR U17096 ( .A(n139), .B(n57), .Z(n16801) );
  IV U17097 ( .A(n16801), .Z(n16798) );
  NOR U17098 ( .A(n16802), .B(n16798), .Z(n16805) );
  XOR U17099 ( .A(n16800), .B(n16799), .Z(n16942) );
  IV U17100 ( .A(n16942), .Z(n16803) );
  XOR U17101 ( .A(n16802), .B(n16801), .Z(n16941) );
  NOR U17102 ( .A(n16803), .B(n16941), .Z(n16804) );
  NOR U17103 ( .A(n16805), .B(n16804), .Z(n16808) );
  XOR U17104 ( .A(n16807), .B(n16806), .Z(n16809) );
  NOR U17105 ( .A(n16808), .B(n16809), .Z(n16813) );
  IV U17106 ( .A(n16808), .Z(n16810) );
  XOR U17107 ( .A(n16810), .B(n16809), .Z(n16937) );
  NOR U17108 ( .A(n141), .B(n57), .Z(n16811) );
  IV U17109 ( .A(n16811), .Z(n16938) );
  NOR U17110 ( .A(n16937), .B(n16938), .Z(n16812) );
  NOR U17111 ( .A(n16813), .B(n16812), .Z(n16816) );
  NOR U17112 ( .A(n143), .B(n57), .Z(n16815) );
  IV U17113 ( .A(n16815), .Z(n16814) );
  NOR U17114 ( .A(n16816), .B(n16814), .Z(n16820) );
  XOR U17115 ( .A(n16816), .B(n16815), .Z(n17350) );
  XOR U17116 ( .A(n16818), .B(n16817), .Z(n17351) );
  NOR U17117 ( .A(n17350), .B(n17351), .Z(n16819) );
  NOR U17118 ( .A(n16820), .B(n16819), .Z(n16823) );
  NOR U17119 ( .A(n145), .B(n57), .Z(n16822) );
  IV U17120 ( .A(n16822), .Z(n16821) );
  NOR U17121 ( .A(n16823), .B(n16821), .Z(n16828) );
  XOR U17122 ( .A(n16823), .B(n16822), .Z(n17355) );
  XOR U17123 ( .A(n16825), .B(n16824), .Z(n17356) );
  IV U17124 ( .A(n17356), .Z(n16826) );
  NOR U17125 ( .A(n17355), .B(n16826), .Z(n16827) );
  NOR U17126 ( .A(n16828), .B(n16827), .Z(n16831) );
  XOR U17127 ( .A(n16830), .B(n16829), .Z(n16832) );
  NOR U17128 ( .A(n16831), .B(n16832), .Z(n16836) );
  IV U17129 ( .A(n16831), .Z(n16833) );
  XOR U17130 ( .A(n16833), .B(n16832), .Z(n16934) );
  NOR U17131 ( .A(n147), .B(n57), .Z(n16935) );
  IV U17132 ( .A(n16935), .Z(n16834) );
  NOR U17133 ( .A(n16934), .B(n16834), .Z(n16835) );
  NOR U17134 ( .A(n16836), .B(n16835), .Z(n16839) );
  NOR U17135 ( .A(n148), .B(n57), .Z(n16838) );
  IV U17136 ( .A(n16838), .Z(n16837) );
  NOR U17137 ( .A(n16839), .B(n16837), .Z(n16843) );
  XOR U17138 ( .A(n16839), .B(n16838), .Z(n17370) );
  XOR U17139 ( .A(n16841), .B(n16840), .Z(n17371) );
  NOR U17140 ( .A(n17370), .B(n17371), .Z(n16842) );
  NOR U17141 ( .A(n16843), .B(n16842), .Z(n16848) );
  NOR U17142 ( .A(n150), .B(n57), .Z(n16847) );
  IV U17143 ( .A(n16847), .Z(n16844) );
  NOR U17144 ( .A(n16848), .B(n16844), .Z(n16851) );
  XOR U17145 ( .A(n16846), .B(n16845), .Z(n17376) );
  IV U17146 ( .A(n17376), .Z(n16849) );
  XOR U17147 ( .A(n16848), .B(n16847), .Z(n17375) );
  NOR U17148 ( .A(n16849), .B(n17375), .Z(n16850) );
  NOR U17149 ( .A(n16851), .B(n16850), .Z(n16854) );
  XOR U17150 ( .A(n16853), .B(n16852), .Z(n16855) );
  NOR U17151 ( .A(n16854), .B(n16855), .Z(n16859) );
  IV U17152 ( .A(n16854), .Z(n16856) );
  XOR U17153 ( .A(n16856), .B(n16855), .Z(n17386) );
  NOR U17154 ( .A(n153), .B(n57), .Z(n17387) );
  IV U17155 ( .A(n17387), .Z(n16857) );
  NOR U17156 ( .A(n17386), .B(n16857), .Z(n16858) );
  NOR U17157 ( .A(n16859), .B(n16858), .Z(n17392) );
  XOR U17158 ( .A(n16861), .B(n16860), .Z(n17391) );
  NOR U17159 ( .A(n17392), .B(n17391), .Z(n16862) );
  NOR U17160 ( .A(n16863), .B(n16862), .Z(n16868) );
  NOR U17161 ( .A(n156), .B(n57), .Z(n16867) );
  IV U17162 ( .A(n16867), .Z(n16864) );
  NOR U17163 ( .A(n16868), .B(n16864), .Z(n16871) );
  XOR U17164 ( .A(n16866), .B(n16865), .Z(n17399) );
  IV U17165 ( .A(n17399), .Z(n16869) );
  XOR U17166 ( .A(n16868), .B(n16867), .Z(n17398) );
  NOR U17167 ( .A(n16869), .B(n17398), .Z(n16870) );
  NOR U17168 ( .A(n16871), .B(n16870), .Z(n16876) );
  XOR U17169 ( .A(n16873), .B(n16872), .Z(n16875) );
  IV U17170 ( .A(n16875), .Z(n16874) );
  NOR U17171 ( .A(n16876), .B(n16874), .Z(n16879) );
  XOR U17172 ( .A(n16876), .B(n16875), .Z(n16931) );
  NOR U17173 ( .A(n158), .B(n57), .Z(n16932) );
  IV U17174 ( .A(n16932), .Z(n16877) );
  NOR U17175 ( .A(n16931), .B(n16877), .Z(n16878) );
  NOR U17176 ( .A(n16879), .B(n16878), .Z(n16882) );
  NOR U17177 ( .A(n161), .B(n57), .Z(n16881) );
  IV U17178 ( .A(n16881), .Z(n16880) );
  NOR U17179 ( .A(n16882), .B(n16880), .Z(n16886) );
  XOR U17180 ( .A(n16882), .B(n16881), .Z(n17413) );
  XOR U17181 ( .A(n16884), .B(n16883), .Z(n17414) );
  NOR U17182 ( .A(n17413), .B(n17414), .Z(n16885) );
  NOR U17183 ( .A(n16886), .B(n16885), .Z(n16893) );
  NOR U17184 ( .A(n163), .B(n57), .Z(n16892) );
  IV U17185 ( .A(n16892), .Z(n16887) );
  NOR U17186 ( .A(n16893), .B(n16887), .Z(n16895) );
  XOR U17187 ( .A(n16889), .B(n16888), .Z(n16890) );
  XOR U17188 ( .A(n16891), .B(n16890), .Z(n17419) );
  XOR U17189 ( .A(n16893), .B(n16892), .Z(n17418) );
  NOR U17190 ( .A(n17419), .B(n17418), .Z(n16894) );
  NOR U17191 ( .A(n16895), .B(n16894), .Z(n16900) );
  XOR U17192 ( .A(n16897), .B(n16896), .Z(n16899) );
  IV U17193 ( .A(n16899), .Z(n16898) );
  NOR U17194 ( .A(n16900), .B(n16898), .Z(n16903) );
  XOR U17195 ( .A(n16900), .B(n16899), .Z(n17429) );
  NOR U17196 ( .A(n165), .B(n57), .Z(n17430) );
  IV U17197 ( .A(n17430), .Z(n16901) );
  NOR U17198 ( .A(n17429), .B(n16901), .Z(n16902) );
  NOR U17199 ( .A(n16903), .B(n16902), .Z(n17434) );
  XOR U17200 ( .A(n16905), .B(n16904), .Z(n17435) );
  NOR U17201 ( .A(n17434), .B(n17435), .Z(n16906) );
  NOR U17202 ( .A(n16907), .B(n16906), .Z(n28566) );
  XOR U17203 ( .A(n16909), .B(n16908), .Z(n16921) );
  NOR U17204 ( .A(n16911), .B(n16910), .Z(n16916) );
  IV U17205 ( .A(n16912), .Z(n16913) );
  NOR U17206 ( .A(n16914), .B(n16913), .Z(n16915) );
  NOR U17207 ( .A(n16916), .B(n16915), .Z(n16920) );
  NOR U17208 ( .A(n167), .B(n56), .Z(n16918) );
  XOR U17209 ( .A(n16920), .B(n16918), .Z(n16922) );
  XOR U17210 ( .A(n16921), .B(n16922), .Z(n28575) );
  IV U17211 ( .A(n28575), .Z(n16917) );
  NOR U17212 ( .A(n28566), .B(n16917), .Z(n31610) );
  IV U17213 ( .A(n16918), .Z(n16919) );
  NOR U17214 ( .A(n16920), .B(n16919), .Z(n16924) );
  NOR U17215 ( .A(n16922), .B(n16921), .Z(n16923) );
  NOR U17216 ( .A(n16924), .B(n16923), .Z(n16928) );
  XOR U17217 ( .A(n16926), .B(n16925), .Z(n16930) );
  IV U17218 ( .A(n16930), .Z(n16927) );
  NOR U17219 ( .A(n16928), .B(n16927), .Z(n31611) );
  IV U17220 ( .A(n16928), .Z(n16929) );
  NOR U17221 ( .A(n16930), .B(n16929), .Z(n31606) );
  NOR U17222 ( .A(n31611), .B(n31606), .Z(n31602) );
  NOR U17223 ( .A(n31610), .B(n31602), .Z(n17944) );
  XOR U17224 ( .A(n16932), .B(n16931), .Z(n17406) );
  NOR U17225 ( .A(n161), .B(n58), .Z(n17407) );
  IV U17226 ( .A(n17407), .Z(n16933) );
  NOR U17227 ( .A(n17406), .B(n16933), .Z(n17409) );
  XOR U17228 ( .A(n16935), .B(n16934), .Z(n17363) );
  NOR U17229 ( .A(n148), .B(n58), .Z(n17364) );
  IV U17230 ( .A(n17364), .Z(n16936) );
  NOR U17231 ( .A(n17363), .B(n16936), .Z(n17366) );
  XOR U17232 ( .A(n16938), .B(n16937), .Z(n17857) );
  IV U17233 ( .A(n17857), .Z(n16940) );
  NOR U17234 ( .A(n143), .B(n58), .Z(n17855) );
  IV U17235 ( .A(n17855), .Z(n16939) );
  NOR U17236 ( .A(n16940), .B(n16939), .Z(n17346) );
  NOR U17237 ( .A(n17857), .B(n17855), .Z(n17344) );
  XOR U17238 ( .A(n16942), .B(n16941), .Z(n17341) );
  NOR U17239 ( .A(n141), .B(n58), .Z(n17340) );
  IV U17240 ( .A(n17340), .Z(n16943) );
  NOR U17241 ( .A(n17341), .B(n16943), .Z(n17343) );
  NOR U17242 ( .A(n135), .B(n58), .Z(n17311) );
  XOR U17243 ( .A(n16945), .B(n16944), .Z(n17306) );
  NOR U17244 ( .A(n131), .B(n58), .Z(n17302) );
  NOR U17245 ( .A(n128), .B(n58), .Z(n17290) );
  NOR U17246 ( .A(n125), .B(n58), .Z(n17279) );
  IV U17247 ( .A(n17279), .Z(n16948) );
  XOR U17248 ( .A(n16947), .B(n16946), .Z(n17278) );
  NOR U17249 ( .A(n16948), .B(n17278), .Z(n17281) );
  NOR U17250 ( .A(n120), .B(n58), .Z(n17265) );
  IV U17251 ( .A(n17265), .Z(n17770) );
  XOR U17252 ( .A(n16950), .B(n16949), .Z(n17264) );
  IV U17253 ( .A(n17264), .Z(n17769) );
  NOR U17254 ( .A(n17770), .B(n17769), .Z(n17268) );
  NOR U17255 ( .A(n79), .B(n58), .Z(n16953) );
  XOR U17256 ( .A(n16952), .B(n16951), .Z(n16954) );
  NOR U17257 ( .A(n16953), .B(n16954), .Z(n17253) );
  IV U17258 ( .A(n16953), .Z(n17757) );
  IV U17259 ( .A(n16954), .Z(n17756) );
  NOR U17260 ( .A(n17757), .B(n17756), .Z(n17251) );
  XOR U17261 ( .A(n16956), .B(n16955), .Z(n17237) );
  IV U17262 ( .A(n17237), .Z(n17743) );
  NOR U17263 ( .A(n80), .B(n58), .Z(n17236) );
  IV U17264 ( .A(n17236), .Z(n17742) );
  NOR U17265 ( .A(n17743), .B(n17742), .Z(n17240) );
  XOR U17266 ( .A(n16958), .B(n16957), .Z(n16959) );
  NOR U17267 ( .A(n81), .B(n58), .Z(n16960) );
  NOR U17268 ( .A(n16959), .B(n16960), .Z(n17225) );
  IV U17269 ( .A(n16959), .Z(n17729) );
  IV U17270 ( .A(n16960), .Z(n17728) );
  NOR U17271 ( .A(n17729), .B(n17728), .Z(n17223) );
  XOR U17272 ( .A(n16962), .B(n16961), .Z(n16963) );
  NOR U17273 ( .A(n82), .B(n58), .Z(n16964) );
  NOR U17274 ( .A(n16963), .B(n16964), .Z(n17211) );
  IV U17275 ( .A(n16963), .Z(n17464) );
  IV U17276 ( .A(n16964), .Z(n17463) );
  NOR U17277 ( .A(n17464), .B(n17463), .Z(n17209) );
  XOR U17278 ( .A(n16966), .B(n16965), .Z(n16967) );
  XOR U17279 ( .A(n16968), .B(n16967), .Z(n17204) );
  NOR U17280 ( .A(n114), .B(n58), .Z(n17203) );
  IV U17281 ( .A(n17203), .Z(n16969) );
  NOR U17282 ( .A(n17204), .B(n16969), .Z(n17207) );
  NOR U17283 ( .A(n83), .B(n58), .Z(n17199) );
  XOR U17284 ( .A(n16971), .B(n16970), .Z(n17198) );
  NOR U17285 ( .A(n17199), .B(n17198), .Z(n17202) );
  NOR U17286 ( .A(n84), .B(n58), .Z(n16974) );
  XOR U17287 ( .A(n16973), .B(n16972), .Z(n16975) );
  NOR U17288 ( .A(n16974), .B(n16975), .Z(n17187) );
  IV U17289 ( .A(n16974), .Z(n17474) );
  IV U17290 ( .A(n16975), .Z(n17473) );
  NOR U17291 ( .A(n17474), .B(n17473), .Z(n17185) );
  XOR U17292 ( .A(n16977), .B(n16976), .Z(n16978) );
  XOR U17293 ( .A(n16979), .B(n16978), .Z(n17181) );
  NOR U17294 ( .A(n112), .B(n58), .Z(n17180) );
  IV U17295 ( .A(n17180), .Z(n16980) );
  NOR U17296 ( .A(n17181), .B(n16980), .Z(n17183) );
  NOR U17297 ( .A(n85), .B(n58), .Z(n17175) );
  XOR U17298 ( .A(n16982), .B(n16981), .Z(n17174) );
  NOR U17299 ( .A(n17175), .B(n17174), .Z(n17178) );
  XOR U17300 ( .A(n16984), .B(n16983), .Z(n17170) );
  NOR U17301 ( .A(n111), .B(n58), .Z(n17169) );
  IV U17302 ( .A(n17169), .Z(n16985) );
  NOR U17303 ( .A(n17170), .B(n16985), .Z(n17172) );
  IV U17304 ( .A(n16986), .Z(n16988) );
  XOR U17305 ( .A(n16988), .B(n16987), .Z(n17165) );
  NOR U17306 ( .A(n86), .B(n58), .Z(n17166) );
  IV U17307 ( .A(n17166), .Z(n16989) );
  NOR U17308 ( .A(n17165), .B(n16989), .Z(n17168) );
  IV U17309 ( .A(n16990), .Z(n16992) );
  XOR U17310 ( .A(n16992), .B(n16991), .Z(n17161) );
  NOR U17311 ( .A(n110), .B(n58), .Z(n17162) );
  IV U17312 ( .A(n17162), .Z(n16993) );
  NOR U17313 ( .A(n17161), .B(n16993), .Z(n17164) );
  XOR U17314 ( .A(n16995), .B(n16994), .Z(n17157) );
  NOR U17315 ( .A(n109), .B(n58), .Z(n17158) );
  IV U17316 ( .A(n17158), .Z(n16996) );
  NOR U17317 ( .A(n17157), .B(n16996), .Z(n17160) );
  IV U17318 ( .A(n16997), .Z(n16999) );
  XOR U17319 ( .A(n16999), .B(n16998), .Z(n17153) );
  NOR U17320 ( .A(n108), .B(n58), .Z(n17154) );
  IV U17321 ( .A(n17154), .Z(n17000) );
  NOR U17322 ( .A(n17153), .B(n17000), .Z(n17156) );
  XOR U17323 ( .A(n17002), .B(n17001), .Z(n17149) );
  NOR U17324 ( .A(n87), .B(n58), .Z(n17150) );
  IV U17325 ( .A(n17150), .Z(n17003) );
  NOR U17326 ( .A(n17149), .B(n17003), .Z(n17152) );
  IV U17327 ( .A(n17004), .Z(n17006) );
  XOR U17328 ( .A(n17006), .B(n17005), .Z(n17145) );
  NOR U17329 ( .A(n107), .B(n58), .Z(n17146) );
  IV U17330 ( .A(n17146), .Z(n17007) );
  NOR U17331 ( .A(n17145), .B(n17007), .Z(n17148) );
  XOR U17332 ( .A(n17009), .B(n17008), .Z(n17141) );
  NOR U17333 ( .A(n88), .B(n58), .Z(n17142) );
  IV U17334 ( .A(n17142), .Z(n17010) );
  NOR U17335 ( .A(n17141), .B(n17010), .Z(n17144) );
  IV U17336 ( .A(n17011), .Z(n17013) );
  XOR U17337 ( .A(n17013), .B(n17012), .Z(n17137) );
  NOR U17338 ( .A(n106), .B(n58), .Z(n17138) );
  IV U17339 ( .A(n17138), .Z(n17014) );
  NOR U17340 ( .A(n17137), .B(n17014), .Z(n17140) );
  XOR U17341 ( .A(n17016), .B(n17015), .Z(n17133) );
  IV U17342 ( .A(n17133), .Z(n17018) );
  NOR U17343 ( .A(n105), .B(n58), .Z(n17017) );
  IV U17344 ( .A(n17017), .Z(n17134) );
  NOR U17345 ( .A(n17018), .B(n17134), .Z(n17136) );
  IV U17346 ( .A(n17019), .Z(n17021) );
  XOR U17347 ( .A(n17021), .B(n17020), .Z(n17121) );
  NOR U17348 ( .A(n89), .B(n58), .Z(n17122) );
  IV U17349 ( .A(n17122), .Z(n17022) );
  NOR U17350 ( .A(n17121), .B(n17022), .Z(n17124) );
  IV U17351 ( .A(n17023), .Z(n17025) );
  XOR U17352 ( .A(n17025), .B(n17024), .Z(n17117) );
  NOR U17353 ( .A(n103), .B(n58), .Z(n17118) );
  IV U17354 ( .A(n17118), .Z(n17026) );
  NOR U17355 ( .A(n17117), .B(n17026), .Z(n17120) );
  IV U17356 ( .A(n17027), .Z(n17029) );
  XOR U17357 ( .A(n17029), .B(n17028), .Z(n17113) );
  NOR U17358 ( .A(n90), .B(n58), .Z(n17114) );
  IV U17359 ( .A(n17114), .Z(n17030) );
  NOR U17360 ( .A(n17113), .B(n17030), .Z(n17116) );
  IV U17361 ( .A(n17031), .Z(n17033) );
  XOR U17362 ( .A(n17033), .B(n17032), .Z(n17109) );
  NOR U17363 ( .A(n102), .B(n58), .Z(n17110) );
  IV U17364 ( .A(n17110), .Z(n17034) );
  NOR U17365 ( .A(n17109), .B(n17034), .Z(n17112) );
  IV U17366 ( .A(n17035), .Z(n17037) );
  XOR U17367 ( .A(n17037), .B(n17036), .Z(n17105) );
  NOR U17368 ( .A(n101), .B(n58), .Z(n17106) );
  IV U17369 ( .A(n17106), .Z(n17038) );
  NOR U17370 ( .A(n17105), .B(n17038), .Z(n17108) );
  IV U17371 ( .A(n17039), .Z(n17041) );
  XOR U17372 ( .A(n17041), .B(n17040), .Z(n17101) );
  NOR U17373 ( .A(n100), .B(n58), .Z(n17102) );
  IV U17374 ( .A(n17102), .Z(n17042) );
  NOR U17375 ( .A(n17101), .B(n17042), .Z(n17104) );
  IV U17376 ( .A(n17043), .Z(n17045) );
  XOR U17377 ( .A(n17045), .B(n17044), .Z(n17097) );
  NOR U17378 ( .A(n99), .B(n58), .Z(n17098) );
  IV U17379 ( .A(n17098), .Z(n17046) );
  NOR U17380 ( .A(n17097), .B(n17046), .Z(n17100) );
  IV U17381 ( .A(n17047), .Z(n17049) );
  XOR U17382 ( .A(n17049), .B(n17048), .Z(n17093) );
  NOR U17383 ( .A(n98), .B(n58), .Z(n17094) );
  IV U17384 ( .A(n17094), .Z(n17050) );
  NOR U17385 ( .A(n17093), .B(n17050), .Z(n17096) );
  XOR U17386 ( .A(n17052), .B(n17051), .Z(n17089) );
  NOR U17387 ( .A(n91), .B(n58), .Z(n17090) );
  IV U17388 ( .A(n17090), .Z(n17053) );
  NOR U17389 ( .A(n17089), .B(n17053), .Z(n17092) );
  XOR U17390 ( .A(n17055), .B(n17054), .Z(n17077) );
  IV U17391 ( .A(n17077), .Z(n17057) );
  NOR U17392 ( .A(n96), .B(n58), .Z(n17056) );
  IV U17393 ( .A(n17056), .Z(n17078) );
  NOR U17394 ( .A(n17057), .B(n17078), .Z(n17080) );
  NOR U17395 ( .A(n95), .B(n58), .Z(n17074) );
  IV U17396 ( .A(n17074), .Z(n17060) );
  XOR U17397 ( .A(n17059), .B(n17058), .Z(n17073) );
  NOR U17398 ( .A(n17060), .B(n17073), .Z(n17076) );
  NOR U17399 ( .A(n58), .B(n93), .Z(n18079) );
  IV U17400 ( .A(n18079), .Z(n17061) );
  NOR U17401 ( .A(n57), .B(n168), .Z(n17069) );
  IV U17402 ( .A(n17069), .Z(n17064) );
  NOR U17403 ( .A(n17061), .B(n17064), .Z(n17062) );
  IV U17404 ( .A(n17062), .Z(n17063) );
  NOR U17405 ( .A(n94), .B(n17063), .Z(n17072) );
  NOR U17406 ( .A(n17064), .B(n93), .Z(n17065) );
  XOR U17407 ( .A(n94), .B(n17065), .Z(n17066) );
  NOR U17408 ( .A(n58), .B(n17066), .Z(n17067) );
  IV U17409 ( .A(n17067), .Z(n17562) );
  XOR U17410 ( .A(n17069), .B(n17068), .Z(n17561) );
  IV U17411 ( .A(n17561), .Z(n17070) );
  NOR U17412 ( .A(n17562), .B(n17070), .Z(n17071) );
  NOR U17413 ( .A(n17072), .B(n17071), .Z(n17558) );
  XOR U17414 ( .A(n17074), .B(n17073), .Z(n17557) );
  NOR U17415 ( .A(n17558), .B(n17557), .Z(n17075) );
  NOR U17416 ( .A(n17076), .B(n17075), .Z(n17585) );
  XOR U17417 ( .A(n17078), .B(n17077), .Z(n17584) );
  NOR U17418 ( .A(n17585), .B(n17584), .Z(n17079) );
  NOR U17419 ( .A(n17080), .B(n17079), .Z(n17085) );
  XOR U17420 ( .A(n17082), .B(n17081), .Z(n17084) );
  IV U17421 ( .A(n17084), .Z(n17083) );
  NOR U17422 ( .A(n17085), .B(n17083), .Z(n17088) );
  XOR U17423 ( .A(n17085), .B(n17084), .Z(n17554) );
  NOR U17424 ( .A(n97), .B(n58), .Z(n17555) );
  IV U17425 ( .A(n17555), .Z(n17086) );
  NOR U17426 ( .A(n17554), .B(n17086), .Z(n17087) );
  NOR U17427 ( .A(n17088), .B(n17087), .Z(n17550) );
  XOR U17428 ( .A(n17090), .B(n17089), .Z(n17551) );
  NOR U17429 ( .A(n17550), .B(n17551), .Z(n17091) );
  NOR U17430 ( .A(n17092), .B(n17091), .Z(n17546) );
  XOR U17431 ( .A(n17094), .B(n17093), .Z(n17547) );
  NOR U17432 ( .A(n17546), .B(n17547), .Z(n17095) );
  NOR U17433 ( .A(n17096), .B(n17095), .Z(n17542) );
  XOR U17434 ( .A(n17098), .B(n17097), .Z(n17543) );
  NOR U17435 ( .A(n17542), .B(n17543), .Z(n17099) );
  NOR U17436 ( .A(n17100), .B(n17099), .Z(n17538) );
  XOR U17437 ( .A(n17102), .B(n17101), .Z(n17539) );
  NOR U17438 ( .A(n17538), .B(n17539), .Z(n17103) );
  NOR U17439 ( .A(n17104), .B(n17103), .Z(n17534) );
  XOR U17440 ( .A(n17106), .B(n17105), .Z(n17535) );
  NOR U17441 ( .A(n17534), .B(n17535), .Z(n17107) );
  NOR U17442 ( .A(n17108), .B(n17107), .Z(n17530) );
  XOR U17443 ( .A(n17110), .B(n17109), .Z(n17531) );
  NOR U17444 ( .A(n17530), .B(n17531), .Z(n17111) );
  NOR U17445 ( .A(n17112), .B(n17111), .Z(n17526) );
  XOR U17446 ( .A(n17114), .B(n17113), .Z(n17527) );
  NOR U17447 ( .A(n17526), .B(n17527), .Z(n17115) );
  NOR U17448 ( .A(n17116), .B(n17115), .Z(n17523) );
  XOR U17449 ( .A(n17118), .B(n17117), .Z(n17522) );
  NOR U17450 ( .A(n17523), .B(n17522), .Z(n17119) );
  NOR U17451 ( .A(n17120), .B(n17119), .Z(n17518) );
  XOR U17452 ( .A(n17122), .B(n17121), .Z(n17519) );
  NOR U17453 ( .A(n17518), .B(n17519), .Z(n17123) );
  NOR U17454 ( .A(n17124), .B(n17123), .Z(n17129) );
  XOR U17455 ( .A(n17126), .B(n17125), .Z(n17128) );
  IV U17456 ( .A(n17128), .Z(n17127) );
  NOR U17457 ( .A(n17129), .B(n17127), .Z(n17132) );
  XOR U17458 ( .A(n17129), .B(n17128), .Z(n17515) );
  NOR U17459 ( .A(n104), .B(n58), .Z(n17516) );
  IV U17460 ( .A(n17516), .Z(n17130) );
  NOR U17461 ( .A(n17515), .B(n17130), .Z(n17131) );
  NOR U17462 ( .A(n17132), .B(n17131), .Z(n17637) );
  XOR U17463 ( .A(n17134), .B(n17133), .Z(n17636) );
  NOR U17464 ( .A(n17637), .B(n17636), .Z(n17135) );
  NOR U17465 ( .A(n17136), .B(n17135), .Z(n17512) );
  XOR U17466 ( .A(n17138), .B(n17137), .Z(n17511) );
  NOR U17467 ( .A(n17512), .B(n17511), .Z(n17139) );
  NOR U17468 ( .A(n17140), .B(n17139), .Z(n17507) );
  XOR U17469 ( .A(n17142), .B(n17141), .Z(n17508) );
  NOR U17470 ( .A(n17507), .B(n17508), .Z(n17143) );
  NOR U17471 ( .A(n17144), .B(n17143), .Z(n17504) );
  XOR U17472 ( .A(n17146), .B(n17145), .Z(n17503) );
  NOR U17473 ( .A(n17504), .B(n17503), .Z(n17147) );
  NOR U17474 ( .A(n17148), .B(n17147), .Z(n17499) );
  XOR U17475 ( .A(n17150), .B(n17149), .Z(n17500) );
  NOR U17476 ( .A(n17499), .B(n17500), .Z(n17151) );
  NOR U17477 ( .A(n17152), .B(n17151), .Z(n17495) );
  XOR U17478 ( .A(n17154), .B(n17153), .Z(n17496) );
  NOR U17479 ( .A(n17495), .B(n17496), .Z(n17155) );
  NOR U17480 ( .A(n17156), .B(n17155), .Z(n17491) );
  XOR U17481 ( .A(n17158), .B(n17157), .Z(n17492) );
  NOR U17482 ( .A(n17491), .B(n17492), .Z(n17159) );
  NOR U17483 ( .A(n17160), .B(n17159), .Z(n17490) );
  XOR U17484 ( .A(n17162), .B(n17161), .Z(n17489) );
  NOR U17485 ( .A(n17490), .B(n17489), .Z(n17163) );
  NOR U17486 ( .A(n17164), .B(n17163), .Z(n17486) );
  XOR U17487 ( .A(n17166), .B(n17165), .Z(n17485) );
  NOR U17488 ( .A(n17486), .B(n17485), .Z(n17167) );
  NOR U17489 ( .A(n17168), .B(n17167), .Z(n17484) );
  XOR U17490 ( .A(n17170), .B(n17169), .Z(n17483) );
  NOR U17491 ( .A(n17484), .B(n17483), .Z(n17171) );
  NOR U17492 ( .A(n17172), .B(n17171), .Z(n17173) );
  IV U17493 ( .A(n17173), .Z(n17481) );
  XOR U17494 ( .A(n17175), .B(n17174), .Z(n17176) );
  IV U17495 ( .A(n17176), .Z(n17480) );
  NOR U17496 ( .A(n17481), .B(n17480), .Z(n17177) );
  NOR U17497 ( .A(n17178), .B(n17177), .Z(n17179) );
  IV U17498 ( .A(n17179), .Z(n17479) );
  XOR U17499 ( .A(n17181), .B(n17180), .Z(n17478) );
  NOR U17500 ( .A(n17479), .B(n17478), .Z(n17182) );
  NOR U17501 ( .A(n17183), .B(n17182), .Z(n17476) );
  IV U17502 ( .A(n17476), .Z(n17184) );
  NOR U17503 ( .A(n17185), .B(n17184), .Z(n17186) );
  NOR U17504 ( .A(n17187), .B(n17186), .Z(n17194) );
  IV U17505 ( .A(n17194), .Z(n17189) );
  NOR U17506 ( .A(n113), .B(n58), .Z(n17188) );
  IV U17507 ( .A(n17188), .Z(n17193) );
  NOR U17508 ( .A(n17189), .B(n17193), .Z(n17196) );
  XOR U17509 ( .A(n17191), .B(n17190), .Z(n17192) );
  IV U17510 ( .A(n17192), .Z(n17471) );
  XOR U17511 ( .A(n17194), .B(n17193), .Z(n17472) );
  NOR U17512 ( .A(n17471), .B(n17472), .Z(n17195) );
  NOR U17513 ( .A(n17196), .B(n17195), .Z(n17197) );
  IV U17514 ( .A(n17197), .Z(n17708) );
  XOR U17515 ( .A(n17199), .B(n17198), .Z(n17200) );
  IV U17516 ( .A(n17200), .Z(n17707) );
  NOR U17517 ( .A(n17708), .B(n17707), .Z(n17201) );
  NOR U17518 ( .A(n17202), .B(n17201), .Z(n17469) );
  IV U17519 ( .A(n17469), .Z(n17205) );
  XOR U17520 ( .A(n17204), .B(n17203), .Z(n17468) );
  NOR U17521 ( .A(n17205), .B(n17468), .Z(n17206) );
  NOR U17522 ( .A(n17207), .B(n17206), .Z(n17466) );
  IV U17523 ( .A(n17466), .Z(n17208) );
  NOR U17524 ( .A(n17209), .B(n17208), .Z(n17210) );
  NOR U17525 ( .A(n17211), .B(n17210), .Z(n17219) );
  IV U17526 ( .A(n17219), .Z(n17213) );
  NOR U17527 ( .A(n115), .B(n58), .Z(n17212) );
  IV U17528 ( .A(n17212), .Z(n17218) );
  NOR U17529 ( .A(n17213), .B(n17218), .Z(n17221) );
  XOR U17530 ( .A(n17215), .B(n17214), .Z(n17216) );
  XOR U17531 ( .A(n17217), .B(n17216), .Z(n17462) );
  XOR U17532 ( .A(n17219), .B(n17218), .Z(n17461) );
  NOR U17533 ( .A(n17462), .B(n17461), .Z(n17220) );
  NOR U17534 ( .A(n17221), .B(n17220), .Z(n17731) );
  IV U17535 ( .A(n17731), .Z(n17222) );
  NOR U17536 ( .A(n17223), .B(n17222), .Z(n17224) );
  NOR U17537 ( .A(n17225), .B(n17224), .Z(n17226) );
  IV U17538 ( .A(n17226), .Z(n17233) );
  NOR U17539 ( .A(n116), .B(n58), .Z(n17232) );
  IV U17540 ( .A(n17232), .Z(n17227) );
  NOR U17541 ( .A(n17233), .B(n17227), .Z(n17235) );
  XOR U17542 ( .A(n17229), .B(n17228), .Z(n17230) );
  XOR U17543 ( .A(n17231), .B(n17230), .Z(n17457) );
  XOR U17544 ( .A(n17233), .B(n17232), .Z(n17458) );
  NOR U17545 ( .A(n17457), .B(n17458), .Z(n17234) );
  NOR U17546 ( .A(n17235), .B(n17234), .Z(n17745) );
  NOR U17547 ( .A(n17237), .B(n17236), .Z(n17238) );
  NOR U17548 ( .A(n17745), .B(n17238), .Z(n17239) );
  NOR U17549 ( .A(n17240), .B(n17239), .Z(n17246) );
  NOR U17550 ( .A(n117), .B(n58), .Z(n17247) );
  IV U17551 ( .A(n17247), .Z(n17241) );
  NOR U17552 ( .A(n17246), .B(n17241), .Z(n17249) );
  XOR U17553 ( .A(n17243), .B(n17242), .Z(n17244) );
  XOR U17554 ( .A(n17245), .B(n17244), .Z(n17454) );
  XOR U17555 ( .A(n17247), .B(n17246), .Z(n17453) );
  NOR U17556 ( .A(n17454), .B(n17453), .Z(n17248) );
  NOR U17557 ( .A(n17249), .B(n17248), .Z(n17759) );
  IV U17558 ( .A(n17759), .Z(n17250) );
  NOR U17559 ( .A(n17251), .B(n17250), .Z(n17252) );
  NOR U17560 ( .A(n17253), .B(n17252), .Z(n17254) );
  IV U17561 ( .A(n17254), .Z(n17261) );
  NOR U17562 ( .A(n119), .B(n58), .Z(n17260) );
  IV U17563 ( .A(n17260), .Z(n17255) );
  NOR U17564 ( .A(n17261), .B(n17255), .Z(n17263) );
  XOR U17565 ( .A(n17257), .B(n17256), .Z(n17258) );
  XOR U17566 ( .A(n17259), .B(n17258), .Z(n17449) );
  XOR U17567 ( .A(n17261), .B(n17260), .Z(n17450) );
  NOR U17568 ( .A(n17449), .B(n17450), .Z(n17262) );
  NOR U17569 ( .A(n17263), .B(n17262), .Z(n17772) );
  NOR U17570 ( .A(n17265), .B(n17264), .Z(n17266) );
  NOR U17571 ( .A(n17772), .B(n17266), .Z(n17267) );
  NOR U17572 ( .A(n17268), .B(n17267), .Z(n17275) );
  NOR U17573 ( .A(n123), .B(n58), .Z(n17274) );
  IV U17574 ( .A(n17274), .Z(n17269) );
  NOR U17575 ( .A(n17275), .B(n17269), .Z(n17277) );
  XOR U17576 ( .A(n17271), .B(n17270), .Z(n17272) );
  XOR U17577 ( .A(n17273), .B(n17272), .Z(n17447) );
  XOR U17578 ( .A(n17275), .B(n17274), .Z(n17446) );
  NOR U17579 ( .A(n17447), .B(n17446), .Z(n17276) );
  NOR U17580 ( .A(n17277), .B(n17276), .Z(n17783) );
  XOR U17581 ( .A(n17279), .B(n17278), .Z(n17784) );
  NOR U17582 ( .A(n17783), .B(n17784), .Z(n17280) );
  NOR U17583 ( .A(n17281), .B(n17280), .Z(n17286) );
  XOR U17584 ( .A(n17283), .B(n17282), .Z(n17285) );
  IV U17585 ( .A(n17285), .Z(n17284) );
  NOR U17586 ( .A(n17286), .B(n17284), .Z(n17289) );
  XOR U17587 ( .A(n17286), .B(n17285), .Z(n17791) );
  NOR U17588 ( .A(n126), .B(n58), .Z(n17792) );
  IV U17589 ( .A(n17792), .Z(n17287) );
  NOR U17590 ( .A(n17791), .B(n17287), .Z(n17288) );
  NOR U17591 ( .A(n17289), .B(n17288), .Z(n17291) );
  IV U17592 ( .A(n17291), .Z(n17798) );
  NOR U17593 ( .A(n17290), .B(n17798), .Z(n17296) );
  IV U17594 ( .A(n17290), .Z(n17799) );
  NOR U17595 ( .A(n17291), .B(n17799), .Z(n17294) );
  XOR U17596 ( .A(n17293), .B(n17292), .Z(n17801) );
  NOR U17597 ( .A(n17294), .B(n17801), .Z(n17295) );
  NOR U17598 ( .A(n17296), .B(n17295), .Z(n17301) );
  NOR U17599 ( .A(n17302), .B(n17301), .Z(n17305) );
  XOR U17600 ( .A(n17298), .B(n17297), .Z(n17299) );
  XOR U17601 ( .A(n17300), .B(n17299), .Z(n17807) );
  XOR U17602 ( .A(n17302), .B(n17301), .Z(n17806) );
  IV U17603 ( .A(n17806), .Z(n17303) );
  NOR U17604 ( .A(n17807), .B(n17303), .Z(n17304) );
  NOR U17605 ( .A(n17305), .B(n17304), .Z(n17307) );
  NOR U17606 ( .A(n17306), .B(n17307), .Z(n17310) );
  IV U17607 ( .A(n17306), .Z(n17817) );
  IV U17608 ( .A(n17307), .Z(n17816) );
  NOR U17609 ( .A(n17817), .B(n17816), .Z(n17308) );
  NOR U17610 ( .A(n133), .B(n58), .Z(n17819) );
  NOR U17611 ( .A(n17308), .B(n17819), .Z(n17309) );
  NOR U17612 ( .A(n17310), .B(n17309), .Z(n17312) );
  NOR U17613 ( .A(n17311), .B(n17312), .Z(n17320) );
  IV U17614 ( .A(n17311), .Z(n17826) );
  IV U17615 ( .A(n17312), .Z(n17825) );
  NOR U17616 ( .A(n17826), .B(n17825), .Z(n17318) );
  XOR U17617 ( .A(n17314), .B(n17313), .Z(n17315) );
  XOR U17618 ( .A(n17316), .B(n17315), .Z(n17828) );
  IV U17619 ( .A(n17828), .Z(n17317) );
  NOR U17620 ( .A(n17318), .B(n17317), .Z(n17319) );
  NOR U17621 ( .A(n17320), .B(n17319), .Z(n17328) );
  IV U17622 ( .A(n17328), .Z(n17322) );
  NOR U17623 ( .A(n137), .B(n58), .Z(n17321) );
  IV U17624 ( .A(n17321), .Z(n17327) );
  NOR U17625 ( .A(n17322), .B(n17327), .Z(n17331) );
  XOR U17626 ( .A(n17324), .B(n17323), .Z(n17325) );
  XOR U17627 ( .A(n17326), .B(n17325), .Z(n17834) );
  IV U17628 ( .A(n17834), .Z(n17329) );
  XOR U17629 ( .A(n17328), .B(n17327), .Z(n17833) );
  NOR U17630 ( .A(n17329), .B(n17833), .Z(n17330) );
  NOR U17631 ( .A(n17331), .B(n17330), .Z(n17336) );
  XOR U17632 ( .A(n17333), .B(n17332), .Z(n17335) );
  IV U17633 ( .A(n17335), .Z(n17334) );
  NOR U17634 ( .A(n17336), .B(n17334), .Z(n17339) );
  XOR U17635 ( .A(n17336), .B(n17335), .Z(n17444) );
  NOR U17636 ( .A(n139), .B(n58), .Z(n17443) );
  IV U17637 ( .A(n17443), .Z(n17337) );
  NOR U17638 ( .A(n17444), .B(n17337), .Z(n17338) );
  NOR U17639 ( .A(n17339), .B(n17338), .Z(n17846) );
  XOR U17640 ( .A(n17341), .B(n17340), .Z(n17845) );
  NOR U17641 ( .A(n17846), .B(n17845), .Z(n17342) );
  NOR U17642 ( .A(n17343), .B(n17342), .Z(n17854) );
  NOR U17643 ( .A(n17344), .B(n17854), .Z(n17345) );
  NOR U17644 ( .A(n17346), .B(n17345), .Z(n17349) );
  NOR U17645 ( .A(n145), .B(n58), .Z(n17348) );
  IV U17646 ( .A(n17348), .Z(n17347) );
  NOR U17647 ( .A(n17349), .B(n17347), .Z(n17354) );
  XOR U17648 ( .A(n17349), .B(n17348), .Z(n17863) );
  XOR U17649 ( .A(n17351), .B(n17350), .Z(n17862) );
  IV U17650 ( .A(n17862), .Z(n17352) );
  NOR U17651 ( .A(n17863), .B(n17352), .Z(n17353) );
  NOR U17652 ( .A(n17354), .B(n17353), .Z(n17358) );
  XOR U17653 ( .A(n17356), .B(n17355), .Z(n17357) );
  NOR U17654 ( .A(n17358), .B(n17357), .Z(n17362) );
  XOR U17655 ( .A(n17358), .B(n17357), .Z(n17359) );
  IV U17656 ( .A(n17359), .Z(n17874) );
  NOR U17657 ( .A(n147), .B(n58), .Z(n17360) );
  IV U17658 ( .A(n17360), .Z(n17873) );
  NOR U17659 ( .A(n17874), .B(n17873), .Z(n17361) );
  NOR U17660 ( .A(n17362), .B(n17361), .Z(n17882) );
  XOR U17661 ( .A(n17364), .B(n17363), .Z(n17881) );
  NOR U17662 ( .A(n17882), .B(n17881), .Z(n17365) );
  NOR U17663 ( .A(n17366), .B(n17365), .Z(n17369) );
  NOR U17664 ( .A(n150), .B(n58), .Z(n17368) );
  IV U17665 ( .A(n17368), .Z(n17367) );
  NOR U17666 ( .A(n17369), .B(n17367), .Z(n17374) );
  XOR U17667 ( .A(n17369), .B(n17368), .Z(n17887) );
  XOR U17668 ( .A(n17371), .B(n17370), .Z(n17886) );
  IV U17669 ( .A(n17886), .Z(n17372) );
  NOR U17670 ( .A(n17887), .B(n17372), .Z(n17373) );
  NOR U17671 ( .A(n17374), .B(n17373), .Z(n17378) );
  XOR U17672 ( .A(n17376), .B(n17375), .Z(n17377) );
  NOR U17673 ( .A(n17378), .B(n17377), .Z(n17382) );
  XOR U17674 ( .A(n17378), .B(n17377), .Z(n17441) );
  IV U17675 ( .A(n17441), .Z(n17380) );
  NOR U17676 ( .A(n153), .B(n58), .Z(n17379) );
  IV U17677 ( .A(n17379), .Z(n17440) );
  NOR U17678 ( .A(n17380), .B(n17440), .Z(n17381) );
  NOR U17679 ( .A(n17382), .B(n17381), .Z(n17385) );
  NOR U17680 ( .A(n155), .B(n58), .Z(n17384) );
  IV U17681 ( .A(n17384), .Z(n17383) );
  NOR U17682 ( .A(n17385), .B(n17383), .Z(n17389) );
  XOR U17683 ( .A(n17385), .B(n17384), .Z(n17902) );
  XOR U17684 ( .A(n17387), .B(n17386), .Z(n17901) );
  NOR U17685 ( .A(n17902), .B(n17901), .Z(n17388) );
  NOR U17686 ( .A(n17389), .B(n17388), .Z(n17394) );
  NOR U17687 ( .A(n156), .B(n58), .Z(n17393) );
  IV U17688 ( .A(n17393), .Z(n17390) );
  NOR U17689 ( .A(n17394), .B(n17390), .Z(n17397) );
  XOR U17690 ( .A(n17392), .B(n17391), .Z(n17907) );
  IV U17691 ( .A(n17907), .Z(n17395) );
  XOR U17692 ( .A(n17394), .B(n17393), .Z(n17906) );
  NOR U17693 ( .A(n17395), .B(n17906), .Z(n17396) );
  NOR U17694 ( .A(n17397), .B(n17396), .Z(n17401) );
  XOR U17695 ( .A(n17399), .B(n17398), .Z(n17400) );
  NOR U17696 ( .A(n17401), .B(n17400), .Z(n17405) );
  XOR U17697 ( .A(n17401), .B(n17400), .Z(n17918) );
  IV U17698 ( .A(n17918), .Z(n17403) );
  NOR U17699 ( .A(n158), .B(n58), .Z(n17402) );
  IV U17700 ( .A(n17402), .Z(n17917) );
  NOR U17701 ( .A(n17403), .B(n17917), .Z(n17404) );
  NOR U17702 ( .A(n17405), .B(n17404), .Z(n17925) );
  XOR U17703 ( .A(n17407), .B(n17406), .Z(n17924) );
  NOR U17704 ( .A(n17925), .B(n17924), .Z(n17408) );
  NOR U17705 ( .A(n17409), .B(n17408), .Z(n17412) );
  NOR U17706 ( .A(n163), .B(n58), .Z(n17411) );
  IV U17707 ( .A(n17411), .Z(n17410) );
  NOR U17708 ( .A(n17412), .B(n17410), .Z(n17417) );
  XOR U17709 ( .A(n17412), .B(n17411), .Z(n17930) );
  XOR U17710 ( .A(n17414), .B(n17413), .Z(n17929) );
  IV U17711 ( .A(n17929), .Z(n17415) );
  NOR U17712 ( .A(n17930), .B(n17415), .Z(n17416) );
  NOR U17713 ( .A(n17417), .B(n17416), .Z(n17422) );
  XOR U17714 ( .A(n17419), .B(n17418), .Z(n17421) );
  IV U17715 ( .A(n17421), .Z(n17420) );
  NOR U17716 ( .A(n17422), .B(n17420), .Z(n17425) );
  XOR U17717 ( .A(n17422), .B(n17421), .Z(n17438) );
  NOR U17718 ( .A(n165), .B(n58), .Z(n17437) );
  IV U17719 ( .A(n17437), .Z(n17423) );
  NOR U17720 ( .A(n17438), .B(n17423), .Z(n17424) );
  NOR U17721 ( .A(n17425), .B(n17424), .Z(n17428) );
  NOR U17722 ( .A(n167), .B(n58), .Z(n17426) );
  IV U17723 ( .A(n17426), .Z(n17427) );
  NOR U17724 ( .A(n17428), .B(n17427), .Z(n17433) );
  XOR U17725 ( .A(n17428), .B(n17427), .Z(n17942) );
  IV U17726 ( .A(n17942), .Z(n17431) );
  XOR U17727 ( .A(n17430), .B(n17429), .Z(n17941) );
  NOR U17728 ( .A(n17431), .B(n17941), .Z(n17432) );
  NOR U17729 ( .A(n17433), .B(n17432), .Z(n28565) );
  IV U17730 ( .A(n17434), .Z(n17436) );
  XOR U17731 ( .A(n17436), .B(n17435), .Z(n28564) );
  XOR U17732 ( .A(n28565), .B(n28564), .Z(n28570) );
  XOR U17733 ( .A(n17438), .B(n17437), .Z(n17938) );
  NOR U17734 ( .A(n167), .B(n59), .Z(n17937) );
  IV U17735 ( .A(n17937), .Z(n17439) );
  NOR U17736 ( .A(n17938), .B(n17439), .Z(n17940) );
  XOR U17737 ( .A(n17441), .B(n17440), .Z(n17895) );
  NOR U17738 ( .A(n155), .B(n59), .Z(n17894) );
  IV U17739 ( .A(n17894), .Z(n17442) );
  NOR U17740 ( .A(n17895), .B(n17442), .Z(n17897) );
  XOR U17741 ( .A(n17444), .B(n17443), .Z(n17842) );
  NOR U17742 ( .A(n141), .B(n59), .Z(n17841) );
  IV U17743 ( .A(n17841), .Z(n17445) );
  NOR U17744 ( .A(n17842), .B(n17445), .Z(n17844) );
  NOR U17745 ( .A(n135), .B(n59), .Z(n17814) );
  XOR U17746 ( .A(n17447), .B(n17446), .Z(n17778) );
  IV U17747 ( .A(n17778), .Z(n18292) );
  NOR U17748 ( .A(n125), .B(n59), .Z(n17777) );
  IV U17749 ( .A(n17777), .Z(n18291) );
  NOR U17750 ( .A(n18292), .B(n18291), .Z(n17781) );
  NOR U17751 ( .A(n123), .B(n59), .Z(n17448) );
  IV U17752 ( .A(n17448), .Z(n17774) );
  NOR U17753 ( .A(n120), .B(n59), .Z(n17451) );
  XOR U17754 ( .A(n17450), .B(n17449), .Z(n17452) );
  NOR U17755 ( .A(n17451), .B(n17452), .Z(n17767) );
  IV U17756 ( .A(n17451), .Z(n18278) );
  IV U17757 ( .A(n17452), .Z(n18277) );
  NOR U17758 ( .A(n18278), .B(n18277), .Z(n17765) );
  NOR U17759 ( .A(n79), .B(n59), .Z(n17455) );
  XOR U17760 ( .A(n17454), .B(n17453), .Z(n17456) );
  NOR U17761 ( .A(n17455), .B(n17456), .Z(n17753) );
  IV U17762 ( .A(n17455), .Z(n18265) );
  IV U17763 ( .A(n17456), .Z(n18264) );
  NOR U17764 ( .A(n18265), .B(n18264), .Z(n17751) );
  XOR U17765 ( .A(n17458), .B(n17457), .Z(n17459) );
  NOR U17766 ( .A(n80), .B(n59), .Z(n17460) );
  NOR U17767 ( .A(n17459), .B(n17460), .Z(n17739) );
  IV U17768 ( .A(n17459), .Z(n18252) );
  IV U17769 ( .A(n17460), .Z(n18251) );
  NOR U17770 ( .A(n18252), .B(n18251), .Z(n17737) );
  XOR U17771 ( .A(n17462), .B(n17461), .Z(n17723) );
  IV U17772 ( .A(n17723), .Z(n17972) );
  NOR U17773 ( .A(n81), .B(n59), .Z(n17722) );
  IV U17774 ( .A(n17722), .Z(n17971) );
  NOR U17775 ( .A(n17972), .B(n17971), .Z(n17726) );
  XOR U17776 ( .A(n17464), .B(n17463), .Z(n17465) );
  XOR U17777 ( .A(n17466), .B(n17465), .Z(n17719) );
  NOR U17778 ( .A(n115), .B(n59), .Z(n17718) );
  IV U17779 ( .A(n17718), .Z(n17467) );
  NOR U17780 ( .A(n17719), .B(n17467), .Z(n17721) );
  XOR U17781 ( .A(n17469), .B(n17468), .Z(n17713) );
  NOR U17782 ( .A(n82), .B(n59), .Z(n17470) );
  IV U17783 ( .A(n17470), .Z(n17714) );
  NOR U17784 ( .A(n17713), .B(n17714), .Z(n17717) );
  XOR U17785 ( .A(n17472), .B(n17471), .Z(n17702) );
  IV U17786 ( .A(n17702), .Z(n17983) );
  NOR U17787 ( .A(n83), .B(n59), .Z(n17701) );
  IV U17788 ( .A(n17701), .Z(n17982) );
  NOR U17789 ( .A(n17983), .B(n17982), .Z(n17705) );
  XOR U17790 ( .A(n17474), .B(n17473), .Z(n17475) );
  XOR U17791 ( .A(n17476), .B(n17475), .Z(n17698) );
  NOR U17792 ( .A(n113), .B(n59), .Z(n17697) );
  IV U17793 ( .A(n17697), .Z(n17477) );
  NOR U17794 ( .A(n17698), .B(n17477), .Z(n17700) );
  NOR U17795 ( .A(n84), .B(n59), .Z(n17692) );
  XOR U17796 ( .A(n17479), .B(n17478), .Z(n17691) );
  NOR U17797 ( .A(n17692), .B(n17691), .Z(n17695) );
  XOR U17798 ( .A(n17481), .B(n17480), .Z(n17687) );
  NOR U17799 ( .A(n112), .B(n59), .Z(n17686) );
  IV U17800 ( .A(n17686), .Z(n17482) );
  NOR U17801 ( .A(n17687), .B(n17482), .Z(n17689) );
  NOR U17802 ( .A(n85), .B(n59), .Z(n17681) );
  XOR U17803 ( .A(n17484), .B(n17483), .Z(n17680) );
  NOR U17804 ( .A(n17681), .B(n17680), .Z(n17684) );
  XOR U17805 ( .A(n17486), .B(n17485), .Z(n17675) );
  IV U17806 ( .A(n17675), .Z(n17488) );
  NOR U17807 ( .A(n111), .B(n59), .Z(n17487) );
  IV U17808 ( .A(n17487), .Z(n17676) );
  NOR U17809 ( .A(n17488), .B(n17676), .Z(n17678) );
  NOR U17810 ( .A(n86), .B(n59), .Z(n17670) );
  XOR U17811 ( .A(n17490), .B(n17489), .Z(n17669) );
  NOR U17812 ( .A(n17670), .B(n17669), .Z(n17673) );
  IV U17813 ( .A(n17491), .Z(n17493) );
  XOR U17814 ( .A(n17493), .B(n17492), .Z(n17664) );
  NOR U17815 ( .A(n110), .B(n59), .Z(n17665) );
  IV U17816 ( .A(n17665), .Z(n17494) );
  NOR U17817 ( .A(n17664), .B(n17494), .Z(n17667) );
  IV U17818 ( .A(n17495), .Z(n17497) );
  XOR U17819 ( .A(n17497), .B(n17496), .Z(n17660) );
  NOR U17820 ( .A(n109), .B(n59), .Z(n17661) );
  IV U17821 ( .A(n17661), .Z(n17498) );
  NOR U17822 ( .A(n17660), .B(n17498), .Z(n17663) );
  IV U17823 ( .A(n17499), .Z(n17501) );
  XOR U17824 ( .A(n17501), .B(n17500), .Z(n17656) );
  NOR U17825 ( .A(n108), .B(n59), .Z(n17657) );
  IV U17826 ( .A(n17657), .Z(n17502) );
  NOR U17827 ( .A(n17656), .B(n17502), .Z(n17659) );
  XOR U17828 ( .A(n17504), .B(n17503), .Z(n17652) );
  IV U17829 ( .A(n17652), .Z(n17506) );
  NOR U17830 ( .A(n87), .B(n59), .Z(n17505) );
  IV U17831 ( .A(n17505), .Z(n17653) );
  NOR U17832 ( .A(n17506), .B(n17653), .Z(n17655) );
  IV U17833 ( .A(n17507), .Z(n17509) );
  XOR U17834 ( .A(n17509), .B(n17508), .Z(n17648) );
  NOR U17835 ( .A(n107), .B(n59), .Z(n17649) );
  IV U17836 ( .A(n17649), .Z(n17510) );
  NOR U17837 ( .A(n17648), .B(n17510), .Z(n17651) );
  XOR U17838 ( .A(n17512), .B(n17511), .Z(n17644) );
  IV U17839 ( .A(n17644), .Z(n17514) );
  NOR U17840 ( .A(n88), .B(n59), .Z(n17513) );
  IV U17841 ( .A(n17513), .Z(n17645) );
  NOR U17842 ( .A(n17514), .B(n17645), .Z(n17647) );
  XOR U17843 ( .A(n17516), .B(n17515), .Z(n17632) );
  NOR U17844 ( .A(n105), .B(n59), .Z(n17633) );
  IV U17845 ( .A(n17633), .Z(n17517) );
  NOR U17846 ( .A(n17632), .B(n17517), .Z(n17635) );
  IV U17847 ( .A(n17518), .Z(n17520) );
  XOR U17848 ( .A(n17520), .B(n17519), .Z(n17628) );
  NOR U17849 ( .A(n104), .B(n59), .Z(n17629) );
  IV U17850 ( .A(n17629), .Z(n17521) );
  NOR U17851 ( .A(n17628), .B(n17521), .Z(n17631) );
  XOR U17852 ( .A(n17523), .B(n17522), .Z(n17624) );
  IV U17853 ( .A(n17624), .Z(n17525) );
  NOR U17854 ( .A(n89), .B(n59), .Z(n17524) );
  IV U17855 ( .A(n17524), .Z(n17625) );
  NOR U17856 ( .A(n17525), .B(n17625), .Z(n17627) );
  IV U17857 ( .A(n17526), .Z(n17528) );
  XOR U17858 ( .A(n17528), .B(n17527), .Z(n17620) );
  NOR U17859 ( .A(n103), .B(n59), .Z(n17621) );
  IV U17860 ( .A(n17621), .Z(n17529) );
  NOR U17861 ( .A(n17620), .B(n17529), .Z(n17623) );
  IV U17862 ( .A(n17530), .Z(n17532) );
  XOR U17863 ( .A(n17532), .B(n17531), .Z(n17616) );
  NOR U17864 ( .A(n90), .B(n59), .Z(n17617) );
  IV U17865 ( .A(n17617), .Z(n17533) );
  NOR U17866 ( .A(n17616), .B(n17533), .Z(n17619) );
  IV U17867 ( .A(n17534), .Z(n17536) );
  XOR U17868 ( .A(n17536), .B(n17535), .Z(n17612) );
  NOR U17869 ( .A(n102), .B(n59), .Z(n17613) );
  IV U17870 ( .A(n17613), .Z(n17537) );
  NOR U17871 ( .A(n17612), .B(n17537), .Z(n17615) );
  IV U17872 ( .A(n17538), .Z(n17540) );
  XOR U17873 ( .A(n17540), .B(n17539), .Z(n17608) );
  NOR U17874 ( .A(n101), .B(n59), .Z(n17609) );
  IV U17875 ( .A(n17609), .Z(n17541) );
  NOR U17876 ( .A(n17608), .B(n17541), .Z(n17611) );
  IV U17877 ( .A(n17542), .Z(n17544) );
  XOR U17878 ( .A(n17544), .B(n17543), .Z(n17604) );
  NOR U17879 ( .A(n100), .B(n59), .Z(n17605) );
  IV U17880 ( .A(n17605), .Z(n17545) );
  NOR U17881 ( .A(n17604), .B(n17545), .Z(n17607) );
  IV U17882 ( .A(n17546), .Z(n17548) );
  XOR U17883 ( .A(n17548), .B(n17547), .Z(n17600) );
  NOR U17884 ( .A(n99), .B(n59), .Z(n17601) );
  IV U17885 ( .A(n17601), .Z(n17549) );
  NOR U17886 ( .A(n17600), .B(n17549), .Z(n17603) );
  IV U17887 ( .A(n17550), .Z(n17552) );
  XOR U17888 ( .A(n17552), .B(n17551), .Z(n17596) );
  NOR U17889 ( .A(n98), .B(n59), .Z(n17597) );
  IV U17890 ( .A(n17597), .Z(n17553) );
  NOR U17891 ( .A(n17596), .B(n17553), .Z(n17599) );
  XOR U17892 ( .A(n17555), .B(n17554), .Z(n17592) );
  NOR U17893 ( .A(n91), .B(n59), .Z(n17593) );
  IV U17894 ( .A(n17593), .Z(n17556) );
  NOR U17895 ( .A(n17592), .B(n17556), .Z(n17595) );
  XOR U17896 ( .A(n17558), .B(n17557), .Z(n17580) );
  IV U17897 ( .A(n17580), .Z(n17560) );
  NOR U17898 ( .A(n96), .B(n59), .Z(n17559) );
  IV U17899 ( .A(n17559), .Z(n17581) );
  NOR U17900 ( .A(n17560), .B(n17581), .Z(n17583) );
  NOR U17901 ( .A(n95), .B(n59), .Z(n17577) );
  IV U17902 ( .A(n17577), .Z(n17563) );
  XOR U17903 ( .A(n17562), .B(n17561), .Z(n17576) );
  NOR U17904 ( .A(n17563), .B(n17576), .Z(n17579) );
  NOR U17905 ( .A(n59), .B(n93), .Z(n18599) );
  IV U17906 ( .A(n18599), .Z(n17564) );
  NOR U17907 ( .A(n58), .B(n168), .Z(n17572) );
  IV U17908 ( .A(n17572), .Z(n17567) );
  NOR U17909 ( .A(n17564), .B(n17567), .Z(n17565) );
  IV U17910 ( .A(n17565), .Z(n17566) );
  NOR U17911 ( .A(n94), .B(n17566), .Z(n17575) );
  NOR U17912 ( .A(n17567), .B(n93), .Z(n17568) );
  XOR U17913 ( .A(n94), .B(n17568), .Z(n17569) );
  NOR U17914 ( .A(n59), .B(n17569), .Z(n17570) );
  IV U17915 ( .A(n17570), .Z(n18070) );
  XOR U17916 ( .A(n17572), .B(n17571), .Z(n18069) );
  IV U17917 ( .A(n18069), .Z(n17573) );
  NOR U17918 ( .A(n18070), .B(n17573), .Z(n17574) );
  NOR U17919 ( .A(n17575), .B(n17574), .Z(n18066) );
  XOR U17920 ( .A(n17577), .B(n17576), .Z(n18065) );
  NOR U17921 ( .A(n18066), .B(n18065), .Z(n17578) );
  NOR U17922 ( .A(n17579), .B(n17578), .Z(n18093) );
  XOR U17923 ( .A(n17581), .B(n17580), .Z(n18092) );
  NOR U17924 ( .A(n18093), .B(n18092), .Z(n17582) );
  NOR U17925 ( .A(n17583), .B(n17582), .Z(n17588) );
  XOR U17926 ( .A(n17585), .B(n17584), .Z(n17587) );
  IV U17927 ( .A(n17587), .Z(n17586) );
  NOR U17928 ( .A(n17588), .B(n17586), .Z(n17591) );
  XOR U17929 ( .A(n17588), .B(n17587), .Z(n18062) );
  NOR U17930 ( .A(n97), .B(n59), .Z(n18063) );
  IV U17931 ( .A(n18063), .Z(n17589) );
  NOR U17932 ( .A(n18062), .B(n17589), .Z(n17590) );
  NOR U17933 ( .A(n17591), .B(n17590), .Z(n18058) );
  XOR U17934 ( .A(n17593), .B(n17592), .Z(n18059) );
  NOR U17935 ( .A(n18058), .B(n18059), .Z(n17594) );
  NOR U17936 ( .A(n17595), .B(n17594), .Z(n18054) );
  XOR U17937 ( .A(n17597), .B(n17596), .Z(n18055) );
  NOR U17938 ( .A(n18054), .B(n18055), .Z(n17598) );
  NOR U17939 ( .A(n17599), .B(n17598), .Z(n18050) );
  XOR U17940 ( .A(n17601), .B(n17600), .Z(n18051) );
  NOR U17941 ( .A(n18050), .B(n18051), .Z(n17602) );
  NOR U17942 ( .A(n17603), .B(n17602), .Z(n18046) );
  XOR U17943 ( .A(n17605), .B(n17604), .Z(n18047) );
  NOR U17944 ( .A(n18046), .B(n18047), .Z(n17606) );
  NOR U17945 ( .A(n17607), .B(n17606), .Z(n18042) );
  XOR U17946 ( .A(n17609), .B(n17608), .Z(n18043) );
  NOR U17947 ( .A(n18042), .B(n18043), .Z(n17610) );
  NOR U17948 ( .A(n17611), .B(n17610), .Z(n18038) );
  XOR U17949 ( .A(n17613), .B(n17612), .Z(n18039) );
  NOR U17950 ( .A(n18038), .B(n18039), .Z(n17614) );
  NOR U17951 ( .A(n17615), .B(n17614), .Z(n18034) );
  XOR U17952 ( .A(n17617), .B(n17616), .Z(n18035) );
  NOR U17953 ( .A(n18034), .B(n18035), .Z(n17618) );
  NOR U17954 ( .A(n17619), .B(n17618), .Z(n18031) );
  XOR U17955 ( .A(n17621), .B(n17620), .Z(n18030) );
  NOR U17956 ( .A(n18031), .B(n18030), .Z(n17622) );
  NOR U17957 ( .A(n17623), .B(n17622), .Z(n18137) );
  XOR U17958 ( .A(n17625), .B(n17624), .Z(n18136) );
  NOR U17959 ( .A(n18137), .B(n18136), .Z(n17626) );
  NOR U17960 ( .A(n17627), .B(n17626), .Z(n18026) );
  XOR U17961 ( .A(n17629), .B(n17628), .Z(n18027) );
  NOR U17962 ( .A(n18026), .B(n18027), .Z(n17630) );
  NOR U17963 ( .A(n17631), .B(n17630), .Z(n18022) );
  XOR U17964 ( .A(n17633), .B(n17632), .Z(n18023) );
  NOR U17965 ( .A(n18022), .B(n18023), .Z(n17634) );
  NOR U17966 ( .A(n17635), .B(n17634), .Z(n17640) );
  XOR U17967 ( .A(n17637), .B(n17636), .Z(n17639) );
  IV U17968 ( .A(n17639), .Z(n17638) );
  NOR U17969 ( .A(n17640), .B(n17638), .Z(n17643) );
  XOR U17970 ( .A(n17640), .B(n17639), .Z(n18019) );
  NOR U17971 ( .A(n106), .B(n59), .Z(n18020) );
  IV U17972 ( .A(n18020), .Z(n17641) );
  NOR U17973 ( .A(n18019), .B(n17641), .Z(n17642) );
  NOR U17974 ( .A(n17643), .B(n17642), .Z(n18157) );
  XOR U17975 ( .A(n17645), .B(n17644), .Z(n18156) );
  NOR U17976 ( .A(n18157), .B(n18156), .Z(n17646) );
  NOR U17977 ( .A(n17647), .B(n17646), .Z(n18015) );
  XOR U17978 ( .A(n17649), .B(n17648), .Z(n18016) );
  NOR U17979 ( .A(n18015), .B(n18016), .Z(n17650) );
  NOR U17980 ( .A(n17651), .B(n17650), .Z(n18172) );
  XOR U17981 ( .A(n17653), .B(n17652), .Z(n18171) );
  NOR U17982 ( .A(n18172), .B(n18171), .Z(n17654) );
  NOR U17983 ( .A(n17655), .B(n17654), .Z(n18011) );
  XOR U17984 ( .A(n17657), .B(n17656), .Z(n18012) );
  NOR U17985 ( .A(n18011), .B(n18012), .Z(n17658) );
  NOR U17986 ( .A(n17659), .B(n17658), .Z(n18007) );
  XOR U17987 ( .A(n17661), .B(n17660), .Z(n18008) );
  NOR U17988 ( .A(n18007), .B(n18008), .Z(n17662) );
  NOR U17989 ( .A(n17663), .B(n17662), .Z(n18006) );
  XOR U17990 ( .A(n17665), .B(n17664), .Z(n18005) );
  NOR U17991 ( .A(n18006), .B(n18005), .Z(n17666) );
  NOR U17992 ( .A(n17667), .B(n17666), .Z(n17668) );
  IV U17993 ( .A(n17668), .Z(n18003) );
  XOR U17994 ( .A(n17670), .B(n17669), .Z(n17671) );
  IV U17995 ( .A(n17671), .Z(n18002) );
  NOR U17996 ( .A(n18003), .B(n18002), .Z(n17672) );
  NOR U17997 ( .A(n17673), .B(n17672), .Z(n17674) );
  IV U17998 ( .A(n17674), .Z(n17998) );
  XOR U17999 ( .A(n17676), .B(n17675), .Z(n17997) );
  NOR U18000 ( .A(n17998), .B(n17997), .Z(n17677) );
  NOR U18001 ( .A(n17678), .B(n17677), .Z(n17679) );
  IV U18002 ( .A(n17679), .Z(n17995) );
  XOR U18003 ( .A(n17681), .B(n17680), .Z(n17682) );
  IV U18004 ( .A(n17682), .Z(n17994) );
  NOR U18005 ( .A(n17995), .B(n17994), .Z(n17683) );
  NOR U18006 ( .A(n17684), .B(n17683), .Z(n17685) );
  IV U18007 ( .A(n17685), .Z(n17993) );
  XOR U18008 ( .A(n17687), .B(n17686), .Z(n17992) );
  NOR U18009 ( .A(n17993), .B(n17992), .Z(n17688) );
  NOR U18010 ( .A(n17689), .B(n17688), .Z(n17690) );
  IV U18011 ( .A(n17690), .Z(n17990) );
  XOR U18012 ( .A(n17692), .B(n17691), .Z(n17693) );
  IV U18013 ( .A(n17693), .Z(n17989) );
  NOR U18014 ( .A(n17990), .B(n17989), .Z(n17694) );
  NOR U18015 ( .A(n17695), .B(n17694), .Z(n17696) );
  IV U18016 ( .A(n17696), .Z(n17988) );
  XOR U18017 ( .A(n17698), .B(n17697), .Z(n17987) );
  NOR U18018 ( .A(n17988), .B(n17987), .Z(n17699) );
  NOR U18019 ( .A(n17700), .B(n17699), .Z(n17985) );
  NOR U18020 ( .A(n17702), .B(n17701), .Z(n17703) );
  NOR U18021 ( .A(n17985), .B(n17703), .Z(n17704) );
  NOR U18022 ( .A(n17705), .B(n17704), .Z(n17710) );
  NOR U18023 ( .A(n114), .B(n59), .Z(n17709) );
  IV U18024 ( .A(n17709), .Z(n17706) );
  NOR U18025 ( .A(n17710), .B(n17706), .Z(n17712) );
  XOR U18026 ( .A(n17708), .B(n17707), .Z(n17981) );
  XOR U18027 ( .A(n17710), .B(n17709), .Z(n17980) );
  NOR U18028 ( .A(n17981), .B(n17980), .Z(n17711) );
  NOR U18029 ( .A(n17712), .B(n17711), .Z(n18231) );
  XOR U18030 ( .A(n17714), .B(n17713), .Z(n18232) );
  IV U18031 ( .A(n18232), .Z(n17715) );
  NOR U18032 ( .A(n18231), .B(n17715), .Z(n17716) );
  NOR U18033 ( .A(n17717), .B(n17716), .Z(n17976) );
  XOR U18034 ( .A(n17719), .B(n17718), .Z(n17977) );
  NOR U18035 ( .A(n17976), .B(n17977), .Z(n17720) );
  NOR U18036 ( .A(n17721), .B(n17720), .Z(n17974) );
  NOR U18037 ( .A(n17723), .B(n17722), .Z(n17724) );
  NOR U18038 ( .A(n17974), .B(n17724), .Z(n17725) );
  NOR U18039 ( .A(n17726), .B(n17725), .Z(n17733) );
  NOR U18040 ( .A(n116), .B(n59), .Z(n17732) );
  IV U18041 ( .A(n17732), .Z(n17727) );
  NOR U18042 ( .A(n17733), .B(n17727), .Z(n17735) );
  XOR U18043 ( .A(n17729), .B(n17728), .Z(n17730) );
  XOR U18044 ( .A(n17731), .B(n17730), .Z(n17970) );
  XOR U18045 ( .A(n17733), .B(n17732), .Z(n17969) );
  NOR U18046 ( .A(n17970), .B(n17969), .Z(n17734) );
  NOR U18047 ( .A(n17735), .B(n17734), .Z(n18254) );
  IV U18048 ( .A(n18254), .Z(n17736) );
  NOR U18049 ( .A(n17737), .B(n17736), .Z(n17738) );
  NOR U18050 ( .A(n17739), .B(n17738), .Z(n17740) );
  IV U18051 ( .A(n17740), .Z(n17747) );
  NOR U18052 ( .A(n117), .B(n59), .Z(n17746) );
  IV U18053 ( .A(n17746), .Z(n17741) );
  NOR U18054 ( .A(n17747), .B(n17741), .Z(n17749) );
  XOR U18055 ( .A(n17743), .B(n17742), .Z(n17744) );
  XOR U18056 ( .A(n17745), .B(n17744), .Z(n17965) );
  XOR U18057 ( .A(n17747), .B(n17746), .Z(n17966) );
  NOR U18058 ( .A(n17965), .B(n17966), .Z(n17748) );
  NOR U18059 ( .A(n17749), .B(n17748), .Z(n18267) );
  IV U18060 ( .A(n18267), .Z(n17750) );
  NOR U18061 ( .A(n17751), .B(n17750), .Z(n17752) );
  NOR U18062 ( .A(n17753), .B(n17752), .Z(n17754) );
  IV U18063 ( .A(n17754), .Z(n17761) );
  NOR U18064 ( .A(n119), .B(n59), .Z(n17760) );
  IV U18065 ( .A(n17760), .Z(n17755) );
  NOR U18066 ( .A(n17761), .B(n17755), .Z(n17763) );
  XOR U18067 ( .A(n17757), .B(n17756), .Z(n17758) );
  XOR U18068 ( .A(n17759), .B(n17758), .Z(n17960) );
  XOR U18069 ( .A(n17761), .B(n17760), .Z(n17961) );
  NOR U18070 ( .A(n17960), .B(n17961), .Z(n17762) );
  NOR U18071 ( .A(n17763), .B(n17762), .Z(n18280) );
  IV U18072 ( .A(n18280), .Z(n17764) );
  NOR U18073 ( .A(n17765), .B(n17764), .Z(n17766) );
  NOR U18074 ( .A(n17767), .B(n17766), .Z(n17773) );
  IV U18075 ( .A(n17773), .Z(n17768) );
  NOR U18076 ( .A(n17774), .B(n17768), .Z(n17776) );
  XOR U18077 ( .A(n17770), .B(n17769), .Z(n17771) );
  XOR U18078 ( .A(n17772), .B(n17771), .Z(n17955) );
  XOR U18079 ( .A(n17774), .B(n17773), .Z(n17956) );
  NOR U18080 ( .A(n17955), .B(n17956), .Z(n17775) );
  NOR U18081 ( .A(n17776), .B(n17775), .Z(n18294) );
  NOR U18082 ( .A(n17778), .B(n17777), .Z(n17779) );
  NOR U18083 ( .A(n18294), .B(n17779), .Z(n17780) );
  NOR U18084 ( .A(n17781), .B(n17780), .Z(n17786) );
  NOR U18085 ( .A(n126), .B(n59), .Z(n17785) );
  IV U18086 ( .A(n17785), .Z(n17782) );
  NOR U18087 ( .A(n17786), .B(n17782), .Z(n17789) );
  XOR U18088 ( .A(n17784), .B(n17783), .Z(n17953) );
  IV U18089 ( .A(n17953), .Z(n17787) );
  XOR U18090 ( .A(n17786), .B(n17785), .Z(n17952) );
  NOR U18091 ( .A(n17787), .B(n17952), .Z(n17788) );
  NOR U18092 ( .A(n17789), .B(n17788), .Z(n17794) );
  NOR U18093 ( .A(n128), .B(n59), .Z(n17793) );
  IV U18094 ( .A(n17793), .Z(n17790) );
  NOR U18095 ( .A(n17794), .B(n17790), .Z(n17796) );
  XOR U18096 ( .A(n17792), .B(n17791), .Z(n18304) );
  XOR U18097 ( .A(n17794), .B(n17793), .Z(n18303) );
  NOR U18098 ( .A(n18304), .B(n18303), .Z(n17795) );
  NOR U18099 ( .A(n17796), .B(n17795), .Z(n17803) );
  NOR U18100 ( .A(n131), .B(n59), .Z(n17802) );
  IV U18101 ( .A(n17802), .Z(n17797) );
  NOR U18102 ( .A(n17803), .B(n17797), .Z(n17805) );
  XOR U18103 ( .A(n17799), .B(n17798), .Z(n17800) );
  XOR U18104 ( .A(n17801), .B(n17800), .Z(n17948) );
  XOR U18105 ( .A(n17803), .B(n17802), .Z(n17949) );
  NOR U18106 ( .A(n17948), .B(n17949), .Z(n17804) );
  NOR U18107 ( .A(n17805), .B(n17804), .Z(n17809) );
  XOR U18108 ( .A(n17807), .B(n17806), .Z(n18317) );
  IV U18109 ( .A(n18317), .Z(n17808) );
  NOR U18110 ( .A(n17809), .B(n17808), .Z(n17813) );
  IV U18111 ( .A(n17809), .Z(n18318) );
  NOR U18112 ( .A(n18318), .B(n18317), .Z(n17811) );
  NOR U18113 ( .A(n133), .B(n59), .Z(n18320) );
  IV U18114 ( .A(n18320), .Z(n17810) );
  NOR U18115 ( .A(n17811), .B(n17810), .Z(n17812) );
  NOR U18116 ( .A(n17813), .B(n17812), .Z(n17815) );
  IV U18117 ( .A(n17815), .Z(n18326) );
  NOR U18118 ( .A(n17814), .B(n18326), .Z(n17822) );
  IV U18119 ( .A(n17814), .Z(n18327) );
  NOR U18120 ( .A(n17815), .B(n18327), .Z(n17820) );
  XOR U18121 ( .A(n17817), .B(n17816), .Z(n17818) );
  XOR U18122 ( .A(n17819), .B(n17818), .Z(n18329) );
  NOR U18123 ( .A(n17820), .B(n18329), .Z(n17821) );
  NOR U18124 ( .A(n17822), .B(n17821), .Z(n17830) );
  IV U18125 ( .A(n17830), .Z(n17824) );
  NOR U18126 ( .A(n137), .B(n59), .Z(n17823) );
  IV U18127 ( .A(n17823), .Z(n17829) );
  NOR U18128 ( .A(n17824), .B(n17829), .Z(n17832) );
  XOR U18129 ( .A(n17826), .B(n17825), .Z(n17827) );
  XOR U18130 ( .A(n17828), .B(n17827), .Z(n18334) );
  XOR U18131 ( .A(n17830), .B(n17829), .Z(n18335) );
  NOR U18132 ( .A(n18334), .B(n18335), .Z(n17831) );
  NOR U18133 ( .A(n17832), .B(n17831), .Z(n17836) );
  XOR U18134 ( .A(n17834), .B(n17833), .Z(n17835) );
  NOR U18135 ( .A(n17836), .B(n17835), .Z(n17840) );
  XOR U18136 ( .A(n17836), .B(n17835), .Z(n18342) );
  IV U18137 ( .A(n18342), .Z(n17838) );
  NOR U18138 ( .A(n139), .B(n59), .Z(n18343) );
  IV U18139 ( .A(n18343), .Z(n17837) );
  NOR U18140 ( .A(n17838), .B(n17837), .Z(n17839) );
  NOR U18141 ( .A(n17840), .B(n17839), .Z(n18352) );
  XOR U18142 ( .A(n17842), .B(n17841), .Z(n18351) );
  NOR U18143 ( .A(n18352), .B(n18351), .Z(n17843) );
  NOR U18144 ( .A(n17844), .B(n17843), .Z(n17849) );
  XOR U18145 ( .A(n17846), .B(n17845), .Z(n17848) );
  IV U18146 ( .A(n17848), .Z(n17847) );
  NOR U18147 ( .A(n17849), .B(n17847), .Z(n17852) );
  XOR U18148 ( .A(n17849), .B(n17848), .Z(n18359) );
  NOR U18149 ( .A(n143), .B(n59), .Z(n17850) );
  IV U18150 ( .A(n17850), .Z(n18358) );
  NOR U18151 ( .A(n18359), .B(n18358), .Z(n17851) );
  NOR U18152 ( .A(n17852), .B(n17851), .Z(n17859) );
  NOR U18153 ( .A(n145), .B(n59), .Z(n17858) );
  IV U18154 ( .A(n17858), .Z(n17853) );
  NOR U18155 ( .A(n17859), .B(n17853), .Z(n17861) );
  XOR U18156 ( .A(n17855), .B(n17854), .Z(n17856) );
  XOR U18157 ( .A(n17857), .B(n17856), .Z(n18370) );
  XOR U18158 ( .A(n17859), .B(n17858), .Z(n18369) );
  NOR U18159 ( .A(n18370), .B(n18369), .Z(n17860) );
  NOR U18160 ( .A(n17861), .B(n17860), .Z(n17864) );
  XOR U18161 ( .A(n17863), .B(n17862), .Z(n17865) );
  NOR U18162 ( .A(n17864), .B(n17865), .Z(n17869) );
  IV U18163 ( .A(n17864), .Z(n17866) );
  XOR U18164 ( .A(n17866), .B(n17865), .Z(n18377) );
  NOR U18165 ( .A(n147), .B(n59), .Z(n18378) );
  IV U18166 ( .A(n18378), .Z(n17867) );
  NOR U18167 ( .A(n18377), .B(n17867), .Z(n17868) );
  NOR U18168 ( .A(n17869), .B(n17868), .Z(n17872) );
  NOR U18169 ( .A(n148), .B(n59), .Z(n17871) );
  IV U18170 ( .A(n17871), .Z(n17870) );
  NOR U18171 ( .A(n17872), .B(n17870), .Z(n17877) );
  XOR U18172 ( .A(n17872), .B(n17871), .Z(n18382) );
  XOR U18173 ( .A(n17874), .B(n17873), .Z(n18383) );
  IV U18174 ( .A(n18383), .Z(n17875) );
  NOR U18175 ( .A(n18382), .B(n17875), .Z(n17876) );
  NOR U18176 ( .A(n17877), .B(n17876), .Z(n17880) );
  NOR U18177 ( .A(n150), .B(n59), .Z(n17879) );
  IV U18178 ( .A(n17879), .Z(n17878) );
  NOR U18179 ( .A(n17880), .B(n17878), .Z(n17885) );
  XOR U18180 ( .A(n17880), .B(n17879), .Z(n18388) );
  XOR U18181 ( .A(n17882), .B(n17881), .Z(n18389) );
  IV U18182 ( .A(n18389), .Z(n17883) );
  NOR U18183 ( .A(n18388), .B(n17883), .Z(n17884) );
  NOR U18184 ( .A(n17885), .B(n17884), .Z(n17889) );
  XOR U18185 ( .A(n17887), .B(n17886), .Z(n17888) );
  NOR U18186 ( .A(n17889), .B(n17888), .Z(n17893) );
  XOR U18187 ( .A(n17889), .B(n17888), .Z(n18399) );
  IV U18188 ( .A(n18399), .Z(n17891) );
  NOR U18189 ( .A(n153), .B(n59), .Z(n17890) );
  IV U18190 ( .A(n17890), .Z(n18400) );
  NOR U18191 ( .A(n17891), .B(n18400), .Z(n17892) );
  NOR U18192 ( .A(n17893), .B(n17892), .Z(n18405) );
  XOR U18193 ( .A(n17895), .B(n17894), .Z(n18404) );
  NOR U18194 ( .A(n18405), .B(n18404), .Z(n17896) );
  NOR U18195 ( .A(n17897), .B(n17896), .Z(n17900) );
  NOR U18196 ( .A(n156), .B(n59), .Z(n17899) );
  IV U18197 ( .A(n17899), .Z(n17898) );
  NOR U18198 ( .A(n17900), .B(n17898), .Z(n17905) );
  XOR U18199 ( .A(n17900), .B(n17899), .Z(n18411) );
  XOR U18200 ( .A(n17902), .B(n17901), .Z(n18412) );
  IV U18201 ( .A(n18412), .Z(n17903) );
  NOR U18202 ( .A(n18411), .B(n17903), .Z(n17904) );
  NOR U18203 ( .A(n17905), .B(n17904), .Z(n17909) );
  XOR U18204 ( .A(n17907), .B(n17906), .Z(n17908) );
  NOR U18205 ( .A(n17909), .B(n17908), .Z(n17913) );
  XOR U18206 ( .A(n17909), .B(n17908), .Z(n18422) );
  IV U18207 ( .A(n18422), .Z(n17911) );
  NOR U18208 ( .A(n158), .B(n59), .Z(n17910) );
  IV U18209 ( .A(n17910), .Z(n18423) );
  NOR U18210 ( .A(n17911), .B(n18423), .Z(n17912) );
  NOR U18211 ( .A(n17913), .B(n17912), .Z(n17916) );
  NOR U18212 ( .A(n161), .B(n59), .Z(n17915) );
  IV U18213 ( .A(n17915), .Z(n17914) );
  NOR U18214 ( .A(n17916), .B(n17914), .Z(n17920) );
  XOR U18215 ( .A(n17916), .B(n17915), .Z(n18427) );
  XOR U18216 ( .A(n17918), .B(n17917), .Z(n18428) );
  NOR U18217 ( .A(n18427), .B(n18428), .Z(n17919) );
  NOR U18218 ( .A(n17920), .B(n17919), .Z(n17923) );
  NOR U18219 ( .A(n163), .B(n59), .Z(n17922) );
  IV U18220 ( .A(n17922), .Z(n17921) );
  NOR U18221 ( .A(n17923), .B(n17921), .Z(n17928) );
  XOR U18222 ( .A(n17923), .B(n17922), .Z(n18434) );
  XOR U18223 ( .A(n17925), .B(n17924), .Z(n18435) );
  IV U18224 ( .A(n18435), .Z(n17926) );
  NOR U18225 ( .A(n18434), .B(n17926), .Z(n17927) );
  NOR U18226 ( .A(n17928), .B(n17927), .Z(n17932) );
  XOR U18227 ( .A(n17930), .B(n17929), .Z(n17931) );
  NOR U18228 ( .A(n17932), .B(n17931), .Z(n17936) );
  XOR U18229 ( .A(n17932), .B(n17931), .Z(n18445) );
  IV U18230 ( .A(n18445), .Z(n17934) );
  NOR U18231 ( .A(n165), .B(n59), .Z(n17933) );
  IV U18232 ( .A(n17933), .Z(n18446) );
  NOR U18233 ( .A(n17934), .B(n18446), .Z(n17935) );
  NOR U18234 ( .A(n17936), .B(n17935), .Z(n17947) );
  XOR U18235 ( .A(n17938), .B(n17937), .Z(n17946) );
  NOR U18236 ( .A(n17947), .B(n17946), .Z(n17939) );
  NOR U18237 ( .A(n17940), .B(n17939), .Z(n18450) );
  XOR U18238 ( .A(n17942), .B(n17941), .Z(n18449) );
  NOR U18239 ( .A(n18450), .B(n18449), .Z(n31588) );
  NOR U18240 ( .A(n28570), .B(n31588), .Z(n17943) );
  NOR U18241 ( .A(n17944), .B(n17943), .Z(n17945) );
  IV U18242 ( .A(n17945), .Z(n28569) );
  XOR U18243 ( .A(n17947), .B(n17946), .Z(n31581) );
  IV U18244 ( .A(n31581), .Z(n18452) );
  NOR U18245 ( .A(n145), .B(n60), .Z(n18360) );
  NOR U18246 ( .A(n135), .B(n60), .Z(n18315) );
  IV U18247 ( .A(n17948), .Z(n17950) );
  XOR U18248 ( .A(n17950), .B(n17949), .Z(n18311) );
  NOR U18249 ( .A(n133), .B(n60), .Z(n18312) );
  IV U18250 ( .A(n18312), .Z(n17951) );
  NOR U18251 ( .A(n18311), .B(n17951), .Z(n18314) );
  XOR U18252 ( .A(n17953), .B(n17952), .Z(n18299) );
  NOR U18253 ( .A(n128), .B(n60), .Z(n18300) );
  IV U18254 ( .A(n18300), .Z(n17954) );
  NOR U18255 ( .A(n18299), .B(n17954), .Z(n18302) );
  XOR U18256 ( .A(n17956), .B(n17955), .Z(n17957) );
  NOR U18257 ( .A(n125), .B(n60), .Z(n18811) );
  NOR U18258 ( .A(n17957), .B(n18811), .Z(n18288) );
  IV U18259 ( .A(n17957), .Z(n18808) );
  IV U18260 ( .A(n18811), .Z(n17958) );
  NOR U18261 ( .A(n18808), .B(n17958), .Z(n18286) );
  NOR U18262 ( .A(n123), .B(n60), .Z(n17959) );
  IV U18263 ( .A(n17959), .Z(n18282) );
  NOR U18264 ( .A(n120), .B(n60), .Z(n17962) );
  XOR U18265 ( .A(n17961), .B(n17960), .Z(n17963) );
  NOR U18266 ( .A(n17962), .B(n17963), .Z(n18275) );
  IV U18267 ( .A(n17962), .Z(n18795) );
  IV U18268 ( .A(n17963), .Z(n18794) );
  NOR U18269 ( .A(n18795), .B(n18794), .Z(n18273) );
  NOR U18270 ( .A(n119), .B(n60), .Z(n17964) );
  IV U18271 ( .A(n17964), .Z(n18269) );
  XOR U18272 ( .A(n17966), .B(n17965), .Z(n17967) );
  NOR U18273 ( .A(n79), .B(n60), .Z(n17968) );
  NOR U18274 ( .A(n17967), .B(n17968), .Z(n18262) );
  IV U18275 ( .A(n17967), .Z(n18779) );
  IV U18276 ( .A(n17968), .Z(n18778) );
  NOR U18277 ( .A(n18779), .B(n18778), .Z(n18260) );
  XOR U18278 ( .A(n17970), .B(n17969), .Z(n18246) );
  IV U18279 ( .A(n18246), .Z(n18484) );
  NOR U18280 ( .A(n80), .B(n60), .Z(n18245) );
  IV U18281 ( .A(n18245), .Z(n18483) );
  NOR U18282 ( .A(n18484), .B(n18483), .Z(n18249) );
  XOR U18283 ( .A(n17972), .B(n17971), .Z(n17973) );
  XOR U18284 ( .A(n17974), .B(n17973), .Z(n18242) );
  NOR U18285 ( .A(n116), .B(n60), .Z(n18241) );
  IV U18286 ( .A(n18241), .Z(n17975) );
  NOR U18287 ( .A(n18242), .B(n17975), .Z(n18244) );
  IV U18288 ( .A(n17976), .Z(n17978) );
  XOR U18289 ( .A(n17978), .B(n17977), .Z(n18237) );
  NOR U18290 ( .A(n81), .B(n60), .Z(n18238) );
  IV U18291 ( .A(n18238), .Z(n17979) );
  NOR U18292 ( .A(n18237), .B(n17979), .Z(n18240) );
  XOR U18293 ( .A(n17981), .B(n17980), .Z(n18226) );
  IV U18294 ( .A(n18226), .Z(n18495) );
  NOR U18295 ( .A(n82), .B(n60), .Z(n18225) );
  IV U18296 ( .A(n18225), .Z(n18494) );
  NOR U18297 ( .A(n18495), .B(n18494), .Z(n18229) );
  XOR U18298 ( .A(n17983), .B(n17982), .Z(n17984) );
  XOR U18299 ( .A(n17985), .B(n17984), .Z(n18222) );
  NOR U18300 ( .A(n114), .B(n60), .Z(n18221) );
  IV U18301 ( .A(n18221), .Z(n17986) );
  NOR U18302 ( .A(n18222), .B(n17986), .Z(n18224) );
  NOR U18303 ( .A(n83), .B(n60), .Z(n18216) );
  XOR U18304 ( .A(n17988), .B(n17987), .Z(n18215) );
  NOR U18305 ( .A(n18216), .B(n18215), .Z(n18219) );
  XOR U18306 ( .A(n17990), .B(n17989), .Z(n18211) );
  NOR U18307 ( .A(n113), .B(n60), .Z(n18210) );
  IV U18308 ( .A(n18210), .Z(n17991) );
  NOR U18309 ( .A(n18211), .B(n17991), .Z(n18213) );
  NOR U18310 ( .A(n84), .B(n60), .Z(n18205) );
  XOR U18311 ( .A(n17993), .B(n17992), .Z(n18204) );
  NOR U18312 ( .A(n18205), .B(n18204), .Z(n18208) );
  XOR U18313 ( .A(n17995), .B(n17994), .Z(n18200) );
  NOR U18314 ( .A(n112), .B(n60), .Z(n18199) );
  IV U18315 ( .A(n18199), .Z(n17996) );
  NOR U18316 ( .A(n18200), .B(n17996), .Z(n18202) );
  NOR U18317 ( .A(n85), .B(n60), .Z(n18000) );
  XOR U18318 ( .A(n17998), .B(n17997), .Z(n17999) );
  NOR U18319 ( .A(n18000), .B(n17999), .Z(n18197) );
  XOR U18320 ( .A(n18000), .B(n17999), .Z(n18001) );
  IV U18321 ( .A(n18001), .Z(n18512) );
  XOR U18322 ( .A(n18003), .B(n18002), .Z(n18192) );
  NOR U18323 ( .A(n111), .B(n60), .Z(n18191) );
  IV U18324 ( .A(n18191), .Z(n18004) );
  NOR U18325 ( .A(n18192), .B(n18004), .Z(n18194) );
  NOR U18326 ( .A(n86), .B(n60), .Z(n18186) );
  XOR U18327 ( .A(n18006), .B(n18005), .Z(n18185) );
  NOR U18328 ( .A(n18186), .B(n18185), .Z(n18189) );
  IV U18329 ( .A(n18007), .Z(n18009) );
  XOR U18330 ( .A(n18009), .B(n18008), .Z(n18180) );
  NOR U18331 ( .A(n110), .B(n60), .Z(n18181) );
  IV U18332 ( .A(n18181), .Z(n18010) );
  NOR U18333 ( .A(n18180), .B(n18010), .Z(n18183) );
  IV U18334 ( .A(n18011), .Z(n18013) );
  XOR U18335 ( .A(n18013), .B(n18012), .Z(n18176) );
  NOR U18336 ( .A(n109), .B(n60), .Z(n18177) );
  IV U18337 ( .A(n18177), .Z(n18014) );
  NOR U18338 ( .A(n18176), .B(n18014), .Z(n18179) );
  IV U18339 ( .A(n18015), .Z(n18017) );
  XOR U18340 ( .A(n18017), .B(n18016), .Z(n18164) );
  NOR U18341 ( .A(n87), .B(n60), .Z(n18165) );
  IV U18342 ( .A(n18165), .Z(n18018) );
  NOR U18343 ( .A(n18164), .B(n18018), .Z(n18167) );
  XOR U18344 ( .A(n18020), .B(n18019), .Z(n18152) );
  NOR U18345 ( .A(n88), .B(n60), .Z(n18153) );
  IV U18346 ( .A(n18153), .Z(n18021) );
  NOR U18347 ( .A(n18152), .B(n18021), .Z(n18155) );
  IV U18348 ( .A(n18022), .Z(n18024) );
  XOR U18349 ( .A(n18024), .B(n18023), .Z(n18148) );
  NOR U18350 ( .A(n106), .B(n60), .Z(n18149) );
  IV U18351 ( .A(n18149), .Z(n18025) );
  NOR U18352 ( .A(n18148), .B(n18025), .Z(n18151) );
  IV U18353 ( .A(n18026), .Z(n18028) );
  XOR U18354 ( .A(n18028), .B(n18027), .Z(n18144) );
  NOR U18355 ( .A(n105), .B(n60), .Z(n18145) );
  IV U18356 ( .A(n18145), .Z(n18029) );
  NOR U18357 ( .A(n18144), .B(n18029), .Z(n18147) );
  XOR U18358 ( .A(n18031), .B(n18030), .Z(n18132) );
  IV U18359 ( .A(n18132), .Z(n18033) );
  NOR U18360 ( .A(n89), .B(n60), .Z(n18032) );
  IV U18361 ( .A(n18032), .Z(n18133) );
  NOR U18362 ( .A(n18033), .B(n18133), .Z(n18135) );
  IV U18363 ( .A(n18034), .Z(n18036) );
  XOR U18364 ( .A(n18036), .B(n18035), .Z(n18128) );
  NOR U18365 ( .A(n103), .B(n60), .Z(n18129) );
  IV U18366 ( .A(n18129), .Z(n18037) );
  NOR U18367 ( .A(n18128), .B(n18037), .Z(n18131) );
  IV U18368 ( .A(n18038), .Z(n18040) );
  XOR U18369 ( .A(n18040), .B(n18039), .Z(n18124) );
  NOR U18370 ( .A(n90), .B(n60), .Z(n18125) );
  IV U18371 ( .A(n18125), .Z(n18041) );
  NOR U18372 ( .A(n18124), .B(n18041), .Z(n18127) );
  IV U18373 ( .A(n18042), .Z(n18044) );
  XOR U18374 ( .A(n18044), .B(n18043), .Z(n18120) );
  NOR U18375 ( .A(n102), .B(n60), .Z(n18121) );
  IV U18376 ( .A(n18121), .Z(n18045) );
  NOR U18377 ( .A(n18120), .B(n18045), .Z(n18123) );
  IV U18378 ( .A(n18046), .Z(n18048) );
  XOR U18379 ( .A(n18048), .B(n18047), .Z(n18116) );
  NOR U18380 ( .A(n101), .B(n60), .Z(n18117) );
  IV U18381 ( .A(n18117), .Z(n18049) );
  NOR U18382 ( .A(n18116), .B(n18049), .Z(n18119) );
  IV U18383 ( .A(n18050), .Z(n18052) );
  XOR U18384 ( .A(n18052), .B(n18051), .Z(n18112) );
  NOR U18385 ( .A(n100), .B(n60), .Z(n18113) );
  IV U18386 ( .A(n18113), .Z(n18053) );
  NOR U18387 ( .A(n18112), .B(n18053), .Z(n18115) );
  IV U18388 ( .A(n18054), .Z(n18056) );
  XOR U18389 ( .A(n18056), .B(n18055), .Z(n18108) );
  NOR U18390 ( .A(n99), .B(n60), .Z(n18109) );
  IV U18391 ( .A(n18109), .Z(n18057) );
  NOR U18392 ( .A(n18108), .B(n18057), .Z(n18111) );
  IV U18393 ( .A(n18058), .Z(n18060) );
  XOR U18394 ( .A(n18060), .B(n18059), .Z(n18104) );
  NOR U18395 ( .A(n98), .B(n60), .Z(n18105) );
  IV U18396 ( .A(n18105), .Z(n18061) );
  NOR U18397 ( .A(n18104), .B(n18061), .Z(n18107) );
  XOR U18398 ( .A(n18063), .B(n18062), .Z(n18100) );
  NOR U18399 ( .A(n91), .B(n60), .Z(n18101) );
  IV U18400 ( .A(n18101), .Z(n18064) );
  NOR U18401 ( .A(n18100), .B(n18064), .Z(n18103) );
  XOR U18402 ( .A(n18066), .B(n18065), .Z(n18088) );
  IV U18403 ( .A(n18088), .Z(n18068) );
  NOR U18404 ( .A(n96), .B(n60), .Z(n18067) );
  IV U18405 ( .A(n18067), .Z(n18089) );
  NOR U18406 ( .A(n18068), .B(n18089), .Z(n18091) );
  NOR U18407 ( .A(n95), .B(n60), .Z(n18085) );
  IV U18408 ( .A(n18085), .Z(n18071) );
  XOR U18409 ( .A(n18070), .B(n18069), .Z(n18084) );
  NOR U18410 ( .A(n18071), .B(n18084), .Z(n18087) );
  NOR U18411 ( .A(n60), .B(n93), .Z(n19097) );
  IV U18412 ( .A(n19097), .Z(n18072) );
  NOR U18413 ( .A(n59), .B(n168), .Z(n18080) );
  IV U18414 ( .A(n18080), .Z(n18075) );
  NOR U18415 ( .A(n18072), .B(n18075), .Z(n18073) );
  IV U18416 ( .A(n18073), .Z(n18074) );
  NOR U18417 ( .A(n94), .B(n18074), .Z(n18083) );
  NOR U18418 ( .A(n18075), .B(n93), .Z(n18076) );
  XOR U18419 ( .A(n94), .B(n18076), .Z(n18077) );
  NOR U18420 ( .A(n60), .B(n18077), .Z(n18078) );
  IV U18421 ( .A(n18078), .Z(n18590) );
  XOR U18422 ( .A(n18080), .B(n18079), .Z(n18589) );
  IV U18423 ( .A(n18589), .Z(n18081) );
  NOR U18424 ( .A(n18590), .B(n18081), .Z(n18082) );
  NOR U18425 ( .A(n18083), .B(n18082), .Z(n18586) );
  XOR U18426 ( .A(n18085), .B(n18084), .Z(n18585) );
  NOR U18427 ( .A(n18586), .B(n18585), .Z(n18086) );
  NOR U18428 ( .A(n18087), .B(n18086), .Z(n18613) );
  XOR U18429 ( .A(n18089), .B(n18088), .Z(n18612) );
  NOR U18430 ( .A(n18613), .B(n18612), .Z(n18090) );
  NOR U18431 ( .A(n18091), .B(n18090), .Z(n18096) );
  XOR U18432 ( .A(n18093), .B(n18092), .Z(n18095) );
  IV U18433 ( .A(n18095), .Z(n18094) );
  NOR U18434 ( .A(n18096), .B(n18094), .Z(n18099) );
  XOR U18435 ( .A(n18096), .B(n18095), .Z(n18582) );
  NOR U18436 ( .A(n97), .B(n60), .Z(n18583) );
  IV U18437 ( .A(n18583), .Z(n18097) );
  NOR U18438 ( .A(n18582), .B(n18097), .Z(n18098) );
  NOR U18439 ( .A(n18099), .B(n18098), .Z(n18578) );
  XOR U18440 ( .A(n18101), .B(n18100), .Z(n18579) );
  NOR U18441 ( .A(n18578), .B(n18579), .Z(n18102) );
  NOR U18442 ( .A(n18103), .B(n18102), .Z(n18574) );
  XOR U18443 ( .A(n18105), .B(n18104), .Z(n18575) );
  NOR U18444 ( .A(n18574), .B(n18575), .Z(n18106) );
  NOR U18445 ( .A(n18107), .B(n18106), .Z(n18570) );
  XOR U18446 ( .A(n18109), .B(n18108), .Z(n18571) );
  NOR U18447 ( .A(n18570), .B(n18571), .Z(n18110) );
  NOR U18448 ( .A(n18111), .B(n18110), .Z(n18566) );
  XOR U18449 ( .A(n18113), .B(n18112), .Z(n18567) );
  NOR U18450 ( .A(n18566), .B(n18567), .Z(n18114) );
  NOR U18451 ( .A(n18115), .B(n18114), .Z(n18562) );
  XOR U18452 ( .A(n18117), .B(n18116), .Z(n18563) );
  NOR U18453 ( .A(n18562), .B(n18563), .Z(n18118) );
  NOR U18454 ( .A(n18119), .B(n18118), .Z(n18558) );
  XOR U18455 ( .A(n18121), .B(n18120), .Z(n18559) );
  NOR U18456 ( .A(n18558), .B(n18559), .Z(n18122) );
  NOR U18457 ( .A(n18123), .B(n18122), .Z(n18554) );
  XOR U18458 ( .A(n18125), .B(n18124), .Z(n18555) );
  NOR U18459 ( .A(n18554), .B(n18555), .Z(n18126) );
  NOR U18460 ( .A(n18127), .B(n18126), .Z(n18550) );
  XOR U18461 ( .A(n18129), .B(n18128), .Z(n18551) );
  NOR U18462 ( .A(n18550), .B(n18551), .Z(n18130) );
  NOR U18463 ( .A(n18131), .B(n18130), .Z(n18657) );
  XOR U18464 ( .A(n18133), .B(n18132), .Z(n18656) );
  NOR U18465 ( .A(n18657), .B(n18656), .Z(n18134) );
  NOR U18466 ( .A(n18135), .B(n18134), .Z(n18140) );
  XOR U18467 ( .A(n18137), .B(n18136), .Z(n18139) );
  IV U18468 ( .A(n18139), .Z(n18138) );
  NOR U18469 ( .A(n18140), .B(n18138), .Z(n18143) );
  XOR U18470 ( .A(n18140), .B(n18139), .Z(n18547) );
  NOR U18471 ( .A(n104), .B(n60), .Z(n18548) );
  IV U18472 ( .A(n18548), .Z(n18141) );
  NOR U18473 ( .A(n18547), .B(n18141), .Z(n18142) );
  NOR U18474 ( .A(n18143), .B(n18142), .Z(n18543) );
  XOR U18475 ( .A(n18145), .B(n18144), .Z(n18544) );
  NOR U18476 ( .A(n18543), .B(n18544), .Z(n18146) );
  NOR U18477 ( .A(n18147), .B(n18146), .Z(n18539) );
  XOR U18478 ( .A(n18149), .B(n18148), .Z(n18540) );
  NOR U18479 ( .A(n18539), .B(n18540), .Z(n18150) );
  NOR U18480 ( .A(n18151), .B(n18150), .Z(n18535) );
  XOR U18481 ( .A(n18153), .B(n18152), .Z(n18536) );
  NOR U18482 ( .A(n18535), .B(n18536), .Z(n18154) );
  NOR U18483 ( .A(n18155), .B(n18154), .Z(n18160) );
  XOR U18484 ( .A(n18157), .B(n18156), .Z(n18159) );
  IV U18485 ( .A(n18159), .Z(n18158) );
  NOR U18486 ( .A(n18160), .B(n18158), .Z(n18163) );
  XOR U18487 ( .A(n18160), .B(n18159), .Z(n18532) );
  NOR U18488 ( .A(n107), .B(n60), .Z(n18533) );
  IV U18489 ( .A(n18533), .Z(n18161) );
  NOR U18490 ( .A(n18532), .B(n18161), .Z(n18162) );
  NOR U18491 ( .A(n18163), .B(n18162), .Z(n18528) );
  XOR U18492 ( .A(n18165), .B(n18164), .Z(n18529) );
  NOR U18493 ( .A(n18528), .B(n18529), .Z(n18166) );
  NOR U18494 ( .A(n18167), .B(n18166), .Z(n18170) );
  NOR U18495 ( .A(n108), .B(n60), .Z(n18169) );
  IV U18496 ( .A(n18169), .Z(n18168) );
  NOR U18497 ( .A(n18170), .B(n18168), .Z(n18175) );
  XOR U18498 ( .A(n18170), .B(n18169), .Z(n18525) );
  XOR U18499 ( .A(n18172), .B(n18171), .Z(n18526) );
  IV U18500 ( .A(n18526), .Z(n18173) );
  NOR U18501 ( .A(n18525), .B(n18173), .Z(n18174) );
  NOR U18502 ( .A(n18175), .B(n18174), .Z(n18521) );
  XOR U18503 ( .A(n18177), .B(n18176), .Z(n18522) );
  NOR U18504 ( .A(n18521), .B(n18522), .Z(n18178) );
  NOR U18505 ( .A(n18179), .B(n18178), .Z(n18520) );
  XOR U18506 ( .A(n18181), .B(n18180), .Z(n18519) );
  NOR U18507 ( .A(n18520), .B(n18519), .Z(n18182) );
  NOR U18508 ( .A(n18183), .B(n18182), .Z(n18184) );
  IV U18509 ( .A(n18184), .Z(n18517) );
  XOR U18510 ( .A(n18186), .B(n18185), .Z(n18187) );
  IV U18511 ( .A(n18187), .Z(n18516) );
  NOR U18512 ( .A(n18517), .B(n18516), .Z(n18188) );
  NOR U18513 ( .A(n18189), .B(n18188), .Z(n18190) );
  IV U18514 ( .A(n18190), .Z(n18515) );
  XOR U18515 ( .A(n18192), .B(n18191), .Z(n18514) );
  NOR U18516 ( .A(n18515), .B(n18514), .Z(n18193) );
  NOR U18517 ( .A(n18194), .B(n18193), .Z(n18195) );
  IV U18518 ( .A(n18195), .Z(n18511) );
  NOR U18519 ( .A(n18512), .B(n18511), .Z(n18196) );
  NOR U18520 ( .A(n18197), .B(n18196), .Z(n18198) );
  IV U18521 ( .A(n18198), .Z(n18510) );
  XOR U18522 ( .A(n18200), .B(n18199), .Z(n18509) );
  NOR U18523 ( .A(n18510), .B(n18509), .Z(n18201) );
  NOR U18524 ( .A(n18202), .B(n18201), .Z(n18203) );
  IV U18525 ( .A(n18203), .Z(n18507) );
  XOR U18526 ( .A(n18205), .B(n18204), .Z(n18206) );
  IV U18527 ( .A(n18206), .Z(n18506) );
  NOR U18528 ( .A(n18507), .B(n18506), .Z(n18207) );
  NOR U18529 ( .A(n18208), .B(n18207), .Z(n18209) );
  IV U18530 ( .A(n18209), .Z(n18505) );
  XOR U18531 ( .A(n18211), .B(n18210), .Z(n18504) );
  NOR U18532 ( .A(n18505), .B(n18504), .Z(n18212) );
  NOR U18533 ( .A(n18213), .B(n18212), .Z(n18214) );
  IV U18534 ( .A(n18214), .Z(n18502) );
  XOR U18535 ( .A(n18216), .B(n18215), .Z(n18217) );
  IV U18536 ( .A(n18217), .Z(n18501) );
  NOR U18537 ( .A(n18502), .B(n18501), .Z(n18218) );
  NOR U18538 ( .A(n18219), .B(n18218), .Z(n18220) );
  IV U18539 ( .A(n18220), .Z(n18500) );
  XOR U18540 ( .A(n18222), .B(n18221), .Z(n18499) );
  NOR U18541 ( .A(n18500), .B(n18499), .Z(n18223) );
  NOR U18542 ( .A(n18224), .B(n18223), .Z(n18497) );
  NOR U18543 ( .A(n18226), .B(n18225), .Z(n18227) );
  NOR U18544 ( .A(n18497), .B(n18227), .Z(n18228) );
  NOR U18545 ( .A(n18229), .B(n18228), .Z(n18234) );
  NOR U18546 ( .A(n115), .B(n60), .Z(n18233) );
  IV U18547 ( .A(n18233), .Z(n18230) );
  NOR U18548 ( .A(n18234), .B(n18230), .Z(n18236) );
  XOR U18549 ( .A(n18232), .B(n18231), .Z(n18493) );
  XOR U18550 ( .A(n18234), .B(n18233), .Z(n18492) );
  NOR U18551 ( .A(n18493), .B(n18492), .Z(n18235) );
  NOR U18552 ( .A(n18236), .B(n18235), .Z(n18757) );
  XOR U18553 ( .A(n18238), .B(n18237), .Z(n18758) );
  NOR U18554 ( .A(n18757), .B(n18758), .Z(n18239) );
  NOR U18555 ( .A(n18240), .B(n18239), .Z(n18490) );
  XOR U18556 ( .A(n18242), .B(n18241), .Z(n18489) );
  NOR U18557 ( .A(n18490), .B(n18489), .Z(n18243) );
  NOR U18558 ( .A(n18244), .B(n18243), .Z(n18486) );
  NOR U18559 ( .A(n18246), .B(n18245), .Z(n18247) );
  NOR U18560 ( .A(n18486), .B(n18247), .Z(n18248) );
  NOR U18561 ( .A(n18249), .B(n18248), .Z(n18255) );
  NOR U18562 ( .A(n117), .B(n60), .Z(n18256) );
  IV U18563 ( .A(n18256), .Z(n18250) );
  NOR U18564 ( .A(n18255), .B(n18250), .Z(n18258) );
  XOR U18565 ( .A(n18252), .B(n18251), .Z(n18253) );
  XOR U18566 ( .A(n18254), .B(n18253), .Z(n18482) );
  XOR U18567 ( .A(n18256), .B(n18255), .Z(n18481) );
  NOR U18568 ( .A(n18482), .B(n18481), .Z(n18257) );
  NOR U18569 ( .A(n18258), .B(n18257), .Z(n18781) );
  IV U18570 ( .A(n18781), .Z(n18259) );
  NOR U18571 ( .A(n18260), .B(n18259), .Z(n18261) );
  NOR U18572 ( .A(n18262), .B(n18261), .Z(n18268) );
  IV U18573 ( .A(n18268), .Z(n18263) );
  NOR U18574 ( .A(n18269), .B(n18263), .Z(n18271) );
  XOR U18575 ( .A(n18265), .B(n18264), .Z(n18266) );
  XOR U18576 ( .A(n18267), .B(n18266), .Z(n18479) );
  XOR U18577 ( .A(n18269), .B(n18268), .Z(n18480) );
  NOR U18578 ( .A(n18479), .B(n18480), .Z(n18270) );
  NOR U18579 ( .A(n18271), .B(n18270), .Z(n18797) );
  IV U18580 ( .A(n18797), .Z(n18272) );
  NOR U18581 ( .A(n18273), .B(n18272), .Z(n18274) );
  NOR U18582 ( .A(n18275), .B(n18274), .Z(n18281) );
  IV U18583 ( .A(n18281), .Z(n18276) );
  NOR U18584 ( .A(n18282), .B(n18276), .Z(n18284) );
  XOR U18585 ( .A(n18278), .B(n18277), .Z(n18279) );
  XOR U18586 ( .A(n18280), .B(n18279), .Z(n18475) );
  XOR U18587 ( .A(n18282), .B(n18281), .Z(n18476) );
  NOR U18588 ( .A(n18475), .B(n18476), .Z(n18283) );
  NOR U18589 ( .A(n18284), .B(n18283), .Z(n18285) );
  IV U18590 ( .A(n18285), .Z(n18809) );
  NOR U18591 ( .A(n18286), .B(n18809), .Z(n18287) );
  NOR U18592 ( .A(n18288), .B(n18287), .Z(n18289) );
  IV U18593 ( .A(n18289), .Z(n18296) );
  NOR U18594 ( .A(n126), .B(n60), .Z(n18295) );
  IV U18595 ( .A(n18295), .Z(n18290) );
  NOR U18596 ( .A(n18296), .B(n18290), .Z(n18298) );
  XOR U18597 ( .A(n18292), .B(n18291), .Z(n18293) );
  XOR U18598 ( .A(n18294), .B(n18293), .Z(n18471) );
  XOR U18599 ( .A(n18296), .B(n18295), .Z(n18472) );
  NOR U18600 ( .A(n18471), .B(n18472), .Z(n18297) );
  NOR U18601 ( .A(n18298), .B(n18297), .Z(n18824) );
  XOR U18602 ( .A(n18300), .B(n18299), .Z(n18825) );
  NOR U18603 ( .A(n18824), .B(n18825), .Z(n18301) );
  NOR U18604 ( .A(n18302), .B(n18301), .Z(n18307) );
  XOR U18605 ( .A(n18304), .B(n18303), .Z(n18306) );
  IV U18606 ( .A(n18306), .Z(n18305) );
  NOR U18607 ( .A(n18307), .B(n18305), .Z(n18310) );
  XOR U18608 ( .A(n18307), .B(n18306), .Z(n18830) );
  NOR U18609 ( .A(n131), .B(n60), .Z(n18831) );
  IV U18610 ( .A(n18831), .Z(n18308) );
  NOR U18611 ( .A(n18830), .B(n18308), .Z(n18309) );
  NOR U18612 ( .A(n18310), .B(n18309), .Z(n18837) );
  XOR U18613 ( .A(n18312), .B(n18311), .Z(n18836) );
  NOR U18614 ( .A(n18837), .B(n18836), .Z(n18313) );
  NOR U18615 ( .A(n18314), .B(n18313), .Z(n18316) );
  IV U18616 ( .A(n18316), .Z(n18465) );
  NOR U18617 ( .A(n18315), .B(n18465), .Z(n18323) );
  IV U18618 ( .A(n18315), .Z(n18466) );
  NOR U18619 ( .A(n18316), .B(n18466), .Z(n18321) );
  XOR U18620 ( .A(n18318), .B(n18317), .Z(n18319) );
  XOR U18621 ( .A(n18320), .B(n18319), .Z(n18468) );
  NOR U18622 ( .A(n18321), .B(n18468), .Z(n18322) );
  NOR U18623 ( .A(n18323), .B(n18322), .Z(n18324) );
  IV U18624 ( .A(n18324), .Z(n18331) );
  NOR U18625 ( .A(n137), .B(n60), .Z(n18330) );
  IV U18626 ( .A(n18330), .Z(n18325) );
  NOR U18627 ( .A(n18331), .B(n18325), .Z(n18333) );
  XOR U18628 ( .A(n18327), .B(n18326), .Z(n18328) );
  XOR U18629 ( .A(n18329), .B(n18328), .Z(n18464) );
  XOR U18630 ( .A(n18331), .B(n18330), .Z(n18463) );
  NOR U18631 ( .A(n18464), .B(n18463), .Z(n18332) );
  NOR U18632 ( .A(n18333), .B(n18332), .Z(n18338) );
  XOR U18633 ( .A(n18335), .B(n18334), .Z(n18337) );
  IV U18634 ( .A(n18337), .Z(n18336) );
  NOR U18635 ( .A(n18338), .B(n18336), .Z(n18341) );
  XOR U18636 ( .A(n18338), .B(n18337), .Z(n18849) );
  NOR U18637 ( .A(n139), .B(n60), .Z(n18339) );
  IV U18638 ( .A(n18339), .Z(n18848) );
  NOR U18639 ( .A(n18849), .B(n18848), .Z(n18340) );
  NOR U18640 ( .A(n18341), .B(n18340), .Z(n18345) );
  XOR U18641 ( .A(n18343), .B(n18342), .Z(n18860) );
  IV U18642 ( .A(n18860), .Z(n18344) );
  NOR U18643 ( .A(n18345), .B(n18344), .Z(n18349) );
  IV U18644 ( .A(n18345), .Z(n18857) );
  NOR U18645 ( .A(n18860), .B(n18857), .Z(n18347) );
  NOR U18646 ( .A(n141), .B(n60), .Z(n18346) );
  IV U18647 ( .A(n18346), .Z(n18858) );
  NOR U18648 ( .A(n18347), .B(n18858), .Z(n18348) );
  NOR U18649 ( .A(n18349), .B(n18348), .Z(n18354) );
  NOR U18650 ( .A(n143), .B(n60), .Z(n18353) );
  IV U18651 ( .A(n18353), .Z(n18350) );
  NOR U18652 ( .A(n18354), .B(n18350), .Z(n18357) );
  XOR U18653 ( .A(n18352), .B(n18351), .Z(n18866) );
  IV U18654 ( .A(n18866), .Z(n18355) );
  XOR U18655 ( .A(n18354), .B(n18353), .Z(n18865) );
  NOR U18656 ( .A(n18355), .B(n18865), .Z(n18356) );
  NOR U18657 ( .A(n18357), .B(n18356), .Z(n18361) );
  IV U18658 ( .A(n18361), .Z(n18459) );
  NOR U18659 ( .A(n18360), .B(n18459), .Z(n18364) );
  XOR U18660 ( .A(n18359), .B(n18358), .Z(n18462) );
  IV U18661 ( .A(n18360), .Z(n18460) );
  NOR U18662 ( .A(n18361), .B(n18460), .Z(n18362) );
  NOR U18663 ( .A(n18462), .B(n18362), .Z(n18363) );
  NOR U18664 ( .A(n18364), .B(n18363), .Z(n18368) );
  IV U18665 ( .A(n18368), .Z(n18366) );
  NOR U18666 ( .A(n147), .B(n60), .Z(n18365) );
  IV U18667 ( .A(n18365), .Z(n18367) );
  NOR U18668 ( .A(n18366), .B(n18367), .Z(n18373) );
  XOR U18669 ( .A(n18368), .B(n18367), .Z(n18883) );
  XOR U18670 ( .A(n18370), .B(n18369), .Z(n18882) );
  IV U18671 ( .A(n18882), .Z(n18371) );
  NOR U18672 ( .A(n18883), .B(n18371), .Z(n18372) );
  NOR U18673 ( .A(n18373), .B(n18372), .Z(n18376) );
  NOR U18674 ( .A(n148), .B(n60), .Z(n18375) );
  IV U18675 ( .A(n18375), .Z(n18374) );
  NOR U18676 ( .A(n18376), .B(n18374), .Z(n18380) );
  XOR U18677 ( .A(n18376), .B(n18375), .Z(n18886) );
  XOR U18678 ( .A(n18378), .B(n18377), .Z(n18887) );
  NOR U18679 ( .A(n18886), .B(n18887), .Z(n18379) );
  NOR U18680 ( .A(n18380), .B(n18379), .Z(n18385) );
  NOR U18681 ( .A(n150), .B(n60), .Z(n18384) );
  IV U18682 ( .A(n18384), .Z(n18381) );
  NOR U18683 ( .A(n18385), .B(n18381), .Z(n18387) );
  XOR U18684 ( .A(n18383), .B(n18382), .Z(n18898) );
  XOR U18685 ( .A(n18385), .B(n18384), .Z(n18897) );
  NOR U18686 ( .A(n18898), .B(n18897), .Z(n18386) );
  NOR U18687 ( .A(n18387), .B(n18386), .Z(n18391) );
  XOR U18688 ( .A(n18389), .B(n18388), .Z(n18390) );
  NOR U18689 ( .A(n18391), .B(n18390), .Z(n18395) );
  XOR U18690 ( .A(n18391), .B(n18390), .Z(n18457) );
  IV U18691 ( .A(n18457), .Z(n18393) );
  NOR U18692 ( .A(n153), .B(n60), .Z(n18392) );
  IV U18693 ( .A(n18392), .Z(n18456) );
  NOR U18694 ( .A(n18393), .B(n18456), .Z(n18394) );
  NOR U18695 ( .A(n18395), .B(n18394), .Z(n18398) );
  NOR U18696 ( .A(n155), .B(n60), .Z(n18397) );
  IV U18697 ( .A(n18397), .Z(n18396) );
  NOR U18698 ( .A(n18398), .B(n18396), .Z(n18402) );
  XOR U18699 ( .A(n18398), .B(n18397), .Z(n18910) );
  XOR U18700 ( .A(n18400), .B(n18399), .Z(n18909) );
  NOR U18701 ( .A(n18910), .B(n18909), .Z(n18401) );
  NOR U18702 ( .A(n18402), .B(n18401), .Z(n18407) );
  NOR U18703 ( .A(n156), .B(n60), .Z(n18406) );
  IV U18704 ( .A(n18406), .Z(n18403) );
  NOR U18705 ( .A(n18407), .B(n18403), .Z(n18410) );
  XOR U18706 ( .A(n18405), .B(n18404), .Z(n18915) );
  IV U18707 ( .A(n18915), .Z(n18408) );
  XOR U18708 ( .A(n18407), .B(n18406), .Z(n18914) );
  NOR U18709 ( .A(n18408), .B(n18914), .Z(n18409) );
  NOR U18710 ( .A(n18410), .B(n18409), .Z(n18414) );
  XOR U18711 ( .A(n18412), .B(n18411), .Z(n18413) );
  NOR U18712 ( .A(n18414), .B(n18413), .Z(n18418) );
  XOR U18713 ( .A(n18414), .B(n18413), .Z(n18415) );
  IV U18714 ( .A(n18415), .Z(n18926) );
  NOR U18715 ( .A(n158), .B(n60), .Z(n18925) );
  IV U18716 ( .A(n18925), .Z(n18416) );
  NOR U18717 ( .A(n18926), .B(n18416), .Z(n18417) );
  NOR U18718 ( .A(n18418), .B(n18417), .Z(n18421) );
  NOR U18719 ( .A(n161), .B(n60), .Z(n18420) );
  IV U18720 ( .A(n18420), .Z(n18419) );
  NOR U18721 ( .A(n18421), .B(n18419), .Z(n18425) );
  XOR U18722 ( .A(n18421), .B(n18420), .Z(n18933) );
  XOR U18723 ( .A(n18423), .B(n18422), .Z(n18932) );
  NOR U18724 ( .A(n18933), .B(n18932), .Z(n18424) );
  NOR U18725 ( .A(n18425), .B(n18424), .Z(n18430) );
  NOR U18726 ( .A(n163), .B(n60), .Z(n18429) );
  IV U18727 ( .A(n18429), .Z(n18426) );
  NOR U18728 ( .A(n18430), .B(n18426), .Z(n18433) );
  XOR U18729 ( .A(n18428), .B(n18427), .Z(n18938) );
  IV U18730 ( .A(n18938), .Z(n18431) );
  XOR U18731 ( .A(n18430), .B(n18429), .Z(n18937) );
  NOR U18732 ( .A(n18431), .B(n18937), .Z(n18432) );
  NOR U18733 ( .A(n18433), .B(n18432), .Z(n18437) );
  XOR U18734 ( .A(n18435), .B(n18434), .Z(n18436) );
  NOR U18735 ( .A(n18437), .B(n18436), .Z(n18441) );
  XOR U18736 ( .A(n18437), .B(n18436), .Z(n18454) );
  IV U18737 ( .A(n18454), .Z(n18439) );
  NOR U18738 ( .A(n165), .B(n60), .Z(n18438) );
  IV U18739 ( .A(n18438), .Z(n18453) );
  NOR U18740 ( .A(n18439), .B(n18453), .Z(n18440) );
  NOR U18741 ( .A(n18441), .B(n18440), .Z(n18444) );
  NOR U18742 ( .A(n167), .B(n60), .Z(n18443) );
  IV U18743 ( .A(n18443), .Z(n18442) );
  NOR U18744 ( .A(n18444), .B(n18442), .Z(n18448) );
  XOR U18745 ( .A(n18444), .B(n18443), .Z(n18949) );
  XOR U18746 ( .A(n18446), .B(n18445), .Z(n18950) );
  NOR U18747 ( .A(n18949), .B(n18950), .Z(n18447) );
  NOR U18748 ( .A(n18448), .B(n18447), .Z(n31580) );
  NOR U18749 ( .A(n18452), .B(n31580), .Z(n31578) );
  IV U18750 ( .A(n31578), .Z(n18451) );
  XOR U18751 ( .A(n18450), .B(n18449), .Z(n28556) );
  IV U18752 ( .A(n28556), .Z(n31587) );
  NOR U18753 ( .A(n18451), .B(n31587), .Z(n28563) );
  XOR U18754 ( .A(n31580), .B(n18452), .Z(n31577) );
  IV U18755 ( .A(n31577), .Z(n18952) );
  NOR U18756 ( .A(n167), .B(n61), .Z(n18946) );
  IV U18757 ( .A(n18946), .Z(n18455) );
  XOR U18758 ( .A(n18454), .B(n18453), .Z(n18945) );
  NOR U18759 ( .A(n18455), .B(n18945), .Z(n18948) );
  XOR U18760 ( .A(n18457), .B(n18456), .Z(n18902) );
  NOR U18761 ( .A(n155), .B(n61), .Z(n19873) );
  IV U18762 ( .A(n19873), .Z(n18458) );
  NOR U18763 ( .A(n18902), .B(n18458), .Z(n18905) );
  XOR U18764 ( .A(n18460), .B(n18459), .Z(n18461) );
  XOR U18765 ( .A(n18462), .B(n18461), .Z(n18874) );
  IV U18766 ( .A(n18874), .Z(n19807) );
  NOR U18767 ( .A(n141), .B(n61), .Z(n18850) );
  XOR U18768 ( .A(n18464), .B(n18463), .Z(n18955) );
  XOR U18769 ( .A(n18466), .B(n18465), .Z(n18467) );
  XOR U18770 ( .A(n18468), .B(n18467), .Z(n19341) );
  IV U18771 ( .A(n19341), .Z(n18469) );
  NOR U18772 ( .A(n137), .B(n61), .Z(n19344) );
  NOR U18773 ( .A(n18469), .B(n19344), .Z(n18847) );
  IV U18774 ( .A(n19344), .Z(n18470) );
  NOR U18775 ( .A(n19341), .B(n18470), .Z(n18845) );
  NOR U18776 ( .A(n128), .B(n61), .Z(n18473) );
  XOR U18777 ( .A(n18472), .B(n18471), .Z(n19313) );
  NOR U18778 ( .A(n18473), .B(n19313), .Z(n18819) );
  IV U18779 ( .A(n18473), .Z(n19310) );
  IV U18780 ( .A(n19313), .Z(n18474) );
  NOR U18781 ( .A(n19310), .B(n18474), .Z(n18817) );
  XOR U18782 ( .A(n18476), .B(n18475), .Z(n18477) );
  NOR U18783 ( .A(n125), .B(n61), .Z(n18478) );
  NOR U18784 ( .A(n18477), .B(n18478), .Z(n18805) );
  IV U18785 ( .A(n18477), .Z(n19297) );
  IV U18786 ( .A(n18478), .Z(n19296) );
  NOR U18787 ( .A(n19297), .B(n19296), .Z(n18803) );
  XOR U18788 ( .A(n18480), .B(n18479), .Z(n18786) );
  NOR U18789 ( .A(n120), .B(n61), .Z(n18787) );
  NOR U18790 ( .A(n18786), .B(n18787), .Z(n18791) );
  XOR U18791 ( .A(n18482), .B(n18481), .Z(n18773) );
  IV U18792 ( .A(n18773), .Z(n18970) );
  NOR U18793 ( .A(n79), .B(n61), .Z(n18772) );
  IV U18794 ( .A(n18772), .Z(n18969) );
  NOR U18795 ( .A(n18970), .B(n18969), .Z(n18776) );
  XOR U18796 ( .A(n18484), .B(n18483), .Z(n18485) );
  XOR U18797 ( .A(n18486), .B(n18485), .Z(n18769) );
  NOR U18798 ( .A(n117), .B(n61), .Z(n18768) );
  IV U18799 ( .A(n18768), .Z(n18487) );
  NOR U18800 ( .A(n18769), .B(n18487), .Z(n18771) );
  NOR U18801 ( .A(n80), .B(n61), .Z(n18488) );
  IV U18802 ( .A(n18488), .Z(n18765) );
  XOR U18803 ( .A(n18490), .B(n18489), .Z(n18764) );
  IV U18804 ( .A(n18764), .Z(n18491) );
  NOR U18805 ( .A(n18765), .B(n18491), .Z(n18767) );
  XOR U18806 ( .A(n18493), .B(n18492), .Z(n18752) );
  IV U18807 ( .A(n18752), .Z(n18981) );
  NOR U18808 ( .A(n81), .B(n61), .Z(n18751) );
  IV U18809 ( .A(n18751), .Z(n18980) );
  NOR U18810 ( .A(n18981), .B(n18980), .Z(n18755) );
  XOR U18811 ( .A(n18495), .B(n18494), .Z(n18496) );
  XOR U18812 ( .A(n18497), .B(n18496), .Z(n18748) );
  NOR U18813 ( .A(n115), .B(n61), .Z(n18747) );
  IV U18814 ( .A(n18747), .Z(n18498) );
  NOR U18815 ( .A(n18748), .B(n18498), .Z(n18750) );
  NOR U18816 ( .A(n82), .B(n61), .Z(n18742) );
  XOR U18817 ( .A(n18500), .B(n18499), .Z(n18741) );
  NOR U18818 ( .A(n18742), .B(n18741), .Z(n18745) );
  XOR U18819 ( .A(n18502), .B(n18501), .Z(n18737) );
  NOR U18820 ( .A(n114), .B(n61), .Z(n18736) );
  IV U18821 ( .A(n18736), .Z(n18503) );
  NOR U18822 ( .A(n18737), .B(n18503), .Z(n18739) );
  NOR U18823 ( .A(n83), .B(n61), .Z(n18731) );
  XOR U18824 ( .A(n18505), .B(n18504), .Z(n18730) );
  NOR U18825 ( .A(n18731), .B(n18730), .Z(n18734) );
  XOR U18826 ( .A(n18507), .B(n18506), .Z(n18726) );
  NOR U18827 ( .A(n113), .B(n61), .Z(n18725) );
  IV U18828 ( .A(n18725), .Z(n18508) );
  NOR U18829 ( .A(n18726), .B(n18508), .Z(n18728) );
  NOR U18830 ( .A(n84), .B(n61), .Z(n18720) );
  XOR U18831 ( .A(n18510), .B(n18509), .Z(n18719) );
  NOR U18832 ( .A(n18720), .B(n18719), .Z(n18723) );
  XOR U18833 ( .A(n18512), .B(n18511), .Z(n18715) );
  NOR U18834 ( .A(n112), .B(n61), .Z(n18714) );
  IV U18835 ( .A(n18714), .Z(n18513) );
  NOR U18836 ( .A(n18715), .B(n18513), .Z(n18717) );
  NOR U18837 ( .A(n85), .B(n61), .Z(n18709) );
  XOR U18838 ( .A(n18515), .B(n18514), .Z(n18708) );
  NOR U18839 ( .A(n18709), .B(n18708), .Z(n18712) );
  XOR U18840 ( .A(n18517), .B(n18516), .Z(n18704) );
  NOR U18841 ( .A(n111), .B(n61), .Z(n18703) );
  IV U18842 ( .A(n18703), .Z(n18518) );
  NOR U18843 ( .A(n18704), .B(n18518), .Z(n18706) );
  NOR U18844 ( .A(n86), .B(n61), .Z(n18698) );
  XOR U18845 ( .A(n18520), .B(n18519), .Z(n18697) );
  NOR U18846 ( .A(n18698), .B(n18697), .Z(n18701) );
  IV U18847 ( .A(n18521), .Z(n18523) );
  XOR U18848 ( .A(n18523), .B(n18522), .Z(n18692) );
  NOR U18849 ( .A(n110), .B(n61), .Z(n18693) );
  IV U18850 ( .A(n18693), .Z(n18524) );
  NOR U18851 ( .A(n18692), .B(n18524), .Z(n18695) );
  XOR U18852 ( .A(n18526), .B(n18525), .Z(n18688) );
  NOR U18853 ( .A(n109), .B(n61), .Z(n18689) );
  IV U18854 ( .A(n18689), .Z(n18527) );
  NOR U18855 ( .A(n18688), .B(n18527), .Z(n18691) );
  IV U18856 ( .A(n18528), .Z(n18530) );
  XOR U18857 ( .A(n18530), .B(n18529), .Z(n18684) );
  NOR U18858 ( .A(n108), .B(n61), .Z(n18685) );
  IV U18859 ( .A(n18685), .Z(n18531) );
  NOR U18860 ( .A(n18684), .B(n18531), .Z(n18687) );
  XOR U18861 ( .A(n18533), .B(n18532), .Z(n18680) );
  NOR U18862 ( .A(n87), .B(n61), .Z(n18681) );
  IV U18863 ( .A(n18681), .Z(n18534) );
  NOR U18864 ( .A(n18680), .B(n18534), .Z(n18683) );
  IV U18865 ( .A(n18535), .Z(n18537) );
  XOR U18866 ( .A(n18537), .B(n18536), .Z(n18676) );
  NOR U18867 ( .A(n107), .B(n61), .Z(n18677) );
  IV U18868 ( .A(n18677), .Z(n18538) );
  NOR U18869 ( .A(n18676), .B(n18538), .Z(n18679) );
  IV U18870 ( .A(n18539), .Z(n18541) );
  XOR U18871 ( .A(n18541), .B(n18540), .Z(n18672) );
  NOR U18872 ( .A(n88), .B(n61), .Z(n18673) );
  IV U18873 ( .A(n18673), .Z(n18542) );
  NOR U18874 ( .A(n18672), .B(n18542), .Z(n18675) );
  IV U18875 ( .A(n18543), .Z(n18545) );
  XOR U18876 ( .A(n18545), .B(n18544), .Z(n18668) );
  NOR U18877 ( .A(n106), .B(n61), .Z(n18669) );
  IV U18878 ( .A(n18669), .Z(n18546) );
  NOR U18879 ( .A(n18668), .B(n18546), .Z(n18671) );
  XOR U18880 ( .A(n18548), .B(n18547), .Z(n18664) );
  NOR U18881 ( .A(n105), .B(n61), .Z(n18665) );
  IV U18882 ( .A(n18665), .Z(n18549) );
  NOR U18883 ( .A(n18664), .B(n18549), .Z(n18667) );
  IV U18884 ( .A(n18550), .Z(n18552) );
  XOR U18885 ( .A(n18552), .B(n18551), .Z(n18652) );
  NOR U18886 ( .A(n89), .B(n61), .Z(n18653) );
  IV U18887 ( .A(n18653), .Z(n18553) );
  NOR U18888 ( .A(n18652), .B(n18553), .Z(n18655) );
  IV U18889 ( .A(n18554), .Z(n18556) );
  XOR U18890 ( .A(n18556), .B(n18555), .Z(n18648) );
  NOR U18891 ( .A(n103), .B(n61), .Z(n18649) );
  IV U18892 ( .A(n18649), .Z(n18557) );
  NOR U18893 ( .A(n18648), .B(n18557), .Z(n18651) );
  IV U18894 ( .A(n18558), .Z(n18560) );
  XOR U18895 ( .A(n18560), .B(n18559), .Z(n18644) );
  NOR U18896 ( .A(n90), .B(n61), .Z(n18645) );
  IV U18897 ( .A(n18645), .Z(n18561) );
  NOR U18898 ( .A(n18644), .B(n18561), .Z(n18647) );
  IV U18899 ( .A(n18562), .Z(n18564) );
  XOR U18900 ( .A(n18564), .B(n18563), .Z(n18640) );
  NOR U18901 ( .A(n102), .B(n61), .Z(n18641) );
  IV U18902 ( .A(n18641), .Z(n18565) );
  NOR U18903 ( .A(n18640), .B(n18565), .Z(n18643) );
  IV U18904 ( .A(n18566), .Z(n18568) );
  XOR U18905 ( .A(n18568), .B(n18567), .Z(n18636) );
  NOR U18906 ( .A(n101), .B(n61), .Z(n18637) );
  IV U18907 ( .A(n18637), .Z(n18569) );
  NOR U18908 ( .A(n18636), .B(n18569), .Z(n18639) );
  IV U18909 ( .A(n18570), .Z(n18572) );
  XOR U18910 ( .A(n18572), .B(n18571), .Z(n18632) );
  NOR U18911 ( .A(n100), .B(n61), .Z(n18633) );
  IV U18912 ( .A(n18633), .Z(n18573) );
  NOR U18913 ( .A(n18632), .B(n18573), .Z(n18635) );
  IV U18914 ( .A(n18574), .Z(n18576) );
  XOR U18915 ( .A(n18576), .B(n18575), .Z(n18628) );
  NOR U18916 ( .A(n99), .B(n61), .Z(n18629) );
  IV U18917 ( .A(n18629), .Z(n18577) );
  NOR U18918 ( .A(n18628), .B(n18577), .Z(n18631) );
  IV U18919 ( .A(n18578), .Z(n18580) );
  XOR U18920 ( .A(n18580), .B(n18579), .Z(n18624) );
  NOR U18921 ( .A(n98), .B(n61), .Z(n18625) );
  IV U18922 ( .A(n18625), .Z(n18581) );
  NOR U18923 ( .A(n18624), .B(n18581), .Z(n18627) );
  XOR U18924 ( .A(n18583), .B(n18582), .Z(n18620) );
  NOR U18925 ( .A(n91), .B(n61), .Z(n18621) );
  IV U18926 ( .A(n18621), .Z(n18584) );
  NOR U18927 ( .A(n18620), .B(n18584), .Z(n18623) );
  XOR U18928 ( .A(n18586), .B(n18585), .Z(n18608) );
  IV U18929 ( .A(n18608), .Z(n18588) );
  NOR U18930 ( .A(n96), .B(n61), .Z(n18587) );
  IV U18931 ( .A(n18587), .Z(n18609) );
  NOR U18932 ( .A(n18588), .B(n18609), .Z(n18611) );
  NOR U18933 ( .A(n95), .B(n61), .Z(n18605) );
  IV U18934 ( .A(n18605), .Z(n18591) );
  XOR U18935 ( .A(n18590), .B(n18589), .Z(n18604) );
  NOR U18936 ( .A(n18591), .B(n18604), .Z(n18607) );
  NOR U18937 ( .A(n93), .B(n61), .Z(n19493) );
  IV U18938 ( .A(n19493), .Z(n18592) );
  NOR U18939 ( .A(n60), .B(n168), .Z(n18600) );
  IV U18940 ( .A(n18600), .Z(n18595) );
  NOR U18941 ( .A(n18592), .B(n18595), .Z(n18593) );
  IV U18942 ( .A(n18593), .Z(n18594) );
  NOR U18943 ( .A(n94), .B(n18594), .Z(n18603) );
  NOR U18944 ( .A(n18595), .B(n93), .Z(n18596) );
  XOR U18945 ( .A(n94), .B(n18596), .Z(n18597) );
  NOR U18946 ( .A(n61), .B(n18597), .Z(n18598) );
  IV U18947 ( .A(n18598), .Z(n19088) );
  XOR U18948 ( .A(n18600), .B(n18599), .Z(n19087) );
  IV U18949 ( .A(n19087), .Z(n18601) );
  NOR U18950 ( .A(n19088), .B(n18601), .Z(n18602) );
  NOR U18951 ( .A(n18603), .B(n18602), .Z(n19084) );
  XOR U18952 ( .A(n18605), .B(n18604), .Z(n19083) );
  NOR U18953 ( .A(n19084), .B(n19083), .Z(n18606) );
  NOR U18954 ( .A(n18607), .B(n18606), .Z(n19111) );
  XOR U18955 ( .A(n18609), .B(n18608), .Z(n19110) );
  NOR U18956 ( .A(n19111), .B(n19110), .Z(n18610) );
  NOR U18957 ( .A(n18611), .B(n18610), .Z(n18616) );
  XOR U18958 ( .A(n18613), .B(n18612), .Z(n18615) );
  IV U18959 ( .A(n18615), .Z(n18614) );
  NOR U18960 ( .A(n18616), .B(n18614), .Z(n18619) );
  XOR U18961 ( .A(n18616), .B(n18615), .Z(n19080) );
  NOR U18962 ( .A(n97), .B(n61), .Z(n19081) );
  IV U18963 ( .A(n19081), .Z(n18617) );
  NOR U18964 ( .A(n19080), .B(n18617), .Z(n18618) );
  NOR U18965 ( .A(n18619), .B(n18618), .Z(n19076) );
  XOR U18966 ( .A(n18621), .B(n18620), .Z(n19077) );
  NOR U18967 ( .A(n19076), .B(n19077), .Z(n18622) );
  NOR U18968 ( .A(n18623), .B(n18622), .Z(n19072) );
  XOR U18969 ( .A(n18625), .B(n18624), .Z(n19073) );
  NOR U18970 ( .A(n19072), .B(n19073), .Z(n18626) );
  NOR U18971 ( .A(n18627), .B(n18626), .Z(n19068) );
  XOR U18972 ( .A(n18629), .B(n18628), .Z(n19069) );
  NOR U18973 ( .A(n19068), .B(n19069), .Z(n18630) );
  NOR U18974 ( .A(n18631), .B(n18630), .Z(n19064) );
  XOR U18975 ( .A(n18633), .B(n18632), .Z(n19065) );
  NOR U18976 ( .A(n19064), .B(n19065), .Z(n18634) );
  NOR U18977 ( .A(n18635), .B(n18634), .Z(n19060) );
  XOR U18978 ( .A(n18637), .B(n18636), .Z(n19061) );
  NOR U18979 ( .A(n19060), .B(n19061), .Z(n18638) );
  NOR U18980 ( .A(n18639), .B(n18638), .Z(n19056) );
  XOR U18981 ( .A(n18641), .B(n18640), .Z(n19057) );
  NOR U18982 ( .A(n19056), .B(n19057), .Z(n18642) );
  NOR U18983 ( .A(n18643), .B(n18642), .Z(n19052) );
  XOR U18984 ( .A(n18645), .B(n18644), .Z(n19053) );
  NOR U18985 ( .A(n19052), .B(n19053), .Z(n18646) );
  NOR U18986 ( .A(n18647), .B(n18646), .Z(n19049) );
  XOR U18987 ( .A(n18649), .B(n18648), .Z(n19048) );
  NOR U18988 ( .A(n19049), .B(n19048), .Z(n18650) );
  NOR U18989 ( .A(n18651), .B(n18650), .Z(n19044) );
  XOR U18990 ( .A(n18653), .B(n18652), .Z(n19045) );
  NOR U18991 ( .A(n19044), .B(n19045), .Z(n18654) );
  NOR U18992 ( .A(n18655), .B(n18654), .Z(n18660) );
  XOR U18993 ( .A(n18657), .B(n18656), .Z(n18659) );
  IV U18994 ( .A(n18659), .Z(n18658) );
  NOR U18995 ( .A(n18660), .B(n18658), .Z(n18663) );
  XOR U18996 ( .A(n18660), .B(n18659), .Z(n19041) );
  NOR U18997 ( .A(n104), .B(n61), .Z(n19042) );
  IV U18998 ( .A(n19042), .Z(n18661) );
  NOR U18999 ( .A(n19041), .B(n18661), .Z(n18662) );
  NOR U19000 ( .A(n18663), .B(n18662), .Z(n19037) );
  XOR U19001 ( .A(n18665), .B(n18664), .Z(n19038) );
  NOR U19002 ( .A(n19037), .B(n19038), .Z(n18666) );
  NOR U19003 ( .A(n18667), .B(n18666), .Z(n19033) );
  XOR U19004 ( .A(n18669), .B(n18668), .Z(n19034) );
  NOR U19005 ( .A(n19033), .B(n19034), .Z(n18670) );
  NOR U19006 ( .A(n18671), .B(n18670), .Z(n19029) );
  XOR U19007 ( .A(n18673), .B(n18672), .Z(n19030) );
  NOR U19008 ( .A(n19029), .B(n19030), .Z(n18674) );
  NOR U19009 ( .A(n18675), .B(n18674), .Z(n19025) );
  XOR U19010 ( .A(n18677), .B(n18676), .Z(n19026) );
  NOR U19011 ( .A(n19025), .B(n19026), .Z(n18678) );
  NOR U19012 ( .A(n18679), .B(n18678), .Z(n19179) );
  XOR U19013 ( .A(n18681), .B(n18680), .Z(n19178) );
  NOR U19014 ( .A(n19179), .B(n19178), .Z(n18682) );
  NOR U19015 ( .A(n18683), .B(n18682), .Z(n19021) );
  XOR U19016 ( .A(n18685), .B(n18684), .Z(n19022) );
  NOR U19017 ( .A(n19021), .B(n19022), .Z(n18686) );
  NOR U19018 ( .A(n18687), .B(n18686), .Z(n19017) );
  XOR U19019 ( .A(n18689), .B(n18688), .Z(n19018) );
  NOR U19020 ( .A(n19017), .B(n19018), .Z(n18690) );
  NOR U19021 ( .A(n18691), .B(n18690), .Z(n19013) );
  XOR U19022 ( .A(n18693), .B(n18692), .Z(n19014) );
  NOR U19023 ( .A(n19013), .B(n19014), .Z(n18694) );
  NOR U19024 ( .A(n18695), .B(n18694), .Z(n18696) );
  IV U19025 ( .A(n18696), .Z(n19011) );
  XOR U19026 ( .A(n18698), .B(n18697), .Z(n18699) );
  IV U19027 ( .A(n18699), .Z(n19010) );
  NOR U19028 ( .A(n19011), .B(n19010), .Z(n18700) );
  NOR U19029 ( .A(n18701), .B(n18700), .Z(n18702) );
  IV U19030 ( .A(n18702), .Z(n19009) );
  XOR U19031 ( .A(n18704), .B(n18703), .Z(n19008) );
  NOR U19032 ( .A(n19009), .B(n19008), .Z(n18705) );
  NOR U19033 ( .A(n18706), .B(n18705), .Z(n18707) );
  IV U19034 ( .A(n18707), .Z(n19006) );
  XOR U19035 ( .A(n18709), .B(n18708), .Z(n18710) );
  IV U19036 ( .A(n18710), .Z(n19005) );
  NOR U19037 ( .A(n19006), .B(n19005), .Z(n18711) );
  NOR U19038 ( .A(n18712), .B(n18711), .Z(n18713) );
  IV U19039 ( .A(n18713), .Z(n19001) );
  XOR U19040 ( .A(n18715), .B(n18714), .Z(n19000) );
  NOR U19041 ( .A(n19001), .B(n19000), .Z(n18716) );
  NOR U19042 ( .A(n18717), .B(n18716), .Z(n18718) );
  IV U19043 ( .A(n18718), .Z(n18998) );
  XOR U19044 ( .A(n18720), .B(n18719), .Z(n18721) );
  IV U19045 ( .A(n18721), .Z(n18997) );
  NOR U19046 ( .A(n18998), .B(n18997), .Z(n18722) );
  NOR U19047 ( .A(n18723), .B(n18722), .Z(n18724) );
  IV U19048 ( .A(n18724), .Z(n18996) );
  XOR U19049 ( .A(n18726), .B(n18725), .Z(n18995) );
  NOR U19050 ( .A(n18996), .B(n18995), .Z(n18727) );
  NOR U19051 ( .A(n18728), .B(n18727), .Z(n18729) );
  IV U19052 ( .A(n18729), .Z(n18993) );
  XOR U19053 ( .A(n18731), .B(n18730), .Z(n18732) );
  IV U19054 ( .A(n18732), .Z(n18992) );
  NOR U19055 ( .A(n18993), .B(n18992), .Z(n18733) );
  NOR U19056 ( .A(n18734), .B(n18733), .Z(n18735) );
  IV U19057 ( .A(n18735), .Z(n18991) );
  XOR U19058 ( .A(n18737), .B(n18736), .Z(n18990) );
  NOR U19059 ( .A(n18991), .B(n18990), .Z(n18738) );
  NOR U19060 ( .A(n18739), .B(n18738), .Z(n18740) );
  IV U19061 ( .A(n18740), .Z(n18988) );
  XOR U19062 ( .A(n18742), .B(n18741), .Z(n18743) );
  IV U19063 ( .A(n18743), .Z(n18987) );
  NOR U19064 ( .A(n18988), .B(n18987), .Z(n18744) );
  NOR U19065 ( .A(n18745), .B(n18744), .Z(n18746) );
  IV U19066 ( .A(n18746), .Z(n18986) );
  XOR U19067 ( .A(n18748), .B(n18747), .Z(n18985) );
  NOR U19068 ( .A(n18986), .B(n18985), .Z(n18749) );
  NOR U19069 ( .A(n18750), .B(n18749), .Z(n18983) );
  NOR U19070 ( .A(n18752), .B(n18751), .Z(n18753) );
  NOR U19071 ( .A(n18983), .B(n18753), .Z(n18754) );
  NOR U19072 ( .A(n18755), .B(n18754), .Z(n18761) );
  NOR U19073 ( .A(n116), .B(n61), .Z(n18760) );
  IV U19074 ( .A(n18760), .Z(n18756) );
  NOR U19075 ( .A(n18761), .B(n18756), .Z(n18763) );
  XOR U19076 ( .A(n18758), .B(n18757), .Z(n18759) );
  IV U19077 ( .A(n18759), .Z(n18977) );
  XOR U19078 ( .A(n18761), .B(n18760), .Z(n18976) );
  NOR U19079 ( .A(n18977), .B(n18976), .Z(n18762) );
  NOR U19080 ( .A(n18763), .B(n18762), .Z(n19261) );
  XOR U19081 ( .A(n18765), .B(n18764), .Z(n19260) );
  NOR U19082 ( .A(n19261), .B(n19260), .Z(n18766) );
  NOR U19083 ( .A(n18767), .B(n18766), .Z(n18975) );
  XOR U19084 ( .A(n18769), .B(n18768), .Z(n18974) );
  NOR U19085 ( .A(n18975), .B(n18974), .Z(n18770) );
  NOR U19086 ( .A(n18771), .B(n18770), .Z(n18972) );
  NOR U19087 ( .A(n18773), .B(n18772), .Z(n18774) );
  NOR U19088 ( .A(n18972), .B(n18774), .Z(n18775) );
  NOR U19089 ( .A(n18776), .B(n18775), .Z(n18782) );
  NOR U19090 ( .A(n119), .B(n61), .Z(n18783) );
  IV U19091 ( .A(n18783), .Z(n18777) );
  NOR U19092 ( .A(n18782), .B(n18777), .Z(n18785) );
  XOR U19093 ( .A(n18779), .B(n18778), .Z(n18780) );
  XOR U19094 ( .A(n18781), .B(n18780), .Z(n18966) );
  XOR U19095 ( .A(n18783), .B(n18782), .Z(n18965) );
  NOR U19096 ( .A(n18966), .B(n18965), .Z(n18784) );
  NOR U19097 ( .A(n18785), .B(n18784), .Z(n19285) );
  IV U19098 ( .A(n19285), .Z(n18789) );
  IV U19099 ( .A(n18786), .Z(n19283) );
  IV U19100 ( .A(n18787), .Z(n19282) );
  NOR U19101 ( .A(n19283), .B(n19282), .Z(n18788) );
  NOR U19102 ( .A(n18789), .B(n18788), .Z(n18790) );
  NOR U19103 ( .A(n18791), .B(n18790), .Z(n18799) );
  IV U19104 ( .A(n18799), .Z(n18793) );
  NOR U19105 ( .A(n123), .B(n61), .Z(n18792) );
  IV U19106 ( .A(n18792), .Z(n18798) );
  NOR U19107 ( .A(n18793), .B(n18798), .Z(n18801) );
  XOR U19108 ( .A(n18795), .B(n18794), .Z(n18796) );
  XOR U19109 ( .A(n18797), .B(n18796), .Z(n18964) );
  XOR U19110 ( .A(n18799), .B(n18798), .Z(n18963) );
  NOR U19111 ( .A(n18964), .B(n18963), .Z(n18800) );
  NOR U19112 ( .A(n18801), .B(n18800), .Z(n19299) );
  IV U19113 ( .A(n19299), .Z(n18802) );
  NOR U19114 ( .A(n18803), .B(n18802), .Z(n18804) );
  NOR U19115 ( .A(n18805), .B(n18804), .Z(n18806) );
  IV U19116 ( .A(n18806), .Z(n18813) );
  NOR U19117 ( .A(n126), .B(n61), .Z(n18812) );
  IV U19118 ( .A(n18812), .Z(n18807) );
  NOR U19119 ( .A(n18813), .B(n18807), .Z(n18815) );
  XOR U19120 ( .A(n18809), .B(n18808), .Z(n18810) );
  XOR U19121 ( .A(n18811), .B(n18810), .Z(n18959) );
  XOR U19122 ( .A(n18813), .B(n18812), .Z(n18960) );
  NOR U19123 ( .A(n18959), .B(n18960), .Z(n18814) );
  NOR U19124 ( .A(n18815), .B(n18814), .Z(n18816) );
  IV U19125 ( .A(n18816), .Z(n19311) );
  NOR U19126 ( .A(n18817), .B(n19311), .Z(n18818) );
  NOR U19127 ( .A(n18819), .B(n18818), .Z(n18823) );
  IV U19128 ( .A(n18823), .Z(n18821) );
  NOR U19129 ( .A(n131), .B(n61), .Z(n18820) );
  IV U19130 ( .A(n18820), .Z(n18822) );
  NOR U19131 ( .A(n18821), .B(n18822), .Z(n18828) );
  XOR U19132 ( .A(n18823), .B(n18822), .Z(n19322) );
  XOR U19133 ( .A(n18825), .B(n18824), .Z(n19321) );
  IV U19134 ( .A(n19321), .Z(n18826) );
  NOR U19135 ( .A(n19322), .B(n18826), .Z(n18827) );
  NOR U19136 ( .A(n18828), .B(n18827), .Z(n18833) );
  NOR U19137 ( .A(n133), .B(n61), .Z(n18832) );
  IV U19138 ( .A(n18832), .Z(n18829) );
  NOR U19139 ( .A(n18833), .B(n18829), .Z(n18835) );
  XOR U19140 ( .A(n18831), .B(n18830), .Z(n19326) );
  XOR U19141 ( .A(n18833), .B(n18832), .Z(n19325) );
  NOR U19142 ( .A(n19326), .B(n19325), .Z(n18834) );
  NOR U19143 ( .A(n18835), .B(n18834), .Z(n18840) );
  XOR U19144 ( .A(n18837), .B(n18836), .Z(n18839) );
  IV U19145 ( .A(n18839), .Z(n18838) );
  NOR U19146 ( .A(n18840), .B(n18838), .Z(n18843) );
  XOR U19147 ( .A(n18840), .B(n18839), .Z(n19336) );
  NOR U19148 ( .A(n135), .B(n61), .Z(n19337) );
  IV U19149 ( .A(n19337), .Z(n18841) );
  NOR U19150 ( .A(n19336), .B(n18841), .Z(n18842) );
  NOR U19151 ( .A(n18843), .B(n18842), .Z(n18844) );
  IV U19152 ( .A(n18844), .Z(n19342) );
  NOR U19153 ( .A(n18845), .B(n19342), .Z(n18846) );
  NOR U19154 ( .A(n18847), .B(n18846), .Z(n18958) );
  NOR U19155 ( .A(n139), .B(n61), .Z(n18956) );
  NOR U19156 ( .A(n18850), .B(n18851), .Z(n18854) );
  XOR U19157 ( .A(n18849), .B(n18848), .Z(n19765) );
  IV U19158 ( .A(n18850), .Z(n19763) );
  IV U19159 ( .A(n18851), .Z(n19762) );
  NOR U19160 ( .A(n19763), .B(n19762), .Z(n18852) );
  NOR U19161 ( .A(n19765), .B(n18852), .Z(n18853) );
  NOR U19162 ( .A(n18854), .B(n18853), .Z(n18862) );
  IV U19163 ( .A(n18862), .Z(n18856) );
  NOR U19164 ( .A(n143), .B(n61), .Z(n18855) );
  IV U19165 ( .A(n18855), .Z(n18861) );
  NOR U19166 ( .A(n18856), .B(n18861), .Z(n18864) );
  XOR U19167 ( .A(n18858), .B(n18857), .Z(n18859) );
  XOR U19168 ( .A(n18860), .B(n18859), .Z(n19781) );
  XOR U19169 ( .A(n18862), .B(n18861), .Z(n19782) );
  NOR U19170 ( .A(n19781), .B(n19782), .Z(n18863) );
  NOR U19171 ( .A(n18864), .B(n18863), .Z(n18868) );
  XOR U19172 ( .A(n18866), .B(n18865), .Z(n18867) );
  NOR U19173 ( .A(n18868), .B(n18867), .Z(n18872) );
  XOR U19174 ( .A(n18868), .B(n18867), .Z(n18869) );
  IV U19175 ( .A(n18869), .Z(n19790) );
  NOR U19176 ( .A(n145), .B(n61), .Z(n19791) );
  IV U19177 ( .A(n19791), .Z(n18870) );
  NOR U19178 ( .A(n19790), .B(n18870), .Z(n18871) );
  NOR U19179 ( .A(n18872), .B(n18871), .Z(n19810) );
  IV U19180 ( .A(n19810), .Z(n18873) );
  NOR U19181 ( .A(n19807), .B(n18873), .Z(n18877) );
  NOR U19182 ( .A(n147), .B(n61), .Z(n19808) );
  NOR U19183 ( .A(n19810), .B(n18874), .Z(n18875) );
  NOR U19184 ( .A(n19808), .B(n18875), .Z(n18876) );
  NOR U19185 ( .A(n18877), .B(n18876), .Z(n18878) );
  IV U19186 ( .A(n18878), .Z(n18881) );
  NOR U19187 ( .A(n148), .B(n61), .Z(n18880) );
  IV U19188 ( .A(n18880), .Z(n18879) );
  NOR U19189 ( .A(n18881), .B(n18879), .Z(n18885) );
  XOR U19190 ( .A(n18881), .B(n18880), .Z(n19828) );
  XOR U19191 ( .A(n18883), .B(n18882), .Z(n19829) );
  NOR U19192 ( .A(n19828), .B(n19829), .Z(n18884) );
  NOR U19193 ( .A(n18885), .B(n18884), .Z(n18889) );
  XOR U19194 ( .A(n18887), .B(n18886), .Z(n19850) );
  IV U19195 ( .A(n19850), .Z(n18888) );
  NOR U19196 ( .A(n18889), .B(n18888), .Z(n18893) );
  IV U19197 ( .A(n18889), .Z(n19847) );
  NOR U19198 ( .A(n19850), .B(n19847), .Z(n18891) );
  NOR U19199 ( .A(n150), .B(n61), .Z(n18890) );
  IV U19200 ( .A(n18890), .Z(n19848) );
  NOR U19201 ( .A(n18891), .B(n19848), .Z(n18892) );
  NOR U19202 ( .A(n18893), .B(n18892), .Z(n18896) );
  NOR U19203 ( .A(n153), .B(n61), .Z(n18895) );
  IV U19204 ( .A(n18895), .Z(n18894) );
  NOR U19205 ( .A(n18896), .B(n18894), .Z(n18901) );
  XOR U19206 ( .A(n18896), .B(n18895), .Z(n19861) );
  XOR U19207 ( .A(n18898), .B(n18897), .Z(n19862) );
  IV U19208 ( .A(n19862), .Z(n18899) );
  NOR U19209 ( .A(n19861), .B(n18899), .Z(n18900) );
  NOR U19210 ( .A(n18901), .B(n18900), .Z(n19871) );
  IV U19211 ( .A(n18902), .Z(n19870) );
  NOR U19212 ( .A(n19870), .B(n19873), .Z(n18903) );
  NOR U19213 ( .A(n19871), .B(n18903), .Z(n18904) );
  NOR U19214 ( .A(n18905), .B(n18904), .Z(n18908) );
  NOR U19215 ( .A(n156), .B(n61), .Z(n18907) );
  IV U19216 ( .A(n18907), .Z(n18906) );
  NOR U19217 ( .A(n18908), .B(n18906), .Z(n18913) );
  XOR U19218 ( .A(n18908), .B(n18907), .Z(n19897) );
  XOR U19219 ( .A(n18910), .B(n18909), .Z(n19898) );
  IV U19220 ( .A(n19898), .Z(n18911) );
  NOR U19221 ( .A(n19897), .B(n18911), .Z(n18912) );
  NOR U19222 ( .A(n18913), .B(n18912), .Z(n18917) );
  XOR U19223 ( .A(n18915), .B(n18914), .Z(n18916) );
  NOR U19224 ( .A(n18917), .B(n18916), .Z(n18921) );
  XOR U19225 ( .A(n18917), .B(n18916), .Z(n19909) );
  IV U19226 ( .A(n19909), .Z(n18919) );
  NOR U19227 ( .A(n158), .B(n61), .Z(n18918) );
  IV U19228 ( .A(n18918), .Z(n19910) );
  NOR U19229 ( .A(n18919), .B(n19910), .Z(n18920) );
  NOR U19230 ( .A(n18921), .B(n18920), .Z(n18924) );
  NOR U19231 ( .A(n161), .B(n61), .Z(n18923) );
  IV U19232 ( .A(n18923), .Z(n18922) );
  NOR U19233 ( .A(n18924), .B(n18922), .Z(n18928) );
  XOR U19234 ( .A(n18924), .B(n18923), .Z(n19916) );
  XOR U19235 ( .A(n18926), .B(n18925), .Z(n19917) );
  NOR U19236 ( .A(n19916), .B(n19917), .Z(n18927) );
  NOR U19237 ( .A(n18928), .B(n18927), .Z(n18931) );
  NOR U19238 ( .A(n163), .B(n61), .Z(n18930) );
  IV U19239 ( .A(n18930), .Z(n18929) );
  NOR U19240 ( .A(n18931), .B(n18929), .Z(n18936) );
  XOR U19241 ( .A(n18931), .B(n18930), .Z(n19942) );
  XOR U19242 ( .A(n18933), .B(n18932), .Z(n19943) );
  IV U19243 ( .A(n19943), .Z(n18934) );
  NOR U19244 ( .A(n19942), .B(n18934), .Z(n18935) );
  NOR U19245 ( .A(n18936), .B(n18935), .Z(n18939) );
  XOR U19246 ( .A(n18938), .B(n18937), .Z(n18940) );
  NOR U19247 ( .A(n18939), .B(n18940), .Z(n18944) );
  IV U19248 ( .A(n18939), .Z(n18941) );
  XOR U19249 ( .A(n18941), .B(n18940), .Z(n19947) );
  NOR U19250 ( .A(n165), .B(n61), .Z(n19948) );
  IV U19251 ( .A(n19948), .Z(n18942) );
  NOR U19252 ( .A(n19947), .B(n18942), .Z(n18943) );
  NOR U19253 ( .A(n18944), .B(n18943), .Z(n19966) );
  XOR U19254 ( .A(n18946), .B(n18945), .Z(n19965) );
  NOR U19255 ( .A(n19966), .B(n19965), .Z(n18947) );
  NOR U19256 ( .A(n18948), .B(n18947), .Z(n18954) );
  XOR U19257 ( .A(n18950), .B(n18949), .Z(n18951) );
  IV U19258 ( .A(n18951), .Z(n18953) );
  NOR U19259 ( .A(n18954), .B(n18953), .Z(n31570) );
  IV U19260 ( .A(n31570), .Z(n31571) );
  NOR U19261 ( .A(n18952), .B(n31571), .Z(n19976) );
  XOR U19262 ( .A(n18954), .B(n18953), .Z(n31563) );
  IV U19263 ( .A(n31563), .Z(n19972) );
  XOR U19264 ( .A(n18956), .B(n18955), .Z(n18957) );
  XOR U19265 ( .A(n18958), .B(n18957), .Z(n19757) );
  NOR U19266 ( .A(n141), .B(n62), .Z(n19754) );
  IV U19267 ( .A(n19754), .Z(n19755) );
  NOR U19268 ( .A(n128), .B(n62), .Z(n18961) );
  XOR U19269 ( .A(n18960), .B(n18959), .Z(n18962) );
  NOR U19270 ( .A(n18961), .B(n18962), .Z(n19307) );
  IV U19271 ( .A(n18961), .Z(n19706) );
  IV U19272 ( .A(n18962), .Z(n19705) );
  NOR U19273 ( .A(n19706), .B(n19705), .Z(n19305) );
  NOR U19274 ( .A(n125), .B(n62), .Z(n19291) );
  IV U19275 ( .A(n19291), .Z(n19692) );
  XOR U19276 ( .A(n18964), .B(n18963), .Z(n19290) );
  IV U19277 ( .A(n19290), .Z(n19691) );
  NOR U19278 ( .A(n19692), .B(n19691), .Z(n19294) );
  NOR U19279 ( .A(n123), .B(n62), .Z(n19287) );
  IV U19280 ( .A(n19287), .Z(n19281) );
  XOR U19281 ( .A(n18966), .B(n18965), .Z(n18967) );
  NOR U19282 ( .A(n120), .B(n62), .Z(n18968) );
  NOR U19283 ( .A(n18967), .B(n18968), .Z(n19279) );
  IV U19284 ( .A(n18967), .Z(n19363) );
  IV U19285 ( .A(n18968), .Z(n19362) );
  NOR U19286 ( .A(n19363), .B(n19362), .Z(n19277) );
  XOR U19287 ( .A(n18970), .B(n18969), .Z(n18971) );
  XOR U19288 ( .A(n18972), .B(n18971), .Z(n19273) );
  NOR U19289 ( .A(n119), .B(n62), .Z(n19272) );
  IV U19290 ( .A(n19272), .Z(n18973) );
  NOR U19291 ( .A(n19273), .B(n18973), .Z(n19275) );
  NOR U19292 ( .A(n79), .B(n62), .Z(n19268) );
  IV U19293 ( .A(n19268), .Z(n19671) );
  XOR U19294 ( .A(n18975), .B(n18974), .Z(n19267) );
  IV U19295 ( .A(n19267), .Z(n19670) );
  NOR U19296 ( .A(n19671), .B(n19670), .Z(n19271) );
  NOR U19297 ( .A(n80), .B(n62), .Z(n18978) );
  XOR U19298 ( .A(n18977), .B(n18976), .Z(n18979) );
  NOR U19299 ( .A(n18978), .B(n18979), .Z(n19257) );
  IV U19300 ( .A(n18978), .Z(n19374) );
  IV U19301 ( .A(n18979), .Z(n19373) );
  NOR U19302 ( .A(n19374), .B(n19373), .Z(n19255) );
  XOR U19303 ( .A(n18981), .B(n18980), .Z(n18982) );
  XOR U19304 ( .A(n18983), .B(n18982), .Z(n19251) );
  NOR U19305 ( .A(n116), .B(n62), .Z(n19250) );
  IV U19306 ( .A(n19250), .Z(n18984) );
  NOR U19307 ( .A(n19251), .B(n18984), .Z(n19253) );
  NOR U19308 ( .A(n81), .B(n62), .Z(n19245) );
  XOR U19309 ( .A(n18986), .B(n18985), .Z(n19244) );
  NOR U19310 ( .A(n19245), .B(n19244), .Z(n19248) );
  XOR U19311 ( .A(n18988), .B(n18987), .Z(n19240) );
  NOR U19312 ( .A(n115), .B(n62), .Z(n19239) );
  IV U19313 ( .A(n19239), .Z(n18989) );
  NOR U19314 ( .A(n19240), .B(n18989), .Z(n19242) );
  NOR U19315 ( .A(n82), .B(n62), .Z(n19234) );
  XOR U19316 ( .A(n18991), .B(n18990), .Z(n19233) );
  NOR U19317 ( .A(n19234), .B(n19233), .Z(n19237) );
  XOR U19318 ( .A(n18993), .B(n18992), .Z(n19229) );
  NOR U19319 ( .A(n114), .B(n62), .Z(n19228) );
  IV U19320 ( .A(n19228), .Z(n18994) );
  NOR U19321 ( .A(n19229), .B(n18994), .Z(n19231) );
  NOR U19322 ( .A(n83), .B(n62), .Z(n19223) );
  XOR U19323 ( .A(n18996), .B(n18995), .Z(n19222) );
  NOR U19324 ( .A(n19223), .B(n19222), .Z(n19226) );
  XOR U19325 ( .A(n18998), .B(n18997), .Z(n19218) );
  NOR U19326 ( .A(n113), .B(n62), .Z(n19217) );
  IV U19327 ( .A(n19217), .Z(n18999) );
  NOR U19328 ( .A(n19218), .B(n18999), .Z(n19220) );
  NOR U19329 ( .A(n84), .B(n62), .Z(n19003) );
  XOR U19330 ( .A(n19001), .B(n19000), .Z(n19002) );
  NOR U19331 ( .A(n19003), .B(n19002), .Z(n19215) );
  XOR U19332 ( .A(n19003), .B(n19002), .Z(n19004) );
  IV U19333 ( .A(n19004), .Z(n19396) );
  XOR U19334 ( .A(n19006), .B(n19005), .Z(n19210) );
  NOR U19335 ( .A(n112), .B(n62), .Z(n19209) );
  IV U19336 ( .A(n19209), .Z(n19007) );
  NOR U19337 ( .A(n19210), .B(n19007), .Z(n19212) );
  NOR U19338 ( .A(n85), .B(n62), .Z(n19204) );
  XOR U19339 ( .A(n19009), .B(n19008), .Z(n19203) );
  NOR U19340 ( .A(n19204), .B(n19203), .Z(n19207) );
  XOR U19341 ( .A(n19011), .B(n19010), .Z(n19199) );
  NOR U19342 ( .A(n111), .B(n62), .Z(n19198) );
  IV U19343 ( .A(n19198), .Z(n19012) );
  NOR U19344 ( .A(n19199), .B(n19012), .Z(n19201) );
  IV U19345 ( .A(n19013), .Z(n19015) );
  XOR U19346 ( .A(n19015), .B(n19014), .Z(n19194) );
  NOR U19347 ( .A(n86), .B(n62), .Z(n19195) );
  IV U19348 ( .A(n19195), .Z(n19016) );
  NOR U19349 ( .A(n19194), .B(n19016), .Z(n19197) );
  IV U19350 ( .A(n19017), .Z(n19019) );
  XOR U19351 ( .A(n19019), .B(n19018), .Z(n19190) );
  NOR U19352 ( .A(n110), .B(n62), .Z(n19191) );
  IV U19353 ( .A(n19191), .Z(n19020) );
  NOR U19354 ( .A(n19190), .B(n19020), .Z(n19193) );
  IV U19355 ( .A(n19021), .Z(n19023) );
  XOR U19356 ( .A(n19023), .B(n19022), .Z(n19186) );
  NOR U19357 ( .A(n109), .B(n62), .Z(n19187) );
  IV U19358 ( .A(n19187), .Z(n19024) );
  NOR U19359 ( .A(n19186), .B(n19024), .Z(n19189) );
  IV U19360 ( .A(n19025), .Z(n19027) );
  XOR U19361 ( .A(n19027), .B(n19026), .Z(n19174) );
  NOR U19362 ( .A(n87), .B(n62), .Z(n19175) );
  IV U19363 ( .A(n19175), .Z(n19028) );
  NOR U19364 ( .A(n19174), .B(n19028), .Z(n19177) );
  IV U19365 ( .A(n19029), .Z(n19031) );
  XOR U19366 ( .A(n19031), .B(n19030), .Z(n19170) );
  NOR U19367 ( .A(n107), .B(n62), .Z(n19171) );
  IV U19368 ( .A(n19171), .Z(n19032) );
  NOR U19369 ( .A(n19170), .B(n19032), .Z(n19173) );
  IV U19370 ( .A(n19033), .Z(n19035) );
  XOR U19371 ( .A(n19035), .B(n19034), .Z(n19166) );
  NOR U19372 ( .A(n88), .B(n62), .Z(n19167) );
  IV U19373 ( .A(n19167), .Z(n19036) );
  NOR U19374 ( .A(n19166), .B(n19036), .Z(n19169) );
  IV U19375 ( .A(n19037), .Z(n19039) );
  XOR U19376 ( .A(n19039), .B(n19038), .Z(n19162) );
  NOR U19377 ( .A(n106), .B(n62), .Z(n19163) );
  IV U19378 ( .A(n19163), .Z(n19040) );
  NOR U19379 ( .A(n19162), .B(n19040), .Z(n19165) );
  XOR U19380 ( .A(n19042), .B(n19041), .Z(n19158) );
  NOR U19381 ( .A(n105), .B(n62), .Z(n19159) );
  IV U19382 ( .A(n19159), .Z(n19043) );
  NOR U19383 ( .A(n19158), .B(n19043), .Z(n19161) );
  IV U19384 ( .A(n19044), .Z(n19046) );
  XOR U19385 ( .A(n19046), .B(n19045), .Z(n19154) );
  NOR U19386 ( .A(n104), .B(n62), .Z(n19155) );
  IV U19387 ( .A(n19155), .Z(n19047) );
  NOR U19388 ( .A(n19154), .B(n19047), .Z(n19157) );
  XOR U19389 ( .A(n19049), .B(n19048), .Z(n19150) );
  IV U19390 ( .A(n19150), .Z(n19051) );
  NOR U19391 ( .A(n89), .B(n62), .Z(n19050) );
  IV U19392 ( .A(n19050), .Z(n19151) );
  NOR U19393 ( .A(n19051), .B(n19151), .Z(n19153) );
  IV U19394 ( .A(n19052), .Z(n19054) );
  XOR U19395 ( .A(n19054), .B(n19053), .Z(n19146) );
  NOR U19396 ( .A(n103), .B(n62), .Z(n19147) );
  IV U19397 ( .A(n19147), .Z(n19055) );
  NOR U19398 ( .A(n19146), .B(n19055), .Z(n19149) );
  IV U19399 ( .A(n19056), .Z(n19058) );
  XOR U19400 ( .A(n19058), .B(n19057), .Z(n19142) );
  NOR U19401 ( .A(n90), .B(n62), .Z(n19143) );
  IV U19402 ( .A(n19143), .Z(n19059) );
  NOR U19403 ( .A(n19142), .B(n19059), .Z(n19145) );
  IV U19404 ( .A(n19060), .Z(n19062) );
  XOR U19405 ( .A(n19062), .B(n19061), .Z(n19138) );
  NOR U19406 ( .A(n102), .B(n62), .Z(n19139) );
  IV U19407 ( .A(n19139), .Z(n19063) );
  NOR U19408 ( .A(n19138), .B(n19063), .Z(n19141) );
  IV U19409 ( .A(n19064), .Z(n19066) );
  XOR U19410 ( .A(n19066), .B(n19065), .Z(n19134) );
  NOR U19411 ( .A(n101), .B(n62), .Z(n19135) );
  IV U19412 ( .A(n19135), .Z(n19067) );
  NOR U19413 ( .A(n19134), .B(n19067), .Z(n19137) );
  IV U19414 ( .A(n19068), .Z(n19070) );
  XOR U19415 ( .A(n19070), .B(n19069), .Z(n19130) );
  NOR U19416 ( .A(n100), .B(n62), .Z(n19131) );
  IV U19417 ( .A(n19131), .Z(n19071) );
  NOR U19418 ( .A(n19130), .B(n19071), .Z(n19133) );
  IV U19419 ( .A(n19072), .Z(n19074) );
  XOR U19420 ( .A(n19074), .B(n19073), .Z(n19126) );
  NOR U19421 ( .A(n99), .B(n62), .Z(n19127) );
  IV U19422 ( .A(n19127), .Z(n19075) );
  NOR U19423 ( .A(n19126), .B(n19075), .Z(n19129) );
  IV U19424 ( .A(n19076), .Z(n19078) );
  XOR U19425 ( .A(n19078), .B(n19077), .Z(n19122) );
  NOR U19426 ( .A(n98), .B(n62), .Z(n19123) );
  IV U19427 ( .A(n19123), .Z(n19079) );
  NOR U19428 ( .A(n19122), .B(n19079), .Z(n19125) );
  XOR U19429 ( .A(n19081), .B(n19080), .Z(n19118) );
  NOR U19430 ( .A(n91), .B(n62), .Z(n19119) );
  IV U19431 ( .A(n19119), .Z(n19082) );
  NOR U19432 ( .A(n19118), .B(n19082), .Z(n19121) );
  XOR U19433 ( .A(n19084), .B(n19083), .Z(n19106) );
  IV U19434 ( .A(n19106), .Z(n19086) );
  NOR U19435 ( .A(n96), .B(n62), .Z(n19085) );
  IV U19436 ( .A(n19085), .Z(n19107) );
  NOR U19437 ( .A(n19086), .B(n19107), .Z(n19109) );
  NOR U19438 ( .A(n95), .B(n62), .Z(n19103) );
  IV U19439 ( .A(n19103), .Z(n19089) );
  XOR U19440 ( .A(n19088), .B(n19087), .Z(n19102) );
  NOR U19441 ( .A(n19089), .B(n19102), .Z(n19105) );
  NOR U19442 ( .A(n62), .B(n93), .Z(n20165) );
  IV U19443 ( .A(n20165), .Z(n19090) );
  NOR U19444 ( .A(n61), .B(n168), .Z(n19098) );
  IV U19445 ( .A(n19098), .Z(n19093) );
  NOR U19446 ( .A(n19090), .B(n19093), .Z(n19091) );
  IV U19447 ( .A(n19091), .Z(n19092) );
  NOR U19448 ( .A(n94), .B(n19092), .Z(n19101) );
  NOR U19449 ( .A(n19093), .B(n93), .Z(n19094) );
  XOR U19450 ( .A(n94), .B(n19094), .Z(n19095) );
  NOR U19451 ( .A(n62), .B(n19095), .Z(n19096) );
  IV U19452 ( .A(n19096), .Z(n19484) );
  XOR U19453 ( .A(n19098), .B(n19097), .Z(n19483) );
  IV U19454 ( .A(n19483), .Z(n19099) );
  NOR U19455 ( .A(n19484), .B(n19099), .Z(n19100) );
  NOR U19456 ( .A(n19101), .B(n19100), .Z(n19479) );
  XOR U19457 ( .A(n19103), .B(n19102), .Z(n19480) );
  NOR U19458 ( .A(n19479), .B(n19480), .Z(n19104) );
  NOR U19459 ( .A(n19105), .B(n19104), .Z(n19507) );
  XOR U19460 ( .A(n19107), .B(n19106), .Z(n19506) );
  NOR U19461 ( .A(n19507), .B(n19506), .Z(n19108) );
  NOR U19462 ( .A(n19109), .B(n19108), .Z(n19114) );
  XOR U19463 ( .A(n19111), .B(n19110), .Z(n19113) );
  IV U19464 ( .A(n19113), .Z(n19112) );
  NOR U19465 ( .A(n19114), .B(n19112), .Z(n19117) );
  XOR U19466 ( .A(n19114), .B(n19113), .Z(n19476) );
  NOR U19467 ( .A(n97), .B(n62), .Z(n19477) );
  IV U19468 ( .A(n19477), .Z(n19115) );
  NOR U19469 ( .A(n19476), .B(n19115), .Z(n19116) );
  NOR U19470 ( .A(n19117), .B(n19116), .Z(n19472) );
  XOR U19471 ( .A(n19119), .B(n19118), .Z(n19473) );
  NOR U19472 ( .A(n19472), .B(n19473), .Z(n19120) );
  NOR U19473 ( .A(n19121), .B(n19120), .Z(n19468) );
  XOR U19474 ( .A(n19123), .B(n19122), .Z(n19469) );
  NOR U19475 ( .A(n19468), .B(n19469), .Z(n19124) );
  NOR U19476 ( .A(n19125), .B(n19124), .Z(n19464) );
  XOR U19477 ( .A(n19127), .B(n19126), .Z(n19465) );
  NOR U19478 ( .A(n19464), .B(n19465), .Z(n19128) );
  NOR U19479 ( .A(n19129), .B(n19128), .Z(n19460) );
  XOR U19480 ( .A(n19131), .B(n19130), .Z(n19461) );
  NOR U19481 ( .A(n19460), .B(n19461), .Z(n19132) );
  NOR U19482 ( .A(n19133), .B(n19132), .Z(n19456) );
  XOR U19483 ( .A(n19135), .B(n19134), .Z(n19457) );
  NOR U19484 ( .A(n19456), .B(n19457), .Z(n19136) );
  NOR U19485 ( .A(n19137), .B(n19136), .Z(n19452) );
  XOR U19486 ( .A(n19139), .B(n19138), .Z(n19453) );
  NOR U19487 ( .A(n19452), .B(n19453), .Z(n19140) );
  NOR U19488 ( .A(n19141), .B(n19140), .Z(n19448) );
  XOR U19489 ( .A(n19143), .B(n19142), .Z(n19449) );
  NOR U19490 ( .A(n19448), .B(n19449), .Z(n19144) );
  NOR U19491 ( .A(n19145), .B(n19144), .Z(n19445) );
  XOR U19492 ( .A(n19147), .B(n19146), .Z(n19444) );
  NOR U19493 ( .A(n19445), .B(n19444), .Z(n19148) );
  NOR U19494 ( .A(n19149), .B(n19148), .Z(n19551) );
  XOR U19495 ( .A(n19151), .B(n19150), .Z(n19550) );
  NOR U19496 ( .A(n19551), .B(n19550), .Z(n19152) );
  NOR U19497 ( .A(n19153), .B(n19152), .Z(n19440) );
  XOR U19498 ( .A(n19155), .B(n19154), .Z(n19441) );
  NOR U19499 ( .A(n19440), .B(n19441), .Z(n19156) );
  NOR U19500 ( .A(n19157), .B(n19156), .Z(n19436) );
  XOR U19501 ( .A(n19159), .B(n19158), .Z(n19437) );
  NOR U19502 ( .A(n19436), .B(n19437), .Z(n19160) );
  NOR U19503 ( .A(n19161), .B(n19160), .Z(n19432) );
  XOR U19504 ( .A(n19163), .B(n19162), .Z(n19433) );
  NOR U19505 ( .A(n19432), .B(n19433), .Z(n19164) );
  NOR U19506 ( .A(n19165), .B(n19164), .Z(n19428) );
  XOR U19507 ( .A(n19167), .B(n19166), .Z(n19429) );
  NOR U19508 ( .A(n19428), .B(n19429), .Z(n19168) );
  NOR U19509 ( .A(n19169), .B(n19168), .Z(n19425) );
  XOR U19510 ( .A(n19171), .B(n19170), .Z(n19424) );
  NOR U19511 ( .A(n19425), .B(n19424), .Z(n19172) );
  NOR U19512 ( .A(n19173), .B(n19172), .Z(n19420) );
  XOR U19513 ( .A(n19175), .B(n19174), .Z(n19421) );
  NOR U19514 ( .A(n19420), .B(n19421), .Z(n19176) );
  NOR U19515 ( .A(n19177), .B(n19176), .Z(n19182) );
  XOR U19516 ( .A(n19179), .B(n19178), .Z(n19181) );
  IV U19517 ( .A(n19181), .Z(n19180) );
  NOR U19518 ( .A(n19182), .B(n19180), .Z(n19185) );
  XOR U19519 ( .A(n19182), .B(n19181), .Z(n19417) );
  NOR U19520 ( .A(n108), .B(n62), .Z(n19418) );
  IV U19521 ( .A(n19418), .Z(n19183) );
  NOR U19522 ( .A(n19417), .B(n19183), .Z(n19184) );
  NOR U19523 ( .A(n19185), .B(n19184), .Z(n19413) );
  XOR U19524 ( .A(n19187), .B(n19186), .Z(n19414) );
  NOR U19525 ( .A(n19413), .B(n19414), .Z(n19188) );
  NOR U19526 ( .A(n19189), .B(n19188), .Z(n19409) );
  XOR U19527 ( .A(n19191), .B(n19190), .Z(n19410) );
  NOR U19528 ( .A(n19409), .B(n19410), .Z(n19192) );
  NOR U19529 ( .A(n19193), .B(n19192), .Z(n19405) );
  XOR U19530 ( .A(n19195), .B(n19194), .Z(n19406) );
  NOR U19531 ( .A(n19405), .B(n19406), .Z(n19196) );
  NOR U19532 ( .A(n19197), .B(n19196), .Z(n19404) );
  XOR U19533 ( .A(n19199), .B(n19198), .Z(n19403) );
  NOR U19534 ( .A(n19404), .B(n19403), .Z(n19200) );
  NOR U19535 ( .A(n19201), .B(n19200), .Z(n19202) );
  IV U19536 ( .A(n19202), .Z(n19401) );
  XOR U19537 ( .A(n19204), .B(n19203), .Z(n19205) );
  IV U19538 ( .A(n19205), .Z(n19400) );
  NOR U19539 ( .A(n19401), .B(n19400), .Z(n19206) );
  NOR U19540 ( .A(n19207), .B(n19206), .Z(n19208) );
  IV U19541 ( .A(n19208), .Z(n19399) );
  XOR U19542 ( .A(n19210), .B(n19209), .Z(n19398) );
  NOR U19543 ( .A(n19399), .B(n19398), .Z(n19211) );
  NOR U19544 ( .A(n19212), .B(n19211), .Z(n19213) );
  IV U19545 ( .A(n19213), .Z(n19395) );
  NOR U19546 ( .A(n19396), .B(n19395), .Z(n19214) );
  NOR U19547 ( .A(n19215), .B(n19214), .Z(n19216) );
  IV U19548 ( .A(n19216), .Z(n19394) );
  XOR U19549 ( .A(n19218), .B(n19217), .Z(n19393) );
  NOR U19550 ( .A(n19394), .B(n19393), .Z(n19219) );
  NOR U19551 ( .A(n19220), .B(n19219), .Z(n19221) );
  IV U19552 ( .A(n19221), .Z(n19391) );
  XOR U19553 ( .A(n19223), .B(n19222), .Z(n19224) );
  IV U19554 ( .A(n19224), .Z(n19390) );
  NOR U19555 ( .A(n19391), .B(n19390), .Z(n19225) );
  NOR U19556 ( .A(n19226), .B(n19225), .Z(n19227) );
  IV U19557 ( .A(n19227), .Z(n19389) );
  XOR U19558 ( .A(n19229), .B(n19228), .Z(n19388) );
  NOR U19559 ( .A(n19389), .B(n19388), .Z(n19230) );
  NOR U19560 ( .A(n19231), .B(n19230), .Z(n19232) );
  IV U19561 ( .A(n19232), .Z(n19386) );
  XOR U19562 ( .A(n19234), .B(n19233), .Z(n19235) );
  IV U19563 ( .A(n19235), .Z(n19385) );
  NOR U19564 ( .A(n19386), .B(n19385), .Z(n19236) );
  NOR U19565 ( .A(n19237), .B(n19236), .Z(n19238) );
  IV U19566 ( .A(n19238), .Z(n19384) );
  XOR U19567 ( .A(n19240), .B(n19239), .Z(n19383) );
  NOR U19568 ( .A(n19384), .B(n19383), .Z(n19241) );
  NOR U19569 ( .A(n19242), .B(n19241), .Z(n19243) );
  IV U19570 ( .A(n19243), .Z(n19381) );
  XOR U19571 ( .A(n19245), .B(n19244), .Z(n19246) );
  IV U19572 ( .A(n19246), .Z(n19380) );
  NOR U19573 ( .A(n19381), .B(n19380), .Z(n19247) );
  NOR U19574 ( .A(n19248), .B(n19247), .Z(n19249) );
  IV U19575 ( .A(n19249), .Z(n19379) );
  XOR U19576 ( .A(n19251), .B(n19250), .Z(n19378) );
  NOR U19577 ( .A(n19379), .B(n19378), .Z(n19252) );
  NOR U19578 ( .A(n19253), .B(n19252), .Z(n19376) );
  IV U19579 ( .A(n19376), .Z(n19254) );
  NOR U19580 ( .A(n19255), .B(n19254), .Z(n19256) );
  NOR U19581 ( .A(n19257), .B(n19256), .Z(n19264) );
  IV U19582 ( .A(n19264), .Z(n19259) );
  NOR U19583 ( .A(n117), .B(n62), .Z(n19258) );
  IV U19584 ( .A(n19258), .Z(n19263) );
  NOR U19585 ( .A(n19259), .B(n19263), .Z(n19266) );
  IV U19586 ( .A(n19260), .Z(n19262) );
  XOR U19587 ( .A(n19262), .B(n19261), .Z(n19370) );
  XOR U19588 ( .A(n19264), .B(n19263), .Z(n19369) );
  NOR U19589 ( .A(n19370), .B(n19369), .Z(n19265) );
  NOR U19590 ( .A(n19266), .B(n19265), .Z(n19673) );
  NOR U19591 ( .A(n19268), .B(n19267), .Z(n19269) );
  NOR U19592 ( .A(n19673), .B(n19269), .Z(n19270) );
  NOR U19593 ( .A(n19271), .B(n19270), .Z(n19368) );
  XOR U19594 ( .A(n19273), .B(n19272), .Z(n19367) );
  NOR U19595 ( .A(n19368), .B(n19367), .Z(n19274) );
  NOR U19596 ( .A(n19275), .B(n19274), .Z(n19365) );
  IV U19597 ( .A(n19365), .Z(n19276) );
  NOR U19598 ( .A(n19277), .B(n19276), .Z(n19278) );
  NOR U19599 ( .A(n19279), .B(n19278), .Z(n19280) );
  IV U19600 ( .A(n19280), .Z(n19286) );
  NOR U19601 ( .A(n19281), .B(n19286), .Z(n19289) );
  XOR U19602 ( .A(n19283), .B(n19282), .Z(n19284) );
  XOR U19603 ( .A(n19285), .B(n19284), .Z(n19359) );
  XOR U19604 ( .A(n19287), .B(n19286), .Z(n19358) );
  NOR U19605 ( .A(n19359), .B(n19358), .Z(n19288) );
  NOR U19606 ( .A(n19289), .B(n19288), .Z(n19694) );
  NOR U19607 ( .A(n19291), .B(n19290), .Z(n19292) );
  NOR U19608 ( .A(n19694), .B(n19292), .Z(n19293) );
  NOR U19609 ( .A(n19294), .B(n19293), .Z(n19300) );
  NOR U19610 ( .A(n126), .B(n62), .Z(n19301) );
  IV U19611 ( .A(n19301), .Z(n19295) );
  NOR U19612 ( .A(n19300), .B(n19295), .Z(n19303) );
  XOR U19613 ( .A(n19297), .B(n19296), .Z(n19298) );
  XOR U19614 ( .A(n19299), .B(n19298), .Z(n19355) );
  XOR U19615 ( .A(n19301), .B(n19300), .Z(n19354) );
  NOR U19616 ( .A(n19355), .B(n19354), .Z(n19302) );
  NOR U19617 ( .A(n19303), .B(n19302), .Z(n19708) );
  IV U19618 ( .A(n19708), .Z(n19304) );
  NOR U19619 ( .A(n19305), .B(n19304), .Z(n19306) );
  NOR U19620 ( .A(n19307), .B(n19306), .Z(n19308) );
  IV U19621 ( .A(n19308), .Z(n19315) );
  NOR U19622 ( .A(n131), .B(n62), .Z(n19314) );
  IV U19623 ( .A(n19314), .Z(n19309) );
  NOR U19624 ( .A(n19315), .B(n19309), .Z(n19317) );
  XOR U19625 ( .A(n19311), .B(n19310), .Z(n19312) );
  XOR U19626 ( .A(n19313), .B(n19312), .Z(n19351) );
  XOR U19627 ( .A(n19315), .B(n19314), .Z(n19350) );
  NOR U19628 ( .A(n19351), .B(n19350), .Z(n19316) );
  NOR U19629 ( .A(n19317), .B(n19316), .Z(n19320) );
  NOR U19630 ( .A(n133), .B(n62), .Z(n19319) );
  IV U19631 ( .A(n19319), .Z(n19318) );
  NOR U19632 ( .A(n19320), .B(n19318), .Z(n19324) );
  XOR U19633 ( .A(n19320), .B(n19319), .Z(n19720) );
  XOR U19634 ( .A(n19322), .B(n19321), .Z(n19721) );
  NOR U19635 ( .A(n19720), .B(n19721), .Z(n19323) );
  NOR U19636 ( .A(n19324), .B(n19323), .Z(n19329) );
  XOR U19637 ( .A(n19326), .B(n19325), .Z(n19328) );
  IV U19638 ( .A(n19328), .Z(n19327) );
  NOR U19639 ( .A(n19329), .B(n19327), .Z(n19332) );
  XOR U19640 ( .A(n19329), .B(n19328), .Z(n19728) );
  NOR U19641 ( .A(n135), .B(n62), .Z(n19729) );
  IV U19642 ( .A(n19729), .Z(n19330) );
  NOR U19643 ( .A(n19728), .B(n19330), .Z(n19331) );
  NOR U19644 ( .A(n19332), .B(n19331), .Z(n19335) );
  NOR U19645 ( .A(n137), .B(n62), .Z(n19334) );
  IV U19646 ( .A(n19334), .Z(n19333) );
  NOR U19647 ( .A(n19335), .B(n19333), .Z(n19339) );
  XOR U19648 ( .A(n19335), .B(n19334), .Z(n19735) );
  XOR U19649 ( .A(n19337), .B(n19336), .Z(n19736) );
  NOR U19650 ( .A(n19735), .B(n19736), .Z(n19338) );
  NOR U19651 ( .A(n19339), .B(n19338), .Z(n19346) );
  NOR U19652 ( .A(n139), .B(n62), .Z(n19345) );
  IV U19653 ( .A(n19345), .Z(n19340) );
  NOR U19654 ( .A(n19346), .B(n19340), .Z(n19348) );
  XOR U19655 ( .A(n19342), .B(n19341), .Z(n19343) );
  XOR U19656 ( .A(n19344), .B(n19343), .Z(n19741) );
  XOR U19657 ( .A(n19346), .B(n19345), .Z(n19740) );
  NOR U19658 ( .A(n19741), .B(n19740), .Z(n19347) );
  NOR U19659 ( .A(n19348), .B(n19347), .Z(n19756) );
  IV U19660 ( .A(n19756), .Z(n19753) );
  XOR U19661 ( .A(n19755), .B(n19753), .Z(n19349) );
  XOR U19662 ( .A(n19757), .B(n19349), .Z(n20415) );
  IV U19663 ( .A(n20415), .Z(n19748) );
  NOR U19664 ( .A(n133), .B(n63), .Z(n19714) );
  IV U19665 ( .A(n19714), .Z(n19353) );
  XOR U19666 ( .A(n19351), .B(n19350), .Z(n19352) );
  IV U19667 ( .A(n19352), .Z(n19713) );
  NOR U19668 ( .A(n19353), .B(n19713), .Z(n19716) );
  NOR U19669 ( .A(n128), .B(n63), .Z(n19356) );
  XOR U19670 ( .A(n19355), .B(n19354), .Z(n19357) );
  NOR U19671 ( .A(n19356), .B(n19357), .Z(n19702) );
  IV U19672 ( .A(n19356), .Z(n20372) );
  IV U19673 ( .A(n19357), .Z(n20371) );
  NOR U19674 ( .A(n20372), .B(n20371), .Z(n19700) );
  XOR U19675 ( .A(n19359), .B(n19358), .Z(n19361) );
  IV U19676 ( .A(n19361), .Z(n20025) );
  NOR U19677 ( .A(n125), .B(n63), .Z(n19360) );
  IV U19678 ( .A(n19360), .Z(n20024) );
  NOR U19679 ( .A(n20025), .B(n20024), .Z(n19689) );
  NOR U19680 ( .A(n19361), .B(n19360), .Z(n19687) );
  XOR U19681 ( .A(n19363), .B(n19362), .Z(n19364) );
  XOR U19682 ( .A(n19365), .B(n19364), .Z(n19684) );
  NOR U19683 ( .A(n123), .B(n63), .Z(n19683) );
  IV U19684 ( .A(n19683), .Z(n19366) );
  NOR U19685 ( .A(n19684), .B(n19366), .Z(n19686) );
  XOR U19686 ( .A(n19368), .B(n19367), .Z(n19679) );
  IV U19687 ( .A(n19679), .Z(n20351) );
  NOR U19688 ( .A(n120), .B(n63), .Z(n19678) );
  IV U19689 ( .A(n19678), .Z(n20350) );
  NOR U19690 ( .A(n20351), .B(n20350), .Z(n19682) );
  NOR U19691 ( .A(n79), .B(n63), .Z(n19371) );
  XOR U19692 ( .A(n19370), .B(n19369), .Z(n19372) );
  NOR U19693 ( .A(n19371), .B(n19372), .Z(n19667) );
  IV U19694 ( .A(n19371), .Z(n20038) );
  IV U19695 ( .A(n19372), .Z(n20037) );
  NOR U19696 ( .A(n20038), .B(n20037), .Z(n19665) );
  XOR U19697 ( .A(n19374), .B(n19373), .Z(n19375) );
  XOR U19698 ( .A(n19376), .B(n19375), .Z(n19661) );
  NOR U19699 ( .A(n117), .B(n63), .Z(n19660) );
  IV U19700 ( .A(n19660), .Z(n19377) );
  NOR U19701 ( .A(n19661), .B(n19377), .Z(n19663) );
  NOR U19702 ( .A(n80), .B(n63), .Z(n19655) );
  XOR U19703 ( .A(n19379), .B(n19378), .Z(n19654) );
  NOR U19704 ( .A(n19655), .B(n19654), .Z(n19658) );
  XOR U19705 ( .A(n19381), .B(n19380), .Z(n19650) );
  NOR U19706 ( .A(n116), .B(n63), .Z(n19649) );
  IV U19707 ( .A(n19649), .Z(n19382) );
  NOR U19708 ( .A(n19650), .B(n19382), .Z(n19652) );
  NOR U19709 ( .A(n81), .B(n63), .Z(n19644) );
  XOR U19710 ( .A(n19384), .B(n19383), .Z(n19643) );
  NOR U19711 ( .A(n19644), .B(n19643), .Z(n19647) );
  XOR U19712 ( .A(n19386), .B(n19385), .Z(n19639) );
  NOR U19713 ( .A(n115), .B(n63), .Z(n19638) );
  IV U19714 ( .A(n19638), .Z(n19387) );
  NOR U19715 ( .A(n19639), .B(n19387), .Z(n19641) );
  NOR U19716 ( .A(n82), .B(n63), .Z(n19633) );
  XOR U19717 ( .A(n19389), .B(n19388), .Z(n19632) );
  NOR U19718 ( .A(n19633), .B(n19632), .Z(n19636) );
  XOR U19719 ( .A(n19391), .B(n19390), .Z(n19628) );
  NOR U19720 ( .A(n114), .B(n63), .Z(n19627) );
  IV U19721 ( .A(n19627), .Z(n19392) );
  NOR U19722 ( .A(n19628), .B(n19392), .Z(n19630) );
  NOR U19723 ( .A(n83), .B(n63), .Z(n19622) );
  XOR U19724 ( .A(n19394), .B(n19393), .Z(n19621) );
  NOR U19725 ( .A(n19622), .B(n19621), .Z(n19625) );
  XOR U19726 ( .A(n19396), .B(n19395), .Z(n19617) );
  NOR U19727 ( .A(n113), .B(n63), .Z(n19616) );
  IV U19728 ( .A(n19616), .Z(n19397) );
  NOR U19729 ( .A(n19617), .B(n19397), .Z(n19619) );
  NOR U19730 ( .A(n84), .B(n63), .Z(n19611) );
  XOR U19731 ( .A(n19399), .B(n19398), .Z(n19610) );
  NOR U19732 ( .A(n19611), .B(n19610), .Z(n19614) );
  XOR U19733 ( .A(n19401), .B(n19400), .Z(n19606) );
  NOR U19734 ( .A(n112), .B(n63), .Z(n19605) );
  IV U19735 ( .A(n19605), .Z(n19402) );
  NOR U19736 ( .A(n19606), .B(n19402), .Z(n19608) );
  NOR U19737 ( .A(n85), .B(n63), .Z(n19600) );
  XOR U19738 ( .A(n19404), .B(n19403), .Z(n19599) );
  NOR U19739 ( .A(n19600), .B(n19599), .Z(n19603) );
  IV U19740 ( .A(n19405), .Z(n19407) );
  XOR U19741 ( .A(n19407), .B(n19406), .Z(n19594) );
  NOR U19742 ( .A(n111), .B(n63), .Z(n19595) );
  IV U19743 ( .A(n19595), .Z(n19408) );
  NOR U19744 ( .A(n19594), .B(n19408), .Z(n19597) );
  IV U19745 ( .A(n19409), .Z(n19411) );
  XOR U19746 ( .A(n19411), .B(n19410), .Z(n19590) );
  NOR U19747 ( .A(n86), .B(n63), .Z(n19591) );
  IV U19748 ( .A(n19591), .Z(n19412) );
  NOR U19749 ( .A(n19590), .B(n19412), .Z(n19593) );
  IV U19750 ( .A(n19413), .Z(n19415) );
  XOR U19751 ( .A(n19415), .B(n19414), .Z(n19586) );
  NOR U19752 ( .A(n110), .B(n63), .Z(n19587) );
  IV U19753 ( .A(n19587), .Z(n19416) );
  NOR U19754 ( .A(n19586), .B(n19416), .Z(n19589) );
  XOR U19755 ( .A(n19418), .B(n19417), .Z(n19582) );
  NOR U19756 ( .A(n109), .B(n63), .Z(n19583) );
  IV U19757 ( .A(n19583), .Z(n19419) );
  NOR U19758 ( .A(n19582), .B(n19419), .Z(n19585) );
  IV U19759 ( .A(n19420), .Z(n19422) );
  XOR U19760 ( .A(n19422), .B(n19421), .Z(n19578) );
  NOR U19761 ( .A(n108), .B(n63), .Z(n19579) );
  IV U19762 ( .A(n19579), .Z(n19423) );
  NOR U19763 ( .A(n19578), .B(n19423), .Z(n19581) );
  XOR U19764 ( .A(n19425), .B(n19424), .Z(n19574) );
  IV U19765 ( .A(n19574), .Z(n19427) );
  NOR U19766 ( .A(n87), .B(n63), .Z(n19426) );
  IV U19767 ( .A(n19426), .Z(n19575) );
  NOR U19768 ( .A(n19427), .B(n19575), .Z(n19577) );
  IV U19769 ( .A(n19428), .Z(n19430) );
  XOR U19770 ( .A(n19430), .B(n19429), .Z(n19570) );
  NOR U19771 ( .A(n107), .B(n63), .Z(n19571) );
  IV U19772 ( .A(n19571), .Z(n19431) );
  NOR U19773 ( .A(n19570), .B(n19431), .Z(n19573) );
  IV U19774 ( .A(n19432), .Z(n19434) );
  XOR U19775 ( .A(n19434), .B(n19433), .Z(n19566) );
  NOR U19776 ( .A(n88), .B(n63), .Z(n19567) );
  IV U19777 ( .A(n19567), .Z(n19435) );
  NOR U19778 ( .A(n19566), .B(n19435), .Z(n19569) );
  IV U19779 ( .A(n19436), .Z(n19438) );
  XOR U19780 ( .A(n19438), .B(n19437), .Z(n19562) );
  NOR U19781 ( .A(n106), .B(n63), .Z(n19563) );
  IV U19782 ( .A(n19563), .Z(n19439) );
  NOR U19783 ( .A(n19562), .B(n19439), .Z(n19565) );
  IV U19784 ( .A(n19440), .Z(n19442) );
  XOR U19785 ( .A(n19442), .B(n19441), .Z(n19558) );
  NOR U19786 ( .A(n105), .B(n63), .Z(n19559) );
  IV U19787 ( .A(n19559), .Z(n19443) );
  NOR U19788 ( .A(n19558), .B(n19443), .Z(n19561) );
  XOR U19789 ( .A(n19445), .B(n19444), .Z(n19546) );
  IV U19790 ( .A(n19546), .Z(n19447) );
  NOR U19791 ( .A(n89), .B(n63), .Z(n19446) );
  IV U19792 ( .A(n19446), .Z(n19547) );
  NOR U19793 ( .A(n19447), .B(n19547), .Z(n19549) );
  IV U19794 ( .A(n19448), .Z(n19450) );
  XOR U19795 ( .A(n19450), .B(n19449), .Z(n19542) );
  NOR U19796 ( .A(n103), .B(n63), .Z(n19543) );
  IV U19797 ( .A(n19543), .Z(n19451) );
  NOR U19798 ( .A(n19542), .B(n19451), .Z(n19545) );
  IV U19799 ( .A(n19452), .Z(n19454) );
  XOR U19800 ( .A(n19454), .B(n19453), .Z(n19538) );
  NOR U19801 ( .A(n90), .B(n63), .Z(n19539) );
  IV U19802 ( .A(n19539), .Z(n19455) );
  NOR U19803 ( .A(n19538), .B(n19455), .Z(n19541) );
  IV U19804 ( .A(n19456), .Z(n19458) );
  XOR U19805 ( .A(n19458), .B(n19457), .Z(n19534) );
  NOR U19806 ( .A(n102), .B(n63), .Z(n19535) );
  IV U19807 ( .A(n19535), .Z(n19459) );
  NOR U19808 ( .A(n19534), .B(n19459), .Z(n19537) );
  IV U19809 ( .A(n19460), .Z(n19462) );
  XOR U19810 ( .A(n19462), .B(n19461), .Z(n19530) );
  NOR U19811 ( .A(n101), .B(n63), .Z(n19531) );
  IV U19812 ( .A(n19531), .Z(n19463) );
  NOR U19813 ( .A(n19530), .B(n19463), .Z(n19533) );
  IV U19814 ( .A(n19464), .Z(n19466) );
  XOR U19815 ( .A(n19466), .B(n19465), .Z(n19526) );
  NOR U19816 ( .A(n100), .B(n63), .Z(n19527) );
  IV U19817 ( .A(n19527), .Z(n19467) );
  NOR U19818 ( .A(n19526), .B(n19467), .Z(n19529) );
  IV U19819 ( .A(n19468), .Z(n19470) );
  XOR U19820 ( .A(n19470), .B(n19469), .Z(n19522) );
  NOR U19821 ( .A(n99), .B(n63), .Z(n19523) );
  IV U19822 ( .A(n19523), .Z(n19471) );
  NOR U19823 ( .A(n19522), .B(n19471), .Z(n19525) );
  IV U19824 ( .A(n19472), .Z(n19474) );
  XOR U19825 ( .A(n19474), .B(n19473), .Z(n19518) );
  NOR U19826 ( .A(n98), .B(n63), .Z(n19519) );
  IV U19827 ( .A(n19519), .Z(n19475) );
  NOR U19828 ( .A(n19518), .B(n19475), .Z(n19521) );
  XOR U19829 ( .A(n19477), .B(n19476), .Z(n19514) );
  NOR U19830 ( .A(n91), .B(n63), .Z(n19515) );
  IV U19831 ( .A(n19515), .Z(n19478) );
  NOR U19832 ( .A(n19514), .B(n19478), .Z(n19517) );
  IV U19833 ( .A(n19479), .Z(n19481) );
  XOR U19834 ( .A(n19481), .B(n19480), .Z(n19502) );
  NOR U19835 ( .A(n96), .B(n63), .Z(n19503) );
  IV U19836 ( .A(n19503), .Z(n19482) );
  NOR U19837 ( .A(n19502), .B(n19482), .Z(n19505) );
  NOR U19838 ( .A(n95), .B(n63), .Z(n19499) );
  IV U19839 ( .A(n19499), .Z(n19485) );
  XOR U19840 ( .A(n19484), .B(n19483), .Z(n19498) );
  NOR U19841 ( .A(n19485), .B(n19498), .Z(n19501) );
  NOR U19842 ( .A(n63), .B(n93), .Z(n20649) );
  IV U19843 ( .A(n20649), .Z(n19486) );
  NOR U19844 ( .A(n62), .B(n168), .Z(n19494) );
  IV U19845 ( .A(n19494), .Z(n19489) );
  NOR U19846 ( .A(n19486), .B(n19489), .Z(n19487) );
  IV U19847 ( .A(n19487), .Z(n19488) );
  NOR U19848 ( .A(n94), .B(n19488), .Z(n19497) );
  NOR U19849 ( .A(n19489), .B(n93), .Z(n19490) );
  XOR U19850 ( .A(n94), .B(n19490), .Z(n19491) );
  NOR U19851 ( .A(n63), .B(n19491), .Z(n19492) );
  IV U19852 ( .A(n19492), .Z(n20156) );
  XOR U19853 ( .A(n19494), .B(n19493), .Z(n20155) );
  IV U19854 ( .A(n20155), .Z(n19495) );
  NOR U19855 ( .A(n20156), .B(n19495), .Z(n19496) );
  NOR U19856 ( .A(n19497), .B(n19496), .Z(n20152) );
  XOR U19857 ( .A(n19499), .B(n19498), .Z(n20151) );
  NOR U19858 ( .A(n20152), .B(n20151), .Z(n19500) );
  NOR U19859 ( .A(n19501), .B(n19500), .Z(n20147) );
  XOR U19860 ( .A(n19503), .B(n19502), .Z(n20148) );
  NOR U19861 ( .A(n20147), .B(n20148), .Z(n19504) );
  NOR U19862 ( .A(n19505), .B(n19504), .Z(n19510) );
  XOR U19863 ( .A(n19507), .B(n19506), .Z(n19509) );
  IV U19864 ( .A(n19509), .Z(n19508) );
  NOR U19865 ( .A(n19510), .B(n19508), .Z(n19513) );
  XOR U19866 ( .A(n19510), .B(n19509), .Z(n20144) );
  NOR U19867 ( .A(n97), .B(n63), .Z(n20145) );
  IV U19868 ( .A(n20145), .Z(n19511) );
  NOR U19869 ( .A(n20144), .B(n19511), .Z(n19512) );
  NOR U19870 ( .A(n19513), .B(n19512), .Z(n20140) );
  XOR U19871 ( .A(n19515), .B(n19514), .Z(n20141) );
  NOR U19872 ( .A(n20140), .B(n20141), .Z(n19516) );
  NOR U19873 ( .A(n19517), .B(n19516), .Z(n20136) );
  XOR U19874 ( .A(n19519), .B(n19518), .Z(n20137) );
  NOR U19875 ( .A(n20136), .B(n20137), .Z(n19520) );
  NOR U19876 ( .A(n19521), .B(n19520), .Z(n20132) );
  XOR U19877 ( .A(n19523), .B(n19522), .Z(n20133) );
  NOR U19878 ( .A(n20132), .B(n20133), .Z(n19524) );
  NOR U19879 ( .A(n19525), .B(n19524), .Z(n20128) );
  XOR U19880 ( .A(n19527), .B(n19526), .Z(n20129) );
  NOR U19881 ( .A(n20128), .B(n20129), .Z(n19528) );
  NOR U19882 ( .A(n19529), .B(n19528), .Z(n20124) );
  XOR U19883 ( .A(n19531), .B(n19530), .Z(n20125) );
  NOR U19884 ( .A(n20124), .B(n20125), .Z(n19532) );
  NOR U19885 ( .A(n19533), .B(n19532), .Z(n20120) );
  XOR U19886 ( .A(n19535), .B(n19534), .Z(n20121) );
  NOR U19887 ( .A(n20120), .B(n20121), .Z(n19536) );
  NOR U19888 ( .A(n19537), .B(n19536), .Z(n20116) );
  XOR U19889 ( .A(n19539), .B(n19538), .Z(n20117) );
  NOR U19890 ( .A(n20116), .B(n20117), .Z(n19540) );
  NOR U19891 ( .A(n19541), .B(n19540), .Z(n20113) );
  XOR U19892 ( .A(n19543), .B(n19542), .Z(n20112) );
  NOR U19893 ( .A(n20113), .B(n20112), .Z(n19544) );
  NOR U19894 ( .A(n19545), .B(n19544), .Z(n20219) );
  XOR U19895 ( .A(n19547), .B(n19546), .Z(n20218) );
  NOR U19896 ( .A(n20219), .B(n20218), .Z(n19548) );
  NOR U19897 ( .A(n19549), .B(n19548), .Z(n19554) );
  XOR U19898 ( .A(n19551), .B(n19550), .Z(n19553) );
  IV U19899 ( .A(n19553), .Z(n19552) );
  NOR U19900 ( .A(n19554), .B(n19552), .Z(n19557) );
  XOR U19901 ( .A(n19554), .B(n19553), .Z(n20109) );
  NOR U19902 ( .A(n104), .B(n63), .Z(n20110) );
  IV U19903 ( .A(n20110), .Z(n19555) );
  NOR U19904 ( .A(n20109), .B(n19555), .Z(n19556) );
  NOR U19905 ( .A(n19557), .B(n19556), .Z(n20105) );
  XOR U19906 ( .A(n19559), .B(n19558), .Z(n20106) );
  NOR U19907 ( .A(n20105), .B(n20106), .Z(n19560) );
  NOR U19908 ( .A(n19561), .B(n19560), .Z(n20101) );
  XOR U19909 ( .A(n19563), .B(n19562), .Z(n20102) );
  NOR U19910 ( .A(n20101), .B(n20102), .Z(n19564) );
  NOR U19911 ( .A(n19565), .B(n19564), .Z(n20097) );
  XOR U19912 ( .A(n19567), .B(n19566), .Z(n20098) );
  NOR U19913 ( .A(n20097), .B(n20098), .Z(n19568) );
  NOR U19914 ( .A(n19569), .B(n19568), .Z(n20093) );
  XOR U19915 ( .A(n19571), .B(n19570), .Z(n20094) );
  NOR U19916 ( .A(n20093), .B(n20094), .Z(n19572) );
  NOR U19917 ( .A(n19573), .B(n19572), .Z(n20250) );
  XOR U19918 ( .A(n19575), .B(n19574), .Z(n20249) );
  NOR U19919 ( .A(n20250), .B(n20249), .Z(n19576) );
  NOR U19920 ( .A(n19577), .B(n19576), .Z(n20092) );
  XOR U19921 ( .A(n19579), .B(n19578), .Z(n20091) );
  NOR U19922 ( .A(n20092), .B(n20091), .Z(n19580) );
  NOR U19923 ( .A(n19581), .B(n19580), .Z(n20087) );
  XOR U19924 ( .A(n19583), .B(n19582), .Z(n20088) );
  NOR U19925 ( .A(n20087), .B(n20088), .Z(n19584) );
  NOR U19926 ( .A(n19585), .B(n19584), .Z(n20083) );
  XOR U19927 ( .A(n19587), .B(n19586), .Z(n20084) );
  NOR U19928 ( .A(n20083), .B(n20084), .Z(n19588) );
  NOR U19929 ( .A(n19589), .B(n19588), .Z(n20079) );
  XOR U19930 ( .A(n19591), .B(n19590), .Z(n20080) );
  NOR U19931 ( .A(n20079), .B(n20080), .Z(n19592) );
  NOR U19932 ( .A(n19593), .B(n19592), .Z(n20075) );
  XOR U19933 ( .A(n19595), .B(n19594), .Z(n20076) );
  NOR U19934 ( .A(n20075), .B(n20076), .Z(n19596) );
  NOR U19935 ( .A(n19597), .B(n19596), .Z(n19598) );
  IV U19936 ( .A(n19598), .Z(n20073) );
  XOR U19937 ( .A(n19600), .B(n19599), .Z(n19601) );
  IV U19938 ( .A(n19601), .Z(n20072) );
  NOR U19939 ( .A(n20073), .B(n20072), .Z(n19602) );
  NOR U19940 ( .A(n19603), .B(n19602), .Z(n19604) );
  IV U19941 ( .A(n19604), .Z(n20071) );
  XOR U19942 ( .A(n19606), .B(n19605), .Z(n20070) );
  NOR U19943 ( .A(n20071), .B(n20070), .Z(n19607) );
  NOR U19944 ( .A(n19608), .B(n19607), .Z(n19609) );
  IV U19945 ( .A(n19609), .Z(n20068) );
  XOR U19946 ( .A(n19611), .B(n19610), .Z(n19612) );
  IV U19947 ( .A(n19612), .Z(n20067) );
  NOR U19948 ( .A(n20068), .B(n20067), .Z(n19613) );
  NOR U19949 ( .A(n19614), .B(n19613), .Z(n19615) );
  IV U19950 ( .A(n19615), .Z(n20063) );
  XOR U19951 ( .A(n19617), .B(n19616), .Z(n20062) );
  NOR U19952 ( .A(n20063), .B(n20062), .Z(n19618) );
  NOR U19953 ( .A(n19619), .B(n19618), .Z(n19620) );
  IV U19954 ( .A(n19620), .Z(n20060) );
  XOR U19955 ( .A(n19622), .B(n19621), .Z(n19623) );
  IV U19956 ( .A(n19623), .Z(n20059) );
  NOR U19957 ( .A(n20060), .B(n20059), .Z(n19624) );
  NOR U19958 ( .A(n19625), .B(n19624), .Z(n19626) );
  IV U19959 ( .A(n19626), .Z(n20058) );
  XOR U19960 ( .A(n19628), .B(n19627), .Z(n20057) );
  NOR U19961 ( .A(n20058), .B(n20057), .Z(n19629) );
  NOR U19962 ( .A(n19630), .B(n19629), .Z(n19631) );
  IV U19963 ( .A(n19631), .Z(n20055) );
  XOR U19964 ( .A(n19633), .B(n19632), .Z(n19634) );
  IV U19965 ( .A(n19634), .Z(n20054) );
  NOR U19966 ( .A(n20055), .B(n20054), .Z(n19635) );
  NOR U19967 ( .A(n19636), .B(n19635), .Z(n19637) );
  IV U19968 ( .A(n19637), .Z(n20053) );
  XOR U19969 ( .A(n19639), .B(n19638), .Z(n20052) );
  NOR U19970 ( .A(n20053), .B(n20052), .Z(n19640) );
  NOR U19971 ( .A(n19641), .B(n19640), .Z(n19642) );
  IV U19972 ( .A(n19642), .Z(n20050) );
  XOR U19973 ( .A(n19644), .B(n19643), .Z(n19645) );
  IV U19974 ( .A(n19645), .Z(n20049) );
  NOR U19975 ( .A(n20050), .B(n20049), .Z(n19646) );
  NOR U19976 ( .A(n19647), .B(n19646), .Z(n19648) );
  IV U19977 ( .A(n19648), .Z(n20048) );
  XOR U19978 ( .A(n19650), .B(n19649), .Z(n20047) );
  NOR U19979 ( .A(n20048), .B(n20047), .Z(n19651) );
  NOR U19980 ( .A(n19652), .B(n19651), .Z(n19653) );
  IV U19981 ( .A(n19653), .Z(n20045) );
  XOR U19982 ( .A(n19655), .B(n19654), .Z(n19656) );
  IV U19983 ( .A(n19656), .Z(n20044) );
  NOR U19984 ( .A(n20045), .B(n20044), .Z(n19657) );
  NOR U19985 ( .A(n19658), .B(n19657), .Z(n19659) );
  IV U19986 ( .A(n19659), .Z(n20043) );
  XOR U19987 ( .A(n19661), .B(n19660), .Z(n20042) );
  NOR U19988 ( .A(n20043), .B(n20042), .Z(n19662) );
  NOR U19989 ( .A(n19663), .B(n19662), .Z(n20040) );
  IV U19990 ( .A(n20040), .Z(n19664) );
  NOR U19991 ( .A(n19665), .B(n19664), .Z(n19666) );
  NOR U19992 ( .A(n19667), .B(n19666), .Z(n19668) );
  IV U19993 ( .A(n19668), .Z(n19675) );
  NOR U19994 ( .A(n119), .B(n63), .Z(n19674) );
  IV U19995 ( .A(n19674), .Z(n19669) );
  NOR U19996 ( .A(n19675), .B(n19669), .Z(n19677) );
  XOR U19997 ( .A(n19671), .B(n19670), .Z(n19672) );
  XOR U19998 ( .A(n19673), .B(n19672), .Z(n20033) );
  XOR U19999 ( .A(n19675), .B(n19674), .Z(n20034) );
  NOR U20000 ( .A(n20033), .B(n20034), .Z(n19676) );
  NOR U20001 ( .A(n19677), .B(n19676), .Z(n20353) );
  NOR U20002 ( .A(n19679), .B(n19678), .Z(n19680) );
  NOR U20003 ( .A(n20353), .B(n19680), .Z(n19681) );
  NOR U20004 ( .A(n19682), .B(n19681), .Z(n20031) );
  XOR U20005 ( .A(n19684), .B(n19683), .Z(n20030) );
  NOR U20006 ( .A(n20031), .B(n20030), .Z(n19685) );
  NOR U20007 ( .A(n19686), .B(n19685), .Z(n20027) );
  NOR U20008 ( .A(n19687), .B(n20027), .Z(n19688) );
  NOR U20009 ( .A(n19689), .B(n19688), .Z(n19695) );
  NOR U20010 ( .A(n126), .B(n63), .Z(n19696) );
  IV U20011 ( .A(n19696), .Z(n19690) );
  NOR U20012 ( .A(n19695), .B(n19690), .Z(n19698) );
  XOR U20013 ( .A(n19692), .B(n19691), .Z(n19693) );
  XOR U20014 ( .A(n19694), .B(n19693), .Z(n20021) );
  XOR U20015 ( .A(n19696), .B(n19695), .Z(n20020) );
  NOR U20016 ( .A(n20021), .B(n20020), .Z(n19697) );
  NOR U20017 ( .A(n19698), .B(n19697), .Z(n20374) );
  IV U20018 ( .A(n20374), .Z(n19699) );
  NOR U20019 ( .A(n19700), .B(n19699), .Z(n19701) );
  NOR U20020 ( .A(n19702), .B(n19701), .Z(n19703) );
  IV U20021 ( .A(n19703), .Z(n19710) );
  NOR U20022 ( .A(n131), .B(n63), .Z(n19709) );
  IV U20023 ( .A(n19709), .Z(n19704) );
  NOR U20024 ( .A(n19710), .B(n19704), .Z(n19712) );
  XOR U20025 ( .A(n19706), .B(n19705), .Z(n19707) );
  XOR U20026 ( .A(n19708), .B(n19707), .Z(n20016) );
  XOR U20027 ( .A(n19710), .B(n19709), .Z(n20017) );
  NOR U20028 ( .A(n20016), .B(n20017), .Z(n19711) );
  NOR U20029 ( .A(n19712), .B(n19711), .Z(n20386) );
  XOR U20030 ( .A(n19714), .B(n19713), .Z(n20387) );
  NOR U20031 ( .A(n20386), .B(n20387), .Z(n19715) );
  NOR U20032 ( .A(n19716), .B(n19715), .Z(n19719) );
  NOR U20033 ( .A(n135), .B(n63), .Z(n19718) );
  IV U20034 ( .A(n19718), .Z(n19717) );
  NOR U20035 ( .A(n19719), .B(n19717), .Z(n19724) );
  XOR U20036 ( .A(n19719), .B(n19718), .Z(n20012) );
  XOR U20037 ( .A(n19721), .B(n19720), .Z(n20013) );
  IV U20038 ( .A(n20013), .Z(n19722) );
  NOR U20039 ( .A(n20012), .B(n19722), .Z(n19723) );
  NOR U20040 ( .A(n19724), .B(n19723), .Z(n19727) );
  NOR U20041 ( .A(n137), .B(n63), .Z(n19726) );
  IV U20042 ( .A(n19726), .Z(n19725) );
  NOR U20043 ( .A(n19727), .B(n19725), .Z(n19731) );
  XOR U20044 ( .A(n19727), .B(n19726), .Z(n20395) );
  XOR U20045 ( .A(n19729), .B(n19728), .Z(n20396) );
  NOR U20046 ( .A(n20395), .B(n20396), .Z(n19730) );
  NOR U20047 ( .A(n19731), .B(n19730), .Z(n19734) );
  NOR U20048 ( .A(n139), .B(n63), .Z(n19733) );
  IV U20049 ( .A(n19733), .Z(n19732) );
  NOR U20050 ( .A(n19734), .B(n19732), .Z(n19739) );
  XOR U20051 ( .A(n19734), .B(n19733), .Z(n20009) );
  XOR U20052 ( .A(n19736), .B(n19735), .Z(n20010) );
  IV U20053 ( .A(n20010), .Z(n19737) );
  NOR U20054 ( .A(n20009), .B(n19737), .Z(n19738) );
  NOR U20055 ( .A(n19739), .B(n19738), .Z(n19744) );
  XOR U20056 ( .A(n19741), .B(n19740), .Z(n19743) );
  IV U20057 ( .A(n19743), .Z(n19742) );
  NOR U20058 ( .A(n19744), .B(n19742), .Z(n19747) );
  XOR U20059 ( .A(n19744), .B(n19743), .Z(n20410) );
  NOR U20060 ( .A(n141), .B(n63), .Z(n20411) );
  IV U20061 ( .A(n20411), .Z(n19745) );
  NOR U20062 ( .A(n20410), .B(n19745), .Z(n19746) );
  NOR U20063 ( .A(n19747), .B(n19746), .Z(n19749) );
  IV U20064 ( .A(n19749), .Z(n20414) );
  NOR U20065 ( .A(n19748), .B(n20414), .Z(n19752) );
  NOR U20066 ( .A(n19749), .B(n20415), .Z(n19750) );
  NOR U20067 ( .A(n143), .B(n63), .Z(n20417) );
  NOR U20068 ( .A(n19750), .B(n20417), .Z(n19751) );
  NOR U20069 ( .A(n19752), .B(n19751), .Z(n19768) );
  IV U20070 ( .A(n19768), .Z(n19766) );
  NOR U20071 ( .A(n19754), .B(n19753), .Z(n19760) );
  NOR U20072 ( .A(n19756), .B(n19755), .Z(n19758) );
  NOR U20073 ( .A(n19758), .B(n19757), .Z(n19759) );
  NOR U20074 ( .A(n19760), .B(n19759), .Z(n19761) );
  IV U20075 ( .A(n19761), .Z(n19775) );
  NOR U20076 ( .A(n143), .B(n62), .Z(n19773) );
  XOR U20077 ( .A(n19775), .B(n19773), .Z(n19777) );
  XOR U20078 ( .A(n19763), .B(n19762), .Z(n19764) );
  XOR U20079 ( .A(n19765), .B(n19764), .Z(n19776) );
  XOR U20080 ( .A(n19777), .B(n19776), .Z(n19767) );
  NOR U20081 ( .A(n19766), .B(n19767), .Z(n19771) );
  XOR U20082 ( .A(n19768), .B(n19767), .Z(n20005) );
  NOR U20083 ( .A(n145), .B(n63), .Z(n19769) );
  IV U20084 ( .A(n19769), .Z(n20004) );
  NOR U20085 ( .A(n20005), .B(n20004), .Z(n19770) );
  NOR U20086 ( .A(n19771), .B(n19770), .Z(n19783) );
  NOR U20087 ( .A(n145), .B(n62), .Z(n19772) );
  IV U20088 ( .A(n19772), .Z(n19795) );
  IV U20089 ( .A(n19773), .Z(n19774) );
  NOR U20090 ( .A(n19775), .B(n19774), .Z(n19780) );
  IV U20091 ( .A(n19776), .Z(n19778) );
  NOR U20092 ( .A(n19778), .B(n19777), .Z(n19779) );
  NOR U20093 ( .A(n19780), .B(n19779), .Z(n19794) );
  XOR U20094 ( .A(n19782), .B(n19781), .Z(n19792) );
  XOR U20095 ( .A(n19794), .B(n19792), .Z(n19796) );
  XOR U20096 ( .A(n19795), .B(n19796), .Z(n19784) );
  IV U20097 ( .A(n19784), .Z(n20429) );
  NOR U20098 ( .A(n19783), .B(n20429), .Z(n19788) );
  IV U20099 ( .A(n19783), .Z(n20430) );
  NOR U20100 ( .A(n19784), .B(n20430), .Z(n19786) );
  NOR U20101 ( .A(n147), .B(n63), .Z(n20432) );
  IV U20102 ( .A(n20432), .Z(n19785) );
  NOR U20103 ( .A(n19786), .B(n19785), .Z(n19787) );
  NOR U20104 ( .A(n19788), .B(n19787), .Z(n19800) );
  NOR U20105 ( .A(n148), .B(n63), .Z(n19799) );
  IV U20106 ( .A(n19799), .Z(n19789) );
  NOR U20107 ( .A(n19800), .B(n19789), .Z(n19803) );
  XOR U20108 ( .A(n19791), .B(n19790), .Z(n19815) );
  IV U20109 ( .A(n19792), .Z(n19793) );
  NOR U20110 ( .A(n19794), .B(n19793), .Z(n19798) );
  NOR U20111 ( .A(n19796), .B(n19795), .Z(n19797) );
  NOR U20112 ( .A(n19798), .B(n19797), .Z(n19813) );
  NOR U20113 ( .A(n147), .B(n62), .Z(n19811) );
  XOR U20114 ( .A(n19813), .B(n19811), .Z(n19814) );
  XOR U20115 ( .A(n19815), .B(n19814), .Z(n20438) );
  IV U20116 ( .A(n20438), .Z(n19801) );
  XOR U20117 ( .A(n19800), .B(n19799), .Z(n20437) );
  NOR U20118 ( .A(n19801), .B(n20437), .Z(n19802) );
  NOR U20119 ( .A(n19803), .B(n19802), .Z(n19806) );
  NOR U20120 ( .A(n150), .B(n63), .Z(n19805) );
  IV U20121 ( .A(n19805), .Z(n19804) );
  NOR U20122 ( .A(n19806), .B(n19804), .Z(n19820) );
  XOR U20123 ( .A(n19806), .B(n19805), .Z(n20001) );
  NOR U20124 ( .A(n148), .B(n62), .Z(n19823) );
  XOR U20125 ( .A(n19808), .B(n19807), .Z(n19809) );
  XOR U20126 ( .A(n19810), .B(n19809), .Z(n19821) );
  IV U20127 ( .A(n19811), .Z(n19812) );
  NOR U20128 ( .A(n19813), .B(n19812), .Z(n19817) );
  NOR U20129 ( .A(n19815), .B(n19814), .Z(n19816) );
  NOR U20130 ( .A(n19817), .B(n19816), .Z(n19822) );
  XOR U20131 ( .A(n19821), .B(n19822), .Z(n19818) );
  IV U20132 ( .A(n19818), .Z(n19825) );
  XOR U20133 ( .A(n19823), .B(n19825), .Z(n20000) );
  NOR U20134 ( .A(n20001), .B(n20000), .Z(n19819) );
  NOR U20135 ( .A(n19820), .B(n19819), .Z(n19831) );
  NOR U20136 ( .A(n19822), .B(n19821), .Z(n19827) );
  IV U20137 ( .A(n19823), .Z(n19824) );
  NOR U20138 ( .A(n19825), .B(n19824), .Z(n19826) );
  NOR U20139 ( .A(n19827), .B(n19826), .Z(n19844) );
  NOR U20140 ( .A(n150), .B(n62), .Z(n19840) );
  IV U20141 ( .A(n19828), .Z(n19830) );
  XOR U20142 ( .A(n19830), .B(n19829), .Z(n19842) );
  XOR U20143 ( .A(n19840), .B(n19842), .Z(n19843) );
  XOR U20144 ( .A(n19844), .B(n19843), .Z(n19832) );
  IV U20145 ( .A(n19832), .Z(n19995) );
  NOR U20146 ( .A(n19831), .B(n19995), .Z(n19836) );
  IV U20147 ( .A(n19831), .Z(n19996) );
  NOR U20148 ( .A(n19832), .B(n19996), .Z(n19834) );
  NOR U20149 ( .A(n153), .B(n63), .Z(n19998) );
  IV U20150 ( .A(n19998), .Z(n19833) );
  NOR U20151 ( .A(n19834), .B(n19833), .Z(n19835) );
  NOR U20152 ( .A(n19836), .B(n19835), .Z(n19839) );
  NOR U20153 ( .A(n155), .B(n63), .Z(n19838) );
  IV U20154 ( .A(n19838), .Z(n19837) );
  NOR U20155 ( .A(n19839), .B(n19837), .Z(n19853) );
  XOR U20156 ( .A(n19839), .B(n19838), .Z(n20453) );
  IV U20157 ( .A(n19840), .Z(n19841) );
  NOR U20158 ( .A(n19842), .B(n19841), .Z(n19846) );
  NOR U20159 ( .A(n19844), .B(n19843), .Z(n19845) );
  NOR U20160 ( .A(n19846), .B(n19845), .Z(n19858) );
  NOR U20161 ( .A(n153), .B(n62), .Z(n19854) );
  XOR U20162 ( .A(n19848), .B(n19847), .Z(n19849) );
  XOR U20163 ( .A(n19850), .B(n19849), .Z(n19856) );
  XOR U20164 ( .A(n19854), .B(n19856), .Z(n19857) );
  XOR U20165 ( .A(n19858), .B(n19857), .Z(n20454) );
  IV U20166 ( .A(n20454), .Z(n19851) );
  NOR U20167 ( .A(n20453), .B(n19851), .Z(n19852) );
  NOR U20168 ( .A(n19853), .B(n19852), .Z(n19863) );
  IV U20169 ( .A(n19854), .Z(n19855) );
  NOR U20170 ( .A(n19856), .B(n19855), .Z(n19860) );
  NOR U20171 ( .A(n19858), .B(n19857), .Z(n19859) );
  NOR U20172 ( .A(n19860), .B(n19859), .Z(n19878) );
  NOR U20173 ( .A(n155), .B(n62), .Z(n19874) );
  XOR U20174 ( .A(n19862), .B(n19861), .Z(n19876) );
  XOR U20175 ( .A(n19874), .B(n19876), .Z(n19877) );
  XOR U20176 ( .A(n19878), .B(n19877), .Z(n19864) );
  IV U20177 ( .A(n19864), .Z(n19990) );
  NOR U20178 ( .A(n19863), .B(n19990), .Z(n19868) );
  IV U20179 ( .A(n19863), .Z(n19991) );
  NOR U20180 ( .A(n19864), .B(n19991), .Z(n19866) );
  NOR U20181 ( .A(n156), .B(n63), .Z(n19993) );
  IV U20182 ( .A(n19993), .Z(n19865) );
  NOR U20183 ( .A(n19866), .B(n19865), .Z(n19867) );
  NOR U20184 ( .A(n19868), .B(n19867), .Z(n19882) );
  NOR U20185 ( .A(n158), .B(n63), .Z(n19881) );
  IV U20186 ( .A(n19881), .Z(n19869) );
  NOR U20187 ( .A(n19882), .B(n19869), .Z(n19885) );
  XOR U20188 ( .A(n19871), .B(n19870), .Z(n19872) );
  XOR U20189 ( .A(n19873), .B(n19872), .Z(n19894) );
  IV U20190 ( .A(n19874), .Z(n19875) );
  NOR U20191 ( .A(n19876), .B(n19875), .Z(n19880) );
  NOR U20192 ( .A(n19878), .B(n19877), .Z(n19879) );
  NOR U20193 ( .A(n19880), .B(n19879), .Z(n19892) );
  NOR U20194 ( .A(n156), .B(n62), .Z(n19890) );
  XOR U20195 ( .A(n19892), .B(n19890), .Z(n19893) );
  XOR U20196 ( .A(n19894), .B(n19893), .Z(n19988) );
  IV U20197 ( .A(n19988), .Z(n19883) );
  XOR U20198 ( .A(n19882), .B(n19881), .Z(n19987) );
  NOR U20199 ( .A(n19883), .B(n19987), .Z(n19884) );
  NOR U20200 ( .A(n19885), .B(n19884), .Z(n19888) );
  NOR U20201 ( .A(n161), .B(n63), .Z(n19887) );
  IV U20202 ( .A(n19887), .Z(n19886) );
  NOR U20203 ( .A(n19888), .B(n19886), .Z(n19900) );
  XOR U20204 ( .A(n19888), .B(n19887), .Z(n20469) );
  NOR U20205 ( .A(n158), .B(n62), .Z(n19889) );
  IV U20206 ( .A(n19889), .Z(n19905) );
  IV U20207 ( .A(n19890), .Z(n19891) );
  NOR U20208 ( .A(n19892), .B(n19891), .Z(n19896) );
  NOR U20209 ( .A(n19894), .B(n19893), .Z(n19895) );
  NOR U20210 ( .A(n19896), .B(n19895), .Z(n19903) );
  XOR U20211 ( .A(n19898), .B(n19897), .Z(n19902) );
  XOR U20212 ( .A(n19903), .B(n19902), .Z(n19904) );
  XOR U20213 ( .A(n19905), .B(n19904), .Z(n20470) );
  NOR U20214 ( .A(n20469), .B(n20470), .Z(n19899) );
  NOR U20215 ( .A(n19900), .B(n19899), .Z(n19913) );
  NOR U20216 ( .A(n163), .B(n63), .Z(n19912) );
  IV U20217 ( .A(n19912), .Z(n19901) );
  NOR U20218 ( .A(n19913), .B(n19901), .Z(n19915) );
  NOR U20219 ( .A(n161), .B(n62), .Z(n19920) );
  NOR U20220 ( .A(n19903), .B(n19902), .Z(n19908) );
  IV U20221 ( .A(n19904), .Z(n19906) );
  NOR U20222 ( .A(n19906), .B(n19905), .Z(n19907) );
  NOR U20223 ( .A(n19908), .B(n19907), .Z(n19919) );
  IV U20224 ( .A(n19919), .Z(n19911) );
  XOR U20225 ( .A(n19910), .B(n19909), .Z(n19918) );
  XOR U20226 ( .A(n19911), .B(n19918), .Z(n19922) );
  XOR U20227 ( .A(n19920), .B(n19922), .Z(n19983) );
  XOR U20228 ( .A(n19913), .B(n19912), .Z(n19984) );
  NOR U20229 ( .A(n19983), .B(n19984), .Z(n19914) );
  NOR U20230 ( .A(n19915), .B(n19914), .Z(n19926) );
  XOR U20231 ( .A(n19917), .B(n19916), .Z(n19937) );
  NOR U20232 ( .A(n19919), .B(n19918), .Z(n19924) );
  IV U20233 ( .A(n19920), .Z(n19921) );
  NOR U20234 ( .A(n19922), .B(n19921), .Z(n19923) );
  NOR U20235 ( .A(n19924), .B(n19923), .Z(n19936) );
  NOR U20236 ( .A(n163), .B(n62), .Z(n19934) );
  XOR U20237 ( .A(n19936), .B(n19934), .Z(n19938) );
  XOR U20238 ( .A(n19937), .B(n19938), .Z(n19925) );
  NOR U20239 ( .A(n19926), .B(n19925), .Z(n19930) );
  XOR U20240 ( .A(n19926), .B(n19925), .Z(n19980) );
  IV U20241 ( .A(n19980), .Z(n19928) );
  NOR U20242 ( .A(n165), .B(n63), .Z(n19927) );
  IV U20243 ( .A(n19927), .Z(n19981) );
  NOR U20244 ( .A(n19928), .B(n19981), .Z(n19929) );
  NOR U20245 ( .A(n19930), .B(n19929), .Z(n19933) );
  NOR U20246 ( .A(n167), .B(n63), .Z(n19932) );
  IV U20247 ( .A(n19932), .Z(n19931) );
  NOR U20248 ( .A(n19933), .B(n19931), .Z(n19946) );
  XOR U20249 ( .A(n19933), .B(n19932), .Z(n20485) );
  NOR U20250 ( .A(n165), .B(n62), .Z(n19952) );
  IV U20251 ( .A(n19934), .Z(n19935) );
  NOR U20252 ( .A(n19936), .B(n19935), .Z(n19941) );
  IV U20253 ( .A(n19937), .Z(n19939) );
  NOR U20254 ( .A(n19939), .B(n19938), .Z(n19940) );
  NOR U20255 ( .A(n19941), .B(n19940), .Z(n19950) );
  XOR U20256 ( .A(n19943), .B(n19942), .Z(n19949) );
  XOR U20257 ( .A(n19950), .B(n19949), .Z(n19951) );
  XOR U20258 ( .A(n19952), .B(n19951), .Z(n20486) );
  IV U20259 ( .A(n20486), .Z(n19944) );
  NOR U20260 ( .A(n20485), .B(n19944), .Z(n19945) );
  NOR U20261 ( .A(n19946), .B(n19945), .Z(n20488) );
  XOR U20262 ( .A(n19948), .B(n19947), .Z(n19961) );
  NOR U20263 ( .A(n167), .B(n62), .Z(n19958) );
  NOR U20264 ( .A(n19950), .B(n19949), .Z(n19956) );
  IV U20265 ( .A(n19951), .Z(n19954) );
  IV U20266 ( .A(n19952), .Z(n19953) );
  NOR U20267 ( .A(n19954), .B(n19953), .Z(n19955) );
  NOR U20268 ( .A(n19956), .B(n19955), .Z(n19960) );
  XOR U20269 ( .A(n19958), .B(n19960), .Z(n19962) );
  XOR U20270 ( .A(n19961), .B(n19962), .Z(n20487) );
  IV U20271 ( .A(n20487), .Z(n19957) );
  NOR U20272 ( .A(n20488), .B(n19957), .Z(n19979) );
  IV U20273 ( .A(n19979), .Z(n31558) );
  IV U20274 ( .A(n19958), .Z(n19959) );
  NOR U20275 ( .A(n19960), .B(n19959), .Z(n19964) );
  NOR U20276 ( .A(n19962), .B(n19961), .Z(n19963) );
  NOR U20277 ( .A(n19964), .B(n19963), .Z(n19971) );
  IV U20278 ( .A(n19965), .Z(n19967) );
  XOR U20279 ( .A(n19967), .B(n19966), .Z(n19970) );
  XOR U20280 ( .A(n19971), .B(n19970), .Z(n31557) );
  IV U20281 ( .A(n31557), .Z(n19968) );
  NOR U20282 ( .A(n31558), .B(n19968), .Z(n31561) );
  IV U20283 ( .A(n31561), .Z(n19969) );
  NOR U20284 ( .A(n19972), .B(n19969), .Z(n19973) );
  NOR U20285 ( .A(n19971), .B(n19970), .Z(n19978) );
  IV U20286 ( .A(n19978), .Z(n31575) );
  NOR U20287 ( .A(n31575), .B(n19972), .Z(n31567) );
  NOR U20288 ( .A(n19973), .B(n31567), .Z(n19974) );
  IV U20289 ( .A(n19974), .Z(n19975) );
  NOR U20290 ( .A(n19976), .B(n19975), .Z(n19977) );
  IV U20291 ( .A(n19977), .Z(n28555) );
  NOR U20292 ( .A(n19978), .B(n31563), .Z(n28553) );
  NOR U20293 ( .A(n19979), .B(n31557), .Z(n28552) );
  XOR U20294 ( .A(n19981), .B(n19980), .Z(n20481) );
  NOR U20295 ( .A(n167), .B(n64), .Z(n20482) );
  IV U20296 ( .A(n20482), .Z(n19982) );
  NOR U20297 ( .A(n20481), .B(n19982), .Z(n20484) );
  IV U20298 ( .A(n19983), .Z(n19985) );
  XOR U20299 ( .A(n19985), .B(n19984), .Z(n20477) );
  NOR U20300 ( .A(n165), .B(n64), .Z(n20478) );
  IV U20301 ( .A(n20478), .Z(n19986) );
  NOR U20302 ( .A(n20477), .B(n19986), .Z(n20480) );
  XOR U20303 ( .A(n19988), .B(n19987), .Z(n20465) );
  NOR U20304 ( .A(n161), .B(n64), .Z(n20466) );
  IV U20305 ( .A(n20466), .Z(n19989) );
  NOR U20306 ( .A(n20465), .B(n19989), .Z(n20468) );
  XOR U20307 ( .A(n19991), .B(n19990), .Z(n19992) );
  XOR U20308 ( .A(n19993), .B(n19992), .Z(n20461) );
  NOR U20309 ( .A(n158), .B(n64), .Z(n20462) );
  IV U20310 ( .A(n20462), .Z(n19994) );
  NOR U20311 ( .A(n20461), .B(n19994), .Z(n20464) );
  XOR U20312 ( .A(n19996), .B(n19995), .Z(n19997) );
  XOR U20313 ( .A(n19998), .B(n19997), .Z(n20449) );
  NOR U20314 ( .A(n155), .B(n64), .Z(n20450) );
  IV U20315 ( .A(n20450), .Z(n19999) );
  NOR U20316 ( .A(n20449), .B(n19999), .Z(n20452) );
  IV U20317 ( .A(n20000), .Z(n20002) );
  XOR U20318 ( .A(n20002), .B(n20001), .Z(n20445) );
  NOR U20319 ( .A(n153), .B(n64), .Z(n20446) );
  IV U20320 ( .A(n20446), .Z(n20003) );
  NOR U20321 ( .A(n20445), .B(n20003), .Z(n20448) );
  NOR U20322 ( .A(n147), .B(n64), .Z(n20006) );
  XOR U20323 ( .A(n20005), .B(n20004), .Z(n20007) );
  NOR U20324 ( .A(n20006), .B(n20007), .Z(n20426) );
  IV U20325 ( .A(n20006), .Z(n20008) );
  XOR U20326 ( .A(n20008), .B(n20007), .Z(n20491) );
  XOR U20327 ( .A(n20010), .B(n20009), .Z(n20403) );
  NOR U20328 ( .A(n141), .B(n64), .Z(n20404) );
  IV U20329 ( .A(n20404), .Z(n20011) );
  NOR U20330 ( .A(n20403), .B(n20011), .Z(n20406) );
  NOR U20331 ( .A(n137), .B(n64), .Z(n20392) );
  IV U20332 ( .A(n20392), .Z(n20014) );
  XOR U20333 ( .A(n20013), .B(n20012), .Z(n20391) );
  NOR U20334 ( .A(n20014), .B(n20391), .Z(n20394) );
  NOR U20335 ( .A(n135), .B(n64), .Z(n20015) );
  IV U20336 ( .A(n20015), .Z(n20385) );
  NOR U20337 ( .A(n133), .B(n64), .Z(n20018) );
  XOR U20338 ( .A(n20017), .B(n20016), .Z(n20019) );
  NOR U20339 ( .A(n20018), .B(n20019), .Z(n20382) );
  IV U20340 ( .A(n20018), .Z(n20865) );
  IV U20341 ( .A(n20019), .Z(n20864) );
  NOR U20342 ( .A(n20865), .B(n20864), .Z(n20380) );
  XOR U20343 ( .A(n20021), .B(n20020), .Z(n20023) );
  IV U20344 ( .A(n20023), .Z(n20505) );
  NOR U20345 ( .A(n128), .B(n64), .Z(n20022) );
  IV U20346 ( .A(n20022), .Z(n20504) );
  NOR U20347 ( .A(n20505), .B(n20504), .Z(n20369) );
  NOR U20348 ( .A(n20023), .B(n20022), .Z(n20367) );
  XOR U20349 ( .A(n20025), .B(n20024), .Z(n20026) );
  XOR U20350 ( .A(n20027), .B(n20026), .Z(n20364) );
  NOR U20351 ( .A(n126), .B(n64), .Z(n20363) );
  IV U20352 ( .A(n20363), .Z(n20028) );
  NOR U20353 ( .A(n20364), .B(n20028), .Z(n20366) );
  NOR U20354 ( .A(n125), .B(n64), .Z(n20029) );
  IV U20355 ( .A(n20029), .Z(n20359) );
  IV U20356 ( .A(n20030), .Z(n20032) );
  XOR U20357 ( .A(n20032), .B(n20031), .Z(n20358) );
  NOR U20358 ( .A(n20359), .B(n20358), .Z(n20362) );
  NOR U20359 ( .A(n120), .B(n64), .Z(n20035) );
  XOR U20360 ( .A(n20034), .B(n20033), .Z(n20036) );
  NOR U20361 ( .A(n20035), .B(n20036), .Z(n20347) );
  IV U20362 ( .A(n20035), .Z(n20519) );
  IV U20363 ( .A(n20036), .Z(n20518) );
  NOR U20364 ( .A(n20519), .B(n20518), .Z(n20345) );
  XOR U20365 ( .A(n20038), .B(n20037), .Z(n20039) );
  XOR U20366 ( .A(n20040), .B(n20039), .Z(n20341) );
  NOR U20367 ( .A(n119), .B(n64), .Z(n20340) );
  IV U20368 ( .A(n20340), .Z(n20041) );
  NOR U20369 ( .A(n20341), .B(n20041), .Z(n20343) );
  NOR U20370 ( .A(n79), .B(n64), .Z(n20335) );
  XOR U20371 ( .A(n20043), .B(n20042), .Z(n20334) );
  NOR U20372 ( .A(n20335), .B(n20334), .Z(n20338) );
  XOR U20373 ( .A(n20045), .B(n20044), .Z(n20330) );
  NOR U20374 ( .A(n117), .B(n64), .Z(n20329) );
  IV U20375 ( .A(n20329), .Z(n20046) );
  NOR U20376 ( .A(n20330), .B(n20046), .Z(n20332) );
  NOR U20377 ( .A(n80), .B(n64), .Z(n20324) );
  XOR U20378 ( .A(n20048), .B(n20047), .Z(n20323) );
  NOR U20379 ( .A(n20324), .B(n20323), .Z(n20327) );
  XOR U20380 ( .A(n20050), .B(n20049), .Z(n20319) );
  NOR U20381 ( .A(n116), .B(n64), .Z(n20318) );
  IV U20382 ( .A(n20318), .Z(n20051) );
  NOR U20383 ( .A(n20319), .B(n20051), .Z(n20321) );
  NOR U20384 ( .A(n81), .B(n64), .Z(n20313) );
  XOR U20385 ( .A(n20053), .B(n20052), .Z(n20312) );
  NOR U20386 ( .A(n20313), .B(n20312), .Z(n20316) );
  XOR U20387 ( .A(n20055), .B(n20054), .Z(n20308) );
  NOR U20388 ( .A(n115), .B(n64), .Z(n20307) );
  IV U20389 ( .A(n20307), .Z(n20056) );
  NOR U20390 ( .A(n20308), .B(n20056), .Z(n20310) );
  NOR U20391 ( .A(n82), .B(n64), .Z(n20302) );
  XOR U20392 ( .A(n20058), .B(n20057), .Z(n20301) );
  NOR U20393 ( .A(n20302), .B(n20301), .Z(n20305) );
  XOR U20394 ( .A(n20060), .B(n20059), .Z(n20297) );
  NOR U20395 ( .A(n114), .B(n64), .Z(n20296) );
  IV U20396 ( .A(n20296), .Z(n20061) );
  NOR U20397 ( .A(n20297), .B(n20061), .Z(n20299) );
  NOR U20398 ( .A(n83), .B(n64), .Z(n20065) );
  XOR U20399 ( .A(n20063), .B(n20062), .Z(n20064) );
  NOR U20400 ( .A(n20065), .B(n20064), .Z(n20294) );
  XOR U20401 ( .A(n20065), .B(n20064), .Z(n20066) );
  IV U20402 ( .A(n20066), .Z(n20546) );
  XOR U20403 ( .A(n20068), .B(n20067), .Z(n20289) );
  NOR U20404 ( .A(n113), .B(n64), .Z(n20288) );
  IV U20405 ( .A(n20288), .Z(n20069) );
  NOR U20406 ( .A(n20289), .B(n20069), .Z(n20291) );
  NOR U20407 ( .A(n84), .B(n64), .Z(n20283) );
  XOR U20408 ( .A(n20071), .B(n20070), .Z(n20282) );
  NOR U20409 ( .A(n20283), .B(n20282), .Z(n20286) );
  XOR U20410 ( .A(n20073), .B(n20072), .Z(n20278) );
  NOR U20411 ( .A(n112), .B(n64), .Z(n20277) );
  IV U20412 ( .A(n20277), .Z(n20074) );
  NOR U20413 ( .A(n20278), .B(n20074), .Z(n20280) );
  IV U20414 ( .A(n20075), .Z(n20077) );
  XOR U20415 ( .A(n20077), .B(n20076), .Z(n20273) );
  NOR U20416 ( .A(n85), .B(n64), .Z(n20274) );
  IV U20417 ( .A(n20274), .Z(n20078) );
  NOR U20418 ( .A(n20273), .B(n20078), .Z(n20276) );
  IV U20419 ( .A(n20079), .Z(n20081) );
  XOR U20420 ( .A(n20081), .B(n20080), .Z(n20269) );
  NOR U20421 ( .A(n111), .B(n64), .Z(n20270) );
  IV U20422 ( .A(n20270), .Z(n20082) );
  NOR U20423 ( .A(n20269), .B(n20082), .Z(n20272) );
  IV U20424 ( .A(n20083), .Z(n20085) );
  XOR U20425 ( .A(n20085), .B(n20084), .Z(n20265) );
  NOR U20426 ( .A(n86), .B(n64), .Z(n20266) );
  IV U20427 ( .A(n20266), .Z(n20086) );
  NOR U20428 ( .A(n20265), .B(n20086), .Z(n20268) );
  IV U20429 ( .A(n20087), .Z(n20089) );
  XOR U20430 ( .A(n20089), .B(n20088), .Z(n20260) );
  NOR U20431 ( .A(n110), .B(n64), .Z(n20261) );
  IV U20432 ( .A(n20261), .Z(n20090) );
  NOR U20433 ( .A(n20260), .B(n20090), .Z(n20264) );
  NOR U20434 ( .A(n109), .B(n64), .Z(n20256) );
  XOR U20435 ( .A(n20092), .B(n20091), .Z(n20255) );
  NOR U20436 ( .A(n20256), .B(n20255), .Z(n20259) );
  IV U20437 ( .A(n20093), .Z(n20095) );
  XOR U20438 ( .A(n20095), .B(n20094), .Z(n20242) );
  NOR U20439 ( .A(n87), .B(n64), .Z(n20243) );
  IV U20440 ( .A(n20243), .Z(n20096) );
  NOR U20441 ( .A(n20242), .B(n20096), .Z(n20245) );
  IV U20442 ( .A(n20097), .Z(n20099) );
  XOR U20443 ( .A(n20099), .B(n20098), .Z(n20238) );
  NOR U20444 ( .A(n107), .B(n64), .Z(n20239) );
  IV U20445 ( .A(n20239), .Z(n20100) );
  NOR U20446 ( .A(n20238), .B(n20100), .Z(n20241) );
  IV U20447 ( .A(n20101), .Z(n20103) );
  XOR U20448 ( .A(n20103), .B(n20102), .Z(n20234) );
  NOR U20449 ( .A(n88), .B(n64), .Z(n20235) );
  IV U20450 ( .A(n20235), .Z(n20104) );
  NOR U20451 ( .A(n20234), .B(n20104), .Z(n20237) );
  IV U20452 ( .A(n20105), .Z(n20107) );
  XOR U20453 ( .A(n20107), .B(n20106), .Z(n20230) );
  NOR U20454 ( .A(n106), .B(n64), .Z(n20231) );
  IV U20455 ( .A(n20231), .Z(n20108) );
  NOR U20456 ( .A(n20230), .B(n20108), .Z(n20233) );
  XOR U20457 ( .A(n20110), .B(n20109), .Z(n20226) );
  NOR U20458 ( .A(n105), .B(n64), .Z(n20227) );
  IV U20459 ( .A(n20227), .Z(n20111) );
  NOR U20460 ( .A(n20226), .B(n20111), .Z(n20229) );
  XOR U20461 ( .A(n20113), .B(n20112), .Z(n20214) );
  IV U20462 ( .A(n20214), .Z(n20115) );
  NOR U20463 ( .A(n89), .B(n64), .Z(n20114) );
  IV U20464 ( .A(n20114), .Z(n20215) );
  NOR U20465 ( .A(n20115), .B(n20215), .Z(n20217) );
  IV U20466 ( .A(n20116), .Z(n20118) );
  XOR U20467 ( .A(n20118), .B(n20117), .Z(n20210) );
  NOR U20468 ( .A(n103), .B(n64), .Z(n20211) );
  IV U20469 ( .A(n20211), .Z(n20119) );
  NOR U20470 ( .A(n20210), .B(n20119), .Z(n20213) );
  IV U20471 ( .A(n20120), .Z(n20122) );
  XOR U20472 ( .A(n20122), .B(n20121), .Z(n20206) );
  NOR U20473 ( .A(n90), .B(n64), .Z(n20207) );
  IV U20474 ( .A(n20207), .Z(n20123) );
  NOR U20475 ( .A(n20206), .B(n20123), .Z(n20209) );
  IV U20476 ( .A(n20124), .Z(n20126) );
  XOR U20477 ( .A(n20126), .B(n20125), .Z(n20202) );
  NOR U20478 ( .A(n102), .B(n64), .Z(n20203) );
  IV U20479 ( .A(n20203), .Z(n20127) );
  NOR U20480 ( .A(n20202), .B(n20127), .Z(n20205) );
  IV U20481 ( .A(n20128), .Z(n20130) );
  XOR U20482 ( .A(n20130), .B(n20129), .Z(n20198) );
  NOR U20483 ( .A(n101), .B(n64), .Z(n20199) );
  IV U20484 ( .A(n20199), .Z(n20131) );
  NOR U20485 ( .A(n20198), .B(n20131), .Z(n20201) );
  IV U20486 ( .A(n20132), .Z(n20134) );
  XOR U20487 ( .A(n20134), .B(n20133), .Z(n20194) );
  NOR U20488 ( .A(n100), .B(n64), .Z(n20195) );
  IV U20489 ( .A(n20195), .Z(n20135) );
  NOR U20490 ( .A(n20194), .B(n20135), .Z(n20197) );
  IV U20491 ( .A(n20136), .Z(n20138) );
  XOR U20492 ( .A(n20138), .B(n20137), .Z(n20190) );
  NOR U20493 ( .A(n99), .B(n64), .Z(n20191) );
  IV U20494 ( .A(n20191), .Z(n20139) );
  NOR U20495 ( .A(n20190), .B(n20139), .Z(n20193) );
  IV U20496 ( .A(n20140), .Z(n20142) );
  XOR U20497 ( .A(n20142), .B(n20141), .Z(n20186) );
  NOR U20498 ( .A(n98), .B(n64), .Z(n20187) );
  IV U20499 ( .A(n20187), .Z(n20143) );
  NOR U20500 ( .A(n20186), .B(n20143), .Z(n20189) );
  XOR U20501 ( .A(n20145), .B(n20144), .Z(n20182) );
  NOR U20502 ( .A(n91), .B(n64), .Z(n20183) );
  IV U20503 ( .A(n20183), .Z(n20146) );
  NOR U20504 ( .A(n20182), .B(n20146), .Z(n20185) );
  IV U20505 ( .A(n20147), .Z(n20149) );
  XOR U20506 ( .A(n20149), .B(n20148), .Z(n20178) );
  NOR U20507 ( .A(n97), .B(n64), .Z(n20179) );
  IV U20508 ( .A(n20179), .Z(n20150) );
  NOR U20509 ( .A(n20178), .B(n20150), .Z(n20181) );
  XOR U20510 ( .A(n20152), .B(n20151), .Z(n20174) );
  IV U20511 ( .A(n20174), .Z(n20154) );
  NOR U20512 ( .A(n96), .B(n64), .Z(n20153) );
  IV U20513 ( .A(n20153), .Z(n20175) );
  NOR U20514 ( .A(n20154), .B(n20175), .Z(n20177) );
  NOR U20515 ( .A(n95), .B(n64), .Z(n20171) );
  IV U20516 ( .A(n20171), .Z(n20157) );
  XOR U20517 ( .A(n20156), .B(n20155), .Z(n20170) );
  NOR U20518 ( .A(n20157), .B(n20170), .Z(n20173) );
  NOR U20519 ( .A(n64), .B(n93), .Z(n21148) );
  IV U20520 ( .A(n21148), .Z(n20158) );
  NOR U20521 ( .A(n63), .B(n168), .Z(n20166) );
  IV U20522 ( .A(n20166), .Z(n20161) );
  NOR U20523 ( .A(n20158), .B(n20161), .Z(n20159) );
  IV U20524 ( .A(n20159), .Z(n20160) );
  NOR U20525 ( .A(n94), .B(n20160), .Z(n20169) );
  NOR U20526 ( .A(n20161), .B(n93), .Z(n20162) );
  XOR U20527 ( .A(n94), .B(n20162), .Z(n20163) );
  NOR U20528 ( .A(n64), .B(n20163), .Z(n20164) );
  IV U20529 ( .A(n20164), .Z(n20640) );
  XOR U20530 ( .A(n20166), .B(n20165), .Z(n20639) );
  IV U20531 ( .A(n20639), .Z(n20167) );
  NOR U20532 ( .A(n20640), .B(n20167), .Z(n20168) );
  NOR U20533 ( .A(n20169), .B(n20168), .Z(n20636) );
  XOR U20534 ( .A(n20171), .B(n20170), .Z(n20635) );
  NOR U20535 ( .A(n20636), .B(n20635), .Z(n20172) );
  NOR U20536 ( .A(n20173), .B(n20172), .Z(n20663) );
  XOR U20537 ( .A(n20175), .B(n20174), .Z(n20662) );
  NOR U20538 ( .A(n20663), .B(n20662), .Z(n20176) );
  NOR U20539 ( .A(n20177), .B(n20176), .Z(n20631) );
  XOR U20540 ( .A(n20179), .B(n20178), .Z(n20632) );
  NOR U20541 ( .A(n20631), .B(n20632), .Z(n20180) );
  NOR U20542 ( .A(n20181), .B(n20180), .Z(n20627) );
  XOR U20543 ( .A(n20183), .B(n20182), .Z(n20628) );
  NOR U20544 ( .A(n20627), .B(n20628), .Z(n20184) );
  NOR U20545 ( .A(n20185), .B(n20184), .Z(n20623) );
  XOR U20546 ( .A(n20187), .B(n20186), .Z(n20624) );
  NOR U20547 ( .A(n20623), .B(n20624), .Z(n20188) );
  NOR U20548 ( .A(n20189), .B(n20188), .Z(n20619) );
  XOR U20549 ( .A(n20191), .B(n20190), .Z(n20620) );
  NOR U20550 ( .A(n20619), .B(n20620), .Z(n20192) );
  NOR U20551 ( .A(n20193), .B(n20192), .Z(n20615) );
  XOR U20552 ( .A(n20195), .B(n20194), .Z(n20616) );
  NOR U20553 ( .A(n20615), .B(n20616), .Z(n20196) );
  NOR U20554 ( .A(n20197), .B(n20196), .Z(n20611) );
  XOR U20555 ( .A(n20199), .B(n20198), .Z(n20612) );
  NOR U20556 ( .A(n20611), .B(n20612), .Z(n20200) );
  NOR U20557 ( .A(n20201), .B(n20200), .Z(n20607) );
  XOR U20558 ( .A(n20203), .B(n20202), .Z(n20608) );
  NOR U20559 ( .A(n20607), .B(n20608), .Z(n20204) );
  NOR U20560 ( .A(n20205), .B(n20204), .Z(n20603) );
  XOR U20561 ( .A(n20207), .B(n20206), .Z(n20604) );
  NOR U20562 ( .A(n20603), .B(n20604), .Z(n20208) );
  NOR U20563 ( .A(n20209), .B(n20208), .Z(n20600) );
  XOR U20564 ( .A(n20211), .B(n20210), .Z(n20599) );
  NOR U20565 ( .A(n20600), .B(n20599), .Z(n20212) );
  NOR U20566 ( .A(n20213), .B(n20212), .Z(n20707) );
  XOR U20567 ( .A(n20215), .B(n20214), .Z(n20706) );
  NOR U20568 ( .A(n20707), .B(n20706), .Z(n20216) );
  NOR U20569 ( .A(n20217), .B(n20216), .Z(n20222) );
  XOR U20570 ( .A(n20219), .B(n20218), .Z(n20221) );
  IV U20571 ( .A(n20221), .Z(n20220) );
  NOR U20572 ( .A(n20222), .B(n20220), .Z(n20225) );
  XOR U20573 ( .A(n20222), .B(n20221), .Z(n20596) );
  NOR U20574 ( .A(n104), .B(n64), .Z(n20597) );
  IV U20575 ( .A(n20597), .Z(n20223) );
  NOR U20576 ( .A(n20596), .B(n20223), .Z(n20224) );
  NOR U20577 ( .A(n20225), .B(n20224), .Z(n20592) );
  XOR U20578 ( .A(n20227), .B(n20226), .Z(n20593) );
  NOR U20579 ( .A(n20592), .B(n20593), .Z(n20228) );
  NOR U20580 ( .A(n20229), .B(n20228), .Z(n20588) );
  XOR U20581 ( .A(n20231), .B(n20230), .Z(n20589) );
  NOR U20582 ( .A(n20588), .B(n20589), .Z(n20232) );
  NOR U20583 ( .A(n20233), .B(n20232), .Z(n20584) );
  XOR U20584 ( .A(n20235), .B(n20234), .Z(n20585) );
  NOR U20585 ( .A(n20584), .B(n20585), .Z(n20236) );
  NOR U20586 ( .A(n20237), .B(n20236), .Z(n20581) );
  XOR U20587 ( .A(n20239), .B(n20238), .Z(n20580) );
  NOR U20588 ( .A(n20581), .B(n20580), .Z(n20240) );
  NOR U20589 ( .A(n20241), .B(n20240), .Z(n20576) );
  XOR U20590 ( .A(n20243), .B(n20242), .Z(n20577) );
  NOR U20591 ( .A(n20576), .B(n20577), .Z(n20244) );
  NOR U20592 ( .A(n20245), .B(n20244), .Z(n20248) );
  NOR U20593 ( .A(n108), .B(n64), .Z(n20247) );
  IV U20594 ( .A(n20247), .Z(n20246) );
  NOR U20595 ( .A(n20248), .B(n20246), .Z(n20253) );
  XOR U20596 ( .A(n20248), .B(n20247), .Z(n20573) );
  XOR U20597 ( .A(n20250), .B(n20249), .Z(n20574) );
  IV U20598 ( .A(n20574), .Z(n20251) );
  NOR U20599 ( .A(n20573), .B(n20251), .Z(n20252) );
  NOR U20600 ( .A(n20253), .B(n20252), .Z(n20254) );
  IV U20601 ( .A(n20254), .Z(n20571) );
  XOR U20602 ( .A(n20256), .B(n20255), .Z(n20257) );
  IV U20603 ( .A(n20257), .Z(n20570) );
  NOR U20604 ( .A(n20571), .B(n20570), .Z(n20258) );
  NOR U20605 ( .A(n20259), .B(n20258), .Z(n20568) );
  IV U20606 ( .A(n20568), .Z(n20262) );
  XOR U20607 ( .A(n20261), .B(n20260), .Z(n20567) );
  NOR U20608 ( .A(n20262), .B(n20567), .Z(n20263) );
  NOR U20609 ( .A(n20264), .B(n20263), .Z(n20563) );
  XOR U20610 ( .A(n20266), .B(n20265), .Z(n20564) );
  NOR U20611 ( .A(n20563), .B(n20564), .Z(n20267) );
  NOR U20612 ( .A(n20268), .B(n20267), .Z(n20559) );
  XOR U20613 ( .A(n20270), .B(n20269), .Z(n20560) );
  NOR U20614 ( .A(n20559), .B(n20560), .Z(n20271) );
  NOR U20615 ( .A(n20272), .B(n20271), .Z(n20555) );
  XOR U20616 ( .A(n20274), .B(n20273), .Z(n20556) );
  NOR U20617 ( .A(n20555), .B(n20556), .Z(n20275) );
  NOR U20618 ( .A(n20276), .B(n20275), .Z(n20554) );
  XOR U20619 ( .A(n20278), .B(n20277), .Z(n20553) );
  NOR U20620 ( .A(n20554), .B(n20553), .Z(n20279) );
  NOR U20621 ( .A(n20280), .B(n20279), .Z(n20281) );
  IV U20622 ( .A(n20281), .Z(n20551) );
  XOR U20623 ( .A(n20283), .B(n20282), .Z(n20284) );
  IV U20624 ( .A(n20284), .Z(n20550) );
  NOR U20625 ( .A(n20551), .B(n20550), .Z(n20285) );
  NOR U20626 ( .A(n20286), .B(n20285), .Z(n20287) );
  IV U20627 ( .A(n20287), .Z(n20549) );
  XOR U20628 ( .A(n20289), .B(n20288), .Z(n20548) );
  NOR U20629 ( .A(n20549), .B(n20548), .Z(n20290) );
  NOR U20630 ( .A(n20291), .B(n20290), .Z(n20292) );
  IV U20631 ( .A(n20292), .Z(n20545) );
  NOR U20632 ( .A(n20546), .B(n20545), .Z(n20293) );
  NOR U20633 ( .A(n20294), .B(n20293), .Z(n20295) );
  IV U20634 ( .A(n20295), .Z(n20544) );
  XOR U20635 ( .A(n20297), .B(n20296), .Z(n20543) );
  NOR U20636 ( .A(n20544), .B(n20543), .Z(n20298) );
  NOR U20637 ( .A(n20299), .B(n20298), .Z(n20300) );
  IV U20638 ( .A(n20300), .Z(n20541) );
  XOR U20639 ( .A(n20302), .B(n20301), .Z(n20303) );
  IV U20640 ( .A(n20303), .Z(n20540) );
  NOR U20641 ( .A(n20541), .B(n20540), .Z(n20304) );
  NOR U20642 ( .A(n20305), .B(n20304), .Z(n20306) );
  IV U20643 ( .A(n20306), .Z(n20539) );
  XOR U20644 ( .A(n20308), .B(n20307), .Z(n20538) );
  NOR U20645 ( .A(n20539), .B(n20538), .Z(n20309) );
  NOR U20646 ( .A(n20310), .B(n20309), .Z(n20311) );
  IV U20647 ( .A(n20311), .Z(n20536) );
  XOR U20648 ( .A(n20313), .B(n20312), .Z(n20314) );
  IV U20649 ( .A(n20314), .Z(n20535) );
  NOR U20650 ( .A(n20536), .B(n20535), .Z(n20315) );
  NOR U20651 ( .A(n20316), .B(n20315), .Z(n20317) );
  IV U20652 ( .A(n20317), .Z(n20534) );
  XOR U20653 ( .A(n20319), .B(n20318), .Z(n20533) );
  NOR U20654 ( .A(n20534), .B(n20533), .Z(n20320) );
  NOR U20655 ( .A(n20321), .B(n20320), .Z(n20322) );
  IV U20656 ( .A(n20322), .Z(n20531) );
  XOR U20657 ( .A(n20324), .B(n20323), .Z(n20325) );
  IV U20658 ( .A(n20325), .Z(n20530) );
  NOR U20659 ( .A(n20531), .B(n20530), .Z(n20326) );
  NOR U20660 ( .A(n20327), .B(n20326), .Z(n20328) );
  IV U20661 ( .A(n20328), .Z(n20529) );
  XOR U20662 ( .A(n20330), .B(n20329), .Z(n20528) );
  NOR U20663 ( .A(n20529), .B(n20528), .Z(n20331) );
  NOR U20664 ( .A(n20332), .B(n20331), .Z(n20333) );
  IV U20665 ( .A(n20333), .Z(n20526) );
  XOR U20666 ( .A(n20335), .B(n20334), .Z(n20336) );
  IV U20667 ( .A(n20336), .Z(n20525) );
  NOR U20668 ( .A(n20526), .B(n20525), .Z(n20337) );
  NOR U20669 ( .A(n20338), .B(n20337), .Z(n20339) );
  IV U20670 ( .A(n20339), .Z(n20524) );
  XOR U20671 ( .A(n20341), .B(n20340), .Z(n20523) );
  NOR U20672 ( .A(n20524), .B(n20523), .Z(n20342) );
  NOR U20673 ( .A(n20343), .B(n20342), .Z(n20521) );
  IV U20674 ( .A(n20521), .Z(n20344) );
  NOR U20675 ( .A(n20345), .B(n20344), .Z(n20346) );
  NOR U20676 ( .A(n20347), .B(n20346), .Z(n20348) );
  IV U20677 ( .A(n20348), .Z(n20355) );
  NOR U20678 ( .A(n123), .B(n64), .Z(n20354) );
  IV U20679 ( .A(n20354), .Z(n20349) );
  NOR U20680 ( .A(n20355), .B(n20349), .Z(n20357) );
  XOR U20681 ( .A(n20351), .B(n20350), .Z(n20352) );
  XOR U20682 ( .A(n20353), .B(n20352), .Z(n20514) );
  XOR U20683 ( .A(n20355), .B(n20354), .Z(n20515) );
  NOR U20684 ( .A(n20514), .B(n20515), .Z(n20356) );
  NOR U20685 ( .A(n20357), .B(n20356), .Z(n20846) );
  XOR U20686 ( .A(n20359), .B(n20358), .Z(n20847) );
  IV U20687 ( .A(n20847), .Z(n20360) );
  NOR U20688 ( .A(n20846), .B(n20360), .Z(n20361) );
  NOR U20689 ( .A(n20362), .B(n20361), .Z(n20510) );
  XOR U20690 ( .A(n20364), .B(n20363), .Z(n20509) );
  NOR U20691 ( .A(n20510), .B(n20509), .Z(n20365) );
  NOR U20692 ( .A(n20366), .B(n20365), .Z(n20507) );
  NOR U20693 ( .A(n20367), .B(n20507), .Z(n20368) );
  NOR U20694 ( .A(n20369), .B(n20368), .Z(n20375) );
  NOR U20695 ( .A(n131), .B(n64), .Z(n20376) );
  IV U20696 ( .A(n20376), .Z(n20370) );
  NOR U20697 ( .A(n20375), .B(n20370), .Z(n20378) );
  XOR U20698 ( .A(n20372), .B(n20371), .Z(n20373) );
  XOR U20699 ( .A(n20374), .B(n20373), .Z(n20501) );
  XOR U20700 ( .A(n20376), .B(n20375), .Z(n20500) );
  NOR U20701 ( .A(n20501), .B(n20500), .Z(n20377) );
  NOR U20702 ( .A(n20378), .B(n20377), .Z(n20867) );
  IV U20703 ( .A(n20867), .Z(n20379) );
  NOR U20704 ( .A(n20380), .B(n20379), .Z(n20381) );
  NOR U20705 ( .A(n20382), .B(n20381), .Z(n20384) );
  IV U20706 ( .A(n20384), .Z(n20383) );
  NOR U20707 ( .A(n20385), .B(n20383), .Z(n20390) );
  XOR U20708 ( .A(n20385), .B(n20384), .Z(n20499) );
  XOR U20709 ( .A(n20387), .B(n20386), .Z(n20498) );
  IV U20710 ( .A(n20498), .Z(n20388) );
  NOR U20711 ( .A(n20499), .B(n20388), .Z(n20389) );
  NOR U20712 ( .A(n20390), .B(n20389), .Z(n20880) );
  XOR U20713 ( .A(n20392), .B(n20391), .Z(n20881) );
  NOR U20714 ( .A(n20880), .B(n20881), .Z(n20393) );
  NOR U20715 ( .A(n20394), .B(n20393), .Z(n20399) );
  XOR U20716 ( .A(n20396), .B(n20395), .Z(n20398) );
  IV U20717 ( .A(n20398), .Z(n20397) );
  NOR U20718 ( .A(n20399), .B(n20397), .Z(n20402) );
  XOR U20719 ( .A(n20399), .B(n20398), .Z(n20886) );
  NOR U20720 ( .A(n139), .B(n64), .Z(n20887) );
  IV U20721 ( .A(n20887), .Z(n20400) );
  NOR U20722 ( .A(n20886), .B(n20400), .Z(n20401) );
  NOR U20723 ( .A(n20402), .B(n20401), .Z(n20894) );
  XOR U20724 ( .A(n20404), .B(n20403), .Z(n20893) );
  NOR U20725 ( .A(n20894), .B(n20893), .Z(n20405) );
  NOR U20726 ( .A(n20406), .B(n20405), .Z(n20409) );
  NOR U20727 ( .A(n143), .B(n64), .Z(n20408) );
  IV U20728 ( .A(n20408), .Z(n20407) );
  NOR U20729 ( .A(n20409), .B(n20407), .Z(n20413) );
  XOR U20730 ( .A(n20409), .B(n20408), .Z(n20493) );
  XOR U20731 ( .A(n20411), .B(n20410), .Z(n20494) );
  NOR U20732 ( .A(n20493), .B(n20494), .Z(n20412) );
  NOR U20733 ( .A(n20413), .B(n20412), .Z(n20419) );
  XOR U20734 ( .A(n20415), .B(n20414), .Z(n20416) );
  XOR U20735 ( .A(n20417), .B(n20416), .Z(n20418) );
  NOR U20736 ( .A(n20419), .B(n20418), .Z(n20423) );
  IV U20737 ( .A(n20418), .Z(n20420) );
  XOR U20738 ( .A(n20420), .B(n20419), .Z(n20907) );
  NOR U20739 ( .A(n145), .B(n64), .Z(n20908) );
  IV U20740 ( .A(n20908), .Z(n20421) );
  NOR U20741 ( .A(n20907), .B(n20421), .Z(n20422) );
  NOR U20742 ( .A(n20423), .B(n20422), .Z(n20424) );
  IV U20743 ( .A(n20424), .Z(n20492) );
  NOR U20744 ( .A(n20491), .B(n20492), .Z(n20425) );
  NOR U20745 ( .A(n20426), .B(n20425), .Z(n20434) );
  IV U20746 ( .A(n20434), .Z(n20428) );
  NOR U20747 ( .A(n148), .B(n64), .Z(n20427) );
  IV U20748 ( .A(n20427), .Z(n20433) );
  NOR U20749 ( .A(n20428), .B(n20433), .Z(n20436) );
  XOR U20750 ( .A(n20430), .B(n20429), .Z(n20431) );
  XOR U20751 ( .A(n20432), .B(n20431), .Z(n20917) );
  XOR U20752 ( .A(n20434), .B(n20433), .Z(n20916) );
  NOR U20753 ( .A(n20917), .B(n20916), .Z(n20435) );
  NOR U20754 ( .A(n20436), .B(n20435), .Z(n20440) );
  XOR U20755 ( .A(n20438), .B(n20437), .Z(n20439) );
  NOR U20756 ( .A(n20440), .B(n20439), .Z(n20444) );
  XOR U20757 ( .A(n20440), .B(n20439), .Z(n20927) );
  IV U20758 ( .A(n20927), .Z(n20442) );
  NOR U20759 ( .A(n150), .B(n64), .Z(n20441) );
  IV U20760 ( .A(n20441), .Z(n20928) );
  NOR U20761 ( .A(n20442), .B(n20928), .Z(n20443) );
  NOR U20762 ( .A(n20444), .B(n20443), .Z(n20932) );
  XOR U20763 ( .A(n20446), .B(n20445), .Z(n20931) );
  NOR U20764 ( .A(n20932), .B(n20931), .Z(n20447) );
  NOR U20765 ( .A(n20448), .B(n20447), .Z(n20943) );
  XOR U20766 ( .A(n20450), .B(n20449), .Z(n20942) );
  NOR U20767 ( .A(n20943), .B(n20942), .Z(n20451) );
  NOR U20768 ( .A(n20452), .B(n20451), .Z(n20456) );
  XOR U20769 ( .A(n20454), .B(n20453), .Z(n20455) );
  NOR U20770 ( .A(n20456), .B(n20455), .Z(n20460) );
  XOR U20771 ( .A(n20456), .B(n20455), .Z(n20457) );
  IV U20772 ( .A(n20457), .Z(n20950) );
  NOR U20773 ( .A(n156), .B(n64), .Z(n20951) );
  IV U20774 ( .A(n20951), .Z(n20458) );
  NOR U20775 ( .A(n20950), .B(n20458), .Z(n20459) );
  NOR U20776 ( .A(n20460), .B(n20459), .Z(n20955) );
  XOR U20777 ( .A(n20462), .B(n20461), .Z(n20954) );
  NOR U20778 ( .A(n20955), .B(n20954), .Z(n20463) );
  NOR U20779 ( .A(n20464), .B(n20463), .Z(n20490) );
  XOR U20780 ( .A(n20466), .B(n20465), .Z(n20489) );
  NOR U20781 ( .A(n20490), .B(n20489), .Z(n20467) );
  NOR U20782 ( .A(n20468), .B(n20467), .Z(n20473) );
  XOR U20783 ( .A(n20470), .B(n20469), .Z(n20472) );
  IV U20784 ( .A(n20472), .Z(n20471) );
  NOR U20785 ( .A(n20473), .B(n20471), .Z(n20476) );
  XOR U20786 ( .A(n20473), .B(n20472), .Z(n20971) );
  NOR U20787 ( .A(n163), .B(n64), .Z(n20972) );
  IV U20788 ( .A(n20972), .Z(n20474) );
  NOR U20789 ( .A(n20971), .B(n20474), .Z(n20475) );
  NOR U20790 ( .A(n20476), .B(n20475), .Z(n20976) );
  XOR U20791 ( .A(n20478), .B(n20477), .Z(n20975) );
  NOR U20792 ( .A(n20976), .B(n20975), .Z(n20479) );
  NOR U20793 ( .A(n20480), .B(n20479), .Z(n20983) );
  XOR U20794 ( .A(n20482), .B(n20481), .Z(n20984) );
  NOR U20795 ( .A(n20983), .B(n20984), .Z(n20483) );
  NOR U20796 ( .A(n20484), .B(n20483), .Z(n20987) );
  XOR U20797 ( .A(n20486), .B(n20485), .Z(n20986) );
  NOR U20798 ( .A(n20987), .B(n20986), .Z(n31548) );
  XOR U20799 ( .A(n20488), .B(n20487), .Z(n31555) );
  XOR U20800 ( .A(n31548), .B(n31555), .Z(n28549) );
  XOR U20801 ( .A(n20490), .B(n20489), .Z(n20962) );
  NOR U20802 ( .A(n150), .B(n65), .Z(n20919) );
  XOR U20803 ( .A(n20492), .B(n20491), .Z(n21415) );
  IV U20804 ( .A(n21415), .Z(n20912) );
  XOR U20805 ( .A(n20494), .B(n20493), .Z(n20495) );
  IV U20806 ( .A(n20495), .Z(n20899) );
  NOR U20807 ( .A(n145), .B(n65), .Z(n20900) );
  IV U20808 ( .A(n20900), .Z(n20496) );
  NOR U20809 ( .A(n20899), .B(n20496), .Z(n20903) );
  NOR U20810 ( .A(n143), .B(n65), .Z(n20896) );
  NOR U20811 ( .A(n137), .B(n65), .Z(n20497) );
  IV U20812 ( .A(n20497), .Z(n20873) );
  XOR U20813 ( .A(n20499), .B(n20498), .Z(n20872) );
  NOR U20814 ( .A(n20873), .B(n20872), .Z(n20876) );
  NOR U20815 ( .A(n135), .B(n65), .Z(n20869) );
  IV U20816 ( .A(n20869), .Z(n20863) );
  XOR U20817 ( .A(n20501), .B(n20500), .Z(n20502) );
  NOR U20818 ( .A(n133), .B(n65), .Z(n20503) );
  NOR U20819 ( .A(n20502), .B(n20503), .Z(n20861) );
  IV U20820 ( .A(n20502), .Z(n20996) );
  IV U20821 ( .A(n20503), .Z(n20995) );
  NOR U20822 ( .A(n20996), .B(n20995), .Z(n20859) );
  XOR U20823 ( .A(n20505), .B(n20504), .Z(n20506) );
  XOR U20824 ( .A(n20507), .B(n20506), .Z(n20854) );
  NOR U20825 ( .A(n131), .B(n65), .Z(n20855) );
  IV U20826 ( .A(n20855), .Z(n20508) );
  NOR U20827 ( .A(n20854), .B(n20508), .Z(n20857) );
  NOR U20828 ( .A(n128), .B(n65), .Z(n20851) );
  IV U20829 ( .A(n20851), .Z(n20512) );
  IV U20830 ( .A(n20509), .Z(n20511) );
  XOR U20831 ( .A(n20511), .B(n20510), .Z(n20850) );
  NOR U20832 ( .A(n20512), .B(n20850), .Z(n20853) );
  NOR U20833 ( .A(n126), .B(n65), .Z(n20513) );
  IV U20834 ( .A(n20513), .Z(n20845) );
  NOR U20835 ( .A(n125), .B(n65), .Z(n20516) );
  XOR U20836 ( .A(n20515), .B(n20514), .Z(n20517) );
  NOR U20837 ( .A(n20516), .B(n20517), .Z(n20842) );
  IV U20838 ( .A(n20516), .Z(n21010) );
  IV U20839 ( .A(n20517), .Z(n21009) );
  NOR U20840 ( .A(n21010), .B(n21009), .Z(n20840) );
  XOR U20841 ( .A(n20519), .B(n20518), .Z(n20520) );
  XOR U20842 ( .A(n20521), .B(n20520), .Z(n20836) );
  NOR U20843 ( .A(n123), .B(n65), .Z(n20835) );
  IV U20844 ( .A(n20835), .Z(n20522) );
  NOR U20845 ( .A(n20836), .B(n20522), .Z(n20838) );
  NOR U20846 ( .A(n120), .B(n65), .Z(n20830) );
  XOR U20847 ( .A(n20524), .B(n20523), .Z(n20829) );
  NOR U20848 ( .A(n20830), .B(n20829), .Z(n20833) );
  XOR U20849 ( .A(n20526), .B(n20525), .Z(n20825) );
  NOR U20850 ( .A(n119), .B(n65), .Z(n20824) );
  IV U20851 ( .A(n20824), .Z(n20527) );
  NOR U20852 ( .A(n20825), .B(n20527), .Z(n20827) );
  NOR U20853 ( .A(n79), .B(n65), .Z(n20819) );
  XOR U20854 ( .A(n20529), .B(n20528), .Z(n20818) );
  NOR U20855 ( .A(n20819), .B(n20818), .Z(n20822) );
  XOR U20856 ( .A(n20531), .B(n20530), .Z(n20814) );
  NOR U20857 ( .A(n117), .B(n65), .Z(n20813) );
  IV U20858 ( .A(n20813), .Z(n20532) );
  NOR U20859 ( .A(n20814), .B(n20532), .Z(n20816) );
  NOR U20860 ( .A(n80), .B(n65), .Z(n20808) );
  XOR U20861 ( .A(n20534), .B(n20533), .Z(n20807) );
  NOR U20862 ( .A(n20808), .B(n20807), .Z(n20811) );
  XOR U20863 ( .A(n20536), .B(n20535), .Z(n20803) );
  NOR U20864 ( .A(n116), .B(n65), .Z(n20802) );
  IV U20865 ( .A(n20802), .Z(n20537) );
  NOR U20866 ( .A(n20803), .B(n20537), .Z(n20805) );
  NOR U20867 ( .A(n81), .B(n65), .Z(n20797) );
  XOR U20868 ( .A(n20539), .B(n20538), .Z(n20796) );
  NOR U20869 ( .A(n20797), .B(n20796), .Z(n20800) );
  XOR U20870 ( .A(n20541), .B(n20540), .Z(n20792) );
  NOR U20871 ( .A(n115), .B(n65), .Z(n20791) );
  IV U20872 ( .A(n20791), .Z(n20542) );
  NOR U20873 ( .A(n20792), .B(n20542), .Z(n20794) );
  NOR U20874 ( .A(n82), .B(n65), .Z(n20786) );
  XOR U20875 ( .A(n20544), .B(n20543), .Z(n20785) );
  NOR U20876 ( .A(n20786), .B(n20785), .Z(n20789) );
  XOR U20877 ( .A(n20546), .B(n20545), .Z(n20781) );
  NOR U20878 ( .A(n114), .B(n65), .Z(n20780) );
  IV U20879 ( .A(n20780), .Z(n20547) );
  NOR U20880 ( .A(n20781), .B(n20547), .Z(n20783) );
  NOR U20881 ( .A(n83), .B(n65), .Z(n20775) );
  XOR U20882 ( .A(n20549), .B(n20548), .Z(n20774) );
  NOR U20883 ( .A(n20775), .B(n20774), .Z(n20778) );
  XOR U20884 ( .A(n20551), .B(n20550), .Z(n20770) );
  NOR U20885 ( .A(n113), .B(n65), .Z(n20769) );
  IV U20886 ( .A(n20769), .Z(n20552) );
  NOR U20887 ( .A(n20770), .B(n20552), .Z(n20772) );
  NOR U20888 ( .A(n84), .B(n65), .Z(n20764) );
  XOR U20889 ( .A(n20554), .B(n20553), .Z(n20763) );
  NOR U20890 ( .A(n20764), .B(n20763), .Z(n20767) );
  IV U20891 ( .A(n20555), .Z(n20557) );
  XOR U20892 ( .A(n20557), .B(n20556), .Z(n20758) );
  NOR U20893 ( .A(n112), .B(n65), .Z(n20759) );
  IV U20894 ( .A(n20759), .Z(n20558) );
  NOR U20895 ( .A(n20758), .B(n20558), .Z(n20761) );
  IV U20896 ( .A(n20559), .Z(n20561) );
  XOR U20897 ( .A(n20561), .B(n20560), .Z(n20754) );
  NOR U20898 ( .A(n85), .B(n65), .Z(n20755) );
  IV U20899 ( .A(n20755), .Z(n20562) );
  NOR U20900 ( .A(n20754), .B(n20562), .Z(n20757) );
  IV U20901 ( .A(n20563), .Z(n20565) );
  XOR U20902 ( .A(n20565), .B(n20564), .Z(n20750) );
  NOR U20903 ( .A(n111), .B(n65), .Z(n20751) );
  IV U20904 ( .A(n20751), .Z(n20566) );
  NOR U20905 ( .A(n20750), .B(n20566), .Z(n20753) );
  XOR U20906 ( .A(n20568), .B(n20567), .Z(n20746) );
  NOR U20907 ( .A(n86), .B(n65), .Z(n20747) );
  IV U20908 ( .A(n20747), .Z(n20569) );
  NOR U20909 ( .A(n20746), .B(n20569), .Z(n20749) );
  XOR U20910 ( .A(n20571), .B(n20570), .Z(n20743) );
  NOR U20911 ( .A(n110), .B(n65), .Z(n20742) );
  IV U20912 ( .A(n20742), .Z(n20572) );
  NOR U20913 ( .A(n20743), .B(n20572), .Z(n20745) );
  XOR U20914 ( .A(n20574), .B(n20573), .Z(n20738) );
  NOR U20915 ( .A(n109), .B(n65), .Z(n20739) );
  IV U20916 ( .A(n20739), .Z(n20575) );
  NOR U20917 ( .A(n20738), .B(n20575), .Z(n20741) );
  IV U20918 ( .A(n20576), .Z(n20578) );
  XOR U20919 ( .A(n20578), .B(n20577), .Z(n20734) );
  NOR U20920 ( .A(n108), .B(n65), .Z(n20735) );
  IV U20921 ( .A(n20735), .Z(n20579) );
  NOR U20922 ( .A(n20734), .B(n20579), .Z(n20737) );
  XOR U20923 ( .A(n20581), .B(n20580), .Z(n20730) );
  IV U20924 ( .A(n20730), .Z(n20583) );
  NOR U20925 ( .A(n87), .B(n65), .Z(n20582) );
  IV U20926 ( .A(n20582), .Z(n20731) );
  NOR U20927 ( .A(n20583), .B(n20731), .Z(n20733) );
  IV U20928 ( .A(n20584), .Z(n20586) );
  XOR U20929 ( .A(n20586), .B(n20585), .Z(n20726) );
  NOR U20930 ( .A(n107), .B(n65), .Z(n20727) );
  IV U20931 ( .A(n20727), .Z(n20587) );
  NOR U20932 ( .A(n20726), .B(n20587), .Z(n20729) );
  IV U20933 ( .A(n20588), .Z(n20590) );
  XOR U20934 ( .A(n20590), .B(n20589), .Z(n20722) );
  NOR U20935 ( .A(n88), .B(n65), .Z(n20723) );
  IV U20936 ( .A(n20723), .Z(n20591) );
  NOR U20937 ( .A(n20722), .B(n20591), .Z(n20725) );
  IV U20938 ( .A(n20592), .Z(n20594) );
  XOR U20939 ( .A(n20594), .B(n20593), .Z(n20718) );
  NOR U20940 ( .A(n106), .B(n65), .Z(n20719) );
  IV U20941 ( .A(n20719), .Z(n20595) );
  NOR U20942 ( .A(n20718), .B(n20595), .Z(n20721) );
  XOR U20943 ( .A(n20597), .B(n20596), .Z(n20714) );
  NOR U20944 ( .A(n105), .B(n65), .Z(n20715) );
  IV U20945 ( .A(n20715), .Z(n20598) );
  NOR U20946 ( .A(n20714), .B(n20598), .Z(n20717) );
  XOR U20947 ( .A(n20600), .B(n20599), .Z(n20702) );
  IV U20948 ( .A(n20702), .Z(n20602) );
  NOR U20949 ( .A(n89), .B(n65), .Z(n20601) );
  IV U20950 ( .A(n20601), .Z(n20703) );
  NOR U20951 ( .A(n20602), .B(n20703), .Z(n20705) );
  IV U20952 ( .A(n20603), .Z(n20605) );
  XOR U20953 ( .A(n20605), .B(n20604), .Z(n20698) );
  NOR U20954 ( .A(n103), .B(n65), .Z(n20699) );
  IV U20955 ( .A(n20699), .Z(n20606) );
  NOR U20956 ( .A(n20698), .B(n20606), .Z(n20701) );
  IV U20957 ( .A(n20607), .Z(n20609) );
  XOR U20958 ( .A(n20609), .B(n20608), .Z(n20694) );
  NOR U20959 ( .A(n90), .B(n65), .Z(n20695) );
  IV U20960 ( .A(n20695), .Z(n20610) );
  NOR U20961 ( .A(n20694), .B(n20610), .Z(n20697) );
  IV U20962 ( .A(n20611), .Z(n20613) );
  XOR U20963 ( .A(n20613), .B(n20612), .Z(n20690) );
  NOR U20964 ( .A(n102), .B(n65), .Z(n20691) );
  IV U20965 ( .A(n20691), .Z(n20614) );
  NOR U20966 ( .A(n20690), .B(n20614), .Z(n20693) );
  IV U20967 ( .A(n20615), .Z(n20617) );
  XOR U20968 ( .A(n20617), .B(n20616), .Z(n20686) );
  NOR U20969 ( .A(n101), .B(n65), .Z(n20687) );
  IV U20970 ( .A(n20687), .Z(n20618) );
  NOR U20971 ( .A(n20686), .B(n20618), .Z(n20689) );
  IV U20972 ( .A(n20619), .Z(n20621) );
  XOR U20973 ( .A(n20621), .B(n20620), .Z(n20682) );
  NOR U20974 ( .A(n100), .B(n65), .Z(n20683) );
  IV U20975 ( .A(n20683), .Z(n20622) );
  NOR U20976 ( .A(n20682), .B(n20622), .Z(n20685) );
  IV U20977 ( .A(n20623), .Z(n20625) );
  XOR U20978 ( .A(n20625), .B(n20624), .Z(n20678) );
  NOR U20979 ( .A(n99), .B(n65), .Z(n20679) );
  IV U20980 ( .A(n20679), .Z(n20626) );
  NOR U20981 ( .A(n20678), .B(n20626), .Z(n20681) );
  IV U20982 ( .A(n20627), .Z(n20629) );
  XOR U20983 ( .A(n20629), .B(n20628), .Z(n20674) );
  NOR U20984 ( .A(n98), .B(n65), .Z(n20675) );
  IV U20985 ( .A(n20675), .Z(n20630) );
  NOR U20986 ( .A(n20674), .B(n20630), .Z(n20677) );
  IV U20987 ( .A(n20631), .Z(n20633) );
  XOR U20988 ( .A(n20633), .B(n20632), .Z(n20670) );
  NOR U20989 ( .A(n91), .B(n65), .Z(n20671) );
  IV U20990 ( .A(n20671), .Z(n20634) );
  NOR U20991 ( .A(n20670), .B(n20634), .Z(n20673) );
  XOR U20992 ( .A(n20636), .B(n20635), .Z(n20658) );
  IV U20993 ( .A(n20658), .Z(n20638) );
  NOR U20994 ( .A(n96), .B(n65), .Z(n20637) );
  IV U20995 ( .A(n20637), .Z(n20659) );
  NOR U20996 ( .A(n20638), .B(n20659), .Z(n20661) );
  NOR U20997 ( .A(n95), .B(n65), .Z(n20655) );
  IV U20998 ( .A(n20655), .Z(n20641) );
  XOR U20999 ( .A(n20640), .B(n20639), .Z(n20654) );
  NOR U21000 ( .A(n20641), .B(n20654), .Z(n20657) );
  NOR U21001 ( .A(n65), .B(n93), .Z(n21650) );
  IV U21002 ( .A(n21650), .Z(n20642) );
  NOR U21003 ( .A(n64), .B(n168), .Z(n20650) );
  IV U21004 ( .A(n20650), .Z(n20645) );
  NOR U21005 ( .A(n20642), .B(n20645), .Z(n20643) );
  IV U21006 ( .A(n20643), .Z(n20644) );
  NOR U21007 ( .A(n94), .B(n20644), .Z(n20653) );
  NOR U21008 ( .A(n20645), .B(n93), .Z(n20646) );
  XOR U21009 ( .A(n94), .B(n20646), .Z(n20647) );
  NOR U21010 ( .A(n65), .B(n20647), .Z(n20648) );
  IV U21011 ( .A(n20648), .Z(n21139) );
  XOR U21012 ( .A(n20650), .B(n20649), .Z(n21138) );
  IV U21013 ( .A(n21138), .Z(n20651) );
  NOR U21014 ( .A(n21139), .B(n20651), .Z(n20652) );
  NOR U21015 ( .A(n20653), .B(n20652), .Z(n21135) );
  XOR U21016 ( .A(n20655), .B(n20654), .Z(n21134) );
  NOR U21017 ( .A(n21135), .B(n21134), .Z(n20656) );
  NOR U21018 ( .A(n20657), .B(n20656), .Z(n21162) );
  XOR U21019 ( .A(n20659), .B(n20658), .Z(n21161) );
  NOR U21020 ( .A(n21162), .B(n21161), .Z(n20660) );
  NOR U21021 ( .A(n20661), .B(n20660), .Z(n20666) );
  XOR U21022 ( .A(n20663), .B(n20662), .Z(n20665) );
  IV U21023 ( .A(n20665), .Z(n20664) );
  NOR U21024 ( .A(n20666), .B(n20664), .Z(n20669) );
  XOR U21025 ( .A(n20666), .B(n20665), .Z(n21131) );
  NOR U21026 ( .A(n97), .B(n65), .Z(n21132) );
  IV U21027 ( .A(n21132), .Z(n20667) );
  NOR U21028 ( .A(n21131), .B(n20667), .Z(n20668) );
  NOR U21029 ( .A(n20669), .B(n20668), .Z(n21127) );
  XOR U21030 ( .A(n20671), .B(n20670), .Z(n21128) );
  NOR U21031 ( .A(n21127), .B(n21128), .Z(n20672) );
  NOR U21032 ( .A(n20673), .B(n20672), .Z(n21123) );
  XOR U21033 ( .A(n20675), .B(n20674), .Z(n21124) );
  NOR U21034 ( .A(n21123), .B(n21124), .Z(n20676) );
  NOR U21035 ( .A(n20677), .B(n20676), .Z(n21119) );
  XOR U21036 ( .A(n20679), .B(n20678), .Z(n21120) );
  NOR U21037 ( .A(n21119), .B(n21120), .Z(n20680) );
  NOR U21038 ( .A(n20681), .B(n20680), .Z(n21115) );
  XOR U21039 ( .A(n20683), .B(n20682), .Z(n21116) );
  NOR U21040 ( .A(n21115), .B(n21116), .Z(n20684) );
  NOR U21041 ( .A(n20685), .B(n20684), .Z(n21111) );
  XOR U21042 ( .A(n20687), .B(n20686), .Z(n21112) );
  NOR U21043 ( .A(n21111), .B(n21112), .Z(n20688) );
  NOR U21044 ( .A(n20689), .B(n20688), .Z(n21107) );
  XOR U21045 ( .A(n20691), .B(n20690), .Z(n21108) );
  NOR U21046 ( .A(n21107), .B(n21108), .Z(n20692) );
  NOR U21047 ( .A(n20693), .B(n20692), .Z(n21103) );
  XOR U21048 ( .A(n20695), .B(n20694), .Z(n21104) );
  NOR U21049 ( .A(n21103), .B(n21104), .Z(n20696) );
  NOR U21050 ( .A(n20697), .B(n20696), .Z(n21100) );
  XOR U21051 ( .A(n20699), .B(n20698), .Z(n21099) );
  NOR U21052 ( .A(n21100), .B(n21099), .Z(n20700) );
  NOR U21053 ( .A(n20701), .B(n20700), .Z(n21206) );
  XOR U21054 ( .A(n20703), .B(n20702), .Z(n21205) );
  NOR U21055 ( .A(n21206), .B(n21205), .Z(n20704) );
  NOR U21056 ( .A(n20705), .B(n20704), .Z(n20710) );
  XOR U21057 ( .A(n20707), .B(n20706), .Z(n20709) );
  IV U21058 ( .A(n20709), .Z(n20708) );
  NOR U21059 ( .A(n20710), .B(n20708), .Z(n20713) );
  XOR U21060 ( .A(n20710), .B(n20709), .Z(n21096) );
  NOR U21061 ( .A(n104), .B(n65), .Z(n21097) );
  IV U21062 ( .A(n21097), .Z(n20711) );
  NOR U21063 ( .A(n21096), .B(n20711), .Z(n20712) );
  NOR U21064 ( .A(n20713), .B(n20712), .Z(n21092) );
  XOR U21065 ( .A(n20715), .B(n20714), .Z(n21093) );
  NOR U21066 ( .A(n21092), .B(n21093), .Z(n20716) );
  NOR U21067 ( .A(n20717), .B(n20716), .Z(n21088) );
  XOR U21068 ( .A(n20719), .B(n20718), .Z(n21089) );
  NOR U21069 ( .A(n21088), .B(n21089), .Z(n20720) );
  NOR U21070 ( .A(n20721), .B(n20720), .Z(n21084) );
  XOR U21071 ( .A(n20723), .B(n20722), .Z(n21085) );
  NOR U21072 ( .A(n21084), .B(n21085), .Z(n20724) );
  NOR U21073 ( .A(n20725), .B(n20724), .Z(n21081) );
  XOR U21074 ( .A(n20727), .B(n20726), .Z(n21080) );
  NOR U21075 ( .A(n21081), .B(n21080), .Z(n20728) );
  NOR U21076 ( .A(n20729), .B(n20728), .Z(n21234) );
  XOR U21077 ( .A(n20731), .B(n20730), .Z(n21233) );
  NOR U21078 ( .A(n21234), .B(n21233), .Z(n20732) );
  NOR U21079 ( .A(n20733), .B(n20732), .Z(n21076) );
  XOR U21080 ( .A(n20735), .B(n20734), .Z(n21077) );
  NOR U21081 ( .A(n21076), .B(n21077), .Z(n20736) );
  NOR U21082 ( .A(n20737), .B(n20736), .Z(n21072) );
  XOR U21083 ( .A(n20739), .B(n20738), .Z(n21073) );
  NOR U21084 ( .A(n21072), .B(n21073), .Z(n20740) );
  NOR U21085 ( .A(n20741), .B(n20740), .Z(n21068) );
  XOR U21086 ( .A(n20743), .B(n20742), .Z(n21069) );
  NOR U21087 ( .A(n21068), .B(n21069), .Z(n20744) );
  NOR U21088 ( .A(n20745), .B(n20744), .Z(n21064) );
  XOR U21089 ( .A(n20747), .B(n20746), .Z(n21065) );
  NOR U21090 ( .A(n21064), .B(n21065), .Z(n20748) );
  NOR U21091 ( .A(n20749), .B(n20748), .Z(n21060) );
  XOR U21092 ( .A(n20751), .B(n20750), .Z(n21061) );
  NOR U21093 ( .A(n21060), .B(n21061), .Z(n20752) );
  NOR U21094 ( .A(n20753), .B(n20752), .Z(n21056) );
  XOR U21095 ( .A(n20755), .B(n20754), .Z(n21057) );
  NOR U21096 ( .A(n21056), .B(n21057), .Z(n20756) );
  NOR U21097 ( .A(n20757), .B(n20756), .Z(n21052) );
  XOR U21098 ( .A(n20759), .B(n20758), .Z(n21053) );
  NOR U21099 ( .A(n21052), .B(n21053), .Z(n20760) );
  NOR U21100 ( .A(n20761), .B(n20760), .Z(n20762) );
  IV U21101 ( .A(n20762), .Z(n21050) );
  XOR U21102 ( .A(n20764), .B(n20763), .Z(n20765) );
  IV U21103 ( .A(n20765), .Z(n21049) );
  NOR U21104 ( .A(n21050), .B(n21049), .Z(n20766) );
  NOR U21105 ( .A(n20767), .B(n20766), .Z(n20768) );
  IV U21106 ( .A(n20768), .Z(n21048) );
  XOR U21107 ( .A(n20770), .B(n20769), .Z(n21047) );
  NOR U21108 ( .A(n21048), .B(n21047), .Z(n20771) );
  NOR U21109 ( .A(n20772), .B(n20771), .Z(n20773) );
  IV U21110 ( .A(n20773), .Z(n21045) );
  XOR U21111 ( .A(n20775), .B(n20774), .Z(n20776) );
  IV U21112 ( .A(n20776), .Z(n21044) );
  NOR U21113 ( .A(n21045), .B(n21044), .Z(n20777) );
  NOR U21114 ( .A(n20778), .B(n20777), .Z(n20779) );
  IV U21115 ( .A(n20779), .Z(n21040) );
  XOR U21116 ( .A(n20781), .B(n20780), .Z(n21039) );
  NOR U21117 ( .A(n21040), .B(n21039), .Z(n20782) );
  NOR U21118 ( .A(n20783), .B(n20782), .Z(n20784) );
  IV U21119 ( .A(n20784), .Z(n21037) );
  XOR U21120 ( .A(n20786), .B(n20785), .Z(n20787) );
  IV U21121 ( .A(n20787), .Z(n21036) );
  NOR U21122 ( .A(n21037), .B(n21036), .Z(n20788) );
  NOR U21123 ( .A(n20789), .B(n20788), .Z(n20790) );
  IV U21124 ( .A(n20790), .Z(n21035) );
  XOR U21125 ( .A(n20792), .B(n20791), .Z(n21034) );
  NOR U21126 ( .A(n21035), .B(n21034), .Z(n20793) );
  NOR U21127 ( .A(n20794), .B(n20793), .Z(n20795) );
  IV U21128 ( .A(n20795), .Z(n21032) );
  XOR U21129 ( .A(n20797), .B(n20796), .Z(n20798) );
  IV U21130 ( .A(n20798), .Z(n21031) );
  NOR U21131 ( .A(n21032), .B(n21031), .Z(n20799) );
  NOR U21132 ( .A(n20800), .B(n20799), .Z(n20801) );
  IV U21133 ( .A(n20801), .Z(n21030) );
  XOR U21134 ( .A(n20803), .B(n20802), .Z(n21029) );
  NOR U21135 ( .A(n21030), .B(n21029), .Z(n20804) );
  NOR U21136 ( .A(n20805), .B(n20804), .Z(n20806) );
  IV U21137 ( .A(n20806), .Z(n21027) );
  XOR U21138 ( .A(n20808), .B(n20807), .Z(n20809) );
  IV U21139 ( .A(n20809), .Z(n21026) );
  NOR U21140 ( .A(n21027), .B(n21026), .Z(n20810) );
  NOR U21141 ( .A(n20811), .B(n20810), .Z(n20812) );
  IV U21142 ( .A(n20812), .Z(n21025) );
  XOR U21143 ( .A(n20814), .B(n20813), .Z(n21024) );
  NOR U21144 ( .A(n21025), .B(n21024), .Z(n20815) );
  NOR U21145 ( .A(n20816), .B(n20815), .Z(n20817) );
  IV U21146 ( .A(n20817), .Z(n21022) );
  XOR U21147 ( .A(n20819), .B(n20818), .Z(n20820) );
  IV U21148 ( .A(n20820), .Z(n21021) );
  NOR U21149 ( .A(n21022), .B(n21021), .Z(n20821) );
  NOR U21150 ( .A(n20822), .B(n20821), .Z(n20823) );
  IV U21151 ( .A(n20823), .Z(n21020) );
  XOR U21152 ( .A(n20825), .B(n20824), .Z(n21019) );
  NOR U21153 ( .A(n21020), .B(n21019), .Z(n20826) );
  NOR U21154 ( .A(n20827), .B(n20826), .Z(n20828) );
  IV U21155 ( .A(n20828), .Z(n21017) );
  XOR U21156 ( .A(n20830), .B(n20829), .Z(n20831) );
  IV U21157 ( .A(n20831), .Z(n21016) );
  NOR U21158 ( .A(n21017), .B(n21016), .Z(n20832) );
  NOR U21159 ( .A(n20833), .B(n20832), .Z(n20834) );
  IV U21160 ( .A(n20834), .Z(n21015) );
  XOR U21161 ( .A(n20836), .B(n20835), .Z(n21014) );
  NOR U21162 ( .A(n21015), .B(n21014), .Z(n20837) );
  NOR U21163 ( .A(n20838), .B(n20837), .Z(n21012) );
  IV U21164 ( .A(n21012), .Z(n20839) );
  NOR U21165 ( .A(n20840), .B(n20839), .Z(n20841) );
  NOR U21166 ( .A(n20842), .B(n20841), .Z(n20844) );
  IV U21167 ( .A(n20844), .Z(n20843) );
  NOR U21168 ( .A(n20845), .B(n20843), .Z(n20849) );
  XOR U21169 ( .A(n20845), .B(n20844), .Z(n21006) );
  XOR U21170 ( .A(n20847), .B(n20846), .Z(n21005) );
  NOR U21171 ( .A(n21006), .B(n21005), .Z(n20848) );
  NOR U21172 ( .A(n20849), .B(n20848), .Z(n21354) );
  XOR U21173 ( .A(n20851), .B(n20850), .Z(n21355) );
  NOR U21174 ( .A(n21354), .B(n21355), .Z(n20852) );
  NOR U21175 ( .A(n20853), .B(n20852), .Z(n21000) );
  XOR U21176 ( .A(n20855), .B(n20854), .Z(n21001) );
  NOR U21177 ( .A(n21000), .B(n21001), .Z(n20856) );
  NOR U21178 ( .A(n20857), .B(n20856), .Z(n20998) );
  IV U21179 ( .A(n20998), .Z(n20858) );
  NOR U21180 ( .A(n20859), .B(n20858), .Z(n20860) );
  NOR U21181 ( .A(n20861), .B(n20860), .Z(n20862) );
  IV U21182 ( .A(n20862), .Z(n20868) );
  NOR U21183 ( .A(n20863), .B(n20868), .Z(n20871) );
  XOR U21184 ( .A(n20865), .B(n20864), .Z(n20866) );
  XOR U21185 ( .A(n20867), .B(n20866), .Z(n20992) );
  XOR U21186 ( .A(n20869), .B(n20868), .Z(n20991) );
  NOR U21187 ( .A(n20992), .B(n20991), .Z(n20870) );
  NOR U21188 ( .A(n20871), .B(n20870), .Z(n21373) );
  XOR U21189 ( .A(n20873), .B(n20872), .Z(n21374) );
  IV U21190 ( .A(n21374), .Z(n20874) );
  NOR U21191 ( .A(n21373), .B(n20874), .Z(n20875) );
  NOR U21192 ( .A(n20876), .B(n20875), .Z(n20879) );
  NOR U21193 ( .A(n139), .B(n65), .Z(n20878) );
  IV U21194 ( .A(n20878), .Z(n20877) );
  NOR U21195 ( .A(n20879), .B(n20877), .Z(n20884) );
  XOR U21196 ( .A(n20879), .B(n20878), .Z(n20988) );
  XOR U21197 ( .A(n20881), .B(n20880), .Z(n20989) );
  IV U21198 ( .A(n20989), .Z(n20882) );
  NOR U21199 ( .A(n20988), .B(n20882), .Z(n20883) );
  NOR U21200 ( .A(n20884), .B(n20883), .Z(n20889) );
  NOR U21201 ( .A(n141), .B(n65), .Z(n20888) );
  IV U21202 ( .A(n20888), .Z(n20885) );
  NOR U21203 ( .A(n20889), .B(n20885), .Z(n20891) );
  XOR U21204 ( .A(n20887), .B(n20886), .Z(n21382) );
  XOR U21205 ( .A(n20889), .B(n20888), .Z(n21381) );
  NOR U21206 ( .A(n21382), .B(n21381), .Z(n20890) );
  NOR U21207 ( .A(n20891), .B(n20890), .Z(n20895) );
  IV U21208 ( .A(n20895), .Z(n20892) );
  NOR U21209 ( .A(n20896), .B(n20892), .Z(n20898) );
  XOR U21210 ( .A(n20894), .B(n20893), .Z(n21391) );
  XOR U21211 ( .A(n20896), .B(n20895), .Z(n21390) );
  NOR U21212 ( .A(n21391), .B(n21390), .Z(n20897) );
  NOR U21213 ( .A(n20898), .B(n20897), .Z(n21400) );
  IV U21214 ( .A(n21400), .Z(n20901) );
  XOR U21215 ( .A(n20900), .B(n20899), .Z(n21399) );
  NOR U21216 ( .A(n20901), .B(n21399), .Z(n20902) );
  NOR U21217 ( .A(n20903), .B(n20902), .Z(n20906) );
  NOR U21218 ( .A(n147), .B(n65), .Z(n20905) );
  IV U21219 ( .A(n20905), .Z(n20904) );
  NOR U21220 ( .A(n20906), .B(n20904), .Z(n20910) );
  XOR U21221 ( .A(n20906), .B(n20905), .Z(n21406) );
  XOR U21222 ( .A(n20908), .B(n20907), .Z(n21407) );
  NOR U21223 ( .A(n21406), .B(n21407), .Z(n20909) );
  NOR U21224 ( .A(n20910), .B(n20909), .Z(n21413) );
  IV U21225 ( .A(n21413), .Z(n20911) );
  NOR U21226 ( .A(n20912), .B(n20911), .Z(n20915) );
  NOR U21227 ( .A(n21415), .B(n21413), .Z(n20913) );
  NOR U21228 ( .A(n148), .B(n65), .Z(n21412) );
  NOR U21229 ( .A(n20913), .B(n21412), .Z(n20914) );
  NOR U21230 ( .A(n20915), .B(n20914), .Z(n20918) );
  NOR U21231 ( .A(n20919), .B(n20918), .Z(n20922) );
  XOR U21232 ( .A(n20917), .B(n20916), .Z(n21422) );
  XOR U21233 ( .A(n20919), .B(n20918), .Z(n20920) );
  IV U21234 ( .A(n20920), .Z(n21423) );
  NOR U21235 ( .A(n21422), .B(n21423), .Z(n20921) );
  NOR U21236 ( .A(n20922), .B(n20921), .Z(n20926) );
  IV U21237 ( .A(n20926), .Z(n20924) );
  NOR U21238 ( .A(n153), .B(n65), .Z(n20923) );
  IV U21239 ( .A(n20923), .Z(n20925) );
  NOR U21240 ( .A(n20924), .B(n20925), .Z(n20930) );
  XOR U21241 ( .A(n20926), .B(n20925), .Z(n21429) );
  XOR U21242 ( .A(n20928), .B(n20927), .Z(n21428) );
  NOR U21243 ( .A(n21429), .B(n21428), .Z(n20929) );
  NOR U21244 ( .A(n20930), .B(n20929), .Z(n20935) );
  XOR U21245 ( .A(n20932), .B(n20931), .Z(n20934) );
  IV U21246 ( .A(n20934), .Z(n20933) );
  NOR U21247 ( .A(n20935), .B(n20933), .Z(n20938) );
  XOR U21248 ( .A(n20935), .B(n20934), .Z(n21439) );
  NOR U21249 ( .A(n155), .B(n65), .Z(n20936) );
  IV U21250 ( .A(n20936), .Z(n21438) );
  NOR U21251 ( .A(n21439), .B(n21438), .Z(n20937) );
  NOR U21252 ( .A(n20938), .B(n20937), .Z(n20941) );
  NOR U21253 ( .A(n156), .B(n65), .Z(n20940) );
  IV U21254 ( .A(n20940), .Z(n20939) );
  NOR U21255 ( .A(n20941), .B(n20939), .Z(n20946) );
  XOR U21256 ( .A(n20941), .B(n20940), .Z(n21447) );
  XOR U21257 ( .A(n20943), .B(n20942), .Z(n21448) );
  IV U21258 ( .A(n21448), .Z(n20944) );
  NOR U21259 ( .A(n21447), .B(n20944), .Z(n20945) );
  NOR U21260 ( .A(n20946), .B(n20945), .Z(n20949) );
  NOR U21261 ( .A(n158), .B(n65), .Z(n20948) );
  IV U21262 ( .A(n20948), .Z(n20947) );
  NOR U21263 ( .A(n20949), .B(n20947), .Z(n20953) );
  XOR U21264 ( .A(n20949), .B(n20948), .Z(n21451) );
  XOR U21265 ( .A(n20951), .B(n20950), .Z(n21452) );
  NOR U21266 ( .A(n21451), .B(n21452), .Z(n20952) );
  NOR U21267 ( .A(n20953), .B(n20952), .Z(n20958) );
  XOR U21268 ( .A(n20955), .B(n20954), .Z(n20957) );
  IV U21269 ( .A(n20957), .Z(n20956) );
  NOR U21270 ( .A(n20958), .B(n20956), .Z(n20961) );
  XOR U21271 ( .A(n20958), .B(n20957), .Z(n21462) );
  NOR U21272 ( .A(n161), .B(n65), .Z(n20959) );
  IV U21273 ( .A(n20959), .Z(n21461) );
  NOR U21274 ( .A(n21462), .B(n21461), .Z(n20960) );
  NOR U21275 ( .A(n20961), .B(n20960), .Z(n20963) );
  IV U21276 ( .A(n20963), .Z(n21468) );
  NOR U21277 ( .A(n20962), .B(n21468), .Z(n20966) );
  IV U21278 ( .A(n20962), .Z(n21469) );
  NOR U21279 ( .A(n20963), .B(n21469), .Z(n20964) );
  NOR U21280 ( .A(n163), .B(n65), .Z(n21471) );
  NOR U21281 ( .A(n20964), .B(n21471), .Z(n20965) );
  NOR U21282 ( .A(n20966), .B(n20965), .Z(n20970) );
  IV U21283 ( .A(n20970), .Z(n20968) );
  NOR U21284 ( .A(n165), .B(n65), .Z(n20967) );
  IV U21285 ( .A(n20967), .Z(n20969) );
  NOR U21286 ( .A(n20968), .B(n20969), .Z(n20974) );
  XOR U21287 ( .A(n20970), .B(n20969), .Z(n21477) );
  XOR U21288 ( .A(n20972), .B(n20971), .Z(n21476) );
  NOR U21289 ( .A(n21477), .B(n21476), .Z(n20973) );
  NOR U21290 ( .A(n20974), .B(n20973), .Z(n20979) );
  XOR U21291 ( .A(n20976), .B(n20975), .Z(n20978) );
  IV U21292 ( .A(n20978), .Z(n20977) );
  NOR U21293 ( .A(n20979), .B(n20977), .Z(n20982) );
  XOR U21294 ( .A(n20979), .B(n20978), .Z(n21484) );
  NOR U21295 ( .A(n167), .B(n65), .Z(n21485) );
  IV U21296 ( .A(n21485), .Z(n20980) );
  NOR U21297 ( .A(n21484), .B(n20980), .Z(n20981) );
  NOR U21298 ( .A(n20982), .B(n20981), .Z(n21487) );
  IV U21299 ( .A(n20983), .Z(n20985) );
  XOR U21300 ( .A(n20985), .B(n20984), .Z(n21486) );
  NOR U21301 ( .A(n21487), .B(n21486), .Z(n28544) );
  XOR U21302 ( .A(n20987), .B(n20986), .Z(n28545) );
  NOR U21303 ( .A(n28544), .B(n28545), .Z(n28547) );
  NOR U21304 ( .A(n163), .B(n66), .Z(n21459) );
  NOR U21305 ( .A(n156), .B(n66), .Z(n21436) );
  NOR U21306 ( .A(n141), .B(n66), .Z(n21378) );
  IV U21307 ( .A(n21378), .Z(n20990) );
  XOR U21308 ( .A(n20989), .B(n20988), .Z(n21377) );
  NOR U21309 ( .A(n20990), .B(n21377), .Z(n21380) );
  XOR U21310 ( .A(n20992), .B(n20991), .Z(n20994) );
  IV U21311 ( .A(n20994), .Z(n21493) );
  NOR U21312 ( .A(n137), .B(n66), .Z(n20993) );
  IV U21313 ( .A(n20993), .Z(n21492) );
  NOR U21314 ( .A(n21493), .B(n21492), .Z(n21369) );
  NOR U21315 ( .A(n20994), .B(n20993), .Z(n21367) );
  XOR U21316 ( .A(n20996), .B(n20995), .Z(n20997) );
  XOR U21317 ( .A(n20998), .B(n20997), .Z(n21364) );
  NOR U21318 ( .A(n135), .B(n66), .Z(n21363) );
  IV U21319 ( .A(n21363), .Z(n20999) );
  NOR U21320 ( .A(n21364), .B(n20999), .Z(n21366) );
  NOR U21321 ( .A(n133), .B(n66), .Z(n21360) );
  IV U21322 ( .A(n21360), .Z(n21003) );
  XOR U21323 ( .A(n21001), .B(n21000), .Z(n21002) );
  IV U21324 ( .A(n21002), .Z(n21359) );
  NOR U21325 ( .A(n21003), .B(n21359), .Z(n21362) );
  NOR U21326 ( .A(n131), .B(n66), .Z(n21004) );
  IV U21327 ( .A(n21004), .Z(n21353) );
  NOR U21328 ( .A(n128), .B(n66), .Z(n21007) );
  XOR U21329 ( .A(n21006), .B(n21005), .Z(n21008) );
  NOR U21330 ( .A(n21007), .B(n21008), .Z(n21350) );
  IV U21331 ( .A(n21007), .Z(n21510) );
  IV U21332 ( .A(n21008), .Z(n21509) );
  NOR U21333 ( .A(n21510), .B(n21509), .Z(n21348) );
  XOR U21334 ( .A(n21010), .B(n21009), .Z(n21011) );
  XOR U21335 ( .A(n21012), .B(n21011), .Z(n21344) );
  NOR U21336 ( .A(n126), .B(n66), .Z(n21343) );
  IV U21337 ( .A(n21343), .Z(n21013) );
  NOR U21338 ( .A(n21344), .B(n21013), .Z(n21346) );
  NOR U21339 ( .A(n125), .B(n66), .Z(n21338) );
  XOR U21340 ( .A(n21015), .B(n21014), .Z(n21337) );
  NOR U21341 ( .A(n21338), .B(n21337), .Z(n21341) );
  XOR U21342 ( .A(n21017), .B(n21016), .Z(n21333) );
  NOR U21343 ( .A(n123), .B(n66), .Z(n21332) );
  IV U21344 ( .A(n21332), .Z(n21018) );
  NOR U21345 ( .A(n21333), .B(n21018), .Z(n21335) );
  NOR U21346 ( .A(n120), .B(n66), .Z(n21327) );
  XOR U21347 ( .A(n21020), .B(n21019), .Z(n21326) );
  NOR U21348 ( .A(n21327), .B(n21326), .Z(n21330) );
  XOR U21349 ( .A(n21022), .B(n21021), .Z(n21322) );
  NOR U21350 ( .A(n119), .B(n66), .Z(n21321) );
  IV U21351 ( .A(n21321), .Z(n21023) );
  NOR U21352 ( .A(n21322), .B(n21023), .Z(n21324) );
  NOR U21353 ( .A(n79), .B(n66), .Z(n21316) );
  XOR U21354 ( .A(n21025), .B(n21024), .Z(n21315) );
  NOR U21355 ( .A(n21316), .B(n21315), .Z(n21319) );
  XOR U21356 ( .A(n21027), .B(n21026), .Z(n21311) );
  NOR U21357 ( .A(n117), .B(n66), .Z(n21310) );
  IV U21358 ( .A(n21310), .Z(n21028) );
  NOR U21359 ( .A(n21311), .B(n21028), .Z(n21313) );
  NOR U21360 ( .A(n80), .B(n66), .Z(n21305) );
  XOR U21361 ( .A(n21030), .B(n21029), .Z(n21304) );
  NOR U21362 ( .A(n21305), .B(n21304), .Z(n21308) );
  XOR U21363 ( .A(n21032), .B(n21031), .Z(n21300) );
  NOR U21364 ( .A(n116), .B(n66), .Z(n21299) );
  IV U21365 ( .A(n21299), .Z(n21033) );
  NOR U21366 ( .A(n21300), .B(n21033), .Z(n21302) );
  NOR U21367 ( .A(n81), .B(n66), .Z(n21294) );
  XOR U21368 ( .A(n21035), .B(n21034), .Z(n21293) );
  NOR U21369 ( .A(n21294), .B(n21293), .Z(n21297) );
  XOR U21370 ( .A(n21037), .B(n21036), .Z(n21289) );
  NOR U21371 ( .A(n115), .B(n66), .Z(n21288) );
  IV U21372 ( .A(n21288), .Z(n21038) );
  NOR U21373 ( .A(n21289), .B(n21038), .Z(n21291) );
  NOR U21374 ( .A(n82), .B(n66), .Z(n21042) );
  XOR U21375 ( .A(n21040), .B(n21039), .Z(n21041) );
  NOR U21376 ( .A(n21042), .B(n21041), .Z(n21286) );
  XOR U21377 ( .A(n21042), .B(n21041), .Z(n21043) );
  IV U21378 ( .A(n21043), .Z(n21542) );
  XOR U21379 ( .A(n21045), .B(n21044), .Z(n21281) );
  NOR U21380 ( .A(n114), .B(n66), .Z(n21280) );
  IV U21381 ( .A(n21280), .Z(n21046) );
  NOR U21382 ( .A(n21281), .B(n21046), .Z(n21283) );
  NOR U21383 ( .A(n83), .B(n66), .Z(n21275) );
  XOR U21384 ( .A(n21048), .B(n21047), .Z(n21274) );
  NOR U21385 ( .A(n21275), .B(n21274), .Z(n21278) );
  XOR U21386 ( .A(n21050), .B(n21049), .Z(n21270) );
  NOR U21387 ( .A(n113), .B(n66), .Z(n21269) );
  IV U21388 ( .A(n21269), .Z(n21051) );
  NOR U21389 ( .A(n21270), .B(n21051), .Z(n21272) );
  IV U21390 ( .A(n21052), .Z(n21054) );
  XOR U21391 ( .A(n21054), .B(n21053), .Z(n21265) );
  NOR U21392 ( .A(n84), .B(n66), .Z(n21266) );
  IV U21393 ( .A(n21266), .Z(n21055) );
  NOR U21394 ( .A(n21265), .B(n21055), .Z(n21268) );
  IV U21395 ( .A(n21056), .Z(n21058) );
  XOR U21396 ( .A(n21058), .B(n21057), .Z(n21261) );
  NOR U21397 ( .A(n112), .B(n66), .Z(n21262) );
  IV U21398 ( .A(n21262), .Z(n21059) );
  NOR U21399 ( .A(n21261), .B(n21059), .Z(n21264) );
  IV U21400 ( .A(n21060), .Z(n21062) );
  XOR U21401 ( .A(n21062), .B(n21061), .Z(n21257) );
  NOR U21402 ( .A(n85), .B(n66), .Z(n21258) );
  IV U21403 ( .A(n21258), .Z(n21063) );
  NOR U21404 ( .A(n21257), .B(n21063), .Z(n21260) );
  IV U21405 ( .A(n21064), .Z(n21066) );
  XOR U21406 ( .A(n21066), .B(n21065), .Z(n21253) );
  NOR U21407 ( .A(n111), .B(n66), .Z(n21254) );
  IV U21408 ( .A(n21254), .Z(n21067) );
  NOR U21409 ( .A(n21253), .B(n21067), .Z(n21256) );
  IV U21410 ( .A(n21068), .Z(n21070) );
  XOR U21411 ( .A(n21070), .B(n21069), .Z(n21249) );
  NOR U21412 ( .A(n86), .B(n66), .Z(n21250) );
  IV U21413 ( .A(n21250), .Z(n21071) );
  NOR U21414 ( .A(n21249), .B(n21071), .Z(n21252) );
  IV U21415 ( .A(n21072), .Z(n21074) );
  XOR U21416 ( .A(n21074), .B(n21073), .Z(n21245) );
  NOR U21417 ( .A(n110), .B(n66), .Z(n21246) );
  IV U21418 ( .A(n21246), .Z(n21075) );
  NOR U21419 ( .A(n21245), .B(n21075), .Z(n21248) );
  IV U21420 ( .A(n21076), .Z(n21078) );
  XOR U21421 ( .A(n21078), .B(n21077), .Z(n21241) );
  NOR U21422 ( .A(n109), .B(n66), .Z(n21242) );
  IV U21423 ( .A(n21242), .Z(n21079) );
  NOR U21424 ( .A(n21241), .B(n21079), .Z(n21244) );
  XOR U21425 ( .A(n21081), .B(n21080), .Z(n21229) );
  IV U21426 ( .A(n21229), .Z(n21083) );
  NOR U21427 ( .A(n87), .B(n66), .Z(n21082) );
  IV U21428 ( .A(n21082), .Z(n21230) );
  NOR U21429 ( .A(n21083), .B(n21230), .Z(n21232) );
  IV U21430 ( .A(n21084), .Z(n21086) );
  XOR U21431 ( .A(n21086), .B(n21085), .Z(n21225) );
  NOR U21432 ( .A(n107), .B(n66), .Z(n21226) );
  IV U21433 ( .A(n21226), .Z(n21087) );
  NOR U21434 ( .A(n21225), .B(n21087), .Z(n21228) );
  IV U21435 ( .A(n21088), .Z(n21090) );
  XOR U21436 ( .A(n21090), .B(n21089), .Z(n21221) );
  NOR U21437 ( .A(n88), .B(n66), .Z(n21222) );
  IV U21438 ( .A(n21222), .Z(n21091) );
  NOR U21439 ( .A(n21221), .B(n21091), .Z(n21224) );
  IV U21440 ( .A(n21092), .Z(n21094) );
  XOR U21441 ( .A(n21094), .B(n21093), .Z(n21217) );
  NOR U21442 ( .A(n106), .B(n66), .Z(n21218) );
  IV U21443 ( .A(n21218), .Z(n21095) );
  NOR U21444 ( .A(n21217), .B(n21095), .Z(n21220) );
  XOR U21445 ( .A(n21097), .B(n21096), .Z(n21213) );
  NOR U21446 ( .A(n105), .B(n66), .Z(n21214) );
  IV U21447 ( .A(n21214), .Z(n21098) );
  NOR U21448 ( .A(n21213), .B(n21098), .Z(n21216) );
  XOR U21449 ( .A(n21100), .B(n21099), .Z(n21201) );
  IV U21450 ( .A(n21201), .Z(n21102) );
  NOR U21451 ( .A(n89), .B(n66), .Z(n21101) );
  IV U21452 ( .A(n21101), .Z(n21202) );
  NOR U21453 ( .A(n21102), .B(n21202), .Z(n21204) );
  IV U21454 ( .A(n21103), .Z(n21105) );
  XOR U21455 ( .A(n21105), .B(n21104), .Z(n21197) );
  NOR U21456 ( .A(n103), .B(n66), .Z(n21198) );
  IV U21457 ( .A(n21198), .Z(n21106) );
  NOR U21458 ( .A(n21197), .B(n21106), .Z(n21200) );
  IV U21459 ( .A(n21107), .Z(n21109) );
  XOR U21460 ( .A(n21109), .B(n21108), .Z(n21193) );
  NOR U21461 ( .A(n90), .B(n66), .Z(n21194) );
  IV U21462 ( .A(n21194), .Z(n21110) );
  NOR U21463 ( .A(n21193), .B(n21110), .Z(n21196) );
  IV U21464 ( .A(n21111), .Z(n21113) );
  XOR U21465 ( .A(n21113), .B(n21112), .Z(n21189) );
  NOR U21466 ( .A(n102), .B(n66), .Z(n21190) );
  IV U21467 ( .A(n21190), .Z(n21114) );
  NOR U21468 ( .A(n21189), .B(n21114), .Z(n21192) );
  IV U21469 ( .A(n21115), .Z(n21117) );
  XOR U21470 ( .A(n21117), .B(n21116), .Z(n21185) );
  NOR U21471 ( .A(n101), .B(n66), .Z(n21186) );
  IV U21472 ( .A(n21186), .Z(n21118) );
  NOR U21473 ( .A(n21185), .B(n21118), .Z(n21188) );
  IV U21474 ( .A(n21119), .Z(n21121) );
  XOR U21475 ( .A(n21121), .B(n21120), .Z(n21181) );
  NOR U21476 ( .A(n100), .B(n66), .Z(n21182) );
  IV U21477 ( .A(n21182), .Z(n21122) );
  NOR U21478 ( .A(n21181), .B(n21122), .Z(n21184) );
  IV U21479 ( .A(n21123), .Z(n21125) );
  XOR U21480 ( .A(n21125), .B(n21124), .Z(n21177) );
  NOR U21481 ( .A(n99), .B(n66), .Z(n21178) );
  IV U21482 ( .A(n21178), .Z(n21126) );
  NOR U21483 ( .A(n21177), .B(n21126), .Z(n21180) );
  IV U21484 ( .A(n21127), .Z(n21129) );
  XOR U21485 ( .A(n21129), .B(n21128), .Z(n21173) );
  NOR U21486 ( .A(n98), .B(n66), .Z(n21174) );
  IV U21487 ( .A(n21174), .Z(n21130) );
  NOR U21488 ( .A(n21173), .B(n21130), .Z(n21176) );
  XOR U21489 ( .A(n21132), .B(n21131), .Z(n21169) );
  NOR U21490 ( .A(n91), .B(n66), .Z(n21170) );
  IV U21491 ( .A(n21170), .Z(n21133) );
  NOR U21492 ( .A(n21169), .B(n21133), .Z(n21172) );
  XOR U21493 ( .A(n21135), .B(n21134), .Z(n21157) );
  IV U21494 ( .A(n21157), .Z(n21137) );
  NOR U21495 ( .A(n96), .B(n66), .Z(n21136) );
  IV U21496 ( .A(n21136), .Z(n21158) );
  NOR U21497 ( .A(n21137), .B(n21158), .Z(n21160) );
  NOR U21498 ( .A(n95), .B(n66), .Z(n21154) );
  IV U21499 ( .A(n21154), .Z(n21140) );
  XOR U21500 ( .A(n21139), .B(n21138), .Z(n21153) );
  NOR U21501 ( .A(n21140), .B(n21153), .Z(n21156) );
  NOR U21502 ( .A(n66), .B(n93), .Z(n22161) );
  IV U21503 ( .A(n22161), .Z(n21141) );
  NOR U21504 ( .A(n65), .B(n168), .Z(n21149) );
  IV U21505 ( .A(n21149), .Z(n21144) );
  NOR U21506 ( .A(n21141), .B(n21144), .Z(n21142) );
  IV U21507 ( .A(n21142), .Z(n21143) );
  NOR U21508 ( .A(n94), .B(n21143), .Z(n21152) );
  NOR U21509 ( .A(n21144), .B(n93), .Z(n21145) );
  XOR U21510 ( .A(n94), .B(n21145), .Z(n21146) );
  NOR U21511 ( .A(n66), .B(n21146), .Z(n21147) );
  IV U21512 ( .A(n21147), .Z(n21641) );
  XOR U21513 ( .A(n21149), .B(n21148), .Z(n21640) );
  IV U21514 ( .A(n21640), .Z(n21150) );
  NOR U21515 ( .A(n21641), .B(n21150), .Z(n21151) );
  NOR U21516 ( .A(n21152), .B(n21151), .Z(n21637) );
  XOR U21517 ( .A(n21154), .B(n21153), .Z(n21636) );
  NOR U21518 ( .A(n21637), .B(n21636), .Z(n21155) );
  NOR U21519 ( .A(n21156), .B(n21155), .Z(n21664) );
  XOR U21520 ( .A(n21158), .B(n21157), .Z(n21663) );
  NOR U21521 ( .A(n21664), .B(n21663), .Z(n21159) );
  NOR U21522 ( .A(n21160), .B(n21159), .Z(n21165) );
  XOR U21523 ( .A(n21162), .B(n21161), .Z(n21164) );
  IV U21524 ( .A(n21164), .Z(n21163) );
  NOR U21525 ( .A(n21165), .B(n21163), .Z(n21168) );
  XOR U21526 ( .A(n21165), .B(n21164), .Z(n21633) );
  NOR U21527 ( .A(n97), .B(n66), .Z(n21634) );
  IV U21528 ( .A(n21634), .Z(n21166) );
  NOR U21529 ( .A(n21633), .B(n21166), .Z(n21167) );
  NOR U21530 ( .A(n21168), .B(n21167), .Z(n21629) );
  XOR U21531 ( .A(n21170), .B(n21169), .Z(n21630) );
  NOR U21532 ( .A(n21629), .B(n21630), .Z(n21171) );
  NOR U21533 ( .A(n21172), .B(n21171), .Z(n21625) );
  XOR U21534 ( .A(n21174), .B(n21173), .Z(n21626) );
  NOR U21535 ( .A(n21625), .B(n21626), .Z(n21175) );
  NOR U21536 ( .A(n21176), .B(n21175), .Z(n21621) );
  XOR U21537 ( .A(n21178), .B(n21177), .Z(n21622) );
  NOR U21538 ( .A(n21621), .B(n21622), .Z(n21179) );
  NOR U21539 ( .A(n21180), .B(n21179), .Z(n21617) );
  XOR U21540 ( .A(n21182), .B(n21181), .Z(n21618) );
  NOR U21541 ( .A(n21617), .B(n21618), .Z(n21183) );
  NOR U21542 ( .A(n21184), .B(n21183), .Z(n21613) );
  XOR U21543 ( .A(n21186), .B(n21185), .Z(n21614) );
  NOR U21544 ( .A(n21613), .B(n21614), .Z(n21187) );
  NOR U21545 ( .A(n21188), .B(n21187), .Z(n21609) );
  XOR U21546 ( .A(n21190), .B(n21189), .Z(n21610) );
  NOR U21547 ( .A(n21609), .B(n21610), .Z(n21191) );
  NOR U21548 ( .A(n21192), .B(n21191), .Z(n21605) );
  XOR U21549 ( .A(n21194), .B(n21193), .Z(n21606) );
  NOR U21550 ( .A(n21605), .B(n21606), .Z(n21195) );
  NOR U21551 ( .A(n21196), .B(n21195), .Z(n21602) );
  XOR U21552 ( .A(n21198), .B(n21197), .Z(n21601) );
  NOR U21553 ( .A(n21602), .B(n21601), .Z(n21199) );
  NOR U21554 ( .A(n21200), .B(n21199), .Z(n21708) );
  XOR U21555 ( .A(n21202), .B(n21201), .Z(n21707) );
  NOR U21556 ( .A(n21708), .B(n21707), .Z(n21203) );
  NOR U21557 ( .A(n21204), .B(n21203), .Z(n21209) );
  XOR U21558 ( .A(n21206), .B(n21205), .Z(n21208) );
  IV U21559 ( .A(n21208), .Z(n21207) );
  NOR U21560 ( .A(n21209), .B(n21207), .Z(n21212) );
  XOR U21561 ( .A(n21209), .B(n21208), .Z(n21598) );
  NOR U21562 ( .A(n104), .B(n66), .Z(n21599) );
  IV U21563 ( .A(n21599), .Z(n21210) );
  NOR U21564 ( .A(n21598), .B(n21210), .Z(n21211) );
  NOR U21565 ( .A(n21212), .B(n21211), .Z(n21594) );
  XOR U21566 ( .A(n21214), .B(n21213), .Z(n21595) );
  NOR U21567 ( .A(n21594), .B(n21595), .Z(n21215) );
  NOR U21568 ( .A(n21216), .B(n21215), .Z(n21590) );
  XOR U21569 ( .A(n21218), .B(n21217), .Z(n21591) );
  NOR U21570 ( .A(n21590), .B(n21591), .Z(n21219) );
  NOR U21571 ( .A(n21220), .B(n21219), .Z(n21586) );
  XOR U21572 ( .A(n21222), .B(n21221), .Z(n21587) );
  NOR U21573 ( .A(n21586), .B(n21587), .Z(n21223) );
  NOR U21574 ( .A(n21224), .B(n21223), .Z(n21583) );
  XOR U21575 ( .A(n21226), .B(n21225), .Z(n21582) );
  NOR U21576 ( .A(n21583), .B(n21582), .Z(n21227) );
  NOR U21577 ( .A(n21228), .B(n21227), .Z(n21739) );
  XOR U21578 ( .A(n21230), .B(n21229), .Z(n21738) );
  NOR U21579 ( .A(n21739), .B(n21738), .Z(n21231) );
  NOR U21580 ( .A(n21232), .B(n21231), .Z(n21237) );
  XOR U21581 ( .A(n21234), .B(n21233), .Z(n21236) );
  IV U21582 ( .A(n21236), .Z(n21235) );
  NOR U21583 ( .A(n21237), .B(n21235), .Z(n21240) );
  XOR U21584 ( .A(n21237), .B(n21236), .Z(n21579) );
  NOR U21585 ( .A(n108), .B(n66), .Z(n21580) );
  IV U21586 ( .A(n21580), .Z(n21238) );
  NOR U21587 ( .A(n21579), .B(n21238), .Z(n21239) );
  NOR U21588 ( .A(n21240), .B(n21239), .Z(n21575) );
  XOR U21589 ( .A(n21242), .B(n21241), .Z(n21576) );
  NOR U21590 ( .A(n21575), .B(n21576), .Z(n21243) );
  NOR U21591 ( .A(n21244), .B(n21243), .Z(n21571) );
  XOR U21592 ( .A(n21246), .B(n21245), .Z(n21572) );
  NOR U21593 ( .A(n21571), .B(n21572), .Z(n21247) );
  NOR U21594 ( .A(n21248), .B(n21247), .Z(n21567) );
  XOR U21595 ( .A(n21250), .B(n21249), .Z(n21568) );
  NOR U21596 ( .A(n21567), .B(n21568), .Z(n21251) );
  NOR U21597 ( .A(n21252), .B(n21251), .Z(n21563) );
  XOR U21598 ( .A(n21254), .B(n21253), .Z(n21564) );
  NOR U21599 ( .A(n21563), .B(n21564), .Z(n21255) );
  NOR U21600 ( .A(n21256), .B(n21255), .Z(n21559) );
  XOR U21601 ( .A(n21258), .B(n21257), .Z(n21560) );
  NOR U21602 ( .A(n21559), .B(n21560), .Z(n21259) );
  NOR U21603 ( .A(n21260), .B(n21259), .Z(n21555) );
  XOR U21604 ( .A(n21262), .B(n21261), .Z(n21556) );
  NOR U21605 ( .A(n21555), .B(n21556), .Z(n21263) );
  NOR U21606 ( .A(n21264), .B(n21263), .Z(n21551) );
  XOR U21607 ( .A(n21266), .B(n21265), .Z(n21552) );
  NOR U21608 ( .A(n21551), .B(n21552), .Z(n21267) );
  NOR U21609 ( .A(n21268), .B(n21267), .Z(n21550) );
  XOR U21610 ( .A(n21270), .B(n21269), .Z(n21549) );
  NOR U21611 ( .A(n21550), .B(n21549), .Z(n21271) );
  NOR U21612 ( .A(n21272), .B(n21271), .Z(n21273) );
  IV U21613 ( .A(n21273), .Z(n21547) );
  XOR U21614 ( .A(n21275), .B(n21274), .Z(n21276) );
  IV U21615 ( .A(n21276), .Z(n21546) );
  NOR U21616 ( .A(n21547), .B(n21546), .Z(n21277) );
  NOR U21617 ( .A(n21278), .B(n21277), .Z(n21279) );
  IV U21618 ( .A(n21279), .Z(n21545) );
  XOR U21619 ( .A(n21281), .B(n21280), .Z(n21544) );
  NOR U21620 ( .A(n21545), .B(n21544), .Z(n21282) );
  NOR U21621 ( .A(n21283), .B(n21282), .Z(n21284) );
  IV U21622 ( .A(n21284), .Z(n21541) );
  NOR U21623 ( .A(n21542), .B(n21541), .Z(n21285) );
  NOR U21624 ( .A(n21286), .B(n21285), .Z(n21287) );
  IV U21625 ( .A(n21287), .Z(n21540) );
  XOR U21626 ( .A(n21289), .B(n21288), .Z(n21539) );
  NOR U21627 ( .A(n21540), .B(n21539), .Z(n21290) );
  NOR U21628 ( .A(n21291), .B(n21290), .Z(n21292) );
  IV U21629 ( .A(n21292), .Z(n21537) );
  XOR U21630 ( .A(n21294), .B(n21293), .Z(n21295) );
  IV U21631 ( .A(n21295), .Z(n21536) );
  NOR U21632 ( .A(n21537), .B(n21536), .Z(n21296) );
  NOR U21633 ( .A(n21297), .B(n21296), .Z(n21298) );
  IV U21634 ( .A(n21298), .Z(n21535) );
  XOR U21635 ( .A(n21300), .B(n21299), .Z(n21534) );
  NOR U21636 ( .A(n21535), .B(n21534), .Z(n21301) );
  NOR U21637 ( .A(n21302), .B(n21301), .Z(n21303) );
  IV U21638 ( .A(n21303), .Z(n21532) );
  XOR U21639 ( .A(n21305), .B(n21304), .Z(n21306) );
  IV U21640 ( .A(n21306), .Z(n21531) );
  NOR U21641 ( .A(n21532), .B(n21531), .Z(n21307) );
  NOR U21642 ( .A(n21308), .B(n21307), .Z(n21309) );
  IV U21643 ( .A(n21309), .Z(n21530) );
  XOR U21644 ( .A(n21311), .B(n21310), .Z(n21529) );
  NOR U21645 ( .A(n21530), .B(n21529), .Z(n21312) );
  NOR U21646 ( .A(n21313), .B(n21312), .Z(n21314) );
  IV U21647 ( .A(n21314), .Z(n21527) );
  XOR U21648 ( .A(n21316), .B(n21315), .Z(n21317) );
  IV U21649 ( .A(n21317), .Z(n21526) );
  NOR U21650 ( .A(n21527), .B(n21526), .Z(n21318) );
  NOR U21651 ( .A(n21319), .B(n21318), .Z(n21320) );
  IV U21652 ( .A(n21320), .Z(n21525) );
  XOR U21653 ( .A(n21322), .B(n21321), .Z(n21524) );
  NOR U21654 ( .A(n21525), .B(n21524), .Z(n21323) );
  NOR U21655 ( .A(n21324), .B(n21323), .Z(n21325) );
  IV U21656 ( .A(n21325), .Z(n21522) );
  XOR U21657 ( .A(n21327), .B(n21326), .Z(n21328) );
  IV U21658 ( .A(n21328), .Z(n21521) );
  NOR U21659 ( .A(n21522), .B(n21521), .Z(n21329) );
  NOR U21660 ( .A(n21330), .B(n21329), .Z(n21331) );
  IV U21661 ( .A(n21331), .Z(n21520) );
  XOR U21662 ( .A(n21333), .B(n21332), .Z(n21519) );
  NOR U21663 ( .A(n21520), .B(n21519), .Z(n21334) );
  NOR U21664 ( .A(n21335), .B(n21334), .Z(n21336) );
  IV U21665 ( .A(n21336), .Z(n21517) );
  XOR U21666 ( .A(n21338), .B(n21337), .Z(n21339) );
  IV U21667 ( .A(n21339), .Z(n21516) );
  NOR U21668 ( .A(n21517), .B(n21516), .Z(n21340) );
  NOR U21669 ( .A(n21341), .B(n21340), .Z(n21342) );
  IV U21670 ( .A(n21342), .Z(n21515) );
  XOR U21671 ( .A(n21344), .B(n21343), .Z(n21514) );
  NOR U21672 ( .A(n21515), .B(n21514), .Z(n21345) );
  NOR U21673 ( .A(n21346), .B(n21345), .Z(n21512) );
  IV U21674 ( .A(n21512), .Z(n21347) );
  NOR U21675 ( .A(n21348), .B(n21347), .Z(n21349) );
  NOR U21676 ( .A(n21350), .B(n21349), .Z(n21352) );
  IV U21677 ( .A(n21352), .Z(n21351) );
  NOR U21678 ( .A(n21353), .B(n21351), .Z(n21358) );
  XOR U21679 ( .A(n21353), .B(n21352), .Z(n21508) );
  XOR U21680 ( .A(n21355), .B(n21354), .Z(n21356) );
  IV U21681 ( .A(n21356), .Z(n21507) );
  NOR U21682 ( .A(n21508), .B(n21507), .Z(n21357) );
  NOR U21683 ( .A(n21358), .B(n21357), .Z(n21501) );
  XOR U21684 ( .A(n21360), .B(n21359), .Z(n21502) );
  NOR U21685 ( .A(n21501), .B(n21502), .Z(n21361) );
  NOR U21686 ( .A(n21362), .B(n21361), .Z(n21500) );
  XOR U21687 ( .A(n21364), .B(n21363), .Z(n21499) );
  NOR U21688 ( .A(n21500), .B(n21499), .Z(n21365) );
  NOR U21689 ( .A(n21366), .B(n21365), .Z(n21495) );
  NOR U21690 ( .A(n21367), .B(n21495), .Z(n21368) );
  NOR U21691 ( .A(n21369), .B(n21368), .Z(n21371) );
  NOR U21692 ( .A(n139), .B(n66), .Z(n21372) );
  IV U21693 ( .A(n21372), .Z(n21370) );
  NOR U21694 ( .A(n21371), .B(n21370), .Z(n21376) );
  XOR U21695 ( .A(n21372), .B(n21371), .Z(n21491) );
  XOR U21696 ( .A(n21374), .B(n21373), .Z(n21490) );
  NOR U21697 ( .A(n21491), .B(n21490), .Z(n21375) );
  NOR U21698 ( .A(n21376), .B(n21375), .Z(n21889) );
  XOR U21699 ( .A(n21378), .B(n21377), .Z(n21890) );
  NOR U21700 ( .A(n21889), .B(n21890), .Z(n21379) );
  NOR U21701 ( .A(n21380), .B(n21379), .Z(n21385) );
  XOR U21702 ( .A(n21382), .B(n21381), .Z(n21384) );
  IV U21703 ( .A(n21384), .Z(n21383) );
  NOR U21704 ( .A(n21385), .B(n21383), .Z(n21388) );
  XOR U21705 ( .A(n21385), .B(n21384), .Z(n21897) );
  NOR U21706 ( .A(n143), .B(n66), .Z(n21898) );
  IV U21707 ( .A(n21898), .Z(n21386) );
  NOR U21708 ( .A(n21897), .B(n21386), .Z(n21387) );
  NOR U21709 ( .A(n21388), .B(n21387), .Z(n21393) );
  NOR U21710 ( .A(n145), .B(n66), .Z(n21392) );
  IV U21711 ( .A(n21392), .Z(n21389) );
  NOR U21712 ( .A(n21393), .B(n21389), .Z(n21395) );
  XOR U21713 ( .A(n21391), .B(n21390), .Z(n21907) );
  XOR U21714 ( .A(n21393), .B(n21392), .Z(n21906) );
  NOR U21715 ( .A(n21907), .B(n21906), .Z(n21394) );
  NOR U21716 ( .A(n21395), .B(n21394), .Z(n21398) );
  NOR U21717 ( .A(n147), .B(n66), .Z(n21397) );
  IV U21718 ( .A(n21397), .Z(n21396) );
  NOR U21719 ( .A(n21398), .B(n21396), .Z(n21402) );
  XOR U21720 ( .A(n21398), .B(n21397), .Z(n21911) );
  XOR U21721 ( .A(n21400), .B(n21399), .Z(n21912) );
  NOR U21722 ( .A(n21911), .B(n21912), .Z(n21401) );
  NOR U21723 ( .A(n21402), .B(n21401), .Z(n21405) );
  NOR U21724 ( .A(n148), .B(n66), .Z(n21404) );
  IV U21725 ( .A(n21404), .Z(n21403) );
  NOR U21726 ( .A(n21405), .B(n21403), .Z(n21410) );
  XOR U21727 ( .A(n21405), .B(n21404), .Z(n21922) );
  XOR U21728 ( .A(n21407), .B(n21406), .Z(n21923) );
  IV U21729 ( .A(n21923), .Z(n21408) );
  NOR U21730 ( .A(n21922), .B(n21408), .Z(n21409) );
  NOR U21731 ( .A(n21410), .B(n21409), .Z(n21417) );
  NOR U21732 ( .A(n150), .B(n66), .Z(n21416) );
  IV U21733 ( .A(n21416), .Z(n21411) );
  NOR U21734 ( .A(n21417), .B(n21411), .Z(n21420) );
  XOR U21735 ( .A(n21413), .B(n21412), .Z(n21414) );
  XOR U21736 ( .A(n21415), .B(n21414), .Z(n21928) );
  IV U21737 ( .A(n21928), .Z(n21418) );
  XOR U21738 ( .A(n21417), .B(n21416), .Z(n21927) );
  NOR U21739 ( .A(n21418), .B(n21927), .Z(n21419) );
  NOR U21740 ( .A(n21420), .B(n21419), .Z(n21425) );
  NOR U21741 ( .A(n153), .B(n66), .Z(n21424) );
  IV U21742 ( .A(n21424), .Z(n21421) );
  NOR U21743 ( .A(n21425), .B(n21421), .Z(n21427) );
  XOR U21744 ( .A(n21423), .B(n21422), .Z(n21489) );
  XOR U21745 ( .A(n21425), .B(n21424), .Z(n21488) );
  NOR U21746 ( .A(n21489), .B(n21488), .Z(n21426) );
  NOR U21747 ( .A(n21427), .B(n21426), .Z(n21432) );
  XOR U21748 ( .A(n21429), .B(n21428), .Z(n21431) );
  IV U21749 ( .A(n21431), .Z(n21430) );
  NOR U21750 ( .A(n21432), .B(n21430), .Z(n21435) );
  XOR U21751 ( .A(n21432), .B(n21431), .Z(n21941) );
  NOR U21752 ( .A(n155), .B(n66), .Z(n21433) );
  IV U21753 ( .A(n21433), .Z(n21940) );
  NOR U21754 ( .A(n21941), .B(n21940), .Z(n21434) );
  NOR U21755 ( .A(n21435), .B(n21434), .Z(n21437) );
  IV U21756 ( .A(n21437), .Z(n21947) );
  NOR U21757 ( .A(n21436), .B(n21947), .Z(n21442) );
  IV U21758 ( .A(n21436), .Z(n21948) );
  NOR U21759 ( .A(n21437), .B(n21948), .Z(n21440) );
  XOR U21760 ( .A(n21439), .B(n21438), .Z(n21950) );
  NOR U21761 ( .A(n21440), .B(n21950), .Z(n21441) );
  NOR U21762 ( .A(n21442), .B(n21441), .Z(n21446) );
  IV U21763 ( .A(n21446), .Z(n21444) );
  NOR U21764 ( .A(n158), .B(n66), .Z(n21443) );
  IV U21765 ( .A(n21443), .Z(n21445) );
  NOR U21766 ( .A(n21444), .B(n21445), .Z(n21450) );
  XOR U21767 ( .A(n21446), .B(n21445), .Z(n21956) );
  XOR U21768 ( .A(n21448), .B(n21447), .Z(n21955) );
  NOR U21769 ( .A(n21956), .B(n21955), .Z(n21449) );
  NOR U21770 ( .A(n21450), .B(n21449), .Z(n21455) );
  XOR U21771 ( .A(n21452), .B(n21451), .Z(n21454) );
  IV U21772 ( .A(n21454), .Z(n21453) );
  NOR U21773 ( .A(n21455), .B(n21453), .Z(n21458) );
  XOR U21774 ( .A(n21455), .B(n21454), .Z(n21966) );
  NOR U21775 ( .A(n161), .B(n66), .Z(n21967) );
  IV U21776 ( .A(n21967), .Z(n21456) );
  NOR U21777 ( .A(n21966), .B(n21456), .Z(n21457) );
  NOR U21778 ( .A(n21458), .B(n21457), .Z(n21460) );
  IV U21779 ( .A(n21460), .Z(n21971) );
  NOR U21780 ( .A(n21459), .B(n21971), .Z(n21465) );
  IV U21781 ( .A(n21459), .Z(n21972) );
  NOR U21782 ( .A(n21460), .B(n21972), .Z(n21463) );
  XOR U21783 ( .A(n21462), .B(n21461), .Z(n21974) );
  NOR U21784 ( .A(n21463), .B(n21974), .Z(n21464) );
  NOR U21785 ( .A(n21465), .B(n21464), .Z(n21473) );
  IV U21786 ( .A(n21473), .Z(n21467) );
  NOR U21787 ( .A(n165), .B(n66), .Z(n21466) );
  IV U21788 ( .A(n21466), .Z(n21472) );
  NOR U21789 ( .A(n21467), .B(n21472), .Z(n21475) );
  XOR U21790 ( .A(n21469), .B(n21468), .Z(n21470) );
  XOR U21791 ( .A(n21471), .B(n21470), .Z(n21979) );
  XOR U21792 ( .A(n21473), .B(n21472), .Z(n21980) );
  NOR U21793 ( .A(n21979), .B(n21980), .Z(n21474) );
  NOR U21794 ( .A(n21475), .B(n21474), .Z(n21480) );
  XOR U21795 ( .A(n21477), .B(n21476), .Z(n21479) );
  IV U21796 ( .A(n21479), .Z(n21478) );
  NOR U21797 ( .A(n21480), .B(n21478), .Z(n21483) );
  XOR U21798 ( .A(n21480), .B(n21479), .Z(n21987) );
  NOR U21799 ( .A(n167), .B(n66), .Z(n21988) );
  IV U21800 ( .A(n21988), .Z(n21481) );
  NOR U21801 ( .A(n21987), .B(n21481), .Z(n21482) );
  NOR U21802 ( .A(n21483), .B(n21482), .Z(n21990) );
  XOR U21803 ( .A(n21485), .B(n21484), .Z(n21989) );
  NOR U21804 ( .A(n21990), .B(n21989), .Z(n28540) );
  XOR U21805 ( .A(n21487), .B(n21486), .Z(n28539) );
  NOR U21806 ( .A(n28540), .B(n28539), .Z(n28543) );
  NOR U21807 ( .A(n156), .B(n67), .Z(n21938) );
  XOR U21808 ( .A(n21489), .B(n21488), .Z(n21935) );
  XOR U21809 ( .A(n21491), .B(n21490), .Z(n21882) );
  NOR U21810 ( .A(n141), .B(n67), .Z(n21883) );
  NOR U21811 ( .A(n21882), .B(n21883), .Z(n21886) );
  XOR U21812 ( .A(n21493), .B(n21492), .Z(n21494) );
  XOR U21813 ( .A(n21495), .B(n21494), .Z(n21498) );
  NOR U21814 ( .A(n139), .B(n67), .Z(n21497) );
  IV U21815 ( .A(n21497), .Z(n21496) );
  NOR U21816 ( .A(n21498), .B(n21496), .Z(n21880) );
  XOR U21817 ( .A(n21498), .B(n21497), .Z(n22000) );
  XOR U21818 ( .A(n21500), .B(n21499), .Z(n21873) );
  NOR U21819 ( .A(n137), .B(n67), .Z(n21874) );
  NOR U21820 ( .A(n21873), .B(n21874), .Z(n21877) );
  XOR U21821 ( .A(n21502), .B(n21501), .Z(n21503) );
  IV U21822 ( .A(n21503), .Z(n21505) );
  NOR U21823 ( .A(n135), .B(n67), .Z(n21506) );
  IV U21824 ( .A(n21506), .Z(n21504) );
  NOR U21825 ( .A(n21505), .B(n21504), .Z(n21871) );
  XOR U21826 ( .A(n21506), .B(n21505), .Z(n22006) );
  XOR U21827 ( .A(n21508), .B(n21507), .Z(n21864) );
  NOR U21828 ( .A(n133), .B(n67), .Z(n21865) );
  NOR U21829 ( .A(n21864), .B(n21865), .Z(n21868) );
  XOR U21830 ( .A(n21510), .B(n21509), .Z(n21511) );
  XOR U21831 ( .A(n21512), .B(n21511), .Z(n21860) );
  NOR U21832 ( .A(n131), .B(n67), .Z(n21859) );
  IV U21833 ( .A(n21859), .Z(n21513) );
  NOR U21834 ( .A(n21860), .B(n21513), .Z(n21862) );
  NOR U21835 ( .A(n128), .B(n67), .Z(n21854) );
  XOR U21836 ( .A(n21515), .B(n21514), .Z(n21853) );
  NOR U21837 ( .A(n21854), .B(n21853), .Z(n21857) );
  XOR U21838 ( .A(n21517), .B(n21516), .Z(n21849) );
  NOR U21839 ( .A(n126), .B(n67), .Z(n21848) );
  IV U21840 ( .A(n21848), .Z(n21518) );
  NOR U21841 ( .A(n21849), .B(n21518), .Z(n21851) );
  NOR U21842 ( .A(n125), .B(n67), .Z(n21843) );
  XOR U21843 ( .A(n21520), .B(n21519), .Z(n21842) );
  NOR U21844 ( .A(n21843), .B(n21842), .Z(n21846) );
  XOR U21845 ( .A(n21522), .B(n21521), .Z(n21838) );
  NOR U21846 ( .A(n123), .B(n67), .Z(n21837) );
  IV U21847 ( .A(n21837), .Z(n21523) );
  NOR U21848 ( .A(n21838), .B(n21523), .Z(n21840) );
  NOR U21849 ( .A(n120), .B(n67), .Z(n21832) );
  XOR U21850 ( .A(n21525), .B(n21524), .Z(n21831) );
  NOR U21851 ( .A(n21832), .B(n21831), .Z(n21835) );
  XOR U21852 ( .A(n21527), .B(n21526), .Z(n21827) );
  NOR U21853 ( .A(n119), .B(n67), .Z(n21826) );
  IV U21854 ( .A(n21826), .Z(n21528) );
  NOR U21855 ( .A(n21827), .B(n21528), .Z(n21829) );
  NOR U21856 ( .A(n79), .B(n67), .Z(n21821) );
  XOR U21857 ( .A(n21530), .B(n21529), .Z(n21820) );
  NOR U21858 ( .A(n21821), .B(n21820), .Z(n21824) );
  XOR U21859 ( .A(n21532), .B(n21531), .Z(n21816) );
  NOR U21860 ( .A(n117), .B(n67), .Z(n21815) );
  IV U21861 ( .A(n21815), .Z(n21533) );
  NOR U21862 ( .A(n21816), .B(n21533), .Z(n21818) );
  NOR U21863 ( .A(n80), .B(n67), .Z(n21810) );
  XOR U21864 ( .A(n21535), .B(n21534), .Z(n21809) );
  NOR U21865 ( .A(n21810), .B(n21809), .Z(n21813) );
  XOR U21866 ( .A(n21537), .B(n21536), .Z(n21805) );
  NOR U21867 ( .A(n116), .B(n67), .Z(n21804) );
  IV U21868 ( .A(n21804), .Z(n21538) );
  NOR U21869 ( .A(n21805), .B(n21538), .Z(n21807) );
  NOR U21870 ( .A(n81), .B(n67), .Z(n21799) );
  XOR U21871 ( .A(n21540), .B(n21539), .Z(n21798) );
  NOR U21872 ( .A(n21799), .B(n21798), .Z(n21802) );
  XOR U21873 ( .A(n21542), .B(n21541), .Z(n21794) );
  NOR U21874 ( .A(n115), .B(n67), .Z(n21793) );
  IV U21875 ( .A(n21793), .Z(n21543) );
  NOR U21876 ( .A(n21794), .B(n21543), .Z(n21796) );
  NOR U21877 ( .A(n82), .B(n67), .Z(n21788) );
  XOR U21878 ( .A(n21545), .B(n21544), .Z(n21787) );
  NOR U21879 ( .A(n21788), .B(n21787), .Z(n21791) );
  XOR U21880 ( .A(n21547), .B(n21546), .Z(n21783) );
  NOR U21881 ( .A(n114), .B(n67), .Z(n21782) );
  IV U21882 ( .A(n21782), .Z(n21548) );
  NOR U21883 ( .A(n21783), .B(n21548), .Z(n21785) );
  NOR U21884 ( .A(n83), .B(n67), .Z(n21777) );
  XOR U21885 ( .A(n21550), .B(n21549), .Z(n21776) );
  NOR U21886 ( .A(n21777), .B(n21776), .Z(n21780) );
  IV U21887 ( .A(n21551), .Z(n21553) );
  XOR U21888 ( .A(n21553), .B(n21552), .Z(n21771) );
  NOR U21889 ( .A(n113), .B(n67), .Z(n21772) );
  IV U21890 ( .A(n21772), .Z(n21554) );
  NOR U21891 ( .A(n21771), .B(n21554), .Z(n21774) );
  IV U21892 ( .A(n21555), .Z(n21557) );
  XOR U21893 ( .A(n21557), .B(n21556), .Z(n21767) );
  NOR U21894 ( .A(n84), .B(n67), .Z(n21768) );
  IV U21895 ( .A(n21768), .Z(n21558) );
  NOR U21896 ( .A(n21767), .B(n21558), .Z(n21770) );
  IV U21897 ( .A(n21559), .Z(n21561) );
  XOR U21898 ( .A(n21561), .B(n21560), .Z(n21763) );
  NOR U21899 ( .A(n112), .B(n67), .Z(n21764) );
  IV U21900 ( .A(n21764), .Z(n21562) );
  NOR U21901 ( .A(n21763), .B(n21562), .Z(n21766) );
  IV U21902 ( .A(n21563), .Z(n21565) );
  XOR U21903 ( .A(n21565), .B(n21564), .Z(n21759) );
  NOR U21904 ( .A(n85), .B(n67), .Z(n21760) );
  IV U21905 ( .A(n21760), .Z(n21566) );
  NOR U21906 ( .A(n21759), .B(n21566), .Z(n21762) );
  IV U21907 ( .A(n21567), .Z(n21569) );
  XOR U21908 ( .A(n21569), .B(n21568), .Z(n21755) );
  NOR U21909 ( .A(n111), .B(n67), .Z(n21756) );
  IV U21910 ( .A(n21756), .Z(n21570) );
  NOR U21911 ( .A(n21755), .B(n21570), .Z(n21758) );
  IV U21912 ( .A(n21571), .Z(n21573) );
  XOR U21913 ( .A(n21573), .B(n21572), .Z(n21751) );
  NOR U21914 ( .A(n86), .B(n67), .Z(n21752) );
  IV U21915 ( .A(n21752), .Z(n21574) );
  NOR U21916 ( .A(n21751), .B(n21574), .Z(n21754) );
  IV U21917 ( .A(n21575), .Z(n21577) );
  XOR U21918 ( .A(n21577), .B(n21576), .Z(n21747) );
  NOR U21919 ( .A(n110), .B(n67), .Z(n21748) );
  IV U21920 ( .A(n21748), .Z(n21578) );
  NOR U21921 ( .A(n21747), .B(n21578), .Z(n21750) );
  XOR U21922 ( .A(n21580), .B(n21579), .Z(n21743) );
  NOR U21923 ( .A(n109), .B(n67), .Z(n21744) );
  IV U21924 ( .A(n21744), .Z(n21581) );
  NOR U21925 ( .A(n21743), .B(n21581), .Z(n21746) );
  XOR U21926 ( .A(n21583), .B(n21582), .Z(n21731) );
  IV U21927 ( .A(n21731), .Z(n21585) );
  NOR U21928 ( .A(n87), .B(n67), .Z(n21584) );
  IV U21929 ( .A(n21584), .Z(n21732) );
  NOR U21930 ( .A(n21585), .B(n21732), .Z(n21734) );
  IV U21931 ( .A(n21586), .Z(n21588) );
  XOR U21932 ( .A(n21588), .B(n21587), .Z(n21727) );
  NOR U21933 ( .A(n107), .B(n67), .Z(n21728) );
  IV U21934 ( .A(n21728), .Z(n21589) );
  NOR U21935 ( .A(n21727), .B(n21589), .Z(n21730) );
  IV U21936 ( .A(n21590), .Z(n21592) );
  XOR U21937 ( .A(n21592), .B(n21591), .Z(n21723) );
  NOR U21938 ( .A(n88), .B(n67), .Z(n21724) );
  IV U21939 ( .A(n21724), .Z(n21593) );
  NOR U21940 ( .A(n21723), .B(n21593), .Z(n21726) );
  IV U21941 ( .A(n21594), .Z(n21596) );
  XOR U21942 ( .A(n21596), .B(n21595), .Z(n21719) );
  NOR U21943 ( .A(n106), .B(n67), .Z(n21720) );
  IV U21944 ( .A(n21720), .Z(n21597) );
  NOR U21945 ( .A(n21719), .B(n21597), .Z(n21722) );
  XOR U21946 ( .A(n21599), .B(n21598), .Z(n21715) );
  NOR U21947 ( .A(n105), .B(n67), .Z(n21716) );
  IV U21948 ( .A(n21716), .Z(n21600) );
  NOR U21949 ( .A(n21715), .B(n21600), .Z(n21718) );
  XOR U21950 ( .A(n21602), .B(n21601), .Z(n21703) );
  IV U21951 ( .A(n21703), .Z(n21604) );
  NOR U21952 ( .A(n89), .B(n67), .Z(n21603) );
  IV U21953 ( .A(n21603), .Z(n21704) );
  NOR U21954 ( .A(n21604), .B(n21704), .Z(n21706) );
  IV U21955 ( .A(n21605), .Z(n21607) );
  XOR U21956 ( .A(n21607), .B(n21606), .Z(n21699) );
  NOR U21957 ( .A(n103), .B(n67), .Z(n21700) );
  IV U21958 ( .A(n21700), .Z(n21608) );
  NOR U21959 ( .A(n21699), .B(n21608), .Z(n21702) );
  IV U21960 ( .A(n21609), .Z(n21611) );
  XOR U21961 ( .A(n21611), .B(n21610), .Z(n21695) );
  NOR U21962 ( .A(n90), .B(n67), .Z(n21696) );
  IV U21963 ( .A(n21696), .Z(n21612) );
  NOR U21964 ( .A(n21695), .B(n21612), .Z(n21698) );
  IV U21965 ( .A(n21613), .Z(n21615) );
  XOR U21966 ( .A(n21615), .B(n21614), .Z(n21691) );
  NOR U21967 ( .A(n102), .B(n67), .Z(n21692) );
  IV U21968 ( .A(n21692), .Z(n21616) );
  NOR U21969 ( .A(n21691), .B(n21616), .Z(n21694) );
  IV U21970 ( .A(n21617), .Z(n21619) );
  XOR U21971 ( .A(n21619), .B(n21618), .Z(n21687) );
  NOR U21972 ( .A(n101), .B(n67), .Z(n21688) );
  IV U21973 ( .A(n21688), .Z(n21620) );
  NOR U21974 ( .A(n21687), .B(n21620), .Z(n21690) );
  IV U21975 ( .A(n21621), .Z(n21623) );
  XOR U21976 ( .A(n21623), .B(n21622), .Z(n21683) );
  NOR U21977 ( .A(n100), .B(n67), .Z(n21684) );
  IV U21978 ( .A(n21684), .Z(n21624) );
  NOR U21979 ( .A(n21683), .B(n21624), .Z(n21686) );
  IV U21980 ( .A(n21625), .Z(n21627) );
  XOR U21981 ( .A(n21627), .B(n21626), .Z(n21679) );
  NOR U21982 ( .A(n99), .B(n67), .Z(n21680) );
  IV U21983 ( .A(n21680), .Z(n21628) );
  NOR U21984 ( .A(n21679), .B(n21628), .Z(n21682) );
  IV U21985 ( .A(n21629), .Z(n21631) );
  XOR U21986 ( .A(n21631), .B(n21630), .Z(n21675) );
  NOR U21987 ( .A(n98), .B(n67), .Z(n21676) );
  IV U21988 ( .A(n21676), .Z(n21632) );
  NOR U21989 ( .A(n21675), .B(n21632), .Z(n21678) );
  XOR U21990 ( .A(n21634), .B(n21633), .Z(n21671) );
  NOR U21991 ( .A(n91), .B(n67), .Z(n21672) );
  IV U21992 ( .A(n21672), .Z(n21635) );
  NOR U21993 ( .A(n21671), .B(n21635), .Z(n21674) );
  XOR U21994 ( .A(n21637), .B(n21636), .Z(n21659) );
  IV U21995 ( .A(n21659), .Z(n21639) );
  NOR U21996 ( .A(n96), .B(n67), .Z(n21638) );
  IV U21997 ( .A(n21638), .Z(n21660) );
  NOR U21998 ( .A(n21639), .B(n21660), .Z(n21662) );
  NOR U21999 ( .A(n95), .B(n67), .Z(n21656) );
  IV U22000 ( .A(n21656), .Z(n21642) );
  XOR U22001 ( .A(n21641), .B(n21640), .Z(n21655) );
  NOR U22002 ( .A(n21642), .B(n21655), .Z(n21658) );
  NOR U22003 ( .A(n67), .B(n93), .Z(n22670) );
  IV U22004 ( .A(n22670), .Z(n21643) );
  NOR U22005 ( .A(n66), .B(n168), .Z(n21651) );
  IV U22006 ( .A(n21651), .Z(n21646) );
  NOR U22007 ( .A(n21643), .B(n21646), .Z(n21644) );
  IV U22008 ( .A(n21644), .Z(n21645) );
  NOR U22009 ( .A(n94), .B(n21645), .Z(n21654) );
  NOR U22010 ( .A(n21646), .B(n93), .Z(n21647) );
  XOR U22011 ( .A(n94), .B(n21647), .Z(n21648) );
  NOR U22012 ( .A(n67), .B(n21648), .Z(n21649) );
  IV U22013 ( .A(n21649), .Z(n22152) );
  XOR U22014 ( .A(n21651), .B(n21650), .Z(n22151) );
  IV U22015 ( .A(n22151), .Z(n21652) );
  NOR U22016 ( .A(n22152), .B(n21652), .Z(n21653) );
  NOR U22017 ( .A(n21654), .B(n21653), .Z(n22148) );
  XOR U22018 ( .A(n21656), .B(n21655), .Z(n22147) );
  NOR U22019 ( .A(n22148), .B(n22147), .Z(n21657) );
  NOR U22020 ( .A(n21658), .B(n21657), .Z(n22175) );
  XOR U22021 ( .A(n21660), .B(n21659), .Z(n22174) );
  NOR U22022 ( .A(n22175), .B(n22174), .Z(n21661) );
  NOR U22023 ( .A(n21662), .B(n21661), .Z(n21667) );
  XOR U22024 ( .A(n21664), .B(n21663), .Z(n21666) );
  IV U22025 ( .A(n21666), .Z(n21665) );
  NOR U22026 ( .A(n21667), .B(n21665), .Z(n21670) );
  XOR U22027 ( .A(n21667), .B(n21666), .Z(n22144) );
  NOR U22028 ( .A(n97), .B(n67), .Z(n22145) );
  IV U22029 ( .A(n22145), .Z(n21668) );
  NOR U22030 ( .A(n22144), .B(n21668), .Z(n21669) );
  NOR U22031 ( .A(n21670), .B(n21669), .Z(n22140) );
  XOR U22032 ( .A(n21672), .B(n21671), .Z(n22141) );
  NOR U22033 ( .A(n22140), .B(n22141), .Z(n21673) );
  NOR U22034 ( .A(n21674), .B(n21673), .Z(n22136) );
  XOR U22035 ( .A(n21676), .B(n21675), .Z(n22137) );
  NOR U22036 ( .A(n22136), .B(n22137), .Z(n21677) );
  NOR U22037 ( .A(n21678), .B(n21677), .Z(n22132) );
  XOR U22038 ( .A(n21680), .B(n21679), .Z(n22133) );
  NOR U22039 ( .A(n22132), .B(n22133), .Z(n21681) );
  NOR U22040 ( .A(n21682), .B(n21681), .Z(n22128) );
  XOR U22041 ( .A(n21684), .B(n21683), .Z(n22129) );
  NOR U22042 ( .A(n22128), .B(n22129), .Z(n21685) );
  NOR U22043 ( .A(n21686), .B(n21685), .Z(n22124) );
  XOR U22044 ( .A(n21688), .B(n21687), .Z(n22125) );
  NOR U22045 ( .A(n22124), .B(n22125), .Z(n21689) );
  NOR U22046 ( .A(n21690), .B(n21689), .Z(n22120) );
  XOR U22047 ( .A(n21692), .B(n21691), .Z(n22121) );
  NOR U22048 ( .A(n22120), .B(n22121), .Z(n21693) );
  NOR U22049 ( .A(n21694), .B(n21693), .Z(n22116) );
  XOR U22050 ( .A(n21696), .B(n21695), .Z(n22117) );
  NOR U22051 ( .A(n22116), .B(n22117), .Z(n21697) );
  NOR U22052 ( .A(n21698), .B(n21697), .Z(n22113) );
  XOR U22053 ( .A(n21700), .B(n21699), .Z(n22112) );
  NOR U22054 ( .A(n22113), .B(n22112), .Z(n21701) );
  NOR U22055 ( .A(n21702), .B(n21701), .Z(n22219) );
  XOR U22056 ( .A(n21704), .B(n21703), .Z(n22218) );
  NOR U22057 ( .A(n22219), .B(n22218), .Z(n21705) );
  NOR U22058 ( .A(n21706), .B(n21705), .Z(n21711) );
  XOR U22059 ( .A(n21708), .B(n21707), .Z(n21710) );
  IV U22060 ( .A(n21710), .Z(n21709) );
  NOR U22061 ( .A(n21711), .B(n21709), .Z(n21714) );
  XOR U22062 ( .A(n21711), .B(n21710), .Z(n22109) );
  NOR U22063 ( .A(n104), .B(n67), .Z(n22110) );
  IV U22064 ( .A(n22110), .Z(n21712) );
  NOR U22065 ( .A(n22109), .B(n21712), .Z(n21713) );
  NOR U22066 ( .A(n21714), .B(n21713), .Z(n22105) );
  XOR U22067 ( .A(n21716), .B(n21715), .Z(n22106) );
  NOR U22068 ( .A(n22105), .B(n22106), .Z(n21717) );
  NOR U22069 ( .A(n21718), .B(n21717), .Z(n22101) );
  XOR U22070 ( .A(n21720), .B(n21719), .Z(n22102) );
  NOR U22071 ( .A(n22101), .B(n22102), .Z(n21721) );
  NOR U22072 ( .A(n21722), .B(n21721), .Z(n22097) );
  XOR U22073 ( .A(n21724), .B(n21723), .Z(n22098) );
  NOR U22074 ( .A(n22097), .B(n22098), .Z(n21725) );
  NOR U22075 ( .A(n21726), .B(n21725), .Z(n22094) );
  XOR U22076 ( .A(n21728), .B(n21727), .Z(n22093) );
  NOR U22077 ( .A(n22094), .B(n22093), .Z(n21729) );
  NOR U22078 ( .A(n21730), .B(n21729), .Z(n22247) );
  XOR U22079 ( .A(n21732), .B(n21731), .Z(n22246) );
  NOR U22080 ( .A(n22247), .B(n22246), .Z(n21733) );
  NOR U22081 ( .A(n21734), .B(n21733), .Z(n21737) );
  NOR U22082 ( .A(n108), .B(n67), .Z(n21736) );
  IV U22083 ( .A(n21736), .Z(n21735) );
  NOR U22084 ( .A(n21737), .B(n21735), .Z(n21742) );
  XOR U22085 ( .A(n21737), .B(n21736), .Z(n22090) );
  XOR U22086 ( .A(n21739), .B(n21738), .Z(n22091) );
  IV U22087 ( .A(n22091), .Z(n21740) );
  NOR U22088 ( .A(n22090), .B(n21740), .Z(n21741) );
  NOR U22089 ( .A(n21742), .B(n21741), .Z(n22086) );
  XOR U22090 ( .A(n21744), .B(n21743), .Z(n22087) );
  NOR U22091 ( .A(n22086), .B(n22087), .Z(n21745) );
  NOR U22092 ( .A(n21746), .B(n21745), .Z(n22082) );
  XOR U22093 ( .A(n21748), .B(n21747), .Z(n22083) );
  NOR U22094 ( .A(n22082), .B(n22083), .Z(n21749) );
  NOR U22095 ( .A(n21750), .B(n21749), .Z(n22078) );
  XOR U22096 ( .A(n21752), .B(n21751), .Z(n22079) );
  NOR U22097 ( .A(n22078), .B(n22079), .Z(n21753) );
  NOR U22098 ( .A(n21754), .B(n21753), .Z(n22074) );
  XOR U22099 ( .A(n21756), .B(n21755), .Z(n22075) );
  NOR U22100 ( .A(n22074), .B(n22075), .Z(n21757) );
  NOR U22101 ( .A(n21758), .B(n21757), .Z(n22070) );
  XOR U22102 ( .A(n21760), .B(n21759), .Z(n22071) );
  NOR U22103 ( .A(n22070), .B(n22071), .Z(n21761) );
  NOR U22104 ( .A(n21762), .B(n21761), .Z(n22066) );
  XOR U22105 ( .A(n21764), .B(n21763), .Z(n22067) );
  NOR U22106 ( .A(n22066), .B(n22067), .Z(n21765) );
  NOR U22107 ( .A(n21766), .B(n21765), .Z(n22062) );
  XOR U22108 ( .A(n21768), .B(n21767), .Z(n22063) );
  NOR U22109 ( .A(n22062), .B(n22063), .Z(n21769) );
  NOR U22110 ( .A(n21770), .B(n21769), .Z(n22058) );
  XOR U22111 ( .A(n21772), .B(n21771), .Z(n22059) );
  NOR U22112 ( .A(n22058), .B(n22059), .Z(n21773) );
  NOR U22113 ( .A(n21774), .B(n21773), .Z(n21775) );
  IV U22114 ( .A(n21775), .Z(n22056) );
  XOR U22115 ( .A(n21777), .B(n21776), .Z(n21778) );
  IV U22116 ( .A(n21778), .Z(n22055) );
  NOR U22117 ( .A(n22056), .B(n22055), .Z(n21779) );
  NOR U22118 ( .A(n21780), .B(n21779), .Z(n21781) );
  IV U22119 ( .A(n21781), .Z(n22054) );
  XOR U22120 ( .A(n21783), .B(n21782), .Z(n22053) );
  NOR U22121 ( .A(n22054), .B(n22053), .Z(n21784) );
  NOR U22122 ( .A(n21785), .B(n21784), .Z(n21786) );
  IV U22123 ( .A(n21786), .Z(n22051) );
  XOR U22124 ( .A(n21788), .B(n21787), .Z(n21789) );
  IV U22125 ( .A(n21789), .Z(n22050) );
  NOR U22126 ( .A(n22051), .B(n22050), .Z(n21790) );
  NOR U22127 ( .A(n21791), .B(n21790), .Z(n21792) );
  IV U22128 ( .A(n21792), .Z(n22046) );
  XOR U22129 ( .A(n21794), .B(n21793), .Z(n22045) );
  NOR U22130 ( .A(n22046), .B(n22045), .Z(n21795) );
  NOR U22131 ( .A(n21796), .B(n21795), .Z(n21797) );
  IV U22132 ( .A(n21797), .Z(n22043) );
  XOR U22133 ( .A(n21799), .B(n21798), .Z(n21800) );
  IV U22134 ( .A(n21800), .Z(n22042) );
  NOR U22135 ( .A(n22043), .B(n22042), .Z(n21801) );
  NOR U22136 ( .A(n21802), .B(n21801), .Z(n21803) );
  IV U22137 ( .A(n21803), .Z(n22041) );
  XOR U22138 ( .A(n21805), .B(n21804), .Z(n22040) );
  NOR U22139 ( .A(n22041), .B(n22040), .Z(n21806) );
  NOR U22140 ( .A(n21807), .B(n21806), .Z(n21808) );
  IV U22141 ( .A(n21808), .Z(n22038) );
  XOR U22142 ( .A(n21810), .B(n21809), .Z(n21811) );
  IV U22143 ( .A(n21811), .Z(n22037) );
  NOR U22144 ( .A(n22038), .B(n22037), .Z(n21812) );
  NOR U22145 ( .A(n21813), .B(n21812), .Z(n21814) );
  IV U22146 ( .A(n21814), .Z(n22036) );
  XOR U22147 ( .A(n21816), .B(n21815), .Z(n22035) );
  NOR U22148 ( .A(n22036), .B(n22035), .Z(n21817) );
  NOR U22149 ( .A(n21818), .B(n21817), .Z(n21819) );
  IV U22150 ( .A(n21819), .Z(n22033) );
  XOR U22151 ( .A(n21821), .B(n21820), .Z(n21822) );
  IV U22152 ( .A(n21822), .Z(n22032) );
  NOR U22153 ( .A(n22033), .B(n22032), .Z(n21823) );
  NOR U22154 ( .A(n21824), .B(n21823), .Z(n21825) );
  IV U22155 ( .A(n21825), .Z(n22031) );
  XOR U22156 ( .A(n21827), .B(n21826), .Z(n22030) );
  NOR U22157 ( .A(n22031), .B(n22030), .Z(n21828) );
  NOR U22158 ( .A(n21829), .B(n21828), .Z(n21830) );
  IV U22159 ( .A(n21830), .Z(n22028) );
  XOR U22160 ( .A(n21832), .B(n21831), .Z(n21833) );
  IV U22161 ( .A(n21833), .Z(n22027) );
  NOR U22162 ( .A(n22028), .B(n22027), .Z(n21834) );
  NOR U22163 ( .A(n21835), .B(n21834), .Z(n21836) );
  IV U22164 ( .A(n21836), .Z(n22026) );
  XOR U22165 ( .A(n21838), .B(n21837), .Z(n22025) );
  NOR U22166 ( .A(n22026), .B(n22025), .Z(n21839) );
  NOR U22167 ( .A(n21840), .B(n21839), .Z(n21841) );
  IV U22168 ( .A(n21841), .Z(n22023) );
  XOR U22169 ( .A(n21843), .B(n21842), .Z(n21844) );
  IV U22170 ( .A(n21844), .Z(n22022) );
  NOR U22171 ( .A(n22023), .B(n22022), .Z(n21845) );
  NOR U22172 ( .A(n21846), .B(n21845), .Z(n21847) );
  IV U22173 ( .A(n21847), .Z(n22021) );
  XOR U22174 ( .A(n21849), .B(n21848), .Z(n22020) );
  NOR U22175 ( .A(n22021), .B(n22020), .Z(n21850) );
  NOR U22176 ( .A(n21851), .B(n21850), .Z(n21852) );
  IV U22177 ( .A(n21852), .Z(n22018) );
  XOR U22178 ( .A(n21854), .B(n21853), .Z(n21855) );
  IV U22179 ( .A(n21855), .Z(n22017) );
  NOR U22180 ( .A(n22018), .B(n22017), .Z(n21856) );
  NOR U22181 ( .A(n21857), .B(n21856), .Z(n21858) );
  IV U22182 ( .A(n21858), .Z(n22013) );
  XOR U22183 ( .A(n21860), .B(n21859), .Z(n22012) );
  NOR U22184 ( .A(n22013), .B(n22012), .Z(n21861) );
  NOR U22185 ( .A(n21862), .B(n21861), .Z(n21863) );
  IV U22186 ( .A(n21863), .Z(n22010) );
  XOR U22187 ( .A(n21865), .B(n21864), .Z(n21866) );
  IV U22188 ( .A(n21866), .Z(n22009) );
  NOR U22189 ( .A(n22010), .B(n22009), .Z(n21867) );
  NOR U22190 ( .A(n21868), .B(n21867), .Z(n22007) );
  IV U22191 ( .A(n22007), .Z(n21869) );
  NOR U22192 ( .A(n22006), .B(n21869), .Z(n21870) );
  NOR U22193 ( .A(n21871), .B(n21870), .Z(n21872) );
  IV U22194 ( .A(n21872), .Z(n22004) );
  XOR U22195 ( .A(n21874), .B(n21873), .Z(n21875) );
  IV U22196 ( .A(n21875), .Z(n22003) );
  NOR U22197 ( .A(n22004), .B(n22003), .Z(n21876) );
  NOR U22198 ( .A(n21877), .B(n21876), .Z(n22001) );
  IV U22199 ( .A(n22001), .Z(n21878) );
  NOR U22200 ( .A(n22000), .B(n21878), .Z(n21879) );
  NOR U22201 ( .A(n21880), .B(n21879), .Z(n21881) );
  IV U22202 ( .A(n21881), .Z(n21998) );
  XOR U22203 ( .A(n21883), .B(n21882), .Z(n21884) );
  IV U22204 ( .A(n21884), .Z(n21997) );
  NOR U22205 ( .A(n21998), .B(n21997), .Z(n21885) );
  NOR U22206 ( .A(n21886), .B(n21885), .Z(n21887) );
  IV U22207 ( .A(n21887), .Z(n21892) );
  NOR U22208 ( .A(n143), .B(n67), .Z(n21891) );
  IV U22209 ( .A(n21891), .Z(n21888) );
  NOR U22210 ( .A(n21892), .B(n21888), .Z(n21895) );
  XOR U22211 ( .A(n21890), .B(n21889), .Z(n22395) );
  IV U22212 ( .A(n22395), .Z(n21893) );
  XOR U22213 ( .A(n21892), .B(n21891), .Z(n22396) );
  NOR U22214 ( .A(n21893), .B(n22396), .Z(n21894) );
  NOR U22215 ( .A(n21895), .B(n21894), .Z(n21900) );
  NOR U22216 ( .A(n145), .B(n67), .Z(n21899) );
  IV U22217 ( .A(n21899), .Z(n21896) );
  NOR U22218 ( .A(n21900), .B(n21896), .Z(n21902) );
  XOR U22219 ( .A(n21898), .B(n21897), .Z(n22401) );
  XOR U22220 ( .A(n21900), .B(n21899), .Z(n22400) );
  NOR U22221 ( .A(n22401), .B(n22400), .Z(n21901) );
  NOR U22222 ( .A(n21902), .B(n21901), .Z(n21905) );
  NOR U22223 ( .A(n147), .B(n67), .Z(n21904) );
  IV U22224 ( .A(n21904), .Z(n21903) );
  NOR U22225 ( .A(n21905), .B(n21903), .Z(n21910) );
  XOR U22226 ( .A(n21905), .B(n21904), .Z(n21994) );
  XOR U22227 ( .A(n21907), .B(n21906), .Z(n21995) );
  IV U22228 ( .A(n21995), .Z(n21908) );
  NOR U22229 ( .A(n21994), .B(n21908), .Z(n21909) );
  NOR U22230 ( .A(n21910), .B(n21909), .Z(n21915) );
  XOR U22231 ( .A(n21912), .B(n21911), .Z(n21914) );
  IV U22232 ( .A(n21914), .Z(n21913) );
  NOR U22233 ( .A(n21915), .B(n21913), .Z(n21918) );
  XOR U22234 ( .A(n21915), .B(n21914), .Z(n22415) );
  NOR U22235 ( .A(n148), .B(n67), .Z(n22416) );
  IV U22236 ( .A(n22416), .Z(n21916) );
  NOR U22237 ( .A(n22415), .B(n21916), .Z(n21917) );
  NOR U22238 ( .A(n21918), .B(n21917), .Z(n21921) );
  NOR U22239 ( .A(n150), .B(n67), .Z(n21920) );
  IV U22240 ( .A(n21920), .Z(n21919) );
  NOR U22241 ( .A(n21921), .B(n21919), .Z(n21925) );
  XOR U22242 ( .A(n21921), .B(n21920), .Z(n22420) );
  XOR U22243 ( .A(n21923), .B(n21922), .Z(n22421) );
  NOR U22244 ( .A(n22420), .B(n22421), .Z(n21924) );
  NOR U22245 ( .A(n21925), .B(n21924), .Z(n21930) );
  NOR U22246 ( .A(n153), .B(n67), .Z(n21929) );
  IV U22247 ( .A(n21929), .Z(n21926) );
  NOR U22248 ( .A(n21930), .B(n21926), .Z(n21932) );
  XOR U22249 ( .A(n21928), .B(n21927), .Z(n22429) );
  XOR U22250 ( .A(n21930), .B(n21929), .Z(n22428) );
  NOR U22251 ( .A(n22429), .B(n22428), .Z(n21931) );
  NOR U22252 ( .A(n21932), .B(n21931), .Z(n21934) );
  IV U22253 ( .A(n21934), .Z(n21933) );
  NOR U22254 ( .A(n21935), .B(n21933), .Z(n21937) );
  NOR U22255 ( .A(n155), .B(n67), .Z(n22437) );
  XOR U22256 ( .A(n21935), .B(n21934), .Z(n22436) );
  NOR U22257 ( .A(n22437), .B(n22436), .Z(n21936) );
  NOR U22258 ( .A(n21937), .B(n21936), .Z(n21939) );
  NOR U22259 ( .A(n21938), .B(n21939), .Z(n21944) );
  IV U22260 ( .A(n21938), .Z(n22444) );
  IV U22261 ( .A(n21939), .Z(n22443) );
  NOR U22262 ( .A(n22444), .B(n22443), .Z(n21942) );
  XOR U22263 ( .A(n21941), .B(n21940), .Z(n22446) );
  NOR U22264 ( .A(n21942), .B(n22446), .Z(n21943) );
  NOR U22265 ( .A(n21944), .B(n21943), .Z(n21952) );
  IV U22266 ( .A(n21952), .Z(n21946) );
  NOR U22267 ( .A(n158), .B(n67), .Z(n21945) );
  IV U22268 ( .A(n21945), .Z(n21951) );
  NOR U22269 ( .A(n21946), .B(n21951), .Z(n21954) );
  XOR U22270 ( .A(n21948), .B(n21947), .Z(n21949) );
  XOR U22271 ( .A(n21950), .B(n21949), .Z(n22452) );
  XOR U22272 ( .A(n21952), .B(n21951), .Z(n22453) );
  NOR U22273 ( .A(n22452), .B(n22453), .Z(n21953) );
  NOR U22274 ( .A(n21954), .B(n21953), .Z(n21959) );
  XOR U22275 ( .A(n21956), .B(n21955), .Z(n21958) );
  IV U22276 ( .A(n21958), .Z(n21957) );
  NOR U22277 ( .A(n21959), .B(n21957), .Z(n21962) );
  XOR U22278 ( .A(n21959), .B(n21958), .Z(n22463) );
  NOR U22279 ( .A(n161), .B(n67), .Z(n22464) );
  IV U22280 ( .A(n22464), .Z(n21960) );
  NOR U22281 ( .A(n22463), .B(n21960), .Z(n21961) );
  NOR U22282 ( .A(n21962), .B(n21961), .Z(n21965) );
  NOR U22283 ( .A(n163), .B(n67), .Z(n21964) );
  IV U22284 ( .A(n21964), .Z(n21963) );
  NOR U22285 ( .A(n21965), .B(n21963), .Z(n21969) );
  XOR U22286 ( .A(n21965), .B(n21964), .Z(n22470) );
  XOR U22287 ( .A(n21967), .B(n21966), .Z(n22471) );
  NOR U22288 ( .A(n22470), .B(n22471), .Z(n21968) );
  NOR U22289 ( .A(n21969), .B(n21968), .Z(n21976) );
  NOR U22290 ( .A(n165), .B(n67), .Z(n21975) );
  IV U22291 ( .A(n21975), .Z(n21970) );
  NOR U22292 ( .A(n21976), .B(n21970), .Z(n21978) );
  XOR U22293 ( .A(n21972), .B(n21971), .Z(n21973) );
  XOR U22294 ( .A(n21974), .B(n21973), .Z(n22476) );
  XOR U22295 ( .A(n21976), .B(n21975), .Z(n22475) );
  NOR U22296 ( .A(n22476), .B(n22475), .Z(n21977) );
  NOR U22297 ( .A(n21978), .B(n21977), .Z(n21983) );
  XOR U22298 ( .A(n21980), .B(n21979), .Z(n21982) );
  IV U22299 ( .A(n21982), .Z(n21981) );
  NOR U22300 ( .A(n21983), .B(n21981), .Z(n21986) );
  XOR U22301 ( .A(n21983), .B(n21982), .Z(n22483) );
  NOR U22302 ( .A(n167), .B(n67), .Z(n22484) );
  IV U22303 ( .A(n22484), .Z(n21984) );
  NOR U22304 ( .A(n22483), .B(n21984), .Z(n21985) );
  NOR U22305 ( .A(n21986), .B(n21985), .Z(n22486) );
  XOR U22306 ( .A(n21988), .B(n21987), .Z(n22485) );
  NOR U22307 ( .A(n22486), .B(n22485), .Z(n21992) );
  XOR U22308 ( .A(n21990), .B(n21989), .Z(n21991) );
  NOR U22309 ( .A(n21992), .B(n21991), .Z(n28538) );
  XOR U22310 ( .A(n21992), .B(n21991), .Z(n21993) );
  IV U22311 ( .A(n21993), .Z(n31542) );
  NOR U22312 ( .A(n155), .B(n68), .Z(n22431) );
  XOR U22313 ( .A(n21995), .B(n21994), .Z(n22408) );
  NOR U22314 ( .A(n148), .B(n68), .Z(n22409) );
  IV U22315 ( .A(n22409), .Z(n21996) );
  NOR U22316 ( .A(n22408), .B(n21996), .Z(n22411) );
  XOR U22317 ( .A(n21998), .B(n21997), .Z(n22389) );
  NOR U22318 ( .A(n143), .B(n68), .Z(n22388) );
  IV U22319 ( .A(n22388), .Z(n21999) );
  NOR U22320 ( .A(n22389), .B(n21999), .Z(n22391) );
  NOR U22321 ( .A(n141), .B(n68), .Z(n22385) );
  IV U22322 ( .A(n22385), .Z(n22002) );
  XOR U22323 ( .A(n22001), .B(n22000), .Z(n22384) );
  NOR U22324 ( .A(n22002), .B(n22384), .Z(n22387) );
  XOR U22325 ( .A(n22004), .B(n22003), .Z(n22381) );
  NOR U22326 ( .A(n139), .B(n68), .Z(n22380) );
  IV U22327 ( .A(n22380), .Z(n22005) );
  NOR U22328 ( .A(n22381), .B(n22005), .Z(n22383) );
  NOR U22329 ( .A(n137), .B(n68), .Z(n22377) );
  IV U22330 ( .A(n22377), .Z(n22008) );
  XOR U22331 ( .A(n22007), .B(n22006), .Z(n22376) );
  NOR U22332 ( .A(n22008), .B(n22376), .Z(n22379) );
  XOR U22333 ( .A(n22010), .B(n22009), .Z(n22373) );
  NOR U22334 ( .A(n135), .B(n68), .Z(n22372) );
  IV U22335 ( .A(n22372), .Z(n22011) );
  NOR U22336 ( .A(n22373), .B(n22011), .Z(n22375) );
  NOR U22337 ( .A(n133), .B(n68), .Z(n22015) );
  XOR U22338 ( .A(n22013), .B(n22012), .Z(n22014) );
  NOR U22339 ( .A(n22015), .B(n22014), .Z(n22370) );
  XOR U22340 ( .A(n22015), .B(n22014), .Z(n22016) );
  IV U22341 ( .A(n22016), .Z(n22523) );
  XOR U22342 ( .A(n22018), .B(n22017), .Z(n22365) );
  NOR U22343 ( .A(n131), .B(n68), .Z(n22364) );
  IV U22344 ( .A(n22364), .Z(n22019) );
  NOR U22345 ( .A(n22365), .B(n22019), .Z(n22367) );
  NOR U22346 ( .A(n128), .B(n68), .Z(n22359) );
  XOR U22347 ( .A(n22021), .B(n22020), .Z(n22358) );
  NOR U22348 ( .A(n22359), .B(n22358), .Z(n22362) );
  XOR U22349 ( .A(n22023), .B(n22022), .Z(n22354) );
  NOR U22350 ( .A(n126), .B(n68), .Z(n22353) );
  IV U22351 ( .A(n22353), .Z(n22024) );
  NOR U22352 ( .A(n22354), .B(n22024), .Z(n22356) );
  NOR U22353 ( .A(n125), .B(n68), .Z(n22348) );
  XOR U22354 ( .A(n22026), .B(n22025), .Z(n22347) );
  NOR U22355 ( .A(n22348), .B(n22347), .Z(n22351) );
  XOR U22356 ( .A(n22028), .B(n22027), .Z(n22343) );
  NOR U22357 ( .A(n123), .B(n68), .Z(n22342) );
  IV U22358 ( .A(n22342), .Z(n22029) );
  NOR U22359 ( .A(n22343), .B(n22029), .Z(n22345) );
  NOR U22360 ( .A(n120), .B(n68), .Z(n22337) );
  XOR U22361 ( .A(n22031), .B(n22030), .Z(n22336) );
  NOR U22362 ( .A(n22337), .B(n22336), .Z(n22340) );
  XOR U22363 ( .A(n22033), .B(n22032), .Z(n22332) );
  NOR U22364 ( .A(n119), .B(n68), .Z(n22331) );
  IV U22365 ( .A(n22331), .Z(n22034) );
  NOR U22366 ( .A(n22332), .B(n22034), .Z(n22334) );
  NOR U22367 ( .A(n79), .B(n68), .Z(n22326) );
  XOR U22368 ( .A(n22036), .B(n22035), .Z(n22325) );
  NOR U22369 ( .A(n22326), .B(n22325), .Z(n22329) );
  XOR U22370 ( .A(n22038), .B(n22037), .Z(n22321) );
  NOR U22371 ( .A(n117), .B(n68), .Z(n22320) );
  IV U22372 ( .A(n22320), .Z(n22039) );
  NOR U22373 ( .A(n22321), .B(n22039), .Z(n22323) );
  NOR U22374 ( .A(n80), .B(n68), .Z(n22315) );
  XOR U22375 ( .A(n22041), .B(n22040), .Z(n22314) );
  NOR U22376 ( .A(n22315), .B(n22314), .Z(n22318) );
  XOR U22377 ( .A(n22043), .B(n22042), .Z(n22310) );
  NOR U22378 ( .A(n116), .B(n68), .Z(n22309) );
  IV U22379 ( .A(n22309), .Z(n22044) );
  NOR U22380 ( .A(n22310), .B(n22044), .Z(n22312) );
  NOR U22381 ( .A(n81), .B(n68), .Z(n22048) );
  XOR U22382 ( .A(n22046), .B(n22045), .Z(n22047) );
  NOR U22383 ( .A(n22048), .B(n22047), .Z(n22307) );
  XOR U22384 ( .A(n22048), .B(n22047), .Z(n22049) );
  IV U22385 ( .A(n22049), .Z(n22554) );
  XOR U22386 ( .A(n22051), .B(n22050), .Z(n22302) );
  NOR U22387 ( .A(n115), .B(n68), .Z(n22301) );
  IV U22388 ( .A(n22301), .Z(n22052) );
  NOR U22389 ( .A(n22302), .B(n22052), .Z(n22304) );
  NOR U22390 ( .A(n82), .B(n68), .Z(n22296) );
  XOR U22391 ( .A(n22054), .B(n22053), .Z(n22295) );
  NOR U22392 ( .A(n22296), .B(n22295), .Z(n22299) );
  XOR U22393 ( .A(n22056), .B(n22055), .Z(n22291) );
  NOR U22394 ( .A(n114), .B(n68), .Z(n22290) );
  IV U22395 ( .A(n22290), .Z(n22057) );
  NOR U22396 ( .A(n22291), .B(n22057), .Z(n22293) );
  IV U22397 ( .A(n22058), .Z(n22060) );
  XOR U22398 ( .A(n22060), .B(n22059), .Z(n22286) );
  NOR U22399 ( .A(n83), .B(n68), .Z(n22287) );
  IV U22400 ( .A(n22287), .Z(n22061) );
  NOR U22401 ( .A(n22286), .B(n22061), .Z(n22289) );
  IV U22402 ( .A(n22062), .Z(n22064) );
  XOR U22403 ( .A(n22064), .B(n22063), .Z(n22282) );
  NOR U22404 ( .A(n113), .B(n68), .Z(n22283) );
  IV U22405 ( .A(n22283), .Z(n22065) );
  NOR U22406 ( .A(n22282), .B(n22065), .Z(n22285) );
  IV U22407 ( .A(n22066), .Z(n22068) );
  XOR U22408 ( .A(n22068), .B(n22067), .Z(n22278) );
  NOR U22409 ( .A(n84), .B(n68), .Z(n22279) );
  IV U22410 ( .A(n22279), .Z(n22069) );
  NOR U22411 ( .A(n22278), .B(n22069), .Z(n22281) );
  IV U22412 ( .A(n22070), .Z(n22072) );
  XOR U22413 ( .A(n22072), .B(n22071), .Z(n22274) );
  NOR U22414 ( .A(n112), .B(n68), .Z(n22275) );
  IV U22415 ( .A(n22275), .Z(n22073) );
  NOR U22416 ( .A(n22274), .B(n22073), .Z(n22277) );
  IV U22417 ( .A(n22074), .Z(n22076) );
  XOR U22418 ( .A(n22076), .B(n22075), .Z(n22270) );
  NOR U22419 ( .A(n85), .B(n68), .Z(n22271) );
  IV U22420 ( .A(n22271), .Z(n22077) );
  NOR U22421 ( .A(n22270), .B(n22077), .Z(n22273) );
  IV U22422 ( .A(n22078), .Z(n22080) );
  XOR U22423 ( .A(n22080), .B(n22079), .Z(n22266) );
  NOR U22424 ( .A(n111), .B(n68), .Z(n22267) );
  IV U22425 ( .A(n22267), .Z(n22081) );
  NOR U22426 ( .A(n22266), .B(n22081), .Z(n22269) );
  IV U22427 ( .A(n22082), .Z(n22084) );
  XOR U22428 ( .A(n22084), .B(n22083), .Z(n22262) );
  NOR U22429 ( .A(n86), .B(n68), .Z(n22263) );
  IV U22430 ( .A(n22263), .Z(n22085) );
  NOR U22431 ( .A(n22262), .B(n22085), .Z(n22265) );
  IV U22432 ( .A(n22086), .Z(n22088) );
  XOR U22433 ( .A(n22088), .B(n22087), .Z(n22258) );
  NOR U22434 ( .A(n110), .B(n68), .Z(n22259) );
  IV U22435 ( .A(n22259), .Z(n22089) );
  NOR U22436 ( .A(n22258), .B(n22089), .Z(n22261) );
  XOR U22437 ( .A(n22091), .B(n22090), .Z(n22254) );
  NOR U22438 ( .A(n109), .B(n68), .Z(n22255) );
  IV U22439 ( .A(n22255), .Z(n22092) );
  NOR U22440 ( .A(n22254), .B(n22092), .Z(n22257) );
  XOR U22441 ( .A(n22094), .B(n22093), .Z(n22242) );
  IV U22442 ( .A(n22242), .Z(n22096) );
  NOR U22443 ( .A(n87), .B(n68), .Z(n22095) );
  IV U22444 ( .A(n22095), .Z(n22243) );
  NOR U22445 ( .A(n22096), .B(n22243), .Z(n22245) );
  IV U22446 ( .A(n22097), .Z(n22099) );
  XOR U22447 ( .A(n22099), .B(n22098), .Z(n22238) );
  NOR U22448 ( .A(n107), .B(n68), .Z(n22239) );
  IV U22449 ( .A(n22239), .Z(n22100) );
  NOR U22450 ( .A(n22238), .B(n22100), .Z(n22241) );
  IV U22451 ( .A(n22101), .Z(n22103) );
  XOR U22452 ( .A(n22103), .B(n22102), .Z(n22234) );
  NOR U22453 ( .A(n88), .B(n68), .Z(n22235) );
  IV U22454 ( .A(n22235), .Z(n22104) );
  NOR U22455 ( .A(n22234), .B(n22104), .Z(n22237) );
  IV U22456 ( .A(n22105), .Z(n22107) );
  XOR U22457 ( .A(n22107), .B(n22106), .Z(n22230) );
  NOR U22458 ( .A(n106), .B(n68), .Z(n22231) );
  IV U22459 ( .A(n22231), .Z(n22108) );
  NOR U22460 ( .A(n22230), .B(n22108), .Z(n22233) );
  XOR U22461 ( .A(n22110), .B(n22109), .Z(n22226) );
  NOR U22462 ( .A(n105), .B(n68), .Z(n22227) );
  IV U22463 ( .A(n22227), .Z(n22111) );
  NOR U22464 ( .A(n22226), .B(n22111), .Z(n22229) );
  XOR U22465 ( .A(n22113), .B(n22112), .Z(n22214) );
  IV U22466 ( .A(n22214), .Z(n22115) );
  NOR U22467 ( .A(n89), .B(n68), .Z(n22114) );
  IV U22468 ( .A(n22114), .Z(n22215) );
  NOR U22469 ( .A(n22115), .B(n22215), .Z(n22217) );
  IV U22470 ( .A(n22116), .Z(n22118) );
  XOR U22471 ( .A(n22118), .B(n22117), .Z(n22210) );
  NOR U22472 ( .A(n103), .B(n68), .Z(n22211) );
  IV U22473 ( .A(n22211), .Z(n22119) );
  NOR U22474 ( .A(n22210), .B(n22119), .Z(n22213) );
  IV U22475 ( .A(n22120), .Z(n22122) );
  XOR U22476 ( .A(n22122), .B(n22121), .Z(n22206) );
  NOR U22477 ( .A(n90), .B(n68), .Z(n22207) );
  IV U22478 ( .A(n22207), .Z(n22123) );
  NOR U22479 ( .A(n22206), .B(n22123), .Z(n22209) );
  IV U22480 ( .A(n22124), .Z(n22126) );
  XOR U22481 ( .A(n22126), .B(n22125), .Z(n22202) );
  NOR U22482 ( .A(n102), .B(n68), .Z(n22203) );
  IV U22483 ( .A(n22203), .Z(n22127) );
  NOR U22484 ( .A(n22202), .B(n22127), .Z(n22205) );
  IV U22485 ( .A(n22128), .Z(n22130) );
  XOR U22486 ( .A(n22130), .B(n22129), .Z(n22198) );
  NOR U22487 ( .A(n101), .B(n68), .Z(n22199) );
  IV U22488 ( .A(n22199), .Z(n22131) );
  NOR U22489 ( .A(n22198), .B(n22131), .Z(n22201) );
  IV U22490 ( .A(n22132), .Z(n22134) );
  XOR U22491 ( .A(n22134), .B(n22133), .Z(n22194) );
  NOR U22492 ( .A(n100), .B(n68), .Z(n22195) );
  IV U22493 ( .A(n22195), .Z(n22135) );
  NOR U22494 ( .A(n22194), .B(n22135), .Z(n22197) );
  IV U22495 ( .A(n22136), .Z(n22138) );
  XOR U22496 ( .A(n22138), .B(n22137), .Z(n22190) );
  NOR U22497 ( .A(n99), .B(n68), .Z(n22191) );
  IV U22498 ( .A(n22191), .Z(n22139) );
  NOR U22499 ( .A(n22190), .B(n22139), .Z(n22193) );
  IV U22500 ( .A(n22140), .Z(n22142) );
  XOR U22501 ( .A(n22142), .B(n22141), .Z(n22186) );
  NOR U22502 ( .A(n98), .B(n68), .Z(n22187) );
  IV U22503 ( .A(n22187), .Z(n22143) );
  NOR U22504 ( .A(n22186), .B(n22143), .Z(n22189) );
  XOR U22505 ( .A(n22145), .B(n22144), .Z(n22182) );
  NOR U22506 ( .A(n91), .B(n68), .Z(n22183) );
  IV U22507 ( .A(n22183), .Z(n22146) );
  NOR U22508 ( .A(n22182), .B(n22146), .Z(n22185) );
  XOR U22509 ( .A(n22148), .B(n22147), .Z(n22170) );
  IV U22510 ( .A(n22170), .Z(n22150) );
  NOR U22511 ( .A(n96), .B(n68), .Z(n22149) );
  IV U22512 ( .A(n22149), .Z(n22171) );
  NOR U22513 ( .A(n22150), .B(n22171), .Z(n22173) );
  NOR U22514 ( .A(n95), .B(n68), .Z(n22167) );
  IV U22515 ( .A(n22167), .Z(n22153) );
  XOR U22516 ( .A(n22152), .B(n22151), .Z(n22166) );
  NOR U22517 ( .A(n22153), .B(n22166), .Z(n22169) );
  NOR U22518 ( .A(n68), .B(n93), .Z(n23170) );
  IV U22519 ( .A(n23170), .Z(n22154) );
  NOR U22520 ( .A(n67), .B(n168), .Z(n22162) );
  IV U22521 ( .A(n22162), .Z(n22157) );
  NOR U22522 ( .A(n22154), .B(n22157), .Z(n22155) );
  IV U22523 ( .A(n22155), .Z(n22156) );
  NOR U22524 ( .A(n94), .B(n22156), .Z(n22165) );
  NOR U22525 ( .A(n22157), .B(n93), .Z(n22158) );
  XOR U22526 ( .A(n94), .B(n22158), .Z(n22159) );
  NOR U22527 ( .A(n68), .B(n22159), .Z(n22160) );
  IV U22528 ( .A(n22160), .Z(n22661) );
  XOR U22529 ( .A(n22162), .B(n22161), .Z(n22660) );
  IV U22530 ( .A(n22660), .Z(n22163) );
  NOR U22531 ( .A(n22661), .B(n22163), .Z(n22164) );
  NOR U22532 ( .A(n22165), .B(n22164), .Z(n22657) );
  XOR U22533 ( .A(n22167), .B(n22166), .Z(n22656) );
  NOR U22534 ( .A(n22657), .B(n22656), .Z(n22168) );
  NOR U22535 ( .A(n22169), .B(n22168), .Z(n22684) );
  XOR U22536 ( .A(n22171), .B(n22170), .Z(n22683) );
  NOR U22537 ( .A(n22684), .B(n22683), .Z(n22172) );
  NOR U22538 ( .A(n22173), .B(n22172), .Z(n22178) );
  XOR U22539 ( .A(n22175), .B(n22174), .Z(n22177) );
  IV U22540 ( .A(n22177), .Z(n22176) );
  NOR U22541 ( .A(n22178), .B(n22176), .Z(n22181) );
  XOR U22542 ( .A(n22178), .B(n22177), .Z(n22653) );
  NOR U22543 ( .A(n97), .B(n68), .Z(n22654) );
  IV U22544 ( .A(n22654), .Z(n22179) );
  NOR U22545 ( .A(n22653), .B(n22179), .Z(n22180) );
  NOR U22546 ( .A(n22181), .B(n22180), .Z(n22649) );
  XOR U22547 ( .A(n22183), .B(n22182), .Z(n22650) );
  NOR U22548 ( .A(n22649), .B(n22650), .Z(n22184) );
  NOR U22549 ( .A(n22185), .B(n22184), .Z(n22645) );
  XOR U22550 ( .A(n22187), .B(n22186), .Z(n22646) );
  NOR U22551 ( .A(n22645), .B(n22646), .Z(n22188) );
  NOR U22552 ( .A(n22189), .B(n22188), .Z(n22641) );
  XOR U22553 ( .A(n22191), .B(n22190), .Z(n22642) );
  NOR U22554 ( .A(n22641), .B(n22642), .Z(n22192) );
  NOR U22555 ( .A(n22193), .B(n22192), .Z(n22637) );
  XOR U22556 ( .A(n22195), .B(n22194), .Z(n22638) );
  NOR U22557 ( .A(n22637), .B(n22638), .Z(n22196) );
  NOR U22558 ( .A(n22197), .B(n22196), .Z(n22633) );
  XOR U22559 ( .A(n22199), .B(n22198), .Z(n22634) );
  NOR U22560 ( .A(n22633), .B(n22634), .Z(n22200) );
  NOR U22561 ( .A(n22201), .B(n22200), .Z(n22629) );
  XOR U22562 ( .A(n22203), .B(n22202), .Z(n22630) );
  NOR U22563 ( .A(n22629), .B(n22630), .Z(n22204) );
  NOR U22564 ( .A(n22205), .B(n22204), .Z(n22625) );
  XOR U22565 ( .A(n22207), .B(n22206), .Z(n22626) );
  NOR U22566 ( .A(n22625), .B(n22626), .Z(n22208) );
  NOR U22567 ( .A(n22209), .B(n22208), .Z(n22622) );
  XOR U22568 ( .A(n22211), .B(n22210), .Z(n22621) );
  NOR U22569 ( .A(n22622), .B(n22621), .Z(n22212) );
  NOR U22570 ( .A(n22213), .B(n22212), .Z(n22728) );
  XOR U22571 ( .A(n22215), .B(n22214), .Z(n22727) );
  NOR U22572 ( .A(n22728), .B(n22727), .Z(n22216) );
  NOR U22573 ( .A(n22217), .B(n22216), .Z(n22222) );
  XOR U22574 ( .A(n22219), .B(n22218), .Z(n22221) );
  IV U22575 ( .A(n22221), .Z(n22220) );
  NOR U22576 ( .A(n22222), .B(n22220), .Z(n22225) );
  XOR U22577 ( .A(n22222), .B(n22221), .Z(n22618) );
  NOR U22578 ( .A(n104), .B(n68), .Z(n22619) );
  IV U22579 ( .A(n22619), .Z(n22223) );
  NOR U22580 ( .A(n22618), .B(n22223), .Z(n22224) );
  NOR U22581 ( .A(n22225), .B(n22224), .Z(n22614) );
  XOR U22582 ( .A(n22227), .B(n22226), .Z(n22615) );
  NOR U22583 ( .A(n22614), .B(n22615), .Z(n22228) );
  NOR U22584 ( .A(n22229), .B(n22228), .Z(n22610) );
  XOR U22585 ( .A(n22231), .B(n22230), .Z(n22611) );
  NOR U22586 ( .A(n22610), .B(n22611), .Z(n22232) );
  NOR U22587 ( .A(n22233), .B(n22232), .Z(n22606) );
  XOR U22588 ( .A(n22235), .B(n22234), .Z(n22607) );
  NOR U22589 ( .A(n22606), .B(n22607), .Z(n22236) );
  NOR U22590 ( .A(n22237), .B(n22236), .Z(n22602) );
  XOR U22591 ( .A(n22239), .B(n22238), .Z(n22603) );
  NOR U22592 ( .A(n22602), .B(n22603), .Z(n22240) );
  NOR U22593 ( .A(n22241), .B(n22240), .Z(n22759) );
  XOR U22594 ( .A(n22243), .B(n22242), .Z(n22758) );
  NOR U22595 ( .A(n22759), .B(n22758), .Z(n22244) );
  NOR U22596 ( .A(n22245), .B(n22244), .Z(n22250) );
  XOR U22597 ( .A(n22247), .B(n22246), .Z(n22249) );
  IV U22598 ( .A(n22249), .Z(n22248) );
  NOR U22599 ( .A(n22250), .B(n22248), .Z(n22253) );
  XOR U22600 ( .A(n22250), .B(n22249), .Z(n22599) );
  NOR U22601 ( .A(n108), .B(n68), .Z(n22600) );
  IV U22602 ( .A(n22600), .Z(n22251) );
  NOR U22603 ( .A(n22599), .B(n22251), .Z(n22252) );
  NOR U22604 ( .A(n22253), .B(n22252), .Z(n22595) );
  XOR U22605 ( .A(n22255), .B(n22254), .Z(n22596) );
  NOR U22606 ( .A(n22595), .B(n22596), .Z(n22256) );
  NOR U22607 ( .A(n22257), .B(n22256), .Z(n22591) );
  XOR U22608 ( .A(n22259), .B(n22258), .Z(n22592) );
  NOR U22609 ( .A(n22591), .B(n22592), .Z(n22260) );
  NOR U22610 ( .A(n22261), .B(n22260), .Z(n22587) );
  XOR U22611 ( .A(n22263), .B(n22262), .Z(n22588) );
  NOR U22612 ( .A(n22587), .B(n22588), .Z(n22264) );
  NOR U22613 ( .A(n22265), .B(n22264), .Z(n22583) );
  XOR U22614 ( .A(n22267), .B(n22266), .Z(n22584) );
  NOR U22615 ( .A(n22583), .B(n22584), .Z(n22268) );
  NOR U22616 ( .A(n22269), .B(n22268), .Z(n22579) );
  XOR U22617 ( .A(n22271), .B(n22270), .Z(n22580) );
  NOR U22618 ( .A(n22579), .B(n22580), .Z(n22272) );
  NOR U22619 ( .A(n22273), .B(n22272), .Z(n22575) );
  XOR U22620 ( .A(n22275), .B(n22274), .Z(n22576) );
  NOR U22621 ( .A(n22575), .B(n22576), .Z(n22276) );
  NOR U22622 ( .A(n22277), .B(n22276), .Z(n22571) );
  XOR U22623 ( .A(n22279), .B(n22278), .Z(n22572) );
  NOR U22624 ( .A(n22571), .B(n22572), .Z(n22280) );
  NOR U22625 ( .A(n22281), .B(n22280), .Z(n22567) );
  XOR U22626 ( .A(n22283), .B(n22282), .Z(n22568) );
  NOR U22627 ( .A(n22567), .B(n22568), .Z(n22284) );
  NOR U22628 ( .A(n22285), .B(n22284), .Z(n22563) );
  XOR U22629 ( .A(n22287), .B(n22286), .Z(n22564) );
  NOR U22630 ( .A(n22563), .B(n22564), .Z(n22288) );
  NOR U22631 ( .A(n22289), .B(n22288), .Z(n22562) );
  XOR U22632 ( .A(n22291), .B(n22290), .Z(n22561) );
  NOR U22633 ( .A(n22562), .B(n22561), .Z(n22292) );
  NOR U22634 ( .A(n22293), .B(n22292), .Z(n22294) );
  IV U22635 ( .A(n22294), .Z(n22559) );
  XOR U22636 ( .A(n22296), .B(n22295), .Z(n22297) );
  IV U22637 ( .A(n22297), .Z(n22558) );
  NOR U22638 ( .A(n22559), .B(n22558), .Z(n22298) );
  NOR U22639 ( .A(n22299), .B(n22298), .Z(n22300) );
  IV U22640 ( .A(n22300), .Z(n22557) );
  XOR U22641 ( .A(n22302), .B(n22301), .Z(n22556) );
  NOR U22642 ( .A(n22557), .B(n22556), .Z(n22303) );
  NOR U22643 ( .A(n22304), .B(n22303), .Z(n22305) );
  IV U22644 ( .A(n22305), .Z(n22553) );
  NOR U22645 ( .A(n22554), .B(n22553), .Z(n22306) );
  NOR U22646 ( .A(n22307), .B(n22306), .Z(n22308) );
  IV U22647 ( .A(n22308), .Z(n22552) );
  XOR U22648 ( .A(n22310), .B(n22309), .Z(n22551) );
  NOR U22649 ( .A(n22552), .B(n22551), .Z(n22311) );
  NOR U22650 ( .A(n22312), .B(n22311), .Z(n22313) );
  IV U22651 ( .A(n22313), .Z(n22549) );
  XOR U22652 ( .A(n22315), .B(n22314), .Z(n22316) );
  IV U22653 ( .A(n22316), .Z(n22548) );
  NOR U22654 ( .A(n22549), .B(n22548), .Z(n22317) );
  NOR U22655 ( .A(n22318), .B(n22317), .Z(n22319) );
  IV U22656 ( .A(n22319), .Z(n22547) );
  XOR U22657 ( .A(n22321), .B(n22320), .Z(n22546) );
  NOR U22658 ( .A(n22547), .B(n22546), .Z(n22322) );
  NOR U22659 ( .A(n22323), .B(n22322), .Z(n22324) );
  IV U22660 ( .A(n22324), .Z(n22544) );
  XOR U22661 ( .A(n22326), .B(n22325), .Z(n22327) );
  IV U22662 ( .A(n22327), .Z(n22543) );
  NOR U22663 ( .A(n22544), .B(n22543), .Z(n22328) );
  NOR U22664 ( .A(n22329), .B(n22328), .Z(n22330) );
  IV U22665 ( .A(n22330), .Z(n22542) );
  XOR U22666 ( .A(n22332), .B(n22331), .Z(n22541) );
  NOR U22667 ( .A(n22542), .B(n22541), .Z(n22333) );
  NOR U22668 ( .A(n22334), .B(n22333), .Z(n22335) );
  IV U22669 ( .A(n22335), .Z(n22539) );
  XOR U22670 ( .A(n22337), .B(n22336), .Z(n22338) );
  IV U22671 ( .A(n22338), .Z(n22538) );
  NOR U22672 ( .A(n22539), .B(n22538), .Z(n22339) );
  NOR U22673 ( .A(n22340), .B(n22339), .Z(n22341) );
  IV U22674 ( .A(n22341), .Z(n22537) );
  XOR U22675 ( .A(n22343), .B(n22342), .Z(n22536) );
  NOR U22676 ( .A(n22537), .B(n22536), .Z(n22344) );
  NOR U22677 ( .A(n22345), .B(n22344), .Z(n22346) );
  IV U22678 ( .A(n22346), .Z(n22534) );
  XOR U22679 ( .A(n22348), .B(n22347), .Z(n22349) );
  IV U22680 ( .A(n22349), .Z(n22533) );
  NOR U22681 ( .A(n22534), .B(n22533), .Z(n22350) );
  NOR U22682 ( .A(n22351), .B(n22350), .Z(n22352) );
  IV U22683 ( .A(n22352), .Z(n22532) );
  XOR U22684 ( .A(n22354), .B(n22353), .Z(n22531) );
  NOR U22685 ( .A(n22532), .B(n22531), .Z(n22355) );
  NOR U22686 ( .A(n22356), .B(n22355), .Z(n22357) );
  IV U22687 ( .A(n22357), .Z(n22527) );
  XOR U22688 ( .A(n22359), .B(n22358), .Z(n22360) );
  IV U22689 ( .A(n22360), .Z(n22526) );
  NOR U22690 ( .A(n22527), .B(n22526), .Z(n22361) );
  NOR U22691 ( .A(n22362), .B(n22361), .Z(n22363) );
  IV U22692 ( .A(n22363), .Z(n22525) );
  XOR U22693 ( .A(n22365), .B(n22364), .Z(n22524) );
  NOR U22694 ( .A(n22525), .B(n22524), .Z(n22366) );
  NOR U22695 ( .A(n22367), .B(n22366), .Z(n22368) );
  IV U22696 ( .A(n22368), .Z(n22522) );
  NOR U22697 ( .A(n22523), .B(n22522), .Z(n22369) );
  NOR U22698 ( .A(n22370), .B(n22369), .Z(n22371) );
  IV U22699 ( .A(n22371), .Z(n22518) );
  XOR U22700 ( .A(n22373), .B(n22372), .Z(n22517) );
  NOR U22701 ( .A(n22518), .B(n22517), .Z(n22374) );
  NOR U22702 ( .A(n22375), .B(n22374), .Z(n22514) );
  XOR U22703 ( .A(n22377), .B(n22376), .Z(n22513) );
  NOR U22704 ( .A(n22514), .B(n22513), .Z(n22378) );
  NOR U22705 ( .A(n22379), .B(n22378), .Z(n22509) );
  XOR U22706 ( .A(n22381), .B(n22380), .Z(n22508) );
  NOR U22707 ( .A(n22509), .B(n22508), .Z(n22382) );
  NOR U22708 ( .A(n22383), .B(n22382), .Z(n22502) );
  XOR U22709 ( .A(n22385), .B(n22384), .Z(n22503) );
  NOR U22710 ( .A(n22502), .B(n22503), .Z(n22386) );
  NOR U22711 ( .A(n22387), .B(n22386), .Z(n22499) );
  XOR U22712 ( .A(n22389), .B(n22388), .Z(n22498) );
  NOR U22713 ( .A(n22499), .B(n22498), .Z(n22390) );
  NOR U22714 ( .A(n22391), .B(n22390), .Z(n22394) );
  NOR U22715 ( .A(n145), .B(n68), .Z(n22392) );
  IV U22716 ( .A(n22392), .Z(n22393) );
  NOR U22717 ( .A(n22394), .B(n22393), .Z(n22399) );
  XOR U22718 ( .A(n22394), .B(n22393), .Z(n22911) );
  IV U22719 ( .A(n22911), .Z(n22397) );
  XOR U22720 ( .A(n22396), .B(n22395), .Z(n22910) );
  NOR U22721 ( .A(n22397), .B(n22910), .Z(n22398) );
  NOR U22722 ( .A(n22399), .B(n22398), .Z(n22404) );
  XOR U22723 ( .A(n22401), .B(n22400), .Z(n22403) );
  IV U22724 ( .A(n22403), .Z(n22402) );
  NOR U22725 ( .A(n22404), .B(n22402), .Z(n22407) );
  XOR U22726 ( .A(n22404), .B(n22403), .Z(n22920) );
  NOR U22727 ( .A(n147), .B(n68), .Z(n22919) );
  IV U22728 ( .A(n22919), .Z(n22405) );
  NOR U22729 ( .A(n22920), .B(n22405), .Z(n22406) );
  NOR U22730 ( .A(n22407), .B(n22406), .Z(n22924) );
  XOR U22731 ( .A(n22409), .B(n22408), .Z(n22923) );
  NOR U22732 ( .A(n22924), .B(n22923), .Z(n22410) );
  NOR U22733 ( .A(n22411), .B(n22410), .Z(n22414) );
  NOR U22734 ( .A(n150), .B(n68), .Z(n22413) );
  IV U22735 ( .A(n22413), .Z(n22412) );
  NOR U22736 ( .A(n22414), .B(n22412), .Z(n22418) );
  XOR U22737 ( .A(n22414), .B(n22413), .Z(n22494) );
  XOR U22738 ( .A(n22416), .B(n22415), .Z(n22495) );
  NOR U22739 ( .A(n22494), .B(n22495), .Z(n22417) );
  NOR U22740 ( .A(n22418), .B(n22417), .Z(n22423) );
  NOR U22741 ( .A(n153), .B(n68), .Z(n22422) );
  IV U22742 ( .A(n22422), .Z(n22419) );
  NOR U22743 ( .A(n22423), .B(n22419), .Z(n22426) );
  XOR U22744 ( .A(n22421), .B(n22420), .Z(n22936) );
  IV U22745 ( .A(n22936), .Z(n22424) );
  XOR U22746 ( .A(n22423), .B(n22422), .Z(n22935) );
  NOR U22747 ( .A(n22424), .B(n22935), .Z(n22425) );
  NOR U22748 ( .A(n22426), .B(n22425), .Z(n22430) );
  IV U22749 ( .A(n22430), .Z(n22427) );
  NOR U22750 ( .A(n22431), .B(n22427), .Z(n22433) );
  XOR U22751 ( .A(n22429), .B(n22428), .Z(n22945) );
  XOR U22752 ( .A(n22431), .B(n22430), .Z(n22944) );
  NOR U22753 ( .A(n22945), .B(n22944), .Z(n22432) );
  NOR U22754 ( .A(n22433), .B(n22432), .Z(n22434) );
  IV U22755 ( .A(n22434), .Z(n22439) );
  NOR U22756 ( .A(n156), .B(n68), .Z(n22438) );
  IV U22757 ( .A(n22438), .Z(n22435) );
  NOR U22758 ( .A(n22439), .B(n22435), .Z(n22441) );
  XOR U22759 ( .A(n22437), .B(n22436), .Z(n22951) );
  XOR U22760 ( .A(n22439), .B(n22438), .Z(n22952) );
  NOR U22761 ( .A(n22951), .B(n22952), .Z(n22440) );
  NOR U22762 ( .A(n22441), .B(n22440), .Z(n22448) );
  NOR U22763 ( .A(n158), .B(n68), .Z(n22447) );
  IV U22764 ( .A(n22447), .Z(n22442) );
  NOR U22765 ( .A(n22448), .B(n22442), .Z(n22451) );
  XOR U22766 ( .A(n22444), .B(n22443), .Z(n22445) );
  XOR U22767 ( .A(n22446), .B(n22445), .Z(n22959) );
  IV U22768 ( .A(n22959), .Z(n22449) );
  XOR U22769 ( .A(n22448), .B(n22447), .Z(n22958) );
  NOR U22770 ( .A(n22449), .B(n22958), .Z(n22450) );
  NOR U22771 ( .A(n22451), .B(n22450), .Z(n22456) );
  XOR U22772 ( .A(n22453), .B(n22452), .Z(n22455) );
  IV U22773 ( .A(n22455), .Z(n22454) );
  NOR U22774 ( .A(n22456), .B(n22454), .Z(n22459) );
  XOR U22775 ( .A(n22456), .B(n22455), .Z(n22491) );
  NOR U22776 ( .A(n161), .B(n68), .Z(n22492) );
  IV U22777 ( .A(n22492), .Z(n22457) );
  NOR U22778 ( .A(n22491), .B(n22457), .Z(n22458) );
  NOR U22779 ( .A(n22459), .B(n22458), .Z(n22462) );
  NOR U22780 ( .A(n163), .B(n68), .Z(n22461) );
  IV U22781 ( .A(n22461), .Z(n22460) );
  NOR U22782 ( .A(n22462), .B(n22460), .Z(n22466) );
  XOR U22783 ( .A(n22462), .B(n22461), .Z(n22971) );
  XOR U22784 ( .A(n22464), .B(n22463), .Z(n22972) );
  NOR U22785 ( .A(n22971), .B(n22972), .Z(n22465) );
  NOR U22786 ( .A(n22466), .B(n22465), .Z(n22469) );
  NOR U22787 ( .A(n165), .B(n68), .Z(n22468) );
  IV U22788 ( .A(n22468), .Z(n22467) );
  NOR U22789 ( .A(n22469), .B(n22467), .Z(n22474) );
  XOR U22790 ( .A(n22469), .B(n22468), .Z(n22979) );
  XOR U22791 ( .A(n22471), .B(n22470), .Z(n22978) );
  IV U22792 ( .A(n22978), .Z(n22472) );
  NOR U22793 ( .A(n22979), .B(n22472), .Z(n22473) );
  NOR U22794 ( .A(n22474), .B(n22473), .Z(n22479) );
  XOR U22795 ( .A(n22476), .B(n22475), .Z(n22478) );
  IV U22796 ( .A(n22478), .Z(n22477) );
  NOR U22797 ( .A(n22479), .B(n22477), .Z(n22482) );
  XOR U22798 ( .A(n22479), .B(n22478), .Z(n22489) );
  NOR U22799 ( .A(n167), .B(n68), .Z(n22480) );
  IV U22800 ( .A(n22480), .Z(n22490) );
  NOR U22801 ( .A(n22489), .B(n22490), .Z(n22481) );
  NOR U22802 ( .A(n22482), .B(n22481), .Z(n23976) );
  XOR U22803 ( .A(n22484), .B(n22483), .Z(n23975) );
  NOR U22804 ( .A(n23976), .B(n23975), .Z(n31538) );
  IV U22805 ( .A(n31538), .Z(n22487) );
  XOR U22806 ( .A(n22486), .B(n22485), .Z(n22488) );
  IV U22807 ( .A(n22488), .Z(n31537) );
  NOR U22808 ( .A(n22487), .B(n31537), .Z(n28535) );
  NOR U22809 ( .A(n31538), .B(n22488), .Z(n28533) );
  XOR U22810 ( .A(n22490), .B(n22489), .Z(n28520) );
  XOR U22811 ( .A(n22492), .B(n22491), .Z(n22966) );
  NOR U22812 ( .A(n163), .B(n69), .Z(n22967) );
  IV U22813 ( .A(n22967), .Z(n22493) );
  NOR U22814 ( .A(n22966), .B(n22493), .Z(n22969) );
  IV U22815 ( .A(n22494), .Z(n22496) );
  XOR U22816 ( .A(n22496), .B(n22495), .Z(n22932) );
  NOR U22817 ( .A(n153), .B(n69), .Z(n22931) );
  IV U22818 ( .A(n22931), .Z(n22497) );
  NOR U22819 ( .A(n22932), .B(n22497), .Z(n22934) );
  XOR U22820 ( .A(n22499), .B(n22498), .Z(n22500) );
  NOR U22821 ( .A(n145), .B(n69), .Z(n23399) );
  NOR U22822 ( .A(n22500), .B(n23399), .Z(n22907) );
  IV U22823 ( .A(n22500), .Z(n23396) );
  IV U22824 ( .A(n23399), .Z(n22501) );
  NOR U22825 ( .A(n23396), .B(n22501), .Z(n22905) );
  XOR U22826 ( .A(n22503), .B(n22502), .Z(n22504) );
  IV U22827 ( .A(n22504), .Z(n22506) );
  NOR U22828 ( .A(n143), .B(n69), .Z(n22507) );
  IV U22829 ( .A(n22507), .Z(n22505) );
  NOR U22830 ( .A(n22506), .B(n22505), .Z(n22903) );
  XOR U22831 ( .A(n22507), .B(n22506), .Z(n22992) );
  XOR U22832 ( .A(n22509), .B(n22508), .Z(n22510) );
  NOR U22833 ( .A(n141), .B(n69), .Z(n22511) );
  NOR U22834 ( .A(n22510), .B(n22511), .Z(n22900) );
  XOR U22835 ( .A(n22511), .B(n22510), .Z(n22512) );
  IV U22836 ( .A(n22512), .Z(n22997) );
  IV U22837 ( .A(n22513), .Z(n22515) );
  XOR U22838 ( .A(n22515), .B(n22514), .Z(n22894) );
  NOR U22839 ( .A(n139), .B(n69), .Z(n22895) );
  IV U22840 ( .A(n22895), .Z(n22516) );
  NOR U22841 ( .A(n22894), .B(n22516), .Z(n22897) );
  NOR U22842 ( .A(n137), .B(n69), .Z(n22520) );
  XOR U22843 ( .A(n22518), .B(n22517), .Z(n22519) );
  NOR U22844 ( .A(n22520), .B(n22519), .Z(n22892) );
  XOR U22845 ( .A(n22520), .B(n22519), .Z(n22521) );
  IV U22846 ( .A(n22521), .Z(n23004) );
  XOR U22847 ( .A(n22523), .B(n22522), .Z(n22886) );
  NOR U22848 ( .A(n133), .B(n69), .Z(n22880) );
  XOR U22849 ( .A(n22525), .B(n22524), .Z(n22879) );
  NOR U22850 ( .A(n22880), .B(n22879), .Z(n22883) );
  XOR U22851 ( .A(n22527), .B(n22526), .Z(n22530) );
  NOR U22852 ( .A(n131), .B(n69), .Z(n22529) );
  IV U22853 ( .A(n22529), .Z(n22528) );
  NOR U22854 ( .A(n22530), .B(n22528), .Z(n22877) );
  XOR U22855 ( .A(n22530), .B(n22529), .Z(n23013) );
  NOR U22856 ( .A(n128), .B(n69), .Z(n22871) );
  XOR U22857 ( .A(n22532), .B(n22531), .Z(n22870) );
  NOR U22858 ( .A(n22871), .B(n22870), .Z(n22874) );
  XOR U22859 ( .A(n22534), .B(n22533), .Z(n22866) );
  NOR U22860 ( .A(n126), .B(n69), .Z(n22865) );
  IV U22861 ( .A(n22865), .Z(n22535) );
  NOR U22862 ( .A(n22866), .B(n22535), .Z(n22868) );
  NOR U22863 ( .A(n125), .B(n69), .Z(n22860) );
  XOR U22864 ( .A(n22537), .B(n22536), .Z(n22859) );
  NOR U22865 ( .A(n22860), .B(n22859), .Z(n22863) );
  XOR U22866 ( .A(n22539), .B(n22538), .Z(n22855) );
  NOR U22867 ( .A(n123), .B(n69), .Z(n22854) );
  IV U22868 ( .A(n22854), .Z(n22540) );
  NOR U22869 ( .A(n22855), .B(n22540), .Z(n22857) );
  NOR U22870 ( .A(n120), .B(n69), .Z(n22849) );
  XOR U22871 ( .A(n22542), .B(n22541), .Z(n22848) );
  NOR U22872 ( .A(n22849), .B(n22848), .Z(n22852) );
  XOR U22873 ( .A(n22544), .B(n22543), .Z(n22844) );
  NOR U22874 ( .A(n119), .B(n69), .Z(n22843) );
  IV U22875 ( .A(n22843), .Z(n22545) );
  NOR U22876 ( .A(n22844), .B(n22545), .Z(n22846) );
  NOR U22877 ( .A(n79), .B(n69), .Z(n22838) );
  XOR U22878 ( .A(n22547), .B(n22546), .Z(n22837) );
  NOR U22879 ( .A(n22838), .B(n22837), .Z(n22841) );
  XOR U22880 ( .A(n22549), .B(n22548), .Z(n22833) );
  NOR U22881 ( .A(n117), .B(n69), .Z(n22832) );
  IV U22882 ( .A(n22832), .Z(n22550) );
  NOR U22883 ( .A(n22833), .B(n22550), .Z(n22835) );
  NOR U22884 ( .A(n80), .B(n69), .Z(n22827) );
  XOR U22885 ( .A(n22552), .B(n22551), .Z(n22826) );
  NOR U22886 ( .A(n22827), .B(n22826), .Z(n22830) );
  XOR U22887 ( .A(n22554), .B(n22553), .Z(n22822) );
  NOR U22888 ( .A(n116), .B(n69), .Z(n22821) );
  IV U22889 ( .A(n22821), .Z(n22555) );
  NOR U22890 ( .A(n22822), .B(n22555), .Z(n22824) );
  NOR U22891 ( .A(n81), .B(n69), .Z(n22816) );
  XOR U22892 ( .A(n22557), .B(n22556), .Z(n22815) );
  NOR U22893 ( .A(n22816), .B(n22815), .Z(n22819) );
  XOR U22894 ( .A(n22559), .B(n22558), .Z(n22811) );
  NOR U22895 ( .A(n115), .B(n69), .Z(n22810) );
  IV U22896 ( .A(n22810), .Z(n22560) );
  NOR U22897 ( .A(n22811), .B(n22560), .Z(n22813) );
  NOR U22898 ( .A(n82), .B(n69), .Z(n22805) );
  XOR U22899 ( .A(n22562), .B(n22561), .Z(n22804) );
  NOR U22900 ( .A(n22805), .B(n22804), .Z(n22808) );
  IV U22901 ( .A(n22563), .Z(n22565) );
  XOR U22902 ( .A(n22565), .B(n22564), .Z(n22799) );
  NOR U22903 ( .A(n114), .B(n69), .Z(n22800) );
  IV U22904 ( .A(n22800), .Z(n22566) );
  NOR U22905 ( .A(n22799), .B(n22566), .Z(n22802) );
  IV U22906 ( .A(n22567), .Z(n22569) );
  XOR U22907 ( .A(n22569), .B(n22568), .Z(n22795) );
  NOR U22908 ( .A(n83), .B(n69), .Z(n22796) );
  IV U22909 ( .A(n22796), .Z(n22570) );
  NOR U22910 ( .A(n22795), .B(n22570), .Z(n22798) );
  IV U22911 ( .A(n22571), .Z(n22573) );
  XOR U22912 ( .A(n22573), .B(n22572), .Z(n22791) );
  NOR U22913 ( .A(n113), .B(n69), .Z(n22792) );
  IV U22914 ( .A(n22792), .Z(n22574) );
  NOR U22915 ( .A(n22791), .B(n22574), .Z(n22794) );
  IV U22916 ( .A(n22575), .Z(n22577) );
  XOR U22917 ( .A(n22577), .B(n22576), .Z(n22787) );
  NOR U22918 ( .A(n84), .B(n69), .Z(n22788) );
  IV U22919 ( .A(n22788), .Z(n22578) );
  NOR U22920 ( .A(n22787), .B(n22578), .Z(n22790) );
  IV U22921 ( .A(n22579), .Z(n22581) );
  XOR U22922 ( .A(n22581), .B(n22580), .Z(n22783) );
  NOR U22923 ( .A(n112), .B(n69), .Z(n22784) );
  IV U22924 ( .A(n22784), .Z(n22582) );
  NOR U22925 ( .A(n22783), .B(n22582), .Z(n22786) );
  IV U22926 ( .A(n22583), .Z(n22585) );
  XOR U22927 ( .A(n22585), .B(n22584), .Z(n22779) );
  NOR U22928 ( .A(n85), .B(n69), .Z(n22780) );
  IV U22929 ( .A(n22780), .Z(n22586) );
  NOR U22930 ( .A(n22779), .B(n22586), .Z(n22782) );
  IV U22931 ( .A(n22587), .Z(n22589) );
  XOR U22932 ( .A(n22589), .B(n22588), .Z(n22775) );
  NOR U22933 ( .A(n111), .B(n69), .Z(n22776) );
  IV U22934 ( .A(n22776), .Z(n22590) );
  NOR U22935 ( .A(n22775), .B(n22590), .Z(n22778) );
  IV U22936 ( .A(n22591), .Z(n22593) );
  XOR U22937 ( .A(n22593), .B(n22592), .Z(n22771) );
  NOR U22938 ( .A(n86), .B(n69), .Z(n22772) );
  IV U22939 ( .A(n22772), .Z(n22594) );
  NOR U22940 ( .A(n22771), .B(n22594), .Z(n22774) );
  IV U22941 ( .A(n22595), .Z(n22597) );
  XOR U22942 ( .A(n22597), .B(n22596), .Z(n22767) );
  NOR U22943 ( .A(n110), .B(n69), .Z(n22768) );
  IV U22944 ( .A(n22768), .Z(n22598) );
  NOR U22945 ( .A(n22767), .B(n22598), .Z(n22770) );
  XOR U22946 ( .A(n22600), .B(n22599), .Z(n22763) );
  NOR U22947 ( .A(n109), .B(n69), .Z(n22764) );
  IV U22948 ( .A(n22764), .Z(n22601) );
  NOR U22949 ( .A(n22763), .B(n22601), .Z(n22766) );
  IV U22950 ( .A(n22602), .Z(n22604) );
  XOR U22951 ( .A(n22604), .B(n22603), .Z(n22751) );
  NOR U22952 ( .A(n87), .B(n69), .Z(n22752) );
  IV U22953 ( .A(n22752), .Z(n22605) );
  NOR U22954 ( .A(n22751), .B(n22605), .Z(n22754) );
  IV U22955 ( .A(n22606), .Z(n22608) );
  XOR U22956 ( .A(n22608), .B(n22607), .Z(n22747) );
  NOR U22957 ( .A(n107), .B(n69), .Z(n22748) );
  IV U22958 ( .A(n22748), .Z(n22609) );
  NOR U22959 ( .A(n22747), .B(n22609), .Z(n22750) );
  IV U22960 ( .A(n22610), .Z(n22612) );
  XOR U22961 ( .A(n22612), .B(n22611), .Z(n22743) );
  NOR U22962 ( .A(n88), .B(n69), .Z(n22744) );
  IV U22963 ( .A(n22744), .Z(n22613) );
  NOR U22964 ( .A(n22743), .B(n22613), .Z(n22746) );
  IV U22965 ( .A(n22614), .Z(n22616) );
  XOR U22966 ( .A(n22616), .B(n22615), .Z(n22739) );
  NOR U22967 ( .A(n106), .B(n69), .Z(n22740) );
  IV U22968 ( .A(n22740), .Z(n22617) );
  NOR U22969 ( .A(n22739), .B(n22617), .Z(n22742) );
  XOR U22970 ( .A(n22619), .B(n22618), .Z(n22735) );
  NOR U22971 ( .A(n105), .B(n69), .Z(n22736) );
  IV U22972 ( .A(n22736), .Z(n22620) );
  NOR U22973 ( .A(n22735), .B(n22620), .Z(n22738) );
  XOR U22974 ( .A(n22622), .B(n22621), .Z(n22723) );
  IV U22975 ( .A(n22723), .Z(n22624) );
  NOR U22976 ( .A(n89), .B(n69), .Z(n22623) );
  IV U22977 ( .A(n22623), .Z(n22724) );
  NOR U22978 ( .A(n22624), .B(n22724), .Z(n22726) );
  IV U22979 ( .A(n22625), .Z(n22627) );
  XOR U22980 ( .A(n22627), .B(n22626), .Z(n22719) );
  NOR U22981 ( .A(n103), .B(n69), .Z(n22720) );
  IV U22982 ( .A(n22720), .Z(n22628) );
  NOR U22983 ( .A(n22719), .B(n22628), .Z(n22722) );
  IV U22984 ( .A(n22629), .Z(n22631) );
  XOR U22985 ( .A(n22631), .B(n22630), .Z(n22715) );
  NOR U22986 ( .A(n90), .B(n69), .Z(n22716) );
  IV U22987 ( .A(n22716), .Z(n22632) );
  NOR U22988 ( .A(n22715), .B(n22632), .Z(n22718) );
  IV U22989 ( .A(n22633), .Z(n22635) );
  XOR U22990 ( .A(n22635), .B(n22634), .Z(n22711) );
  NOR U22991 ( .A(n102), .B(n69), .Z(n22712) );
  IV U22992 ( .A(n22712), .Z(n22636) );
  NOR U22993 ( .A(n22711), .B(n22636), .Z(n22714) );
  IV U22994 ( .A(n22637), .Z(n22639) );
  XOR U22995 ( .A(n22639), .B(n22638), .Z(n22707) );
  NOR U22996 ( .A(n101), .B(n69), .Z(n22708) );
  IV U22997 ( .A(n22708), .Z(n22640) );
  NOR U22998 ( .A(n22707), .B(n22640), .Z(n22710) );
  IV U22999 ( .A(n22641), .Z(n22643) );
  XOR U23000 ( .A(n22643), .B(n22642), .Z(n22703) );
  NOR U23001 ( .A(n100), .B(n69), .Z(n22704) );
  IV U23002 ( .A(n22704), .Z(n22644) );
  NOR U23003 ( .A(n22703), .B(n22644), .Z(n22706) );
  IV U23004 ( .A(n22645), .Z(n22647) );
  XOR U23005 ( .A(n22647), .B(n22646), .Z(n22699) );
  NOR U23006 ( .A(n99), .B(n69), .Z(n22700) );
  IV U23007 ( .A(n22700), .Z(n22648) );
  NOR U23008 ( .A(n22699), .B(n22648), .Z(n22702) );
  IV U23009 ( .A(n22649), .Z(n22651) );
  XOR U23010 ( .A(n22651), .B(n22650), .Z(n22695) );
  NOR U23011 ( .A(n98), .B(n69), .Z(n22696) );
  IV U23012 ( .A(n22696), .Z(n22652) );
  NOR U23013 ( .A(n22695), .B(n22652), .Z(n22698) );
  XOR U23014 ( .A(n22654), .B(n22653), .Z(n22691) );
  NOR U23015 ( .A(n91), .B(n69), .Z(n22692) );
  IV U23016 ( .A(n22692), .Z(n22655) );
  NOR U23017 ( .A(n22691), .B(n22655), .Z(n22694) );
  XOR U23018 ( .A(n22657), .B(n22656), .Z(n22679) );
  IV U23019 ( .A(n22679), .Z(n22659) );
  NOR U23020 ( .A(n96), .B(n69), .Z(n22658) );
  IV U23021 ( .A(n22658), .Z(n22680) );
  NOR U23022 ( .A(n22659), .B(n22680), .Z(n22682) );
  NOR U23023 ( .A(n95), .B(n69), .Z(n22676) );
  IV U23024 ( .A(n22676), .Z(n22662) );
  XOR U23025 ( .A(n22661), .B(n22660), .Z(n22675) );
  NOR U23026 ( .A(n22662), .B(n22675), .Z(n22678) );
  NOR U23027 ( .A(n93), .B(n69), .Z(n23628) );
  IV U23028 ( .A(n23628), .Z(n22663) );
  NOR U23029 ( .A(n68), .B(n168), .Z(n22671) );
  IV U23030 ( .A(n22671), .Z(n22666) );
  NOR U23031 ( .A(n22663), .B(n22666), .Z(n22664) );
  IV U23032 ( .A(n22664), .Z(n22665) );
  NOR U23033 ( .A(n94), .B(n22665), .Z(n22674) );
  NOR U23034 ( .A(n22666), .B(n93), .Z(n22667) );
  XOR U23035 ( .A(n94), .B(n22667), .Z(n22668) );
  NOR U23036 ( .A(n69), .B(n22668), .Z(n22669) );
  IV U23037 ( .A(n22669), .Z(n23161) );
  XOR U23038 ( .A(n22671), .B(n22670), .Z(n23160) );
  IV U23039 ( .A(n23160), .Z(n22672) );
  NOR U23040 ( .A(n23161), .B(n22672), .Z(n22673) );
  NOR U23041 ( .A(n22674), .B(n22673), .Z(n23157) );
  XOR U23042 ( .A(n22676), .B(n22675), .Z(n23156) );
  NOR U23043 ( .A(n23157), .B(n23156), .Z(n22677) );
  NOR U23044 ( .A(n22678), .B(n22677), .Z(n23184) );
  XOR U23045 ( .A(n22680), .B(n22679), .Z(n23183) );
  NOR U23046 ( .A(n23184), .B(n23183), .Z(n22681) );
  NOR U23047 ( .A(n22682), .B(n22681), .Z(n22687) );
  XOR U23048 ( .A(n22684), .B(n22683), .Z(n22686) );
  IV U23049 ( .A(n22686), .Z(n22685) );
  NOR U23050 ( .A(n22687), .B(n22685), .Z(n22690) );
  XOR U23051 ( .A(n22687), .B(n22686), .Z(n23153) );
  NOR U23052 ( .A(n97), .B(n69), .Z(n23154) );
  IV U23053 ( .A(n23154), .Z(n22688) );
  NOR U23054 ( .A(n23153), .B(n22688), .Z(n22689) );
  NOR U23055 ( .A(n22690), .B(n22689), .Z(n23149) );
  XOR U23056 ( .A(n22692), .B(n22691), .Z(n23150) );
  NOR U23057 ( .A(n23149), .B(n23150), .Z(n22693) );
  NOR U23058 ( .A(n22694), .B(n22693), .Z(n23145) );
  XOR U23059 ( .A(n22696), .B(n22695), .Z(n23146) );
  NOR U23060 ( .A(n23145), .B(n23146), .Z(n22697) );
  NOR U23061 ( .A(n22698), .B(n22697), .Z(n23141) );
  XOR U23062 ( .A(n22700), .B(n22699), .Z(n23142) );
  NOR U23063 ( .A(n23141), .B(n23142), .Z(n22701) );
  NOR U23064 ( .A(n22702), .B(n22701), .Z(n23137) );
  XOR U23065 ( .A(n22704), .B(n22703), .Z(n23138) );
  NOR U23066 ( .A(n23137), .B(n23138), .Z(n22705) );
  NOR U23067 ( .A(n22706), .B(n22705), .Z(n23133) );
  XOR U23068 ( .A(n22708), .B(n22707), .Z(n23134) );
  NOR U23069 ( .A(n23133), .B(n23134), .Z(n22709) );
  NOR U23070 ( .A(n22710), .B(n22709), .Z(n23129) );
  XOR U23071 ( .A(n22712), .B(n22711), .Z(n23130) );
  NOR U23072 ( .A(n23129), .B(n23130), .Z(n22713) );
  NOR U23073 ( .A(n22714), .B(n22713), .Z(n23125) );
  XOR U23074 ( .A(n22716), .B(n22715), .Z(n23126) );
  NOR U23075 ( .A(n23125), .B(n23126), .Z(n22717) );
  NOR U23076 ( .A(n22718), .B(n22717), .Z(n23122) );
  XOR U23077 ( .A(n22720), .B(n22719), .Z(n23121) );
  NOR U23078 ( .A(n23122), .B(n23121), .Z(n22721) );
  NOR U23079 ( .A(n22722), .B(n22721), .Z(n23228) );
  XOR U23080 ( .A(n22724), .B(n22723), .Z(n23227) );
  NOR U23081 ( .A(n23228), .B(n23227), .Z(n22725) );
  NOR U23082 ( .A(n22726), .B(n22725), .Z(n22731) );
  XOR U23083 ( .A(n22728), .B(n22727), .Z(n22730) );
  IV U23084 ( .A(n22730), .Z(n22729) );
  NOR U23085 ( .A(n22731), .B(n22729), .Z(n22734) );
  XOR U23086 ( .A(n22731), .B(n22730), .Z(n23118) );
  NOR U23087 ( .A(n104), .B(n69), .Z(n23119) );
  IV U23088 ( .A(n23119), .Z(n22732) );
  NOR U23089 ( .A(n23118), .B(n22732), .Z(n22733) );
  NOR U23090 ( .A(n22734), .B(n22733), .Z(n23114) );
  XOR U23091 ( .A(n22736), .B(n22735), .Z(n23115) );
  NOR U23092 ( .A(n23114), .B(n23115), .Z(n22737) );
  NOR U23093 ( .A(n22738), .B(n22737), .Z(n23110) );
  XOR U23094 ( .A(n22740), .B(n22739), .Z(n23111) );
  NOR U23095 ( .A(n23110), .B(n23111), .Z(n22741) );
  NOR U23096 ( .A(n22742), .B(n22741), .Z(n23106) );
  XOR U23097 ( .A(n22744), .B(n22743), .Z(n23107) );
  NOR U23098 ( .A(n23106), .B(n23107), .Z(n22745) );
  NOR U23099 ( .A(n22746), .B(n22745), .Z(n23103) );
  XOR U23100 ( .A(n22748), .B(n22747), .Z(n23102) );
  NOR U23101 ( .A(n23103), .B(n23102), .Z(n22749) );
  NOR U23102 ( .A(n22750), .B(n22749), .Z(n23098) );
  XOR U23103 ( .A(n22752), .B(n22751), .Z(n23099) );
  NOR U23104 ( .A(n23098), .B(n23099), .Z(n22753) );
  NOR U23105 ( .A(n22754), .B(n22753), .Z(n22757) );
  NOR U23106 ( .A(n108), .B(n69), .Z(n22756) );
  IV U23107 ( .A(n22756), .Z(n22755) );
  NOR U23108 ( .A(n22757), .B(n22755), .Z(n22762) );
  XOR U23109 ( .A(n22757), .B(n22756), .Z(n23095) );
  XOR U23110 ( .A(n22759), .B(n22758), .Z(n23096) );
  IV U23111 ( .A(n23096), .Z(n22760) );
  NOR U23112 ( .A(n23095), .B(n22760), .Z(n22761) );
  NOR U23113 ( .A(n22762), .B(n22761), .Z(n23091) );
  XOR U23114 ( .A(n22764), .B(n22763), .Z(n23092) );
  NOR U23115 ( .A(n23091), .B(n23092), .Z(n22765) );
  NOR U23116 ( .A(n22766), .B(n22765), .Z(n23087) );
  XOR U23117 ( .A(n22768), .B(n22767), .Z(n23088) );
  NOR U23118 ( .A(n23087), .B(n23088), .Z(n22769) );
  NOR U23119 ( .A(n22770), .B(n22769), .Z(n23083) );
  XOR U23120 ( .A(n22772), .B(n22771), .Z(n23084) );
  NOR U23121 ( .A(n23083), .B(n23084), .Z(n22773) );
  NOR U23122 ( .A(n22774), .B(n22773), .Z(n23079) );
  XOR U23123 ( .A(n22776), .B(n22775), .Z(n23080) );
  NOR U23124 ( .A(n23079), .B(n23080), .Z(n22777) );
  NOR U23125 ( .A(n22778), .B(n22777), .Z(n23075) );
  XOR U23126 ( .A(n22780), .B(n22779), .Z(n23076) );
  NOR U23127 ( .A(n23075), .B(n23076), .Z(n22781) );
  NOR U23128 ( .A(n22782), .B(n22781), .Z(n23071) );
  XOR U23129 ( .A(n22784), .B(n22783), .Z(n23072) );
  NOR U23130 ( .A(n23071), .B(n23072), .Z(n22785) );
  NOR U23131 ( .A(n22786), .B(n22785), .Z(n23067) );
  XOR U23132 ( .A(n22788), .B(n22787), .Z(n23068) );
  NOR U23133 ( .A(n23067), .B(n23068), .Z(n22789) );
  NOR U23134 ( .A(n22790), .B(n22789), .Z(n23063) );
  XOR U23135 ( .A(n22792), .B(n22791), .Z(n23064) );
  NOR U23136 ( .A(n23063), .B(n23064), .Z(n22793) );
  NOR U23137 ( .A(n22794), .B(n22793), .Z(n23059) );
  XOR U23138 ( .A(n22796), .B(n22795), .Z(n23060) );
  NOR U23139 ( .A(n23059), .B(n23060), .Z(n22797) );
  NOR U23140 ( .A(n22798), .B(n22797), .Z(n23055) );
  XOR U23141 ( .A(n22800), .B(n22799), .Z(n23056) );
  NOR U23142 ( .A(n23055), .B(n23056), .Z(n22801) );
  NOR U23143 ( .A(n22802), .B(n22801), .Z(n22803) );
  IV U23144 ( .A(n22803), .Z(n23053) );
  XOR U23145 ( .A(n22805), .B(n22804), .Z(n22806) );
  IV U23146 ( .A(n22806), .Z(n23052) );
  NOR U23147 ( .A(n23053), .B(n23052), .Z(n22807) );
  NOR U23148 ( .A(n22808), .B(n22807), .Z(n22809) );
  IV U23149 ( .A(n22809), .Z(n23051) );
  XOR U23150 ( .A(n22811), .B(n22810), .Z(n23050) );
  NOR U23151 ( .A(n23051), .B(n23050), .Z(n22812) );
  NOR U23152 ( .A(n22813), .B(n22812), .Z(n22814) );
  IV U23153 ( .A(n22814), .Z(n23048) );
  XOR U23154 ( .A(n22816), .B(n22815), .Z(n22817) );
  IV U23155 ( .A(n22817), .Z(n23047) );
  NOR U23156 ( .A(n23048), .B(n23047), .Z(n22818) );
  NOR U23157 ( .A(n22819), .B(n22818), .Z(n22820) );
  IV U23158 ( .A(n22820), .Z(n23043) );
  XOR U23159 ( .A(n22822), .B(n22821), .Z(n23042) );
  NOR U23160 ( .A(n23043), .B(n23042), .Z(n22823) );
  NOR U23161 ( .A(n22824), .B(n22823), .Z(n22825) );
  IV U23162 ( .A(n22825), .Z(n23040) );
  XOR U23163 ( .A(n22827), .B(n22826), .Z(n22828) );
  IV U23164 ( .A(n22828), .Z(n23039) );
  NOR U23165 ( .A(n23040), .B(n23039), .Z(n22829) );
  NOR U23166 ( .A(n22830), .B(n22829), .Z(n22831) );
  IV U23167 ( .A(n22831), .Z(n23038) );
  XOR U23168 ( .A(n22833), .B(n22832), .Z(n23037) );
  NOR U23169 ( .A(n23038), .B(n23037), .Z(n22834) );
  NOR U23170 ( .A(n22835), .B(n22834), .Z(n22836) );
  IV U23171 ( .A(n22836), .Z(n23035) );
  XOR U23172 ( .A(n22838), .B(n22837), .Z(n22839) );
  IV U23173 ( .A(n22839), .Z(n23034) );
  NOR U23174 ( .A(n23035), .B(n23034), .Z(n22840) );
  NOR U23175 ( .A(n22841), .B(n22840), .Z(n22842) );
  IV U23176 ( .A(n22842), .Z(n23033) );
  XOR U23177 ( .A(n22844), .B(n22843), .Z(n23032) );
  NOR U23178 ( .A(n23033), .B(n23032), .Z(n22845) );
  NOR U23179 ( .A(n22846), .B(n22845), .Z(n22847) );
  IV U23180 ( .A(n22847), .Z(n23030) );
  XOR U23181 ( .A(n22849), .B(n22848), .Z(n22850) );
  IV U23182 ( .A(n22850), .Z(n23029) );
  NOR U23183 ( .A(n23030), .B(n23029), .Z(n22851) );
  NOR U23184 ( .A(n22852), .B(n22851), .Z(n22853) );
  IV U23185 ( .A(n22853), .Z(n23028) );
  XOR U23186 ( .A(n22855), .B(n22854), .Z(n23027) );
  NOR U23187 ( .A(n23028), .B(n23027), .Z(n22856) );
  NOR U23188 ( .A(n22857), .B(n22856), .Z(n22858) );
  IV U23189 ( .A(n22858), .Z(n23025) );
  XOR U23190 ( .A(n22860), .B(n22859), .Z(n22861) );
  IV U23191 ( .A(n22861), .Z(n23024) );
  NOR U23192 ( .A(n23025), .B(n23024), .Z(n22862) );
  NOR U23193 ( .A(n22863), .B(n22862), .Z(n22864) );
  IV U23194 ( .A(n22864), .Z(n23023) );
  XOR U23195 ( .A(n22866), .B(n22865), .Z(n23022) );
  NOR U23196 ( .A(n23023), .B(n23022), .Z(n22867) );
  NOR U23197 ( .A(n22868), .B(n22867), .Z(n22869) );
  IV U23198 ( .A(n22869), .Z(n23018) );
  XOR U23199 ( .A(n22871), .B(n22870), .Z(n22872) );
  IV U23200 ( .A(n22872), .Z(n23017) );
  NOR U23201 ( .A(n23018), .B(n23017), .Z(n22873) );
  NOR U23202 ( .A(n22874), .B(n22873), .Z(n22875) );
  IV U23203 ( .A(n22875), .Z(n23012) );
  NOR U23204 ( .A(n23013), .B(n23012), .Z(n22876) );
  NOR U23205 ( .A(n22877), .B(n22876), .Z(n22878) );
  IV U23206 ( .A(n22878), .Z(n23010) );
  XOR U23207 ( .A(n22880), .B(n22879), .Z(n22881) );
  IV U23208 ( .A(n22881), .Z(n23009) );
  NOR U23209 ( .A(n23010), .B(n23009), .Z(n22882) );
  NOR U23210 ( .A(n22883), .B(n22882), .Z(n22885) );
  IV U23211 ( .A(n22885), .Z(n22884) );
  NOR U23212 ( .A(n22886), .B(n22884), .Z(n22889) );
  XOR U23213 ( .A(n22886), .B(n22885), .Z(n23006) );
  NOR U23214 ( .A(n135), .B(n69), .Z(n23007) );
  IV U23215 ( .A(n23007), .Z(n22887) );
  NOR U23216 ( .A(n23006), .B(n22887), .Z(n22888) );
  NOR U23217 ( .A(n22889), .B(n22888), .Z(n22890) );
  IV U23218 ( .A(n22890), .Z(n23003) );
  NOR U23219 ( .A(n23004), .B(n23003), .Z(n22891) );
  NOR U23220 ( .A(n22892), .B(n22891), .Z(n22893) );
  IV U23221 ( .A(n22893), .Z(n23002) );
  XOR U23222 ( .A(n22895), .B(n22894), .Z(n23001) );
  NOR U23223 ( .A(n23002), .B(n23001), .Z(n22896) );
  NOR U23224 ( .A(n22897), .B(n22896), .Z(n22898) );
  IV U23225 ( .A(n22898), .Z(n22996) );
  NOR U23226 ( .A(n22997), .B(n22996), .Z(n22899) );
  NOR U23227 ( .A(n22900), .B(n22899), .Z(n22901) );
  IV U23228 ( .A(n22901), .Z(n22993) );
  NOR U23229 ( .A(n22992), .B(n22993), .Z(n22902) );
  NOR U23230 ( .A(n22903), .B(n22902), .Z(n22904) );
  IV U23231 ( .A(n22904), .Z(n23397) );
  NOR U23232 ( .A(n22905), .B(n23397), .Z(n22906) );
  NOR U23233 ( .A(n22907), .B(n22906), .Z(n22913) );
  IV U23234 ( .A(n22913), .Z(n22909) );
  NOR U23235 ( .A(n147), .B(n69), .Z(n22908) );
  IV U23236 ( .A(n22908), .Z(n22912) );
  NOR U23237 ( .A(n22909), .B(n22912), .Z(n22915) );
  XOR U23238 ( .A(n22911), .B(n22910), .Z(n22988) );
  XOR U23239 ( .A(n22913), .B(n22912), .Z(n22987) );
  NOR U23240 ( .A(n22988), .B(n22987), .Z(n22914) );
  NOR U23241 ( .A(n22915), .B(n22914), .Z(n22918) );
  NOR U23242 ( .A(n148), .B(n69), .Z(n22917) );
  IV U23243 ( .A(n22917), .Z(n22916) );
  NOR U23244 ( .A(n22918), .B(n22916), .Z(n22922) );
  XOR U23245 ( .A(n22918), .B(n22917), .Z(n23410) );
  XOR U23246 ( .A(n22920), .B(n22919), .Z(n23409) );
  NOR U23247 ( .A(n23410), .B(n23409), .Z(n22921) );
  NOR U23248 ( .A(n22922), .B(n22921), .Z(n22927) );
  XOR U23249 ( .A(n22924), .B(n22923), .Z(n22926) );
  IV U23250 ( .A(n22926), .Z(n22925) );
  NOR U23251 ( .A(n22927), .B(n22925), .Z(n22930) );
  XOR U23252 ( .A(n22927), .B(n22926), .Z(n23421) );
  NOR U23253 ( .A(n150), .B(n69), .Z(n22928) );
  IV U23254 ( .A(n22928), .Z(n23422) );
  NOR U23255 ( .A(n23421), .B(n23422), .Z(n22929) );
  NOR U23256 ( .A(n22930), .B(n22929), .Z(n23430) );
  XOR U23257 ( .A(n22932), .B(n22931), .Z(n23429) );
  NOR U23258 ( .A(n23430), .B(n23429), .Z(n22933) );
  NOR U23259 ( .A(n22934), .B(n22933), .Z(n22938) );
  XOR U23260 ( .A(n22936), .B(n22935), .Z(n22937) );
  NOR U23261 ( .A(n22938), .B(n22937), .Z(n22942) );
  XOR U23262 ( .A(n22938), .B(n22937), .Z(n23435) );
  IV U23263 ( .A(n23435), .Z(n22940) );
  NOR U23264 ( .A(n155), .B(n69), .Z(n22939) );
  IV U23265 ( .A(n22939), .Z(n23436) );
  NOR U23266 ( .A(n22940), .B(n23436), .Z(n22941) );
  NOR U23267 ( .A(n22942), .B(n22941), .Z(n22947) );
  NOR U23268 ( .A(n156), .B(n69), .Z(n22946) );
  IV U23269 ( .A(n22946), .Z(n22943) );
  NOR U23270 ( .A(n22947), .B(n22943), .Z(n22949) );
  XOR U23271 ( .A(n22945), .B(n22944), .Z(n23443) );
  XOR U23272 ( .A(n22947), .B(n22946), .Z(n23442) );
  NOR U23273 ( .A(n23443), .B(n23442), .Z(n22948) );
  NOR U23274 ( .A(n22949), .B(n22948), .Z(n22954) );
  NOR U23275 ( .A(n158), .B(n69), .Z(n22953) );
  IV U23276 ( .A(n22953), .Z(n22950) );
  NOR U23277 ( .A(n22954), .B(n22950), .Z(n22957) );
  XOR U23278 ( .A(n22952), .B(n22951), .Z(n23450) );
  IV U23279 ( .A(n23450), .Z(n22955) );
  XOR U23280 ( .A(n22954), .B(n22953), .Z(n23449) );
  NOR U23281 ( .A(n22955), .B(n23449), .Z(n22956) );
  NOR U23282 ( .A(n22957), .B(n22956), .Z(n22961) );
  XOR U23283 ( .A(n22959), .B(n22958), .Z(n22960) );
  NOR U23284 ( .A(n22961), .B(n22960), .Z(n22965) );
  XOR U23285 ( .A(n22961), .B(n22960), .Z(n22962) );
  IV U23286 ( .A(n22962), .Z(n23921) );
  NOR U23287 ( .A(n161), .B(n69), .Z(n23920) );
  IV U23288 ( .A(n23920), .Z(n22963) );
  NOR U23289 ( .A(n23921), .B(n22963), .Z(n22964) );
  NOR U23290 ( .A(n22965), .B(n22964), .Z(n23935) );
  XOR U23291 ( .A(n22967), .B(n22966), .Z(n23934) );
  NOR U23292 ( .A(n23935), .B(n23934), .Z(n22968) );
  NOR U23293 ( .A(n22969), .B(n22968), .Z(n22974) );
  NOR U23294 ( .A(n165), .B(n69), .Z(n22973) );
  IV U23295 ( .A(n22973), .Z(n22970) );
  NOR U23296 ( .A(n22974), .B(n22970), .Z(n22977) );
  XOR U23297 ( .A(n22972), .B(n22971), .Z(n23950) );
  IV U23298 ( .A(n23950), .Z(n22975) );
  XOR U23299 ( .A(n22974), .B(n22973), .Z(n23949) );
  NOR U23300 ( .A(n22975), .B(n23949), .Z(n22976) );
  NOR U23301 ( .A(n22977), .B(n22976), .Z(n22980) );
  XOR U23302 ( .A(n22979), .B(n22978), .Z(n22981) );
  NOR U23303 ( .A(n22980), .B(n22981), .Z(n22985) );
  IV U23304 ( .A(n22980), .Z(n22982) );
  XOR U23305 ( .A(n22982), .B(n22981), .Z(n23967) );
  NOR U23306 ( .A(n167), .B(n69), .Z(n23968) );
  IV U23307 ( .A(n23968), .Z(n22983) );
  NOR U23308 ( .A(n23967), .B(n22983), .Z(n22984) );
  NOR U23309 ( .A(n22985), .B(n22984), .Z(n28521) );
  IV U23310 ( .A(n28521), .Z(n22986) );
  NOR U23311 ( .A(n28520), .B(n22986), .Z(n23980) );
  NOR U23312 ( .A(n158), .B(n70), .Z(n23445) );
  NOR U23313 ( .A(n148), .B(n70), .Z(n22990) );
  XOR U23314 ( .A(n22988), .B(n22987), .Z(n22989) );
  NOR U23315 ( .A(n22990), .B(n22989), .Z(n23408) );
  XOR U23316 ( .A(n22990), .B(n22989), .Z(n22991) );
  IV U23317 ( .A(n22991), .Z(n23873) );
  XOR U23318 ( .A(n22993), .B(n22992), .Z(n22995) );
  IV U23319 ( .A(n22995), .Z(n23456) );
  NOR U23320 ( .A(n145), .B(n70), .Z(n22994) );
  IV U23321 ( .A(n22994), .Z(n23455) );
  NOR U23322 ( .A(n23456), .B(n23455), .Z(n23395) );
  NOR U23323 ( .A(n22995), .B(n22994), .Z(n23393) );
  XOR U23324 ( .A(n22997), .B(n22996), .Z(n23000) );
  NOR U23325 ( .A(n143), .B(n70), .Z(n22999) );
  IV U23326 ( .A(n22999), .Z(n22998) );
  NOR U23327 ( .A(n23000), .B(n22998), .Z(n23392) );
  XOR U23328 ( .A(n23000), .B(n22999), .Z(n23460) );
  XOR U23329 ( .A(n23002), .B(n23001), .Z(n23385) );
  NOR U23330 ( .A(n141), .B(n70), .Z(n23386) );
  NOR U23331 ( .A(n23385), .B(n23386), .Z(n23389) );
  XOR U23332 ( .A(n23004), .B(n23003), .Z(n23381) );
  NOR U23333 ( .A(n139), .B(n70), .Z(n23380) );
  IV U23334 ( .A(n23380), .Z(n23005) );
  NOR U23335 ( .A(n23381), .B(n23005), .Z(n23383) );
  XOR U23336 ( .A(n23007), .B(n23006), .Z(n23376) );
  NOR U23337 ( .A(n137), .B(n70), .Z(n23377) );
  IV U23338 ( .A(n23377), .Z(n23008) );
  NOR U23339 ( .A(n23376), .B(n23008), .Z(n23379) );
  XOR U23340 ( .A(n23010), .B(n23009), .Z(n23372) );
  NOR U23341 ( .A(n135), .B(n70), .Z(n23371) );
  IV U23342 ( .A(n23371), .Z(n23011) );
  NOR U23343 ( .A(n23372), .B(n23011), .Z(n23375) );
  NOR U23344 ( .A(n133), .B(n70), .Z(n23015) );
  XOR U23345 ( .A(n23013), .B(n23012), .Z(n23014) );
  NOR U23346 ( .A(n23015), .B(n23014), .Z(n23370) );
  XOR U23347 ( .A(n23015), .B(n23014), .Z(n23016) );
  IV U23348 ( .A(n23016), .Z(n23475) );
  XOR U23349 ( .A(n23018), .B(n23017), .Z(n23021) );
  NOR U23350 ( .A(n131), .B(n70), .Z(n23020) );
  IV U23351 ( .A(n23020), .Z(n23019) );
  NOR U23352 ( .A(n23021), .B(n23019), .Z(n23367) );
  XOR U23353 ( .A(n23021), .B(n23020), .Z(n23478) );
  NOR U23354 ( .A(n128), .B(n70), .Z(n23361) );
  XOR U23355 ( .A(n23023), .B(n23022), .Z(n23360) );
  NOR U23356 ( .A(n23361), .B(n23360), .Z(n23364) );
  XOR U23357 ( .A(n23025), .B(n23024), .Z(n23356) );
  NOR U23358 ( .A(n126), .B(n70), .Z(n23355) );
  IV U23359 ( .A(n23355), .Z(n23026) );
  NOR U23360 ( .A(n23356), .B(n23026), .Z(n23358) );
  NOR U23361 ( .A(n125), .B(n70), .Z(n23350) );
  XOR U23362 ( .A(n23028), .B(n23027), .Z(n23349) );
  NOR U23363 ( .A(n23350), .B(n23349), .Z(n23353) );
  XOR U23364 ( .A(n23030), .B(n23029), .Z(n23345) );
  NOR U23365 ( .A(n123), .B(n70), .Z(n23344) );
  IV U23366 ( .A(n23344), .Z(n23031) );
  NOR U23367 ( .A(n23345), .B(n23031), .Z(n23347) );
  NOR U23368 ( .A(n120), .B(n70), .Z(n23339) );
  XOR U23369 ( .A(n23033), .B(n23032), .Z(n23338) );
  NOR U23370 ( .A(n23339), .B(n23338), .Z(n23342) );
  XOR U23371 ( .A(n23035), .B(n23034), .Z(n23334) );
  NOR U23372 ( .A(n119), .B(n70), .Z(n23333) );
  IV U23373 ( .A(n23333), .Z(n23036) );
  NOR U23374 ( .A(n23334), .B(n23036), .Z(n23336) );
  NOR U23375 ( .A(n79), .B(n70), .Z(n23328) );
  XOR U23376 ( .A(n23038), .B(n23037), .Z(n23327) );
  NOR U23377 ( .A(n23328), .B(n23327), .Z(n23331) );
  XOR U23378 ( .A(n23040), .B(n23039), .Z(n23323) );
  NOR U23379 ( .A(n117), .B(n70), .Z(n23322) );
  IV U23380 ( .A(n23322), .Z(n23041) );
  NOR U23381 ( .A(n23323), .B(n23041), .Z(n23325) );
  NOR U23382 ( .A(n80), .B(n70), .Z(n23045) );
  XOR U23383 ( .A(n23043), .B(n23042), .Z(n23044) );
  NOR U23384 ( .A(n23045), .B(n23044), .Z(n23320) );
  XOR U23385 ( .A(n23045), .B(n23044), .Z(n23046) );
  IV U23386 ( .A(n23046), .Z(n23503) );
  XOR U23387 ( .A(n23048), .B(n23047), .Z(n23315) );
  NOR U23388 ( .A(n116), .B(n70), .Z(n23314) );
  IV U23389 ( .A(n23314), .Z(n23049) );
  NOR U23390 ( .A(n23315), .B(n23049), .Z(n23317) );
  NOR U23391 ( .A(n81), .B(n70), .Z(n23309) );
  XOR U23392 ( .A(n23051), .B(n23050), .Z(n23308) );
  NOR U23393 ( .A(n23309), .B(n23308), .Z(n23312) );
  XOR U23394 ( .A(n23053), .B(n23052), .Z(n23304) );
  NOR U23395 ( .A(n115), .B(n70), .Z(n23303) );
  IV U23396 ( .A(n23303), .Z(n23054) );
  NOR U23397 ( .A(n23304), .B(n23054), .Z(n23306) );
  IV U23398 ( .A(n23055), .Z(n23057) );
  XOR U23399 ( .A(n23057), .B(n23056), .Z(n23299) );
  NOR U23400 ( .A(n82), .B(n70), .Z(n23300) );
  IV U23401 ( .A(n23300), .Z(n23058) );
  NOR U23402 ( .A(n23299), .B(n23058), .Z(n23302) );
  IV U23403 ( .A(n23059), .Z(n23061) );
  XOR U23404 ( .A(n23061), .B(n23060), .Z(n23295) );
  NOR U23405 ( .A(n114), .B(n70), .Z(n23296) );
  IV U23406 ( .A(n23296), .Z(n23062) );
  NOR U23407 ( .A(n23295), .B(n23062), .Z(n23298) );
  IV U23408 ( .A(n23063), .Z(n23065) );
  XOR U23409 ( .A(n23065), .B(n23064), .Z(n23291) );
  NOR U23410 ( .A(n83), .B(n70), .Z(n23292) );
  IV U23411 ( .A(n23292), .Z(n23066) );
  NOR U23412 ( .A(n23291), .B(n23066), .Z(n23294) );
  IV U23413 ( .A(n23067), .Z(n23069) );
  XOR U23414 ( .A(n23069), .B(n23068), .Z(n23287) );
  NOR U23415 ( .A(n113), .B(n70), .Z(n23288) );
  IV U23416 ( .A(n23288), .Z(n23070) );
  NOR U23417 ( .A(n23287), .B(n23070), .Z(n23290) );
  IV U23418 ( .A(n23071), .Z(n23073) );
  XOR U23419 ( .A(n23073), .B(n23072), .Z(n23283) );
  NOR U23420 ( .A(n84), .B(n70), .Z(n23284) );
  IV U23421 ( .A(n23284), .Z(n23074) );
  NOR U23422 ( .A(n23283), .B(n23074), .Z(n23286) );
  IV U23423 ( .A(n23075), .Z(n23077) );
  XOR U23424 ( .A(n23077), .B(n23076), .Z(n23279) );
  NOR U23425 ( .A(n112), .B(n70), .Z(n23280) );
  IV U23426 ( .A(n23280), .Z(n23078) );
  NOR U23427 ( .A(n23279), .B(n23078), .Z(n23282) );
  IV U23428 ( .A(n23079), .Z(n23081) );
  XOR U23429 ( .A(n23081), .B(n23080), .Z(n23275) );
  NOR U23430 ( .A(n85), .B(n70), .Z(n23276) );
  IV U23431 ( .A(n23276), .Z(n23082) );
  NOR U23432 ( .A(n23275), .B(n23082), .Z(n23278) );
  IV U23433 ( .A(n23083), .Z(n23085) );
  XOR U23434 ( .A(n23085), .B(n23084), .Z(n23271) );
  NOR U23435 ( .A(n111), .B(n70), .Z(n23272) );
  IV U23436 ( .A(n23272), .Z(n23086) );
  NOR U23437 ( .A(n23271), .B(n23086), .Z(n23274) );
  IV U23438 ( .A(n23087), .Z(n23089) );
  XOR U23439 ( .A(n23089), .B(n23088), .Z(n23267) );
  NOR U23440 ( .A(n86), .B(n70), .Z(n23268) );
  IV U23441 ( .A(n23268), .Z(n23090) );
  NOR U23442 ( .A(n23267), .B(n23090), .Z(n23270) );
  IV U23443 ( .A(n23091), .Z(n23093) );
  XOR U23444 ( .A(n23093), .B(n23092), .Z(n23263) );
  NOR U23445 ( .A(n110), .B(n70), .Z(n23264) );
  IV U23446 ( .A(n23264), .Z(n23094) );
  NOR U23447 ( .A(n23263), .B(n23094), .Z(n23266) );
  XOR U23448 ( .A(n23096), .B(n23095), .Z(n23259) );
  NOR U23449 ( .A(n109), .B(n70), .Z(n23260) );
  IV U23450 ( .A(n23260), .Z(n23097) );
  NOR U23451 ( .A(n23259), .B(n23097), .Z(n23262) );
  IV U23452 ( .A(n23098), .Z(n23100) );
  XOR U23453 ( .A(n23100), .B(n23099), .Z(n23255) );
  NOR U23454 ( .A(n108), .B(n70), .Z(n23256) );
  IV U23455 ( .A(n23256), .Z(n23101) );
  NOR U23456 ( .A(n23255), .B(n23101), .Z(n23258) );
  XOR U23457 ( .A(n23103), .B(n23102), .Z(n23251) );
  IV U23458 ( .A(n23251), .Z(n23105) );
  NOR U23459 ( .A(n87), .B(n70), .Z(n23104) );
  IV U23460 ( .A(n23104), .Z(n23252) );
  NOR U23461 ( .A(n23105), .B(n23252), .Z(n23254) );
  IV U23462 ( .A(n23106), .Z(n23108) );
  XOR U23463 ( .A(n23108), .B(n23107), .Z(n23247) );
  NOR U23464 ( .A(n107), .B(n70), .Z(n23248) );
  IV U23465 ( .A(n23248), .Z(n23109) );
  NOR U23466 ( .A(n23247), .B(n23109), .Z(n23250) );
  IV U23467 ( .A(n23110), .Z(n23112) );
  XOR U23468 ( .A(n23112), .B(n23111), .Z(n23243) );
  NOR U23469 ( .A(n88), .B(n70), .Z(n23244) );
  IV U23470 ( .A(n23244), .Z(n23113) );
  NOR U23471 ( .A(n23243), .B(n23113), .Z(n23246) );
  IV U23472 ( .A(n23114), .Z(n23116) );
  XOR U23473 ( .A(n23116), .B(n23115), .Z(n23239) );
  NOR U23474 ( .A(n106), .B(n70), .Z(n23240) );
  IV U23475 ( .A(n23240), .Z(n23117) );
  NOR U23476 ( .A(n23239), .B(n23117), .Z(n23242) );
  XOR U23477 ( .A(n23119), .B(n23118), .Z(n23235) );
  NOR U23478 ( .A(n105), .B(n70), .Z(n23236) );
  IV U23479 ( .A(n23236), .Z(n23120) );
  NOR U23480 ( .A(n23235), .B(n23120), .Z(n23238) );
  XOR U23481 ( .A(n23122), .B(n23121), .Z(n23223) );
  IV U23482 ( .A(n23223), .Z(n23124) );
  NOR U23483 ( .A(n89), .B(n70), .Z(n23123) );
  IV U23484 ( .A(n23123), .Z(n23224) );
  NOR U23485 ( .A(n23124), .B(n23224), .Z(n23226) );
  IV U23486 ( .A(n23125), .Z(n23127) );
  XOR U23487 ( .A(n23127), .B(n23126), .Z(n23219) );
  NOR U23488 ( .A(n103), .B(n70), .Z(n23220) );
  IV U23489 ( .A(n23220), .Z(n23128) );
  NOR U23490 ( .A(n23219), .B(n23128), .Z(n23222) );
  IV U23491 ( .A(n23129), .Z(n23131) );
  XOR U23492 ( .A(n23131), .B(n23130), .Z(n23215) );
  NOR U23493 ( .A(n90), .B(n70), .Z(n23216) );
  IV U23494 ( .A(n23216), .Z(n23132) );
  NOR U23495 ( .A(n23215), .B(n23132), .Z(n23218) );
  IV U23496 ( .A(n23133), .Z(n23135) );
  XOR U23497 ( .A(n23135), .B(n23134), .Z(n23211) );
  NOR U23498 ( .A(n102), .B(n70), .Z(n23212) );
  IV U23499 ( .A(n23212), .Z(n23136) );
  NOR U23500 ( .A(n23211), .B(n23136), .Z(n23214) );
  IV U23501 ( .A(n23137), .Z(n23139) );
  XOR U23502 ( .A(n23139), .B(n23138), .Z(n23207) );
  NOR U23503 ( .A(n101), .B(n70), .Z(n23208) );
  IV U23504 ( .A(n23208), .Z(n23140) );
  NOR U23505 ( .A(n23207), .B(n23140), .Z(n23210) );
  IV U23506 ( .A(n23141), .Z(n23143) );
  XOR U23507 ( .A(n23143), .B(n23142), .Z(n23203) );
  NOR U23508 ( .A(n100), .B(n70), .Z(n23204) );
  IV U23509 ( .A(n23204), .Z(n23144) );
  NOR U23510 ( .A(n23203), .B(n23144), .Z(n23206) );
  IV U23511 ( .A(n23145), .Z(n23147) );
  XOR U23512 ( .A(n23147), .B(n23146), .Z(n23199) );
  NOR U23513 ( .A(n99), .B(n70), .Z(n23200) );
  IV U23514 ( .A(n23200), .Z(n23148) );
  NOR U23515 ( .A(n23199), .B(n23148), .Z(n23202) );
  IV U23516 ( .A(n23149), .Z(n23151) );
  XOR U23517 ( .A(n23151), .B(n23150), .Z(n23195) );
  NOR U23518 ( .A(n98), .B(n70), .Z(n23196) );
  IV U23519 ( .A(n23196), .Z(n23152) );
  NOR U23520 ( .A(n23195), .B(n23152), .Z(n23198) );
  XOR U23521 ( .A(n23154), .B(n23153), .Z(n23191) );
  NOR U23522 ( .A(n91), .B(n70), .Z(n23192) );
  IV U23523 ( .A(n23192), .Z(n23155) );
  NOR U23524 ( .A(n23191), .B(n23155), .Z(n23194) );
  XOR U23525 ( .A(n23157), .B(n23156), .Z(n23179) );
  IV U23526 ( .A(n23179), .Z(n23159) );
  NOR U23527 ( .A(n96), .B(n70), .Z(n23158) );
  IV U23528 ( .A(n23158), .Z(n23180) );
  NOR U23529 ( .A(n23159), .B(n23180), .Z(n23182) );
  NOR U23530 ( .A(n95), .B(n70), .Z(n23176) );
  IV U23531 ( .A(n23176), .Z(n23162) );
  XOR U23532 ( .A(n23161), .B(n23160), .Z(n23175) );
  NOR U23533 ( .A(n23162), .B(n23175), .Z(n23178) );
  NOR U23534 ( .A(n93), .B(n70), .Z(n24181) );
  IV U23535 ( .A(n24181), .Z(n23163) );
  NOR U23536 ( .A(n69), .B(n168), .Z(n23171) );
  IV U23537 ( .A(n23171), .Z(n23166) );
  NOR U23538 ( .A(n23163), .B(n23166), .Z(n23164) );
  IV U23539 ( .A(n23164), .Z(n23165) );
  NOR U23540 ( .A(n94), .B(n23165), .Z(n23174) );
  NOR U23541 ( .A(n23166), .B(n93), .Z(n23167) );
  XOR U23542 ( .A(n94), .B(n23167), .Z(n23168) );
  NOR U23543 ( .A(n70), .B(n23168), .Z(n23169) );
  IV U23544 ( .A(n23169), .Z(n23619) );
  XOR U23545 ( .A(n23171), .B(n23170), .Z(n23618) );
  IV U23546 ( .A(n23618), .Z(n23172) );
  NOR U23547 ( .A(n23619), .B(n23172), .Z(n23173) );
  NOR U23548 ( .A(n23174), .B(n23173), .Z(n23615) );
  XOR U23549 ( .A(n23176), .B(n23175), .Z(n23614) );
  NOR U23550 ( .A(n23615), .B(n23614), .Z(n23177) );
  NOR U23551 ( .A(n23178), .B(n23177), .Z(n23642) );
  XOR U23552 ( .A(n23180), .B(n23179), .Z(n23641) );
  NOR U23553 ( .A(n23642), .B(n23641), .Z(n23181) );
  NOR U23554 ( .A(n23182), .B(n23181), .Z(n23187) );
  XOR U23555 ( .A(n23184), .B(n23183), .Z(n23186) );
  IV U23556 ( .A(n23186), .Z(n23185) );
  NOR U23557 ( .A(n23187), .B(n23185), .Z(n23190) );
  XOR U23558 ( .A(n23187), .B(n23186), .Z(n23611) );
  NOR U23559 ( .A(n97), .B(n70), .Z(n23612) );
  IV U23560 ( .A(n23612), .Z(n23188) );
  NOR U23561 ( .A(n23611), .B(n23188), .Z(n23189) );
  NOR U23562 ( .A(n23190), .B(n23189), .Z(n23607) );
  XOR U23563 ( .A(n23192), .B(n23191), .Z(n23608) );
  NOR U23564 ( .A(n23607), .B(n23608), .Z(n23193) );
  NOR U23565 ( .A(n23194), .B(n23193), .Z(n23603) );
  XOR U23566 ( .A(n23196), .B(n23195), .Z(n23604) );
  NOR U23567 ( .A(n23603), .B(n23604), .Z(n23197) );
  NOR U23568 ( .A(n23198), .B(n23197), .Z(n23599) );
  XOR U23569 ( .A(n23200), .B(n23199), .Z(n23600) );
  NOR U23570 ( .A(n23599), .B(n23600), .Z(n23201) );
  NOR U23571 ( .A(n23202), .B(n23201), .Z(n23595) );
  XOR U23572 ( .A(n23204), .B(n23203), .Z(n23596) );
  NOR U23573 ( .A(n23595), .B(n23596), .Z(n23205) );
  NOR U23574 ( .A(n23206), .B(n23205), .Z(n23591) );
  XOR U23575 ( .A(n23208), .B(n23207), .Z(n23592) );
  NOR U23576 ( .A(n23591), .B(n23592), .Z(n23209) );
  NOR U23577 ( .A(n23210), .B(n23209), .Z(n23587) );
  XOR U23578 ( .A(n23212), .B(n23211), .Z(n23588) );
  NOR U23579 ( .A(n23587), .B(n23588), .Z(n23213) );
  NOR U23580 ( .A(n23214), .B(n23213), .Z(n23583) );
  XOR U23581 ( .A(n23216), .B(n23215), .Z(n23584) );
  NOR U23582 ( .A(n23583), .B(n23584), .Z(n23217) );
  NOR U23583 ( .A(n23218), .B(n23217), .Z(n23579) );
  XOR U23584 ( .A(n23220), .B(n23219), .Z(n23580) );
  NOR U23585 ( .A(n23579), .B(n23580), .Z(n23221) );
  NOR U23586 ( .A(n23222), .B(n23221), .Z(n23686) );
  XOR U23587 ( .A(n23224), .B(n23223), .Z(n23685) );
  NOR U23588 ( .A(n23686), .B(n23685), .Z(n23225) );
  NOR U23589 ( .A(n23226), .B(n23225), .Z(n23231) );
  XOR U23590 ( .A(n23228), .B(n23227), .Z(n23230) );
  IV U23591 ( .A(n23230), .Z(n23229) );
  NOR U23592 ( .A(n23231), .B(n23229), .Z(n23234) );
  XOR U23593 ( .A(n23231), .B(n23230), .Z(n23576) );
  NOR U23594 ( .A(n104), .B(n70), .Z(n23577) );
  IV U23595 ( .A(n23577), .Z(n23232) );
  NOR U23596 ( .A(n23576), .B(n23232), .Z(n23233) );
  NOR U23597 ( .A(n23234), .B(n23233), .Z(n23572) );
  XOR U23598 ( .A(n23236), .B(n23235), .Z(n23573) );
  NOR U23599 ( .A(n23572), .B(n23573), .Z(n23237) );
  NOR U23600 ( .A(n23238), .B(n23237), .Z(n23568) );
  XOR U23601 ( .A(n23240), .B(n23239), .Z(n23569) );
  NOR U23602 ( .A(n23568), .B(n23569), .Z(n23241) );
  NOR U23603 ( .A(n23242), .B(n23241), .Z(n23564) );
  XOR U23604 ( .A(n23244), .B(n23243), .Z(n23565) );
  NOR U23605 ( .A(n23564), .B(n23565), .Z(n23245) );
  NOR U23606 ( .A(n23246), .B(n23245), .Z(n23561) );
  XOR U23607 ( .A(n23248), .B(n23247), .Z(n23560) );
  NOR U23608 ( .A(n23561), .B(n23560), .Z(n23249) );
  NOR U23609 ( .A(n23250), .B(n23249), .Z(n23714) );
  XOR U23610 ( .A(n23252), .B(n23251), .Z(n23713) );
  NOR U23611 ( .A(n23714), .B(n23713), .Z(n23253) );
  NOR U23612 ( .A(n23254), .B(n23253), .Z(n23556) );
  XOR U23613 ( .A(n23256), .B(n23255), .Z(n23557) );
  NOR U23614 ( .A(n23556), .B(n23557), .Z(n23257) );
  NOR U23615 ( .A(n23258), .B(n23257), .Z(n23552) );
  XOR U23616 ( .A(n23260), .B(n23259), .Z(n23553) );
  NOR U23617 ( .A(n23552), .B(n23553), .Z(n23261) );
  NOR U23618 ( .A(n23262), .B(n23261), .Z(n23548) );
  XOR U23619 ( .A(n23264), .B(n23263), .Z(n23549) );
  NOR U23620 ( .A(n23548), .B(n23549), .Z(n23265) );
  NOR U23621 ( .A(n23266), .B(n23265), .Z(n23544) );
  XOR U23622 ( .A(n23268), .B(n23267), .Z(n23545) );
  NOR U23623 ( .A(n23544), .B(n23545), .Z(n23269) );
  NOR U23624 ( .A(n23270), .B(n23269), .Z(n23540) );
  XOR U23625 ( .A(n23272), .B(n23271), .Z(n23541) );
  NOR U23626 ( .A(n23540), .B(n23541), .Z(n23273) );
  NOR U23627 ( .A(n23274), .B(n23273), .Z(n23536) );
  XOR U23628 ( .A(n23276), .B(n23275), .Z(n23537) );
  NOR U23629 ( .A(n23536), .B(n23537), .Z(n23277) );
  NOR U23630 ( .A(n23278), .B(n23277), .Z(n23532) );
  XOR U23631 ( .A(n23280), .B(n23279), .Z(n23533) );
  NOR U23632 ( .A(n23532), .B(n23533), .Z(n23281) );
  NOR U23633 ( .A(n23282), .B(n23281), .Z(n23528) );
  XOR U23634 ( .A(n23284), .B(n23283), .Z(n23529) );
  NOR U23635 ( .A(n23528), .B(n23529), .Z(n23285) );
  NOR U23636 ( .A(n23286), .B(n23285), .Z(n23524) );
  XOR U23637 ( .A(n23288), .B(n23287), .Z(n23525) );
  NOR U23638 ( .A(n23524), .B(n23525), .Z(n23289) );
  NOR U23639 ( .A(n23290), .B(n23289), .Z(n23520) );
  XOR U23640 ( .A(n23292), .B(n23291), .Z(n23521) );
  NOR U23641 ( .A(n23520), .B(n23521), .Z(n23293) );
  NOR U23642 ( .A(n23294), .B(n23293), .Z(n23516) );
  XOR U23643 ( .A(n23296), .B(n23295), .Z(n23517) );
  NOR U23644 ( .A(n23516), .B(n23517), .Z(n23297) );
  NOR U23645 ( .A(n23298), .B(n23297), .Z(n23512) );
  XOR U23646 ( .A(n23300), .B(n23299), .Z(n23513) );
  NOR U23647 ( .A(n23512), .B(n23513), .Z(n23301) );
  NOR U23648 ( .A(n23302), .B(n23301), .Z(n23511) );
  XOR U23649 ( .A(n23304), .B(n23303), .Z(n23510) );
  NOR U23650 ( .A(n23511), .B(n23510), .Z(n23305) );
  NOR U23651 ( .A(n23306), .B(n23305), .Z(n23307) );
  IV U23652 ( .A(n23307), .Z(n23508) );
  XOR U23653 ( .A(n23309), .B(n23308), .Z(n23310) );
  IV U23654 ( .A(n23310), .Z(n23507) );
  NOR U23655 ( .A(n23508), .B(n23507), .Z(n23311) );
  NOR U23656 ( .A(n23312), .B(n23311), .Z(n23313) );
  IV U23657 ( .A(n23313), .Z(n23506) );
  XOR U23658 ( .A(n23315), .B(n23314), .Z(n23505) );
  NOR U23659 ( .A(n23506), .B(n23505), .Z(n23316) );
  NOR U23660 ( .A(n23317), .B(n23316), .Z(n23318) );
  IV U23661 ( .A(n23318), .Z(n23502) );
  NOR U23662 ( .A(n23503), .B(n23502), .Z(n23319) );
  NOR U23663 ( .A(n23320), .B(n23319), .Z(n23321) );
  IV U23664 ( .A(n23321), .Z(n23501) );
  XOR U23665 ( .A(n23323), .B(n23322), .Z(n23500) );
  NOR U23666 ( .A(n23501), .B(n23500), .Z(n23324) );
  NOR U23667 ( .A(n23325), .B(n23324), .Z(n23326) );
  IV U23668 ( .A(n23326), .Z(n23498) );
  XOR U23669 ( .A(n23328), .B(n23327), .Z(n23329) );
  IV U23670 ( .A(n23329), .Z(n23497) );
  NOR U23671 ( .A(n23498), .B(n23497), .Z(n23330) );
  NOR U23672 ( .A(n23331), .B(n23330), .Z(n23332) );
  IV U23673 ( .A(n23332), .Z(n23496) );
  XOR U23674 ( .A(n23334), .B(n23333), .Z(n23495) );
  NOR U23675 ( .A(n23496), .B(n23495), .Z(n23335) );
  NOR U23676 ( .A(n23336), .B(n23335), .Z(n23337) );
  IV U23677 ( .A(n23337), .Z(n23493) );
  XOR U23678 ( .A(n23339), .B(n23338), .Z(n23340) );
  IV U23679 ( .A(n23340), .Z(n23492) );
  NOR U23680 ( .A(n23493), .B(n23492), .Z(n23341) );
  NOR U23681 ( .A(n23342), .B(n23341), .Z(n23343) );
  IV U23682 ( .A(n23343), .Z(n23491) );
  XOR U23683 ( .A(n23345), .B(n23344), .Z(n23490) );
  NOR U23684 ( .A(n23491), .B(n23490), .Z(n23346) );
  NOR U23685 ( .A(n23347), .B(n23346), .Z(n23348) );
  IV U23686 ( .A(n23348), .Z(n23488) );
  XOR U23687 ( .A(n23350), .B(n23349), .Z(n23351) );
  IV U23688 ( .A(n23351), .Z(n23487) );
  NOR U23689 ( .A(n23488), .B(n23487), .Z(n23352) );
  NOR U23690 ( .A(n23353), .B(n23352), .Z(n23354) );
  IV U23691 ( .A(n23354), .Z(n23486) );
  XOR U23692 ( .A(n23356), .B(n23355), .Z(n23485) );
  NOR U23693 ( .A(n23486), .B(n23485), .Z(n23357) );
  NOR U23694 ( .A(n23358), .B(n23357), .Z(n23359) );
  IV U23695 ( .A(n23359), .Z(n23483) );
  XOR U23696 ( .A(n23361), .B(n23360), .Z(n23362) );
  IV U23697 ( .A(n23362), .Z(n23482) );
  NOR U23698 ( .A(n23483), .B(n23482), .Z(n23363) );
  NOR U23699 ( .A(n23364), .B(n23363), .Z(n23365) );
  IV U23700 ( .A(n23365), .Z(n23477) );
  NOR U23701 ( .A(n23478), .B(n23477), .Z(n23366) );
  NOR U23702 ( .A(n23367), .B(n23366), .Z(n23368) );
  IV U23703 ( .A(n23368), .Z(n23474) );
  NOR U23704 ( .A(n23475), .B(n23474), .Z(n23369) );
  NOR U23705 ( .A(n23370), .B(n23369), .Z(n23472) );
  IV U23706 ( .A(n23472), .Z(n23373) );
  XOR U23707 ( .A(n23372), .B(n23371), .Z(n23471) );
  NOR U23708 ( .A(n23373), .B(n23471), .Z(n23374) );
  NOR U23709 ( .A(n23375), .B(n23374), .Z(n23468) );
  XOR U23710 ( .A(n23377), .B(n23376), .Z(n23467) );
  NOR U23711 ( .A(n23468), .B(n23467), .Z(n23378) );
  NOR U23712 ( .A(n23379), .B(n23378), .Z(n23464) );
  XOR U23713 ( .A(n23381), .B(n23380), .Z(n23463) );
  NOR U23714 ( .A(n23464), .B(n23463), .Z(n23382) );
  NOR U23715 ( .A(n23383), .B(n23382), .Z(n23384) );
  IV U23716 ( .A(n23384), .Z(n23857) );
  XOR U23717 ( .A(n23386), .B(n23385), .Z(n23387) );
  IV U23718 ( .A(n23387), .Z(n23856) );
  NOR U23719 ( .A(n23857), .B(n23856), .Z(n23388) );
  NOR U23720 ( .A(n23389), .B(n23388), .Z(n23461) );
  IV U23721 ( .A(n23461), .Z(n23390) );
  NOR U23722 ( .A(n23460), .B(n23390), .Z(n23391) );
  NOR U23723 ( .A(n23392), .B(n23391), .Z(n23458) );
  NOR U23724 ( .A(n23393), .B(n23458), .Z(n23394) );
  NOR U23725 ( .A(n23395), .B(n23394), .Z(n23401) );
  XOR U23726 ( .A(n23397), .B(n23396), .Z(n23398) );
  XOR U23727 ( .A(n23399), .B(n23398), .Z(n23400) );
  NOR U23728 ( .A(n23401), .B(n23400), .Z(n23405) );
  NOR U23729 ( .A(n147), .B(n70), .Z(n23454) );
  IV U23730 ( .A(n23454), .Z(n23403) );
  XOR U23731 ( .A(n23401), .B(n23400), .Z(n23402) );
  IV U23732 ( .A(n23402), .Z(n23453) );
  NOR U23733 ( .A(n23403), .B(n23453), .Z(n23404) );
  NOR U23734 ( .A(n23405), .B(n23404), .Z(n23406) );
  IV U23735 ( .A(n23406), .Z(n23872) );
  NOR U23736 ( .A(n23873), .B(n23872), .Z(n23407) );
  NOR U23737 ( .A(n23408), .B(n23407), .Z(n23414) );
  IV U23738 ( .A(n23414), .Z(n23412) );
  IV U23739 ( .A(n23409), .Z(n23411) );
  XOR U23740 ( .A(n23411), .B(n23410), .Z(n23413) );
  NOR U23741 ( .A(n23412), .B(n23413), .Z(n23417) );
  XOR U23742 ( .A(n23414), .B(n23413), .Z(n23879) );
  NOR U23743 ( .A(n150), .B(n70), .Z(n23880) );
  IV U23744 ( .A(n23880), .Z(n23415) );
  NOR U23745 ( .A(n23879), .B(n23415), .Z(n23416) );
  NOR U23746 ( .A(n23417), .B(n23416), .Z(n23420) );
  NOR U23747 ( .A(n153), .B(n70), .Z(n23419) );
  IV U23748 ( .A(n23419), .Z(n23418) );
  NOR U23749 ( .A(n23420), .B(n23418), .Z(n23425) );
  XOR U23750 ( .A(n23420), .B(n23419), .Z(n23886) );
  XOR U23751 ( .A(n23422), .B(n23421), .Z(n23887) );
  IV U23752 ( .A(n23887), .Z(n23423) );
  NOR U23753 ( .A(n23886), .B(n23423), .Z(n23424) );
  NOR U23754 ( .A(n23425), .B(n23424), .Z(n23428) );
  NOR U23755 ( .A(n155), .B(n70), .Z(n23427) );
  IV U23756 ( .A(n23427), .Z(n23426) );
  NOR U23757 ( .A(n23428), .B(n23426), .Z(n23433) );
  XOR U23758 ( .A(n23428), .B(n23427), .Z(n23892) );
  XOR U23759 ( .A(n23430), .B(n23429), .Z(n23893) );
  IV U23760 ( .A(n23893), .Z(n23431) );
  NOR U23761 ( .A(n23892), .B(n23431), .Z(n23432) );
  NOR U23762 ( .A(n23433), .B(n23432), .Z(n23438) );
  NOR U23763 ( .A(n156), .B(n70), .Z(n23437) );
  IV U23764 ( .A(n23437), .Z(n23434) );
  NOR U23765 ( .A(n23438), .B(n23434), .Z(n23440) );
  XOR U23766 ( .A(n23436), .B(n23435), .Z(n23904) );
  XOR U23767 ( .A(n23438), .B(n23437), .Z(n23903) );
  NOR U23768 ( .A(n23904), .B(n23903), .Z(n23439) );
  NOR U23769 ( .A(n23440), .B(n23439), .Z(n23444) );
  IV U23770 ( .A(n23444), .Z(n23441) );
  NOR U23771 ( .A(n23445), .B(n23441), .Z(n23447) );
  XOR U23772 ( .A(n23443), .B(n23442), .Z(n23910) );
  XOR U23773 ( .A(n23445), .B(n23444), .Z(n23909) );
  NOR U23774 ( .A(n23910), .B(n23909), .Z(n23446) );
  NOR U23775 ( .A(n23447), .B(n23446), .Z(n23922) );
  NOR U23776 ( .A(n161), .B(n70), .Z(n23448) );
  IV U23777 ( .A(n23448), .Z(n23923) );
  XOR U23778 ( .A(n23922), .B(n23923), .Z(n23926) );
  XOR U23779 ( .A(n23450), .B(n23449), .Z(n23925) );
  XOR U23780 ( .A(n23926), .B(n23925), .Z(n23451) );
  IV U23781 ( .A(n23451), .Z(n23915) );
  NOR U23782 ( .A(n163), .B(n71), .Z(n23916) );
  IV U23783 ( .A(n23916), .Z(n23452) );
  NOR U23784 ( .A(n23915), .B(n23452), .Z(n23918) );
  XOR U23785 ( .A(n23454), .B(n23453), .Z(n23989) );
  NOR U23786 ( .A(n148), .B(n71), .Z(n23992) );
  XOR U23787 ( .A(n23456), .B(n23455), .Z(n23457) );
  XOR U23788 ( .A(n23458), .B(n23457), .Z(n23867) );
  NOR U23789 ( .A(n147), .B(n71), .Z(n23866) );
  IV U23790 ( .A(n23866), .Z(n23459) );
  NOR U23791 ( .A(n23867), .B(n23459), .Z(n23869) );
  XOR U23792 ( .A(n23461), .B(n23460), .Z(n23862) );
  NOR U23793 ( .A(n145), .B(n71), .Z(n23863) );
  IV U23794 ( .A(n23863), .Z(n23462) );
  NOR U23795 ( .A(n23862), .B(n23462), .Z(n23865) );
  NOR U23796 ( .A(n143), .B(n71), .Z(n23859) );
  IV U23797 ( .A(n23859), .Z(n23855) );
  NOR U23798 ( .A(n141), .B(n71), .Z(n24003) );
  XOR U23799 ( .A(n23464), .B(n23463), .Z(n23465) );
  NOR U23800 ( .A(n24003), .B(n23465), .Z(n23853) );
  IV U23801 ( .A(n24003), .Z(n23466) );
  IV U23802 ( .A(n23465), .Z(n24005) );
  NOR U23803 ( .A(n23466), .B(n24005), .Z(n23851) );
  NOR U23804 ( .A(n139), .B(n71), .Z(n23469) );
  XOR U23805 ( .A(n23468), .B(n23467), .Z(n24010) );
  NOR U23806 ( .A(n23469), .B(n24010), .Z(n23850) );
  IV U23807 ( .A(n23469), .Z(n24007) );
  IV U23808 ( .A(n24010), .Z(n23470) );
  NOR U23809 ( .A(n24007), .B(n23470), .Z(n23848) );
  XOR U23810 ( .A(n23472), .B(n23471), .Z(n23843) );
  NOR U23811 ( .A(n137), .B(n71), .Z(n23844) );
  IV U23812 ( .A(n23844), .Z(n23473) );
  NOR U23813 ( .A(n23843), .B(n23473), .Z(n23846) );
  XOR U23814 ( .A(n23475), .B(n23474), .Z(n23839) );
  NOR U23815 ( .A(n135), .B(n71), .Z(n23838) );
  IV U23816 ( .A(n23838), .Z(n23476) );
  NOR U23817 ( .A(n23839), .B(n23476), .Z(n23842) );
  NOR U23818 ( .A(n133), .B(n71), .Z(n23480) );
  XOR U23819 ( .A(n23478), .B(n23477), .Z(n23479) );
  NOR U23820 ( .A(n23480), .B(n23479), .Z(n23837) );
  XOR U23821 ( .A(n23480), .B(n23479), .Z(n23481) );
  IV U23822 ( .A(n23481), .Z(n24020) );
  XOR U23823 ( .A(n23483), .B(n23482), .Z(n23832) );
  NOR U23824 ( .A(n131), .B(n71), .Z(n23831) );
  IV U23825 ( .A(n23831), .Z(n23484) );
  NOR U23826 ( .A(n23832), .B(n23484), .Z(n23834) );
  NOR U23827 ( .A(n128), .B(n71), .Z(n23826) );
  XOR U23828 ( .A(n23486), .B(n23485), .Z(n23825) );
  NOR U23829 ( .A(n23826), .B(n23825), .Z(n23829) );
  XOR U23830 ( .A(n23488), .B(n23487), .Z(n23821) );
  NOR U23831 ( .A(n126), .B(n71), .Z(n23820) );
  IV U23832 ( .A(n23820), .Z(n23489) );
  NOR U23833 ( .A(n23821), .B(n23489), .Z(n23823) );
  NOR U23834 ( .A(n125), .B(n71), .Z(n23815) );
  XOR U23835 ( .A(n23491), .B(n23490), .Z(n23814) );
  NOR U23836 ( .A(n23815), .B(n23814), .Z(n23818) );
  XOR U23837 ( .A(n23493), .B(n23492), .Z(n23810) );
  NOR U23838 ( .A(n123), .B(n71), .Z(n23809) );
  IV U23839 ( .A(n23809), .Z(n23494) );
  NOR U23840 ( .A(n23810), .B(n23494), .Z(n23812) );
  NOR U23841 ( .A(n120), .B(n71), .Z(n23804) );
  XOR U23842 ( .A(n23496), .B(n23495), .Z(n23803) );
  NOR U23843 ( .A(n23804), .B(n23803), .Z(n23807) );
  XOR U23844 ( .A(n23498), .B(n23497), .Z(n23799) );
  NOR U23845 ( .A(n119), .B(n71), .Z(n23798) );
  IV U23846 ( .A(n23798), .Z(n23499) );
  NOR U23847 ( .A(n23799), .B(n23499), .Z(n23801) );
  NOR U23848 ( .A(n79), .B(n71), .Z(n23793) );
  XOR U23849 ( .A(n23501), .B(n23500), .Z(n23792) );
  NOR U23850 ( .A(n23793), .B(n23792), .Z(n23796) );
  XOR U23851 ( .A(n23503), .B(n23502), .Z(n23788) );
  NOR U23852 ( .A(n117), .B(n71), .Z(n23787) );
  IV U23853 ( .A(n23787), .Z(n23504) );
  NOR U23854 ( .A(n23788), .B(n23504), .Z(n23790) );
  NOR U23855 ( .A(n80), .B(n71), .Z(n23782) );
  XOR U23856 ( .A(n23506), .B(n23505), .Z(n23781) );
  NOR U23857 ( .A(n23782), .B(n23781), .Z(n23785) );
  XOR U23858 ( .A(n23508), .B(n23507), .Z(n23777) );
  NOR U23859 ( .A(n116), .B(n71), .Z(n23776) );
  IV U23860 ( .A(n23776), .Z(n23509) );
  NOR U23861 ( .A(n23777), .B(n23509), .Z(n23779) );
  NOR U23862 ( .A(n81), .B(n71), .Z(n23771) );
  XOR U23863 ( .A(n23511), .B(n23510), .Z(n23770) );
  NOR U23864 ( .A(n23771), .B(n23770), .Z(n23774) );
  IV U23865 ( .A(n23512), .Z(n23514) );
  XOR U23866 ( .A(n23514), .B(n23513), .Z(n23765) );
  NOR U23867 ( .A(n115), .B(n71), .Z(n23766) );
  IV U23868 ( .A(n23766), .Z(n23515) );
  NOR U23869 ( .A(n23765), .B(n23515), .Z(n23768) );
  IV U23870 ( .A(n23516), .Z(n23518) );
  XOR U23871 ( .A(n23518), .B(n23517), .Z(n23761) );
  NOR U23872 ( .A(n82), .B(n71), .Z(n23762) );
  IV U23873 ( .A(n23762), .Z(n23519) );
  NOR U23874 ( .A(n23761), .B(n23519), .Z(n23764) );
  IV U23875 ( .A(n23520), .Z(n23522) );
  XOR U23876 ( .A(n23522), .B(n23521), .Z(n23757) );
  NOR U23877 ( .A(n114), .B(n71), .Z(n23758) );
  IV U23878 ( .A(n23758), .Z(n23523) );
  NOR U23879 ( .A(n23757), .B(n23523), .Z(n23760) );
  IV U23880 ( .A(n23524), .Z(n23526) );
  XOR U23881 ( .A(n23526), .B(n23525), .Z(n23753) );
  NOR U23882 ( .A(n83), .B(n71), .Z(n23754) );
  IV U23883 ( .A(n23754), .Z(n23527) );
  NOR U23884 ( .A(n23753), .B(n23527), .Z(n23756) );
  IV U23885 ( .A(n23528), .Z(n23530) );
  XOR U23886 ( .A(n23530), .B(n23529), .Z(n23749) );
  NOR U23887 ( .A(n113), .B(n71), .Z(n23750) );
  IV U23888 ( .A(n23750), .Z(n23531) );
  NOR U23889 ( .A(n23749), .B(n23531), .Z(n23752) );
  IV U23890 ( .A(n23532), .Z(n23534) );
  XOR U23891 ( .A(n23534), .B(n23533), .Z(n23745) );
  NOR U23892 ( .A(n84), .B(n71), .Z(n23746) );
  IV U23893 ( .A(n23746), .Z(n23535) );
  NOR U23894 ( .A(n23745), .B(n23535), .Z(n23748) );
  IV U23895 ( .A(n23536), .Z(n23538) );
  XOR U23896 ( .A(n23538), .B(n23537), .Z(n23741) );
  NOR U23897 ( .A(n112), .B(n71), .Z(n23742) );
  IV U23898 ( .A(n23742), .Z(n23539) );
  NOR U23899 ( .A(n23741), .B(n23539), .Z(n23744) );
  IV U23900 ( .A(n23540), .Z(n23542) );
  XOR U23901 ( .A(n23542), .B(n23541), .Z(n23737) );
  NOR U23902 ( .A(n85), .B(n71), .Z(n23738) );
  IV U23903 ( .A(n23738), .Z(n23543) );
  NOR U23904 ( .A(n23737), .B(n23543), .Z(n23740) );
  IV U23905 ( .A(n23544), .Z(n23546) );
  XOR U23906 ( .A(n23546), .B(n23545), .Z(n23733) );
  NOR U23907 ( .A(n111), .B(n71), .Z(n23734) );
  IV U23908 ( .A(n23734), .Z(n23547) );
  NOR U23909 ( .A(n23733), .B(n23547), .Z(n23736) );
  IV U23910 ( .A(n23548), .Z(n23550) );
  XOR U23911 ( .A(n23550), .B(n23549), .Z(n23729) );
  NOR U23912 ( .A(n86), .B(n71), .Z(n23730) );
  IV U23913 ( .A(n23730), .Z(n23551) );
  NOR U23914 ( .A(n23729), .B(n23551), .Z(n23732) );
  IV U23915 ( .A(n23552), .Z(n23554) );
  XOR U23916 ( .A(n23554), .B(n23553), .Z(n23725) );
  NOR U23917 ( .A(n110), .B(n71), .Z(n23726) );
  IV U23918 ( .A(n23726), .Z(n23555) );
  NOR U23919 ( .A(n23725), .B(n23555), .Z(n23728) );
  IV U23920 ( .A(n23556), .Z(n23558) );
  XOR U23921 ( .A(n23558), .B(n23557), .Z(n23721) );
  NOR U23922 ( .A(n109), .B(n71), .Z(n23722) );
  IV U23923 ( .A(n23722), .Z(n23559) );
  NOR U23924 ( .A(n23721), .B(n23559), .Z(n23724) );
  XOR U23925 ( .A(n23561), .B(n23560), .Z(n23709) );
  IV U23926 ( .A(n23709), .Z(n23563) );
  NOR U23927 ( .A(n87), .B(n71), .Z(n23562) );
  IV U23928 ( .A(n23562), .Z(n23710) );
  NOR U23929 ( .A(n23563), .B(n23710), .Z(n23712) );
  IV U23930 ( .A(n23564), .Z(n23566) );
  XOR U23931 ( .A(n23566), .B(n23565), .Z(n23705) );
  NOR U23932 ( .A(n107), .B(n71), .Z(n23706) );
  IV U23933 ( .A(n23706), .Z(n23567) );
  NOR U23934 ( .A(n23705), .B(n23567), .Z(n23708) );
  IV U23935 ( .A(n23568), .Z(n23570) );
  XOR U23936 ( .A(n23570), .B(n23569), .Z(n23701) );
  NOR U23937 ( .A(n88), .B(n71), .Z(n23702) );
  IV U23938 ( .A(n23702), .Z(n23571) );
  NOR U23939 ( .A(n23701), .B(n23571), .Z(n23704) );
  IV U23940 ( .A(n23572), .Z(n23574) );
  XOR U23941 ( .A(n23574), .B(n23573), .Z(n23697) );
  NOR U23942 ( .A(n106), .B(n71), .Z(n23698) );
  IV U23943 ( .A(n23698), .Z(n23575) );
  NOR U23944 ( .A(n23697), .B(n23575), .Z(n23700) );
  XOR U23945 ( .A(n23577), .B(n23576), .Z(n23693) );
  NOR U23946 ( .A(n105), .B(n71), .Z(n23694) );
  IV U23947 ( .A(n23694), .Z(n23578) );
  NOR U23948 ( .A(n23693), .B(n23578), .Z(n23696) );
  IV U23949 ( .A(n23579), .Z(n23581) );
  XOR U23950 ( .A(n23581), .B(n23580), .Z(n23681) );
  NOR U23951 ( .A(n89), .B(n71), .Z(n23682) );
  IV U23952 ( .A(n23682), .Z(n23582) );
  NOR U23953 ( .A(n23681), .B(n23582), .Z(n23684) );
  IV U23954 ( .A(n23583), .Z(n23585) );
  XOR U23955 ( .A(n23585), .B(n23584), .Z(n23677) );
  NOR U23956 ( .A(n103), .B(n71), .Z(n23678) );
  IV U23957 ( .A(n23678), .Z(n23586) );
  NOR U23958 ( .A(n23677), .B(n23586), .Z(n23680) );
  IV U23959 ( .A(n23587), .Z(n23589) );
  XOR U23960 ( .A(n23589), .B(n23588), .Z(n23673) );
  NOR U23961 ( .A(n90), .B(n71), .Z(n23674) );
  IV U23962 ( .A(n23674), .Z(n23590) );
  NOR U23963 ( .A(n23673), .B(n23590), .Z(n23676) );
  IV U23964 ( .A(n23591), .Z(n23593) );
  XOR U23965 ( .A(n23593), .B(n23592), .Z(n23669) );
  NOR U23966 ( .A(n102), .B(n71), .Z(n23670) );
  IV U23967 ( .A(n23670), .Z(n23594) );
  NOR U23968 ( .A(n23669), .B(n23594), .Z(n23672) );
  IV U23969 ( .A(n23595), .Z(n23597) );
  XOR U23970 ( .A(n23597), .B(n23596), .Z(n23665) );
  NOR U23971 ( .A(n101), .B(n71), .Z(n23666) );
  IV U23972 ( .A(n23666), .Z(n23598) );
  NOR U23973 ( .A(n23665), .B(n23598), .Z(n23668) );
  IV U23974 ( .A(n23599), .Z(n23601) );
  XOR U23975 ( .A(n23601), .B(n23600), .Z(n23661) );
  NOR U23976 ( .A(n100), .B(n71), .Z(n23662) );
  IV U23977 ( .A(n23662), .Z(n23602) );
  NOR U23978 ( .A(n23661), .B(n23602), .Z(n23664) );
  IV U23979 ( .A(n23603), .Z(n23605) );
  XOR U23980 ( .A(n23605), .B(n23604), .Z(n23657) );
  NOR U23981 ( .A(n99), .B(n71), .Z(n23658) );
  IV U23982 ( .A(n23658), .Z(n23606) );
  NOR U23983 ( .A(n23657), .B(n23606), .Z(n23660) );
  IV U23984 ( .A(n23607), .Z(n23609) );
  XOR U23985 ( .A(n23609), .B(n23608), .Z(n23653) );
  NOR U23986 ( .A(n98), .B(n71), .Z(n23654) );
  IV U23987 ( .A(n23654), .Z(n23610) );
  NOR U23988 ( .A(n23653), .B(n23610), .Z(n23656) );
  XOR U23989 ( .A(n23612), .B(n23611), .Z(n23649) );
  NOR U23990 ( .A(n91), .B(n71), .Z(n23650) );
  IV U23991 ( .A(n23650), .Z(n23613) );
  NOR U23992 ( .A(n23649), .B(n23613), .Z(n23652) );
  XOR U23993 ( .A(n23615), .B(n23614), .Z(n23637) );
  IV U23994 ( .A(n23637), .Z(n23617) );
  NOR U23995 ( .A(n96), .B(n71), .Z(n23616) );
  IV U23996 ( .A(n23616), .Z(n23638) );
  NOR U23997 ( .A(n23617), .B(n23638), .Z(n23640) );
  NOR U23998 ( .A(n95), .B(n71), .Z(n23634) );
  IV U23999 ( .A(n23634), .Z(n23620) );
  XOR U24000 ( .A(n23619), .B(n23618), .Z(n23633) );
  NOR U24001 ( .A(n23620), .B(n23633), .Z(n23636) );
  NOR U24002 ( .A(n93), .B(n71), .Z(n24675) );
  IV U24003 ( .A(n24675), .Z(n23621) );
  NOR U24004 ( .A(n70), .B(n168), .Z(n23629) );
  IV U24005 ( .A(n23629), .Z(n23624) );
  NOR U24006 ( .A(n23621), .B(n23624), .Z(n23622) );
  IV U24007 ( .A(n23622), .Z(n23623) );
  NOR U24008 ( .A(n94), .B(n23623), .Z(n23632) );
  NOR U24009 ( .A(n23624), .B(n93), .Z(n23625) );
  XOR U24010 ( .A(n94), .B(n23625), .Z(n23626) );
  NOR U24011 ( .A(n71), .B(n23626), .Z(n23627) );
  IV U24012 ( .A(n23627), .Z(n24172) );
  XOR U24013 ( .A(n23629), .B(n23628), .Z(n24171) );
  IV U24014 ( .A(n24171), .Z(n23630) );
  NOR U24015 ( .A(n24172), .B(n23630), .Z(n23631) );
  NOR U24016 ( .A(n23632), .B(n23631), .Z(n24168) );
  XOR U24017 ( .A(n23634), .B(n23633), .Z(n24167) );
  NOR U24018 ( .A(n24168), .B(n24167), .Z(n23635) );
  NOR U24019 ( .A(n23636), .B(n23635), .Z(n24195) );
  XOR U24020 ( .A(n23638), .B(n23637), .Z(n24194) );
  NOR U24021 ( .A(n24195), .B(n24194), .Z(n23639) );
  NOR U24022 ( .A(n23640), .B(n23639), .Z(n23645) );
  XOR U24023 ( .A(n23642), .B(n23641), .Z(n23644) );
  IV U24024 ( .A(n23644), .Z(n23643) );
  NOR U24025 ( .A(n23645), .B(n23643), .Z(n23648) );
  XOR U24026 ( .A(n23645), .B(n23644), .Z(n24164) );
  NOR U24027 ( .A(n97), .B(n71), .Z(n24165) );
  IV U24028 ( .A(n24165), .Z(n23646) );
  NOR U24029 ( .A(n24164), .B(n23646), .Z(n23647) );
  NOR U24030 ( .A(n23648), .B(n23647), .Z(n24160) );
  XOR U24031 ( .A(n23650), .B(n23649), .Z(n24161) );
  NOR U24032 ( .A(n24160), .B(n24161), .Z(n23651) );
  NOR U24033 ( .A(n23652), .B(n23651), .Z(n24156) );
  XOR U24034 ( .A(n23654), .B(n23653), .Z(n24157) );
  NOR U24035 ( .A(n24156), .B(n24157), .Z(n23655) );
  NOR U24036 ( .A(n23656), .B(n23655), .Z(n24152) );
  XOR U24037 ( .A(n23658), .B(n23657), .Z(n24153) );
  NOR U24038 ( .A(n24152), .B(n24153), .Z(n23659) );
  NOR U24039 ( .A(n23660), .B(n23659), .Z(n24148) );
  XOR U24040 ( .A(n23662), .B(n23661), .Z(n24149) );
  NOR U24041 ( .A(n24148), .B(n24149), .Z(n23663) );
  NOR U24042 ( .A(n23664), .B(n23663), .Z(n24144) );
  XOR U24043 ( .A(n23666), .B(n23665), .Z(n24145) );
  NOR U24044 ( .A(n24144), .B(n24145), .Z(n23667) );
  NOR U24045 ( .A(n23668), .B(n23667), .Z(n24140) );
  XOR U24046 ( .A(n23670), .B(n23669), .Z(n24141) );
  NOR U24047 ( .A(n24140), .B(n24141), .Z(n23671) );
  NOR U24048 ( .A(n23672), .B(n23671), .Z(n24136) );
  XOR U24049 ( .A(n23674), .B(n23673), .Z(n24137) );
  NOR U24050 ( .A(n24136), .B(n24137), .Z(n23675) );
  NOR U24051 ( .A(n23676), .B(n23675), .Z(n24133) );
  XOR U24052 ( .A(n23678), .B(n23677), .Z(n24132) );
  NOR U24053 ( .A(n24133), .B(n24132), .Z(n23679) );
  NOR U24054 ( .A(n23680), .B(n23679), .Z(n24128) );
  XOR U24055 ( .A(n23682), .B(n23681), .Z(n24129) );
  NOR U24056 ( .A(n24128), .B(n24129), .Z(n23683) );
  NOR U24057 ( .A(n23684), .B(n23683), .Z(n23689) );
  XOR U24058 ( .A(n23686), .B(n23685), .Z(n23688) );
  IV U24059 ( .A(n23688), .Z(n23687) );
  NOR U24060 ( .A(n23689), .B(n23687), .Z(n23692) );
  XOR U24061 ( .A(n23689), .B(n23688), .Z(n24125) );
  NOR U24062 ( .A(n104), .B(n71), .Z(n24126) );
  IV U24063 ( .A(n24126), .Z(n23690) );
  NOR U24064 ( .A(n24125), .B(n23690), .Z(n23691) );
  NOR U24065 ( .A(n23692), .B(n23691), .Z(n24121) );
  XOR U24066 ( .A(n23694), .B(n23693), .Z(n24122) );
  NOR U24067 ( .A(n24121), .B(n24122), .Z(n23695) );
  NOR U24068 ( .A(n23696), .B(n23695), .Z(n24117) );
  XOR U24069 ( .A(n23698), .B(n23697), .Z(n24118) );
  NOR U24070 ( .A(n24117), .B(n24118), .Z(n23699) );
  NOR U24071 ( .A(n23700), .B(n23699), .Z(n24113) );
  XOR U24072 ( .A(n23702), .B(n23701), .Z(n24114) );
  NOR U24073 ( .A(n24113), .B(n24114), .Z(n23703) );
  NOR U24074 ( .A(n23704), .B(n23703), .Z(n24110) );
  XOR U24075 ( .A(n23706), .B(n23705), .Z(n24109) );
  NOR U24076 ( .A(n24110), .B(n24109), .Z(n23707) );
  NOR U24077 ( .A(n23708), .B(n23707), .Z(n24263) );
  XOR U24078 ( .A(n23710), .B(n23709), .Z(n24262) );
  NOR U24079 ( .A(n24263), .B(n24262), .Z(n23711) );
  NOR U24080 ( .A(n23712), .B(n23711), .Z(n23717) );
  XOR U24081 ( .A(n23714), .B(n23713), .Z(n23716) );
  IV U24082 ( .A(n23716), .Z(n23715) );
  NOR U24083 ( .A(n23717), .B(n23715), .Z(n23720) );
  XOR U24084 ( .A(n23717), .B(n23716), .Z(n24106) );
  NOR U24085 ( .A(n108), .B(n71), .Z(n24107) );
  IV U24086 ( .A(n24107), .Z(n23718) );
  NOR U24087 ( .A(n24106), .B(n23718), .Z(n23719) );
  NOR U24088 ( .A(n23720), .B(n23719), .Z(n24102) );
  XOR U24089 ( .A(n23722), .B(n23721), .Z(n24103) );
  NOR U24090 ( .A(n24102), .B(n24103), .Z(n23723) );
  NOR U24091 ( .A(n23724), .B(n23723), .Z(n24098) );
  XOR U24092 ( .A(n23726), .B(n23725), .Z(n24099) );
  NOR U24093 ( .A(n24098), .B(n24099), .Z(n23727) );
  NOR U24094 ( .A(n23728), .B(n23727), .Z(n24094) );
  XOR U24095 ( .A(n23730), .B(n23729), .Z(n24095) );
  NOR U24096 ( .A(n24094), .B(n24095), .Z(n23731) );
  NOR U24097 ( .A(n23732), .B(n23731), .Z(n24090) );
  XOR U24098 ( .A(n23734), .B(n23733), .Z(n24091) );
  NOR U24099 ( .A(n24090), .B(n24091), .Z(n23735) );
  NOR U24100 ( .A(n23736), .B(n23735), .Z(n24086) );
  XOR U24101 ( .A(n23738), .B(n23737), .Z(n24087) );
  NOR U24102 ( .A(n24086), .B(n24087), .Z(n23739) );
  NOR U24103 ( .A(n23740), .B(n23739), .Z(n24082) );
  XOR U24104 ( .A(n23742), .B(n23741), .Z(n24083) );
  NOR U24105 ( .A(n24082), .B(n24083), .Z(n23743) );
  NOR U24106 ( .A(n23744), .B(n23743), .Z(n24078) );
  XOR U24107 ( .A(n23746), .B(n23745), .Z(n24079) );
  NOR U24108 ( .A(n24078), .B(n24079), .Z(n23747) );
  NOR U24109 ( .A(n23748), .B(n23747), .Z(n24074) );
  XOR U24110 ( .A(n23750), .B(n23749), .Z(n24075) );
  NOR U24111 ( .A(n24074), .B(n24075), .Z(n23751) );
  NOR U24112 ( .A(n23752), .B(n23751), .Z(n24070) );
  XOR U24113 ( .A(n23754), .B(n23753), .Z(n24071) );
  NOR U24114 ( .A(n24070), .B(n24071), .Z(n23755) );
  NOR U24115 ( .A(n23756), .B(n23755), .Z(n24066) );
  XOR U24116 ( .A(n23758), .B(n23757), .Z(n24067) );
  NOR U24117 ( .A(n24066), .B(n24067), .Z(n23759) );
  NOR U24118 ( .A(n23760), .B(n23759), .Z(n24062) );
  XOR U24119 ( .A(n23762), .B(n23761), .Z(n24063) );
  NOR U24120 ( .A(n24062), .B(n24063), .Z(n23763) );
  NOR U24121 ( .A(n23764), .B(n23763), .Z(n24058) );
  XOR U24122 ( .A(n23766), .B(n23765), .Z(n24059) );
  NOR U24123 ( .A(n24058), .B(n24059), .Z(n23767) );
  NOR U24124 ( .A(n23768), .B(n23767), .Z(n23769) );
  IV U24125 ( .A(n23769), .Z(n24056) );
  XOR U24126 ( .A(n23771), .B(n23770), .Z(n23772) );
  IV U24127 ( .A(n23772), .Z(n24055) );
  NOR U24128 ( .A(n24056), .B(n24055), .Z(n23773) );
  NOR U24129 ( .A(n23774), .B(n23773), .Z(n23775) );
  IV U24130 ( .A(n23775), .Z(n24054) );
  XOR U24131 ( .A(n23777), .B(n23776), .Z(n24053) );
  NOR U24132 ( .A(n24054), .B(n24053), .Z(n23778) );
  NOR U24133 ( .A(n23779), .B(n23778), .Z(n23780) );
  IV U24134 ( .A(n23780), .Z(n24051) );
  XOR U24135 ( .A(n23782), .B(n23781), .Z(n23783) );
  IV U24136 ( .A(n23783), .Z(n24050) );
  NOR U24137 ( .A(n24051), .B(n24050), .Z(n23784) );
  NOR U24138 ( .A(n23785), .B(n23784), .Z(n23786) );
  IV U24139 ( .A(n23786), .Z(n24046) );
  XOR U24140 ( .A(n23788), .B(n23787), .Z(n24045) );
  NOR U24141 ( .A(n24046), .B(n24045), .Z(n23789) );
  NOR U24142 ( .A(n23790), .B(n23789), .Z(n23791) );
  IV U24143 ( .A(n23791), .Z(n24043) );
  XOR U24144 ( .A(n23793), .B(n23792), .Z(n23794) );
  IV U24145 ( .A(n23794), .Z(n24042) );
  NOR U24146 ( .A(n24043), .B(n24042), .Z(n23795) );
  NOR U24147 ( .A(n23796), .B(n23795), .Z(n23797) );
  IV U24148 ( .A(n23797), .Z(n24041) );
  XOR U24149 ( .A(n23799), .B(n23798), .Z(n24040) );
  NOR U24150 ( .A(n24041), .B(n24040), .Z(n23800) );
  NOR U24151 ( .A(n23801), .B(n23800), .Z(n23802) );
  IV U24152 ( .A(n23802), .Z(n24038) );
  XOR U24153 ( .A(n23804), .B(n23803), .Z(n23805) );
  IV U24154 ( .A(n23805), .Z(n24037) );
  NOR U24155 ( .A(n24038), .B(n24037), .Z(n23806) );
  NOR U24156 ( .A(n23807), .B(n23806), .Z(n23808) );
  IV U24157 ( .A(n23808), .Z(n24036) );
  XOR U24158 ( .A(n23810), .B(n23809), .Z(n24035) );
  NOR U24159 ( .A(n24036), .B(n24035), .Z(n23811) );
  NOR U24160 ( .A(n23812), .B(n23811), .Z(n23813) );
  IV U24161 ( .A(n23813), .Z(n24033) );
  XOR U24162 ( .A(n23815), .B(n23814), .Z(n23816) );
  IV U24163 ( .A(n23816), .Z(n24032) );
  NOR U24164 ( .A(n24033), .B(n24032), .Z(n23817) );
  NOR U24165 ( .A(n23818), .B(n23817), .Z(n23819) );
  IV U24166 ( .A(n23819), .Z(n24031) );
  XOR U24167 ( .A(n23821), .B(n23820), .Z(n24030) );
  NOR U24168 ( .A(n24031), .B(n24030), .Z(n23822) );
  NOR U24169 ( .A(n23823), .B(n23822), .Z(n23824) );
  IV U24170 ( .A(n23824), .Z(n24028) );
  XOR U24171 ( .A(n23826), .B(n23825), .Z(n23827) );
  IV U24172 ( .A(n23827), .Z(n24027) );
  NOR U24173 ( .A(n24028), .B(n24027), .Z(n23828) );
  NOR U24174 ( .A(n23829), .B(n23828), .Z(n23830) );
  IV U24175 ( .A(n23830), .Z(n24023) );
  XOR U24176 ( .A(n23832), .B(n23831), .Z(n24022) );
  NOR U24177 ( .A(n24023), .B(n24022), .Z(n23833) );
  NOR U24178 ( .A(n23834), .B(n23833), .Z(n23835) );
  IV U24179 ( .A(n23835), .Z(n24019) );
  NOR U24180 ( .A(n24020), .B(n24019), .Z(n23836) );
  NOR U24181 ( .A(n23837), .B(n23836), .Z(n24017) );
  IV U24182 ( .A(n24017), .Z(n23840) );
  XOR U24183 ( .A(n23839), .B(n23838), .Z(n24016) );
  NOR U24184 ( .A(n23840), .B(n24016), .Z(n23841) );
  NOR U24185 ( .A(n23842), .B(n23841), .Z(n24012) );
  XOR U24186 ( .A(n23844), .B(n23843), .Z(n24013) );
  NOR U24187 ( .A(n24012), .B(n24013), .Z(n23845) );
  NOR U24188 ( .A(n23846), .B(n23845), .Z(n23847) );
  IV U24189 ( .A(n23847), .Z(n24008) );
  NOR U24190 ( .A(n23848), .B(n24008), .Z(n23849) );
  NOR U24191 ( .A(n23850), .B(n23849), .Z(n24002) );
  NOR U24192 ( .A(n23851), .B(n24002), .Z(n23852) );
  NOR U24193 ( .A(n23853), .B(n23852), .Z(n23854) );
  IV U24194 ( .A(n23854), .Z(n23858) );
  NOR U24195 ( .A(n23855), .B(n23858), .Z(n23861) );
  XOR U24196 ( .A(n23857), .B(n23856), .Z(n23999) );
  XOR U24197 ( .A(n23859), .B(n23858), .Z(n23998) );
  NOR U24198 ( .A(n23999), .B(n23998), .Z(n23860) );
  NOR U24199 ( .A(n23861), .B(n23860), .Z(n24408) );
  XOR U24200 ( .A(n23863), .B(n23862), .Z(n24409) );
  NOR U24201 ( .A(n24408), .B(n24409), .Z(n23864) );
  NOR U24202 ( .A(n23865), .B(n23864), .Z(n23995) );
  XOR U24203 ( .A(n23867), .B(n23866), .Z(n23994) );
  NOR U24204 ( .A(n23995), .B(n23994), .Z(n23868) );
  NOR U24205 ( .A(n23869), .B(n23868), .Z(n23870) );
  IV U24206 ( .A(n23870), .Z(n23990) );
  NOR U24207 ( .A(n150), .B(n71), .Z(n23874) );
  IV U24208 ( .A(n23874), .Z(n23871) );
  NOR U24209 ( .A(n23875), .B(n23871), .Z(n23877) );
  XOR U24210 ( .A(n23873), .B(n23872), .Z(n23985) );
  XOR U24211 ( .A(n23875), .B(n23874), .Z(n23986) );
  NOR U24212 ( .A(n23985), .B(n23986), .Z(n23876) );
  NOR U24213 ( .A(n23877), .B(n23876), .Z(n23882) );
  NOR U24214 ( .A(n153), .B(n71), .Z(n23881) );
  IV U24215 ( .A(n23881), .Z(n23878) );
  NOR U24216 ( .A(n23882), .B(n23878), .Z(n23884) );
  XOR U24217 ( .A(n23880), .B(n23879), .Z(n24426) );
  XOR U24218 ( .A(n23882), .B(n23881), .Z(n24425) );
  NOR U24219 ( .A(n24426), .B(n24425), .Z(n23883) );
  NOR U24220 ( .A(n23884), .B(n23883), .Z(n23889) );
  NOR U24221 ( .A(n155), .B(n71), .Z(n23888) );
  IV U24222 ( .A(n23888), .Z(n23885) );
  NOR U24223 ( .A(n23889), .B(n23885), .Z(n23891) );
  XOR U24224 ( .A(n23887), .B(n23886), .Z(n24434) );
  XOR U24225 ( .A(n23889), .B(n23888), .Z(n24433) );
  NOR U24226 ( .A(n24434), .B(n24433), .Z(n23890) );
  NOR U24227 ( .A(n23891), .B(n23890), .Z(n23895) );
  XOR U24228 ( .A(n23893), .B(n23892), .Z(n23894) );
  NOR U24229 ( .A(n23895), .B(n23894), .Z(n23899) );
  XOR U24230 ( .A(n23895), .B(n23894), .Z(n23896) );
  IV U24231 ( .A(n23896), .Z(n24442) );
  NOR U24232 ( .A(n156), .B(n71), .Z(n24443) );
  IV U24233 ( .A(n24443), .Z(n23897) );
  NOR U24234 ( .A(n24442), .B(n23897), .Z(n23898) );
  NOR U24235 ( .A(n23899), .B(n23898), .Z(n23902) );
  NOR U24236 ( .A(n158), .B(n71), .Z(n23901) );
  IV U24237 ( .A(n23901), .Z(n23900) );
  NOR U24238 ( .A(n23902), .B(n23900), .Z(n23907) );
  XOR U24239 ( .A(n23902), .B(n23901), .Z(n24448) );
  XOR U24240 ( .A(n23904), .B(n23903), .Z(n24449) );
  IV U24241 ( .A(n24449), .Z(n23905) );
  NOR U24242 ( .A(n24448), .B(n23905), .Z(n23906) );
  NOR U24243 ( .A(n23907), .B(n23906), .Z(n23912) );
  NOR U24244 ( .A(n161), .B(n71), .Z(n23911) );
  IV U24245 ( .A(n23911), .Z(n23908) );
  NOR U24246 ( .A(n23912), .B(n23908), .Z(n23914) );
  XOR U24247 ( .A(n23910), .B(n23909), .Z(n24457) );
  XOR U24248 ( .A(n23912), .B(n23911), .Z(n24456) );
  NOR U24249 ( .A(n24457), .B(n24456), .Z(n23913) );
  NOR U24250 ( .A(n23914), .B(n23913), .Z(n24468) );
  XOR U24251 ( .A(n23916), .B(n23915), .Z(n24467) );
  NOR U24252 ( .A(n24468), .B(n24467), .Z(n23917) );
  NOR U24253 ( .A(n23918), .B(n23917), .Z(n23931) );
  NOR U24254 ( .A(n165), .B(n71), .Z(n23930) );
  IV U24255 ( .A(n23930), .Z(n23919) );
  NOR U24256 ( .A(n23931), .B(n23919), .Z(n23933) );
  XOR U24257 ( .A(n23921), .B(n23920), .Z(n23939) );
  IV U24258 ( .A(n23922), .Z(n23924) );
  NOR U24259 ( .A(n23924), .B(n23923), .Z(n23928) );
  NOR U24260 ( .A(n23926), .B(n23925), .Z(n23927) );
  NOR U24261 ( .A(n23928), .B(n23927), .Z(n23938) );
  NOR U24262 ( .A(n163), .B(n70), .Z(n23936) );
  XOR U24263 ( .A(n23938), .B(n23936), .Z(n23940) );
  XOR U24264 ( .A(n23939), .B(n23940), .Z(n23929) );
  IV U24265 ( .A(n23929), .Z(n24476) );
  XOR U24266 ( .A(n23931), .B(n23930), .Z(n24475) );
  NOR U24267 ( .A(n24476), .B(n24475), .Z(n23932) );
  NOR U24268 ( .A(n23933), .B(n23932), .Z(n23944) );
  XOR U24269 ( .A(n23935), .B(n23934), .Z(n23954) );
  IV U24270 ( .A(n23936), .Z(n23937) );
  NOR U24271 ( .A(n23938), .B(n23937), .Z(n23942) );
  NOR U24272 ( .A(n23940), .B(n23939), .Z(n23941) );
  NOR U24273 ( .A(n23942), .B(n23941), .Z(n23953) );
  NOR U24274 ( .A(n165), .B(n70), .Z(n23951) );
  XOR U24275 ( .A(n23953), .B(n23951), .Z(n23955) );
  XOR U24276 ( .A(n23954), .B(n23955), .Z(n23943) );
  NOR U24277 ( .A(n23944), .B(n23943), .Z(n23948) );
  XOR U24278 ( .A(n23944), .B(n23943), .Z(n23945) );
  IV U24279 ( .A(n23945), .Z(n23983) );
  NOR U24280 ( .A(n167), .B(n71), .Z(n23946) );
  IV U24281 ( .A(n23946), .Z(n23984) );
  NOR U24282 ( .A(n23983), .B(n23984), .Z(n23947) );
  NOR U24283 ( .A(n23948), .B(n23947), .Z(n24481) );
  XOR U24284 ( .A(n23950), .B(n23949), .Z(n23963) );
  NOR U24285 ( .A(n167), .B(n70), .Z(n23960) );
  IV U24286 ( .A(n23951), .Z(n23952) );
  NOR U24287 ( .A(n23953), .B(n23952), .Z(n23958) );
  IV U24288 ( .A(n23954), .Z(n23956) );
  NOR U24289 ( .A(n23956), .B(n23955), .Z(n23957) );
  NOR U24290 ( .A(n23958), .B(n23957), .Z(n23962) );
  XOR U24291 ( .A(n23960), .B(n23962), .Z(n23964) );
  XOR U24292 ( .A(n23963), .B(n23964), .Z(n23959) );
  IV U24293 ( .A(n23959), .Z(n24480) );
  NOR U24294 ( .A(n24481), .B(n24480), .Z(n23981) );
  IV U24295 ( .A(n23981), .Z(n31515) );
  IV U24296 ( .A(n23960), .Z(n23961) );
  NOR U24297 ( .A(n23962), .B(n23961), .Z(n23966) );
  NOR U24298 ( .A(n23964), .B(n23963), .Z(n23965) );
  NOR U24299 ( .A(n23966), .B(n23965), .Z(n23971) );
  XOR U24300 ( .A(n23968), .B(n23967), .Z(n23970) );
  XOR U24301 ( .A(n23971), .B(n23970), .Z(n31514) );
  IV U24302 ( .A(n31514), .Z(n23969) );
  NOR U24303 ( .A(n31515), .B(n23969), .Z(n31519) );
  NOR U24304 ( .A(n23971), .B(n23970), .Z(n31523) );
  IV U24305 ( .A(n28520), .Z(n23972) );
  NOR U24306 ( .A(n28521), .B(n23972), .Z(n31520) );
  NOR U24307 ( .A(n31523), .B(n31520), .Z(n23973) );
  IV U24308 ( .A(n23973), .Z(n23974) );
  NOR U24309 ( .A(n31519), .B(n23974), .Z(n23977) );
  XOR U24310 ( .A(n23976), .B(n23975), .Z(n23982) );
  IV U24311 ( .A(n23982), .Z(n31534) );
  NOR U24312 ( .A(n23977), .B(n31534), .Z(n23978) );
  IV U24313 ( .A(n23978), .Z(n23979) );
  NOR U24314 ( .A(n23980), .B(n23979), .Z(n28531) );
  NOR U24315 ( .A(n23981), .B(n31514), .Z(n28529) );
  NOR U24316 ( .A(n31520), .B(n23982), .Z(n28526) );
  XOR U24317 ( .A(n23984), .B(n23983), .Z(n31507) );
  IV U24318 ( .A(n31507), .Z(n24483) );
  NOR U24319 ( .A(n153), .B(n72), .Z(n24422) );
  IV U24320 ( .A(n24422), .Z(n23988) );
  XOR U24321 ( .A(n23986), .B(n23985), .Z(n23987) );
  IV U24322 ( .A(n23987), .Z(n24421) );
  NOR U24323 ( .A(n23988), .B(n24421), .Z(n24424) );
  XOR U24324 ( .A(n23990), .B(n23989), .Z(n23991) );
  XOR U24325 ( .A(n23992), .B(n23991), .Z(n24418) );
  NOR U24326 ( .A(n150), .B(n72), .Z(n24417) );
  IV U24327 ( .A(n24417), .Z(n23993) );
  NOR U24328 ( .A(n24418), .B(n23993), .Z(n24420) );
  NOR U24329 ( .A(n148), .B(n72), .Z(n24414) );
  IV U24330 ( .A(n24414), .Z(n23997) );
  IV U24331 ( .A(n23994), .Z(n23996) );
  XOR U24332 ( .A(n23996), .B(n23995), .Z(n24413) );
  NOR U24333 ( .A(n23997), .B(n24413), .Z(n24416) );
  XOR U24334 ( .A(n23999), .B(n23998), .Z(n24001) );
  IV U24335 ( .A(n24001), .Z(n24500) );
  NOR U24336 ( .A(n145), .B(n72), .Z(n24000) );
  IV U24337 ( .A(n24000), .Z(n24499) );
  NOR U24338 ( .A(n24500), .B(n24499), .Z(n24404) );
  NOR U24339 ( .A(n24001), .B(n24000), .Z(n24402) );
  XOR U24340 ( .A(n24003), .B(n24002), .Z(n24004) );
  XOR U24341 ( .A(n24005), .B(n24004), .Z(n24398) );
  NOR U24342 ( .A(n143), .B(n72), .Z(n24399) );
  IV U24343 ( .A(n24399), .Z(n24006) );
  NOR U24344 ( .A(n24398), .B(n24006), .Z(n24401) );
  XOR U24345 ( .A(n24008), .B(n24007), .Z(n24009) );
  XOR U24346 ( .A(n24010), .B(n24009), .Z(n24395) );
  NOR U24347 ( .A(n141), .B(n72), .Z(n24394) );
  IV U24348 ( .A(n24394), .Z(n24011) );
  NOR U24349 ( .A(n24395), .B(n24011), .Z(n24397) );
  IV U24350 ( .A(n24012), .Z(n24014) );
  XOR U24351 ( .A(n24014), .B(n24013), .Z(n24390) );
  NOR U24352 ( .A(n139), .B(n72), .Z(n24391) );
  IV U24353 ( .A(n24391), .Z(n24015) );
  NOR U24354 ( .A(n24390), .B(n24015), .Z(n24393) );
  XOR U24355 ( .A(n24017), .B(n24016), .Z(n24386) );
  NOR U24356 ( .A(n137), .B(n72), .Z(n24387) );
  IV U24357 ( .A(n24387), .Z(n24018) );
  NOR U24358 ( .A(n24386), .B(n24018), .Z(n24389) );
  XOR U24359 ( .A(n24020), .B(n24019), .Z(n24382) );
  NOR U24360 ( .A(n135), .B(n72), .Z(n24381) );
  IV U24361 ( .A(n24381), .Z(n24021) );
  NOR U24362 ( .A(n24382), .B(n24021), .Z(n24385) );
  NOR U24363 ( .A(n133), .B(n72), .Z(n24025) );
  XOR U24364 ( .A(n24023), .B(n24022), .Z(n24024) );
  NOR U24365 ( .A(n24025), .B(n24024), .Z(n24380) );
  XOR U24366 ( .A(n24025), .B(n24024), .Z(n24026) );
  IV U24367 ( .A(n24026), .Z(n24520) );
  XOR U24368 ( .A(n24028), .B(n24027), .Z(n24375) );
  NOR U24369 ( .A(n131), .B(n72), .Z(n24374) );
  IV U24370 ( .A(n24374), .Z(n24029) );
  NOR U24371 ( .A(n24375), .B(n24029), .Z(n24377) );
  NOR U24372 ( .A(n128), .B(n72), .Z(n24369) );
  XOR U24373 ( .A(n24031), .B(n24030), .Z(n24368) );
  NOR U24374 ( .A(n24369), .B(n24368), .Z(n24372) );
  XOR U24375 ( .A(n24033), .B(n24032), .Z(n24364) );
  NOR U24376 ( .A(n126), .B(n72), .Z(n24363) );
  IV U24377 ( .A(n24363), .Z(n24034) );
  NOR U24378 ( .A(n24364), .B(n24034), .Z(n24366) );
  NOR U24379 ( .A(n125), .B(n72), .Z(n24358) );
  XOR U24380 ( .A(n24036), .B(n24035), .Z(n24357) );
  NOR U24381 ( .A(n24358), .B(n24357), .Z(n24361) );
  XOR U24382 ( .A(n24038), .B(n24037), .Z(n24353) );
  NOR U24383 ( .A(n123), .B(n72), .Z(n24352) );
  IV U24384 ( .A(n24352), .Z(n24039) );
  NOR U24385 ( .A(n24353), .B(n24039), .Z(n24355) );
  NOR U24386 ( .A(n120), .B(n72), .Z(n24347) );
  XOR U24387 ( .A(n24041), .B(n24040), .Z(n24346) );
  NOR U24388 ( .A(n24347), .B(n24346), .Z(n24350) );
  XOR U24389 ( .A(n24043), .B(n24042), .Z(n24342) );
  NOR U24390 ( .A(n119), .B(n72), .Z(n24341) );
  IV U24391 ( .A(n24341), .Z(n24044) );
  NOR U24392 ( .A(n24342), .B(n24044), .Z(n24344) );
  NOR U24393 ( .A(n79), .B(n72), .Z(n24048) );
  XOR U24394 ( .A(n24046), .B(n24045), .Z(n24047) );
  NOR U24395 ( .A(n24048), .B(n24047), .Z(n24339) );
  XOR U24396 ( .A(n24048), .B(n24047), .Z(n24049) );
  IV U24397 ( .A(n24049), .Z(n24542) );
  XOR U24398 ( .A(n24051), .B(n24050), .Z(n24334) );
  NOR U24399 ( .A(n117), .B(n72), .Z(n24333) );
  IV U24400 ( .A(n24333), .Z(n24052) );
  NOR U24401 ( .A(n24334), .B(n24052), .Z(n24336) );
  NOR U24402 ( .A(n80), .B(n72), .Z(n24328) );
  XOR U24403 ( .A(n24054), .B(n24053), .Z(n24327) );
  NOR U24404 ( .A(n24328), .B(n24327), .Z(n24331) );
  XOR U24405 ( .A(n24056), .B(n24055), .Z(n24323) );
  NOR U24406 ( .A(n116), .B(n72), .Z(n24322) );
  IV U24407 ( .A(n24322), .Z(n24057) );
  NOR U24408 ( .A(n24323), .B(n24057), .Z(n24325) );
  IV U24409 ( .A(n24058), .Z(n24060) );
  XOR U24410 ( .A(n24060), .B(n24059), .Z(n24318) );
  NOR U24411 ( .A(n81), .B(n72), .Z(n24319) );
  IV U24412 ( .A(n24319), .Z(n24061) );
  NOR U24413 ( .A(n24318), .B(n24061), .Z(n24321) );
  IV U24414 ( .A(n24062), .Z(n24064) );
  XOR U24415 ( .A(n24064), .B(n24063), .Z(n24314) );
  NOR U24416 ( .A(n115), .B(n72), .Z(n24315) );
  IV U24417 ( .A(n24315), .Z(n24065) );
  NOR U24418 ( .A(n24314), .B(n24065), .Z(n24317) );
  IV U24419 ( .A(n24066), .Z(n24068) );
  XOR U24420 ( .A(n24068), .B(n24067), .Z(n24310) );
  NOR U24421 ( .A(n82), .B(n72), .Z(n24311) );
  IV U24422 ( .A(n24311), .Z(n24069) );
  NOR U24423 ( .A(n24310), .B(n24069), .Z(n24313) );
  IV U24424 ( .A(n24070), .Z(n24072) );
  XOR U24425 ( .A(n24072), .B(n24071), .Z(n24306) );
  NOR U24426 ( .A(n114), .B(n72), .Z(n24307) );
  IV U24427 ( .A(n24307), .Z(n24073) );
  NOR U24428 ( .A(n24306), .B(n24073), .Z(n24309) );
  IV U24429 ( .A(n24074), .Z(n24076) );
  XOR U24430 ( .A(n24076), .B(n24075), .Z(n24302) );
  NOR U24431 ( .A(n83), .B(n72), .Z(n24303) );
  IV U24432 ( .A(n24303), .Z(n24077) );
  NOR U24433 ( .A(n24302), .B(n24077), .Z(n24305) );
  IV U24434 ( .A(n24078), .Z(n24080) );
  XOR U24435 ( .A(n24080), .B(n24079), .Z(n24298) );
  NOR U24436 ( .A(n113), .B(n72), .Z(n24299) );
  IV U24437 ( .A(n24299), .Z(n24081) );
  NOR U24438 ( .A(n24298), .B(n24081), .Z(n24301) );
  IV U24439 ( .A(n24082), .Z(n24084) );
  XOR U24440 ( .A(n24084), .B(n24083), .Z(n24294) );
  NOR U24441 ( .A(n84), .B(n72), .Z(n24295) );
  IV U24442 ( .A(n24295), .Z(n24085) );
  NOR U24443 ( .A(n24294), .B(n24085), .Z(n24297) );
  IV U24444 ( .A(n24086), .Z(n24088) );
  XOR U24445 ( .A(n24088), .B(n24087), .Z(n24290) );
  NOR U24446 ( .A(n112), .B(n72), .Z(n24291) );
  IV U24447 ( .A(n24291), .Z(n24089) );
  NOR U24448 ( .A(n24290), .B(n24089), .Z(n24293) );
  IV U24449 ( .A(n24090), .Z(n24092) );
  XOR U24450 ( .A(n24092), .B(n24091), .Z(n24286) );
  NOR U24451 ( .A(n85), .B(n72), .Z(n24287) );
  IV U24452 ( .A(n24287), .Z(n24093) );
  NOR U24453 ( .A(n24286), .B(n24093), .Z(n24289) );
  IV U24454 ( .A(n24094), .Z(n24096) );
  XOR U24455 ( .A(n24096), .B(n24095), .Z(n24282) );
  NOR U24456 ( .A(n111), .B(n72), .Z(n24283) );
  IV U24457 ( .A(n24283), .Z(n24097) );
  NOR U24458 ( .A(n24282), .B(n24097), .Z(n24285) );
  IV U24459 ( .A(n24098), .Z(n24100) );
  XOR U24460 ( .A(n24100), .B(n24099), .Z(n24278) );
  NOR U24461 ( .A(n86), .B(n72), .Z(n24279) );
  IV U24462 ( .A(n24279), .Z(n24101) );
  NOR U24463 ( .A(n24278), .B(n24101), .Z(n24281) );
  IV U24464 ( .A(n24102), .Z(n24104) );
  XOR U24465 ( .A(n24104), .B(n24103), .Z(n24274) );
  NOR U24466 ( .A(n110), .B(n72), .Z(n24275) );
  IV U24467 ( .A(n24275), .Z(n24105) );
  NOR U24468 ( .A(n24274), .B(n24105), .Z(n24277) );
  XOR U24469 ( .A(n24107), .B(n24106), .Z(n24270) );
  NOR U24470 ( .A(n109), .B(n72), .Z(n24271) );
  IV U24471 ( .A(n24271), .Z(n24108) );
  NOR U24472 ( .A(n24270), .B(n24108), .Z(n24273) );
  XOR U24473 ( .A(n24110), .B(n24109), .Z(n24258) );
  IV U24474 ( .A(n24258), .Z(n24112) );
  NOR U24475 ( .A(n87), .B(n72), .Z(n24111) );
  IV U24476 ( .A(n24111), .Z(n24259) );
  NOR U24477 ( .A(n24112), .B(n24259), .Z(n24261) );
  IV U24478 ( .A(n24113), .Z(n24115) );
  XOR U24479 ( .A(n24115), .B(n24114), .Z(n24254) );
  NOR U24480 ( .A(n107), .B(n72), .Z(n24255) );
  IV U24481 ( .A(n24255), .Z(n24116) );
  NOR U24482 ( .A(n24254), .B(n24116), .Z(n24257) );
  IV U24483 ( .A(n24117), .Z(n24119) );
  XOR U24484 ( .A(n24119), .B(n24118), .Z(n24250) );
  NOR U24485 ( .A(n88), .B(n72), .Z(n24251) );
  IV U24486 ( .A(n24251), .Z(n24120) );
  NOR U24487 ( .A(n24250), .B(n24120), .Z(n24253) );
  IV U24488 ( .A(n24121), .Z(n24123) );
  XOR U24489 ( .A(n24123), .B(n24122), .Z(n24246) );
  NOR U24490 ( .A(n106), .B(n72), .Z(n24247) );
  IV U24491 ( .A(n24247), .Z(n24124) );
  NOR U24492 ( .A(n24246), .B(n24124), .Z(n24249) );
  XOR U24493 ( .A(n24126), .B(n24125), .Z(n24242) );
  NOR U24494 ( .A(n105), .B(n72), .Z(n24243) );
  IV U24495 ( .A(n24243), .Z(n24127) );
  NOR U24496 ( .A(n24242), .B(n24127), .Z(n24245) );
  IV U24497 ( .A(n24128), .Z(n24130) );
  XOR U24498 ( .A(n24130), .B(n24129), .Z(n24238) );
  NOR U24499 ( .A(n104), .B(n72), .Z(n24239) );
  IV U24500 ( .A(n24239), .Z(n24131) );
  NOR U24501 ( .A(n24238), .B(n24131), .Z(n24241) );
  XOR U24502 ( .A(n24133), .B(n24132), .Z(n24234) );
  IV U24503 ( .A(n24234), .Z(n24135) );
  NOR U24504 ( .A(n89), .B(n72), .Z(n24134) );
  IV U24505 ( .A(n24134), .Z(n24235) );
  NOR U24506 ( .A(n24135), .B(n24235), .Z(n24237) );
  IV U24507 ( .A(n24136), .Z(n24138) );
  XOR U24508 ( .A(n24138), .B(n24137), .Z(n24230) );
  NOR U24509 ( .A(n103), .B(n72), .Z(n24231) );
  IV U24510 ( .A(n24231), .Z(n24139) );
  NOR U24511 ( .A(n24230), .B(n24139), .Z(n24233) );
  IV U24512 ( .A(n24140), .Z(n24142) );
  XOR U24513 ( .A(n24142), .B(n24141), .Z(n24226) );
  NOR U24514 ( .A(n90), .B(n72), .Z(n24227) );
  IV U24515 ( .A(n24227), .Z(n24143) );
  NOR U24516 ( .A(n24226), .B(n24143), .Z(n24229) );
  IV U24517 ( .A(n24144), .Z(n24146) );
  XOR U24518 ( .A(n24146), .B(n24145), .Z(n24222) );
  NOR U24519 ( .A(n102), .B(n72), .Z(n24223) );
  IV U24520 ( .A(n24223), .Z(n24147) );
  NOR U24521 ( .A(n24222), .B(n24147), .Z(n24225) );
  IV U24522 ( .A(n24148), .Z(n24150) );
  XOR U24523 ( .A(n24150), .B(n24149), .Z(n24218) );
  NOR U24524 ( .A(n101), .B(n72), .Z(n24219) );
  IV U24525 ( .A(n24219), .Z(n24151) );
  NOR U24526 ( .A(n24218), .B(n24151), .Z(n24221) );
  IV U24527 ( .A(n24152), .Z(n24154) );
  XOR U24528 ( .A(n24154), .B(n24153), .Z(n24214) );
  NOR U24529 ( .A(n100), .B(n72), .Z(n24215) );
  IV U24530 ( .A(n24215), .Z(n24155) );
  NOR U24531 ( .A(n24214), .B(n24155), .Z(n24217) );
  IV U24532 ( .A(n24156), .Z(n24158) );
  XOR U24533 ( .A(n24158), .B(n24157), .Z(n24210) );
  NOR U24534 ( .A(n99), .B(n72), .Z(n24211) );
  IV U24535 ( .A(n24211), .Z(n24159) );
  NOR U24536 ( .A(n24210), .B(n24159), .Z(n24213) );
  IV U24537 ( .A(n24160), .Z(n24162) );
  XOR U24538 ( .A(n24162), .B(n24161), .Z(n24206) );
  NOR U24539 ( .A(n98), .B(n72), .Z(n24207) );
  IV U24540 ( .A(n24207), .Z(n24163) );
  NOR U24541 ( .A(n24206), .B(n24163), .Z(n24209) );
  XOR U24542 ( .A(n24165), .B(n24164), .Z(n24202) );
  NOR U24543 ( .A(n91), .B(n72), .Z(n24203) );
  IV U24544 ( .A(n24203), .Z(n24166) );
  NOR U24545 ( .A(n24202), .B(n24166), .Z(n24205) );
  XOR U24546 ( .A(n24168), .B(n24167), .Z(n24190) );
  IV U24547 ( .A(n24190), .Z(n24170) );
  NOR U24548 ( .A(n96), .B(n72), .Z(n24169) );
  IV U24549 ( .A(n24169), .Z(n24191) );
  NOR U24550 ( .A(n24170), .B(n24191), .Z(n24193) );
  NOR U24551 ( .A(n95), .B(n72), .Z(n24187) );
  IV U24552 ( .A(n24187), .Z(n24173) );
  XOR U24553 ( .A(n24172), .B(n24171), .Z(n24186) );
  NOR U24554 ( .A(n24173), .B(n24186), .Z(n24189) );
  NOR U24555 ( .A(n93), .B(n72), .Z(n25175) );
  IV U24556 ( .A(n25175), .Z(n24174) );
  NOR U24557 ( .A(n71), .B(n168), .Z(n24182) );
  IV U24558 ( .A(n24182), .Z(n24177) );
  NOR U24559 ( .A(n24174), .B(n24177), .Z(n24175) );
  IV U24560 ( .A(n24175), .Z(n24176) );
  NOR U24561 ( .A(n94), .B(n24176), .Z(n24185) );
  NOR U24562 ( .A(n24177), .B(n93), .Z(n24178) );
  XOR U24563 ( .A(n94), .B(n24178), .Z(n24179) );
  NOR U24564 ( .A(n72), .B(n24179), .Z(n24180) );
  IV U24565 ( .A(n24180), .Z(n24666) );
  XOR U24566 ( .A(n24182), .B(n24181), .Z(n24665) );
  IV U24567 ( .A(n24665), .Z(n24183) );
  NOR U24568 ( .A(n24666), .B(n24183), .Z(n24184) );
  NOR U24569 ( .A(n24185), .B(n24184), .Z(n24662) );
  XOR U24570 ( .A(n24187), .B(n24186), .Z(n24661) );
  NOR U24571 ( .A(n24662), .B(n24661), .Z(n24188) );
  NOR U24572 ( .A(n24189), .B(n24188), .Z(n24689) );
  XOR U24573 ( .A(n24191), .B(n24190), .Z(n24688) );
  NOR U24574 ( .A(n24689), .B(n24688), .Z(n24192) );
  NOR U24575 ( .A(n24193), .B(n24192), .Z(n24198) );
  XOR U24576 ( .A(n24195), .B(n24194), .Z(n24197) );
  IV U24577 ( .A(n24197), .Z(n24196) );
  NOR U24578 ( .A(n24198), .B(n24196), .Z(n24201) );
  XOR U24579 ( .A(n24198), .B(n24197), .Z(n24658) );
  NOR U24580 ( .A(n97), .B(n72), .Z(n24659) );
  IV U24581 ( .A(n24659), .Z(n24199) );
  NOR U24582 ( .A(n24658), .B(n24199), .Z(n24200) );
  NOR U24583 ( .A(n24201), .B(n24200), .Z(n24654) );
  XOR U24584 ( .A(n24203), .B(n24202), .Z(n24655) );
  NOR U24585 ( .A(n24654), .B(n24655), .Z(n24204) );
  NOR U24586 ( .A(n24205), .B(n24204), .Z(n24650) );
  XOR U24587 ( .A(n24207), .B(n24206), .Z(n24651) );
  NOR U24588 ( .A(n24650), .B(n24651), .Z(n24208) );
  NOR U24589 ( .A(n24209), .B(n24208), .Z(n24646) );
  XOR U24590 ( .A(n24211), .B(n24210), .Z(n24647) );
  NOR U24591 ( .A(n24646), .B(n24647), .Z(n24212) );
  NOR U24592 ( .A(n24213), .B(n24212), .Z(n24642) );
  XOR U24593 ( .A(n24215), .B(n24214), .Z(n24643) );
  NOR U24594 ( .A(n24642), .B(n24643), .Z(n24216) );
  NOR U24595 ( .A(n24217), .B(n24216), .Z(n24638) );
  XOR U24596 ( .A(n24219), .B(n24218), .Z(n24639) );
  NOR U24597 ( .A(n24638), .B(n24639), .Z(n24220) );
  NOR U24598 ( .A(n24221), .B(n24220), .Z(n24634) );
  XOR U24599 ( .A(n24223), .B(n24222), .Z(n24635) );
  NOR U24600 ( .A(n24634), .B(n24635), .Z(n24224) );
  NOR U24601 ( .A(n24225), .B(n24224), .Z(n24630) );
  XOR U24602 ( .A(n24227), .B(n24226), .Z(n24631) );
  NOR U24603 ( .A(n24630), .B(n24631), .Z(n24228) );
  NOR U24604 ( .A(n24229), .B(n24228), .Z(n24627) );
  XOR U24605 ( .A(n24231), .B(n24230), .Z(n24626) );
  NOR U24606 ( .A(n24627), .B(n24626), .Z(n24232) );
  NOR U24607 ( .A(n24233), .B(n24232), .Z(n24733) );
  XOR U24608 ( .A(n24235), .B(n24234), .Z(n24732) );
  NOR U24609 ( .A(n24733), .B(n24732), .Z(n24236) );
  NOR U24610 ( .A(n24237), .B(n24236), .Z(n24622) );
  XOR U24611 ( .A(n24239), .B(n24238), .Z(n24623) );
  NOR U24612 ( .A(n24622), .B(n24623), .Z(n24240) );
  NOR U24613 ( .A(n24241), .B(n24240), .Z(n24618) );
  XOR U24614 ( .A(n24243), .B(n24242), .Z(n24619) );
  NOR U24615 ( .A(n24618), .B(n24619), .Z(n24244) );
  NOR U24616 ( .A(n24245), .B(n24244), .Z(n24614) );
  XOR U24617 ( .A(n24247), .B(n24246), .Z(n24615) );
  NOR U24618 ( .A(n24614), .B(n24615), .Z(n24248) );
  NOR U24619 ( .A(n24249), .B(n24248), .Z(n24610) );
  XOR U24620 ( .A(n24251), .B(n24250), .Z(n24611) );
  NOR U24621 ( .A(n24610), .B(n24611), .Z(n24252) );
  NOR U24622 ( .A(n24253), .B(n24252), .Z(n24607) );
  XOR U24623 ( .A(n24255), .B(n24254), .Z(n24606) );
  NOR U24624 ( .A(n24607), .B(n24606), .Z(n24256) );
  NOR U24625 ( .A(n24257), .B(n24256), .Z(n24761) );
  XOR U24626 ( .A(n24259), .B(n24258), .Z(n24760) );
  NOR U24627 ( .A(n24761), .B(n24760), .Z(n24260) );
  NOR U24628 ( .A(n24261), .B(n24260), .Z(n24266) );
  XOR U24629 ( .A(n24263), .B(n24262), .Z(n24265) );
  IV U24630 ( .A(n24265), .Z(n24264) );
  NOR U24631 ( .A(n24266), .B(n24264), .Z(n24269) );
  XOR U24632 ( .A(n24266), .B(n24265), .Z(n24603) );
  NOR U24633 ( .A(n108), .B(n72), .Z(n24604) );
  IV U24634 ( .A(n24604), .Z(n24267) );
  NOR U24635 ( .A(n24603), .B(n24267), .Z(n24268) );
  NOR U24636 ( .A(n24269), .B(n24268), .Z(n24599) );
  XOR U24637 ( .A(n24271), .B(n24270), .Z(n24600) );
  NOR U24638 ( .A(n24599), .B(n24600), .Z(n24272) );
  NOR U24639 ( .A(n24273), .B(n24272), .Z(n24595) );
  XOR U24640 ( .A(n24275), .B(n24274), .Z(n24596) );
  NOR U24641 ( .A(n24595), .B(n24596), .Z(n24276) );
  NOR U24642 ( .A(n24277), .B(n24276), .Z(n24591) );
  XOR U24643 ( .A(n24279), .B(n24278), .Z(n24592) );
  NOR U24644 ( .A(n24591), .B(n24592), .Z(n24280) );
  NOR U24645 ( .A(n24281), .B(n24280), .Z(n24587) );
  XOR U24646 ( .A(n24283), .B(n24282), .Z(n24588) );
  NOR U24647 ( .A(n24587), .B(n24588), .Z(n24284) );
  NOR U24648 ( .A(n24285), .B(n24284), .Z(n24583) );
  XOR U24649 ( .A(n24287), .B(n24286), .Z(n24584) );
  NOR U24650 ( .A(n24583), .B(n24584), .Z(n24288) );
  NOR U24651 ( .A(n24289), .B(n24288), .Z(n24579) );
  XOR U24652 ( .A(n24291), .B(n24290), .Z(n24580) );
  NOR U24653 ( .A(n24579), .B(n24580), .Z(n24292) );
  NOR U24654 ( .A(n24293), .B(n24292), .Z(n24575) );
  XOR U24655 ( .A(n24295), .B(n24294), .Z(n24576) );
  NOR U24656 ( .A(n24575), .B(n24576), .Z(n24296) );
  NOR U24657 ( .A(n24297), .B(n24296), .Z(n24571) );
  XOR U24658 ( .A(n24299), .B(n24298), .Z(n24572) );
  NOR U24659 ( .A(n24571), .B(n24572), .Z(n24300) );
  NOR U24660 ( .A(n24301), .B(n24300), .Z(n24567) );
  XOR U24661 ( .A(n24303), .B(n24302), .Z(n24568) );
  NOR U24662 ( .A(n24567), .B(n24568), .Z(n24304) );
  NOR U24663 ( .A(n24305), .B(n24304), .Z(n24563) );
  XOR U24664 ( .A(n24307), .B(n24306), .Z(n24564) );
  NOR U24665 ( .A(n24563), .B(n24564), .Z(n24308) );
  NOR U24666 ( .A(n24309), .B(n24308), .Z(n24559) );
  XOR U24667 ( .A(n24311), .B(n24310), .Z(n24560) );
  NOR U24668 ( .A(n24559), .B(n24560), .Z(n24312) );
  NOR U24669 ( .A(n24313), .B(n24312), .Z(n24555) );
  XOR U24670 ( .A(n24315), .B(n24314), .Z(n24556) );
  NOR U24671 ( .A(n24555), .B(n24556), .Z(n24316) );
  NOR U24672 ( .A(n24317), .B(n24316), .Z(n24551) );
  XOR U24673 ( .A(n24319), .B(n24318), .Z(n24552) );
  NOR U24674 ( .A(n24551), .B(n24552), .Z(n24320) );
  NOR U24675 ( .A(n24321), .B(n24320), .Z(n24550) );
  XOR U24676 ( .A(n24323), .B(n24322), .Z(n24549) );
  NOR U24677 ( .A(n24550), .B(n24549), .Z(n24324) );
  NOR U24678 ( .A(n24325), .B(n24324), .Z(n24326) );
  IV U24679 ( .A(n24326), .Z(n24547) );
  XOR U24680 ( .A(n24328), .B(n24327), .Z(n24329) );
  IV U24681 ( .A(n24329), .Z(n24546) );
  NOR U24682 ( .A(n24547), .B(n24546), .Z(n24330) );
  NOR U24683 ( .A(n24331), .B(n24330), .Z(n24332) );
  IV U24684 ( .A(n24332), .Z(n24545) );
  XOR U24685 ( .A(n24334), .B(n24333), .Z(n24544) );
  NOR U24686 ( .A(n24545), .B(n24544), .Z(n24335) );
  NOR U24687 ( .A(n24336), .B(n24335), .Z(n24337) );
  IV U24688 ( .A(n24337), .Z(n24541) );
  NOR U24689 ( .A(n24542), .B(n24541), .Z(n24338) );
  NOR U24690 ( .A(n24339), .B(n24338), .Z(n24340) );
  IV U24691 ( .A(n24340), .Z(n24540) );
  XOR U24692 ( .A(n24342), .B(n24341), .Z(n24539) );
  NOR U24693 ( .A(n24540), .B(n24539), .Z(n24343) );
  NOR U24694 ( .A(n24344), .B(n24343), .Z(n24345) );
  IV U24695 ( .A(n24345), .Z(n24537) );
  XOR U24696 ( .A(n24347), .B(n24346), .Z(n24348) );
  IV U24697 ( .A(n24348), .Z(n24536) );
  NOR U24698 ( .A(n24537), .B(n24536), .Z(n24349) );
  NOR U24699 ( .A(n24350), .B(n24349), .Z(n24351) );
  IV U24700 ( .A(n24351), .Z(n24535) );
  XOR U24701 ( .A(n24353), .B(n24352), .Z(n24534) );
  NOR U24702 ( .A(n24535), .B(n24534), .Z(n24354) );
  NOR U24703 ( .A(n24355), .B(n24354), .Z(n24356) );
  IV U24704 ( .A(n24356), .Z(n24532) );
  XOR U24705 ( .A(n24358), .B(n24357), .Z(n24359) );
  IV U24706 ( .A(n24359), .Z(n24531) );
  NOR U24707 ( .A(n24532), .B(n24531), .Z(n24360) );
  NOR U24708 ( .A(n24361), .B(n24360), .Z(n24362) );
  IV U24709 ( .A(n24362), .Z(n24530) );
  XOR U24710 ( .A(n24364), .B(n24363), .Z(n24529) );
  NOR U24711 ( .A(n24530), .B(n24529), .Z(n24365) );
  NOR U24712 ( .A(n24366), .B(n24365), .Z(n24367) );
  IV U24713 ( .A(n24367), .Z(n24527) );
  XOR U24714 ( .A(n24369), .B(n24368), .Z(n24370) );
  IV U24715 ( .A(n24370), .Z(n24526) );
  NOR U24716 ( .A(n24527), .B(n24526), .Z(n24371) );
  NOR U24717 ( .A(n24372), .B(n24371), .Z(n24373) );
  IV U24718 ( .A(n24373), .Z(n24525) );
  XOR U24719 ( .A(n24375), .B(n24374), .Z(n24524) );
  NOR U24720 ( .A(n24525), .B(n24524), .Z(n24376) );
  NOR U24721 ( .A(n24377), .B(n24376), .Z(n24378) );
  IV U24722 ( .A(n24378), .Z(n24519) );
  NOR U24723 ( .A(n24520), .B(n24519), .Z(n24379) );
  NOR U24724 ( .A(n24380), .B(n24379), .Z(n24517) );
  IV U24725 ( .A(n24517), .Z(n24383) );
  XOR U24726 ( .A(n24382), .B(n24381), .Z(n24516) );
  NOR U24727 ( .A(n24383), .B(n24516), .Z(n24384) );
  NOR U24728 ( .A(n24385), .B(n24384), .Z(n24512) );
  XOR U24729 ( .A(n24387), .B(n24386), .Z(n24513) );
  NOR U24730 ( .A(n24512), .B(n24513), .Z(n24388) );
  NOR U24731 ( .A(n24389), .B(n24388), .Z(n24508) );
  XOR U24732 ( .A(n24391), .B(n24390), .Z(n24509) );
  NOR U24733 ( .A(n24508), .B(n24509), .Z(n24392) );
  NOR U24734 ( .A(n24393), .B(n24392), .Z(n24901) );
  XOR U24735 ( .A(n24395), .B(n24394), .Z(n24900) );
  NOR U24736 ( .A(n24901), .B(n24900), .Z(n24396) );
  NOR U24737 ( .A(n24397), .B(n24396), .Z(n24504) );
  XOR U24738 ( .A(n24399), .B(n24398), .Z(n24505) );
  NOR U24739 ( .A(n24504), .B(n24505), .Z(n24400) );
  NOR U24740 ( .A(n24401), .B(n24400), .Z(n24502) );
  NOR U24741 ( .A(n24402), .B(n24502), .Z(n24403) );
  NOR U24742 ( .A(n24404), .B(n24403), .Z(n24407) );
  NOR U24743 ( .A(n147), .B(n72), .Z(n24406) );
  IV U24744 ( .A(n24406), .Z(n24405) );
  NOR U24745 ( .A(n24407), .B(n24405), .Z(n24412) );
  XOR U24746 ( .A(n24407), .B(n24406), .Z(n24496) );
  XOR U24747 ( .A(n24409), .B(n24408), .Z(n24410) );
  IV U24748 ( .A(n24410), .Z(n24495) );
  NOR U24749 ( .A(n24496), .B(n24495), .Z(n24411) );
  NOR U24750 ( .A(n24412), .B(n24411), .Z(n24924) );
  XOR U24751 ( .A(n24414), .B(n24413), .Z(n24925) );
  NOR U24752 ( .A(n24924), .B(n24925), .Z(n24415) );
  NOR U24753 ( .A(n24416), .B(n24415), .Z(n24491) );
  XOR U24754 ( .A(n24418), .B(n24417), .Z(n24492) );
  NOR U24755 ( .A(n24491), .B(n24492), .Z(n24419) );
  NOR U24756 ( .A(n24420), .B(n24419), .Z(n24934) );
  XOR U24757 ( .A(n24422), .B(n24421), .Z(n24933) );
  NOR U24758 ( .A(n24934), .B(n24933), .Z(n24423) );
  NOR U24759 ( .A(n24424), .B(n24423), .Z(n24429) );
  XOR U24760 ( .A(n24426), .B(n24425), .Z(n24428) );
  IV U24761 ( .A(n24428), .Z(n24427) );
  NOR U24762 ( .A(n24429), .B(n24427), .Z(n24432) );
  XOR U24763 ( .A(n24429), .B(n24428), .Z(n24941) );
  NOR U24764 ( .A(n155), .B(n72), .Z(n24942) );
  IV U24765 ( .A(n24942), .Z(n24430) );
  NOR U24766 ( .A(n24941), .B(n24430), .Z(n24431) );
  NOR U24767 ( .A(n24432), .B(n24431), .Z(n24436) );
  XOR U24768 ( .A(n24434), .B(n24433), .Z(n24950) );
  IV U24769 ( .A(n24950), .Z(n24435) );
  NOR U24770 ( .A(n24436), .B(n24435), .Z(n24440) );
  IV U24771 ( .A(n24436), .Z(n24947) );
  NOR U24772 ( .A(n24950), .B(n24947), .Z(n24438) );
  NOR U24773 ( .A(n156), .B(n72), .Z(n24437) );
  IV U24774 ( .A(n24437), .Z(n24948) );
  NOR U24775 ( .A(n24438), .B(n24948), .Z(n24439) );
  NOR U24776 ( .A(n24440), .B(n24439), .Z(n24445) );
  NOR U24777 ( .A(n158), .B(n72), .Z(n24444) );
  IV U24778 ( .A(n24444), .Z(n24441) );
  NOR U24779 ( .A(n24445), .B(n24441), .Z(n24447) );
  XOR U24780 ( .A(n24443), .B(n24442), .Z(n24488) );
  XOR U24781 ( .A(n24445), .B(n24444), .Z(n24487) );
  NOR U24782 ( .A(n24488), .B(n24487), .Z(n24446) );
  NOR U24783 ( .A(n24447), .B(n24446), .Z(n24451) );
  XOR U24784 ( .A(n24449), .B(n24448), .Z(n24450) );
  NOR U24785 ( .A(n24451), .B(n24450), .Z(n24455) );
  XOR U24786 ( .A(n24451), .B(n24450), .Z(n24962) );
  IV U24787 ( .A(n24962), .Z(n24453) );
  NOR U24788 ( .A(n161), .B(n72), .Z(n24452) );
  IV U24789 ( .A(n24452), .Z(n24963) );
  NOR U24790 ( .A(n24453), .B(n24963), .Z(n24454) );
  NOR U24791 ( .A(n24455), .B(n24454), .Z(n24460) );
  XOR U24792 ( .A(n24457), .B(n24456), .Z(n24459) );
  IV U24793 ( .A(n24459), .Z(n24458) );
  NOR U24794 ( .A(n24460), .B(n24458), .Z(n24463) );
  XOR U24795 ( .A(n24460), .B(n24459), .Z(n24969) );
  NOR U24796 ( .A(n163), .B(n72), .Z(n24968) );
  IV U24797 ( .A(n24968), .Z(n24461) );
  NOR U24798 ( .A(n24969), .B(n24461), .Z(n24462) );
  NOR U24799 ( .A(n24463), .B(n24462), .Z(n24466) );
  NOR U24800 ( .A(n165), .B(n72), .Z(n24465) );
  IV U24801 ( .A(n24465), .Z(n24464) );
  NOR U24802 ( .A(n24466), .B(n24464), .Z(n24471) );
  XOR U24803 ( .A(n24466), .B(n24465), .Z(n24485) );
  XOR U24804 ( .A(n24468), .B(n24467), .Z(n24484) );
  IV U24805 ( .A(n24484), .Z(n24469) );
  NOR U24806 ( .A(n24485), .B(n24469), .Z(n24470) );
  NOR U24807 ( .A(n24471), .B(n24470), .Z(n24474) );
  NOR U24808 ( .A(n167), .B(n72), .Z(n24473) );
  IV U24809 ( .A(n24473), .Z(n24472) );
  NOR U24810 ( .A(n24474), .B(n24472), .Z(n24479) );
  XOR U24811 ( .A(n24474), .B(n24473), .Z(n24980) );
  XOR U24812 ( .A(n24476), .B(n24475), .Z(n24981) );
  IV U24813 ( .A(n24981), .Z(n24477) );
  NOR U24814 ( .A(n24980), .B(n24477), .Z(n24478) );
  NOR U24815 ( .A(n24479), .B(n24478), .Z(n31506) );
  NOR U24816 ( .A(n24483), .B(n31506), .Z(n31504) );
  IV U24817 ( .A(n31504), .Z(n24482) );
  XOR U24818 ( .A(n24481), .B(n24480), .Z(n28512) );
  IV U24819 ( .A(n28512), .Z(n31513) );
  NOR U24820 ( .A(n24482), .B(n31513), .Z(n28519) );
  XOR U24821 ( .A(n31506), .B(n24483), .Z(n31503) );
  IV U24822 ( .A(n31503), .Z(n24982) );
  XOR U24823 ( .A(n24485), .B(n24484), .Z(n24977) );
  NOR U24824 ( .A(n167), .B(n73), .Z(n24976) );
  IV U24825 ( .A(n24976), .Z(n24486) );
  NOR U24826 ( .A(n24977), .B(n24486), .Z(n24979) );
  XOR U24827 ( .A(n24488), .B(n24487), .Z(n24489) );
  IV U24828 ( .A(n24489), .Z(n24957) );
  NOR U24829 ( .A(n161), .B(n73), .Z(n24958) );
  IV U24830 ( .A(n24958), .Z(n24490) );
  NOR U24831 ( .A(n24957), .B(n24490), .Z(n24960) );
  NOR U24832 ( .A(n155), .B(n73), .Z(n24935) );
  XOR U24833 ( .A(n24492), .B(n24491), .Z(n24494) );
  IV U24834 ( .A(n24494), .Z(n25429) );
  NOR U24835 ( .A(n153), .B(n73), .Z(n24493) );
  IV U24836 ( .A(n24493), .Z(n25428) );
  NOR U24837 ( .A(n25429), .B(n25428), .Z(n24931) );
  NOR U24838 ( .A(n24494), .B(n24493), .Z(n24929) );
  NOR U24839 ( .A(n148), .B(n73), .Z(n24497) );
  XOR U24840 ( .A(n24496), .B(n24495), .Z(n25414) );
  NOR U24841 ( .A(n24497), .B(n25414), .Z(n24919) );
  IV U24842 ( .A(n24497), .Z(n25411) );
  IV U24843 ( .A(n25414), .Z(n24498) );
  NOR U24844 ( .A(n25411), .B(n24498), .Z(n24917) );
  XOR U24845 ( .A(n24500), .B(n24499), .Z(n24501) );
  XOR U24846 ( .A(n24502), .B(n24501), .Z(n24912) );
  NOR U24847 ( .A(n147), .B(n73), .Z(n24913) );
  IV U24848 ( .A(n24913), .Z(n24503) );
  NOR U24849 ( .A(n24912), .B(n24503), .Z(n24915) );
  IV U24850 ( .A(n24504), .Z(n24506) );
  XOR U24851 ( .A(n24506), .B(n24505), .Z(n24908) );
  NOR U24852 ( .A(n145), .B(n73), .Z(n24909) );
  IV U24853 ( .A(n24909), .Z(n24507) );
  NOR U24854 ( .A(n24908), .B(n24507), .Z(n24911) );
  IV U24855 ( .A(n24508), .Z(n24510) );
  XOR U24856 ( .A(n24510), .B(n24509), .Z(n24896) );
  NOR U24857 ( .A(n141), .B(n73), .Z(n24897) );
  IV U24858 ( .A(n24897), .Z(n24511) );
  NOR U24859 ( .A(n24896), .B(n24511), .Z(n24899) );
  IV U24860 ( .A(n24512), .Z(n24514) );
  XOR U24861 ( .A(n24514), .B(n24513), .Z(n24892) );
  NOR U24862 ( .A(n139), .B(n73), .Z(n24893) );
  IV U24863 ( .A(n24893), .Z(n24515) );
  NOR U24864 ( .A(n24892), .B(n24515), .Z(n24895) );
  XOR U24865 ( .A(n24517), .B(n24516), .Z(n24888) );
  NOR U24866 ( .A(n137), .B(n73), .Z(n24889) );
  IV U24867 ( .A(n24889), .Z(n24518) );
  NOR U24868 ( .A(n24888), .B(n24518), .Z(n24891) );
  XOR U24869 ( .A(n24520), .B(n24519), .Z(n24523) );
  NOR U24870 ( .A(n135), .B(n73), .Z(n24522) );
  IV U24871 ( .A(n24522), .Z(n24521) );
  NOR U24872 ( .A(n24523), .B(n24521), .Z(n24887) );
  XOR U24873 ( .A(n24523), .B(n24522), .Z(n25014) );
  NOR U24874 ( .A(n133), .B(n73), .Z(n24881) );
  XOR U24875 ( .A(n24525), .B(n24524), .Z(n24880) );
  NOR U24876 ( .A(n24881), .B(n24880), .Z(n24884) );
  XOR U24877 ( .A(n24527), .B(n24526), .Z(n24876) );
  NOR U24878 ( .A(n131), .B(n73), .Z(n24875) );
  IV U24879 ( .A(n24875), .Z(n24528) );
  NOR U24880 ( .A(n24876), .B(n24528), .Z(n24878) );
  NOR U24881 ( .A(n128), .B(n73), .Z(n24870) );
  XOR U24882 ( .A(n24530), .B(n24529), .Z(n24869) );
  NOR U24883 ( .A(n24870), .B(n24869), .Z(n24873) );
  XOR U24884 ( .A(n24532), .B(n24531), .Z(n24865) );
  NOR U24885 ( .A(n126), .B(n73), .Z(n24864) );
  IV U24886 ( .A(n24864), .Z(n24533) );
  NOR U24887 ( .A(n24865), .B(n24533), .Z(n24867) );
  NOR U24888 ( .A(n125), .B(n73), .Z(n24859) );
  XOR U24889 ( .A(n24535), .B(n24534), .Z(n24858) );
  NOR U24890 ( .A(n24859), .B(n24858), .Z(n24862) );
  XOR U24891 ( .A(n24537), .B(n24536), .Z(n24854) );
  NOR U24892 ( .A(n123), .B(n73), .Z(n24853) );
  IV U24893 ( .A(n24853), .Z(n24538) );
  NOR U24894 ( .A(n24854), .B(n24538), .Z(n24856) );
  NOR U24895 ( .A(n120), .B(n73), .Z(n24848) );
  XOR U24896 ( .A(n24540), .B(n24539), .Z(n24847) );
  NOR U24897 ( .A(n24848), .B(n24847), .Z(n24851) );
  XOR U24898 ( .A(n24542), .B(n24541), .Z(n24843) );
  NOR U24899 ( .A(n119), .B(n73), .Z(n24842) );
  IV U24900 ( .A(n24842), .Z(n24543) );
  NOR U24901 ( .A(n24843), .B(n24543), .Z(n24845) );
  NOR U24902 ( .A(n79), .B(n73), .Z(n24837) );
  XOR U24903 ( .A(n24545), .B(n24544), .Z(n24836) );
  NOR U24904 ( .A(n24837), .B(n24836), .Z(n24840) );
  XOR U24905 ( .A(n24547), .B(n24546), .Z(n24832) );
  NOR U24906 ( .A(n117), .B(n73), .Z(n24831) );
  IV U24907 ( .A(n24831), .Z(n24548) );
  NOR U24908 ( .A(n24832), .B(n24548), .Z(n24834) );
  NOR U24909 ( .A(n80), .B(n73), .Z(n24826) );
  XOR U24910 ( .A(n24550), .B(n24549), .Z(n24825) );
  NOR U24911 ( .A(n24826), .B(n24825), .Z(n24829) );
  IV U24912 ( .A(n24551), .Z(n24553) );
  XOR U24913 ( .A(n24553), .B(n24552), .Z(n24820) );
  NOR U24914 ( .A(n116), .B(n73), .Z(n24821) );
  IV U24915 ( .A(n24821), .Z(n24554) );
  NOR U24916 ( .A(n24820), .B(n24554), .Z(n24823) );
  IV U24917 ( .A(n24555), .Z(n24557) );
  XOR U24918 ( .A(n24557), .B(n24556), .Z(n24816) );
  NOR U24919 ( .A(n81), .B(n73), .Z(n24817) );
  IV U24920 ( .A(n24817), .Z(n24558) );
  NOR U24921 ( .A(n24816), .B(n24558), .Z(n24819) );
  IV U24922 ( .A(n24559), .Z(n24561) );
  XOR U24923 ( .A(n24561), .B(n24560), .Z(n24812) );
  NOR U24924 ( .A(n115), .B(n73), .Z(n24813) );
  IV U24925 ( .A(n24813), .Z(n24562) );
  NOR U24926 ( .A(n24812), .B(n24562), .Z(n24815) );
  IV U24927 ( .A(n24563), .Z(n24565) );
  XOR U24928 ( .A(n24565), .B(n24564), .Z(n24808) );
  NOR U24929 ( .A(n82), .B(n73), .Z(n24809) );
  IV U24930 ( .A(n24809), .Z(n24566) );
  NOR U24931 ( .A(n24808), .B(n24566), .Z(n24811) );
  IV U24932 ( .A(n24567), .Z(n24569) );
  XOR U24933 ( .A(n24569), .B(n24568), .Z(n24804) );
  NOR U24934 ( .A(n114), .B(n73), .Z(n24805) );
  IV U24935 ( .A(n24805), .Z(n24570) );
  NOR U24936 ( .A(n24804), .B(n24570), .Z(n24807) );
  IV U24937 ( .A(n24571), .Z(n24573) );
  XOR U24938 ( .A(n24573), .B(n24572), .Z(n24800) );
  NOR U24939 ( .A(n83), .B(n73), .Z(n24801) );
  IV U24940 ( .A(n24801), .Z(n24574) );
  NOR U24941 ( .A(n24800), .B(n24574), .Z(n24803) );
  IV U24942 ( .A(n24575), .Z(n24577) );
  XOR U24943 ( .A(n24577), .B(n24576), .Z(n24796) );
  NOR U24944 ( .A(n113), .B(n73), .Z(n24797) );
  IV U24945 ( .A(n24797), .Z(n24578) );
  NOR U24946 ( .A(n24796), .B(n24578), .Z(n24799) );
  IV U24947 ( .A(n24579), .Z(n24581) );
  XOR U24948 ( .A(n24581), .B(n24580), .Z(n24792) );
  NOR U24949 ( .A(n84), .B(n73), .Z(n24793) );
  IV U24950 ( .A(n24793), .Z(n24582) );
  NOR U24951 ( .A(n24792), .B(n24582), .Z(n24795) );
  IV U24952 ( .A(n24583), .Z(n24585) );
  XOR U24953 ( .A(n24585), .B(n24584), .Z(n24788) );
  NOR U24954 ( .A(n112), .B(n73), .Z(n24789) );
  IV U24955 ( .A(n24789), .Z(n24586) );
  NOR U24956 ( .A(n24788), .B(n24586), .Z(n24791) );
  IV U24957 ( .A(n24587), .Z(n24589) );
  XOR U24958 ( .A(n24589), .B(n24588), .Z(n24784) );
  NOR U24959 ( .A(n85), .B(n73), .Z(n24785) );
  IV U24960 ( .A(n24785), .Z(n24590) );
  NOR U24961 ( .A(n24784), .B(n24590), .Z(n24787) );
  IV U24962 ( .A(n24591), .Z(n24593) );
  XOR U24963 ( .A(n24593), .B(n24592), .Z(n24780) );
  NOR U24964 ( .A(n111), .B(n73), .Z(n24781) );
  IV U24965 ( .A(n24781), .Z(n24594) );
  NOR U24966 ( .A(n24780), .B(n24594), .Z(n24783) );
  IV U24967 ( .A(n24595), .Z(n24597) );
  XOR U24968 ( .A(n24597), .B(n24596), .Z(n24776) );
  NOR U24969 ( .A(n86), .B(n73), .Z(n24777) );
  IV U24970 ( .A(n24777), .Z(n24598) );
  NOR U24971 ( .A(n24776), .B(n24598), .Z(n24779) );
  IV U24972 ( .A(n24599), .Z(n24601) );
  XOR U24973 ( .A(n24601), .B(n24600), .Z(n24772) );
  NOR U24974 ( .A(n110), .B(n73), .Z(n24773) );
  IV U24975 ( .A(n24773), .Z(n24602) );
  NOR U24976 ( .A(n24772), .B(n24602), .Z(n24775) );
  XOR U24977 ( .A(n24604), .B(n24603), .Z(n24768) );
  NOR U24978 ( .A(n109), .B(n73), .Z(n24769) );
  IV U24979 ( .A(n24769), .Z(n24605) );
  NOR U24980 ( .A(n24768), .B(n24605), .Z(n24771) );
  XOR U24981 ( .A(n24607), .B(n24606), .Z(n24756) );
  IV U24982 ( .A(n24756), .Z(n24609) );
  NOR U24983 ( .A(n87), .B(n73), .Z(n24608) );
  IV U24984 ( .A(n24608), .Z(n24757) );
  NOR U24985 ( .A(n24609), .B(n24757), .Z(n24759) );
  IV U24986 ( .A(n24610), .Z(n24612) );
  XOR U24987 ( .A(n24612), .B(n24611), .Z(n24752) );
  NOR U24988 ( .A(n107), .B(n73), .Z(n24753) );
  IV U24989 ( .A(n24753), .Z(n24613) );
  NOR U24990 ( .A(n24752), .B(n24613), .Z(n24755) );
  IV U24991 ( .A(n24614), .Z(n24616) );
  XOR U24992 ( .A(n24616), .B(n24615), .Z(n24748) );
  NOR U24993 ( .A(n88), .B(n73), .Z(n24749) );
  IV U24994 ( .A(n24749), .Z(n24617) );
  NOR U24995 ( .A(n24748), .B(n24617), .Z(n24751) );
  IV U24996 ( .A(n24618), .Z(n24620) );
  XOR U24997 ( .A(n24620), .B(n24619), .Z(n24744) );
  NOR U24998 ( .A(n106), .B(n73), .Z(n24745) );
  IV U24999 ( .A(n24745), .Z(n24621) );
  NOR U25000 ( .A(n24744), .B(n24621), .Z(n24747) );
  IV U25001 ( .A(n24622), .Z(n24624) );
  XOR U25002 ( .A(n24624), .B(n24623), .Z(n24740) );
  NOR U25003 ( .A(n105), .B(n73), .Z(n24741) );
  IV U25004 ( .A(n24741), .Z(n24625) );
  NOR U25005 ( .A(n24740), .B(n24625), .Z(n24743) );
  XOR U25006 ( .A(n24627), .B(n24626), .Z(n24728) );
  IV U25007 ( .A(n24728), .Z(n24629) );
  NOR U25008 ( .A(n89), .B(n73), .Z(n24628) );
  IV U25009 ( .A(n24628), .Z(n24729) );
  NOR U25010 ( .A(n24629), .B(n24729), .Z(n24731) );
  IV U25011 ( .A(n24630), .Z(n24632) );
  XOR U25012 ( .A(n24632), .B(n24631), .Z(n24724) );
  NOR U25013 ( .A(n103), .B(n73), .Z(n24725) );
  IV U25014 ( .A(n24725), .Z(n24633) );
  NOR U25015 ( .A(n24724), .B(n24633), .Z(n24727) );
  IV U25016 ( .A(n24634), .Z(n24636) );
  XOR U25017 ( .A(n24636), .B(n24635), .Z(n24720) );
  NOR U25018 ( .A(n90), .B(n73), .Z(n24721) );
  IV U25019 ( .A(n24721), .Z(n24637) );
  NOR U25020 ( .A(n24720), .B(n24637), .Z(n24723) );
  IV U25021 ( .A(n24638), .Z(n24640) );
  XOR U25022 ( .A(n24640), .B(n24639), .Z(n24716) );
  NOR U25023 ( .A(n102), .B(n73), .Z(n24717) );
  IV U25024 ( .A(n24717), .Z(n24641) );
  NOR U25025 ( .A(n24716), .B(n24641), .Z(n24719) );
  IV U25026 ( .A(n24642), .Z(n24644) );
  XOR U25027 ( .A(n24644), .B(n24643), .Z(n24712) );
  NOR U25028 ( .A(n101), .B(n73), .Z(n24713) );
  IV U25029 ( .A(n24713), .Z(n24645) );
  NOR U25030 ( .A(n24712), .B(n24645), .Z(n24715) );
  IV U25031 ( .A(n24646), .Z(n24648) );
  XOR U25032 ( .A(n24648), .B(n24647), .Z(n24708) );
  NOR U25033 ( .A(n100), .B(n73), .Z(n24709) );
  IV U25034 ( .A(n24709), .Z(n24649) );
  NOR U25035 ( .A(n24708), .B(n24649), .Z(n24711) );
  IV U25036 ( .A(n24650), .Z(n24652) );
  XOR U25037 ( .A(n24652), .B(n24651), .Z(n24704) );
  NOR U25038 ( .A(n99), .B(n73), .Z(n24705) );
  IV U25039 ( .A(n24705), .Z(n24653) );
  NOR U25040 ( .A(n24704), .B(n24653), .Z(n24707) );
  IV U25041 ( .A(n24654), .Z(n24656) );
  XOR U25042 ( .A(n24656), .B(n24655), .Z(n24700) );
  NOR U25043 ( .A(n98), .B(n73), .Z(n24701) );
  IV U25044 ( .A(n24701), .Z(n24657) );
  NOR U25045 ( .A(n24700), .B(n24657), .Z(n24703) );
  XOR U25046 ( .A(n24659), .B(n24658), .Z(n24696) );
  NOR U25047 ( .A(n91), .B(n73), .Z(n24697) );
  IV U25048 ( .A(n24697), .Z(n24660) );
  NOR U25049 ( .A(n24696), .B(n24660), .Z(n24699) );
  IV U25050 ( .A(n24661), .Z(n24663) );
  XOR U25051 ( .A(n24663), .B(n24662), .Z(n24684) );
  NOR U25052 ( .A(n96), .B(n73), .Z(n24685) );
  IV U25053 ( .A(n24685), .Z(n24664) );
  NOR U25054 ( .A(n24684), .B(n24664), .Z(n24687) );
  NOR U25055 ( .A(n95), .B(n73), .Z(n24681) );
  IV U25056 ( .A(n24681), .Z(n24667) );
  XOR U25057 ( .A(n24666), .B(n24665), .Z(n24680) );
  NOR U25058 ( .A(n24667), .B(n24680), .Z(n24683) );
  NOR U25059 ( .A(n93), .B(n73), .Z(n25668) );
  IV U25060 ( .A(n25668), .Z(n24668) );
  NOR U25061 ( .A(n72), .B(n168), .Z(n24676) );
  IV U25062 ( .A(n24676), .Z(n24671) );
  NOR U25063 ( .A(n24668), .B(n24671), .Z(n24669) );
  IV U25064 ( .A(n24669), .Z(n24670) );
  NOR U25065 ( .A(n94), .B(n24670), .Z(n24679) );
  NOR U25066 ( .A(n24671), .B(n93), .Z(n24672) );
  XOR U25067 ( .A(n94), .B(n24672), .Z(n24673) );
  NOR U25068 ( .A(n73), .B(n24673), .Z(n24674) );
  IV U25069 ( .A(n24674), .Z(n25166) );
  XOR U25070 ( .A(n24676), .B(n24675), .Z(n25165) );
  IV U25071 ( .A(n25165), .Z(n24677) );
  NOR U25072 ( .A(n25166), .B(n24677), .Z(n24678) );
  NOR U25073 ( .A(n24679), .B(n24678), .Z(n25162) );
  XOR U25074 ( .A(n24681), .B(n24680), .Z(n25161) );
  NOR U25075 ( .A(n25162), .B(n25161), .Z(n24682) );
  NOR U25076 ( .A(n24683), .B(n24682), .Z(n25189) );
  XOR U25077 ( .A(n24685), .B(n24684), .Z(n25190) );
  NOR U25078 ( .A(n25189), .B(n25190), .Z(n24686) );
  NOR U25079 ( .A(n24687), .B(n24686), .Z(n24692) );
  XOR U25080 ( .A(n24689), .B(n24688), .Z(n24691) );
  IV U25081 ( .A(n24691), .Z(n24690) );
  NOR U25082 ( .A(n24692), .B(n24690), .Z(n24695) );
  XOR U25083 ( .A(n24692), .B(n24691), .Z(n25158) );
  NOR U25084 ( .A(n97), .B(n73), .Z(n25159) );
  IV U25085 ( .A(n25159), .Z(n24693) );
  NOR U25086 ( .A(n25158), .B(n24693), .Z(n24694) );
  NOR U25087 ( .A(n24695), .B(n24694), .Z(n25154) );
  XOR U25088 ( .A(n24697), .B(n24696), .Z(n25155) );
  NOR U25089 ( .A(n25154), .B(n25155), .Z(n24698) );
  NOR U25090 ( .A(n24699), .B(n24698), .Z(n25150) );
  XOR U25091 ( .A(n24701), .B(n24700), .Z(n25151) );
  NOR U25092 ( .A(n25150), .B(n25151), .Z(n24702) );
  NOR U25093 ( .A(n24703), .B(n24702), .Z(n25146) );
  XOR U25094 ( .A(n24705), .B(n24704), .Z(n25147) );
  NOR U25095 ( .A(n25146), .B(n25147), .Z(n24706) );
  NOR U25096 ( .A(n24707), .B(n24706), .Z(n25142) );
  XOR U25097 ( .A(n24709), .B(n24708), .Z(n25143) );
  NOR U25098 ( .A(n25142), .B(n25143), .Z(n24710) );
  NOR U25099 ( .A(n24711), .B(n24710), .Z(n25138) );
  XOR U25100 ( .A(n24713), .B(n24712), .Z(n25139) );
  NOR U25101 ( .A(n25138), .B(n25139), .Z(n24714) );
  NOR U25102 ( .A(n24715), .B(n24714), .Z(n25134) );
  XOR U25103 ( .A(n24717), .B(n24716), .Z(n25135) );
  NOR U25104 ( .A(n25134), .B(n25135), .Z(n24718) );
  NOR U25105 ( .A(n24719), .B(n24718), .Z(n25130) );
  XOR U25106 ( .A(n24721), .B(n24720), .Z(n25131) );
  NOR U25107 ( .A(n25130), .B(n25131), .Z(n24722) );
  NOR U25108 ( .A(n24723), .B(n24722), .Z(n25127) );
  XOR U25109 ( .A(n24725), .B(n24724), .Z(n25126) );
  NOR U25110 ( .A(n25127), .B(n25126), .Z(n24726) );
  NOR U25111 ( .A(n24727), .B(n24726), .Z(n25233) );
  XOR U25112 ( .A(n24729), .B(n24728), .Z(n25232) );
  NOR U25113 ( .A(n25233), .B(n25232), .Z(n24730) );
  NOR U25114 ( .A(n24731), .B(n24730), .Z(n24736) );
  XOR U25115 ( .A(n24733), .B(n24732), .Z(n24735) );
  IV U25116 ( .A(n24735), .Z(n24734) );
  NOR U25117 ( .A(n24736), .B(n24734), .Z(n24739) );
  XOR U25118 ( .A(n24736), .B(n24735), .Z(n25123) );
  NOR U25119 ( .A(n104), .B(n73), .Z(n25124) );
  IV U25120 ( .A(n25124), .Z(n24737) );
  NOR U25121 ( .A(n25123), .B(n24737), .Z(n24738) );
  NOR U25122 ( .A(n24739), .B(n24738), .Z(n25119) );
  XOR U25123 ( .A(n24741), .B(n24740), .Z(n25120) );
  NOR U25124 ( .A(n25119), .B(n25120), .Z(n24742) );
  NOR U25125 ( .A(n24743), .B(n24742), .Z(n25115) );
  XOR U25126 ( .A(n24745), .B(n24744), .Z(n25116) );
  NOR U25127 ( .A(n25115), .B(n25116), .Z(n24746) );
  NOR U25128 ( .A(n24747), .B(n24746), .Z(n25111) );
  XOR U25129 ( .A(n24749), .B(n24748), .Z(n25112) );
  NOR U25130 ( .A(n25111), .B(n25112), .Z(n24750) );
  NOR U25131 ( .A(n24751), .B(n24750), .Z(n25108) );
  XOR U25132 ( .A(n24753), .B(n24752), .Z(n25107) );
  NOR U25133 ( .A(n25108), .B(n25107), .Z(n24754) );
  NOR U25134 ( .A(n24755), .B(n24754), .Z(n25261) );
  XOR U25135 ( .A(n24757), .B(n24756), .Z(n25260) );
  NOR U25136 ( .A(n25261), .B(n25260), .Z(n24758) );
  NOR U25137 ( .A(n24759), .B(n24758), .Z(n24764) );
  XOR U25138 ( .A(n24761), .B(n24760), .Z(n24763) );
  IV U25139 ( .A(n24763), .Z(n24762) );
  NOR U25140 ( .A(n24764), .B(n24762), .Z(n24767) );
  XOR U25141 ( .A(n24764), .B(n24763), .Z(n25104) );
  NOR U25142 ( .A(n108), .B(n73), .Z(n25105) );
  IV U25143 ( .A(n25105), .Z(n24765) );
  NOR U25144 ( .A(n25104), .B(n24765), .Z(n24766) );
  NOR U25145 ( .A(n24767), .B(n24766), .Z(n25100) );
  XOR U25146 ( .A(n24769), .B(n24768), .Z(n25101) );
  NOR U25147 ( .A(n25100), .B(n25101), .Z(n24770) );
  NOR U25148 ( .A(n24771), .B(n24770), .Z(n25096) );
  XOR U25149 ( .A(n24773), .B(n24772), .Z(n25097) );
  NOR U25150 ( .A(n25096), .B(n25097), .Z(n24774) );
  NOR U25151 ( .A(n24775), .B(n24774), .Z(n25092) );
  XOR U25152 ( .A(n24777), .B(n24776), .Z(n25093) );
  NOR U25153 ( .A(n25092), .B(n25093), .Z(n24778) );
  NOR U25154 ( .A(n24779), .B(n24778), .Z(n25088) );
  XOR U25155 ( .A(n24781), .B(n24780), .Z(n25089) );
  NOR U25156 ( .A(n25088), .B(n25089), .Z(n24782) );
  NOR U25157 ( .A(n24783), .B(n24782), .Z(n25084) );
  XOR U25158 ( .A(n24785), .B(n24784), .Z(n25085) );
  NOR U25159 ( .A(n25084), .B(n25085), .Z(n24786) );
  NOR U25160 ( .A(n24787), .B(n24786), .Z(n25080) );
  XOR U25161 ( .A(n24789), .B(n24788), .Z(n25081) );
  NOR U25162 ( .A(n25080), .B(n25081), .Z(n24790) );
  NOR U25163 ( .A(n24791), .B(n24790), .Z(n25076) );
  XOR U25164 ( .A(n24793), .B(n24792), .Z(n25077) );
  NOR U25165 ( .A(n25076), .B(n25077), .Z(n24794) );
  NOR U25166 ( .A(n24795), .B(n24794), .Z(n25072) );
  XOR U25167 ( .A(n24797), .B(n24796), .Z(n25073) );
  NOR U25168 ( .A(n25072), .B(n25073), .Z(n24798) );
  NOR U25169 ( .A(n24799), .B(n24798), .Z(n25068) );
  XOR U25170 ( .A(n24801), .B(n24800), .Z(n25069) );
  NOR U25171 ( .A(n25068), .B(n25069), .Z(n24802) );
  NOR U25172 ( .A(n24803), .B(n24802), .Z(n25064) );
  XOR U25173 ( .A(n24805), .B(n24804), .Z(n25065) );
  NOR U25174 ( .A(n25064), .B(n25065), .Z(n24806) );
  NOR U25175 ( .A(n24807), .B(n24806), .Z(n25060) );
  XOR U25176 ( .A(n24809), .B(n24808), .Z(n25061) );
  NOR U25177 ( .A(n25060), .B(n25061), .Z(n24810) );
  NOR U25178 ( .A(n24811), .B(n24810), .Z(n25056) );
  XOR U25179 ( .A(n24813), .B(n24812), .Z(n25057) );
  NOR U25180 ( .A(n25056), .B(n25057), .Z(n24814) );
  NOR U25181 ( .A(n24815), .B(n24814), .Z(n25052) );
  XOR U25182 ( .A(n24817), .B(n24816), .Z(n25053) );
  NOR U25183 ( .A(n25052), .B(n25053), .Z(n24818) );
  NOR U25184 ( .A(n24819), .B(n24818), .Z(n25048) );
  XOR U25185 ( .A(n24821), .B(n24820), .Z(n25049) );
  NOR U25186 ( .A(n25048), .B(n25049), .Z(n24822) );
  NOR U25187 ( .A(n24823), .B(n24822), .Z(n24824) );
  IV U25188 ( .A(n24824), .Z(n25046) );
  XOR U25189 ( .A(n24826), .B(n24825), .Z(n24827) );
  IV U25190 ( .A(n24827), .Z(n25045) );
  NOR U25191 ( .A(n25046), .B(n25045), .Z(n24828) );
  NOR U25192 ( .A(n24829), .B(n24828), .Z(n24830) );
  IV U25193 ( .A(n24830), .Z(n25044) );
  XOR U25194 ( .A(n24832), .B(n24831), .Z(n25043) );
  NOR U25195 ( .A(n25044), .B(n25043), .Z(n24833) );
  NOR U25196 ( .A(n24834), .B(n24833), .Z(n24835) );
  IV U25197 ( .A(n24835), .Z(n25041) );
  XOR U25198 ( .A(n24837), .B(n24836), .Z(n24838) );
  IV U25199 ( .A(n24838), .Z(n25040) );
  NOR U25200 ( .A(n25041), .B(n25040), .Z(n24839) );
  NOR U25201 ( .A(n24840), .B(n24839), .Z(n24841) );
  IV U25202 ( .A(n24841), .Z(n25036) );
  XOR U25203 ( .A(n24843), .B(n24842), .Z(n25035) );
  NOR U25204 ( .A(n25036), .B(n25035), .Z(n24844) );
  NOR U25205 ( .A(n24845), .B(n24844), .Z(n24846) );
  IV U25206 ( .A(n24846), .Z(n25033) );
  XOR U25207 ( .A(n24848), .B(n24847), .Z(n24849) );
  IV U25208 ( .A(n24849), .Z(n25032) );
  NOR U25209 ( .A(n25033), .B(n25032), .Z(n24850) );
  NOR U25210 ( .A(n24851), .B(n24850), .Z(n24852) );
  IV U25211 ( .A(n24852), .Z(n25031) );
  XOR U25212 ( .A(n24854), .B(n24853), .Z(n25030) );
  NOR U25213 ( .A(n25031), .B(n25030), .Z(n24855) );
  NOR U25214 ( .A(n24856), .B(n24855), .Z(n24857) );
  IV U25215 ( .A(n24857), .Z(n25028) );
  XOR U25216 ( .A(n24859), .B(n24858), .Z(n24860) );
  IV U25217 ( .A(n24860), .Z(n25027) );
  NOR U25218 ( .A(n25028), .B(n25027), .Z(n24861) );
  NOR U25219 ( .A(n24862), .B(n24861), .Z(n24863) );
  IV U25220 ( .A(n24863), .Z(n25026) );
  XOR U25221 ( .A(n24865), .B(n24864), .Z(n25025) );
  NOR U25222 ( .A(n25026), .B(n25025), .Z(n24866) );
  NOR U25223 ( .A(n24867), .B(n24866), .Z(n24868) );
  IV U25224 ( .A(n24868), .Z(n25023) );
  XOR U25225 ( .A(n24870), .B(n24869), .Z(n24871) );
  IV U25226 ( .A(n24871), .Z(n25022) );
  NOR U25227 ( .A(n25023), .B(n25022), .Z(n24872) );
  NOR U25228 ( .A(n24873), .B(n24872), .Z(n24874) );
  IV U25229 ( .A(n24874), .Z(n25021) );
  XOR U25230 ( .A(n24876), .B(n24875), .Z(n25020) );
  NOR U25231 ( .A(n25021), .B(n25020), .Z(n24877) );
  NOR U25232 ( .A(n24878), .B(n24877), .Z(n24879) );
  IV U25233 ( .A(n24879), .Z(n25018) );
  XOR U25234 ( .A(n24881), .B(n24880), .Z(n24882) );
  IV U25235 ( .A(n24882), .Z(n25017) );
  NOR U25236 ( .A(n25018), .B(n25017), .Z(n24883) );
  NOR U25237 ( .A(n24884), .B(n24883), .Z(n25015) );
  IV U25238 ( .A(n25015), .Z(n24885) );
  NOR U25239 ( .A(n25014), .B(n24885), .Z(n24886) );
  NOR U25240 ( .A(n24887), .B(n24886), .Z(n25010) );
  XOR U25241 ( .A(n24889), .B(n24888), .Z(n25011) );
  NOR U25242 ( .A(n25010), .B(n25011), .Z(n24890) );
  NOR U25243 ( .A(n24891), .B(n24890), .Z(n25006) );
  XOR U25244 ( .A(n24893), .B(n24892), .Z(n25007) );
  NOR U25245 ( .A(n25006), .B(n25007), .Z(n24894) );
  NOR U25246 ( .A(n24895), .B(n24894), .Z(n25002) );
  XOR U25247 ( .A(n24897), .B(n24896), .Z(n25003) );
  NOR U25248 ( .A(n25002), .B(n25003), .Z(n24898) );
  NOR U25249 ( .A(n24899), .B(n24898), .Z(n24904) );
  XOR U25250 ( .A(n24901), .B(n24900), .Z(n24903) );
  IV U25251 ( .A(n24903), .Z(n24902) );
  NOR U25252 ( .A(n24904), .B(n24902), .Z(n24907) );
  XOR U25253 ( .A(n24904), .B(n24903), .Z(n24999) );
  NOR U25254 ( .A(n143), .B(n73), .Z(n25000) );
  IV U25255 ( .A(n25000), .Z(n24905) );
  NOR U25256 ( .A(n24999), .B(n24905), .Z(n24906) );
  NOR U25257 ( .A(n24907), .B(n24906), .Z(n24995) );
  XOR U25258 ( .A(n24909), .B(n24908), .Z(n24996) );
  NOR U25259 ( .A(n24995), .B(n24996), .Z(n24910) );
  NOR U25260 ( .A(n24911), .B(n24910), .Z(n24992) );
  XOR U25261 ( .A(n24913), .B(n24912), .Z(n24991) );
  NOR U25262 ( .A(n24992), .B(n24991), .Z(n24914) );
  NOR U25263 ( .A(n24915), .B(n24914), .Z(n24916) );
  IV U25264 ( .A(n24916), .Z(n25412) );
  NOR U25265 ( .A(n24917), .B(n25412), .Z(n24918) );
  NOR U25266 ( .A(n24919), .B(n24918), .Z(n24920) );
  IV U25267 ( .A(n24920), .Z(n24923) );
  NOR U25268 ( .A(n150), .B(n73), .Z(n24922) );
  IV U25269 ( .A(n24922), .Z(n24921) );
  NOR U25270 ( .A(n24923), .B(n24921), .Z(n24928) );
  XOR U25271 ( .A(n24923), .B(n24922), .Z(n24990) );
  XOR U25272 ( .A(n24925), .B(n24924), .Z(n24926) );
  IV U25273 ( .A(n24926), .Z(n24989) );
  NOR U25274 ( .A(n24990), .B(n24989), .Z(n24927) );
  NOR U25275 ( .A(n24928), .B(n24927), .Z(n25431) );
  NOR U25276 ( .A(n24929), .B(n25431), .Z(n24930) );
  NOR U25277 ( .A(n24931), .B(n24930), .Z(n24936) );
  IV U25278 ( .A(n24936), .Z(n24932) );
  NOR U25279 ( .A(n24935), .B(n24932), .Z(n24938) );
  XOR U25280 ( .A(n24934), .B(n24933), .Z(n24986) );
  XOR U25281 ( .A(n24936), .B(n24935), .Z(n24985) );
  NOR U25282 ( .A(n24986), .B(n24985), .Z(n24937) );
  NOR U25283 ( .A(n24938), .B(n24937), .Z(n24944) );
  IV U25284 ( .A(n24944), .Z(n24940) );
  NOR U25285 ( .A(n156), .B(n73), .Z(n24939) );
  IV U25286 ( .A(n24939), .Z(n24943) );
  NOR U25287 ( .A(n24940), .B(n24943), .Z(n24946) );
  XOR U25288 ( .A(n24942), .B(n24941), .Z(n25440) );
  XOR U25289 ( .A(n24944), .B(n24943), .Z(n25441) );
  NOR U25290 ( .A(n25440), .B(n25441), .Z(n24945) );
  NOR U25291 ( .A(n24946), .B(n24945), .Z(n24952) );
  XOR U25292 ( .A(n24948), .B(n24947), .Z(n24949) );
  XOR U25293 ( .A(n24950), .B(n24949), .Z(n24951) );
  NOR U25294 ( .A(n24952), .B(n24951), .Z(n24956) );
  IV U25295 ( .A(n24951), .Z(n24953) );
  XOR U25296 ( .A(n24953), .B(n24952), .Z(n25448) );
  NOR U25297 ( .A(n158), .B(n73), .Z(n24954) );
  IV U25298 ( .A(n24954), .Z(n25449) );
  NOR U25299 ( .A(n25448), .B(n25449), .Z(n24955) );
  NOR U25300 ( .A(n24956), .B(n24955), .Z(n25460) );
  XOR U25301 ( .A(n24958), .B(n24957), .Z(n25459) );
  NOR U25302 ( .A(n25460), .B(n25459), .Z(n24959) );
  NOR U25303 ( .A(n24960), .B(n24959), .Z(n24965) );
  NOR U25304 ( .A(n163), .B(n73), .Z(n24964) );
  IV U25305 ( .A(n24964), .Z(n24961) );
  NOR U25306 ( .A(n24965), .B(n24961), .Z(n24967) );
  XOR U25307 ( .A(n24963), .B(n24962), .Z(n25465) );
  XOR U25308 ( .A(n24965), .B(n24964), .Z(n25464) );
  NOR U25309 ( .A(n25465), .B(n25464), .Z(n24966) );
  NOR U25310 ( .A(n24967), .B(n24966), .Z(n24971) );
  XOR U25311 ( .A(n24969), .B(n24968), .Z(n24970) );
  NOR U25312 ( .A(n24971), .B(n24970), .Z(n24975) );
  XOR U25313 ( .A(n24971), .B(n24970), .Z(n25971) );
  IV U25314 ( .A(n25971), .Z(n24973) );
  NOR U25315 ( .A(n165), .B(n73), .Z(n24972) );
  IV U25316 ( .A(n24972), .Z(n25972) );
  NOR U25317 ( .A(n24973), .B(n25972), .Z(n24974) );
  NOR U25318 ( .A(n24975), .B(n24974), .Z(n25982) );
  XOR U25319 ( .A(n24977), .B(n24976), .Z(n25981) );
  NOR U25320 ( .A(n25982), .B(n25981), .Z(n24978) );
  NOR U25321 ( .A(n24979), .B(n24978), .Z(n24984) );
  XOR U25322 ( .A(n24981), .B(n24980), .Z(n24983) );
  NOR U25323 ( .A(n24984), .B(n24983), .Z(n31501) );
  IV U25324 ( .A(n31501), .Z(n31491) );
  NOR U25325 ( .A(n24982), .B(n31491), .Z(n25991) );
  XOR U25326 ( .A(n24984), .B(n24983), .Z(n31488) );
  IV U25327 ( .A(n31488), .Z(n25987) );
  NOR U25328 ( .A(n165), .B(n74), .Z(n25966) );
  NOR U25329 ( .A(n161), .B(n74), .Z(n25450) );
  XOR U25330 ( .A(n24986), .B(n24985), .Z(n25437) );
  NOR U25331 ( .A(n156), .B(n74), .Z(n25436) );
  IV U25332 ( .A(n25436), .Z(n24987) );
  NOR U25333 ( .A(n25437), .B(n24987), .Z(n25439) );
  NOR U25334 ( .A(n155), .B(n74), .Z(n24988) );
  IV U25335 ( .A(n24988), .Z(n25433) );
  XOR U25336 ( .A(n24990), .B(n24989), .Z(n25422) );
  NOR U25337 ( .A(n153), .B(n74), .Z(n25423) );
  NOR U25338 ( .A(n25422), .B(n25423), .Z(n25426) );
  XOR U25339 ( .A(n24992), .B(n24991), .Z(n25479) );
  IV U25340 ( .A(n25479), .Z(n24994) );
  NOR U25341 ( .A(n148), .B(n74), .Z(n25482) );
  IV U25342 ( .A(n25482), .Z(n24993) );
  NOR U25343 ( .A(n24994), .B(n24993), .Z(n25410) );
  IV U25344 ( .A(n24995), .Z(n24997) );
  XOR U25345 ( .A(n24997), .B(n24996), .Z(n25404) );
  NOR U25346 ( .A(n147), .B(n74), .Z(n25405) );
  IV U25347 ( .A(n25405), .Z(n24998) );
  NOR U25348 ( .A(n25404), .B(n24998), .Z(n25407) );
  XOR U25349 ( .A(n25000), .B(n24999), .Z(n25400) );
  NOR U25350 ( .A(n145), .B(n74), .Z(n25401) );
  IV U25351 ( .A(n25401), .Z(n25001) );
  NOR U25352 ( .A(n25400), .B(n25001), .Z(n25403) );
  IV U25353 ( .A(n25002), .Z(n25004) );
  XOR U25354 ( .A(n25004), .B(n25003), .Z(n25396) );
  NOR U25355 ( .A(n143), .B(n74), .Z(n25397) );
  IV U25356 ( .A(n25397), .Z(n25005) );
  NOR U25357 ( .A(n25396), .B(n25005), .Z(n25399) );
  IV U25358 ( .A(n25006), .Z(n25008) );
  XOR U25359 ( .A(n25008), .B(n25007), .Z(n25392) );
  NOR U25360 ( .A(n141), .B(n74), .Z(n25393) );
  IV U25361 ( .A(n25393), .Z(n25009) );
  NOR U25362 ( .A(n25392), .B(n25009), .Z(n25395) );
  IV U25363 ( .A(n25010), .Z(n25012) );
  XOR U25364 ( .A(n25012), .B(n25011), .Z(n25388) );
  NOR U25365 ( .A(n139), .B(n74), .Z(n25389) );
  IV U25366 ( .A(n25389), .Z(n25013) );
  NOR U25367 ( .A(n25388), .B(n25013), .Z(n25391) );
  XOR U25368 ( .A(n25015), .B(n25014), .Z(n25384) );
  NOR U25369 ( .A(n137), .B(n74), .Z(n25385) );
  IV U25370 ( .A(n25385), .Z(n25016) );
  NOR U25371 ( .A(n25384), .B(n25016), .Z(n25387) );
  XOR U25372 ( .A(n25018), .B(n25017), .Z(n25381) );
  NOR U25373 ( .A(n135), .B(n74), .Z(n25380) );
  IV U25374 ( .A(n25380), .Z(n25019) );
  NOR U25375 ( .A(n25381), .B(n25019), .Z(n25383) );
  NOR U25376 ( .A(n133), .B(n74), .Z(n25375) );
  XOR U25377 ( .A(n25021), .B(n25020), .Z(n25374) );
  NOR U25378 ( .A(n25375), .B(n25374), .Z(n25378) );
  XOR U25379 ( .A(n25023), .B(n25022), .Z(n25370) );
  NOR U25380 ( .A(n131), .B(n74), .Z(n25369) );
  IV U25381 ( .A(n25369), .Z(n25024) );
  NOR U25382 ( .A(n25370), .B(n25024), .Z(n25372) );
  NOR U25383 ( .A(n128), .B(n74), .Z(n25364) );
  XOR U25384 ( .A(n25026), .B(n25025), .Z(n25363) );
  NOR U25385 ( .A(n25364), .B(n25363), .Z(n25367) );
  XOR U25386 ( .A(n25028), .B(n25027), .Z(n25359) );
  NOR U25387 ( .A(n126), .B(n74), .Z(n25358) );
  IV U25388 ( .A(n25358), .Z(n25029) );
  NOR U25389 ( .A(n25359), .B(n25029), .Z(n25361) );
  NOR U25390 ( .A(n125), .B(n74), .Z(n25353) );
  XOR U25391 ( .A(n25031), .B(n25030), .Z(n25352) );
  NOR U25392 ( .A(n25353), .B(n25352), .Z(n25356) );
  XOR U25393 ( .A(n25033), .B(n25032), .Z(n25348) );
  NOR U25394 ( .A(n123), .B(n74), .Z(n25347) );
  IV U25395 ( .A(n25347), .Z(n25034) );
  NOR U25396 ( .A(n25348), .B(n25034), .Z(n25350) );
  NOR U25397 ( .A(n120), .B(n74), .Z(n25038) );
  XOR U25398 ( .A(n25036), .B(n25035), .Z(n25037) );
  NOR U25399 ( .A(n25038), .B(n25037), .Z(n25345) );
  XOR U25400 ( .A(n25038), .B(n25037), .Z(n25039) );
  IV U25401 ( .A(n25039), .Z(n25528) );
  XOR U25402 ( .A(n25041), .B(n25040), .Z(n25340) );
  NOR U25403 ( .A(n119), .B(n74), .Z(n25339) );
  IV U25404 ( .A(n25339), .Z(n25042) );
  NOR U25405 ( .A(n25340), .B(n25042), .Z(n25342) );
  NOR U25406 ( .A(n79), .B(n74), .Z(n25334) );
  XOR U25407 ( .A(n25044), .B(n25043), .Z(n25333) );
  NOR U25408 ( .A(n25334), .B(n25333), .Z(n25337) );
  XOR U25409 ( .A(n25046), .B(n25045), .Z(n25329) );
  NOR U25410 ( .A(n117), .B(n74), .Z(n25328) );
  IV U25411 ( .A(n25328), .Z(n25047) );
  NOR U25412 ( .A(n25329), .B(n25047), .Z(n25331) );
  IV U25413 ( .A(n25048), .Z(n25050) );
  XOR U25414 ( .A(n25050), .B(n25049), .Z(n25324) );
  NOR U25415 ( .A(n80), .B(n74), .Z(n25325) );
  IV U25416 ( .A(n25325), .Z(n25051) );
  NOR U25417 ( .A(n25324), .B(n25051), .Z(n25327) );
  IV U25418 ( .A(n25052), .Z(n25054) );
  XOR U25419 ( .A(n25054), .B(n25053), .Z(n25320) );
  NOR U25420 ( .A(n116), .B(n74), .Z(n25321) );
  IV U25421 ( .A(n25321), .Z(n25055) );
  NOR U25422 ( .A(n25320), .B(n25055), .Z(n25323) );
  IV U25423 ( .A(n25056), .Z(n25058) );
  XOR U25424 ( .A(n25058), .B(n25057), .Z(n25316) );
  NOR U25425 ( .A(n81), .B(n74), .Z(n25317) );
  IV U25426 ( .A(n25317), .Z(n25059) );
  NOR U25427 ( .A(n25316), .B(n25059), .Z(n25319) );
  IV U25428 ( .A(n25060), .Z(n25062) );
  XOR U25429 ( .A(n25062), .B(n25061), .Z(n25312) );
  NOR U25430 ( .A(n115), .B(n74), .Z(n25313) );
  IV U25431 ( .A(n25313), .Z(n25063) );
  NOR U25432 ( .A(n25312), .B(n25063), .Z(n25315) );
  IV U25433 ( .A(n25064), .Z(n25066) );
  XOR U25434 ( .A(n25066), .B(n25065), .Z(n25308) );
  NOR U25435 ( .A(n82), .B(n74), .Z(n25309) );
  IV U25436 ( .A(n25309), .Z(n25067) );
  NOR U25437 ( .A(n25308), .B(n25067), .Z(n25311) );
  IV U25438 ( .A(n25068), .Z(n25070) );
  XOR U25439 ( .A(n25070), .B(n25069), .Z(n25304) );
  NOR U25440 ( .A(n114), .B(n74), .Z(n25305) );
  IV U25441 ( .A(n25305), .Z(n25071) );
  NOR U25442 ( .A(n25304), .B(n25071), .Z(n25307) );
  IV U25443 ( .A(n25072), .Z(n25074) );
  XOR U25444 ( .A(n25074), .B(n25073), .Z(n25300) );
  NOR U25445 ( .A(n83), .B(n74), .Z(n25301) );
  IV U25446 ( .A(n25301), .Z(n25075) );
  NOR U25447 ( .A(n25300), .B(n25075), .Z(n25303) );
  IV U25448 ( .A(n25076), .Z(n25078) );
  XOR U25449 ( .A(n25078), .B(n25077), .Z(n25296) );
  NOR U25450 ( .A(n113), .B(n74), .Z(n25297) );
  IV U25451 ( .A(n25297), .Z(n25079) );
  NOR U25452 ( .A(n25296), .B(n25079), .Z(n25299) );
  IV U25453 ( .A(n25080), .Z(n25082) );
  XOR U25454 ( .A(n25082), .B(n25081), .Z(n25292) );
  NOR U25455 ( .A(n84), .B(n74), .Z(n25293) );
  IV U25456 ( .A(n25293), .Z(n25083) );
  NOR U25457 ( .A(n25292), .B(n25083), .Z(n25295) );
  IV U25458 ( .A(n25084), .Z(n25086) );
  XOR U25459 ( .A(n25086), .B(n25085), .Z(n25288) );
  NOR U25460 ( .A(n112), .B(n74), .Z(n25289) );
  IV U25461 ( .A(n25289), .Z(n25087) );
  NOR U25462 ( .A(n25288), .B(n25087), .Z(n25291) );
  IV U25463 ( .A(n25088), .Z(n25090) );
  XOR U25464 ( .A(n25090), .B(n25089), .Z(n25284) );
  NOR U25465 ( .A(n85), .B(n74), .Z(n25285) );
  IV U25466 ( .A(n25285), .Z(n25091) );
  NOR U25467 ( .A(n25284), .B(n25091), .Z(n25287) );
  IV U25468 ( .A(n25092), .Z(n25094) );
  XOR U25469 ( .A(n25094), .B(n25093), .Z(n25280) );
  NOR U25470 ( .A(n111), .B(n74), .Z(n25281) );
  IV U25471 ( .A(n25281), .Z(n25095) );
  NOR U25472 ( .A(n25280), .B(n25095), .Z(n25283) );
  IV U25473 ( .A(n25096), .Z(n25098) );
  XOR U25474 ( .A(n25098), .B(n25097), .Z(n25276) );
  NOR U25475 ( .A(n86), .B(n74), .Z(n25277) );
  IV U25476 ( .A(n25277), .Z(n25099) );
  NOR U25477 ( .A(n25276), .B(n25099), .Z(n25279) );
  IV U25478 ( .A(n25100), .Z(n25102) );
  XOR U25479 ( .A(n25102), .B(n25101), .Z(n25272) );
  NOR U25480 ( .A(n110), .B(n74), .Z(n25273) );
  IV U25481 ( .A(n25273), .Z(n25103) );
  NOR U25482 ( .A(n25272), .B(n25103), .Z(n25275) );
  XOR U25483 ( .A(n25105), .B(n25104), .Z(n25268) );
  NOR U25484 ( .A(n109), .B(n74), .Z(n25269) );
  IV U25485 ( .A(n25269), .Z(n25106) );
  NOR U25486 ( .A(n25268), .B(n25106), .Z(n25271) );
  XOR U25487 ( .A(n25108), .B(n25107), .Z(n25256) );
  IV U25488 ( .A(n25256), .Z(n25110) );
  NOR U25489 ( .A(n87), .B(n74), .Z(n25109) );
  IV U25490 ( .A(n25109), .Z(n25257) );
  NOR U25491 ( .A(n25110), .B(n25257), .Z(n25259) );
  IV U25492 ( .A(n25111), .Z(n25113) );
  XOR U25493 ( .A(n25113), .B(n25112), .Z(n25252) );
  NOR U25494 ( .A(n107), .B(n74), .Z(n25253) );
  IV U25495 ( .A(n25253), .Z(n25114) );
  NOR U25496 ( .A(n25252), .B(n25114), .Z(n25255) );
  IV U25497 ( .A(n25115), .Z(n25117) );
  XOR U25498 ( .A(n25117), .B(n25116), .Z(n25248) );
  NOR U25499 ( .A(n88), .B(n74), .Z(n25249) );
  IV U25500 ( .A(n25249), .Z(n25118) );
  NOR U25501 ( .A(n25248), .B(n25118), .Z(n25251) );
  IV U25502 ( .A(n25119), .Z(n25121) );
  XOR U25503 ( .A(n25121), .B(n25120), .Z(n25244) );
  NOR U25504 ( .A(n106), .B(n74), .Z(n25245) );
  IV U25505 ( .A(n25245), .Z(n25122) );
  NOR U25506 ( .A(n25244), .B(n25122), .Z(n25247) );
  XOR U25507 ( .A(n25124), .B(n25123), .Z(n25240) );
  NOR U25508 ( .A(n105), .B(n74), .Z(n25241) );
  IV U25509 ( .A(n25241), .Z(n25125) );
  NOR U25510 ( .A(n25240), .B(n25125), .Z(n25243) );
  XOR U25511 ( .A(n25127), .B(n25126), .Z(n25228) );
  IV U25512 ( .A(n25228), .Z(n25129) );
  NOR U25513 ( .A(n89), .B(n74), .Z(n25128) );
  IV U25514 ( .A(n25128), .Z(n25229) );
  NOR U25515 ( .A(n25129), .B(n25229), .Z(n25231) );
  IV U25516 ( .A(n25130), .Z(n25132) );
  XOR U25517 ( .A(n25132), .B(n25131), .Z(n25224) );
  NOR U25518 ( .A(n103), .B(n74), .Z(n25225) );
  IV U25519 ( .A(n25225), .Z(n25133) );
  NOR U25520 ( .A(n25224), .B(n25133), .Z(n25227) );
  IV U25521 ( .A(n25134), .Z(n25136) );
  XOR U25522 ( .A(n25136), .B(n25135), .Z(n25220) );
  NOR U25523 ( .A(n90), .B(n74), .Z(n25221) );
  IV U25524 ( .A(n25221), .Z(n25137) );
  NOR U25525 ( .A(n25220), .B(n25137), .Z(n25223) );
  IV U25526 ( .A(n25138), .Z(n25140) );
  XOR U25527 ( .A(n25140), .B(n25139), .Z(n25216) );
  NOR U25528 ( .A(n102), .B(n74), .Z(n25217) );
  IV U25529 ( .A(n25217), .Z(n25141) );
  NOR U25530 ( .A(n25216), .B(n25141), .Z(n25219) );
  IV U25531 ( .A(n25142), .Z(n25144) );
  XOR U25532 ( .A(n25144), .B(n25143), .Z(n25212) );
  NOR U25533 ( .A(n101), .B(n74), .Z(n25213) );
  IV U25534 ( .A(n25213), .Z(n25145) );
  NOR U25535 ( .A(n25212), .B(n25145), .Z(n25215) );
  IV U25536 ( .A(n25146), .Z(n25148) );
  XOR U25537 ( .A(n25148), .B(n25147), .Z(n25208) );
  NOR U25538 ( .A(n100), .B(n74), .Z(n25209) );
  IV U25539 ( .A(n25209), .Z(n25149) );
  NOR U25540 ( .A(n25208), .B(n25149), .Z(n25211) );
  IV U25541 ( .A(n25150), .Z(n25152) );
  XOR U25542 ( .A(n25152), .B(n25151), .Z(n25204) );
  NOR U25543 ( .A(n99), .B(n74), .Z(n25205) );
  IV U25544 ( .A(n25205), .Z(n25153) );
  NOR U25545 ( .A(n25204), .B(n25153), .Z(n25207) );
  IV U25546 ( .A(n25154), .Z(n25156) );
  XOR U25547 ( .A(n25156), .B(n25155), .Z(n25200) );
  NOR U25548 ( .A(n98), .B(n74), .Z(n25201) );
  IV U25549 ( .A(n25201), .Z(n25157) );
  NOR U25550 ( .A(n25200), .B(n25157), .Z(n25203) );
  XOR U25551 ( .A(n25159), .B(n25158), .Z(n25196) );
  NOR U25552 ( .A(n91), .B(n74), .Z(n25197) );
  IV U25553 ( .A(n25197), .Z(n25160) );
  NOR U25554 ( .A(n25196), .B(n25160), .Z(n25199) );
  XOR U25555 ( .A(n25162), .B(n25161), .Z(n25184) );
  IV U25556 ( .A(n25184), .Z(n25164) );
  NOR U25557 ( .A(n96), .B(n74), .Z(n25163) );
  IV U25558 ( .A(n25163), .Z(n25185) );
  NOR U25559 ( .A(n25164), .B(n25185), .Z(n25187) );
  NOR U25560 ( .A(n95), .B(n74), .Z(n25181) );
  IV U25561 ( .A(n25181), .Z(n25167) );
  XOR U25562 ( .A(n25166), .B(n25165), .Z(n25180) );
  NOR U25563 ( .A(n25167), .B(n25180), .Z(n25183) );
  NOR U25564 ( .A(n93), .B(n74), .Z(n26196) );
  IV U25565 ( .A(n26196), .Z(n25168) );
  NOR U25566 ( .A(n73), .B(n168), .Z(n25176) );
  IV U25567 ( .A(n25176), .Z(n25171) );
  NOR U25568 ( .A(n25168), .B(n25171), .Z(n25169) );
  IV U25569 ( .A(n25169), .Z(n25170) );
  NOR U25570 ( .A(n94), .B(n25170), .Z(n25179) );
  NOR U25571 ( .A(n25171), .B(n93), .Z(n25172) );
  XOR U25572 ( .A(n94), .B(n25172), .Z(n25173) );
  NOR U25573 ( .A(n74), .B(n25173), .Z(n25174) );
  IV U25574 ( .A(n25174), .Z(n25659) );
  XOR U25575 ( .A(n25176), .B(n25175), .Z(n25658) );
  IV U25576 ( .A(n25658), .Z(n25177) );
  NOR U25577 ( .A(n25659), .B(n25177), .Z(n25178) );
  NOR U25578 ( .A(n25179), .B(n25178), .Z(n25655) );
  XOR U25579 ( .A(n25181), .B(n25180), .Z(n25654) );
  NOR U25580 ( .A(n25655), .B(n25654), .Z(n25182) );
  NOR U25581 ( .A(n25183), .B(n25182), .Z(n25685) );
  XOR U25582 ( .A(n25185), .B(n25184), .Z(n25684) );
  NOR U25583 ( .A(n25685), .B(n25684), .Z(n25186) );
  NOR U25584 ( .A(n25187), .B(n25186), .Z(n25192) );
  NOR U25585 ( .A(n97), .B(n74), .Z(n25191) );
  IV U25586 ( .A(n25191), .Z(n25188) );
  NOR U25587 ( .A(n25192), .B(n25188), .Z(n25195) );
  XOR U25588 ( .A(n25190), .B(n25189), .Z(n25652) );
  IV U25589 ( .A(n25652), .Z(n25193) );
  XOR U25590 ( .A(n25192), .B(n25191), .Z(n25651) );
  NOR U25591 ( .A(n25193), .B(n25651), .Z(n25194) );
  NOR U25592 ( .A(n25195), .B(n25194), .Z(n25647) );
  XOR U25593 ( .A(n25197), .B(n25196), .Z(n25648) );
  NOR U25594 ( .A(n25647), .B(n25648), .Z(n25198) );
  NOR U25595 ( .A(n25199), .B(n25198), .Z(n25643) );
  XOR U25596 ( .A(n25201), .B(n25200), .Z(n25644) );
  NOR U25597 ( .A(n25643), .B(n25644), .Z(n25202) );
  NOR U25598 ( .A(n25203), .B(n25202), .Z(n25639) );
  XOR U25599 ( .A(n25205), .B(n25204), .Z(n25640) );
  NOR U25600 ( .A(n25639), .B(n25640), .Z(n25206) );
  NOR U25601 ( .A(n25207), .B(n25206), .Z(n25635) );
  XOR U25602 ( .A(n25209), .B(n25208), .Z(n25636) );
  NOR U25603 ( .A(n25635), .B(n25636), .Z(n25210) );
  NOR U25604 ( .A(n25211), .B(n25210), .Z(n25631) );
  XOR U25605 ( .A(n25213), .B(n25212), .Z(n25632) );
  NOR U25606 ( .A(n25631), .B(n25632), .Z(n25214) );
  NOR U25607 ( .A(n25215), .B(n25214), .Z(n25627) );
  XOR U25608 ( .A(n25217), .B(n25216), .Z(n25628) );
  NOR U25609 ( .A(n25627), .B(n25628), .Z(n25218) );
  NOR U25610 ( .A(n25219), .B(n25218), .Z(n25623) );
  XOR U25611 ( .A(n25221), .B(n25220), .Z(n25624) );
  NOR U25612 ( .A(n25623), .B(n25624), .Z(n25222) );
  NOR U25613 ( .A(n25223), .B(n25222), .Z(n25620) );
  XOR U25614 ( .A(n25225), .B(n25224), .Z(n25619) );
  NOR U25615 ( .A(n25620), .B(n25619), .Z(n25226) );
  NOR U25616 ( .A(n25227), .B(n25226), .Z(n25726) );
  XOR U25617 ( .A(n25229), .B(n25228), .Z(n25725) );
  NOR U25618 ( .A(n25726), .B(n25725), .Z(n25230) );
  NOR U25619 ( .A(n25231), .B(n25230), .Z(n25236) );
  XOR U25620 ( .A(n25233), .B(n25232), .Z(n25235) );
  IV U25621 ( .A(n25235), .Z(n25234) );
  NOR U25622 ( .A(n25236), .B(n25234), .Z(n25239) );
  XOR U25623 ( .A(n25236), .B(n25235), .Z(n25616) );
  NOR U25624 ( .A(n104), .B(n74), .Z(n25617) );
  IV U25625 ( .A(n25617), .Z(n25237) );
  NOR U25626 ( .A(n25616), .B(n25237), .Z(n25238) );
  NOR U25627 ( .A(n25239), .B(n25238), .Z(n25612) );
  XOR U25628 ( .A(n25241), .B(n25240), .Z(n25613) );
  NOR U25629 ( .A(n25612), .B(n25613), .Z(n25242) );
  NOR U25630 ( .A(n25243), .B(n25242), .Z(n25608) );
  XOR U25631 ( .A(n25245), .B(n25244), .Z(n25609) );
  NOR U25632 ( .A(n25608), .B(n25609), .Z(n25246) );
  NOR U25633 ( .A(n25247), .B(n25246), .Z(n25604) );
  XOR U25634 ( .A(n25249), .B(n25248), .Z(n25605) );
  NOR U25635 ( .A(n25604), .B(n25605), .Z(n25250) );
  NOR U25636 ( .A(n25251), .B(n25250), .Z(n25601) );
  XOR U25637 ( .A(n25253), .B(n25252), .Z(n25600) );
  NOR U25638 ( .A(n25601), .B(n25600), .Z(n25254) );
  NOR U25639 ( .A(n25255), .B(n25254), .Z(n25754) );
  XOR U25640 ( .A(n25257), .B(n25256), .Z(n25753) );
  NOR U25641 ( .A(n25754), .B(n25753), .Z(n25258) );
  NOR U25642 ( .A(n25259), .B(n25258), .Z(n25264) );
  XOR U25643 ( .A(n25261), .B(n25260), .Z(n25263) );
  IV U25644 ( .A(n25263), .Z(n25262) );
  NOR U25645 ( .A(n25264), .B(n25262), .Z(n25267) );
  XOR U25646 ( .A(n25264), .B(n25263), .Z(n25597) );
  NOR U25647 ( .A(n108), .B(n74), .Z(n25598) );
  IV U25648 ( .A(n25598), .Z(n25265) );
  NOR U25649 ( .A(n25597), .B(n25265), .Z(n25266) );
  NOR U25650 ( .A(n25267), .B(n25266), .Z(n25593) );
  XOR U25651 ( .A(n25269), .B(n25268), .Z(n25594) );
  NOR U25652 ( .A(n25593), .B(n25594), .Z(n25270) );
  NOR U25653 ( .A(n25271), .B(n25270), .Z(n25589) );
  XOR U25654 ( .A(n25273), .B(n25272), .Z(n25590) );
  NOR U25655 ( .A(n25589), .B(n25590), .Z(n25274) );
  NOR U25656 ( .A(n25275), .B(n25274), .Z(n25585) );
  XOR U25657 ( .A(n25277), .B(n25276), .Z(n25586) );
  NOR U25658 ( .A(n25585), .B(n25586), .Z(n25278) );
  NOR U25659 ( .A(n25279), .B(n25278), .Z(n25581) );
  XOR U25660 ( .A(n25281), .B(n25280), .Z(n25582) );
  NOR U25661 ( .A(n25581), .B(n25582), .Z(n25282) );
  NOR U25662 ( .A(n25283), .B(n25282), .Z(n25577) );
  XOR U25663 ( .A(n25285), .B(n25284), .Z(n25578) );
  NOR U25664 ( .A(n25577), .B(n25578), .Z(n25286) );
  NOR U25665 ( .A(n25287), .B(n25286), .Z(n25573) );
  XOR U25666 ( .A(n25289), .B(n25288), .Z(n25574) );
  NOR U25667 ( .A(n25573), .B(n25574), .Z(n25290) );
  NOR U25668 ( .A(n25291), .B(n25290), .Z(n25569) );
  XOR U25669 ( .A(n25293), .B(n25292), .Z(n25570) );
  NOR U25670 ( .A(n25569), .B(n25570), .Z(n25294) );
  NOR U25671 ( .A(n25295), .B(n25294), .Z(n25565) );
  XOR U25672 ( .A(n25297), .B(n25296), .Z(n25566) );
  NOR U25673 ( .A(n25565), .B(n25566), .Z(n25298) );
  NOR U25674 ( .A(n25299), .B(n25298), .Z(n25561) );
  XOR U25675 ( .A(n25301), .B(n25300), .Z(n25562) );
  NOR U25676 ( .A(n25561), .B(n25562), .Z(n25302) );
  NOR U25677 ( .A(n25303), .B(n25302), .Z(n25557) );
  XOR U25678 ( .A(n25305), .B(n25304), .Z(n25558) );
  NOR U25679 ( .A(n25557), .B(n25558), .Z(n25306) );
  NOR U25680 ( .A(n25307), .B(n25306), .Z(n25553) );
  XOR U25681 ( .A(n25309), .B(n25308), .Z(n25554) );
  NOR U25682 ( .A(n25553), .B(n25554), .Z(n25310) );
  NOR U25683 ( .A(n25311), .B(n25310), .Z(n25549) );
  XOR U25684 ( .A(n25313), .B(n25312), .Z(n25550) );
  NOR U25685 ( .A(n25549), .B(n25550), .Z(n25314) );
  NOR U25686 ( .A(n25315), .B(n25314), .Z(n25545) );
  XOR U25687 ( .A(n25317), .B(n25316), .Z(n25546) );
  NOR U25688 ( .A(n25545), .B(n25546), .Z(n25318) );
  NOR U25689 ( .A(n25319), .B(n25318), .Z(n25541) );
  XOR U25690 ( .A(n25321), .B(n25320), .Z(n25542) );
  NOR U25691 ( .A(n25541), .B(n25542), .Z(n25322) );
  NOR U25692 ( .A(n25323), .B(n25322), .Z(n25537) );
  XOR U25693 ( .A(n25325), .B(n25324), .Z(n25538) );
  NOR U25694 ( .A(n25537), .B(n25538), .Z(n25326) );
  NOR U25695 ( .A(n25327), .B(n25326), .Z(n25536) );
  XOR U25696 ( .A(n25329), .B(n25328), .Z(n25535) );
  NOR U25697 ( .A(n25536), .B(n25535), .Z(n25330) );
  NOR U25698 ( .A(n25331), .B(n25330), .Z(n25332) );
  IV U25699 ( .A(n25332), .Z(n25533) );
  XOR U25700 ( .A(n25334), .B(n25333), .Z(n25335) );
  IV U25701 ( .A(n25335), .Z(n25532) );
  NOR U25702 ( .A(n25533), .B(n25532), .Z(n25336) );
  NOR U25703 ( .A(n25337), .B(n25336), .Z(n25338) );
  IV U25704 ( .A(n25338), .Z(n25531) );
  XOR U25705 ( .A(n25340), .B(n25339), .Z(n25530) );
  NOR U25706 ( .A(n25531), .B(n25530), .Z(n25341) );
  NOR U25707 ( .A(n25342), .B(n25341), .Z(n25343) );
  IV U25708 ( .A(n25343), .Z(n25527) );
  NOR U25709 ( .A(n25528), .B(n25527), .Z(n25344) );
  NOR U25710 ( .A(n25345), .B(n25344), .Z(n25346) );
  IV U25711 ( .A(n25346), .Z(n25526) );
  XOR U25712 ( .A(n25348), .B(n25347), .Z(n25525) );
  NOR U25713 ( .A(n25526), .B(n25525), .Z(n25349) );
  NOR U25714 ( .A(n25350), .B(n25349), .Z(n25351) );
  IV U25715 ( .A(n25351), .Z(n25523) );
  XOR U25716 ( .A(n25353), .B(n25352), .Z(n25354) );
  IV U25717 ( .A(n25354), .Z(n25522) );
  NOR U25718 ( .A(n25523), .B(n25522), .Z(n25355) );
  NOR U25719 ( .A(n25356), .B(n25355), .Z(n25357) );
  IV U25720 ( .A(n25357), .Z(n25521) );
  XOR U25721 ( .A(n25359), .B(n25358), .Z(n25520) );
  NOR U25722 ( .A(n25521), .B(n25520), .Z(n25360) );
  NOR U25723 ( .A(n25361), .B(n25360), .Z(n25362) );
  IV U25724 ( .A(n25362), .Z(n25518) );
  XOR U25725 ( .A(n25364), .B(n25363), .Z(n25365) );
  IV U25726 ( .A(n25365), .Z(n25517) );
  NOR U25727 ( .A(n25518), .B(n25517), .Z(n25366) );
  NOR U25728 ( .A(n25367), .B(n25366), .Z(n25368) );
  IV U25729 ( .A(n25368), .Z(n25513) );
  XOR U25730 ( .A(n25370), .B(n25369), .Z(n25512) );
  NOR U25731 ( .A(n25513), .B(n25512), .Z(n25371) );
  NOR U25732 ( .A(n25372), .B(n25371), .Z(n25373) );
  IV U25733 ( .A(n25373), .Z(n25510) );
  XOR U25734 ( .A(n25375), .B(n25374), .Z(n25376) );
  IV U25735 ( .A(n25376), .Z(n25509) );
  NOR U25736 ( .A(n25510), .B(n25509), .Z(n25377) );
  NOR U25737 ( .A(n25378), .B(n25377), .Z(n25379) );
  IV U25738 ( .A(n25379), .Z(n25508) );
  XOR U25739 ( .A(n25381), .B(n25380), .Z(n25507) );
  NOR U25740 ( .A(n25508), .B(n25507), .Z(n25382) );
  NOR U25741 ( .A(n25383), .B(n25382), .Z(n25501) );
  XOR U25742 ( .A(n25385), .B(n25384), .Z(n25502) );
  NOR U25743 ( .A(n25501), .B(n25502), .Z(n25386) );
  NOR U25744 ( .A(n25387), .B(n25386), .Z(n25498) );
  XOR U25745 ( .A(n25389), .B(n25388), .Z(n25497) );
  NOR U25746 ( .A(n25498), .B(n25497), .Z(n25390) );
  NOR U25747 ( .A(n25391), .B(n25390), .Z(n25493) );
  XOR U25748 ( .A(n25393), .B(n25392), .Z(n25494) );
  NOR U25749 ( .A(n25493), .B(n25494), .Z(n25394) );
  NOR U25750 ( .A(n25395), .B(n25394), .Z(n25489) );
  XOR U25751 ( .A(n25397), .B(n25396), .Z(n25490) );
  NOR U25752 ( .A(n25489), .B(n25490), .Z(n25398) );
  NOR U25753 ( .A(n25399), .B(n25398), .Z(n25902) );
  XOR U25754 ( .A(n25401), .B(n25400), .Z(n25901) );
  NOR U25755 ( .A(n25902), .B(n25901), .Z(n25402) );
  NOR U25756 ( .A(n25403), .B(n25402), .Z(n25485) );
  XOR U25757 ( .A(n25405), .B(n25404), .Z(n25484) );
  NOR U25758 ( .A(n25485), .B(n25484), .Z(n25406) );
  NOR U25759 ( .A(n25407), .B(n25406), .Z(n25480) );
  NOR U25760 ( .A(n25479), .B(n25482), .Z(n25408) );
  NOR U25761 ( .A(n25480), .B(n25408), .Z(n25409) );
  NOR U25762 ( .A(n25410), .B(n25409), .Z(n25416) );
  XOR U25763 ( .A(n25412), .B(n25411), .Z(n25413) );
  XOR U25764 ( .A(n25414), .B(n25413), .Z(n25415) );
  NOR U25765 ( .A(n25416), .B(n25415), .Z(n25420) );
  XOR U25766 ( .A(n25416), .B(n25415), .Z(n25476) );
  IV U25767 ( .A(n25476), .Z(n25418) );
  NOR U25768 ( .A(n150), .B(n74), .Z(n25417) );
  IV U25769 ( .A(n25417), .Z(n25475) );
  NOR U25770 ( .A(n25418), .B(n25475), .Z(n25419) );
  NOR U25771 ( .A(n25420), .B(n25419), .Z(n25421) );
  IV U25772 ( .A(n25421), .Z(n25474) );
  XOR U25773 ( .A(n25423), .B(n25422), .Z(n25424) );
  IV U25774 ( .A(n25424), .Z(n25473) );
  NOR U25775 ( .A(n25474), .B(n25473), .Z(n25425) );
  NOR U25776 ( .A(n25426), .B(n25425), .Z(n25432) );
  IV U25777 ( .A(n25432), .Z(n25427) );
  NOR U25778 ( .A(n25433), .B(n25427), .Z(n25435) );
  XOR U25779 ( .A(n25429), .B(n25428), .Z(n25430) );
  XOR U25780 ( .A(n25431), .B(n25430), .Z(n25469) );
  XOR U25781 ( .A(n25433), .B(n25432), .Z(n25470) );
  NOR U25782 ( .A(n25469), .B(n25470), .Z(n25434) );
  NOR U25783 ( .A(n25435), .B(n25434), .Z(n25930) );
  XOR U25784 ( .A(n25437), .B(n25436), .Z(n25931) );
  NOR U25785 ( .A(n25930), .B(n25931), .Z(n25438) );
  NOR U25786 ( .A(n25439), .B(n25438), .Z(n25444) );
  XOR U25787 ( .A(n25441), .B(n25440), .Z(n25443) );
  IV U25788 ( .A(n25443), .Z(n25442) );
  NOR U25789 ( .A(n25444), .B(n25442), .Z(n25447) );
  XOR U25790 ( .A(n25444), .B(n25443), .Z(n25938) );
  NOR U25791 ( .A(n158), .B(n74), .Z(n25445) );
  IV U25792 ( .A(n25445), .Z(n25937) );
  NOR U25793 ( .A(n25938), .B(n25937), .Z(n25446) );
  NOR U25794 ( .A(n25447), .B(n25446), .Z(n25451) );
  IV U25795 ( .A(n25451), .Z(n25945) );
  NOR U25796 ( .A(n25450), .B(n25945), .Z(n25454) );
  XOR U25797 ( .A(n25449), .B(n25448), .Z(n25948) );
  IV U25798 ( .A(n25450), .Z(n25946) );
  NOR U25799 ( .A(n25451), .B(n25946), .Z(n25452) );
  NOR U25800 ( .A(n25948), .B(n25452), .Z(n25453) );
  NOR U25801 ( .A(n25454), .B(n25453), .Z(n25458) );
  IV U25802 ( .A(n25458), .Z(n25456) );
  NOR U25803 ( .A(n163), .B(n74), .Z(n25455) );
  IV U25804 ( .A(n25455), .Z(n25457) );
  NOR U25805 ( .A(n25456), .B(n25457), .Z(n25463) );
  XOR U25806 ( .A(n25458), .B(n25457), .Z(n25955) );
  XOR U25807 ( .A(n25460), .B(n25459), .Z(n25461) );
  IV U25808 ( .A(n25461), .Z(n25954) );
  NOR U25809 ( .A(n25955), .B(n25954), .Z(n25462) );
  NOR U25810 ( .A(n25463), .B(n25462), .Z(n25965) );
  XOR U25811 ( .A(n25465), .B(n25464), .Z(n25963) );
  XOR U25812 ( .A(n25965), .B(n25963), .Z(n25968) );
  XOR U25813 ( .A(n25966), .B(n25968), .Z(n25467) );
  NOR U25814 ( .A(n167), .B(n75), .Z(n25468) );
  IV U25815 ( .A(n25468), .Z(n25466) );
  NOR U25816 ( .A(n25467), .B(n25466), .Z(n25962) );
  XOR U25817 ( .A(n25468), .B(n25467), .Z(n26485) );
  NOR U25818 ( .A(n165), .B(n75), .Z(n25957) );
  NOR U25819 ( .A(n161), .B(n75), .Z(n26463) );
  NOR U25820 ( .A(n156), .B(n75), .Z(n25471) );
  XOR U25821 ( .A(n25470), .B(n25469), .Z(n25472) );
  NOR U25822 ( .A(n25471), .B(n25472), .Z(n25927) );
  IV U25823 ( .A(n25471), .Z(n26452) );
  IV U25824 ( .A(n25472), .Z(n26451) );
  NOR U25825 ( .A(n26452), .B(n26451), .Z(n25925) );
  XOR U25826 ( .A(n25474), .B(n25473), .Z(n25920) );
  NOR U25827 ( .A(n153), .B(n75), .Z(n25478) );
  XOR U25828 ( .A(n25476), .B(n25475), .Z(n26442) );
  IV U25829 ( .A(n26442), .Z(n25477) );
  NOR U25830 ( .A(n25478), .B(n25477), .Z(n25917) );
  IV U25831 ( .A(n25478), .Z(n26439) );
  NOR U25832 ( .A(n26439), .B(n26442), .Z(n25915) );
  XOR U25833 ( .A(n25480), .B(n25479), .Z(n25481) );
  XOR U25834 ( .A(n25482), .B(n25481), .Z(n25910) );
  NOR U25835 ( .A(n150), .B(n75), .Z(n25909) );
  IV U25836 ( .A(n25909), .Z(n25483) );
  NOR U25837 ( .A(n25910), .B(n25483), .Z(n25913) );
  NOR U25838 ( .A(n148), .B(n75), .Z(n25487) );
  XOR U25839 ( .A(n25485), .B(n25484), .Z(n25486) );
  NOR U25840 ( .A(n25487), .B(n25486), .Z(n25908) );
  XOR U25841 ( .A(n25487), .B(n25486), .Z(n25488) );
  IV U25842 ( .A(n25488), .Z(n26010) );
  IV U25843 ( .A(n25489), .Z(n25491) );
  XOR U25844 ( .A(n25491), .B(n25490), .Z(n25894) );
  NOR U25845 ( .A(n145), .B(n75), .Z(n25895) );
  IV U25846 ( .A(n25895), .Z(n25492) );
  NOR U25847 ( .A(n25894), .B(n25492), .Z(n25897) );
  IV U25848 ( .A(n25493), .Z(n25495) );
  XOR U25849 ( .A(n25495), .B(n25494), .Z(n25890) );
  NOR U25850 ( .A(n143), .B(n75), .Z(n25891) );
  IV U25851 ( .A(n25891), .Z(n25496) );
  NOR U25852 ( .A(n25890), .B(n25496), .Z(n25893) );
  XOR U25853 ( .A(n25498), .B(n25497), .Z(n25886) );
  IV U25854 ( .A(n25886), .Z(n25500) );
  NOR U25855 ( .A(n141), .B(n75), .Z(n25499) );
  IV U25856 ( .A(n25499), .Z(n25887) );
  NOR U25857 ( .A(n25500), .B(n25887), .Z(n25889) );
  IV U25858 ( .A(n25501), .Z(n25503) );
  XOR U25859 ( .A(n25503), .B(n25502), .Z(n25505) );
  NOR U25860 ( .A(n139), .B(n75), .Z(n25506) );
  IV U25861 ( .A(n25506), .Z(n25504) );
  NOR U25862 ( .A(n25505), .B(n25504), .Z(n25885) );
  XOR U25863 ( .A(n25506), .B(n25505), .Z(n26023) );
  NOR U25864 ( .A(n137), .B(n75), .Z(n25879) );
  XOR U25865 ( .A(n25508), .B(n25507), .Z(n25878) );
  NOR U25866 ( .A(n25879), .B(n25878), .Z(n25882) );
  XOR U25867 ( .A(n25510), .B(n25509), .Z(n25873) );
  NOR U25868 ( .A(n135), .B(n75), .Z(n25872) );
  IV U25869 ( .A(n25872), .Z(n25511) );
  NOR U25870 ( .A(n25873), .B(n25511), .Z(n25876) );
  NOR U25871 ( .A(n133), .B(n75), .Z(n25515) );
  XOR U25872 ( .A(n25513), .B(n25512), .Z(n25514) );
  NOR U25873 ( .A(n25515), .B(n25514), .Z(n25871) );
  XOR U25874 ( .A(n25515), .B(n25514), .Z(n25516) );
  IV U25875 ( .A(n25516), .Z(n26033) );
  XOR U25876 ( .A(n25518), .B(n25517), .Z(n25866) );
  NOR U25877 ( .A(n131), .B(n75), .Z(n25865) );
  IV U25878 ( .A(n25865), .Z(n25519) );
  NOR U25879 ( .A(n25866), .B(n25519), .Z(n25868) );
  NOR U25880 ( .A(n128), .B(n75), .Z(n25860) );
  XOR U25881 ( .A(n25521), .B(n25520), .Z(n25859) );
  NOR U25882 ( .A(n25860), .B(n25859), .Z(n25863) );
  XOR U25883 ( .A(n25523), .B(n25522), .Z(n25854) );
  NOR U25884 ( .A(n126), .B(n75), .Z(n25853) );
  IV U25885 ( .A(n25853), .Z(n25524) );
  NOR U25886 ( .A(n25854), .B(n25524), .Z(n25857) );
  NOR U25887 ( .A(n125), .B(n75), .Z(n25849) );
  XOR U25888 ( .A(n25526), .B(n25525), .Z(n25848) );
  NOR U25889 ( .A(n25849), .B(n25848), .Z(n25852) );
  XOR U25890 ( .A(n25528), .B(n25527), .Z(n25844) );
  NOR U25891 ( .A(n123), .B(n75), .Z(n25843) );
  IV U25892 ( .A(n25843), .Z(n25529) );
  NOR U25893 ( .A(n25844), .B(n25529), .Z(n25846) );
  NOR U25894 ( .A(n120), .B(n75), .Z(n25838) );
  XOR U25895 ( .A(n25531), .B(n25530), .Z(n25837) );
  NOR U25896 ( .A(n25838), .B(n25837), .Z(n25841) );
  XOR U25897 ( .A(n25533), .B(n25532), .Z(n25833) );
  NOR U25898 ( .A(n119), .B(n75), .Z(n25832) );
  IV U25899 ( .A(n25832), .Z(n25534) );
  NOR U25900 ( .A(n25833), .B(n25534), .Z(n25835) );
  NOR U25901 ( .A(n79), .B(n75), .Z(n25827) );
  XOR U25902 ( .A(n25536), .B(n25535), .Z(n25826) );
  NOR U25903 ( .A(n25827), .B(n25826), .Z(n25830) );
  IV U25904 ( .A(n25537), .Z(n25539) );
  XOR U25905 ( .A(n25539), .B(n25538), .Z(n25821) );
  NOR U25906 ( .A(n117), .B(n75), .Z(n25822) );
  IV U25907 ( .A(n25822), .Z(n25540) );
  NOR U25908 ( .A(n25821), .B(n25540), .Z(n25824) );
  IV U25909 ( .A(n25541), .Z(n25543) );
  XOR U25910 ( .A(n25543), .B(n25542), .Z(n25817) );
  NOR U25911 ( .A(n80), .B(n75), .Z(n25818) );
  IV U25912 ( .A(n25818), .Z(n25544) );
  NOR U25913 ( .A(n25817), .B(n25544), .Z(n25820) );
  IV U25914 ( .A(n25545), .Z(n25547) );
  XOR U25915 ( .A(n25547), .B(n25546), .Z(n25813) );
  NOR U25916 ( .A(n116), .B(n75), .Z(n25814) );
  IV U25917 ( .A(n25814), .Z(n25548) );
  NOR U25918 ( .A(n25813), .B(n25548), .Z(n25816) );
  IV U25919 ( .A(n25549), .Z(n25551) );
  XOR U25920 ( .A(n25551), .B(n25550), .Z(n25809) );
  NOR U25921 ( .A(n81), .B(n75), .Z(n25810) );
  IV U25922 ( .A(n25810), .Z(n25552) );
  NOR U25923 ( .A(n25809), .B(n25552), .Z(n25812) );
  IV U25924 ( .A(n25553), .Z(n25555) );
  XOR U25925 ( .A(n25555), .B(n25554), .Z(n25805) );
  NOR U25926 ( .A(n115), .B(n75), .Z(n25806) );
  IV U25927 ( .A(n25806), .Z(n25556) );
  NOR U25928 ( .A(n25805), .B(n25556), .Z(n25808) );
  IV U25929 ( .A(n25557), .Z(n25559) );
  XOR U25930 ( .A(n25559), .B(n25558), .Z(n25801) );
  NOR U25931 ( .A(n82), .B(n75), .Z(n25802) );
  IV U25932 ( .A(n25802), .Z(n25560) );
  NOR U25933 ( .A(n25801), .B(n25560), .Z(n25804) );
  IV U25934 ( .A(n25561), .Z(n25563) );
  XOR U25935 ( .A(n25563), .B(n25562), .Z(n25797) );
  NOR U25936 ( .A(n114), .B(n75), .Z(n25798) );
  IV U25937 ( .A(n25798), .Z(n25564) );
  NOR U25938 ( .A(n25797), .B(n25564), .Z(n25800) );
  IV U25939 ( .A(n25565), .Z(n25567) );
  XOR U25940 ( .A(n25567), .B(n25566), .Z(n25793) );
  NOR U25941 ( .A(n83), .B(n75), .Z(n25794) );
  IV U25942 ( .A(n25794), .Z(n25568) );
  NOR U25943 ( .A(n25793), .B(n25568), .Z(n25796) );
  IV U25944 ( .A(n25569), .Z(n25571) );
  XOR U25945 ( .A(n25571), .B(n25570), .Z(n25789) );
  NOR U25946 ( .A(n113), .B(n75), .Z(n25790) );
  IV U25947 ( .A(n25790), .Z(n25572) );
  NOR U25948 ( .A(n25789), .B(n25572), .Z(n25792) );
  IV U25949 ( .A(n25573), .Z(n25575) );
  XOR U25950 ( .A(n25575), .B(n25574), .Z(n25785) );
  NOR U25951 ( .A(n84), .B(n75), .Z(n25786) );
  IV U25952 ( .A(n25786), .Z(n25576) );
  NOR U25953 ( .A(n25785), .B(n25576), .Z(n25788) );
  IV U25954 ( .A(n25577), .Z(n25579) );
  XOR U25955 ( .A(n25579), .B(n25578), .Z(n25781) );
  NOR U25956 ( .A(n112), .B(n75), .Z(n25782) );
  IV U25957 ( .A(n25782), .Z(n25580) );
  NOR U25958 ( .A(n25781), .B(n25580), .Z(n25784) );
  IV U25959 ( .A(n25581), .Z(n25583) );
  XOR U25960 ( .A(n25583), .B(n25582), .Z(n25777) );
  NOR U25961 ( .A(n85), .B(n75), .Z(n25778) );
  IV U25962 ( .A(n25778), .Z(n25584) );
  NOR U25963 ( .A(n25777), .B(n25584), .Z(n25780) );
  IV U25964 ( .A(n25585), .Z(n25587) );
  XOR U25965 ( .A(n25587), .B(n25586), .Z(n25773) );
  NOR U25966 ( .A(n111), .B(n75), .Z(n25774) );
  IV U25967 ( .A(n25774), .Z(n25588) );
  NOR U25968 ( .A(n25773), .B(n25588), .Z(n25776) );
  IV U25969 ( .A(n25589), .Z(n25591) );
  XOR U25970 ( .A(n25591), .B(n25590), .Z(n25769) );
  NOR U25971 ( .A(n86), .B(n75), .Z(n25770) );
  IV U25972 ( .A(n25770), .Z(n25592) );
  NOR U25973 ( .A(n25769), .B(n25592), .Z(n25772) );
  IV U25974 ( .A(n25593), .Z(n25595) );
  XOR U25975 ( .A(n25595), .B(n25594), .Z(n25765) );
  NOR U25976 ( .A(n110), .B(n75), .Z(n25766) );
  IV U25977 ( .A(n25766), .Z(n25596) );
  NOR U25978 ( .A(n25765), .B(n25596), .Z(n25768) );
  XOR U25979 ( .A(n25598), .B(n25597), .Z(n25761) );
  NOR U25980 ( .A(n109), .B(n75), .Z(n25762) );
  IV U25981 ( .A(n25762), .Z(n25599) );
  NOR U25982 ( .A(n25761), .B(n25599), .Z(n25764) );
  XOR U25983 ( .A(n25601), .B(n25600), .Z(n25749) );
  IV U25984 ( .A(n25749), .Z(n25603) );
  NOR U25985 ( .A(n87), .B(n75), .Z(n25602) );
  IV U25986 ( .A(n25602), .Z(n25750) );
  NOR U25987 ( .A(n25603), .B(n25750), .Z(n25752) );
  IV U25988 ( .A(n25604), .Z(n25606) );
  XOR U25989 ( .A(n25606), .B(n25605), .Z(n25745) );
  NOR U25990 ( .A(n107), .B(n75), .Z(n25746) );
  IV U25991 ( .A(n25746), .Z(n25607) );
  NOR U25992 ( .A(n25745), .B(n25607), .Z(n25748) );
  IV U25993 ( .A(n25608), .Z(n25610) );
  XOR U25994 ( .A(n25610), .B(n25609), .Z(n25741) );
  NOR U25995 ( .A(n88), .B(n75), .Z(n25742) );
  IV U25996 ( .A(n25742), .Z(n25611) );
  NOR U25997 ( .A(n25741), .B(n25611), .Z(n25744) );
  IV U25998 ( .A(n25612), .Z(n25614) );
  XOR U25999 ( .A(n25614), .B(n25613), .Z(n25737) );
  NOR U26000 ( .A(n106), .B(n75), .Z(n25738) );
  IV U26001 ( .A(n25738), .Z(n25615) );
  NOR U26002 ( .A(n25737), .B(n25615), .Z(n25740) );
  XOR U26003 ( .A(n25617), .B(n25616), .Z(n25733) );
  NOR U26004 ( .A(n105), .B(n75), .Z(n25734) );
  IV U26005 ( .A(n25734), .Z(n25618) );
  NOR U26006 ( .A(n25733), .B(n25618), .Z(n25736) );
  XOR U26007 ( .A(n25620), .B(n25619), .Z(n25721) );
  IV U26008 ( .A(n25721), .Z(n25622) );
  NOR U26009 ( .A(n89), .B(n75), .Z(n25621) );
  IV U26010 ( .A(n25621), .Z(n25722) );
  NOR U26011 ( .A(n25622), .B(n25722), .Z(n25724) );
  IV U26012 ( .A(n25623), .Z(n25625) );
  XOR U26013 ( .A(n25625), .B(n25624), .Z(n25717) );
  NOR U26014 ( .A(n103), .B(n75), .Z(n25718) );
  IV U26015 ( .A(n25718), .Z(n25626) );
  NOR U26016 ( .A(n25717), .B(n25626), .Z(n25720) );
  IV U26017 ( .A(n25627), .Z(n25629) );
  XOR U26018 ( .A(n25629), .B(n25628), .Z(n25713) );
  NOR U26019 ( .A(n90), .B(n75), .Z(n25714) );
  IV U26020 ( .A(n25714), .Z(n25630) );
  NOR U26021 ( .A(n25713), .B(n25630), .Z(n25716) );
  IV U26022 ( .A(n25631), .Z(n25633) );
  XOR U26023 ( .A(n25633), .B(n25632), .Z(n25709) );
  NOR U26024 ( .A(n102), .B(n75), .Z(n25710) );
  IV U26025 ( .A(n25710), .Z(n25634) );
  NOR U26026 ( .A(n25709), .B(n25634), .Z(n25712) );
  IV U26027 ( .A(n25635), .Z(n25637) );
  XOR U26028 ( .A(n25637), .B(n25636), .Z(n25705) );
  NOR U26029 ( .A(n101), .B(n75), .Z(n25706) );
  IV U26030 ( .A(n25706), .Z(n25638) );
  NOR U26031 ( .A(n25705), .B(n25638), .Z(n25708) );
  IV U26032 ( .A(n25639), .Z(n25641) );
  XOR U26033 ( .A(n25641), .B(n25640), .Z(n25701) );
  NOR U26034 ( .A(n100), .B(n75), .Z(n25702) );
  IV U26035 ( .A(n25702), .Z(n25642) );
  NOR U26036 ( .A(n25701), .B(n25642), .Z(n25704) );
  IV U26037 ( .A(n25643), .Z(n25645) );
  XOR U26038 ( .A(n25645), .B(n25644), .Z(n25697) );
  NOR U26039 ( .A(n99), .B(n75), .Z(n25698) );
  IV U26040 ( .A(n25698), .Z(n25646) );
  NOR U26041 ( .A(n25697), .B(n25646), .Z(n25700) );
  IV U26042 ( .A(n25647), .Z(n25649) );
  XOR U26043 ( .A(n25649), .B(n25648), .Z(n25693) );
  NOR U26044 ( .A(n98), .B(n75), .Z(n25694) );
  IV U26045 ( .A(n25694), .Z(n25650) );
  NOR U26046 ( .A(n25693), .B(n25650), .Z(n25696) );
  XOR U26047 ( .A(n25652), .B(n25651), .Z(n25689) );
  NOR U26048 ( .A(n91), .B(n75), .Z(n25690) );
  IV U26049 ( .A(n25690), .Z(n25653) );
  NOR U26050 ( .A(n25689), .B(n25653), .Z(n25692) );
  XOR U26051 ( .A(n25655), .B(n25654), .Z(n25677) );
  IV U26052 ( .A(n25677), .Z(n25657) );
  NOR U26053 ( .A(n96), .B(n75), .Z(n25656) );
  IV U26054 ( .A(n25656), .Z(n25678) );
  NOR U26055 ( .A(n25657), .B(n25678), .Z(n25680) );
  NOR U26056 ( .A(n95), .B(n75), .Z(n25674) );
  IV U26057 ( .A(n25674), .Z(n25660) );
  XOR U26058 ( .A(n25659), .B(n25658), .Z(n25673) );
  NOR U26059 ( .A(n25660), .B(n25673), .Z(n25676) );
  NOR U26060 ( .A(n93), .B(n75), .Z(n26707) );
  IV U26061 ( .A(n26707), .Z(n25661) );
  NOR U26062 ( .A(n74), .B(n168), .Z(n25669) );
  IV U26063 ( .A(n25669), .Z(n25664) );
  NOR U26064 ( .A(n25661), .B(n25664), .Z(n25662) );
  IV U26065 ( .A(n25662), .Z(n25663) );
  NOR U26066 ( .A(n94), .B(n25663), .Z(n25672) );
  NOR U26067 ( .A(n25664), .B(n93), .Z(n25665) );
  XOR U26068 ( .A(n94), .B(n25665), .Z(n25666) );
  NOR U26069 ( .A(n75), .B(n25666), .Z(n25667) );
  IV U26070 ( .A(n25667), .Z(n26187) );
  XOR U26071 ( .A(n25669), .B(n25668), .Z(n26186) );
  IV U26072 ( .A(n26186), .Z(n25670) );
  NOR U26073 ( .A(n26187), .B(n25670), .Z(n25671) );
  NOR U26074 ( .A(n25672), .B(n25671), .Z(n26182) );
  XOR U26075 ( .A(n25674), .B(n25673), .Z(n26183) );
  NOR U26076 ( .A(n26182), .B(n26183), .Z(n25675) );
  NOR U26077 ( .A(n25676), .B(n25675), .Z(n26210) );
  XOR U26078 ( .A(n25678), .B(n25677), .Z(n26209) );
  NOR U26079 ( .A(n26210), .B(n26209), .Z(n25679) );
  NOR U26080 ( .A(n25680), .B(n25679), .Z(n25683) );
  NOR U26081 ( .A(n97), .B(n75), .Z(n25682) );
  IV U26082 ( .A(n25682), .Z(n25681) );
  NOR U26083 ( .A(n25683), .B(n25681), .Z(n25688) );
  XOR U26084 ( .A(n25683), .B(n25682), .Z(n26179) );
  XOR U26085 ( .A(n25685), .B(n25684), .Z(n26180) );
  IV U26086 ( .A(n26180), .Z(n25686) );
  NOR U26087 ( .A(n26179), .B(n25686), .Z(n25687) );
  NOR U26088 ( .A(n25688), .B(n25687), .Z(n26175) );
  XOR U26089 ( .A(n25690), .B(n25689), .Z(n26176) );
  NOR U26090 ( .A(n26175), .B(n26176), .Z(n25691) );
  NOR U26091 ( .A(n25692), .B(n25691), .Z(n26171) );
  XOR U26092 ( .A(n25694), .B(n25693), .Z(n26172) );
  NOR U26093 ( .A(n26171), .B(n26172), .Z(n25695) );
  NOR U26094 ( .A(n25696), .B(n25695), .Z(n26167) );
  XOR U26095 ( .A(n25698), .B(n25697), .Z(n26168) );
  NOR U26096 ( .A(n26167), .B(n26168), .Z(n25699) );
  NOR U26097 ( .A(n25700), .B(n25699), .Z(n26163) );
  XOR U26098 ( .A(n25702), .B(n25701), .Z(n26164) );
  NOR U26099 ( .A(n26163), .B(n26164), .Z(n25703) );
  NOR U26100 ( .A(n25704), .B(n25703), .Z(n26159) );
  XOR U26101 ( .A(n25706), .B(n25705), .Z(n26160) );
  NOR U26102 ( .A(n26159), .B(n26160), .Z(n25707) );
  NOR U26103 ( .A(n25708), .B(n25707), .Z(n26155) );
  XOR U26104 ( .A(n25710), .B(n25709), .Z(n26156) );
  NOR U26105 ( .A(n26155), .B(n26156), .Z(n25711) );
  NOR U26106 ( .A(n25712), .B(n25711), .Z(n26151) );
  XOR U26107 ( .A(n25714), .B(n25713), .Z(n26152) );
  NOR U26108 ( .A(n26151), .B(n26152), .Z(n25715) );
  NOR U26109 ( .A(n25716), .B(n25715), .Z(n26148) );
  XOR U26110 ( .A(n25718), .B(n25717), .Z(n26147) );
  NOR U26111 ( .A(n26148), .B(n26147), .Z(n25719) );
  NOR U26112 ( .A(n25720), .B(n25719), .Z(n26254) );
  XOR U26113 ( .A(n25722), .B(n25721), .Z(n26253) );
  NOR U26114 ( .A(n26254), .B(n26253), .Z(n25723) );
  NOR U26115 ( .A(n25724), .B(n25723), .Z(n25729) );
  XOR U26116 ( .A(n25726), .B(n25725), .Z(n25728) );
  IV U26117 ( .A(n25728), .Z(n25727) );
  NOR U26118 ( .A(n25729), .B(n25727), .Z(n25732) );
  XOR U26119 ( .A(n25729), .B(n25728), .Z(n26144) );
  NOR U26120 ( .A(n104), .B(n75), .Z(n26145) );
  IV U26121 ( .A(n26145), .Z(n25730) );
  NOR U26122 ( .A(n26144), .B(n25730), .Z(n25731) );
  NOR U26123 ( .A(n25732), .B(n25731), .Z(n26140) );
  XOR U26124 ( .A(n25734), .B(n25733), .Z(n26141) );
  NOR U26125 ( .A(n26140), .B(n26141), .Z(n25735) );
  NOR U26126 ( .A(n25736), .B(n25735), .Z(n26136) );
  XOR U26127 ( .A(n25738), .B(n25737), .Z(n26137) );
  NOR U26128 ( .A(n26136), .B(n26137), .Z(n25739) );
  NOR U26129 ( .A(n25740), .B(n25739), .Z(n26132) );
  XOR U26130 ( .A(n25742), .B(n25741), .Z(n26133) );
  NOR U26131 ( .A(n26132), .B(n26133), .Z(n25743) );
  NOR U26132 ( .A(n25744), .B(n25743), .Z(n26129) );
  XOR U26133 ( .A(n25746), .B(n25745), .Z(n26128) );
  NOR U26134 ( .A(n26129), .B(n26128), .Z(n25747) );
  NOR U26135 ( .A(n25748), .B(n25747), .Z(n26282) );
  XOR U26136 ( .A(n25750), .B(n25749), .Z(n26281) );
  NOR U26137 ( .A(n26282), .B(n26281), .Z(n25751) );
  NOR U26138 ( .A(n25752), .B(n25751), .Z(n25757) );
  XOR U26139 ( .A(n25754), .B(n25753), .Z(n25756) );
  IV U26140 ( .A(n25756), .Z(n25755) );
  NOR U26141 ( .A(n25757), .B(n25755), .Z(n25760) );
  XOR U26142 ( .A(n25757), .B(n25756), .Z(n26125) );
  NOR U26143 ( .A(n108), .B(n75), .Z(n26126) );
  IV U26144 ( .A(n26126), .Z(n25758) );
  NOR U26145 ( .A(n26125), .B(n25758), .Z(n25759) );
  NOR U26146 ( .A(n25760), .B(n25759), .Z(n26121) );
  XOR U26147 ( .A(n25762), .B(n25761), .Z(n26122) );
  NOR U26148 ( .A(n26121), .B(n26122), .Z(n25763) );
  NOR U26149 ( .A(n25764), .B(n25763), .Z(n26117) );
  XOR U26150 ( .A(n25766), .B(n25765), .Z(n26118) );
  NOR U26151 ( .A(n26117), .B(n26118), .Z(n25767) );
  NOR U26152 ( .A(n25768), .B(n25767), .Z(n26113) );
  XOR U26153 ( .A(n25770), .B(n25769), .Z(n26114) );
  NOR U26154 ( .A(n26113), .B(n26114), .Z(n25771) );
  NOR U26155 ( .A(n25772), .B(n25771), .Z(n26109) );
  XOR U26156 ( .A(n25774), .B(n25773), .Z(n26110) );
  NOR U26157 ( .A(n26109), .B(n26110), .Z(n25775) );
  NOR U26158 ( .A(n25776), .B(n25775), .Z(n26105) );
  XOR U26159 ( .A(n25778), .B(n25777), .Z(n26106) );
  NOR U26160 ( .A(n26105), .B(n26106), .Z(n25779) );
  NOR U26161 ( .A(n25780), .B(n25779), .Z(n26101) );
  XOR U26162 ( .A(n25782), .B(n25781), .Z(n26102) );
  NOR U26163 ( .A(n26101), .B(n26102), .Z(n25783) );
  NOR U26164 ( .A(n25784), .B(n25783), .Z(n26097) );
  XOR U26165 ( .A(n25786), .B(n25785), .Z(n26098) );
  NOR U26166 ( .A(n26097), .B(n26098), .Z(n25787) );
  NOR U26167 ( .A(n25788), .B(n25787), .Z(n26093) );
  XOR U26168 ( .A(n25790), .B(n25789), .Z(n26094) );
  NOR U26169 ( .A(n26093), .B(n26094), .Z(n25791) );
  NOR U26170 ( .A(n25792), .B(n25791), .Z(n26089) );
  XOR U26171 ( .A(n25794), .B(n25793), .Z(n26090) );
  NOR U26172 ( .A(n26089), .B(n26090), .Z(n25795) );
  NOR U26173 ( .A(n25796), .B(n25795), .Z(n26085) );
  XOR U26174 ( .A(n25798), .B(n25797), .Z(n26086) );
  NOR U26175 ( .A(n26085), .B(n26086), .Z(n25799) );
  NOR U26176 ( .A(n25800), .B(n25799), .Z(n26081) );
  XOR U26177 ( .A(n25802), .B(n25801), .Z(n26082) );
  NOR U26178 ( .A(n26081), .B(n26082), .Z(n25803) );
  NOR U26179 ( .A(n25804), .B(n25803), .Z(n26077) );
  XOR U26180 ( .A(n25806), .B(n25805), .Z(n26078) );
  NOR U26181 ( .A(n26077), .B(n26078), .Z(n25807) );
  NOR U26182 ( .A(n25808), .B(n25807), .Z(n26073) );
  XOR U26183 ( .A(n25810), .B(n25809), .Z(n26074) );
  NOR U26184 ( .A(n26073), .B(n26074), .Z(n25811) );
  NOR U26185 ( .A(n25812), .B(n25811), .Z(n26069) );
  XOR U26186 ( .A(n25814), .B(n25813), .Z(n26070) );
  NOR U26187 ( .A(n26069), .B(n26070), .Z(n25815) );
  NOR U26188 ( .A(n25816), .B(n25815), .Z(n26065) );
  XOR U26189 ( .A(n25818), .B(n25817), .Z(n26066) );
  NOR U26190 ( .A(n26065), .B(n26066), .Z(n25819) );
  NOR U26191 ( .A(n25820), .B(n25819), .Z(n26061) );
  XOR U26192 ( .A(n25822), .B(n25821), .Z(n26062) );
  NOR U26193 ( .A(n26061), .B(n26062), .Z(n25823) );
  NOR U26194 ( .A(n25824), .B(n25823), .Z(n25825) );
  IV U26195 ( .A(n25825), .Z(n26059) );
  XOR U26196 ( .A(n25827), .B(n25826), .Z(n25828) );
  IV U26197 ( .A(n25828), .Z(n26058) );
  NOR U26198 ( .A(n26059), .B(n26058), .Z(n25829) );
  NOR U26199 ( .A(n25830), .B(n25829), .Z(n25831) );
  IV U26200 ( .A(n25831), .Z(n26057) );
  XOR U26201 ( .A(n25833), .B(n25832), .Z(n26056) );
  NOR U26202 ( .A(n26057), .B(n26056), .Z(n25834) );
  NOR U26203 ( .A(n25835), .B(n25834), .Z(n25836) );
  IV U26204 ( .A(n25836), .Z(n26054) );
  XOR U26205 ( .A(n25838), .B(n25837), .Z(n25839) );
  IV U26206 ( .A(n25839), .Z(n26053) );
  NOR U26207 ( .A(n26054), .B(n26053), .Z(n25840) );
  NOR U26208 ( .A(n25841), .B(n25840), .Z(n25842) );
  IV U26209 ( .A(n25842), .Z(n26049) );
  XOR U26210 ( .A(n25844), .B(n25843), .Z(n26048) );
  NOR U26211 ( .A(n26049), .B(n26048), .Z(n25845) );
  NOR U26212 ( .A(n25846), .B(n25845), .Z(n25847) );
  IV U26213 ( .A(n25847), .Z(n26046) );
  XOR U26214 ( .A(n25849), .B(n25848), .Z(n25850) );
  IV U26215 ( .A(n25850), .Z(n26045) );
  NOR U26216 ( .A(n26046), .B(n26045), .Z(n25851) );
  NOR U26217 ( .A(n25852), .B(n25851), .Z(n26043) );
  IV U26218 ( .A(n26043), .Z(n25855) );
  XOR U26219 ( .A(n25854), .B(n25853), .Z(n26042) );
  NOR U26220 ( .A(n25855), .B(n26042), .Z(n25856) );
  NOR U26221 ( .A(n25857), .B(n25856), .Z(n25858) );
  IV U26222 ( .A(n25858), .Z(n26040) );
  XOR U26223 ( .A(n25860), .B(n25859), .Z(n25861) );
  IV U26224 ( .A(n25861), .Z(n26039) );
  NOR U26225 ( .A(n26040), .B(n26039), .Z(n25862) );
  NOR U26226 ( .A(n25863), .B(n25862), .Z(n25864) );
  IV U26227 ( .A(n25864), .Z(n26038) );
  XOR U26228 ( .A(n25866), .B(n25865), .Z(n26037) );
  NOR U26229 ( .A(n26038), .B(n26037), .Z(n25867) );
  NOR U26230 ( .A(n25868), .B(n25867), .Z(n25869) );
  IV U26231 ( .A(n25869), .Z(n26032) );
  NOR U26232 ( .A(n26033), .B(n26032), .Z(n25870) );
  NOR U26233 ( .A(n25871), .B(n25870), .Z(n26030) );
  IV U26234 ( .A(n26030), .Z(n25874) );
  XOR U26235 ( .A(n25873), .B(n25872), .Z(n26029) );
  NOR U26236 ( .A(n25874), .B(n26029), .Z(n25875) );
  NOR U26237 ( .A(n25876), .B(n25875), .Z(n25877) );
  IV U26238 ( .A(n25877), .Z(n26027) );
  XOR U26239 ( .A(n25879), .B(n25878), .Z(n25880) );
  IV U26240 ( .A(n25880), .Z(n26026) );
  NOR U26241 ( .A(n26027), .B(n26026), .Z(n25881) );
  NOR U26242 ( .A(n25882), .B(n25881), .Z(n26024) );
  IV U26243 ( .A(n26024), .Z(n25883) );
  NOR U26244 ( .A(n26023), .B(n25883), .Z(n25884) );
  NOR U26245 ( .A(n25885), .B(n25884), .Z(n26410) );
  XOR U26246 ( .A(n25887), .B(n25886), .Z(n26409) );
  NOR U26247 ( .A(n26410), .B(n26409), .Z(n25888) );
  NOR U26248 ( .A(n25889), .B(n25888), .Z(n26019) );
  XOR U26249 ( .A(n25891), .B(n25890), .Z(n26020) );
  NOR U26250 ( .A(n26019), .B(n26020), .Z(n25892) );
  NOR U26251 ( .A(n25893), .B(n25892), .Z(n26015) );
  XOR U26252 ( .A(n25895), .B(n25894), .Z(n26016) );
  NOR U26253 ( .A(n26015), .B(n26016), .Z(n25896) );
  NOR U26254 ( .A(n25897), .B(n25896), .Z(n25900) );
  NOR U26255 ( .A(n147), .B(n75), .Z(n25899) );
  IV U26256 ( .A(n25899), .Z(n25898) );
  NOR U26257 ( .A(n25900), .B(n25898), .Z(n25905) );
  XOR U26258 ( .A(n25900), .B(n25899), .Z(n26012) );
  XOR U26259 ( .A(n25902), .B(n25901), .Z(n26013) );
  IV U26260 ( .A(n26013), .Z(n25903) );
  NOR U26261 ( .A(n26012), .B(n25903), .Z(n25904) );
  NOR U26262 ( .A(n25905), .B(n25904), .Z(n25906) );
  IV U26263 ( .A(n25906), .Z(n26009) );
  NOR U26264 ( .A(n26010), .B(n26009), .Z(n25907) );
  NOR U26265 ( .A(n25908), .B(n25907), .Z(n26007) );
  IV U26266 ( .A(n26007), .Z(n25911) );
  XOR U26267 ( .A(n25910), .B(n25909), .Z(n26006) );
  NOR U26268 ( .A(n25911), .B(n26006), .Z(n25912) );
  NOR U26269 ( .A(n25913), .B(n25912), .Z(n25914) );
  IV U26270 ( .A(n25914), .Z(n26440) );
  NOR U26271 ( .A(n25915), .B(n26440), .Z(n25916) );
  NOR U26272 ( .A(n25917), .B(n25916), .Z(n25921) );
  IV U26273 ( .A(n25921), .Z(n25918) );
  NOR U26274 ( .A(n25920), .B(n25918), .Z(n25923) );
  NOR U26275 ( .A(n155), .B(n75), .Z(n25919) );
  IV U26276 ( .A(n25919), .Z(n26003) );
  XOR U26277 ( .A(n25921), .B(n25920), .Z(n26002) );
  NOR U26278 ( .A(n26003), .B(n26002), .Z(n25922) );
  NOR U26279 ( .A(n25923), .B(n25922), .Z(n26454) );
  IV U26280 ( .A(n26454), .Z(n25924) );
  NOR U26281 ( .A(n25925), .B(n25924), .Z(n25926) );
  NOR U26282 ( .A(n25927), .B(n25926), .Z(n25929) );
  IV U26283 ( .A(n25929), .Z(n25998) );
  NOR U26284 ( .A(n158), .B(n75), .Z(n25928) );
  IV U26285 ( .A(n25928), .Z(n25997) );
  NOR U26286 ( .A(n25998), .B(n25997), .Z(n25935) );
  NOR U26287 ( .A(n25929), .B(n25928), .Z(n25933) );
  IV U26288 ( .A(n25930), .Z(n25932) );
  XOR U26289 ( .A(n25932), .B(n25931), .Z(n26000) );
  NOR U26290 ( .A(n25933), .B(n26000), .Z(n25934) );
  NOR U26291 ( .A(n25935), .B(n25934), .Z(n26466) );
  IV U26292 ( .A(n26466), .Z(n25936) );
  NOR U26293 ( .A(n26463), .B(n25936), .Z(n25942) );
  XOR U26294 ( .A(n25938), .B(n25937), .Z(n26464) );
  IV U26295 ( .A(n26463), .Z(n25939) );
  NOR U26296 ( .A(n26466), .B(n25939), .Z(n25940) );
  NOR U26297 ( .A(n26464), .B(n25940), .Z(n25941) );
  NOR U26298 ( .A(n25942), .B(n25941), .Z(n25950) );
  IV U26299 ( .A(n25950), .Z(n25944) );
  NOR U26300 ( .A(n163), .B(n75), .Z(n25943) );
  IV U26301 ( .A(n25943), .Z(n25949) );
  NOR U26302 ( .A(n25944), .B(n25949), .Z(n25952) );
  XOR U26303 ( .A(n25946), .B(n25945), .Z(n25947) );
  XOR U26304 ( .A(n25948), .B(n25947), .Z(n25994) );
  XOR U26305 ( .A(n25950), .B(n25949), .Z(n25993) );
  NOR U26306 ( .A(n25994), .B(n25993), .Z(n25951) );
  NOR U26307 ( .A(n25952), .B(n25951), .Z(n25956) );
  IV U26308 ( .A(n25956), .Z(n25953) );
  NOR U26309 ( .A(n25957), .B(n25953), .Z(n25959) );
  XOR U26310 ( .A(n25955), .B(n25954), .Z(n26480) );
  XOR U26311 ( .A(n25957), .B(n25956), .Z(n26479) );
  NOR U26312 ( .A(n26480), .B(n26479), .Z(n25958) );
  NOR U26313 ( .A(n25959), .B(n25958), .Z(n26486) );
  IV U26314 ( .A(n26486), .Z(n25960) );
  NOR U26315 ( .A(n26485), .B(n25960), .Z(n25961) );
  NOR U26316 ( .A(n25962), .B(n25961), .Z(n26488) );
  IV U26317 ( .A(n25963), .Z(n25964) );
  NOR U26318 ( .A(n25965), .B(n25964), .Z(n25970) );
  IV U26319 ( .A(n25966), .Z(n25967) );
  NOR U26320 ( .A(n25968), .B(n25967), .Z(n25969) );
  NOR U26321 ( .A(n25970), .B(n25969), .Z(n25976) );
  NOR U26322 ( .A(n167), .B(n74), .Z(n25974) );
  XOR U26323 ( .A(n25976), .B(n25974), .Z(n25978) );
  XOR U26324 ( .A(n25972), .B(n25971), .Z(n25977) );
  XOR U26325 ( .A(n25978), .B(n25977), .Z(n26487) );
  IV U26326 ( .A(n26487), .Z(n25973) );
  NOR U26327 ( .A(n26488), .B(n25973), .Z(n28505) );
  IV U26328 ( .A(n28505), .Z(n31484) );
  IV U26329 ( .A(n25974), .Z(n25975) );
  NOR U26330 ( .A(n25976), .B(n25975), .Z(n25980) );
  NOR U26331 ( .A(n25978), .B(n25977), .Z(n25979) );
  NOR U26332 ( .A(n25980), .B(n25979), .Z(n25986) );
  XOR U26333 ( .A(n25982), .B(n25981), .Z(n25984) );
  XOR U26334 ( .A(n25986), .B(n25984), .Z(n28504) );
  NOR U26335 ( .A(n31484), .B(n28504), .Z(n31487) );
  IV U26336 ( .A(n31487), .Z(n25983) );
  NOR U26337 ( .A(n25987), .B(n25983), .Z(n25988) );
  IV U26338 ( .A(n25984), .Z(n25985) );
  NOR U26339 ( .A(n25986), .B(n25985), .Z(n28503) );
  IV U26340 ( .A(n28503), .Z(n31494) );
  NOR U26341 ( .A(n31494), .B(n25987), .Z(n31498) );
  NOR U26342 ( .A(n25988), .B(n31498), .Z(n25989) );
  IV U26343 ( .A(n25989), .Z(n25990) );
  NOR U26344 ( .A(n25991), .B(n25990), .Z(n25992) );
  IV U26345 ( .A(n25992), .Z(n28511) );
  NOR U26346 ( .A(n165), .B(n76), .Z(n25995) );
  XOR U26347 ( .A(n25994), .B(n25993), .Z(n27478) );
  NOR U26348 ( .A(n25995), .B(n27478), .Z(n26476) );
  IV U26349 ( .A(n25995), .Z(n27475) );
  IV U26350 ( .A(n27478), .Z(n25996) );
  NOR U26351 ( .A(n27475), .B(n25996), .Z(n26474) );
  XOR U26352 ( .A(n25998), .B(n25997), .Z(n25999) );
  XOR U26353 ( .A(n26000), .B(n25999), .Z(n26459) );
  NOR U26354 ( .A(n161), .B(n76), .Z(n26489) );
  IV U26355 ( .A(n26489), .Z(n26001) );
  NOR U26356 ( .A(n26459), .B(n26001), .Z(n26462) );
  XOR U26357 ( .A(n26003), .B(n26002), .Z(n26005) );
  IV U26358 ( .A(n26005), .Z(n26498) );
  NOR U26359 ( .A(n156), .B(n76), .Z(n26004) );
  IV U26360 ( .A(n26004), .Z(n26497) );
  NOR U26361 ( .A(n26498), .B(n26497), .Z(n26449) );
  NOR U26362 ( .A(n26005), .B(n26004), .Z(n26447) );
  NOR U26363 ( .A(n155), .B(n76), .Z(n26437) );
  XOR U26364 ( .A(n26007), .B(n26006), .Z(n26433) );
  NOR U26365 ( .A(n153), .B(n76), .Z(n26434) );
  IV U26366 ( .A(n26434), .Z(n26008) );
  NOR U26367 ( .A(n26433), .B(n26008), .Z(n26436) );
  XOR U26368 ( .A(n26010), .B(n26009), .Z(n26430) );
  NOR U26369 ( .A(n150), .B(n76), .Z(n26429) );
  IV U26370 ( .A(n26429), .Z(n26011) );
  NOR U26371 ( .A(n26430), .B(n26011), .Z(n26432) );
  XOR U26372 ( .A(n26013), .B(n26012), .Z(n26425) );
  NOR U26373 ( .A(n148), .B(n76), .Z(n26426) );
  IV U26374 ( .A(n26426), .Z(n26014) );
  NOR U26375 ( .A(n26425), .B(n26014), .Z(n26428) );
  IV U26376 ( .A(n26015), .Z(n26017) );
  XOR U26377 ( .A(n26017), .B(n26016), .Z(n26421) );
  NOR U26378 ( .A(n147), .B(n76), .Z(n26422) );
  IV U26379 ( .A(n26422), .Z(n26018) );
  NOR U26380 ( .A(n26421), .B(n26018), .Z(n26424) );
  IV U26381 ( .A(n26019), .Z(n26021) );
  XOR U26382 ( .A(n26021), .B(n26020), .Z(n26417) );
  NOR U26383 ( .A(n145), .B(n76), .Z(n26418) );
  IV U26384 ( .A(n26418), .Z(n26022) );
  NOR U26385 ( .A(n26417), .B(n26022), .Z(n26420) );
  XOR U26386 ( .A(n26024), .B(n26023), .Z(n26405) );
  NOR U26387 ( .A(n141), .B(n76), .Z(n26406) );
  IV U26388 ( .A(n26406), .Z(n26025) );
  NOR U26389 ( .A(n26405), .B(n26025), .Z(n26408) );
  XOR U26390 ( .A(n26027), .B(n26026), .Z(n26402) );
  NOR U26391 ( .A(n139), .B(n76), .Z(n26401) );
  IV U26392 ( .A(n26401), .Z(n26028) );
  NOR U26393 ( .A(n26402), .B(n26028), .Z(n26404) );
  XOR U26394 ( .A(n26030), .B(n26029), .Z(n26397) );
  NOR U26395 ( .A(n137), .B(n76), .Z(n26398) );
  IV U26396 ( .A(n26398), .Z(n26031) );
  NOR U26397 ( .A(n26397), .B(n26031), .Z(n26400) );
  XOR U26398 ( .A(n26033), .B(n26032), .Z(n26036) );
  NOR U26399 ( .A(n135), .B(n76), .Z(n26035) );
  IV U26400 ( .A(n26035), .Z(n26034) );
  NOR U26401 ( .A(n26036), .B(n26034), .Z(n26396) );
  XOR U26402 ( .A(n26036), .B(n26035), .Z(n26541) );
  NOR U26403 ( .A(n133), .B(n76), .Z(n26390) );
  XOR U26404 ( .A(n26038), .B(n26037), .Z(n26389) );
  NOR U26405 ( .A(n26390), .B(n26389), .Z(n26393) );
  XOR U26406 ( .A(n26040), .B(n26039), .Z(n26385) );
  NOR U26407 ( .A(n131), .B(n76), .Z(n26384) );
  IV U26408 ( .A(n26384), .Z(n26041) );
  NOR U26409 ( .A(n26385), .B(n26041), .Z(n26387) );
  XOR U26410 ( .A(n26043), .B(n26042), .Z(n26380) );
  NOR U26411 ( .A(n128), .B(n76), .Z(n26381) );
  IV U26412 ( .A(n26381), .Z(n26044) );
  NOR U26413 ( .A(n26380), .B(n26044), .Z(n26383) );
  XOR U26414 ( .A(n26046), .B(n26045), .Z(n26376) );
  NOR U26415 ( .A(n126), .B(n76), .Z(n26375) );
  IV U26416 ( .A(n26375), .Z(n26047) );
  NOR U26417 ( .A(n26376), .B(n26047), .Z(n26379) );
  NOR U26418 ( .A(n125), .B(n76), .Z(n26051) );
  XOR U26419 ( .A(n26049), .B(n26048), .Z(n26050) );
  NOR U26420 ( .A(n26051), .B(n26050), .Z(n26374) );
  XOR U26421 ( .A(n26051), .B(n26050), .Z(n26052) );
  IV U26422 ( .A(n26052), .Z(n26555) );
  XOR U26423 ( .A(n26054), .B(n26053), .Z(n26369) );
  NOR U26424 ( .A(n123), .B(n76), .Z(n26368) );
  IV U26425 ( .A(n26368), .Z(n26055) );
  NOR U26426 ( .A(n26369), .B(n26055), .Z(n26371) );
  NOR U26427 ( .A(n120), .B(n76), .Z(n26363) );
  XOR U26428 ( .A(n26057), .B(n26056), .Z(n26362) );
  NOR U26429 ( .A(n26363), .B(n26362), .Z(n26366) );
  XOR U26430 ( .A(n26059), .B(n26058), .Z(n26358) );
  NOR U26431 ( .A(n119), .B(n76), .Z(n26357) );
  IV U26432 ( .A(n26357), .Z(n26060) );
  NOR U26433 ( .A(n26358), .B(n26060), .Z(n26360) );
  IV U26434 ( .A(n26061), .Z(n26063) );
  XOR U26435 ( .A(n26063), .B(n26062), .Z(n26353) );
  NOR U26436 ( .A(n79), .B(n76), .Z(n26354) );
  IV U26437 ( .A(n26354), .Z(n26064) );
  NOR U26438 ( .A(n26353), .B(n26064), .Z(n26356) );
  IV U26439 ( .A(n26065), .Z(n26067) );
  XOR U26440 ( .A(n26067), .B(n26066), .Z(n26349) );
  NOR U26441 ( .A(n117), .B(n76), .Z(n26350) );
  IV U26442 ( .A(n26350), .Z(n26068) );
  NOR U26443 ( .A(n26349), .B(n26068), .Z(n26352) );
  IV U26444 ( .A(n26069), .Z(n26071) );
  XOR U26445 ( .A(n26071), .B(n26070), .Z(n26345) );
  NOR U26446 ( .A(n80), .B(n76), .Z(n26346) );
  IV U26447 ( .A(n26346), .Z(n26072) );
  NOR U26448 ( .A(n26345), .B(n26072), .Z(n26348) );
  IV U26449 ( .A(n26073), .Z(n26075) );
  XOR U26450 ( .A(n26075), .B(n26074), .Z(n26341) );
  NOR U26451 ( .A(n116), .B(n76), .Z(n26342) );
  IV U26452 ( .A(n26342), .Z(n26076) );
  NOR U26453 ( .A(n26341), .B(n26076), .Z(n26344) );
  IV U26454 ( .A(n26077), .Z(n26079) );
  XOR U26455 ( .A(n26079), .B(n26078), .Z(n26337) );
  NOR U26456 ( .A(n81), .B(n76), .Z(n26338) );
  IV U26457 ( .A(n26338), .Z(n26080) );
  NOR U26458 ( .A(n26337), .B(n26080), .Z(n26340) );
  IV U26459 ( .A(n26081), .Z(n26083) );
  XOR U26460 ( .A(n26083), .B(n26082), .Z(n26333) );
  NOR U26461 ( .A(n115), .B(n76), .Z(n26334) );
  IV U26462 ( .A(n26334), .Z(n26084) );
  NOR U26463 ( .A(n26333), .B(n26084), .Z(n26336) );
  IV U26464 ( .A(n26085), .Z(n26087) );
  XOR U26465 ( .A(n26087), .B(n26086), .Z(n26329) );
  NOR U26466 ( .A(n82), .B(n76), .Z(n26330) );
  IV U26467 ( .A(n26330), .Z(n26088) );
  NOR U26468 ( .A(n26329), .B(n26088), .Z(n26332) );
  IV U26469 ( .A(n26089), .Z(n26091) );
  XOR U26470 ( .A(n26091), .B(n26090), .Z(n26325) );
  NOR U26471 ( .A(n114), .B(n76), .Z(n26326) );
  IV U26472 ( .A(n26326), .Z(n26092) );
  NOR U26473 ( .A(n26325), .B(n26092), .Z(n26328) );
  IV U26474 ( .A(n26093), .Z(n26095) );
  XOR U26475 ( .A(n26095), .B(n26094), .Z(n26321) );
  NOR U26476 ( .A(n83), .B(n76), .Z(n26322) );
  IV U26477 ( .A(n26322), .Z(n26096) );
  NOR U26478 ( .A(n26321), .B(n26096), .Z(n26324) );
  IV U26479 ( .A(n26097), .Z(n26099) );
  XOR U26480 ( .A(n26099), .B(n26098), .Z(n26317) );
  NOR U26481 ( .A(n113), .B(n76), .Z(n26318) );
  IV U26482 ( .A(n26318), .Z(n26100) );
  NOR U26483 ( .A(n26317), .B(n26100), .Z(n26320) );
  IV U26484 ( .A(n26101), .Z(n26103) );
  XOR U26485 ( .A(n26103), .B(n26102), .Z(n26313) );
  NOR U26486 ( .A(n84), .B(n76), .Z(n26314) );
  IV U26487 ( .A(n26314), .Z(n26104) );
  NOR U26488 ( .A(n26313), .B(n26104), .Z(n26316) );
  IV U26489 ( .A(n26105), .Z(n26107) );
  XOR U26490 ( .A(n26107), .B(n26106), .Z(n26309) );
  NOR U26491 ( .A(n112), .B(n76), .Z(n26310) );
  IV U26492 ( .A(n26310), .Z(n26108) );
  NOR U26493 ( .A(n26309), .B(n26108), .Z(n26312) );
  IV U26494 ( .A(n26109), .Z(n26111) );
  XOR U26495 ( .A(n26111), .B(n26110), .Z(n26305) );
  NOR U26496 ( .A(n85), .B(n76), .Z(n26306) );
  IV U26497 ( .A(n26306), .Z(n26112) );
  NOR U26498 ( .A(n26305), .B(n26112), .Z(n26308) );
  IV U26499 ( .A(n26113), .Z(n26115) );
  XOR U26500 ( .A(n26115), .B(n26114), .Z(n26301) );
  NOR U26501 ( .A(n111), .B(n76), .Z(n26302) );
  IV U26502 ( .A(n26302), .Z(n26116) );
  NOR U26503 ( .A(n26301), .B(n26116), .Z(n26304) );
  IV U26504 ( .A(n26117), .Z(n26119) );
  XOR U26505 ( .A(n26119), .B(n26118), .Z(n26297) );
  NOR U26506 ( .A(n86), .B(n76), .Z(n26298) );
  IV U26507 ( .A(n26298), .Z(n26120) );
  NOR U26508 ( .A(n26297), .B(n26120), .Z(n26300) );
  IV U26509 ( .A(n26121), .Z(n26123) );
  XOR U26510 ( .A(n26123), .B(n26122), .Z(n26293) );
  NOR U26511 ( .A(n110), .B(n76), .Z(n26294) );
  IV U26512 ( .A(n26294), .Z(n26124) );
  NOR U26513 ( .A(n26293), .B(n26124), .Z(n26296) );
  XOR U26514 ( .A(n26126), .B(n26125), .Z(n26289) );
  NOR U26515 ( .A(n109), .B(n76), .Z(n26290) );
  IV U26516 ( .A(n26290), .Z(n26127) );
  NOR U26517 ( .A(n26289), .B(n26127), .Z(n26292) );
  XOR U26518 ( .A(n26129), .B(n26128), .Z(n26277) );
  IV U26519 ( .A(n26277), .Z(n26131) );
  NOR U26520 ( .A(n87), .B(n76), .Z(n26130) );
  IV U26521 ( .A(n26130), .Z(n26278) );
  NOR U26522 ( .A(n26131), .B(n26278), .Z(n26280) );
  IV U26523 ( .A(n26132), .Z(n26134) );
  XOR U26524 ( .A(n26134), .B(n26133), .Z(n26273) );
  NOR U26525 ( .A(n107), .B(n76), .Z(n26274) );
  IV U26526 ( .A(n26274), .Z(n26135) );
  NOR U26527 ( .A(n26273), .B(n26135), .Z(n26276) );
  IV U26528 ( .A(n26136), .Z(n26138) );
  XOR U26529 ( .A(n26138), .B(n26137), .Z(n26269) );
  NOR U26530 ( .A(n88), .B(n76), .Z(n26270) );
  IV U26531 ( .A(n26270), .Z(n26139) );
  NOR U26532 ( .A(n26269), .B(n26139), .Z(n26272) );
  IV U26533 ( .A(n26140), .Z(n26142) );
  XOR U26534 ( .A(n26142), .B(n26141), .Z(n26265) );
  NOR U26535 ( .A(n106), .B(n76), .Z(n26266) );
  IV U26536 ( .A(n26266), .Z(n26143) );
  NOR U26537 ( .A(n26265), .B(n26143), .Z(n26268) );
  XOR U26538 ( .A(n26145), .B(n26144), .Z(n26261) );
  NOR U26539 ( .A(n105), .B(n76), .Z(n26262) );
  IV U26540 ( .A(n26262), .Z(n26146) );
  NOR U26541 ( .A(n26261), .B(n26146), .Z(n26264) );
  XOR U26542 ( .A(n26148), .B(n26147), .Z(n26249) );
  IV U26543 ( .A(n26249), .Z(n26150) );
  NOR U26544 ( .A(n89), .B(n76), .Z(n26149) );
  IV U26545 ( .A(n26149), .Z(n26250) );
  NOR U26546 ( .A(n26150), .B(n26250), .Z(n26252) );
  IV U26547 ( .A(n26151), .Z(n26153) );
  XOR U26548 ( .A(n26153), .B(n26152), .Z(n26245) );
  NOR U26549 ( .A(n103), .B(n76), .Z(n26246) );
  IV U26550 ( .A(n26246), .Z(n26154) );
  NOR U26551 ( .A(n26245), .B(n26154), .Z(n26248) );
  IV U26552 ( .A(n26155), .Z(n26157) );
  XOR U26553 ( .A(n26157), .B(n26156), .Z(n26241) );
  NOR U26554 ( .A(n90), .B(n76), .Z(n26242) );
  IV U26555 ( .A(n26242), .Z(n26158) );
  NOR U26556 ( .A(n26241), .B(n26158), .Z(n26244) );
  IV U26557 ( .A(n26159), .Z(n26161) );
  XOR U26558 ( .A(n26161), .B(n26160), .Z(n26237) );
  NOR U26559 ( .A(n102), .B(n76), .Z(n26238) );
  IV U26560 ( .A(n26238), .Z(n26162) );
  NOR U26561 ( .A(n26237), .B(n26162), .Z(n26240) );
  IV U26562 ( .A(n26163), .Z(n26165) );
  XOR U26563 ( .A(n26165), .B(n26164), .Z(n26233) );
  NOR U26564 ( .A(n101), .B(n76), .Z(n26234) );
  IV U26565 ( .A(n26234), .Z(n26166) );
  NOR U26566 ( .A(n26233), .B(n26166), .Z(n26236) );
  IV U26567 ( .A(n26167), .Z(n26169) );
  XOR U26568 ( .A(n26169), .B(n26168), .Z(n26229) );
  NOR U26569 ( .A(n100), .B(n76), .Z(n26230) );
  IV U26570 ( .A(n26230), .Z(n26170) );
  NOR U26571 ( .A(n26229), .B(n26170), .Z(n26232) );
  IV U26572 ( .A(n26171), .Z(n26173) );
  XOR U26573 ( .A(n26173), .B(n26172), .Z(n26225) );
  NOR U26574 ( .A(n99), .B(n76), .Z(n26226) );
  IV U26575 ( .A(n26226), .Z(n26174) );
  NOR U26576 ( .A(n26225), .B(n26174), .Z(n26228) );
  XOR U26577 ( .A(n26176), .B(n26175), .Z(n26177) );
  IV U26578 ( .A(n26177), .Z(n26221) );
  NOR U26579 ( .A(n98), .B(n76), .Z(n26222) );
  IV U26580 ( .A(n26222), .Z(n26178) );
  NOR U26581 ( .A(n26221), .B(n26178), .Z(n26224) );
  XOR U26582 ( .A(n26180), .B(n26179), .Z(n26217) );
  NOR U26583 ( .A(n91), .B(n76), .Z(n26218) );
  IV U26584 ( .A(n26218), .Z(n26181) );
  NOR U26585 ( .A(n26217), .B(n26181), .Z(n26220) );
  IV U26586 ( .A(n26182), .Z(n26184) );
  XOR U26587 ( .A(n26184), .B(n26183), .Z(n26205) );
  NOR U26588 ( .A(n96), .B(n76), .Z(n26206) );
  IV U26589 ( .A(n26206), .Z(n26185) );
  NOR U26590 ( .A(n26205), .B(n26185), .Z(n26208) );
  NOR U26591 ( .A(n95), .B(n76), .Z(n26202) );
  IV U26592 ( .A(n26202), .Z(n26188) );
  XOR U26593 ( .A(n26187), .B(n26186), .Z(n26201) );
  NOR U26594 ( .A(n26188), .B(n26201), .Z(n26204) );
  NOR U26595 ( .A(n93), .B(n76), .Z(n27189) );
  IV U26596 ( .A(n27189), .Z(n26189) );
  NOR U26597 ( .A(n75), .B(n168), .Z(n26197) );
  IV U26598 ( .A(n26197), .Z(n26192) );
  NOR U26599 ( .A(n26189), .B(n26192), .Z(n26190) );
  IV U26600 ( .A(n26190), .Z(n26191) );
  NOR U26601 ( .A(n94), .B(n26191), .Z(n26200) );
  NOR U26602 ( .A(n26192), .B(n93), .Z(n26193) );
  XOR U26603 ( .A(n94), .B(n26193), .Z(n26194) );
  NOR U26604 ( .A(n76), .B(n26194), .Z(n26195) );
  IV U26605 ( .A(n26195), .Z(n26698) );
  XOR U26606 ( .A(n26197), .B(n26196), .Z(n26697) );
  IV U26607 ( .A(n26697), .Z(n26198) );
  NOR U26608 ( .A(n26698), .B(n26198), .Z(n26199) );
  NOR U26609 ( .A(n26200), .B(n26199), .Z(n26693) );
  XOR U26610 ( .A(n26202), .B(n26201), .Z(n26694) );
  NOR U26611 ( .A(n26693), .B(n26694), .Z(n26203) );
  NOR U26612 ( .A(n26204), .B(n26203), .Z(n26689) );
  XOR U26613 ( .A(n26206), .B(n26205), .Z(n26690) );
  NOR U26614 ( .A(n26689), .B(n26690), .Z(n26207) );
  NOR U26615 ( .A(n26208), .B(n26207), .Z(n26213) );
  XOR U26616 ( .A(n26210), .B(n26209), .Z(n26212) );
  IV U26617 ( .A(n26212), .Z(n26211) );
  NOR U26618 ( .A(n26213), .B(n26211), .Z(n26216) );
  XOR U26619 ( .A(n26213), .B(n26212), .Z(n26686) );
  NOR U26620 ( .A(n97), .B(n76), .Z(n26687) );
  IV U26621 ( .A(n26687), .Z(n26214) );
  NOR U26622 ( .A(n26686), .B(n26214), .Z(n26215) );
  NOR U26623 ( .A(n26216), .B(n26215), .Z(n26682) );
  XOR U26624 ( .A(n26218), .B(n26217), .Z(n26683) );
  NOR U26625 ( .A(n26682), .B(n26683), .Z(n26219) );
  NOR U26626 ( .A(n26220), .B(n26219), .Z(n26678) );
  XOR U26627 ( .A(n26222), .B(n26221), .Z(n26679) );
  NOR U26628 ( .A(n26678), .B(n26679), .Z(n26223) );
  NOR U26629 ( .A(n26224), .B(n26223), .Z(n26674) );
  XOR U26630 ( .A(n26226), .B(n26225), .Z(n26675) );
  NOR U26631 ( .A(n26674), .B(n26675), .Z(n26227) );
  NOR U26632 ( .A(n26228), .B(n26227), .Z(n26670) );
  XOR U26633 ( .A(n26230), .B(n26229), .Z(n26671) );
  NOR U26634 ( .A(n26670), .B(n26671), .Z(n26231) );
  NOR U26635 ( .A(n26232), .B(n26231), .Z(n26666) );
  XOR U26636 ( .A(n26234), .B(n26233), .Z(n26667) );
  NOR U26637 ( .A(n26666), .B(n26667), .Z(n26235) );
  NOR U26638 ( .A(n26236), .B(n26235), .Z(n26662) );
  XOR U26639 ( .A(n26238), .B(n26237), .Z(n26663) );
  NOR U26640 ( .A(n26662), .B(n26663), .Z(n26239) );
  NOR U26641 ( .A(n26240), .B(n26239), .Z(n26658) );
  XOR U26642 ( .A(n26242), .B(n26241), .Z(n26659) );
  NOR U26643 ( .A(n26658), .B(n26659), .Z(n26243) );
  NOR U26644 ( .A(n26244), .B(n26243), .Z(n26655) );
  XOR U26645 ( .A(n26246), .B(n26245), .Z(n26654) );
  NOR U26646 ( .A(n26655), .B(n26654), .Z(n26247) );
  NOR U26647 ( .A(n26248), .B(n26247), .Z(n26761) );
  XOR U26648 ( .A(n26250), .B(n26249), .Z(n26760) );
  NOR U26649 ( .A(n26761), .B(n26760), .Z(n26251) );
  NOR U26650 ( .A(n26252), .B(n26251), .Z(n26257) );
  XOR U26651 ( .A(n26254), .B(n26253), .Z(n26256) );
  IV U26652 ( .A(n26256), .Z(n26255) );
  NOR U26653 ( .A(n26257), .B(n26255), .Z(n26260) );
  XOR U26654 ( .A(n26257), .B(n26256), .Z(n26651) );
  NOR U26655 ( .A(n104), .B(n76), .Z(n26652) );
  IV U26656 ( .A(n26652), .Z(n26258) );
  NOR U26657 ( .A(n26651), .B(n26258), .Z(n26259) );
  NOR U26658 ( .A(n26260), .B(n26259), .Z(n26647) );
  XOR U26659 ( .A(n26262), .B(n26261), .Z(n26648) );
  NOR U26660 ( .A(n26647), .B(n26648), .Z(n26263) );
  NOR U26661 ( .A(n26264), .B(n26263), .Z(n26643) );
  XOR U26662 ( .A(n26266), .B(n26265), .Z(n26644) );
  NOR U26663 ( .A(n26643), .B(n26644), .Z(n26267) );
  NOR U26664 ( .A(n26268), .B(n26267), .Z(n26639) );
  XOR U26665 ( .A(n26270), .B(n26269), .Z(n26640) );
  NOR U26666 ( .A(n26639), .B(n26640), .Z(n26271) );
  NOR U26667 ( .A(n26272), .B(n26271), .Z(n26636) );
  XOR U26668 ( .A(n26274), .B(n26273), .Z(n26635) );
  NOR U26669 ( .A(n26636), .B(n26635), .Z(n26275) );
  NOR U26670 ( .A(n26276), .B(n26275), .Z(n26792) );
  XOR U26671 ( .A(n26278), .B(n26277), .Z(n26791) );
  NOR U26672 ( .A(n26792), .B(n26791), .Z(n26279) );
  NOR U26673 ( .A(n26280), .B(n26279), .Z(n26285) );
  XOR U26674 ( .A(n26282), .B(n26281), .Z(n26284) );
  IV U26675 ( .A(n26284), .Z(n26283) );
  NOR U26676 ( .A(n26285), .B(n26283), .Z(n26288) );
  XOR U26677 ( .A(n26285), .B(n26284), .Z(n26632) );
  NOR U26678 ( .A(n108), .B(n76), .Z(n26633) );
  IV U26679 ( .A(n26633), .Z(n26286) );
  NOR U26680 ( .A(n26632), .B(n26286), .Z(n26287) );
  NOR U26681 ( .A(n26288), .B(n26287), .Z(n26628) );
  XOR U26682 ( .A(n26290), .B(n26289), .Z(n26629) );
  NOR U26683 ( .A(n26628), .B(n26629), .Z(n26291) );
  NOR U26684 ( .A(n26292), .B(n26291), .Z(n26624) );
  XOR U26685 ( .A(n26294), .B(n26293), .Z(n26625) );
  NOR U26686 ( .A(n26624), .B(n26625), .Z(n26295) );
  NOR U26687 ( .A(n26296), .B(n26295), .Z(n26620) );
  XOR U26688 ( .A(n26298), .B(n26297), .Z(n26621) );
  NOR U26689 ( .A(n26620), .B(n26621), .Z(n26299) );
  NOR U26690 ( .A(n26300), .B(n26299), .Z(n26616) );
  XOR U26691 ( .A(n26302), .B(n26301), .Z(n26617) );
  NOR U26692 ( .A(n26616), .B(n26617), .Z(n26303) );
  NOR U26693 ( .A(n26304), .B(n26303), .Z(n26612) );
  XOR U26694 ( .A(n26306), .B(n26305), .Z(n26613) );
  NOR U26695 ( .A(n26612), .B(n26613), .Z(n26307) );
  NOR U26696 ( .A(n26308), .B(n26307), .Z(n26608) );
  XOR U26697 ( .A(n26310), .B(n26309), .Z(n26609) );
  NOR U26698 ( .A(n26608), .B(n26609), .Z(n26311) );
  NOR U26699 ( .A(n26312), .B(n26311), .Z(n26604) );
  XOR U26700 ( .A(n26314), .B(n26313), .Z(n26605) );
  NOR U26701 ( .A(n26604), .B(n26605), .Z(n26315) );
  NOR U26702 ( .A(n26316), .B(n26315), .Z(n26600) );
  XOR U26703 ( .A(n26318), .B(n26317), .Z(n26601) );
  NOR U26704 ( .A(n26600), .B(n26601), .Z(n26319) );
  NOR U26705 ( .A(n26320), .B(n26319), .Z(n26596) );
  XOR U26706 ( .A(n26322), .B(n26321), .Z(n26597) );
  NOR U26707 ( .A(n26596), .B(n26597), .Z(n26323) );
  NOR U26708 ( .A(n26324), .B(n26323), .Z(n26592) );
  XOR U26709 ( .A(n26326), .B(n26325), .Z(n26593) );
  NOR U26710 ( .A(n26592), .B(n26593), .Z(n26327) );
  NOR U26711 ( .A(n26328), .B(n26327), .Z(n26588) );
  XOR U26712 ( .A(n26330), .B(n26329), .Z(n26589) );
  NOR U26713 ( .A(n26588), .B(n26589), .Z(n26331) );
  NOR U26714 ( .A(n26332), .B(n26331), .Z(n26584) );
  XOR U26715 ( .A(n26334), .B(n26333), .Z(n26585) );
  NOR U26716 ( .A(n26584), .B(n26585), .Z(n26335) );
  NOR U26717 ( .A(n26336), .B(n26335), .Z(n26580) );
  XOR U26718 ( .A(n26338), .B(n26337), .Z(n26581) );
  NOR U26719 ( .A(n26580), .B(n26581), .Z(n26339) );
  NOR U26720 ( .A(n26340), .B(n26339), .Z(n26576) );
  XOR U26721 ( .A(n26342), .B(n26341), .Z(n26577) );
  NOR U26722 ( .A(n26576), .B(n26577), .Z(n26343) );
  NOR U26723 ( .A(n26344), .B(n26343), .Z(n26572) );
  XOR U26724 ( .A(n26346), .B(n26345), .Z(n26573) );
  NOR U26725 ( .A(n26572), .B(n26573), .Z(n26347) );
  NOR U26726 ( .A(n26348), .B(n26347), .Z(n26568) );
  XOR U26727 ( .A(n26350), .B(n26349), .Z(n26569) );
  NOR U26728 ( .A(n26568), .B(n26569), .Z(n26351) );
  NOR U26729 ( .A(n26352), .B(n26351), .Z(n26564) );
  XOR U26730 ( .A(n26354), .B(n26353), .Z(n26565) );
  NOR U26731 ( .A(n26564), .B(n26565), .Z(n26355) );
  NOR U26732 ( .A(n26356), .B(n26355), .Z(n26563) );
  XOR U26733 ( .A(n26358), .B(n26357), .Z(n26562) );
  NOR U26734 ( .A(n26563), .B(n26562), .Z(n26359) );
  NOR U26735 ( .A(n26360), .B(n26359), .Z(n26361) );
  IV U26736 ( .A(n26361), .Z(n26560) );
  XOR U26737 ( .A(n26363), .B(n26362), .Z(n26364) );
  IV U26738 ( .A(n26364), .Z(n26559) );
  NOR U26739 ( .A(n26560), .B(n26559), .Z(n26365) );
  NOR U26740 ( .A(n26366), .B(n26365), .Z(n26367) );
  IV U26741 ( .A(n26367), .Z(n26558) );
  XOR U26742 ( .A(n26369), .B(n26368), .Z(n26557) );
  NOR U26743 ( .A(n26558), .B(n26557), .Z(n26370) );
  NOR U26744 ( .A(n26371), .B(n26370), .Z(n26372) );
  IV U26745 ( .A(n26372), .Z(n26554) );
  NOR U26746 ( .A(n26555), .B(n26554), .Z(n26373) );
  NOR U26747 ( .A(n26374), .B(n26373), .Z(n26552) );
  IV U26748 ( .A(n26552), .Z(n26377) );
  XOR U26749 ( .A(n26376), .B(n26375), .Z(n26551) );
  NOR U26750 ( .A(n26377), .B(n26551), .Z(n26378) );
  NOR U26751 ( .A(n26379), .B(n26378), .Z(n26895) );
  XOR U26752 ( .A(n26381), .B(n26380), .Z(n26894) );
  NOR U26753 ( .A(n26895), .B(n26894), .Z(n26382) );
  NOR U26754 ( .A(n26383), .B(n26382), .Z(n26547) );
  XOR U26755 ( .A(n26385), .B(n26384), .Z(n26548) );
  NOR U26756 ( .A(n26547), .B(n26548), .Z(n26386) );
  NOR U26757 ( .A(n26387), .B(n26386), .Z(n26388) );
  IV U26758 ( .A(n26388), .Z(n26545) );
  XOR U26759 ( .A(n26390), .B(n26389), .Z(n26391) );
  IV U26760 ( .A(n26391), .Z(n26544) );
  NOR U26761 ( .A(n26545), .B(n26544), .Z(n26392) );
  NOR U26762 ( .A(n26393), .B(n26392), .Z(n26542) );
  IV U26763 ( .A(n26542), .Z(n26394) );
  NOR U26764 ( .A(n26541), .B(n26394), .Z(n26395) );
  NOR U26765 ( .A(n26396), .B(n26395), .Z(n26537) );
  XOR U26766 ( .A(n26398), .B(n26397), .Z(n26538) );
  NOR U26767 ( .A(n26537), .B(n26538), .Z(n26399) );
  NOR U26768 ( .A(n26400), .B(n26399), .Z(n26533) );
  XOR U26769 ( .A(n26402), .B(n26401), .Z(n26534) );
  NOR U26770 ( .A(n26533), .B(n26534), .Z(n26403) );
  NOR U26771 ( .A(n26404), .B(n26403), .Z(n26529) );
  XOR U26772 ( .A(n26406), .B(n26405), .Z(n26530) );
  NOR U26773 ( .A(n26529), .B(n26530), .Z(n26407) );
  NOR U26774 ( .A(n26408), .B(n26407), .Z(n26413) );
  XOR U26775 ( .A(n26410), .B(n26409), .Z(n26412) );
  IV U26776 ( .A(n26412), .Z(n26411) );
  NOR U26777 ( .A(n26413), .B(n26411), .Z(n26416) );
  XOR U26778 ( .A(n26413), .B(n26412), .Z(n26526) );
  NOR U26779 ( .A(n143), .B(n76), .Z(n26527) );
  IV U26780 ( .A(n26527), .Z(n26414) );
  NOR U26781 ( .A(n26526), .B(n26414), .Z(n26415) );
  NOR U26782 ( .A(n26416), .B(n26415), .Z(n26522) );
  XOR U26783 ( .A(n26418), .B(n26417), .Z(n26523) );
  NOR U26784 ( .A(n26522), .B(n26523), .Z(n26419) );
  NOR U26785 ( .A(n26420), .B(n26419), .Z(n26518) );
  XOR U26786 ( .A(n26422), .B(n26421), .Z(n26519) );
  NOR U26787 ( .A(n26518), .B(n26519), .Z(n26423) );
  NOR U26788 ( .A(n26424), .B(n26423), .Z(n26514) );
  XOR U26789 ( .A(n26426), .B(n26425), .Z(n26515) );
  NOR U26790 ( .A(n26514), .B(n26515), .Z(n26427) );
  NOR U26791 ( .A(n26428), .B(n26427), .Z(n26510) );
  XOR U26792 ( .A(n26430), .B(n26429), .Z(n26511) );
  NOR U26793 ( .A(n26510), .B(n26511), .Z(n26431) );
  NOR U26794 ( .A(n26432), .B(n26431), .Z(n26506) );
  XOR U26795 ( .A(n26434), .B(n26433), .Z(n26507) );
  NOR U26796 ( .A(n26506), .B(n26507), .Z(n26435) );
  NOR U26797 ( .A(n26436), .B(n26435), .Z(n26438) );
  IV U26798 ( .A(n26438), .Z(n26502) );
  NOR U26799 ( .A(n26437), .B(n26502), .Z(n26445) );
  IV U26800 ( .A(n26437), .Z(n26501) );
  NOR U26801 ( .A(n26438), .B(n26501), .Z(n26443) );
  XOR U26802 ( .A(n26440), .B(n26439), .Z(n26441) );
  XOR U26803 ( .A(n26442), .B(n26441), .Z(n26504) );
  NOR U26804 ( .A(n26443), .B(n26504), .Z(n26444) );
  NOR U26805 ( .A(n26445), .B(n26444), .Z(n26446) );
  IV U26806 ( .A(n26446), .Z(n26500) );
  NOR U26807 ( .A(n26447), .B(n26500), .Z(n26448) );
  NOR U26808 ( .A(n26449), .B(n26448), .Z(n26456) );
  NOR U26809 ( .A(n158), .B(n76), .Z(n26455) );
  IV U26810 ( .A(n26455), .Z(n26450) );
  NOR U26811 ( .A(n26456), .B(n26450), .Z(n26458) );
  XOR U26812 ( .A(n26452), .B(n26451), .Z(n26453) );
  XOR U26813 ( .A(n26454), .B(n26453), .Z(n26494) );
  XOR U26814 ( .A(n26456), .B(n26455), .Z(n26493) );
  NOR U26815 ( .A(n26494), .B(n26493), .Z(n26457) );
  NOR U26816 ( .A(n26458), .B(n26457), .Z(n26490) );
  IV U26817 ( .A(n26459), .Z(n26492) );
  NOR U26818 ( .A(n26492), .B(n26489), .Z(n26460) );
  NOR U26819 ( .A(n26490), .B(n26460), .Z(n26461) );
  NOR U26820 ( .A(n26462), .B(n26461), .Z(n26467) );
  XOR U26821 ( .A(n26464), .B(n26463), .Z(n26465) );
  XOR U26822 ( .A(n26466), .B(n26465), .Z(n26468) );
  NOR U26823 ( .A(n26467), .B(n26468), .Z(n26472) );
  XOR U26824 ( .A(n26468), .B(n26467), .Z(n26469) );
  IV U26825 ( .A(n26469), .Z(n27454) );
  NOR U26826 ( .A(n163), .B(n76), .Z(n26470) );
  IV U26827 ( .A(n26470), .Z(n27455) );
  NOR U26828 ( .A(n27454), .B(n27455), .Z(n26471) );
  NOR U26829 ( .A(n26472), .B(n26471), .Z(n26473) );
  IV U26830 ( .A(n26473), .Z(n27476) );
  NOR U26831 ( .A(n26474), .B(n27476), .Z(n26475) );
  NOR U26832 ( .A(n26476), .B(n26475), .Z(n26477) );
  IV U26833 ( .A(n26477), .Z(n26482) );
  NOR U26834 ( .A(n167), .B(n76), .Z(n26481) );
  IV U26835 ( .A(n26481), .Z(n26478) );
  NOR U26836 ( .A(n26482), .B(n26478), .Z(n26484) );
  XOR U26837 ( .A(n26480), .B(n26479), .Z(n27486) );
  XOR U26838 ( .A(n26482), .B(n26481), .Z(n27487) );
  NOR U26839 ( .A(n27486), .B(n27487), .Z(n26483) );
  NOR U26840 ( .A(n26484), .B(n26483), .Z(n28001) );
  XOR U26841 ( .A(n26486), .B(n26485), .Z(n28000) );
  NOR U26842 ( .A(n28001), .B(n28000), .Z(n31476) );
  XOR U26843 ( .A(n26488), .B(n26487), .Z(n31481) );
  XOR U26844 ( .A(n26490), .B(n26489), .Z(n26491) );
  XOR U26845 ( .A(n26492), .B(n26491), .Z(n27460) );
  NOR U26846 ( .A(n163), .B(n77), .Z(n27459) );
  IV U26847 ( .A(n27459), .Z(n27456) );
  XOR U26848 ( .A(n26494), .B(n26493), .Z(n26496) );
  IV U26849 ( .A(n26496), .Z(n26965) );
  NOR U26850 ( .A(n161), .B(n77), .Z(n26495) );
  IV U26851 ( .A(n26495), .Z(n26964) );
  NOR U26852 ( .A(n26965), .B(n26964), .Z(n26962) );
  NOR U26853 ( .A(n26496), .B(n26495), .Z(n26960) );
  XOR U26854 ( .A(n26498), .B(n26497), .Z(n26499) );
  XOR U26855 ( .A(n26500), .B(n26499), .Z(n26954) );
  IV U26856 ( .A(n26954), .Z(n26970) );
  XOR U26857 ( .A(n26502), .B(n26501), .Z(n26503) );
  XOR U26858 ( .A(n26504), .B(n26503), .Z(n26950) );
  NOR U26859 ( .A(n156), .B(n77), .Z(n26976) );
  IV U26860 ( .A(n26976), .Z(n26505) );
  NOR U26861 ( .A(n26950), .B(n26505), .Z(n26953) );
  IV U26862 ( .A(n26506), .Z(n26508) );
  XOR U26863 ( .A(n26508), .B(n26507), .Z(n26946) );
  NOR U26864 ( .A(n155), .B(n77), .Z(n26947) );
  IV U26865 ( .A(n26947), .Z(n26509) );
  NOR U26866 ( .A(n26946), .B(n26509), .Z(n26949) );
  IV U26867 ( .A(n26510), .Z(n26512) );
  XOR U26868 ( .A(n26512), .B(n26511), .Z(n26942) );
  NOR U26869 ( .A(n153), .B(n77), .Z(n26943) );
  IV U26870 ( .A(n26943), .Z(n26513) );
  NOR U26871 ( .A(n26942), .B(n26513), .Z(n26945) );
  IV U26872 ( .A(n26514), .Z(n26516) );
  XOR U26873 ( .A(n26516), .B(n26515), .Z(n26938) );
  NOR U26874 ( .A(n150), .B(n77), .Z(n26939) );
  IV U26875 ( .A(n26939), .Z(n26517) );
  NOR U26876 ( .A(n26938), .B(n26517), .Z(n26941) );
  IV U26877 ( .A(n26518), .Z(n26520) );
  XOR U26878 ( .A(n26520), .B(n26519), .Z(n26934) );
  NOR U26879 ( .A(n148), .B(n77), .Z(n26935) );
  IV U26880 ( .A(n26935), .Z(n26521) );
  NOR U26881 ( .A(n26934), .B(n26521), .Z(n26937) );
  IV U26882 ( .A(n26522), .Z(n26524) );
  XOR U26883 ( .A(n26524), .B(n26523), .Z(n26930) );
  NOR U26884 ( .A(n147), .B(n77), .Z(n26931) );
  IV U26885 ( .A(n26931), .Z(n26525) );
  NOR U26886 ( .A(n26930), .B(n26525), .Z(n26933) );
  XOR U26887 ( .A(n26527), .B(n26526), .Z(n26926) );
  NOR U26888 ( .A(n145), .B(n77), .Z(n26927) );
  IV U26889 ( .A(n26927), .Z(n26528) );
  NOR U26890 ( .A(n26926), .B(n26528), .Z(n26929) );
  IV U26891 ( .A(n26529), .Z(n26531) );
  XOR U26892 ( .A(n26531), .B(n26530), .Z(n26922) );
  NOR U26893 ( .A(n143), .B(n77), .Z(n26923) );
  IV U26894 ( .A(n26923), .Z(n26532) );
  NOR U26895 ( .A(n26922), .B(n26532), .Z(n26925) );
  IV U26896 ( .A(n26533), .Z(n26535) );
  XOR U26897 ( .A(n26535), .B(n26534), .Z(n26918) );
  NOR U26898 ( .A(n141), .B(n77), .Z(n26919) );
  IV U26899 ( .A(n26919), .Z(n26536) );
  NOR U26900 ( .A(n26918), .B(n26536), .Z(n26921) );
  IV U26901 ( .A(n26537), .Z(n26539) );
  XOR U26902 ( .A(n26539), .B(n26538), .Z(n26914) );
  NOR U26903 ( .A(n139), .B(n77), .Z(n26915) );
  IV U26904 ( .A(n26915), .Z(n26540) );
  NOR U26905 ( .A(n26914), .B(n26540), .Z(n26917) );
  XOR U26906 ( .A(n26542), .B(n26541), .Z(n26910) );
  NOR U26907 ( .A(n137), .B(n77), .Z(n26911) );
  IV U26908 ( .A(n26911), .Z(n26543) );
  NOR U26909 ( .A(n26910), .B(n26543), .Z(n26913) );
  XOR U26910 ( .A(n26545), .B(n26544), .Z(n26907) );
  NOR U26911 ( .A(n135), .B(n77), .Z(n26906) );
  IV U26912 ( .A(n26906), .Z(n26546) );
  NOR U26913 ( .A(n26907), .B(n26546), .Z(n26909) );
  IV U26914 ( .A(n26547), .Z(n26549) );
  XOR U26915 ( .A(n26549), .B(n26548), .Z(n26902) );
  NOR U26916 ( .A(n133), .B(n77), .Z(n26903) );
  IV U26917 ( .A(n26903), .Z(n26550) );
  NOR U26918 ( .A(n26902), .B(n26550), .Z(n26905) );
  XOR U26919 ( .A(n26552), .B(n26551), .Z(n26890) );
  NOR U26920 ( .A(n128), .B(n77), .Z(n26891) );
  IV U26921 ( .A(n26891), .Z(n26553) );
  NOR U26922 ( .A(n26890), .B(n26553), .Z(n26893) );
  XOR U26923 ( .A(n26555), .B(n26554), .Z(n26886) );
  NOR U26924 ( .A(n126), .B(n77), .Z(n26885) );
  IV U26925 ( .A(n26885), .Z(n26556) );
  NOR U26926 ( .A(n26886), .B(n26556), .Z(n26889) );
  NOR U26927 ( .A(n125), .B(n77), .Z(n26881) );
  XOR U26928 ( .A(n26558), .B(n26557), .Z(n26880) );
  NOR U26929 ( .A(n26881), .B(n26880), .Z(n26884) );
  XOR U26930 ( .A(n26560), .B(n26559), .Z(n26876) );
  NOR U26931 ( .A(n123), .B(n77), .Z(n26875) );
  IV U26932 ( .A(n26875), .Z(n26561) );
  NOR U26933 ( .A(n26876), .B(n26561), .Z(n26878) );
  NOR U26934 ( .A(n120), .B(n77), .Z(n26870) );
  XOR U26935 ( .A(n26563), .B(n26562), .Z(n26869) );
  NOR U26936 ( .A(n26870), .B(n26869), .Z(n26873) );
  IV U26937 ( .A(n26564), .Z(n26566) );
  XOR U26938 ( .A(n26566), .B(n26565), .Z(n26864) );
  NOR U26939 ( .A(n119), .B(n77), .Z(n26865) );
  IV U26940 ( .A(n26865), .Z(n26567) );
  NOR U26941 ( .A(n26864), .B(n26567), .Z(n26867) );
  IV U26942 ( .A(n26568), .Z(n26570) );
  XOR U26943 ( .A(n26570), .B(n26569), .Z(n26860) );
  NOR U26944 ( .A(n79), .B(n77), .Z(n26861) );
  IV U26945 ( .A(n26861), .Z(n26571) );
  NOR U26946 ( .A(n26860), .B(n26571), .Z(n26863) );
  IV U26947 ( .A(n26572), .Z(n26574) );
  XOR U26948 ( .A(n26574), .B(n26573), .Z(n26856) );
  NOR U26949 ( .A(n117), .B(n77), .Z(n26857) );
  IV U26950 ( .A(n26857), .Z(n26575) );
  NOR U26951 ( .A(n26856), .B(n26575), .Z(n26859) );
  IV U26952 ( .A(n26576), .Z(n26578) );
  XOR U26953 ( .A(n26578), .B(n26577), .Z(n26852) );
  NOR U26954 ( .A(n80), .B(n77), .Z(n26853) );
  IV U26955 ( .A(n26853), .Z(n26579) );
  NOR U26956 ( .A(n26852), .B(n26579), .Z(n26855) );
  IV U26957 ( .A(n26580), .Z(n26582) );
  XOR U26958 ( .A(n26582), .B(n26581), .Z(n26848) );
  NOR U26959 ( .A(n116), .B(n77), .Z(n26849) );
  IV U26960 ( .A(n26849), .Z(n26583) );
  NOR U26961 ( .A(n26848), .B(n26583), .Z(n26851) );
  IV U26962 ( .A(n26584), .Z(n26586) );
  XOR U26963 ( .A(n26586), .B(n26585), .Z(n26844) );
  NOR U26964 ( .A(n81), .B(n77), .Z(n26845) );
  IV U26965 ( .A(n26845), .Z(n26587) );
  NOR U26966 ( .A(n26844), .B(n26587), .Z(n26847) );
  IV U26967 ( .A(n26588), .Z(n26590) );
  XOR U26968 ( .A(n26590), .B(n26589), .Z(n26840) );
  NOR U26969 ( .A(n115), .B(n77), .Z(n26841) );
  IV U26970 ( .A(n26841), .Z(n26591) );
  NOR U26971 ( .A(n26840), .B(n26591), .Z(n26843) );
  IV U26972 ( .A(n26592), .Z(n26594) );
  XOR U26973 ( .A(n26594), .B(n26593), .Z(n26836) );
  NOR U26974 ( .A(n82), .B(n77), .Z(n26837) );
  IV U26975 ( .A(n26837), .Z(n26595) );
  NOR U26976 ( .A(n26836), .B(n26595), .Z(n26839) );
  IV U26977 ( .A(n26596), .Z(n26598) );
  XOR U26978 ( .A(n26598), .B(n26597), .Z(n26832) );
  NOR U26979 ( .A(n114), .B(n77), .Z(n26833) );
  IV U26980 ( .A(n26833), .Z(n26599) );
  NOR U26981 ( .A(n26832), .B(n26599), .Z(n26835) );
  IV U26982 ( .A(n26600), .Z(n26602) );
  XOR U26983 ( .A(n26602), .B(n26601), .Z(n26828) );
  NOR U26984 ( .A(n83), .B(n77), .Z(n26829) );
  IV U26985 ( .A(n26829), .Z(n26603) );
  NOR U26986 ( .A(n26828), .B(n26603), .Z(n26831) );
  IV U26987 ( .A(n26604), .Z(n26606) );
  XOR U26988 ( .A(n26606), .B(n26605), .Z(n26824) );
  NOR U26989 ( .A(n113), .B(n77), .Z(n26825) );
  IV U26990 ( .A(n26825), .Z(n26607) );
  NOR U26991 ( .A(n26824), .B(n26607), .Z(n26827) );
  IV U26992 ( .A(n26608), .Z(n26610) );
  XOR U26993 ( .A(n26610), .B(n26609), .Z(n26820) );
  NOR U26994 ( .A(n84), .B(n77), .Z(n26821) );
  IV U26995 ( .A(n26821), .Z(n26611) );
  NOR U26996 ( .A(n26820), .B(n26611), .Z(n26823) );
  IV U26997 ( .A(n26612), .Z(n26614) );
  XOR U26998 ( .A(n26614), .B(n26613), .Z(n26816) );
  NOR U26999 ( .A(n112), .B(n77), .Z(n26817) );
  IV U27000 ( .A(n26817), .Z(n26615) );
  NOR U27001 ( .A(n26816), .B(n26615), .Z(n26819) );
  IV U27002 ( .A(n26616), .Z(n26618) );
  XOR U27003 ( .A(n26618), .B(n26617), .Z(n26812) );
  NOR U27004 ( .A(n85), .B(n77), .Z(n26813) );
  IV U27005 ( .A(n26813), .Z(n26619) );
  NOR U27006 ( .A(n26812), .B(n26619), .Z(n26815) );
  IV U27007 ( .A(n26620), .Z(n26622) );
  XOR U27008 ( .A(n26622), .B(n26621), .Z(n26808) );
  NOR U27009 ( .A(n111), .B(n77), .Z(n26809) );
  IV U27010 ( .A(n26809), .Z(n26623) );
  NOR U27011 ( .A(n26808), .B(n26623), .Z(n26811) );
  IV U27012 ( .A(n26624), .Z(n26626) );
  XOR U27013 ( .A(n26626), .B(n26625), .Z(n26804) );
  NOR U27014 ( .A(n86), .B(n77), .Z(n26805) );
  IV U27015 ( .A(n26805), .Z(n26627) );
  NOR U27016 ( .A(n26804), .B(n26627), .Z(n26807) );
  IV U27017 ( .A(n26628), .Z(n26630) );
  XOR U27018 ( .A(n26630), .B(n26629), .Z(n26800) );
  NOR U27019 ( .A(n110), .B(n77), .Z(n26801) );
  IV U27020 ( .A(n26801), .Z(n26631) );
  NOR U27021 ( .A(n26800), .B(n26631), .Z(n26803) );
  XOR U27022 ( .A(n26633), .B(n26632), .Z(n26796) );
  NOR U27023 ( .A(n109), .B(n77), .Z(n26797) );
  IV U27024 ( .A(n26797), .Z(n26634) );
  NOR U27025 ( .A(n26796), .B(n26634), .Z(n26799) );
  XOR U27026 ( .A(n26636), .B(n26635), .Z(n26784) );
  IV U27027 ( .A(n26784), .Z(n26638) );
  NOR U27028 ( .A(n87), .B(n77), .Z(n26637) );
  IV U27029 ( .A(n26637), .Z(n26785) );
  NOR U27030 ( .A(n26638), .B(n26785), .Z(n26787) );
  IV U27031 ( .A(n26639), .Z(n26641) );
  XOR U27032 ( .A(n26641), .B(n26640), .Z(n26780) );
  NOR U27033 ( .A(n107), .B(n77), .Z(n26781) );
  IV U27034 ( .A(n26781), .Z(n26642) );
  NOR U27035 ( .A(n26780), .B(n26642), .Z(n26783) );
  IV U27036 ( .A(n26643), .Z(n26645) );
  XOR U27037 ( .A(n26645), .B(n26644), .Z(n26776) );
  NOR U27038 ( .A(n88), .B(n77), .Z(n26777) );
  IV U27039 ( .A(n26777), .Z(n26646) );
  NOR U27040 ( .A(n26776), .B(n26646), .Z(n26779) );
  IV U27041 ( .A(n26647), .Z(n26649) );
  XOR U27042 ( .A(n26649), .B(n26648), .Z(n26772) );
  NOR U27043 ( .A(n106), .B(n77), .Z(n26773) );
  IV U27044 ( .A(n26773), .Z(n26650) );
  NOR U27045 ( .A(n26772), .B(n26650), .Z(n26775) );
  XOR U27046 ( .A(n26652), .B(n26651), .Z(n26768) );
  NOR U27047 ( .A(n105), .B(n77), .Z(n26769) );
  IV U27048 ( .A(n26769), .Z(n26653) );
  NOR U27049 ( .A(n26768), .B(n26653), .Z(n26771) );
  XOR U27050 ( .A(n26655), .B(n26654), .Z(n26756) );
  IV U27051 ( .A(n26756), .Z(n26657) );
  NOR U27052 ( .A(n89), .B(n77), .Z(n26656) );
  IV U27053 ( .A(n26656), .Z(n26757) );
  NOR U27054 ( .A(n26657), .B(n26757), .Z(n26759) );
  IV U27055 ( .A(n26658), .Z(n26660) );
  XOR U27056 ( .A(n26660), .B(n26659), .Z(n26752) );
  NOR U27057 ( .A(n103), .B(n77), .Z(n26753) );
  IV U27058 ( .A(n26753), .Z(n26661) );
  NOR U27059 ( .A(n26752), .B(n26661), .Z(n26755) );
  IV U27060 ( .A(n26662), .Z(n26664) );
  XOR U27061 ( .A(n26664), .B(n26663), .Z(n26748) );
  NOR U27062 ( .A(n90), .B(n77), .Z(n26749) );
  IV U27063 ( .A(n26749), .Z(n26665) );
  NOR U27064 ( .A(n26748), .B(n26665), .Z(n26751) );
  IV U27065 ( .A(n26666), .Z(n26668) );
  XOR U27066 ( .A(n26668), .B(n26667), .Z(n26744) );
  NOR U27067 ( .A(n102), .B(n77), .Z(n26745) );
  IV U27068 ( .A(n26745), .Z(n26669) );
  NOR U27069 ( .A(n26744), .B(n26669), .Z(n26747) );
  IV U27070 ( .A(n26670), .Z(n26672) );
  XOR U27071 ( .A(n26672), .B(n26671), .Z(n26740) );
  NOR U27072 ( .A(n101), .B(n77), .Z(n26741) );
  IV U27073 ( .A(n26741), .Z(n26673) );
  NOR U27074 ( .A(n26740), .B(n26673), .Z(n26743) );
  IV U27075 ( .A(n26674), .Z(n26676) );
  XOR U27076 ( .A(n26676), .B(n26675), .Z(n26736) );
  NOR U27077 ( .A(n100), .B(n77), .Z(n26737) );
  IV U27078 ( .A(n26737), .Z(n26677) );
  NOR U27079 ( .A(n26736), .B(n26677), .Z(n26739) );
  XOR U27080 ( .A(n26679), .B(n26678), .Z(n26680) );
  IV U27081 ( .A(n26680), .Z(n26732) );
  NOR U27082 ( .A(n99), .B(n77), .Z(n26733) );
  IV U27083 ( .A(n26733), .Z(n26681) );
  NOR U27084 ( .A(n26732), .B(n26681), .Z(n26735) );
  IV U27085 ( .A(n26682), .Z(n26684) );
  XOR U27086 ( .A(n26684), .B(n26683), .Z(n26728) );
  NOR U27087 ( .A(n98), .B(n77), .Z(n26729) );
  IV U27088 ( .A(n26729), .Z(n26685) );
  NOR U27089 ( .A(n26728), .B(n26685), .Z(n26731) );
  XOR U27090 ( .A(n26687), .B(n26686), .Z(n26724) );
  NOR U27091 ( .A(n91), .B(n77), .Z(n26725) );
  IV U27092 ( .A(n26725), .Z(n26688) );
  NOR U27093 ( .A(n26724), .B(n26688), .Z(n26727) );
  IV U27094 ( .A(n26689), .Z(n26691) );
  XOR U27095 ( .A(n26691), .B(n26690), .Z(n26720) );
  NOR U27096 ( .A(n97), .B(n77), .Z(n26721) );
  IV U27097 ( .A(n26721), .Z(n26692) );
  NOR U27098 ( .A(n26720), .B(n26692), .Z(n26723) );
  IV U27099 ( .A(n26693), .Z(n26695) );
  XOR U27100 ( .A(n26695), .B(n26694), .Z(n26716) );
  NOR U27101 ( .A(n96), .B(n77), .Z(n26717) );
  IV U27102 ( .A(n26717), .Z(n26696) );
  NOR U27103 ( .A(n26716), .B(n26696), .Z(n26719) );
  NOR U27104 ( .A(n95), .B(n77), .Z(n26713) );
  IV U27105 ( .A(n26713), .Z(n26699) );
  XOR U27106 ( .A(n26698), .B(n26697), .Z(n26712) );
  NOR U27107 ( .A(n26699), .B(n26712), .Z(n26715) );
  NOR U27108 ( .A(n77), .B(n93), .Z(n27699) );
  IV U27109 ( .A(n27699), .Z(n26700) );
  NOR U27110 ( .A(n76), .B(n168), .Z(n26708) );
  IV U27111 ( .A(n26708), .Z(n26703) );
  NOR U27112 ( .A(n26700), .B(n26703), .Z(n26701) );
  IV U27113 ( .A(n26701), .Z(n26702) );
  NOR U27114 ( .A(n94), .B(n26702), .Z(n26711) );
  NOR U27115 ( .A(n26703), .B(n93), .Z(n26704) );
  XOR U27116 ( .A(n94), .B(n26704), .Z(n26705) );
  NOR U27117 ( .A(n77), .B(n26705), .Z(n26706) );
  IV U27118 ( .A(n26706), .Z(n27180) );
  XOR U27119 ( .A(n26708), .B(n26707), .Z(n27179) );
  IV U27120 ( .A(n27179), .Z(n26709) );
  NOR U27121 ( .A(n27180), .B(n26709), .Z(n26710) );
  NOR U27122 ( .A(n26711), .B(n26710), .Z(n27176) );
  XOR U27123 ( .A(n26713), .B(n26712), .Z(n27175) );
  NOR U27124 ( .A(n27176), .B(n27175), .Z(n26714) );
  NOR U27125 ( .A(n26715), .B(n26714), .Z(n27171) );
  XOR U27126 ( .A(n26717), .B(n26716), .Z(n27172) );
  NOR U27127 ( .A(n27171), .B(n27172), .Z(n26718) );
  NOR U27128 ( .A(n26719), .B(n26718), .Z(n27169) );
  XOR U27129 ( .A(n26721), .B(n26720), .Z(n27168) );
  NOR U27130 ( .A(n27169), .B(n27168), .Z(n26722) );
  NOR U27131 ( .A(n26723), .B(n26722), .Z(n27163) );
  XOR U27132 ( .A(n26725), .B(n26724), .Z(n27164) );
  NOR U27133 ( .A(n27163), .B(n27164), .Z(n26726) );
  NOR U27134 ( .A(n26727), .B(n26726), .Z(n27160) );
  XOR U27135 ( .A(n26729), .B(n26728), .Z(n27159) );
  NOR U27136 ( .A(n27160), .B(n27159), .Z(n26730) );
  NOR U27137 ( .A(n26731), .B(n26730), .Z(n27155) );
  XOR U27138 ( .A(n26733), .B(n26732), .Z(n27156) );
  NOR U27139 ( .A(n27155), .B(n27156), .Z(n26734) );
  NOR U27140 ( .A(n26735), .B(n26734), .Z(n27151) );
  XOR U27141 ( .A(n26737), .B(n26736), .Z(n27152) );
  NOR U27142 ( .A(n27151), .B(n27152), .Z(n26738) );
  NOR U27143 ( .A(n26739), .B(n26738), .Z(n27147) );
  XOR U27144 ( .A(n26741), .B(n26740), .Z(n27148) );
  NOR U27145 ( .A(n27147), .B(n27148), .Z(n26742) );
  NOR U27146 ( .A(n26743), .B(n26742), .Z(n27143) );
  XOR U27147 ( .A(n26745), .B(n26744), .Z(n27144) );
  NOR U27148 ( .A(n27143), .B(n27144), .Z(n26746) );
  NOR U27149 ( .A(n26747), .B(n26746), .Z(n27139) );
  XOR U27150 ( .A(n26749), .B(n26748), .Z(n27140) );
  NOR U27151 ( .A(n27139), .B(n27140), .Z(n26750) );
  NOR U27152 ( .A(n26751), .B(n26750), .Z(n27136) );
  XOR U27153 ( .A(n26753), .B(n26752), .Z(n27135) );
  NOR U27154 ( .A(n27136), .B(n27135), .Z(n26754) );
  NOR U27155 ( .A(n26755), .B(n26754), .Z(n27243) );
  XOR U27156 ( .A(n26757), .B(n26756), .Z(n27242) );
  NOR U27157 ( .A(n27243), .B(n27242), .Z(n26758) );
  NOR U27158 ( .A(n26759), .B(n26758), .Z(n26764) );
  XOR U27159 ( .A(n26761), .B(n26760), .Z(n26763) );
  IV U27160 ( .A(n26763), .Z(n26762) );
  NOR U27161 ( .A(n26764), .B(n26762), .Z(n26767) );
  XOR U27162 ( .A(n26764), .B(n26763), .Z(n27132) );
  NOR U27163 ( .A(n104), .B(n77), .Z(n27133) );
  IV U27164 ( .A(n27133), .Z(n26765) );
  NOR U27165 ( .A(n27132), .B(n26765), .Z(n26766) );
  NOR U27166 ( .A(n26767), .B(n26766), .Z(n27128) );
  XOR U27167 ( .A(n26769), .B(n26768), .Z(n27129) );
  NOR U27168 ( .A(n27128), .B(n27129), .Z(n26770) );
  NOR U27169 ( .A(n26771), .B(n26770), .Z(n27124) );
  XOR U27170 ( .A(n26773), .B(n26772), .Z(n27125) );
  NOR U27171 ( .A(n27124), .B(n27125), .Z(n26774) );
  NOR U27172 ( .A(n26775), .B(n26774), .Z(n27120) );
  XOR U27173 ( .A(n26777), .B(n26776), .Z(n27121) );
  NOR U27174 ( .A(n27120), .B(n27121), .Z(n26778) );
  NOR U27175 ( .A(n26779), .B(n26778), .Z(n27117) );
  XOR U27176 ( .A(n26781), .B(n26780), .Z(n27116) );
  NOR U27177 ( .A(n27117), .B(n27116), .Z(n26782) );
  NOR U27178 ( .A(n26783), .B(n26782), .Z(n27271) );
  XOR U27179 ( .A(n26785), .B(n26784), .Z(n27270) );
  NOR U27180 ( .A(n27271), .B(n27270), .Z(n26786) );
  NOR U27181 ( .A(n26787), .B(n26786), .Z(n26790) );
  NOR U27182 ( .A(n108), .B(n77), .Z(n26789) );
  IV U27183 ( .A(n26789), .Z(n26788) );
  NOR U27184 ( .A(n26790), .B(n26788), .Z(n26795) );
  XOR U27185 ( .A(n26790), .B(n26789), .Z(n27113) );
  XOR U27186 ( .A(n26792), .B(n26791), .Z(n27114) );
  IV U27187 ( .A(n27114), .Z(n26793) );
  NOR U27188 ( .A(n27113), .B(n26793), .Z(n26794) );
  NOR U27189 ( .A(n26795), .B(n26794), .Z(n27109) );
  XOR U27190 ( .A(n26797), .B(n26796), .Z(n27110) );
  NOR U27191 ( .A(n27109), .B(n27110), .Z(n26798) );
  NOR U27192 ( .A(n26799), .B(n26798), .Z(n27105) );
  XOR U27193 ( .A(n26801), .B(n26800), .Z(n27106) );
  NOR U27194 ( .A(n27105), .B(n27106), .Z(n26802) );
  NOR U27195 ( .A(n26803), .B(n26802), .Z(n27101) );
  XOR U27196 ( .A(n26805), .B(n26804), .Z(n27102) );
  NOR U27197 ( .A(n27101), .B(n27102), .Z(n26806) );
  NOR U27198 ( .A(n26807), .B(n26806), .Z(n27097) );
  XOR U27199 ( .A(n26809), .B(n26808), .Z(n27098) );
  NOR U27200 ( .A(n27097), .B(n27098), .Z(n26810) );
  NOR U27201 ( .A(n26811), .B(n26810), .Z(n27093) );
  XOR U27202 ( .A(n26813), .B(n26812), .Z(n27094) );
  NOR U27203 ( .A(n27093), .B(n27094), .Z(n26814) );
  NOR U27204 ( .A(n26815), .B(n26814), .Z(n27089) );
  XOR U27205 ( .A(n26817), .B(n26816), .Z(n27090) );
  NOR U27206 ( .A(n27089), .B(n27090), .Z(n26818) );
  NOR U27207 ( .A(n26819), .B(n26818), .Z(n27085) );
  XOR U27208 ( .A(n26821), .B(n26820), .Z(n27086) );
  NOR U27209 ( .A(n27085), .B(n27086), .Z(n26822) );
  NOR U27210 ( .A(n26823), .B(n26822), .Z(n27081) );
  XOR U27211 ( .A(n26825), .B(n26824), .Z(n27082) );
  NOR U27212 ( .A(n27081), .B(n27082), .Z(n26826) );
  NOR U27213 ( .A(n26827), .B(n26826), .Z(n27077) );
  XOR U27214 ( .A(n26829), .B(n26828), .Z(n27078) );
  NOR U27215 ( .A(n27077), .B(n27078), .Z(n26830) );
  NOR U27216 ( .A(n26831), .B(n26830), .Z(n27073) );
  XOR U27217 ( .A(n26833), .B(n26832), .Z(n27074) );
  NOR U27218 ( .A(n27073), .B(n27074), .Z(n26834) );
  NOR U27219 ( .A(n26835), .B(n26834), .Z(n27069) );
  XOR U27220 ( .A(n26837), .B(n26836), .Z(n27070) );
  NOR U27221 ( .A(n27069), .B(n27070), .Z(n26838) );
  NOR U27222 ( .A(n26839), .B(n26838), .Z(n27065) );
  XOR U27223 ( .A(n26841), .B(n26840), .Z(n27066) );
  NOR U27224 ( .A(n27065), .B(n27066), .Z(n26842) );
  NOR U27225 ( .A(n26843), .B(n26842), .Z(n27061) );
  XOR U27226 ( .A(n26845), .B(n26844), .Z(n27062) );
  NOR U27227 ( .A(n27061), .B(n27062), .Z(n26846) );
  NOR U27228 ( .A(n26847), .B(n26846), .Z(n27057) );
  XOR U27229 ( .A(n26849), .B(n26848), .Z(n27058) );
  NOR U27230 ( .A(n27057), .B(n27058), .Z(n26850) );
  NOR U27231 ( .A(n26851), .B(n26850), .Z(n27053) );
  XOR U27232 ( .A(n26853), .B(n26852), .Z(n27054) );
  NOR U27233 ( .A(n27053), .B(n27054), .Z(n26854) );
  NOR U27234 ( .A(n26855), .B(n26854), .Z(n27049) );
  XOR U27235 ( .A(n26857), .B(n26856), .Z(n27050) );
  NOR U27236 ( .A(n27049), .B(n27050), .Z(n26858) );
  NOR U27237 ( .A(n26859), .B(n26858), .Z(n27045) );
  XOR U27238 ( .A(n26861), .B(n26860), .Z(n27046) );
  NOR U27239 ( .A(n27045), .B(n27046), .Z(n26862) );
  NOR U27240 ( .A(n26863), .B(n26862), .Z(n27041) );
  XOR U27241 ( .A(n26865), .B(n26864), .Z(n27042) );
  NOR U27242 ( .A(n27041), .B(n27042), .Z(n26866) );
  NOR U27243 ( .A(n26867), .B(n26866), .Z(n26868) );
  IV U27244 ( .A(n26868), .Z(n27039) );
  XOR U27245 ( .A(n26870), .B(n26869), .Z(n26871) );
  IV U27246 ( .A(n26871), .Z(n27038) );
  NOR U27247 ( .A(n27039), .B(n27038), .Z(n26872) );
  NOR U27248 ( .A(n26873), .B(n26872), .Z(n26874) );
  IV U27249 ( .A(n26874), .Z(n27037) );
  XOR U27250 ( .A(n26876), .B(n26875), .Z(n27036) );
  NOR U27251 ( .A(n27037), .B(n27036), .Z(n26877) );
  NOR U27252 ( .A(n26878), .B(n26877), .Z(n26879) );
  IV U27253 ( .A(n26879), .Z(n27034) );
  XOR U27254 ( .A(n26881), .B(n26880), .Z(n26882) );
  IV U27255 ( .A(n26882), .Z(n27033) );
  NOR U27256 ( .A(n27034), .B(n27033), .Z(n26883) );
  NOR U27257 ( .A(n26884), .B(n26883), .Z(n27031) );
  IV U27258 ( .A(n27031), .Z(n26887) );
  XOR U27259 ( .A(n26886), .B(n26885), .Z(n27030) );
  NOR U27260 ( .A(n26887), .B(n27030), .Z(n26888) );
  NOR U27261 ( .A(n26889), .B(n26888), .Z(n27026) );
  XOR U27262 ( .A(n26891), .B(n26890), .Z(n27027) );
  NOR U27263 ( .A(n27026), .B(n27027), .Z(n26892) );
  NOR U27264 ( .A(n26893), .B(n26892), .Z(n26898) );
  XOR U27265 ( .A(n26895), .B(n26894), .Z(n26897) );
  IV U27266 ( .A(n26897), .Z(n26896) );
  NOR U27267 ( .A(n26898), .B(n26896), .Z(n26901) );
  XOR U27268 ( .A(n26898), .B(n26897), .Z(n27023) );
  NOR U27269 ( .A(n131), .B(n77), .Z(n27024) );
  IV U27270 ( .A(n27024), .Z(n26899) );
  NOR U27271 ( .A(n27023), .B(n26899), .Z(n26900) );
  NOR U27272 ( .A(n26901), .B(n26900), .Z(n27019) );
  XOR U27273 ( .A(n26903), .B(n26902), .Z(n27020) );
  NOR U27274 ( .A(n27019), .B(n27020), .Z(n26904) );
  NOR U27275 ( .A(n26905), .B(n26904), .Z(n27018) );
  XOR U27276 ( .A(n26907), .B(n26906), .Z(n27017) );
  NOR U27277 ( .A(n27018), .B(n27017), .Z(n26908) );
  NOR U27278 ( .A(n26909), .B(n26908), .Z(n27391) );
  XOR U27279 ( .A(n26911), .B(n26910), .Z(n27392) );
  NOR U27280 ( .A(n27391), .B(n27392), .Z(n26912) );
  NOR U27281 ( .A(n26913), .B(n26912), .Z(n27013) );
  XOR U27282 ( .A(n26915), .B(n26914), .Z(n27014) );
  NOR U27283 ( .A(n27013), .B(n27014), .Z(n26916) );
  NOR U27284 ( .A(n26917), .B(n26916), .Z(n27009) );
  XOR U27285 ( .A(n26919), .B(n26918), .Z(n27010) );
  NOR U27286 ( .A(n27009), .B(n27010), .Z(n26920) );
  NOR U27287 ( .A(n26921), .B(n26920), .Z(n27005) );
  XOR U27288 ( .A(n26923), .B(n26922), .Z(n27006) );
  NOR U27289 ( .A(n27005), .B(n27006), .Z(n26924) );
  NOR U27290 ( .A(n26925), .B(n26924), .Z(n27001) );
  XOR U27291 ( .A(n26927), .B(n26926), .Z(n27002) );
  NOR U27292 ( .A(n27001), .B(n27002), .Z(n26928) );
  NOR U27293 ( .A(n26929), .B(n26928), .Z(n26998) );
  XOR U27294 ( .A(n26931), .B(n26930), .Z(n26997) );
  NOR U27295 ( .A(n26998), .B(n26997), .Z(n26932) );
  NOR U27296 ( .A(n26933), .B(n26932), .Z(n26993) );
  XOR U27297 ( .A(n26935), .B(n26934), .Z(n26994) );
  NOR U27298 ( .A(n26993), .B(n26994), .Z(n26936) );
  NOR U27299 ( .A(n26937), .B(n26936), .Z(n26990) );
  XOR U27300 ( .A(n26939), .B(n26938), .Z(n26989) );
  NOR U27301 ( .A(n26990), .B(n26989), .Z(n26940) );
  NOR U27302 ( .A(n26941), .B(n26940), .Z(n26985) );
  XOR U27303 ( .A(n26943), .B(n26942), .Z(n26986) );
  NOR U27304 ( .A(n26985), .B(n26986), .Z(n26944) );
  NOR U27305 ( .A(n26945), .B(n26944), .Z(n26981) );
  XOR U27306 ( .A(n26947), .B(n26946), .Z(n26982) );
  NOR U27307 ( .A(n26981), .B(n26982), .Z(n26948) );
  NOR U27308 ( .A(n26949), .B(n26948), .Z(n26977) );
  IV U27309 ( .A(n26950), .Z(n26979) );
  NOR U27310 ( .A(n26976), .B(n26979), .Z(n26951) );
  NOR U27311 ( .A(n26977), .B(n26951), .Z(n26952) );
  NOR U27312 ( .A(n26953), .B(n26952), .Z(n26955) );
  IV U27313 ( .A(n26955), .Z(n26973) );
  NOR U27314 ( .A(n26970), .B(n26973), .Z(n26958) );
  NOR U27315 ( .A(n158), .B(n77), .Z(n26971) );
  NOR U27316 ( .A(n26955), .B(n26954), .Z(n26956) );
  NOR U27317 ( .A(n26971), .B(n26956), .Z(n26957) );
  NOR U27318 ( .A(n26958), .B(n26957), .Z(n26959) );
  IV U27319 ( .A(n26959), .Z(n26967) );
  NOR U27320 ( .A(n26960), .B(n26967), .Z(n26961) );
  NOR U27321 ( .A(n26962), .B(n26961), .Z(n27457) );
  IV U27322 ( .A(n27457), .Z(n27458) );
  XOR U27323 ( .A(n27456), .B(n27458), .Z(n26963) );
  XOR U27324 ( .A(n27460), .B(n26963), .Z(n27989) );
  IV U27325 ( .A(n27989), .Z(n27448) );
  XOR U27326 ( .A(n26965), .B(n26964), .Z(n26966) );
  XOR U27327 ( .A(n26967), .B(n26966), .Z(n27493) );
  NOR U27328 ( .A(n163), .B(n78), .Z(n26968) );
  IV U27329 ( .A(n26968), .Z(n27492) );
  NOR U27330 ( .A(n27493), .B(n27492), .Z(n27447) );
  IV U27331 ( .A(n27493), .Z(n26969) );
  NOR U27332 ( .A(n26969), .B(n26968), .Z(n27445) );
  XOR U27333 ( .A(n26971), .B(n26970), .Z(n26972) );
  XOR U27334 ( .A(n26973), .B(n26972), .Z(n27500) );
  NOR U27335 ( .A(n161), .B(n78), .Z(n26974) );
  NOR U27336 ( .A(n27500), .B(n26974), .Z(n27443) );
  IV U27337 ( .A(n27500), .Z(n26975) );
  IV U27338 ( .A(n26974), .Z(n27497) );
  NOR U27339 ( .A(n26975), .B(n27497), .Z(n27441) );
  XOR U27340 ( .A(n26977), .B(n26976), .Z(n26978) );
  XOR U27341 ( .A(n26979), .B(n26978), .Z(n27437) );
  NOR U27342 ( .A(n158), .B(n78), .Z(n27436) );
  IV U27343 ( .A(n27436), .Z(n26980) );
  NOR U27344 ( .A(n27437), .B(n26980), .Z(n27439) );
  IV U27345 ( .A(n26981), .Z(n26983) );
  XOR U27346 ( .A(n26983), .B(n26982), .Z(n27432) );
  NOR U27347 ( .A(n156), .B(n78), .Z(n27433) );
  IV U27348 ( .A(n27433), .Z(n26984) );
  NOR U27349 ( .A(n27432), .B(n26984), .Z(n27435) );
  IV U27350 ( .A(n26985), .Z(n26987) );
  XOR U27351 ( .A(n26987), .B(n26986), .Z(n27428) );
  NOR U27352 ( .A(n155), .B(n78), .Z(n27429) );
  IV U27353 ( .A(n27429), .Z(n26988) );
  NOR U27354 ( .A(n27428), .B(n26988), .Z(n27431) );
  XOR U27355 ( .A(n26990), .B(n26989), .Z(n27424) );
  IV U27356 ( .A(n27424), .Z(n26992) );
  NOR U27357 ( .A(n153), .B(n78), .Z(n26991) );
  IV U27358 ( .A(n26991), .Z(n27425) );
  NOR U27359 ( .A(n26992), .B(n27425), .Z(n27427) );
  IV U27360 ( .A(n26993), .Z(n26995) );
  XOR U27361 ( .A(n26995), .B(n26994), .Z(n27420) );
  NOR U27362 ( .A(n150), .B(n78), .Z(n27421) );
  IV U27363 ( .A(n27421), .Z(n26996) );
  NOR U27364 ( .A(n27420), .B(n26996), .Z(n27423) );
  XOR U27365 ( .A(n26998), .B(n26997), .Z(n27416) );
  IV U27366 ( .A(n27416), .Z(n27000) );
  NOR U27367 ( .A(n148), .B(n78), .Z(n26999) );
  IV U27368 ( .A(n26999), .Z(n27417) );
  NOR U27369 ( .A(n27000), .B(n27417), .Z(n27419) );
  IV U27370 ( .A(n27001), .Z(n27003) );
  XOR U27371 ( .A(n27003), .B(n27002), .Z(n27412) );
  NOR U27372 ( .A(n147), .B(n78), .Z(n27413) );
  IV U27373 ( .A(n27413), .Z(n27004) );
  NOR U27374 ( .A(n27412), .B(n27004), .Z(n27415) );
  IV U27375 ( .A(n27005), .Z(n27007) );
  XOR U27376 ( .A(n27007), .B(n27006), .Z(n27408) );
  NOR U27377 ( .A(n145), .B(n78), .Z(n27409) );
  IV U27378 ( .A(n27409), .Z(n27008) );
  NOR U27379 ( .A(n27408), .B(n27008), .Z(n27411) );
  IV U27380 ( .A(n27009), .Z(n27011) );
  XOR U27381 ( .A(n27011), .B(n27010), .Z(n27404) );
  NOR U27382 ( .A(n143), .B(n78), .Z(n27405) );
  IV U27383 ( .A(n27405), .Z(n27012) );
  NOR U27384 ( .A(n27404), .B(n27012), .Z(n27407) );
  IV U27385 ( .A(n27013), .Z(n27015) );
  XOR U27386 ( .A(n27015), .B(n27014), .Z(n27400) );
  NOR U27387 ( .A(n141), .B(n78), .Z(n27401) );
  IV U27388 ( .A(n27401), .Z(n27016) );
  NOR U27389 ( .A(n27400), .B(n27016), .Z(n27403) );
  NOR U27390 ( .A(n137), .B(n78), .Z(n27387) );
  XOR U27391 ( .A(n27018), .B(n27017), .Z(n27386) );
  NOR U27392 ( .A(n27387), .B(n27386), .Z(n27390) );
  IV U27393 ( .A(n27019), .Z(n27021) );
  XOR U27394 ( .A(n27021), .B(n27020), .Z(n27381) );
  NOR U27395 ( .A(n135), .B(n78), .Z(n27382) );
  IV U27396 ( .A(n27382), .Z(n27022) );
  NOR U27397 ( .A(n27381), .B(n27022), .Z(n27384) );
  XOR U27398 ( .A(n27024), .B(n27023), .Z(n27377) );
  NOR U27399 ( .A(n133), .B(n78), .Z(n27378) );
  IV U27400 ( .A(n27378), .Z(n27025) );
  NOR U27401 ( .A(n27377), .B(n27025), .Z(n27380) );
  IV U27402 ( .A(n27026), .Z(n27028) );
  XOR U27403 ( .A(n27028), .B(n27027), .Z(n27373) );
  NOR U27404 ( .A(n131), .B(n78), .Z(n27374) );
  IV U27405 ( .A(n27374), .Z(n27029) );
  NOR U27406 ( .A(n27373), .B(n27029), .Z(n27376) );
  XOR U27407 ( .A(n27031), .B(n27030), .Z(n27369) );
  NOR U27408 ( .A(n128), .B(n78), .Z(n27370) );
  IV U27409 ( .A(n27370), .Z(n27032) );
  NOR U27410 ( .A(n27369), .B(n27032), .Z(n27372) );
  XOR U27411 ( .A(n27034), .B(n27033), .Z(n27366) );
  NOR U27412 ( .A(n126), .B(n78), .Z(n27365) );
  IV U27413 ( .A(n27365), .Z(n27035) );
  NOR U27414 ( .A(n27366), .B(n27035), .Z(n27368) );
  NOR U27415 ( .A(n125), .B(n78), .Z(n27360) );
  XOR U27416 ( .A(n27037), .B(n27036), .Z(n27359) );
  NOR U27417 ( .A(n27360), .B(n27359), .Z(n27363) );
  XOR U27418 ( .A(n27039), .B(n27038), .Z(n27355) );
  NOR U27419 ( .A(n123), .B(n78), .Z(n27354) );
  IV U27420 ( .A(n27354), .Z(n27040) );
  NOR U27421 ( .A(n27355), .B(n27040), .Z(n27357) );
  IV U27422 ( .A(n27041), .Z(n27043) );
  XOR U27423 ( .A(n27043), .B(n27042), .Z(n27350) );
  NOR U27424 ( .A(n120), .B(n78), .Z(n27351) );
  IV U27425 ( .A(n27351), .Z(n27044) );
  NOR U27426 ( .A(n27350), .B(n27044), .Z(n27353) );
  IV U27427 ( .A(n27045), .Z(n27047) );
  XOR U27428 ( .A(n27047), .B(n27046), .Z(n27346) );
  NOR U27429 ( .A(n119), .B(n78), .Z(n27347) );
  IV U27430 ( .A(n27347), .Z(n27048) );
  NOR U27431 ( .A(n27346), .B(n27048), .Z(n27349) );
  IV U27432 ( .A(n27049), .Z(n27051) );
  XOR U27433 ( .A(n27051), .B(n27050), .Z(n27342) );
  NOR U27434 ( .A(n79), .B(n78), .Z(n27343) );
  IV U27435 ( .A(n27343), .Z(n27052) );
  NOR U27436 ( .A(n27342), .B(n27052), .Z(n27345) );
  IV U27437 ( .A(n27053), .Z(n27055) );
  XOR U27438 ( .A(n27055), .B(n27054), .Z(n27338) );
  NOR U27439 ( .A(n117), .B(n78), .Z(n27339) );
  IV U27440 ( .A(n27339), .Z(n27056) );
  NOR U27441 ( .A(n27338), .B(n27056), .Z(n27341) );
  IV U27442 ( .A(n27057), .Z(n27059) );
  XOR U27443 ( .A(n27059), .B(n27058), .Z(n27334) );
  NOR U27444 ( .A(n80), .B(n78), .Z(n27335) );
  IV U27445 ( .A(n27335), .Z(n27060) );
  NOR U27446 ( .A(n27334), .B(n27060), .Z(n27337) );
  IV U27447 ( .A(n27061), .Z(n27063) );
  XOR U27448 ( .A(n27063), .B(n27062), .Z(n27330) );
  NOR U27449 ( .A(n116), .B(n78), .Z(n27331) );
  IV U27450 ( .A(n27331), .Z(n27064) );
  NOR U27451 ( .A(n27330), .B(n27064), .Z(n27333) );
  IV U27452 ( .A(n27065), .Z(n27067) );
  XOR U27453 ( .A(n27067), .B(n27066), .Z(n27326) );
  NOR U27454 ( .A(n81), .B(n78), .Z(n27327) );
  IV U27455 ( .A(n27327), .Z(n27068) );
  NOR U27456 ( .A(n27326), .B(n27068), .Z(n27329) );
  IV U27457 ( .A(n27069), .Z(n27071) );
  XOR U27458 ( .A(n27071), .B(n27070), .Z(n27322) );
  NOR U27459 ( .A(n115), .B(n78), .Z(n27323) );
  IV U27460 ( .A(n27323), .Z(n27072) );
  NOR U27461 ( .A(n27322), .B(n27072), .Z(n27325) );
  IV U27462 ( .A(n27073), .Z(n27075) );
  XOR U27463 ( .A(n27075), .B(n27074), .Z(n27318) );
  NOR U27464 ( .A(n82), .B(n78), .Z(n27319) );
  IV U27465 ( .A(n27319), .Z(n27076) );
  NOR U27466 ( .A(n27318), .B(n27076), .Z(n27321) );
  IV U27467 ( .A(n27077), .Z(n27079) );
  XOR U27468 ( .A(n27079), .B(n27078), .Z(n27314) );
  NOR U27469 ( .A(n114), .B(n78), .Z(n27315) );
  IV U27470 ( .A(n27315), .Z(n27080) );
  NOR U27471 ( .A(n27314), .B(n27080), .Z(n27317) );
  IV U27472 ( .A(n27081), .Z(n27083) );
  XOR U27473 ( .A(n27083), .B(n27082), .Z(n27310) );
  NOR U27474 ( .A(n83), .B(n78), .Z(n27311) );
  IV U27475 ( .A(n27311), .Z(n27084) );
  NOR U27476 ( .A(n27310), .B(n27084), .Z(n27313) );
  IV U27477 ( .A(n27085), .Z(n27087) );
  XOR U27478 ( .A(n27087), .B(n27086), .Z(n27306) );
  NOR U27479 ( .A(n113), .B(n78), .Z(n27307) );
  IV U27480 ( .A(n27307), .Z(n27088) );
  NOR U27481 ( .A(n27306), .B(n27088), .Z(n27309) );
  IV U27482 ( .A(n27089), .Z(n27091) );
  XOR U27483 ( .A(n27091), .B(n27090), .Z(n27302) );
  NOR U27484 ( .A(n84), .B(n78), .Z(n27303) );
  IV U27485 ( .A(n27303), .Z(n27092) );
  NOR U27486 ( .A(n27302), .B(n27092), .Z(n27305) );
  IV U27487 ( .A(n27093), .Z(n27095) );
  XOR U27488 ( .A(n27095), .B(n27094), .Z(n27298) );
  NOR U27489 ( .A(n112), .B(n78), .Z(n27299) );
  IV U27490 ( .A(n27299), .Z(n27096) );
  NOR U27491 ( .A(n27298), .B(n27096), .Z(n27301) );
  IV U27492 ( .A(n27097), .Z(n27099) );
  XOR U27493 ( .A(n27099), .B(n27098), .Z(n27294) );
  NOR U27494 ( .A(n85), .B(n78), .Z(n27295) );
  IV U27495 ( .A(n27295), .Z(n27100) );
  NOR U27496 ( .A(n27294), .B(n27100), .Z(n27297) );
  IV U27497 ( .A(n27101), .Z(n27103) );
  XOR U27498 ( .A(n27103), .B(n27102), .Z(n27290) );
  NOR U27499 ( .A(n111), .B(n78), .Z(n27291) );
  IV U27500 ( .A(n27291), .Z(n27104) );
  NOR U27501 ( .A(n27290), .B(n27104), .Z(n27293) );
  IV U27502 ( .A(n27105), .Z(n27107) );
  XOR U27503 ( .A(n27107), .B(n27106), .Z(n27286) );
  NOR U27504 ( .A(n86), .B(n78), .Z(n27287) );
  IV U27505 ( .A(n27287), .Z(n27108) );
  NOR U27506 ( .A(n27286), .B(n27108), .Z(n27289) );
  IV U27507 ( .A(n27109), .Z(n27111) );
  XOR U27508 ( .A(n27111), .B(n27110), .Z(n27282) );
  NOR U27509 ( .A(n110), .B(n78), .Z(n27283) );
  IV U27510 ( .A(n27283), .Z(n27112) );
  NOR U27511 ( .A(n27282), .B(n27112), .Z(n27285) );
  XOR U27512 ( .A(n27114), .B(n27113), .Z(n27278) );
  NOR U27513 ( .A(n109), .B(n78), .Z(n27279) );
  IV U27514 ( .A(n27279), .Z(n27115) );
  NOR U27515 ( .A(n27278), .B(n27115), .Z(n27281) );
  XOR U27516 ( .A(n27117), .B(n27116), .Z(n27266) );
  IV U27517 ( .A(n27266), .Z(n27119) );
  NOR U27518 ( .A(n87), .B(n78), .Z(n27118) );
  IV U27519 ( .A(n27118), .Z(n27267) );
  NOR U27520 ( .A(n27119), .B(n27267), .Z(n27269) );
  IV U27521 ( .A(n27120), .Z(n27122) );
  XOR U27522 ( .A(n27122), .B(n27121), .Z(n27262) );
  NOR U27523 ( .A(n107), .B(n78), .Z(n27263) );
  IV U27524 ( .A(n27263), .Z(n27123) );
  NOR U27525 ( .A(n27262), .B(n27123), .Z(n27265) );
  IV U27526 ( .A(n27124), .Z(n27126) );
  XOR U27527 ( .A(n27126), .B(n27125), .Z(n27258) );
  NOR U27528 ( .A(n88), .B(n78), .Z(n27259) );
  IV U27529 ( .A(n27259), .Z(n27127) );
  NOR U27530 ( .A(n27258), .B(n27127), .Z(n27261) );
  IV U27531 ( .A(n27128), .Z(n27130) );
  XOR U27532 ( .A(n27130), .B(n27129), .Z(n27254) );
  NOR U27533 ( .A(n106), .B(n78), .Z(n27255) );
  IV U27534 ( .A(n27255), .Z(n27131) );
  NOR U27535 ( .A(n27254), .B(n27131), .Z(n27257) );
  XOR U27536 ( .A(n27133), .B(n27132), .Z(n27250) );
  NOR U27537 ( .A(n105), .B(n78), .Z(n27251) );
  IV U27538 ( .A(n27251), .Z(n27134) );
  NOR U27539 ( .A(n27250), .B(n27134), .Z(n27253) );
  XOR U27540 ( .A(n27136), .B(n27135), .Z(n27238) );
  IV U27541 ( .A(n27238), .Z(n27138) );
  NOR U27542 ( .A(n89), .B(n78), .Z(n27137) );
  IV U27543 ( .A(n27137), .Z(n27239) );
  NOR U27544 ( .A(n27138), .B(n27239), .Z(n27241) );
  IV U27545 ( .A(n27139), .Z(n27141) );
  XOR U27546 ( .A(n27141), .B(n27140), .Z(n27234) );
  NOR U27547 ( .A(n103), .B(n78), .Z(n27235) );
  IV U27548 ( .A(n27235), .Z(n27142) );
  NOR U27549 ( .A(n27234), .B(n27142), .Z(n27237) );
  IV U27550 ( .A(n27143), .Z(n27145) );
  XOR U27551 ( .A(n27145), .B(n27144), .Z(n27230) );
  NOR U27552 ( .A(n90), .B(n78), .Z(n27231) );
  IV U27553 ( .A(n27231), .Z(n27146) );
  NOR U27554 ( .A(n27230), .B(n27146), .Z(n27233) );
  IV U27555 ( .A(n27147), .Z(n27149) );
  XOR U27556 ( .A(n27149), .B(n27148), .Z(n27226) );
  NOR U27557 ( .A(n102), .B(n78), .Z(n27227) );
  IV U27558 ( .A(n27227), .Z(n27150) );
  NOR U27559 ( .A(n27226), .B(n27150), .Z(n27229) );
  IV U27560 ( .A(n27151), .Z(n27153) );
  XOR U27561 ( .A(n27153), .B(n27152), .Z(n27222) );
  NOR U27562 ( .A(n101), .B(n78), .Z(n27223) );
  IV U27563 ( .A(n27223), .Z(n27154) );
  NOR U27564 ( .A(n27222), .B(n27154), .Z(n27225) );
  XOR U27565 ( .A(n27156), .B(n27155), .Z(n27157) );
  IV U27566 ( .A(n27157), .Z(n27218) );
  NOR U27567 ( .A(n100), .B(n78), .Z(n27219) );
  IV U27568 ( .A(n27219), .Z(n27158) );
  NOR U27569 ( .A(n27218), .B(n27158), .Z(n27221) );
  XOR U27570 ( .A(n27160), .B(n27159), .Z(n27214) );
  IV U27571 ( .A(n27214), .Z(n27162) );
  NOR U27572 ( .A(n99), .B(n78), .Z(n27161) );
  IV U27573 ( .A(n27161), .Z(n27215) );
  NOR U27574 ( .A(n27162), .B(n27215), .Z(n27217) );
  XOR U27575 ( .A(n27164), .B(n27163), .Z(n27165) );
  IV U27576 ( .A(n27165), .Z(n27210) );
  NOR U27577 ( .A(n98), .B(n78), .Z(n27211) );
  IV U27578 ( .A(n27211), .Z(n27166) );
  NOR U27579 ( .A(n27210), .B(n27166), .Z(n27213) );
  NOR U27580 ( .A(n91), .B(n78), .Z(n27167) );
  IV U27581 ( .A(n27167), .Z(n27207) );
  XOR U27582 ( .A(n27169), .B(n27168), .Z(n27206) );
  IV U27583 ( .A(n27206), .Z(n27170) );
  NOR U27584 ( .A(n27207), .B(n27170), .Z(n27209) );
  IV U27585 ( .A(n27171), .Z(n27173) );
  XOR U27586 ( .A(n27173), .B(n27172), .Z(n27202) );
  NOR U27587 ( .A(n97), .B(n78), .Z(n27203) );
  IV U27588 ( .A(n27203), .Z(n27174) );
  NOR U27589 ( .A(n27202), .B(n27174), .Z(n27205) );
  XOR U27590 ( .A(n27176), .B(n27175), .Z(n27198) );
  IV U27591 ( .A(n27198), .Z(n27178) );
  NOR U27592 ( .A(n96), .B(n78), .Z(n27177) );
  IV U27593 ( .A(n27177), .Z(n27199) );
  NOR U27594 ( .A(n27178), .B(n27199), .Z(n27201) );
  NOR U27595 ( .A(n95), .B(n78), .Z(n27195) );
  IV U27596 ( .A(n27195), .Z(n27181) );
  XOR U27597 ( .A(n27180), .B(n27179), .Z(n27194) );
  NOR U27598 ( .A(n27181), .B(n27194), .Z(n27197) );
  NOR U27599 ( .A(n78), .B(n93), .Z(n28104) );
  IV U27600 ( .A(n28104), .Z(n27182) );
  NOR U27601 ( .A(n77), .B(n168), .Z(n27190) );
  IV U27602 ( .A(n27190), .Z(n27185) );
  NOR U27603 ( .A(n27182), .B(n27185), .Z(n27183) );
  IV U27604 ( .A(n27183), .Z(n27184) );
  NOR U27605 ( .A(n94), .B(n27184), .Z(n27193) );
  NOR U27606 ( .A(n27185), .B(n93), .Z(n27186) );
  XOR U27607 ( .A(n94), .B(n27186), .Z(n27187) );
  NOR U27608 ( .A(n78), .B(n27187), .Z(n27188) );
  IV U27609 ( .A(n27188), .Z(n27694) );
  XOR U27610 ( .A(n27190), .B(n27189), .Z(n27693) );
  IV U27611 ( .A(n27693), .Z(n27191) );
  NOR U27612 ( .A(n27694), .B(n27191), .Z(n27192) );
  NOR U27613 ( .A(n27193), .B(n27192), .Z(n27689) );
  XOR U27614 ( .A(n27195), .B(n27194), .Z(n27690) );
  NOR U27615 ( .A(n27689), .B(n27690), .Z(n27196) );
  NOR U27616 ( .A(n27197), .B(n27196), .Z(n27718) );
  XOR U27617 ( .A(n27199), .B(n27198), .Z(n27717) );
  NOR U27618 ( .A(n27718), .B(n27717), .Z(n27200) );
  NOR U27619 ( .A(n27201), .B(n27200), .Z(n27685) );
  XOR U27620 ( .A(n27203), .B(n27202), .Z(n27686) );
  NOR U27621 ( .A(n27685), .B(n27686), .Z(n27204) );
  NOR U27622 ( .A(n27205), .B(n27204), .Z(n27729) );
  XOR U27623 ( .A(n27207), .B(n27206), .Z(n27730) );
  NOR U27624 ( .A(n27729), .B(n27730), .Z(n27208) );
  NOR U27625 ( .A(n27209), .B(n27208), .Z(n27681) );
  XOR U27626 ( .A(n27211), .B(n27210), .Z(n27682) );
  NOR U27627 ( .A(n27681), .B(n27682), .Z(n27212) );
  NOR U27628 ( .A(n27213), .B(n27212), .Z(n27745) );
  XOR U27629 ( .A(n27215), .B(n27214), .Z(n27744) );
  NOR U27630 ( .A(n27745), .B(n27744), .Z(n27216) );
  NOR U27631 ( .A(n27217), .B(n27216), .Z(n27677) );
  XOR U27632 ( .A(n27219), .B(n27218), .Z(n27678) );
  NOR U27633 ( .A(n27677), .B(n27678), .Z(n27220) );
  NOR U27634 ( .A(n27221), .B(n27220), .Z(n27673) );
  XOR U27635 ( .A(n27223), .B(n27222), .Z(n27674) );
  NOR U27636 ( .A(n27673), .B(n27674), .Z(n27224) );
  NOR U27637 ( .A(n27225), .B(n27224), .Z(n27669) );
  XOR U27638 ( .A(n27227), .B(n27226), .Z(n27670) );
  NOR U27639 ( .A(n27669), .B(n27670), .Z(n27228) );
  NOR U27640 ( .A(n27229), .B(n27228), .Z(n27665) );
  XOR U27641 ( .A(n27231), .B(n27230), .Z(n27666) );
  NOR U27642 ( .A(n27665), .B(n27666), .Z(n27232) );
  NOR U27643 ( .A(n27233), .B(n27232), .Z(n27661) );
  XOR U27644 ( .A(n27235), .B(n27234), .Z(n27662) );
  NOR U27645 ( .A(n27661), .B(n27662), .Z(n27236) );
  NOR U27646 ( .A(n27237), .B(n27236), .Z(n27774) );
  XOR U27647 ( .A(n27239), .B(n27238), .Z(n27773) );
  NOR U27648 ( .A(n27774), .B(n27773), .Z(n27240) );
  NOR U27649 ( .A(n27241), .B(n27240), .Z(n27246) );
  XOR U27650 ( .A(n27243), .B(n27242), .Z(n27245) );
  IV U27651 ( .A(n27245), .Z(n27244) );
  NOR U27652 ( .A(n27246), .B(n27244), .Z(n27249) );
  XOR U27653 ( .A(n27246), .B(n27245), .Z(n27658) );
  NOR U27654 ( .A(n104), .B(n78), .Z(n27659) );
  IV U27655 ( .A(n27659), .Z(n27247) );
  NOR U27656 ( .A(n27658), .B(n27247), .Z(n27248) );
  NOR U27657 ( .A(n27249), .B(n27248), .Z(n27654) );
  XOR U27658 ( .A(n27251), .B(n27250), .Z(n27655) );
  NOR U27659 ( .A(n27654), .B(n27655), .Z(n27252) );
  NOR U27660 ( .A(n27253), .B(n27252), .Z(n27650) );
  XOR U27661 ( .A(n27255), .B(n27254), .Z(n27651) );
  NOR U27662 ( .A(n27650), .B(n27651), .Z(n27256) );
  NOR U27663 ( .A(n27257), .B(n27256), .Z(n27646) );
  XOR U27664 ( .A(n27259), .B(n27258), .Z(n27647) );
  NOR U27665 ( .A(n27646), .B(n27647), .Z(n27260) );
  NOR U27666 ( .A(n27261), .B(n27260), .Z(n27642) );
  XOR U27667 ( .A(n27263), .B(n27262), .Z(n27643) );
  NOR U27668 ( .A(n27642), .B(n27643), .Z(n27264) );
  NOR U27669 ( .A(n27265), .B(n27264), .Z(n27799) );
  XOR U27670 ( .A(n27267), .B(n27266), .Z(n27798) );
  NOR U27671 ( .A(n27799), .B(n27798), .Z(n27268) );
  NOR U27672 ( .A(n27269), .B(n27268), .Z(n27274) );
  XOR U27673 ( .A(n27271), .B(n27270), .Z(n27273) );
  IV U27674 ( .A(n27273), .Z(n27272) );
  NOR U27675 ( .A(n27274), .B(n27272), .Z(n27277) );
  XOR U27676 ( .A(n27274), .B(n27273), .Z(n27639) );
  NOR U27677 ( .A(n108), .B(n78), .Z(n27640) );
  IV U27678 ( .A(n27640), .Z(n27275) );
  NOR U27679 ( .A(n27639), .B(n27275), .Z(n27276) );
  NOR U27680 ( .A(n27277), .B(n27276), .Z(n27635) );
  XOR U27681 ( .A(n27279), .B(n27278), .Z(n27636) );
  NOR U27682 ( .A(n27635), .B(n27636), .Z(n27280) );
  NOR U27683 ( .A(n27281), .B(n27280), .Z(n27631) );
  XOR U27684 ( .A(n27283), .B(n27282), .Z(n27632) );
  NOR U27685 ( .A(n27631), .B(n27632), .Z(n27284) );
  NOR U27686 ( .A(n27285), .B(n27284), .Z(n27627) );
  XOR U27687 ( .A(n27287), .B(n27286), .Z(n27628) );
  NOR U27688 ( .A(n27627), .B(n27628), .Z(n27288) );
  NOR U27689 ( .A(n27289), .B(n27288), .Z(n27623) );
  XOR U27690 ( .A(n27291), .B(n27290), .Z(n27624) );
  NOR U27691 ( .A(n27623), .B(n27624), .Z(n27292) );
  NOR U27692 ( .A(n27293), .B(n27292), .Z(n27619) );
  XOR U27693 ( .A(n27295), .B(n27294), .Z(n27620) );
  NOR U27694 ( .A(n27619), .B(n27620), .Z(n27296) );
  NOR U27695 ( .A(n27297), .B(n27296), .Z(n27615) );
  XOR U27696 ( .A(n27299), .B(n27298), .Z(n27616) );
  NOR U27697 ( .A(n27615), .B(n27616), .Z(n27300) );
  NOR U27698 ( .A(n27301), .B(n27300), .Z(n27611) );
  XOR U27699 ( .A(n27303), .B(n27302), .Z(n27612) );
  NOR U27700 ( .A(n27611), .B(n27612), .Z(n27304) );
  NOR U27701 ( .A(n27305), .B(n27304), .Z(n27607) );
  XOR U27702 ( .A(n27307), .B(n27306), .Z(n27608) );
  NOR U27703 ( .A(n27607), .B(n27608), .Z(n27308) );
  NOR U27704 ( .A(n27309), .B(n27308), .Z(n27603) );
  XOR U27705 ( .A(n27311), .B(n27310), .Z(n27604) );
  NOR U27706 ( .A(n27603), .B(n27604), .Z(n27312) );
  NOR U27707 ( .A(n27313), .B(n27312), .Z(n27599) );
  XOR U27708 ( .A(n27315), .B(n27314), .Z(n27600) );
  NOR U27709 ( .A(n27599), .B(n27600), .Z(n27316) );
  NOR U27710 ( .A(n27317), .B(n27316), .Z(n27595) );
  XOR U27711 ( .A(n27319), .B(n27318), .Z(n27596) );
  NOR U27712 ( .A(n27595), .B(n27596), .Z(n27320) );
  NOR U27713 ( .A(n27321), .B(n27320), .Z(n27591) );
  XOR U27714 ( .A(n27323), .B(n27322), .Z(n27592) );
  NOR U27715 ( .A(n27591), .B(n27592), .Z(n27324) );
  NOR U27716 ( .A(n27325), .B(n27324), .Z(n27587) );
  XOR U27717 ( .A(n27327), .B(n27326), .Z(n27588) );
  NOR U27718 ( .A(n27587), .B(n27588), .Z(n27328) );
  NOR U27719 ( .A(n27329), .B(n27328), .Z(n27583) );
  XOR U27720 ( .A(n27331), .B(n27330), .Z(n27584) );
  NOR U27721 ( .A(n27583), .B(n27584), .Z(n27332) );
  NOR U27722 ( .A(n27333), .B(n27332), .Z(n27579) );
  XOR U27723 ( .A(n27335), .B(n27334), .Z(n27580) );
  NOR U27724 ( .A(n27579), .B(n27580), .Z(n27336) );
  NOR U27725 ( .A(n27337), .B(n27336), .Z(n27575) );
  XOR U27726 ( .A(n27339), .B(n27338), .Z(n27576) );
  NOR U27727 ( .A(n27575), .B(n27576), .Z(n27340) );
  NOR U27728 ( .A(n27341), .B(n27340), .Z(n27571) );
  XOR U27729 ( .A(n27343), .B(n27342), .Z(n27572) );
  NOR U27730 ( .A(n27571), .B(n27572), .Z(n27344) );
  NOR U27731 ( .A(n27345), .B(n27344), .Z(n27567) );
  XOR U27732 ( .A(n27347), .B(n27346), .Z(n27568) );
  NOR U27733 ( .A(n27567), .B(n27568), .Z(n27348) );
  NOR U27734 ( .A(n27349), .B(n27348), .Z(n27563) );
  XOR U27735 ( .A(n27351), .B(n27350), .Z(n27564) );
  NOR U27736 ( .A(n27563), .B(n27564), .Z(n27352) );
  NOR U27737 ( .A(n27353), .B(n27352), .Z(n27562) );
  XOR U27738 ( .A(n27355), .B(n27354), .Z(n27561) );
  NOR U27739 ( .A(n27562), .B(n27561), .Z(n27356) );
  NOR U27740 ( .A(n27357), .B(n27356), .Z(n27358) );
  IV U27741 ( .A(n27358), .Z(n27559) );
  XOR U27742 ( .A(n27360), .B(n27359), .Z(n27361) );
  IV U27743 ( .A(n27361), .Z(n27558) );
  NOR U27744 ( .A(n27559), .B(n27558), .Z(n27362) );
  NOR U27745 ( .A(n27363), .B(n27362), .Z(n27364) );
  IV U27746 ( .A(n27364), .Z(n27557) );
  XOR U27747 ( .A(n27366), .B(n27365), .Z(n27556) );
  NOR U27748 ( .A(n27557), .B(n27556), .Z(n27367) );
  NOR U27749 ( .A(n27368), .B(n27367), .Z(n27551) );
  XOR U27750 ( .A(n27370), .B(n27369), .Z(n27550) );
  NOR U27751 ( .A(n27551), .B(n27550), .Z(n27371) );
  NOR U27752 ( .A(n27372), .B(n27371), .Z(n27546) );
  XOR U27753 ( .A(n27374), .B(n27373), .Z(n27547) );
  NOR U27754 ( .A(n27546), .B(n27547), .Z(n27375) );
  NOR U27755 ( .A(n27376), .B(n27375), .Z(n27542) );
  XOR U27756 ( .A(n27378), .B(n27377), .Z(n27543) );
  NOR U27757 ( .A(n27542), .B(n27543), .Z(n27379) );
  NOR U27758 ( .A(n27380), .B(n27379), .Z(n27541) );
  XOR U27759 ( .A(n27382), .B(n27381), .Z(n27540) );
  NOR U27760 ( .A(n27541), .B(n27540), .Z(n27383) );
  NOR U27761 ( .A(n27384), .B(n27383), .Z(n27385) );
  IV U27762 ( .A(n27385), .Z(n27536) );
  XOR U27763 ( .A(n27387), .B(n27386), .Z(n27388) );
  IV U27764 ( .A(n27388), .Z(n27535) );
  NOR U27765 ( .A(n27536), .B(n27535), .Z(n27389) );
  NOR U27766 ( .A(n27390), .B(n27389), .Z(n27396) );
  IV U27767 ( .A(n27396), .Z(n27394) );
  IV U27768 ( .A(n27391), .Z(n27393) );
  XOR U27769 ( .A(n27393), .B(n27392), .Z(n27395) );
  NOR U27770 ( .A(n27394), .B(n27395), .Z(n27399) );
  XOR U27771 ( .A(n27396), .B(n27395), .Z(n27531) );
  NOR U27772 ( .A(n139), .B(n78), .Z(n27397) );
  IV U27773 ( .A(n27397), .Z(n27530) );
  NOR U27774 ( .A(n27531), .B(n27530), .Z(n27398) );
  NOR U27775 ( .A(n27399), .B(n27398), .Z(n27926) );
  XOR U27776 ( .A(n27401), .B(n27400), .Z(n27927) );
  NOR U27777 ( .A(n27926), .B(n27927), .Z(n27402) );
  NOR U27778 ( .A(n27403), .B(n27402), .Z(n27526) );
  XOR U27779 ( .A(n27405), .B(n27404), .Z(n27527) );
  NOR U27780 ( .A(n27526), .B(n27527), .Z(n27406) );
  NOR U27781 ( .A(n27407), .B(n27406), .Z(n27522) );
  XOR U27782 ( .A(n27409), .B(n27408), .Z(n27523) );
  NOR U27783 ( .A(n27522), .B(n27523), .Z(n27410) );
  NOR U27784 ( .A(n27411), .B(n27410), .Z(n27518) );
  XOR U27785 ( .A(n27413), .B(n27412), .Z(n27519) );
  NOR U27786 ( .A(n27518), .B(n27519), .Z(n27414) );
  NOR U27787 ( .A(n27415), .B(n27414), .Z(n27948) );
  XOR U27788 ( .A(n27417), .B(n27416), .Z(n27947) );
  NOR U27789 ( .A(n27948), .B(n27947), .Z(n27418) );
  NOR U27790 ( .A(n27419), .B(n27418), .Z(n27514) );
  XOR U27791 ( .A(n27421), .B(n27420), .Z(n27515) );
  NOR U27792 ( .A(n27514), .B(n27515), .Z(n27422) );
  NOR U27793 ( .A(n27423), .B(n27422), .Z(n27960) );
  XOR U27794 ( .A(n27425), .B(n27424), .Z(n27959) );
  NOR U27795 ( .A(n27960), .B(n27959), .Z(n27426) );
  NOR U27796 ( .A(n27427), .B(n27426), .Z(n27510) );
  XOR U27797 ( .A(n27429), .B(n27428), .Z(n27511) );
  NOR U27798 ( .A(n27510), .B(n27511), .Z(n27430) );
  NOR U27799 ( .A(n27431), .B(n27430), .Z(n27506) );
  XOR U27800 ( .A(n27433), .B(n27432), .Z(n27507) );
  NOR U27801 ( .A(n27506), .B(n27507), .Z(n27434) );
  NOR U27802 ( .A(n27435), .B(n27434), .Z(n27502) );
  XOR U27803 ( .A(n27437), .B(n27436), .Z(n27503) );
  NOR U27804 ( .A(n27502), .B(n27503), .Z(n27438) );
  NOR U27805 ( .A(n27439), .B(n27438), .Z(n27440) );
  IV U27806 ( .A(n27440), .Z(n27498) );
  NOR U27807 ( .A(n27441), .B(n27498), .Z(n27442) );
  NOR U27808 ( .A(n27443), .B(n27442), .Z(n27444) );
  IV U27809 ( .A(n27444), .Z(n27495) );
  NOR U27810 ( .A(n27445), .B(n27495), .Z(n27446) );
  NOR U27811 ( .A(n27447), .B(n27446), .Z(n27992) );
  NOR U27812 ( .A(n27448), .B(n27992), .Z(n27453) );
  IV U27813 ( .A(n27992), .Z(n27449) );
  NOR U27814 ( .A(n27989), .B(n27449), .Z(n27451) );
  NOR U27815 ( .A(n165), .B(n78), .Z(n27450) );
  IV U27816 ( .A(n27450), .Z(n27990) );
  NOR U27817 ( .A(n27451), .B(n27990), .Z(n27452) );
  NOR U27818 ( .A(n27453), .B(n27452), .Z(n27491) );
  XOR U27819 ( .A(n27455), .B(n27454), .Z(n27471) );
  NOR U27820 ( .A(n165), .B(n77), .Z(n27467) );
  IV U27821 ( .A(n27467), .Z(n27468) );
  NOR U27822 ( .A(n27457), .B(n27456), .Z(n27463) );
  NOR U27823 ( .A(n27459), .B(n27458), .Z(n27461) );
  NOR U27824 ( .A(n27461), .B(n27460), .Z(n27462) );
  NOR U27825 ( .A(n27463), .B(n27462), .Z(n27469) );
  IV U27826 ( .A(n27469), .Z(n27466) );
  XOR U27827 ( .A(n27468), .B(n27466), .Z(n27464) );
  XOR U27828 ( .A(n27471), .B(n27464), .Z(n27488) );
  NOR U27829 ( .A(n167), .B(n78), .Z(n27465) );
  IV U27830 ( .A(n27465), .Z(n27489) );
  NOR U27831 ( .A(n27467), .B(n27466), .Z(n27473) );
  NOR U27832 ( .A(n27469), .B(n27468), .Z(n27470) );
  NOR U27833 ( .A(n27471), .B(n27470), .Z(n27472) );
  NOR U27834 ( .A(n27473), .B(n27472), .Z(n27479) );
  NOR U27835 ( .A(n167), .B(n77), .Z(n27474) );
  IV U27836 ( .A(n27474), .Z(n27480) );
  XOR U27837 ( .A(n27479), .B(n27480), .Z(n27482) );
  XOR U27838 ( .A(n27476), .B(n27475), .Z(n27477) );
  XOR U27839 ( .A(n27478), .B(n27477), .Z(n27483) );
  XOR U27840 ( .A(n27482), .B(n27483), .Z(n28003) );
  XOR U27841 ( .A(n28005), .B(n28003), .Z(n31465) );
  IV U27842 ( .A(n27479), .Z(n27481) );
  NOR U27843 ( .A(n27481), .B(n27480), .Z(n27485) );
  NOR U27844 ( .A(n27483), .B(n27482), .Z(n27484) );
  NOR U27845 ( .A(n27485), .B(n27484), .Z(n27999) );
  XOR U27846 ( .A(n27487), .B(n27486), .Z(n27997) );
  XOR U27847 ( .A(n27999), .B(n27997), .Z(n31469) );
  XOR U27848 ( .A(n27489), .B(n27488), .Z(n27490) );
  XOR U27849 ( .A(n27491), .B(n27490), .Z(n28500) );
  NOR U27850 ( .A(n167), .B(n92), .Z(n27987) );
  NOR U27851 ( .A(n165), .B(n92), .Z(n27984) );
  IV U27852 ( .A(n27984), .Z(n27496) );
  XOR U27853 ( .A(n27493), .B(n27492), .Z(n27494) );
  XOR U27854 ( .A(n27495), .B(n27494), .Z(n27983) );
  NOR U27855 ( .A(n27496), .B(n27983), .Z(n27986) );
  XOR U27856 ( .A(n27498), .B(n27497), .Z(n27499) );
  XOR U27857 ( .A(n27500), .B(n27499), .Z(n27979) );
  NOR U27858 ( .A(n163), .B(n92), .Z(n27980) );
  IV U27859 ( .A(n27980), .Z(n27501) );
  NOR U27860 ( .A(n27979), .B(n27501), .Z(n27982) );
  IV U27861 ( .A(n27502), .Z(n27504) );
  XOR U27862 ( .A(n27504), .B(n27503), .Z(n27975) );
  NOR U27863 ( .A(n161), .B(n92), .Z(n27976) );
  IV U27864 ( .A(n27976), .Z(n27505) );
  NOR U27865 ( .A(n27975), .B(n27505), .Z(n27978) );
  IV U27866 ( .A(n27506), .Z(n27508) );
  XOR U27867 ( .A(n27508), .B(n27507), .Z(n27971) );
  NOR U27868 ( .A(n158), .B(n92), .Z(n27972) );
  IV U27869 ( .A(n27972), .Z(n27509) );
  NOR U27870 ( .A(n27971), .B(n27509), .Z(n27974) );
  IV U27871 ( .A(n27510), .Z(n27512) );
  XOR U27872 ( .A(n27512), .B(n27511), .Z(n27967) );
  NOR U27873 ( .A(n156), .B(n92), .Z(n27968) );
  IV U27874 ( .A(n27968), .Z(n27513) );
  NOR U27875 ( .A(n27967), .B(n27513), .Z(n27970) );
  IV U27876 ( .A(n27514), .Z(n27516) );
  XOR U27877 ( .A(n27516), .B(n27515), .Z(n27955) );
  NOR U27878 ( .A(n153), .B(n92), .Z(n27956) );
  IV U27879 ( .A(n27956), .Z(n27517) );
  NOR U27880 ( .A(n27955), .B(n27517), .Z(n27958) );
  IV U27881 ( .A(n27518), .Z(n27520) );
  XOR U27882 ( .A(n27520), .B(n27519), .Z(n27943) );
  NOR U27883 ( .A(n148), .B(n92), .Z(n27944) );
  IV U27884 ( .A(n27944), .Z(n27521) );
  NOR U27885 ( .A(n27943), .B(n27521), .Z(n27946) );
  IV U27886 ( .A(n27522), .Z(n27524) );
  XOR U27887 ( .A(n27524), .B(n27523), .Z(n27939) );
  NOR U27888 ( .A(n147), .B(n92), .Z(n27940) );
  IV U27889 ( .A(n27940), .Z(n27525) );
  NOR U27890 ( .A(n27939), .B(n27525), .Z(n27942) );
  IV U27891 ( .A(n27526), .Z(n27528) );
  XOR U27892 ( .A(n27528), .B(n27527), .Z(n27935) );
  NOR U27893 ( .A(n145), .B(n92), .Z(n27936) );
  IV U27894 ( .A(n27936), .Z(n27529) );
  NOR U27895 ( .A(n27935), .B(n27529), .Z(n27938) );
  NOR U27896 ( .A(n141), .B(n92), .Z(n27533) );
  XOR U27897 ( .A(n27531), .B(n27530), .Z(n27532) );
  NOR U27898 ( .A(n27533), .B(n27532), .Z(n27925) );
  XOR U27899 ( .A(n27533), .B(n27532), .Z(n27534) );
  IV U27900 ( .A(n27534), .Z(n28024) );
  XOR U27901 ( .A(n27536), .B(n27535), .Z(n27539) );
  NOR U27902 ( .A(n139), .B(n92), .Z(n27538) );
  IV U27903 ( .A(n27538), .Z(n27537) );
  NOR U27904 ( .A(n27539), .B(n27537), .Z(n27922) );
  XOR U27905 ( .A(n27539), .B(n27538), .Z(n28405) );
  NOR U27906 ( .A(n137), .B(n92), .Z(n27916) );
  XOR U27907 ( .A(n27541), .B(n27540), .Z(n27915) );
  NOR U27908 ( .A(n27916), .B(n27915), .Z(n27919) );
  IV U27909 ( .A(n27542), .Z(n27544) );
  XOR U27910 ( .A(n27544), .B(n27543), .Z(n27910) );
  NOR U27911 ( .A(n135), .B(n92), .Z(n27911) );
  IV U27912 ( .A(n27911), .Z(n27545) );
  NOR U27913 ( .A(n27910), .B(n27545), .Z(n27913) );
  IV U27914 ( .A(n27546), .Z(n27548) );
  XOR U27915 ( .A(n27548), .B(n27547), .Z(n27906) );
  NOR U27916 ( .A(n133), .B(n92), .Z(n27907) );
  IV U27917 ( .A(n27907), .Z(n27549) );
  NOR U27918 ( .A(n27906), .B(n27549), .Z(n27909) );
  XOR U27919 ( .A(n27551), .B(n27550), .Z(n27554) );
  IV U27920 ( .A(n27554), .Z(n27553) );
  NOR U27921 ( .A(n131), .B(n92), .Z(n27552) );
  IV U27922 ( .A(n27552), .Z(n27555) );
  NOR U27923 ( .A(n27553), .B(n27555), .Z(n27905) );
  XOR U27924 ( .A(n27555), .B(n27554), .Z(n28031) );
  NOR U27925 ( .A(n128), .B(n92), .Z(n27899) );
  XOR U27926 ( .A(n27557), .B(n27556), .Z(n27898) );
  NOR U27927 ( .A(n27899), .B(n27898), .Z(n27902) );
  XOR U27928 ( .A(n27559), .B(n27558), .Z(n27894) );
  NOR U27929 ( .A(n126), .B(n92), .Z(n27893) );
  IV U27930 ( .A(n27893), .Z(n27560) );
  NOR U27931 ( .A(n27894), .B(n27560), .Z(n27896) );
  NOR U27932 ( .A(n125), .B(n92), .Z(n27888) );
  XOR U27933 ( .A(n27562), .B(n27561), .Z(n27887) );
  NOR U27934 ( .A(n27888), .B(n27887), .Z(n27891) );
  IV U27935 ( .A(n27563), .Z(n27565) );
  XOR U27936 ( .A(n27565), .B(n27564), .Z(n27882) );
  NOR U27937 ( .A(n123), .B(n92), .Z(n27883) );
  IV U27938 ( .A(n27883), .Z(n27566) );
  NOR U27939 ( .A(n27882), .B(n27566), .Z(n27885) );
  IV U27940 ( .A(n27567), .Z(n27569) );
  XOR U27941 ( .A(n27569), .B(n27568), .Z(n27878) );
  NOR U27942 ( .A(n120), .B(n92), .Z(n27879) );
  IV U27943 ( .A(n27879), .Z(n27570) );
  NOR U27944 ( .A(n27878), .B(n27570), .Z(n27881) );
  IV U27945 ( .A(n27571), .Z(n27573) );
  XOR U27946 ( .A(n27573), .B(n27572), .Z(n27874) );
  NOR U27947 ( .A(n119), .B(n92), .Z(n27875) );
  IV U27948 ( .A(n27875), .Z(n27574) );
  NOR U27949 ( .A(n27874), .B(n27574), .Z(n27877) );
  IV U27950 ( .A(n27575), .Z(n27577) );
  XOR U27951 ( .A(n27577), .B(n27576), .Z(n27870) );
  NOR U27952 ( .A(n79), .B(n92), .Z(n27871) );
  IV U27953 ( .A(n27871), .Z(n27578) );
  NOR U27954 ( .A(n27870), .B(n27578), .Z(n27873) );
  IV U27955 ( .A(n27579), .Z(n27581) );
  XOR U27956 ( .A(n27581), .B(n27580), .Z(n27866) );
  NOR U27957 ( .A(n117), .B(n92), .Z(n27867) );
  IV U27958 ( .A(n27867), .Z(n27582) );
  NOR U27959 ( .A(n27866), .B(n27582), .Z(n27869) );
  IV U27960 ( .A(n27583), .Z(n27585) );
  XOR U27961 ( .A(n27585), .B(n27584), .Z(n27862) );
  NOR U27962 ( .A(n80), .B(n92), .Z(n27863) );
  IV U27963 ( .A(n27863), .Z(n27586) );
  NOR U27964 ( .A(n27862), .B(n27586), .Z(n27865) );
  IV U27965 ( .A(n27587), .Z(n27589) );
  XOR U27966 ( .A(n27589), .B(n27588), .Z(n27858) );
  NOR U27967 ( .A(n116), .B(n92), .Z(n27859) );
  IV U27968 ( .A(n27859), .Z(n27590) );
  NOR U27969 ( .A(n27858), .B(n27590), .Z(n27861) );
  IV U27970 ( .A(n27591), .Z(n27593) );
  XOR U27971 ( .A(n27593), .B(n27592), .Z(n27854) );
  NOR U27972 ( .A(n81), .B(n92), .Z(n27855) );
  IV U27973 ( .A(n27855), .Z(n27594) );
  NOR U27974 ( .A(n27854), .B(n27594), .Z(n27857) );
  IV U27975 ( .A(n27595), .Z(n27597) );
  XOR U27976 ( .A(n27597), .B(n27596), .Z(n27850) );
  NOR U27977 ( .A(n115), .B(n92), .Z(n27851) );
  IV U27978 ( .A(n27851), .Z(n27598) );
  NOR U27979 ( .A(n27850), .B(n27598), .Z(n27853) );
  IV U27980 ( .A(n27599), .Z(n27601) );
  XOR U27981 ( .A(n27601), .B(n27600), .Z(n27846) );
  NOR U27982 ( .A(n82), .B(n92), .Z(n27847) );
  IV U27983 ( .A(n27847), .Z(n27602) );
  NOR U27984 ( .A(n27846), .B(n27602), .Z(n27849) );
  IV U27985 ( .A(n27603), .Z(n27605) );
  XOR U27986 ( .A(n27605), .B(n27604), .Z(n27842) );
  NOR U27987 ( .A(n114), .B(n92), .Z(n27843) );
  IV U27988 ( .A(n27843), .Z(n27606) );
  NOR U27989 ( .A(n27842), .B(n27606), .Z(n27845) );
  IV U27990 ( .A(n27607), .Z(n27609) );
  XOR U27991 ( .A(n27609), .B(n27608), .Z(n27838) );
  NOR U27992 ( .A(n83), .B(n92), .Z(n27839) );
  IV U27993 ( .A(n27839), .Z(n27610) );
  NOR U27994 ( .A(n27838), .B(n27610), .Z(n27841) );
  IV U27995 ( .A(n27611), .Z(n27613) );
  XOR U27996 ( .A(n27613), .B(n27612), .Z(n27834) );
  NOR U27997 ( .A(n113), .B(n92), .Z(n27835) );
  IV U27998 ( .A(n27835), .Z(n27614) );
  NOR U27999 ( .A(n27834), .B(n27614), .Z(n27837) );
  IV U28000 ( .A(n27615), .Z(n27617) );
  XOR U28001 ( .A(n27617), .B(n27616), .Z(n27830) );
  NOR U28002 ( .A(n84), .B(n92), .Z(n27831) );
  IV U28003 ( .A(n27831), .Z(n27618) );
  NOR U28004 ( .A(n27830), .B(n27618), .Z(n27833) );
  IV U28005 ( .A(n27619), .Z(n27621) );
  XOR U28006 ( .A(n27621), .B(n27620), .Z(n27826) );
  NOR U28007 ( .A(n112), .B(n92), .Z(n27827) );
  IV U28008 ( .A(n27827), .Z(n27622) );
  NOR U28009 ( .A(n27826), .B(n27622), .Z(n27829) );
  IV U28010 ( .A(n27623), .Z(n27625) );
  XOR U28011 ( .A(n27625), .B(n27624), .Z(n27822) );
  NOR U28012 ( .A(n85), .B(n92), .Z(n27823) );
  IV U28013 ( .A(n27823), .Z(n27626) );
  NOR U28014 ( .A(n27822), .B(n27626), .Z(n27825) );
  IV U28015 ( .A(n27627), .Z(n27629) );
  XOR U28016 ( .A(n27629), .B(n27628), .Z(n27818) );
  NOR U28017 ( .A(n111), .B(n92), .Z(n27819) );
  IV U28018 ( .A(n27819), .Z(n27630) );
  NOR U28019 ( .A(n27818), .B(n27630), .Z(n27821) );
  IV U28020 ( .A(n27631), .Z(n27633) );
  XOR U28021 ( .A(n27633), .B(n27632), .Z(n27814) );
  NOR U28022 ( .A(n86), .B(n92), .Z(n27815) );
  IV U28023 ( .A(n27815), .Z(n27634) );
  NOR U28024 ( .A(n27814), .B(n27634), .Z(n27817) );
  IV U28025 ( .A(n27635), .Z(n27637) );
  XOR U28026 ( .A(n27637), .B(n27636), .Z(n27810) );
  NOR U28027 ( .A(n110), .B(n92), .Z(n27811) );
  IV U28028 ( .A(n27811), .Z(n27638) );
  NOR U28029 ( .A(n27810), .B(n27638), .Z(n27813) );
  XOR U28030 ( .A(n27640), .B(n27639), .Z(n27806) );
  NOR U28031 ( .A(n109), .B(n92), .Z(n27807) );
  IV U28032 ( .A(n27807), .Z(n27641) );
  NOR U28033 ( .A(n27806), .B(n27641), .Z(n27809) );
  IV U28034 ( .A(n27642), .Z(n27644) );
  XOR U28035 ( .A(n27644), .B(n27643), .Z(n27794) );
  NOR U28036 ( .A(n87), .B(n92), .Z(n27795) );
  IV U28037 ( .A(n27795), .Z(n27645) );
  NOR U28038 ( .A(n27794), .B(n27645), .Z(n27797) );
  IV U28039 ( .A(n27646), .Z(n27648) );
  XOR U28040 ( .A(n27648), .B(n27647), .Z(n27790) );
  NOR U28041 ( .A(n107), .B(n92), .Z(n27791) );
  IV U28042 ( .A(n27791), .Z(n27649) );
  NOR U28043 ( .A(n27790), .B(n27649), .Z(n27793) );
  IV U28044 ( .A(n27650), .Z(n27652) );
  XOR U28045 ( .A(n27652), .B(n27651), .Z(n27786) );
  NOR U28046 ( .A(n88), .B(n92), .Z(n27787) );
  IV U28047 ( .A(n27787), .Z(n27653) );
  NOR U28048 ( .A(n27786), .B(n27653), .Z(n27789) );
  IV U28049 ( .A(n27654), .Z(n27656) );
  XOR U28050 ( .A(n27656), .B(n27655), .Z(n27782) );
  NOR U28051 ( .A(n106), .B(n92), .Z(n27783) );
  IV U28052 ( .A(n27783), .Z(n27657) );
  NOR U28053 ( .A(n27782), .B(n27657), .Z(n27785) );
  XOR U28054 ( .A(n27659), .B(n27658), .Z(n27778) );
  NOR U28055 ( .A(n105), .B(n92), .Z(n27779) );
  IV U28056 ( .A(n27779), .Z(n27660) );
  NOR U28057 ( .A(n27778), .B(n27660), .Z(n27781) );
  IV U28058 ( .A(n27661), .Z(n27663) );
  XOR U28059 ( .A(n27663), .B(n27662), .Z(n27766) );
  NOR U28060 ( .A(n89), .B(n92), .Z(n27767) );
  IV U28061 ( .A(n27767), .Z(n27664) );
  NOR U28062 ( .A(n27766), .B(n27664), .Z(n27769) );
  IV U28063 ( .A(n27665), .Z(n27667) );
  XOR U28064 ( .A(n27667), .B(n27666), .Z(n27762) );
  NOR U28065 ( .A(n103), .B(n92), .Z(n27763) );
  IV U28066 ( .A(n27763), .Z(n27668) );
  NOR U28067 ( .A(n27762), .B(n27668), .Z(n27765) );
  IV U28068 ( .A(n27669), .Z(n27671) );
  XOR U28069 ( .A(n27671), .B(n27670), .Z(n27758) );
  NOR U28070 ( .A(n90), .B(n92), .Z(n27759) );
  IV U28071 ( .A(n27759), .Z(n27672) );
  NOR U28072 ( .A(n27758), .B(n27672), .Z(n27761) );
  IV U28073 ( .A(n27673), .Z(n27675) );
  XOR U28074 ( .A(n27675), .B(n27674), .Z(n27754) );
  NOR U28075 ( .A(n102), .B(n92), .Z(n27755) );
  IV U28076 ( .A(n27755), .Z(n27676) );
  NOR U28077 ( .A(n27754), .B(n27676), .Z(n27757) );
  XOR U28078 ( .A(n27678), .B(n27677), .Z(n27679) );
  IV U28079 ( .A(n27679), .Z(n27749) );
  NOR U28080 ( .A(n101), .B(n92), .Z(n27680) );
  IV U28081 ( .A(n27680), .Z(n27750) );
  NOR U28082 ( .A(n27749), .B(n27750), .Z(n27753) );
  IV U28083 ( .A(n27681), .Z(n27683) );
  XOR U28084 ( .A(n27683), .B(n27682), .Z(n27737) );
  NOR U28085 ( .A(n99), .B(n92), .Z(n27738) );
  IV U28086 ( .A(n27738), .Z(n27684) );
  NOR U28087 ( .A(n27737), .B(n27684), .Z(n27740) );
  IV U28088 ( .A(n27685), .Z(n27687) );
  XOR U28089 ( .A(n27687), .B(n27686), .Z(n27724) );
  NOR U28090 ( .A(n91), .B(n92), .Z(n27688) );
  IV U28091 ( .A(n27688), .Z(n27725) );
  NOR U28092 ( .A(n27724), .B(n27725), .Z(n27728) );
  IV U28093 ( .A(n27689), .Z(n27691) );
  XOR U28094 ( .A(n27691), .B(n27690), .Z(n27712) );
  NOR U28095 ( .A(n96), .B(n92), .Z(n27713) );
  IV U28096 ( .A(n27713), .Z(n27692) );
  NOR U28097 ( .A(n27712), .B(n27692), .Z(n27715) );
  XOR U28098 ( .A(n27694), .B(n27693), .Z(n27708) );
  NOR U28099 ( .A(n95), .B(n92), .Z(n27709) );
  IV U28100 ( .A(n27709), .Z(n27695) );
  NOR U28101 ( .A(n27708), .B(n27695), .Z(n27711) );
  NOR U28102 ( .A(n93), .B(n92), .Z(n31831) );
  IV U28103 ( .A(n31831), .Z(n27696) );
  NOR U28104 ( .A(n78), .B(n168), .Z(n27700) );
  IV U28105 ( .A(n27700), .Z(n27701) );
  NOR U28106 ( .A(n27696), .B(n27701), .Z(n27697) );
  IV U28107 ( .A(n27697), .Z(n27698) );
  NOR U28108 ( .A(n94), .B(n27698), .Z(n27707) );
  XOR U28109 ( .A(n27700), .B(n27699), .Z(n28110) );
  IV U28110 ( .A(n28110), .Z(n27705) );
  NOR U28111 ( .A(n27701), .B(n93), .Z(n27702) );
  XOR U28112 ( .A(n94), .B(n27702), .Z(n27703) );
  NOR U28113 ( .A(n92), .B(n27703), .Z(n27704) );
  IV U28114 ( .A(n27704), .Z(n28111) );
  NOR U28115 ( .A(n27705), .B(n28111), .Z(n27706) );
  NOR U28116 ( .A(n27707), .B(n27706), .Z(n28119) );
  XOR U28117 ( .A(n27709), .B(n27708), .Z(n28118) );
  NOR U28118 ( .A(n28119), .B(n28118), .Z(n27710) );
  NOR U28119 ( .A(n27711), .B(n27710), .Z(n28129) );
  XOR U28120 ( .A(n27713), .B(n27712), .Z(n28130) );
  NOR U28121 ( .A(n28129), .B(n28130), .Z(n27714) );
  NOR U28122 ( .A(n27715), .B(n27714), .Z(n27720) );
  NOR U28123 ( .A(n97), .B(n92), .Z(n27719) );
  IV U28124 ( .A(n27719), .Z(n27716) );
  NOR U28125 ( .A(n27720), .B(n27716), .Z(n27723) );
  XOR U28126 ( .A(n27718), .B(n27717), .Z(n28096) );
  IV U28127 ( .A(n28096), .Z(n27721) );
  XOR U28128 ( .A(n27720), .B(n27719), .Z(n28095) );
  NOR U28129 ( .A(n27721), .B(n28095), .Z(n27722) );
  NOR U28130 ( .A(n27723), .B(n27722), .Z(n28139) );
  XOR U28131 ( .A(n27725), .B(n27724), .Z(n28140) );
  IV U28132 ( .A(n28140), .Z(n27726) );
  NOR U28133 ( .A(n28139), .B(n27726), .Z(n27727) );
  NOR U28134 ( .A(n27728), .B(n27727), .Z(n27733) );
  XOR U28135 ( .A(n27730), .B(n27729), .Z(n27732) );
  IV U28136 ( .A(n27732), .Z(n27731) );
  NOR U28137 ( .A(n27733), .B(n27731), .Z(n27736) );
  XOR U28138 ( .A(n27733), .B(n27732), .Z(n28146) );
  NOR U28139 ( .A(n98), .B(n92), .Z(n28147) );
  IV U28140 ( .A(n28147), .Z(n27734) );
  NOR U28141 ( .A(n28146), .B(n27734), .Z(n27735) );
  NOR U28142 ( .A(n27736), .B(n27735), .Z(n28155) );
  XOR U28143 ( .A(n27738), .B(n27737), .Z(n28156) );
  NOR U28144 ( .A(n28155), .B(n28156), .Z(n27739) );
  NOR U28145 ( .A(n27740), .B(n27739), .Z(n27743) );
  NOR U28146 ( .A(n100), .B(n92), .Z(n27742) );
  IV U28147 ( .A(n27742), .Z(n27741) );
  NOR U28148 ( .A(n27743), .B(n27741), .Z(n27748) );
  XOR U28149 ( .A(n27743), .B(n27742), .Z(n28161) );
  XOR U28150 ( .A(n27745), .B(n27744), .Z(n28162) );
  IV U28151 ( .A(n28162), .Z(n27746) );
  NOR U28152 ( .A(n28161), .B(n27746), .Z(n27747) );
  NOR U28153 ( .A(n27748), .B(n27747), .Z(n28170) );
  XOR U28154 ( .A(n27750), .B(n27749), .Z(n28171) );
  IV U28155 ( .A(n28171), .Z(n27751) );
  NOR U28156 ( .A(n28170), .B(n27751), .Z(n27752) );
  NOR U28157 ( .A(n27753), .B(n27752), .Z(n28091) );
  XOR U28158 ( .A(n27755), .B(n27754), .Z(n28092) );
  NOR U28159 ( .A(n28091), .B(n28092), .Z(n27756) );
  NOR U28160 ( .A(n27757), .B(n27756), .Z(n28181) );
  XOR U28161 ( .A(n27759), .B(n27758), .Z(n28182) );
  NOR U28162 ( .A(n28181), .B(n28182), .Z(n27760) );
  NOR U28163 ( .A(n27761), .B(n27760), .Z(n28087) );
  XOR U28164 ( .A(n27763), .B(n27762), .Z(n28088) );
  NOR U28165 ( .A(n28087), .B(n28088), .Z(n27764) );
  NOR U28166 ( .A(n27765), .B(n27764), .Z(n28193) );
  XOR U28167 ( .A(n27767), .B(n27766), .Z(n28194) );
  NOR U28168 ( .A(n28193), .B(n28194), .Z(n27768) );
  NOR U28169 ( .A(n27769), .B(n27768), .Z(n27772) );
  NOR U28170 ( .A(n104), .B(n92), .Z(n27771) );
  IV U28171 ( .A(n27771), .Z(n27770) );
  NOR U28172 ( .A(n27772), .B(n27770), .Z(n27777) );
  XOR U28173 ( .A(n27772), .B(n27771), .Z(n28201) );
  XOR U28174 ( .A(n27774), .B(n27773), .Z(n28202) );
  IV U28175 ( .A(n28202), .Z(n27775) );
  NOR U28176 ( .A(n28201), .B(n27775), .Z(n27776) );
  NOR U28177 ( .A(n27777), .B(n27776), .Z(n28206) );
  XOR U28178 ( .A(n27779), .B(n27778), .Z(n28207) );
  NOR U28179 ( .A(n28206), .B(n28207), .Z(n27780) );
  NOR U28180 ( .A(n27781), .B(n27780), .Z(n28083) );
  XOR U28181 ( .A(n27783), .B(n27782), .Z(n28084) );
  NOR U28182 ( .A(n28083), .B(n28084), .Z(n27784) );
  NOR U28183 ( .A(n27785), .B(n27784), .Z(n28220) );
  XOR U28184 ( .A(n27787), .B(n27786), .Z(n28221) );
  NOR U28185 ( .A(n28220), .B(n28221), .Z(n27788) );
  NOR U28186 ( .A(n27789), .B(n27788), .Z(n28079) );
  XOR U28187 ( .A(n27791), .B(n27790), .Z(n28080) );
  NOR U28188 ( .A(n28079), .B(n28080), .Z(n27792) );
  NOR U28189 ( .A(n27793), .B(n27792), .Z(n28232) );
  XOR U28190 ( .A(n27795), .B(n27794), .Z(n28233) );
  NOR U28191 ( .A(n28232), .B(n28233), .Z(n27796) );
  NOR U28192 ( .A(n27797), .B(n27796), .Z(n27802) );
  XOR U28193 ( .A(n27799), .B(n27798), .Z(n27801) );
  IV U28194 ( .A(n27801), .Z(n27800) );
  NOR U28195 ( .A(n27802), .B(n27800), .Z(n27805) );
  XOR U28196 ( .A(n27802), .B(n27801), .Z(n28240) );
  NOR U28197 ( .A(n108), .B(n92), .Z(n28241) );
  IV U28198 ( .A(n28241), .Z(n27803) );
  NOR U28199 ( .A(n28240), .B(n27803), .Z(n27804) );
  NOR U28200 ( .A(n27805), .B(n27804), .Z(n28245) );
  XOR U28201 ( .A(n27807), .B(n27806), .Z(n28246) );
  NOR U28202 ( .A(n28245), .B(n28246), .Z(n27808) );
  NOR U28203 ( .A(n27809), .B(n27808), .Z(n28075) );
  XOR U28204 ( .A(n27811), .B(n27810), .Z(n28076) );
  NOR U28205 ( .A(n28075), .B(n28076), .Z(n27812) );
  NOR U28206 ( .A(n27813), .B(n27812), .Z(n28259) );
  XOR U28207 ( .A(n27815), .B(n27814), .Z(n28260) );
  NOR U28208 ( .A(n28259), .B(n28260), .Z(n27816) );
  NOR U28209 ( .A(n27817), .B(n27816), .Z(n28071) );
  XOR U28210 ( .A(n27819), .B(n27818), .Z(n28072) );
  NOR U28211 ( .A(n28071), .B(n28072), .Z(n27820) );
  NOR U28212 ( .A(n27821), .B(n27820), .Z(n28271) );
  XOR U28213 ( .A(n27823), .B(n27822), .Z(n28272) );
  NOR U28214 ( .A(n28271), .B(n28272), .Z(n27824) );
  NOR U28215 ( .A(n27825), .B(n27824), .Z(n28067) );
  XOR U28216 ( .A(n27827), .B(n27826), .Z(n28068) );
  NOR U28217 ( .A(n28067), .B(n28068), .Z(n27828) );
  NOR U28218 ( .A(n27829), .B(n27828), .Z(n28283) );
  XOR U28219 ( .A(n27831), .B(n27830), .Z(n28284) );
  NOR U28220 ( .A(n28283), .B(n28284), .Z(n27832) );
  NOR U28221 ( .A(n27833), .B(n27832), .Z(n28063) );
  XOR U28222 ( .A(n27835), .B(n27834), .Z(n28064) );
  NOR U28223 ( .A(n28063), .B(n28064), .Z(n27836) );
  NOR U28224 ( .A(n27837), .B(n27836), .Z(n28295) );
  XOR U28225 ( .A(n27839), .B(n27838), .Z(n28296) );
  NOR U28226 ( .A(n28295), .B(n28296), .Z(n27840) );
  NOR U28227 ( .A(n27841), .B(n27840), .Z(n28059) );
  XOR U28228 ( .A(n27843), .B(n27842), .Z(n28060) );
  NOR U28229 ( .A(n28059), .B(n28060), .Z(n27844) );
  NOR U28230 ( .A(n27845), .B(n27844), .Z(n28307) );
  XOR U28231 ( .A(n27847), .B(n27846), .Z(n28308) );
  NOR U28232 ( .A(n28307), .B(n28308), .Z(n27848) );
  NOR U28233 ( .A(n27849), .B(n27848), .Z(n28055) );
  XOR U28234 ( .A(n27851), .B(n27850), .Z(n28056) );
  NOR U28235 ( .A(n28055), .B(n28056), .Z(n27852) );
  NOR U28236 ( .A(n27853), .B(n27852), .Z(n28319) );
  XOR U28237 ( .A(n27855), .B(n27854), .Z(n28320) );
  NOR U28238 ( .A(n28319), .B(n28320), .Z(n27856) );
  NOR U28239 ( .A(n27857), .B(n27856), .Z(n28051) );
  XOR U28240 ( .A(n27859), .B(n27858), .Z(n28052) );
  NOR U28241 ( .A(n28051), .B(n28052), .Z(n27860) );
  NOR U28242 ( .A(n27861), .B(n27860), .Z(n28331) );
  XOR U28243 ( .A(n27863), .B(n27862), .Z(n28332) );
  NOR U28244 ( .A(n28331), .B(n28332), .Z(n27864) );
  NOR U28245 ( .A(n27865), .B(n27864), .Z(n28047) );
  XOR U28246 ( .A(n27867), .B(n27866), .Z(n28048) );
  NOR U28247 ( .A(n28047), .B(n28048), .Z(n27868) );
  NOR U28248 ( .A(n27869), .B(n27868), .Z(n28343) );
  XOR U28249 ( .A(n27871), .B(n27870), .Z(n28344) );
  NOR U28250 ( .A(n28343), .B(n28344), .Z(n27872) );
  NOR U28251 ( .A(n27873), .B(n27872), .Z(n28043) );
  XOR U28252 ( .A(n27875), .B(n27874), .Z(n28044) );
  NOR U28253 ( .A(n28043), .B(n28044), .Z(n27876) );
  NOR U28254 ( .A(n27877), .B(n27876), .Z(n28355) );
  XOR U28255 ( .A(n27879), .B(n27878), .Z(n28356) );
  NOR U28256 ( .A(n28355), .B(n28356), .Z(n27880) );
  NOR U28257 ( .A(n27881), .B(n27880), .Z(n28039) );
  XOR U28258 ( .A(n27883), .B(n27882), .Z(n28040) );
  NOR U28259 ( .A(n28039), .B(n28040), .Z(n27884) );
  NOR U28260 ( .A(n27885), .B(n27884), .Z(n27886) );
  IV U28261 ( .A(n27886), .Z(n28366) );
  XOR U28262 ( .A(n27888), .B(n27887), .Z(n27889) );
  IV U28263 ( .A(n27889), .Z(n28365) );
  NOR U28264 ( .A(n28366), .B(n28365), .Z(n27890) );
  NOR U28265 ( .A(n27891), .B(n27890), .Z(n27892) );
  IV U28266 ( .A(n27892), .Z(n28038) );
  XOR U28267 ( .A(n27894), .B(n27893), .Z(n28037) );
  NOR U28268 ( .A(n28038), .B(n28037), .Z(n27895) );
  NOR U28269 ( .A(n27896), .B(n27895), .Z(n27897) );
  IV U28270 ( .A(n27897), .Z(n28033) );
  XOR U28271 ( .A(n27899), .B(n27898), .Z(n27900) );
  IV U28272 ( .A(n27900), .Z(n28032) );
  NOR U28273 ( .A(n28033), .B(n28032), .Z(n27901) );
  NOR U28274 ( .A(n27902), .B(n27901), .Z(n27903) );
  IV U28275 ( .A(n27903), .Z(n28030) );
  NOR U28276 ( .A(n28031), .B(n28030), .Z(n27904) );
  NOR U28277 ( .A(n27905), .B(n27904), .Z(n28389) );
  XOR U28278 ( .A(n27907), .B(n27906), .Z(n28390) );
  NOR U28279 ( .A(n28389), .B(n28390), .Z(n27908) );
  NOR U28280 ( .A(n27909), .B(n27908), .Z(n28026) );
  XOR U28281 ( .A(n27911), .B(n27910), .Z(n28027) );
  NOR U28282 ( .A(n28026), .B(n28027), .Z(n27912) );
  NOR U28283 ( .A(n27913), .B(n27912), .Z(n27914) );
  IV U28284 ( .A(n27914), .Z(n28400) );
  XOR U28285 ( .A(n27916), .B(n27915), .Z(n27917) );
  IV U28286 ( .A(n27917), .Z(n28399) );
  NOR U28287 ( .A(n28400), .B(n28399), .Z(n27918) );
  NOR U28288 ( .A(n27919), .B(n27918), .Z(n28406) );
  IV U28289 ( .A(n28406), .Z(n27920) );
  NOR U28290 ( .A(n28405), .B(n27920), .Z(n27921) );
  NOR U28291 ( .A(n27922), .B(n27921), .Z(n27923) );
  IV U28292 ( .A(n27923), .Z(n28023) );
  NOR U28293 ( .A(n28024), .B(n28023), .Z(n27924) );
  NOR U28294 ( .A(n27925), .B(n27924), .Z(n27931) );
  IV U28295 ( .A(n27931), .Z(n27929) );
  IV U28296 ( .A(n27926), .Z(n27928) );
  XOR U28297 ( .A(n27928), .B(n27927), .Z(n27930) );
  NOR U28298 ( .A(n27929), .B(n27930), .Z(n27934) );
  XOR U28299 ( .A(n27931), .B(n27930), .Z(n28417) );
  NOR U28300 ( .A(n143), .B(n92), .Z(n28418) );
  IV U28301 ( .A(n28418), .Z(n27932) );
  NOR U28302 ( .A(n28417), .B(n27932), .Z(n27933) );
  NOR U28303 ( .A(n27934), .B(n27933), .Z(n28428) );
  XOR U28304 ( .A(n27936), .B(n27935), .Z(n28429) );
  NOR U28305 ( .A(n28428), .B(n28429), .Z(n27937) );
  NOR U28306 ( .A(n27938), .B(n27937), .Z(n28022) );
  XOR U28307 ( .A(n27940), .B(n27939), .Z(n28021) );
  NOR U28308 ( .A(n28022), .B(n28021), .Z(n27941) );
  NOR U28309 ( .A(n27942), .B(n27941), .Z(n28443) );
  XOR U28310 ( .A(n27944), .B(n27943), .Z(n28444) );
  NOR U28311 ( .A(n28443), .B(n28444), .Z(n27945) );
  NOR U28312 ( .A(n27946), .B(n27945), .Z(n27951) );
  XOR U28313 ( .A(n27948), .B(n27947), .Z(n27950) );
  IV U28314 ( .A(n27950), .Z(n27949) );
  NOR U28315 ( .A(n27951), .B(n27949), .Z(n27954) );
  XOR U28316 ( .A(n27951), .B(n27950), .Z(n28018) );
  NOR U28317 ( .A(n150), .B(n92), .Z(n28019) );
  IV U28318 ( .A(n28019), .Z(n27952) );
  NOR U28319 ( .A(n28018), .B(n27952), .Z(n27953) );
  NOR U28320 ( .A(n27954), .B(n27953), .Z(n28455) );
  XOR U28321 ( .A(n27956), .B(n27955), .Z(n28454) );
  NOR U28322 ( .A(n28455), .B(n28454), .Z(n27957) );
  NOR U28323 ( .A(n27958), .B(n27957), .Z(n27963) );
  XOR U28324 ( .A(n27960), .B(n27959), .Z(n27962) );
  IV U28325 ( .A(n27962), .Z(n27961) );
  NOR U28326 ( .A(n27963), .B(n27961), .Z(n27966) );
  XOR U28327 ( .A(n27963), .B(n27962), .Z(n28459) );
  NOR U28328 ( .A(n155), .B(n92), .Z(n28460) );
  IV U28329 ( .A(n28460), .Z(n27964) );
  NOR U28330 ( .A(n28459), .B(n27964), .Z(n27965) );
  NOR U28331 ( .A(n27966), .B(n27965), .Z(n28469) );
  XOR U28332 ( .A(n27968), .B(n27967), .Z(n28470) );
  NOR U28333 ( .A(n28469), .B(n28470), .Z(n27969) );
  NOR U28334 ( .A(n27970), .B(n27969), .Z(n28017) );
  XOR U28335 ( .A(n27972), .B(n27971), .Z(n28016) );
  NOR U28336 ( .A(n28017), .B(n28016), .Z(n27973) );
  NOR U28337 ( .A(n27974), .B(n27973), .Z(n28010) );
  XOR U28338 ( .A(n27976), .B(n27975), .Z(n28011) );
  NOR U28339 ( .A(n28010), .B(n28011), .Z(n27977) );
  NOR U28340 ( .A(n27978), .B(n27977), .Z(n28006) );
  XOR U28341 ( .A(n27980), .B(n27979), .Z(n28007) );
  NOR U28342 ( .A(n28006), .B(n28007), .Z(n27981) );
  NOR U28343 ( .A(n27982), .B(n27981), .Z(n28489) );
  XOR U28344 ( .A(n27984), .B(n27983), .Z(n28488) );
  NOR U28345 ( .A(n28489), .B(n28488), .Z(n27985) );
  NOR U28346 ( .A(n27986), .B(n27985), .Z(n27988) );
  IV U28347 ( .A(n27988), .Z(n28496) );
  NOR U28348 ( .A(n27987), .B(n28496), .Z(n27995) );
  IV U28349 ( .A(n27987), .Z(n28495) );
  NOR U28350 ( .A(n27988), .B(n28495), .Z(n27993) );
  XOR U28351 ( .A(n27990), .B(n27989), .Z(n27991) );
  XOR U28352 ( .A(n27992), .B(n27991), .Z(n28498) );
  NOR U28353 ( .A(n27993), .B(n28498), .Z(n27994) );
  NOR U28354 ( .A(n27995), .B(n27994), .Z(n28501) );
  IV U28355 ( .A(n28501), .Z(n27996) );
  NOR U28356 ( .A(n28500), .B(n27996), .Z(n31464) );
  IV U28357 ( .A(n27997), .Z(n27998) );
  NOR U28358 ( .A(n27999), .B(n27998), .Z(n28502) );
  IV U28359 ( .A(n28502), .Z(n31473) );
  XOR U28360 ( .A(n28001), .B(n28000), .Z(n31472) );
  IV U28361 ( .A(n31472), .Z(n28002) );
  NOR U28362 ( .A(n31473), .B(n28002), .Z(n31477) );
  IV U28363 ( .A(n28003), .Z(n28004) );
  NOR U28364 ( .A(n28005), .B(n28004), .Z(n31468) );
  XOR U28365 ( .A(n28007), .B(n28006), .Z(n31815) );
  IV U28366 ( .A(n31815), .Z(n28008) );
  NOR U28367 ( .A(n165), .B(n169), .Z(n28009) );
  IV U28368 ( .A(n28009), .Z(n31817) );
  NOR U28369 ( .A(n28008), .B(n31817), .Z(n28486) );
  NOR U28370 ( .A(n31815), .B(n28009), .Z(n28484) );
  IV U28371 ( .A(n28010), .Z(n28012) );
  XOR U28372 ( .A(n28012), .B(n28011), .Z(n28014) );
  NOR U28373 ( .A(n163), .B(n169), .Z(n28015) );
  IV U28374 ( .A(n28015), .Z(n28013) );
  NOR U28375 ( .A(n28014), .B(n28013), .Z(n28483) );
  XOR U28376 ( .A(n28015), .B(n28014), .Z(n31811) );
  NOR U28377 ( .A(n161), .B(n169), .Z(n28477) );
  XOR U28378 ( .A(n28017), .B(n28016), .Z(n28476) );
  NOR U28379 ( .A(n28477), .B(n28476), .Z(n28480) );
  NOR U28380 ( .A(n155), .B(n169), .Z(n31799) );
  XOR U28381 ( .A(n28019), .B(n28018), .Z(n28448) );
  NOR U28382 ( .A(n153), .B(n169), .Z(n28449) );
  IV U28383 ( .A(n28449), .Z(n28020) );
  NOR U28384 ( .A(n28448), .B(n28020), .Z(n28451) );
  NOR U28385 ( .A(n148), .B(n169), .Z(n28435) );
  XOR U28386 ( .A(n28022), .B(n28021), .Z(n28434) );
  NOR U28387 ( .A(n28435), .B(n28434), .Z(n28438) );
  XOR U28388 ( .A(n28024), .B(n28023), .Z(n28414) );
  NOR U28389 ( .A(n143), .B(n169), .Z(n28413) );
  IV U28390 ( .A(n28413), .Z(n28025) );
  NOR U28391 ( .A(n28414), .B(n28025), .Z(n28416) );
  IV U28392 ( .A(n28026), .Z(n28028) );
  XOR U28393 ( .A(n28028), .B(n28027), .Z(n28394) );
  NOR U28394 ( .A(n137), .B(n169), .Z(n28395) );
  IV U28395 ( .A(n28395), .Z(n28029) );
  NOR U28396 ( .A(n28394), .B(n28029), .Z(n28397) );
  XOR U28397 ( .A(n28031), .B(n28030), .Z(n28382) );
  XOR U28398 ( .A(n28033), .B(n28032), .Z(n28036) );
  NOR U28399 ( .A(n131), .B(n169), .Z(n28035) );
  IV U28400 ( .A(n28035), .Z(n28034) );
  NOR U28401 ( .A(n28036), .B(n28034), .Z(n28379) );
  XOR U28402 ( .A(n28036), .B(n28035), .Z(n31772) );
  NOR U28403 ( .A(n128), .B(n169), .Z(n28371) );
  XOR U28404 ( .A(n28038), .B(n28037), .Z(n28372) );
  NOR U28405 ( .A(n28371), .B(n28372), .Z(n28376) );
  IV U28406 ( .A(n28039), .Z(n28041) );
  XOR U28407 ( .A(n28041), .B(n28040), .Z(n28360) );
  NOR U28408 ( .A(n125), .B(n169), .Z(n28361) );
  IV U28409 ( .A(n28361), .Z(n28042) );
  NOR U28410 ( .A(n28360), .B(n28042), .Z(n28363) );
  IV U28411 ( .A(n28043), .Z(n28045) );
  XOR U28412 ( .A(n28045), .B(n28044), .Z(n28348) );
  NOR U28413 ( .A(n120), .B(n169), .Z(n28349) );
  IV U28414 ( .A(n28349), .Z(n28046) );
  NOR U28415 ( .A(n28348), .B(n28046), .Z(n28351) );
  IV U28416 ( .A(n28047), .Z(n28049) );
  XOR U28417 ( .A(n28049), .B(n28048), .Z(n28336) );
  NOR U28418 ( .A(n79), .B(n169), .Z(n28337) );
  IV U28419 ( .A(n28337), .Z(n28050) );
  NOR U28420 ( .A(n28336), .B(n28050), .Z(n28339) );
  IV U28421 ( .A(n28051), .Z(n28053) );
  XOR U28422 ( .A(n28053), .B(n28052), .Z(n28324) );
  NOR U28423 ( .A(n80), .B(n169), .Z(n28325) );
  IV U28424 ( .A(n28325), .Z(n28054) );
  NOR U28425 ( .A(n28324), .B(n28054), .Z(n28327) );
  IV U28426 ( .A(n28055), .Z(n28057) );
  XOR U28427 ( .A(n28057), .B(n28056), .Z(n28312) );
  NOR U28428 ( .A(n81), .B(n169), .Z(n28313) );
  IV U28429 ( .A(n28313), .Z(n28058) );
  NOR U28430 ( .A(n28312), .B(n28058), .Z(n28315) );
  IV U28431 ( .A(n28059), .Z(n28061) );
  XOR U28432 ( .A(n28061), .B(n28060), .Z(n28300) );
  NOR U28433 ( .A(n82), .B(n169), .Z(n28301) );
  IV U28434 ( .A(n28301), .Z(n28062) );
  NOR U28435 ( .A(n28300), .B(n28062), .Z(n28303) );
  IV U28436 ( .A(n28063), .Z(n28065) );
  XOR U28437 ( .A(n28065), .B(n28064), .Z(n28288) );
  NOR U28438 ( .A(n83), .B(n169), .Z(n28289) );
  IV U28439 ( .A(n28289), .Z(n28066) );
  NOR U28440 ( .A(n28288), .B(n28066), .Z(n28291) );
  IV U28441 ( .A(n28067), .Z(n28069) );
  XOR U28442 ( .A(n28069), .B(n28068), .Z(n28276) );
  NOR U28443 ( .A(n84), .B(n169), .Z(n28277) );
  IV U28444 ( .A(n28277), .Z(n28070) );
  NOR U28445 ( .A(n28276), .B(n28070), .Z(n28279) );
  IV U28446 ( .A(n28071), .Z(n28073) );
  XOR U28447 ( .A(n28073), .B(n28072), .Z(n28264) );
  NOR U28448 ( .A(n85), .B(n169), .Z(n28265) );
  IV U28449 ( .A(n28265), .Z(n28074) );
  NOR U28450 ( .A(n28264), .B(n28074), .Z(n28267) );
  IV U28451 ( .A(n28075), .Z(n28077) );
  XOR U28452 ( .A(n28077), .B(n28076), .Z(n28252) );
  NOR U28453 ( .A(n86), .B(n169), .Z(n28253) );
  IV U28454 ( .A(n28253), .Z(n28078) );
  NOR U28455 ( .A(n28252), .B(n28078), .Z(n28255) );
  IV U28456 ( .A(n28079), .Z(n28081) );
  XOR U28457 ( .A(n28081), .B(n28080), .Z(n28225) );
  NOR U28458 ( .A(n87), .B(n169), .Z(n28226) );
  IV U28459 ( .A(n28226), .Z(n28082) );
  NOR U28460 ( .A(n28225), .B(n28082), .Z(n28228) );
  IV U28461 ( .A(n28083), .Z(n28085) );
  XOR U28462 ( .A(n28085), .B(n28084), .Z(n28213) );
  NOR U28463 ( .A(n88), .B(n169), .Z(n28214) );
  IV U28464 ( .A(n28214), .Z(n28086) );
  NOR U28465 ( .A(n28213), .B(n28086), .Z(n28216) );
  IV U28466 ( .A(n28087), .Z(n28089) );
  XOR U28467 ( .A(n28089), .B(n28088), .Z(n28186) );
  NOR U28468 ( .A(n89), .B(n169), .Z(n28187) );
  IV U28469 ( .A(n28187), .Z(n28090) );
  NOR U28470 ( .A(n28186), .B(n28090), .Z(n28189) );
  IV U28471 ( .A(n28091), .Z(n28093) );
  XOR U28472 ( .A(n28093), .B(n28092), .Z(n28174) );
  NOR U28473 ( .A(n90), .B(n169), .Z(n28175) );
  IV U28474 ( .A(n28175), .Z(n28094) );
  NOR U28475 ( .A(n28174), .B(n28094), .Z(n28177) );
  XOR U28476 ( .A(n28096), .B(n28095), .Z(n28134) );
  NOR U28477 ( .A(n91), .B(n169), .Z(n28135) );
  IV U28478 ( .A(n28135), .Z(n28097) );
  NOR U28479 ( .A(n28134), .B(n28097), .Z(n28137) );
  NOR U28480 ( .A(n92), .B(n168), .Z(n28105) );
  IV U28481 ( .A(n28105), .Z(n28101) );
  NOR U28482 ( .A(n93), .B(n169), .Z(c[0]) );
  IV U28483 ( .A(c[0]), .Z(n28098) );
  NOR U28484 ( .A(n28101), .B(n28098), .Z(n28099) );
  IV U28485 ( .A(n28099), .Z(n28100) );
  NOR U28486 ( .A(n94), .B(n28100), .Z(n28109) );
  NOR U28487 ( .A(n28101), .B(n93), .Z(n28102) );
  XOR U28488 ( .A(n94), .B(n28102), .Z(n28103) );
  NOR U28489 ( .A(n169), .B(n28103), .Z(n31698) );
  IV U28490 ( .A(n31698), .Z(n28107) );
  XOR U28491 ( .A(n28105), .B(n28104), .Z(n31697) );
  IV U28492 ( .A(n31697), .Z(n28106) );
  NOR U28493 ( .A(n28107), .B(n28106), .Z(n28108) );
  NOR U28494 ( .A(n28109), .B(n28108), .Z(n28112) );
  XOR U28495 ( .A(n28111), .B(n28110), .Z(n28113) );
  NOR U28496 ( .A(n28112), .B(n28113), .Z(n28117) );
  IV U28497 ( .A(n28112), .Z(n28114) );
  XOR U28498 ( .A(n28114), .B(n28113), .Z(n31720) );
  NOR U28499 ( .A(n95), .B(n169), .Z(n28115) );
  IV U28500 ( .A(n28115), .Z(n31719) );
  NOR U28501 ( .A(n31720), .B(n31719), .Z(n28116) );
  NOR U28502 ( .A(n28117), .B(n28116), .Z(n28122) );
  XOR U28503 ( .A(n28119), .B(n28118), .Z(n28121) );
  IV U28504 ( .A(n28121), .Z(n28120) );
  NOR U28505 ( .A(n28122), .B(n28120), .Z(n28125) );
  XOR U28506 ( .A(n28122), .B(n28121), .Z(n31742) );
  NOR U28507 ( .A(n96), .B(n169), .Z(n28123) );
  IV U28508 ( .A(n28123), .Z(n31741) );
  NOR U28509 ( .A(n31742), .B(n31741), .Z(n28124) );
  NOR U28510 ( .A(n28125), .B(n28124), .Z(n28128) );
  NOR U28511 ( .A(n97), .B(n169), .Z(n28127) );
  IV U28512 ( .A(n28127), .Z(n28126) );
  NOR U28513 ( .A(n28128), .B(n28126), .Z(n28133) );
  XOR U28514 ( .A(n28128), .B(n28127), .Z(n31764) );
  IV U28515 ( .A(n28129), .Z(n28131) );
  XOR U28516 ( .A(n28131), .B(n28130), .Z(n31763) );
  NOR U28517 ( .A(n31764), .B(n31763), .Z(n28132) );
  NOR U28518 ( .A(n28133), .B(n28132), .Z(n31787) );
  XOR U28519 ( .A(n28135), .B(n28134), .Z(n31786) );
  NOR U28520 ( .A(n31787), .B(n31786), .Z(n28136) );
  NOR U28521 ( .A(n28137), .B(n28136), .Z(n28142) );
  NOR U28522 ( .A(n98), .B(n169), .Z(n28141) );
  IV U28523 ( .A(n28141), .Z(n28138) );
  NOR U28524 ( .A(n28142), .B(n28138), .Z(n28144) );
  XOR U28525 ( .A(n28140), .B(n28139), .Z(n31813) );
  XOR U28526 ( .A(n28142), .B(n28141), .Z(n31812) );
  NOR U28527 ( .A(n31813), .B(n31812), .Z(n28143) );
  NOR U28528 ( .A(n28144), .B(n28143), .Z(n28149) );
  NOR U28529 ( .A(n99), .B(n169), .Z(n28148) );
  IV U28530 ( .A(n28148), .Z(n28145) );
  NOR U28531 ( .A(n28149), .B(n28145), .Z(n28151) );
  XOR U28532 ( .A(n28147), .B(n28146), .Z(n31823) );
  XOR U28533 ( .A(n28149), .B(n28148), .Z(n31822) );
  NOR U28534 ( .A(n31823), .B(n31822), .Z(n28150) );
  NOR U28535 ( .A(n28151), .B(n28150), .Z(n28154) );
  NOR U28536 ( .A(n100), .B(n169), .Z(n28153) );
  IV U28537 ( .A(n28153), .Z(n28152) );
  NOR U28538 ( .A(n28154), .B(n28152), .Z(n28159) );
  XOR U28539 ( .A(n28154), .B(n28153), .Z(n31825) );
  IV U28540 ( .A(n28155), .Z(n28157) );
  XOR U28541 ( .A(n28157), .B(n28156), .Z(n31824) );
  NOR U28542 ( .A(n31825), .B(n31824), .Z(n28158) );
  NOR U28543 ( .A(n28159), .B(n28158), .Z(n28164) );
  NOR U28544 ( .A(n101), .B(n169), .Z(n28163) );
  IV U28545 ( .A(n28163), .Z(n28160) );
  NOR U28546 ( .A(n28164), .B(n28160), .Z(n28166) );
  XOR U28547 ( .A(n28162), .B(n28161), .Z(n31827) );
  XOR U28548 ( .A(n28164), .B(n28163), .Z(n31826) );
  NOR U28549 ( .A(n31827), .B(n31826), .Z(n28165) );
  NOR U28550 ( .A(n28166), .B(n28165), .Z(n28168) );
  NOR U28551 ( .A(n102), .B(n169), .Z(n28169) );
  IV U28552 ( .A(n28169), .Z(n28167) );
  NOR U28553 ( .A(n28168), .B(n28167), .Z(n28173) );
  XOR U28554 ( .A(n28169), .B(n28168), .Z(n31829) );
  XOR U28555 ( .A(n28171), .B(n28170), .Z(n31828) );
  NOR U28556 ( .A(n31829), .B(n31828), .Z(n28172) );
  NOR U28557 ( .A(n28173), .B(n28172), .Z(n31700) );
  XOR U28558 ( .A(n28175), .B(n28174), .Z(n31699) );
  NOR U28559 ( .A(n31700), .B(n31699), .Z(n28176) );
  NOR U28560 ( .A(n28177), .B(n28176), .Z(n28180) );
  NOR U28561 ( .A(n103), .B(n169), .Z(n28179) );
  IV U28562 ( .A(n28179), .Z(n28178) );
  NOR U28563 ( .A(n28180), .B(n28178), .Z(n28185) );
  XOR U28564 ( .A(n28180), .B(n28179), .Z(n31702) );
  IV U28565 ( .A(n28181), .Z(n28183) );
  XOR U28566 ( .A(n28183), .B(n28182), .Z(n31701) );
  NOR U28567 ( .A(n31702), .B(n31701), .Z(n28184) );
  NOR U28568 ( .A(n28185), .B(n28184), .Z(n31704) );
  XOR U28569 ( .A(n28187), .B(n28186), .Z(n31703) );
  NOR U28570 ( .A(n31704), .B(n31703), .Z(n28188) );
  NOR U28571 ( .A(n28189), .B(n28188), .Z(n28192) );
  NOR U28572 ( .A(n104), .B(n169), .Z(n28191) );
  IV U28573 ( .A(n28191), .Z(n28190) );
  NOR U28574 ( .A(n28192), .B(n28190), .Z(n28197) );
  XOR U28575 ( .A(n28192), .B(n28191), .Z(n31706) );
  IV U28576 ( .A(n28193), .Z(n28195) );
  XOR U28577 ( .A(n28195), .B(n28194), .Z(n31705) );
  NOR U28578 ( .A(n31706), .B(n31705), .Z(n28196) );
  NOR U28579 ( .A(n28197), .B(n28196), .Z(n28200) );
  NOR U28580 ( .A(n105), .B(n169), .Z(n28199) );
  IV U28581 ( .A(n28199), .Z(n28198) );
  NOR U28582 ( .A(n28200), .B(n28198), .Z(n28204) );
  XOR U28583 ( .A(n28200), .B(n28199), .Z(n31708) );
  XOR U28584 ( .A(n28202), .B(n28201), .Z(n31707) );
  NOR U28585 ( .A(n31708), .B(n31707), .Z(n28203) );
  NOR U28586 ( .A(n28204), .B(n28203), .Z(n28210) );
  NOR U28587 ( .A(n106), .B(n169), .Z(n28209) );
  IV U28588 ( .A(n28209), .Z(n28205) );
  NOR U28589 ( .A(n28210), .B(n28205), .Z(n28212) );
  IV U28590 ( .A(n28206), .Z(n28208) );
  XOR U28591 ( .A(n28208), .B(n28207), .Z(n31710) );
  XOR U28592 ( .A(n28210), .B(n28209), .Z(n31709) );
  NOR U28593 ( .A(n31710), .B(n31709), .Z(n28211) );
  NOR U28594 ( .A(n28212), .B(n28211), .Z(n31712) );
  XOR U28595 ( .A(n28214), .B(n28213), .Z(n31711) );
  NOR U28596 ( .A(n31712), .B(n31711), .Z(n28215) );
  NOR U28597 ( .A(n28216), .B(n28215), .Z(n28219) );
  NOR U28598 ( .A(n107), .B(n169), .Z(n28218) );
  IV U28599 ( .A(n28218), .Z(n28217) );
  NOR U28600 ( .A(n28219), .B(n28217), .Z(n28224) );
  XOR U28601 ( .A(n28219), .B(n28218), .Z(n31714) );
  IV U28602 ( .A(n28220), .Z(n28222) );
  XOR U28603 ( .A(n28222), .B(n28221), .Z(n31713) );
  NOR U28604 ( .A(n31714), .B(n31713), .Z(n28223) );
  NOR U28605 ( .A(n28224), .B(n28223), .Z(n31716) );
  XOR U28606 ( .A(n28226), .B(n28225), .Z(n31715) );
  NOR U28607 ( .A(n31716), .B(n31715), .Z(n28227) );
  NOR U28608 ( .A(n28228), .B(n28227), .Z(n28231) );
  NOR U28609 ( .A(n108), .B(n169), .Z(n28230) );
  IV U28610 ( .A(n28230), .Z(n28229) );
  NOR U28611 ( .A(n28231), .B(n28229), .Z(n28236) );
  XOR U28612 ( .A(n28231), .B(n28230), .Z(n31718) );
  IV U28613 ( .A(n28232), .Z(n28234) );
  XOR U28614 ( .A(n28234), .B(n28233), .Z(n31717) );
  NOR U28615 ( .A(n31718), .B(n31717), .Z(n28235) );
  NOR U28616 ( .A(n28236), .B(n28235), .Z(n28239) );
  NOR U28617 ( .A(n109), .B(n169), .Z(n28238) );
  IV U28618 ( .A(n28238), .Z(n28237) );
  NOR U28619 ( .A(n28239), .B(n28237), .Z(n28243) );
  XOR U28620 ( .A(n28239), .B(n28238), .Z(n31722) );
  XOR U28621 ( .A(n28241), .B(n28240), .Z(n31721) );
  NOR U28622 ( .A(n31722), .B(n31721), .Z(n28242) );
  NOR U28623 ( .A(n28243), .B(n28242), .Z(n28249) );
  NOR U28624 ( .A(n110), .B(n169), .Z(n28248) );
  IV U28625 ( .A(n28248), .Z(n28244) );
  NOR U28626 ( .A(n28249), .B(n28244), .Z(n28251) );
  IV U28627 ( .A(n28245), .Z(n28247) );
  XOR U28628 ( .A(n28247), .B(n28246), .Z(n31724) );
  XOR U28629 ( .A(n28249), .B(n28248), .Z(n31723) );
  NOR U28630 ( .A(n31724), .B(n31723), .Z(n28250) );
  NOR U28631 ( .A(n28251), .B(n28250), .Z(n31726) );
  XOR U28632 ( .A(n28253), .B(n28252), .Z(n31725) );
  NOR U28633 ( .A(n31726), .B(n31725), .Z(n28254) );
  NOR U28634 ( .A(n28255), .B(n28254), .Z(n28258) );
  NOR U28635 ( .A(n111), .B(n169), .Z(n28257) );
  IV U28636 ( .A(n28257), .Z(n28256) );
  NOR U28637 ( .A(n28258), .B(n28256), .Z(n28263) );
  XOR U28638 ( .A(n28258), .B(n28257), .Z(n31728) );
  IV U28639 ( .A(n28259), .Z(n28261) );
  XOR U28640 ( .A(n28261), .B(n28260), .Z(n31727) );
  NOR U28641 ( .A(n31728), .B(n31727), .Z(n28262) );
  NOR U28642 ( .A(n28263), .B(n28262), .Z(n31730) );
  XOR U28643 ( .A(n28265), .B(n28264), .Z(n31729) );
  NOR U28644 ( .A(n31730), .B(n31729), .Z(n28266) );
  NOR U28645 ( .A(n28267), .B(n28266), .Z(n28270) );
  NOR U28646 ( .A(n112), .B(n169), .Z(n28269) );
  IV U28647 ( .A(n28269), .Z(n28268) );
  NOR U28648 ( .A(n28270), .B(n28268), .Z(n28275) );
  XOR U28649 ( .A(n28270), .B(n28269), .Z(n31732) );
  IV U28650 ( .A(n28271), .Z(n28273) );
  XOR U28651 ( .A(n28273), .B(n28272), .Z(n31731) );
  NOR U28652 ( .A(n31732), .B(n31731), .Z(n28274) );
  NOR U28653 ( .A(n28275), .B(n28274), .Z(n31734) );
  XOR U28654 ( .A(n28277), .B(n28276), .Z(n31733) );
  NOR U28655 ( .A(n31734), .B(n31733), .Z(n28278) );
  NOR U28656 ( .A(n28279), .B(n28278), .Z(n28282) );
  NOR U28657 ( .A(n113), .B(n169), .Z(n28281) );
  IV U28658 ( .A(n28281), .Z(n28280) );
  NOR U28659 ( .A(n28282), .B(n28280), .Z(n28287) );
  XOR U28660 ( .A(n28282), .B(n28281), .Z(n31736) );
  IV U28661 ( .A(n28283), .Z(n28285) );
  XOR U28662 ( .A(n28285), .B(n28284), .Z(n31735) );
  NOR U28663 ( .A(n31736), .B(n31735), .Z(n28286) );
  NOR U28664 ( .A(n28287), .B(n28286), .Z(n31738) );
  XOR U28665 ( .A(n28289), .B(n28288), .Z(n31737) );
  NOR U28666 ( .A(n31738), .B(n31737), .Z(n28290) );
  NOR U28667 ( .A(n28291), .B(n28290), .Z(n28294) );
  NOR U28668 ( .A(n114), .B(n169), .Z(n28293) );
  IV U28669 ( .A(n28293), .Z(n28292) );
  NOR U28670 ( .A(n28294), .B(n28292), .Z(n28299) );
  XOR U28671 ( .A(n28294), .B(n28293), .Z(n31740) );
  IV U28672 ( .A(n28295), .Z(n28297) );
  XOR U28673 ( .A(n28297), .B(n28296), .Z(n31739) );
  NOR U28674 ( .A(n31740), .B(n31739), .Z(n28298) );
  NOR U28675 ( .A(n28299), .B(n28298), .Z(n31744) );
  XOR U28676 ( .A(n28301), .B(n28300), .Z(n31743) );
  NOR U28677 ( .A(n31744), .B(n31743), .Z(n28302) );
  NOR U28678 ( .A(n28303), .B(n28302), .Z(n28306) );
  NOR U28679 ( .A(n115), .B(n169), .Z(n28305) );
  IV U28680 ( .A(n28305), .Z(n28304) );
  NOR U28681 ( .A(n28306), .B(n28304), .Z(n28311) );
  XOR U28682 ( .A(n28306), .B(n28305), .Z(n31746) );
  IV U28683 ( .A(n28307), .Z(n28309) );
  XOR U28684 ( .A(n28309), .B(n28308), .Z(n31745) );
  NOR U28685 ( .A(n31746), .B(n31745), .Z(n28310) );
  NOR U28686 ( .A(n28311), .B(n28310), .Z(n31748) );
  XOR U28687 ( .A(n28313), .B(n28312), .Z(n31747) );
  NOR U28688 ( .A(n31748), .B(n31747), .Z(n28314) );
  NOR U28689 ( .A(n28315), .B(n28314), .Z(n28318) );
  NOR U28690 ( .A(n116), .B(n169), .Z(n28317) );
  IV U28691 ( .A(n28317), .Z(n28316) );
  NOR U28692 ( .A(n28318), .B(n28316), .Z(n28323) );
  XOR U28693 ( .A(n28318), .B(n28317), .Z(n31750) );
  IV U28694 ( .A(n28319), .Z(n28321) );
  XOR U28695 ( .A(n28321), .B(n28320), .Z(n31749) );
  NOR U28696 ( .A(n31750), .B(n31749), .Z(n28322) );
  NOR U28697 ( .A(n28323), .B(n28322), .Z(n31752) );
  XOR U28698 ( .A(n28325), .B(n28324), .Z(n31751) );
  NOR U28699 ( .A(n31752), .B(n31751), .Z(n28326) );
  NOR U28700 ( .A(n28327), .B(n28326), .Z(n28330) );
  NOR U28701 ( .A(n117), .B(n169), .Z(n28329) );
  IV U28702 ( .A(n28329), .Z(n28328) );
  NOR U28703 ( .A(n28330), .B(n28328), .Z(n28335) );
  XOR U28704 ( .A(n28330), .B(n28329), .Z(n31754) );
  IV U28705 ( .A(n28331), .Z(n28333) );
  XOR U28706 ( .A(n28333), .B(n28332), .Z(n31753) );
  NOR U28707 ( .A(n31754), .B(n31753), .Z(n28334) );
  NOR U28708 ( .A(n28335), .B(n28334), .Z(n31756) );
  XOR U28709 ( .A(n28337), .B(n28336), .Z(n31755) );
  NOR U28710 ( .A(n31756), .B(n31755), .Z(n28338) );
  NOR U28711 ( .A(n28339), .B(n28338), .Z(n28342) );
  NOR U28712 ( .A(n119), .B(n169), .Z(n28341) );
  IV U28713 ( .A(n28341), .Z(n28340) );
  NOR U28714 ( .A(n28342), .B(n28340), .Z(n28347) );
  XOR U28715 ( .A(n28342), .B(n28341), .Z(n31758) );
  IV U28716 ( .A(n28343), .Z(n28345) );
  XOR U28717 ( .A(n28345), .B(n28344), .Z(n31757) );
  NOR U28718 ( .A(n31758), .B(n31757), .Z(n28346) );
  NOR U28719 ( .A(n28347), .B(n28346), .Z(n31760) );
  XOR U28720 ( .A(n28349), .B(n28348), .Z(n31759) );
  NOR U28721 ( .A(n31760), .B(n31759), .Z(n28350) );
  NOR U28722 ( .A(n28351), .B(n28350), .Z(n28354) );
  NOR U28723 ( .A(n123), .B(n169), .Z(n28353) );
  IV U28724 ( .A(n28353), .Z(n28352) );
  NOR U28725 ( .A(n28354), .B(n28352), .Z(n28359) );
  XOR U28726 ( .A(n28354), .B(n28353), .Z(n31762) );
  IV U28727 ( .A(n28355), .Z(n28357) );
  XOR U28728 ( .A(n28357), .B(n28356), .Z(n31761) );
  NOR U28729 ( .A(n31762), .B(n31761), .Z(n28358) );
  NOR U28730 ( .A(n28359), .B(n28358), .Z(n31766) );
  XOR U28731 ( .A(n28361), .B(n28360), .Z(n31765) );
  NOR U28732 ( .A(n31766), .B(n31765), .Z(n28362) );
  NOR U28733 ( .A(n28363), .B(n28362), .Z(n28368) );
  NOR U28734 ( .A(n126), .B(n169), .Z(n28367) );
  IV U28735 ( .A(n28367), .Z(n28364) );
  NOR U28736 ( .A(n28368), .B(n28364), .Z(n28370) );
  XOR U28737 ( .A(n28366), .B(n28365), .Z(n31768) );
  XOR U28738 ( .A(n28368), .B(n28367), .Z(n31767) );
  NOR U28739 ( .A(n31768), .B(n31767), .Z(n28369) );
  NOR U28740 ( .A(n28370), .B(n28369), .Z(n31770) );
  IV U28741 ( .A(n31770), .Z(n28374) );
  IV U28742 ( .A(n28371), .Z(n28373) );
  XOR U28743 ( .A(n28373), .B(n28372), .Z(n31769) );
  NOR U28744 ( .A(n28374), .B(n31769), .Z(n28375) );
  NOR U28745 ( .A(n28376), .B(n28375), .Z(n28377) );
  IV U28746 ( .A(n28377), .Z(n31771) );
  NOR U28747 ( .A(n31772), .B(n31771), .Z(n28378) );
  NOR U28748 ( .A(n28379), .B(n28378), .Z(n28381) );
  IV U28749 ( .A(n28381), .Z(n28380) );
  NOR U28750 ( .A(n28382), .B(n28380), .Z(n28384) );
  NOR U28751 ( .A(n133), .B(n169), .Z(n31773) );
  XOR U28752 ( .A(n28382), .B(n28381), .Z(n31774) );
  NOR U28753 ( .A(n31773), .B(n31774), .Z(n28383) );
  NOR U28754 ( .A(n28384), .B(n28383), .Z(n28385) );
  IV U28755 ( .A(n28385), .Z(n28388) );
  NOR U28756 ( .A(n135), .B(n169), .Z(n28387) );
  IV U28757 ( .A(n28387), .Z(n28386) );
  NOR U28758 ( .A(n28388), .B(n28386), .Z(n28393) );
  XOR U28759 ( .A(n28388), .B(n28387), .Z(n31777) );
  IV U28760 ( .A(n28389), .Z(n28391) );
  XOR U28761 ( .A(n28391), .B(n28390), .Z(n31776) );
  NOR U28762 ( .A(n31777), .B(n31776), .Z(n28392) );
  NOR U28763 ( .A(n28393), .B(n28392), .Z(n31779) );
  XOR U28764 ( .A(n28395), .B(n28394), .Z(n31778) );
  NOR U28765 ( .A(n31779), .B(n31778), .Z(n28396) );
  NOR U28766 ( .A(n28397), .B(n28396), .Z(n28402) );
  NOR U28767 ( .A(n139), .B(n169), .Z(n28401) );
  IV U28768 ( .A(n28401), .Z(n28398) );
  NOR U28769 ( .A(n28402), .B(n28398), .Z(n28404) );
  XOR U28770 ( .A(n28400), .B(n28399), .Z(n31781) );
  XOR U28771 ( .A(n28402), .B(n28401), .Z(n31780) );
  NOR U28772 ( .A(n31781), .B(n31780), .Z(n28403) );
  NOR U28773 ( .A(n28404), .B(n28403), .Z(n28407) );
  XOR U28774 ( .A(n28406), .B(n28405), .Z(n28408) );
  NOR U28775 ( .A(n28407), .B(n28408), .Z(n28412) );
  IV U28776 ( .A(n28407), .Z(n28409) );
  XOR U28777 ( .A(n28409), .B(n28408), .Z(n31783) );
  NOR U28778 ( .A(n141), .B(n169), .Z(n28410) );
  IV U28779 ( .A(n28410), .Z(n31782) );
  NOR U28780 ( .A(n31783), .B(n31782), .Z(n28411) );
  NOR U28781 ( .A(n28412), .B(n28411), .Z(n31785) );
  XOR U28782 ( .A(n28414), .B(n28413), .Z(n31784) );
  NOR U28783 ( .A(n31785), .B(n31784), .Z(n28415) );
  NOR U28784 ( .A(n28416), .B(n28415), .Z(n28419) );
  XOR U28785 ( .A(n28418), .B(n28417), .Z(n28420) );
  NOR U28786 ( .A(n28419), .B(n28420), .Z(n28424) );
  IV U28787 ( .A(n28419), .Z(n28421) );
  XOR U28788 ( .A(n28421), .B(n28420), .Z(n31789) );
  NOR U28789 ( .A(n145), .B(n169), .Z(n28422) );
  IV U28790 ( .A(n28422), .Z(n31788) );
  NOR U28791 ( .A(n31789), .B(n31788), .Z(n28423) );
  NOR U28792 ( .A(n28424), .B(n28423), .Z(n28427) );
  NOR U28793 ( .A(n147), .B(n169), .Z(n28426) );
  IV U28794 ( .A(n28426), .Z(n28425) );
  NOR U28795 ( .A(n28427), .B(n28425), .Z(n28432) );
  XOR U28796 ( .A(n28427), .B(n28426), .Z(n31791) );
  IV U28797 ( .A(n28428), .Z(n28430) );
  XOR U28798 ( .A(n28430), .B(n28429), .Z(n31790) );
  NOR U28799 ( .A(n31791), .B(n31790), .Z(n28431) );
  NOR U28800 ( .A(n28432), .B(n28431), .Z(n28433) );
  IV U28801 ( .A(n28433), .Z(n31793) );
  XOR U28802 ( .A(n28435), .B(n28434), .Z(n31792) );
  IV U28803 ( .A(n31792), .Z(n28436) );
  NOR U28804 ( .A(n31793), .B(n28436), .Z(n28437) );
  NOR U28805 ( .A(n28438), .B(n28437), .Z(n28439) );
  IV U28806 ( .A(n28439), .Z(n28442) );
  NOR U28807 ( .A(n150), .B(n169), .Z(n28441) );
  IV U28808 ( .A(n28441), .Z(n28440) );
  NOR U28809 ( .A(n28442), .B(n28440), .Z(n28447) );
  XOR U28810 ( .A(n28442), .B(n28441), .Z(n31795) );
  IV U28811 ( .A(n28443), .Z(n28445) );
  XOR U28812 ( .A(n28445), .B(n28444), .Z(n31794) );
  NOR U28813 ( .A(n31795), .B(n31794), .Z(n28446) );
  NOR U28814 ( .A(n28447), .B(n28446), .Z(n31797) );
  XOR U28815 ( .A(n28449), .B(n28448), .Z(n31796) );
  NOR U28816 ( .A(n31797), .B(n31796), .Z(n28450) );
  NOR U28817 ( .A(n28451), .B(n28450), .Z(n28453) );
  IV U28818 ( .A(n28453), .Z(n31801) );
  NOR U28819 ( .A(n31799), .B(n31801), .Z(n28458) );
  IV U28820 ( .A(n31799), .Z(n28452) );
  NOR U28821 ( .A(n28453), .B(n28452), .Z(n28456) );
  XOR U28822 ( .A(n28455), .B(n28454), .Z(n31798) );
  NOR U28823 ( .A(n28456), .B(n31798), .Z(n28457) );
  NOR U28824 ( .A(n28458), .B(n28457), .Z(n28463) );
  IV U28825 ( .A(n28463), .Z(n28461) );
  XOR U28826 ( .A(n28460), .B(n28459), .Z(n28462) );
  NOR U28827 ( .A(n28461), .B(n28462), .Z(n28466) );
  XOR U28828 ( .A(n28463), .B(n28462), .Z(n31803) );
  NOR U28829 ( .A(n156), .B(n169), .Z(n28464) );
  IV U28830 ( .A(n28464), .Z(n31802) );
  NOR U28831 ( .A(n31803), .B(n31802), .Z(n28465) );
  NOR U28832 ( .A(n28466), .B(n28465), .Z(n28467) );
  NOR U28833 ( .A(n158), .B(n169), .Z(n28468) );
  IV U28834 ( .A(n28468), .Z(n31804) );
  NOR U28835 ( .A(n28467), .B(n31804), .Z(n28474) );
  IV U28836 ( .A(n28467), .Z(n31805) );
  NOR U28837 ( .A(n28468), .B(n31805), .Z(n28472) );
  IV U28838 ( .A(n28469), .Z(n28471) );
  XOR U28839 ( .A(n28471), .B(n28470), .Z(n31807) );
  NOR U28840 ( .A(n28472), .B(n31807), .Z(n28473) );
  NOR U28841 ( .A(n28474), .B(n28473), .Z(n28475) );
  IV U28842 ( .A(n28475), .Z(n31809) );
  XOR U28843 ( .A(n28477), .B(n28476), .Z(n31808) );
  IV U28844 ( .A(n31808), .Z(n28478) );
  NOR U28845 ( .A(n31809), .B(n28478), .Z(n28479) );
  NOR U28846 ( .A(n28480), .B(n28479), .Z(n28481) );
  IV U28847 ( .A(n28481), .Z(n31810) );
  NOR U28848 ( .A(n31811), .B(n31810), .Z(n28482) );
  NOR U28849 ( .A(n28483), .B(n28482), .Z(n31814) );
  NOR U28850 ( .A(n28484), .B(n31814), .Z(n28485) );
  NOR U28851 ( .A(n28486), .B(n28485), .Z(n28492) );
  NOR U28852 ( .A(n167), .B(n169), .Z(n28491) );
  IV U28853 ( .A(n28491), .Z(n28487) );
  NOR U28854 ( .A(n28492), .B(n28487), .Z(n28494) );
  XOR U28855 ( .A(n28489), .B(n28488), .Z(n28490) );
  IV U28856 ( .A(n28490), .Z(n31819) );
  XOR U28857 ( .A(n28492), .B(n28491), .Z(n31818) );
  NOR U28858 ( .A(n31819), .B(n31818), .Z(n28493) );
  NOR U28859 ( .A(n28494), .B(n28493), .Z(n31821) );
  XOR U28860 ( .A(n28496), .B(n28495), .Z(n28497) );
  XOR U28861 ( .A(n28498), .B(n28497), .Z(n31820) );
  NOR U28862 ( .A(n31821), .B(n31820), .Z(n28499) );
  IV U28863 ( .A(n28499), .Z(n31462) );
  XOR U28864 ( .A(n28501), .B(n28500), .Z(n31461) );
  NOR U28865 ( .A(n31462), .B(n31461), .Z(n31463) );
  NOR U28866 ( .A(n28503), .B(n31488), .Z(n28507) );
  IV U28867 ( .A(n28504), .Z(n31483) );
  NOR U28868 ( .A(n28505), .B(n31483), .Z(n28506) );
  NOR U28869 ( .A(n28507), .B(n28506), .Z(n28508) );
  IV U28870 ( .A(n28508), .Z(n28509) );
  NOR U28871 ( .A(n31486), .B(n28509), .Z(n28510) );
  NOR U28872 ( .A(n28511), .B(n28510), .Z(n28517) );
  NOR U28873 ( .A(n31504), .B(n28512), .Z(n28514) );
  NOR U28874 ( .A(n31501), .B(n31503), .Z(n28513) );
  NOR U28875 ( .A(n28514), .B(n28513), .Z(n28515) );
  IV U28876 ( .A(n28515), .Z(n28516) );
  NOR U28877 ( .A(n28517), .B(n28516), .Z(n28518) );
  NOR U28878 ( .A(n28519), .B(n28518), .Z(n31517) );
  XOR U28879 ( .A(n28521), .B(n28520), .Z(n31524) );
  IV U28880 ( .A(n31524), .Z(n28522) );
  NOR U28881 ( .A(n31523), .B(n28522), .Z(n28523) );
  NOR U28882 ( .A(n31517), .B(n28523), .Z(n28524) );
  IV U28883 ( .A(n28524), .Z(n28525) );
  NOR U28884 ( .A(n28526), .B(n28525), .Z(n28527) );
  IV U28885 ( .A(n28527), .Z(n28528) );
  NOR U28886 ( .A(n28529), .B(n28528), .Z(n28530) );
  NOR U28887 ( .A(n28531), .B(n28530), .Z(n28532) );
  NOR U28888 ( .A(n28533), .B(n28532), .Z(n28534) );
  NOR U28889 ( .A(n28535), .B(n28534), .Z(n31541) );
  IV U28890 ( .A(n31541), .Z(n28536) );
  NOR U28891 ( .A(n31542), .B(n28536), .Z(n28537) );
  NOR U28892 ( .A(n28538), .B(n28537), .Z(n31544) );
  XOR U28893 ( .A(n28540), .B(n28539), .Z(n31543) );
  IV U28894 ( .A(n31543), .Z(n28541) );
  NOR U28895 ( .A(n31544), .B(n28541), .Z(n28542) );
  NOR U28896 ( .A(n28543), .B(n28542), .Z(n31545) );
  IV U28897 ( .A(n28544), .Z(n31549) );
  XOR U28898 ( .A(n31549), .B(n28545), .Z(n31546) );
  NOR U28899 ( .A(n31545), .B(n31546), .Z(n28546) );
  NOR U28900 ( .A(n28547), .B(n28546), .Z(n28548) );
  IV U28901 ( .A(n28548), .Z(n31547) );
  NOR U28902 ( .A(n28549), .B(n31547), .Z(n28551) );
  IV U28903 ( .A(n31548), .Z(n31552) );
  NOR U28904 ( .A(n31552), .B(n31555), .Z(n28550) );
  NOR U28905 ( .A(n28551), .B(n28550), .Z(n31560) );
  NOR U28906 ( .A(n28552), .B(n31560), .Z(n31562) );
  IV U28907 ( .A(n31562), .Z(n31572) );
  NOR U28908 ( .A(n28553), .B(n31572), .Z(n28554) );
  NOR U28909 ( .A(n28555), .B(n28554), .Z(n28561) );
  NOR U28910 ( .A(n31578), .B(n28556), .Z(n28558) );
  NOR U28911 ( .A(n31570), .B(n31577), .Z(n28557) );
  NOR U28912 ( .A(n28558), .B(n28557), .Z(n28559) );
  IV U28913 ( .A(n28559), .Z(n28560) );
  NOR U28914 ( .A(n28561), .B(n28560), .Z(n28562) );
  NOR U28915 ( .A(n28563), .B(n28562), .Z(n31591) );
  NOR U28916 ( .A(n28565), .B(n28564), .Z(n31595) );
  IV U28917 ( .A(n28566), .Z(n28574) );
  XOR U28918 ( .A(n28574), .B(n28575), .Z(n31594) );
  NOR U28919 ( .A(n31595), .B(n31594), .Z(n31601) );
  NOR U28920 ( .A(n31591), .B(n31601), .Z(n28567) );
  IV U28921 ( .A(n28567), .Z(n28568) );
  NOR U28922 ( .A(n28569), .B(n28568), .Z(n28581) );
  NOR U28923 ( .A(n31617), .B(n28581), .Z(n28586) );
  IV U28924 ( .A(n28570), .Z(n31589) );
  IV U28925 ( .A(n31588), .Z(n28571) );
  NOR U28926 ( .A(n31589), .B(n28571), .Z(n31593) );
  NOR U28927 ( .A(n31595), .B(n31593), .Z(n28572) );
  IV U28928 ( .A(n28572), .Z(n28573) );
  NOR U28929 ( .A(n31610), .B(n28573), .Z(n28579) );
  NOR U28930 ( .A(n28575), .B(n28574), .Z(n28576) );
  NOR U28931 ( .A(n31606), .B(n28576), .Z(n28577) );
  IV U28932 ( .A(n28577), .Z(n28578) );
  NOR U28933 ( .A(n28579), .B(n28578), .Z(n28580) );
  NOR U28934 ( .A(n28581), .B(n28580), .Z(n28583) );
  IV U28935 ( .A(n31617), .Z(n28582) );
  NOR U28936 ( .A(n28583), .B(n28582), .Z(n28584) );
  NOR U28937 ( .A(n31611), .B(n28584), .Z(n28585) );
  NOR U28938 ( .A(n28586), .B(n28585), .Z(n31618) );
  IV U28939 ( .A(n31618), .Z(n31628) );
  NOR U28940 ( .A(n28588), .B(n28587), .Z(n31621) );
  XOR U28941 ( .A(n28590), .B(n28589), .Z(n28595) );
  NOR U28942 ( .A(n31621), .B(n28595), .Z(n28591) );
  NOR U28943 ( .A(n31628), .B(n28591), .Z(n28592) );
  IV U28944 ( .A(n28592), .Z(n28593) );
  NOR U28945 ( .A(n28594), .B(n28593), .Z(n28600) );
  IV U28946 ( .A(n31621), .Z(n31631) );
  IV U28947 ( .A(n28595), .Z(n31622) );
  NOR U28948 ( .A(n31631), .B(n31622), .Z(n28596) );
  NOR U28949 ( .A(n31626), .B(n28596), .Z(n28598) );
  IV U28950 ( .A(n28597), .Z(n31633) );
  NOR U28951 ( .A(n28598), .B(n31633), .Z(n28599) );
  NOR U28952 ( .A(n28600), .B(n28599), .Z(n28607) );
  NOR U28953 ( .A(n31643), .B(n28601), .Z(n28604) );
  NOR U28954 ( .A(n28602), .B(n31636), .Z(n28603) );
  NOR U28955 ( .A(n28604), .B(n28603), .Z(n28605) );
  IV U28956 ( .A(n28605), .Z(n28606) );
  NOR U28957 ( .A(n28607), .B(n28606), .Z(n28608) );
  NOR U28958 ( .A(n28609), .B(n28608), .Z(n31650) );
  IV U28959 ( .A(n31650), .Z(n28610) );
  NOR U28960 ( .A(n31646), .B(n28610), .Z(n28611) );
  NOR U28961 ( .A(n28612), .B(n28611), .Z(n28613) );
  IV U28962 ( .A(n28613), .Z(n31647) );
  NOR U28963 ( .A(n28614), .B(n31647), .Z(n28616) );
  IV U28964 ( .A(n31648), .Z(n31652) );
  NOR U28965 ( .A(n31652), .B(n31655), .Z(n28615) );
  NOR U28966 ( .A(n28616), .B(n28615), .Z(n28617) );
  IV U28967 ( .A(n28617), .Z(n31658) );
  XOR U28968 ( .A(n28619), .B(n28618), .Z(n31657) );
  IV U28969 ( .A(n31657), .Z(n28620) );
  NOR U28970 ( .A(n31658), .B(n28620), .Z(n28621) );
  NOR U28971 ( .A(n28622), .B(n28621), .Z(n31660) );
  XOR U28972 ( .A(n28624), .B(n28623), .Z(n31659) );
  IV U28973 ( .A(n31659), .Z(n28625) );
  NOR U28974 ( .A(n31660), .B(n28625), .Z(n28626) );
  NOR U28975 ( .A(n28627), .B(n28626), .Z(n31663) );
  IV U28976 ( .A(n31663), .Z(n31665) );
  NOR U28977 ( .A(n28628), .B(n31665), .Z(n31672) );
  IV U28978 ( .A(n31672), .Z(n28629) );
  NOR U28979 ( .A(n28630), .B(n28629), .Z(n28636) );
  NOR U28980 ( .A(n28632), .B(n28631), .Z(n28641) );
  IV U28981 ( .A(n28641), .Z(n31680) );
  XOR U28982 ( .A(n28634), .B(n28633), .Z(n31679) );
  IV U28983 ( .A(n31679), .Z(n28635) );
  NOR U28984 ( .A(n31680), .B(n28635), .Z(n31684) );
  NOR U28985 ( .A(n28636), .B(n31684), .Z(n28637) );
  IV U28986 ( .A(n28637), .Z(n28638) );
  NOR U28987 ( .A(n28639), .B(n28638), .Z(n28646) );
  NOR U28988 ( .A(n31686), .B(n28640), .Z(n28643) );
  NOR U28989 ( .A(n28641), .B(n31679), .Z(n28642) );
  NOR U28990 ( .A(n28643), .B(n28642), .Z(n28644) );
  IV U28991 ( .A(n28644), .Z(n28645) );
  NOR U28992 ( .A(n28646), .B(n28645), .Z(n28647) );
  NOR U28993 ( .A(n28648), .B(n28647), .Z(n29409) );
  NOR U28994 ( .A(n28650), .B(n28649), .Z(n29022) );
  IV U28995 ( .A(n29022), .Z(n29394) );
  IV U28996 ( .A(n28651), .Z(n28652) );
  NOR U28997 ( .A(n28653), .B(n28652), .Z(n28658) );
  IV U28998 ( .A(n28654), .Z(n28655) );
  NOR U28999 ( .A(n28656), .B(n28655), .Z(n28657) );
  NOR U29000 ( .A(n28658), .B(n28657), .Z(n29028) );
  NOR U29001 ( .A(n167), .B(n118), .Z(n28838) );
  IV U29002 ( .A(n28659), .Z(n28660) );
  NOR U29003 ( .A(n28661), .B(n28660), .Z(n28665) );
  NOR U29004 ( .A(n28663), .B(n28662), .Z(n28664) );
  NOR U29005 ( .A(n28665), .B(n28664), .Z(n28837) );
  NOR U29006 ( .A(n163), .B(n122), .Z(n29016) );
  IV U29007 ( .A(n28666), .Z(n28667) );
  NOR U29008 ( .A(n28668), .B(n28667), .Z(n28673) );
  IV U29009 ( .A(n28669), .Z(n28670) );
  NOR U29010 ( .A(n28671), .B(n28670), .Z(n28672) );
  NOR U29011 ( .A(n28673), .B(n28672), .Z(n29015) );
  NOR U29012 ( .A(n158), .B(n127), .Z(n28854) );
  IV U29013 ( .A(n28674), .Z(n28675) );
  NOR U29014 ( .A(n28676), .B(n28675), .Z(n28681) );
  IV U29015 ( .A(n28677), .Z(n28678) );
  NOR U29016 ( .A(n28679), .B(n28678), .Z(n28680) );
  NOR U29017 ( .A(n28681), .B(n28680), .Z(n28853) );
  NOR U29018 ( .A(n155), .B(n130), .Z(n29001) );
  IV U29019 ( .A(n28682), .Z(n28683) );
  NOR U29020 ( .A(n28684), .B(n28683), .Z(n28689) );
  IV U29021 ( .A(n28685), .Z(n28686) );
  NOR U29022 ( .A(n28687), .B(n28686), .Z(n28688) );
  NOR U29023 ( .A(n28689), .B(n28688), .Z(n29000) );
  NOR U29024 ( .A(n150), .B(n134), .Z(n28986) );
  IV U29025 ( .A(n28690), .Z(n28691) );
  NOR U29026 ( .A(n28692), .B(n28691), .Z(n28697) );
  IV U29027 ( .A(n28693), .Z(n28694) );
  NOR U29028 ( .A(n28695), .B(n28694), .Z(n28696) );
  NOR U29029 ( .A(n28697), .B(n28696), .Z(n28985) );
  NOR U29030 ( .A(n147), .B(n138), .Z(n28978) );
  IV U29031 ( .A(n28698), .Z(n28699) );
  NOR U29032 ( .A(n28700), .B(n28699), .Z(n28705) );
  IV U29033 ( .A(n28701), .Z(n28702) );
  NOR U29034 ( .A(n28703), .B(n28702), .Z(n28704) );
  NOR U29035 ( .A(n28705), .B(n28704), .Z(n28977) );
  NOR U29036 ( .A(n143), .B(n142), .Z(n28877) );
  NOR U29037 ( .A(n28707), .B(n28706), .Z(n28711) );
  NOR U29038 ( .A(n28709), .B(n28708), .Z(n28710) );
  NOR U29039 ( .A(n28711), .B(n28710), .Z(n28882) );
  NOR U29040 ( .A(n141), .B(n144), .Z(n28712) );
  IV U29041 ( .A(n28712), .Z(n28883) );
  XOR U29042 ( .A(n28882), .B(n28883), .Z(n28886) );
  NOR U29043 ( .A(n139), .B(n146), .Z(n28963) );
  NOR U29044 ( .A(n28714), .B(n28713), .Z(n28719) );
  IV U29045 ( .A(n28715), .Z(n28716) );
  NOR U29046 ( .A(n28717), .B(n28716), .Z(n28718) );
  NOR U29047 ( .A(n28719), .B(n28718), .Z(n28960) );
  NOR U29048 ( .A(n135), .B(n151), .Z(n28893) );
  IV U29049 ( .A(n28720), .Z(n28721) );
  NOR U29050 ( .A(n28722), .B(n28721), .Z(n28727) );
  IV U29051 ( .A(n28723), .Z(n28724) );
  NOR U29052 ( .A(n28725), .B(n28724), .Z(n28726) );
  NOR U29053 ( .A(n28727), .B(n28726), .Z(n28892) );
  NOR U29054 ( .A(n131), .B(n154), .Z(n28909) );
  IV U29055 ( .A(n28728), .Z(n28729) );
  NOR U29056 ( .A(n28730), .B(n28729), .Z(n28735) );
  IV U29057 ( .A(n28731), .Z(n28733) );
  NOR U29058 ( .A(n28733), .B(n28732), .Z(n28734) );
  NOR U29059 ( .A(n28735), .B(n28734), .Z(n28908) );
  NOR U29060 ( .A(n126), .B(n159), .Z(n28940) );
  NOR U29061 ( .A(n28737), .B(n28736), .Z(n28741) );
  NOR U29062 ( .A(n28739), .B(n28738), .Z(n28740) );
  NOR U29063 ( .A(n28741), .B(n28740), .Z(n28937) );
  NOR U29064 ( .A(n123), .B(n162), .Z(n28932) );
  NOR U29065 ( .A(n28743), .B(n28742), .Z(n28747) );
  NOR U29066 ( .A(n28745), .B(n28744), .Z(n28746) );
  NOR U29067 ( .A(n28747), .B(n28746), .Z(n28929) );
  IV U29068 ( .A(n28748), .Z(n28921) );
  NOR U29069 ( .A(n28749), .B(n28921), .Z(n28753) );
  NOR U29070 ( .A(n28751), .B(n28750), .Z(n28752) );
  NOR U29071 ( .A(n28753), .B(n28752), .Z(n28925) );
  NOR U29072 ( .A(n164), .B(n120), .Z(n29116) );
  NOR U29073 ( .A(n166), .B(n119), .Z(n28754) );
  XOR U29074 ( .A(n29116), .B(n28754), .Z(n28923) );
  XOR U29075 ( .A(n28925), .B(n28923), .Z(n28931) );
  XOR U29076 ( .A(n28929), .B(n28931), .Z(n28934) );
  XOR U29077 ( .A(n28932), .B(n28934), .Z(n28917) );
  IV U29078 ( .A(n28755), .Z(n28756) );
  NOR U29079 ( .A(n28757), .B(n28756), .Z(n28761) );
  NOR U29080 ( .A(n28759), .B(n28758), .Z(n28760) );
  NOR U29081 ( .A(n28761), .B(n28760), .Z(n28916) );
  NOR U29082 ( .A(n125), .B(n160), .Z(n28914) );
  XOR U29083 ( .A(n28916), .B(n28914), .Z(n28918) );
  XOR U29084 ( .A(n28917), .B(n28918), .Z(n28762) );
  IV U29085 ( .A(n28762), .Z(n28938) );
  XOR U29086 ( .A(n28937), .B(n28938), .Z(n28942) );
  XOR U29087 ( .A(n28940), .B(n28942), .Z(n28949) );
  IV U29088 ( .A(n28763), .Z(n28764) );
  NOR U29089 ( .A(n28765), .B(n28764), .Z(n28769) );
  NOR U29090 ( .A(n28767), .B(n28766), .Z(n28768) );
  NOR U29091 ( .A(n28769), .B(n28768), .Z(n28947) );
  NOR U29092 ( .A(n128), .B(n157), .Z(n28945) );
  XOR U29093 ( .A(n28947), .B(n28945), .Z(n28948) );
  XOR U29094 ( .A(n28949), .B(n28948), .Z(n28906) );
  XOR U29095 ( .A(n28908), .B(n28906), .Z(n28911) );
  XOR U29096 ( .A(n28909), .B(n28911), .Z(n28902) );
  IV U29097 ( .A(n28770), .Z(n28771) );
  NOR U29098 ( .A(n28772), .B(n28771), .Z(n28776) );
  NOR U29099 ( .A(n28774), .B(n28773), .Z(n28775) );
  NOR U29100 ( .A(n28776), .B(n28775), .Z(n28900) );
  NOR U29101 ( .A(n133), .B(n152), .Z(n28898) );
  XOR U29102 ( .A(n28900), .B(n28898), .Z(n28901) );
  XOR U29103 ( .A(n28902), .B(n28901), .Z(n28890) );
  XOR U29104 ( .A(n28892), .B(n28890), .Z(n28895) );
  XOR U29105 ( .A(n28893), .B(n28895), .Z(n28956) );
  IV U29106 ( .A(n28777), .Z(n28778) );
  NOR U29107 ( .A(n28779), .B(n28778), .Z(n28783) );
  NOR U29108 ( .A(n28781), .B(n28780), .Z(n28782) );
  NOR U29109 ( .A(n28783), .B(n28782), .Z(n28955) );
  NOR U29110 ( .A(n137), .B(n149), .Z(n28953) );
  XOR U29111 ( .A(n28955), .B(n28953), .Z(n28957) );
  XOR U29112 ( .A(n28956), .B(n28957), .Z(n28784) );
  IV U29113 ( .A(n28784), .Z(n28961) );
  XOR U29114 ( .A(n28960), .B(n28961), .Z(n28965) );
  XOR U29115 ( .A(n28963), .B(n28965), .Z(n28885) );
  XOR U29116 ( .A(n28886), .B(n28885), .Z(n28875) );
  IV U29117 ( .A(n28785), .Z(n28786) );
  NOR U29118 ( .A(n28787), .B(n28786), .Z(n28792) );
  IV U29119 ( .A(n28788), .Z(n28789) );
  NOR U29120 ( .A(n28790), .B(n28789), .Z(n28791) );
  NOR U29121 ( .A(n28792), .B(n28791), .Z(n28873) );
  XOR U29122 ( .A(n28875), .B(n28873), .Z(n28876) );
  XOR U29123 ( .A(n28877), .B(n28876), .Z(n28972) );
  IV U29124 ( .A(n28793), .Z(n28794) );
  NOR U29125 ( .A(n28795), .B(n28794), .Z(n28799) );
  NOR U29126 ( .A(n28797), .B(n28796), .Z(n28798) );
  NOR U29127 ( .A(n28799), .B(n28798), .Z(n28970) );
  NOR U29128 ( .A(n145), .B(n140), .Z(n28968) );
  XOR U29129 ( .A(n28970), .B(n28968), .Z(n28971) );
  XOR U29130 ( .A(n28972), .B(n28971), .Z(n28975) );
  XOR U29131 ( .A(n28977), .B(n28975), .Z(n28980) );
  XOR U29132 ( .A(n28978), .B(n28980), .Z(n28870) );
  IV U29133 ( .A(n28800), .Z(n28801) );
  NOR U29134 ( .A(n28802), .B(n28801), .Z(n28806) );
  NOR U29135 ( .A(n28804), .B(n28803), .Z(n28805) );
  NOR U29136 ( .A(n28806), .B(n28805), .Z(n28868) );
  NOR U29137 ( .A(n148), .B(n136), .Z(n28866) );
  XOR U29138 ( .A(n28868), .B(n28866), .Z(n28869) );
  XOR U29139 ( .A(n28870), .B(n28869), .Z(n28983) );
  XOR U29140 ( .A(n28985), .B(n28983), .Z(n28988) );
  XOR U29141 ( .A(n28986), .B(n28988), .Z(n28995) );
  IV U29142 ( .A(n28807), .Z(n28808) );
  NOR U29143 ( .A(n28809), .B(n28808), .Z(n28813) );
  NOR U29144 ( .A(n28811), .B(n28810), .Z(n28812) );
  NOR U29145 ( .A(n28813), .B(n28812), .Z(n28993) );
  NOR U29146 ( .A(n153), .B(n132), .Z(n28991) );
  XOR U29147 ( .A(n28993), .B(n28991), .Z(n28994) );
  XOR U29148 ( .A(n28995), .B(n28994), .Z(n28998) );
  XOR U29149 ( .A(n29000), .B(n28998), .Z(n29003) );
  XOR U29150 ( .A(n29001), .B(n29003), .Z(n28862) );
  IV U29151 ( .A(n28814), .Z(n28815) );
  NOR U29152 ( .A(n28816), .B(n28815), .Z(n28820) );
  NOR U29153 ( .A(n28818), .B(n28817), .Z(n28819) );
  NOR U29154 ( .A(n28820), .B(n28819), .Z(n28861) );
  NOR U29155 ( .A(n156), .B(n129), .Z(n28859) );
  XOR U29156 ( .A(n28861), .B(n28859), .Z(n28863) );
  XOR U29157 ( .A(n28862), .B(n28863), .Z(n28851) );
  XOR U29158 ( .A(n28853), .B(n28851), .Z(n28856) );
  XOR U29159 ( .A(n28854), .B(n28856), .Z(n29009) );
  IV U29160 ( .A(n28821), .Z(n28822) );
  NOR U29161 ( .A(n28823), .B(n28822), .Z(n28827) );
  NOR U29162 ( .A(n28825), .B(n28824), .Z(n28826) );
  NOR U29163 ( .A(n28827), .B(n28826), .Z(n29008) );
  NOR U29164 ( .A(n161), .B(n124), .Z(n29006) );
  XOR U29165 ( .A(n29008), .B(n29006), .Z(n29010) );
  XOR U29166 ( .A(n29009), .B(n29010), .Z(n29013) );
  XOR U29167 ( .A(n29015), .B(n29013), .Z(n29018) );
  XOR U29168 ( .A(n29016), .B(n29018), .Z(n28847) );
  IV U29169 ( .A(n28828), .Z(n28829) );
  NOR U29170 ( .A(n28830), .B(n28829), .Z(n28834) );
  NOR U29171 ( .A(n28832), .B(n28831), .Z(n28833) );
  NOR U29172 ( .A(n28834), .B(n28833), .Z(n28845) );
  NOR U29173 ( .A(n165), .B(n121), .Z(n28843) );
  XOR U29174 ( .A(n28845), .B(n28843), .Z(n28846) );
  XOR U29175 ( .A(n28847), .B(n28846), .Z(n28835) );
  XOR U29176 ( .A(n28837), .B(n28835), .Z(n28840) );
  XOR U29177 ( .A(n28838), .B(n28840), .Z(n29027) );
  XOR U29178 ( .A(n29028), .B(n29027), .Z(n29392) );
  XOR U29179 ( .A(n29394), .B(n29392), .Z(n29023) );
  XOR U29180 ( .A(n29409), .B(n29023), .Z(c[102]) );
  IV U29181 ( .A(n28835), .Z(n28836) );
  NOR U29182 ( .A(n28837), .B(n28836), .Z(n28842) );
  IV U29183 ( .A(n28838), .Z(n28839) );
  NOR U29184 ( .A(n28840), .B(n28839), .Z(n28841) );
  NOR U29185 ( .A(n28842), .B(n28841), .Z(n29389) );
  IV U29186 ( .A(n28843), .Z(n28844) );
  NOR U29187 ( .A(n28845), .B(n28844), .Z(n28849) );
  NOR U29188 ( .A(n28847), .B(n28846), .Z(n28848) );
  NOR U29189 ( .A(n28849), .B(n28848), .Z(n29030) );
  NOR U29190 ( .A(n161), .B(n127), .Z(n28850) );
  IV U29191 ( .A(n28850), .Z(n29197) );
  IV U29192 ( .A(n28851), .Z(n28852) );
  NOR U29193 ( .A(n28853), .B(n28852), .Z(n28858) );
  IV U29194 ( .A(n28854), .Z(n28855) );
  NOR U29195 ( .A(n28856), .B(n28855), .Z(n28857) );
  NOR U29196 ( .A(n28858), .B(n28857), .Z(n29195) );
  NOR U29197 ( .A(n158), .B(n129), .Z(n29189) );
  IV U29198 ( .A(n28859), .Z(n28860) );
  NOR U29199 ( .A(n28861), .B(n28860), .Z(n28865) );
  NOR U29200 ( .A(n28863), .B(n28862), .Z(n28864) );
  NOR U29201 ( .A(n28865), .B(n28864), .Z(n29188) );
  NOR U29202 ( .A(n150), .B(n136), .Z(n29062) );
  IV U29203 ( .A(n28866), .Z(n28867) );
  NOR U29204 ( .A(n28868), .B(n28867), .Z(n28872) );
  NOR U29205 ( .A(n28870), .B(n28869), .Z(n28871) );
  NOR U29206 ( .A(n28872), .B(n28871), .Z(n29061) );
  IV U29207 ( .A(n28873), .Z(n28874) );
  NOR U29208 ( .A(n28875), .B(n28874), .Z(n28879) );
  NOR U29209 ( .A(n28877), .B(n28876), .Z(n28878) );
  NOR U29210 ( .A(n28879), .B(n28878), .Z(n28880) );
  IV U29211 ( .A(n28880), .Z(n29160) );
  NOR U29212 ( .A(n145), .B(n142), .Z(n29158) );
  XOR U29213 ( .A(n29160), .B(n29158), .Z(n29162) );
  NOR U29214 ( .A(n143), .B(n144), .Z(n28881) );
  IV U29215 ( .A(n28881), .Z(n29078) );
  IV U29216 ( .A(n28882), .Z(n28884) );
  NOR U29217 ( .A(n28884), .B(n28883), .Z(n28888) );
  NOR U29218 ( .A(n28886), .B(n28885), .Z(n28887) );
  NOR U29219 ( .A(n28888), .B(n28887), .Z(n29076) );
  NOR U29220 ( .A(n137), .B(n151), .Z(n28889) );
  IV U29221 ( .A(n28889), .Z(n29146) );
  IV U29222 ( .A(n28890), .Z(n28891) );
  NOR U29223 ( .A(n28892), .B(n28891), .Z(n28897) );
  IV U29224 ( .A(n28893), .Z(n28894) );
  NOR U29225 ( .A(n28895), .B(n28894), .Z(n28896) );
  NOR U29226 ( .A(n28897), .B(n28896), .Z(n29144) );
  NOR U29227 ( .A(n135), .B(n152), .Z(n29138) );
  IV U29228 ( .A(n28898), .Z(n28899) );
  NOR U29229 ( .A(n28900), .B(n28899), .Z(n28904) );
  NOR U29230 ( .A(n28902), .B(n28901), .Z(n28903) );
  NOR U29231 ( .A(n28904), .B(n28903), .Z(n29137) );
  IV U29232 ( .A(n29137), .Z(n28952) );
  NOR U29233 ( .A(n133), .B(n154), .Z(n28905) );
  IV U29234 ( .A(n28905), .Z(n29092) );
  IV U29235 ( .A(n28906), .Z(n28907) );
  NOR U29236 ( .A(n28908), .B(n28907), .Z(n28913) );
  IV U29237 ( .A(n28909), .Z(n28910) );
  NOR U29238 ( .A(n28911), .B(n28910), .Z(n28912) );
  NOR U29239 ( .A(n28913), .B(n28912), .Z(n29090) );
  NOR U29240 ( .A(n126), .B(n160), .Z(n29107) );
  IV U29241 ( .A(n28914), .Z(n28915) );
  NOR U29242 ( .A(n28916), .B(n28915), .Z(n28920) );
  NOR U29243 ( .A(n28918), .B(n28917), .Z(n28919) );
  NOR U29244 ( .A(n28920), .B(n28919), .Z(n29106) );
  NOR U29245 ( .A(n166), .B(n120), .Z(n29112) );
  IV U29246 ( .A(n29112), .Z(n28922) );
  NOR U29247 ( .A(n28922), .B(n28921), .Z(n28927) );
  IV U29248 ( .A(n28923), .Z(n28924) );
  NOR U29249 ( .A(n28925), .B(n28924), .Z(n28926) );
  NOR U29250 ( .A(n28927), .B(n28926), .Z(n29114) );
  NOR U29251 ( .A(n164), .B(n123), .Z(n29113) );
  XOR U29252 ( .A(n29113), .B(n29112), .Z(n28928) );
  XOR U29253 ( .A(n29114), .B(n28928), .Z(n29126) );
  IV U29254 ( .A(n28929), .Z(n28930) );
  NOR U29255 ( .A(n28931), .B(n28930), .Z(n28936) );
  IV U29256 ( .A(n28932), .Z(n28933) );
  NOR U29257 ( .A(n28934), .B(n28933), .Z(n28935) );
  NOR U29258 ( .A(n28936), .B(n28935), .Z(n29124) );
  NOR U29259 ( .A(n125), .B(n162), .Z(n29122) );
  XOR U29260 ( .A(n29124), .B(n29122), .Z(n29125) );
  XOR U29261 ( .A(n29126), .B(n29125), .Z(n29104) );
  XOR U29262 ( .A(n29106), .B(n29104), .Z(n29109) );
  XOR U29263 ( .A(n29107), .B(n29109), .Z(n29132) );
  IV U29264 ( .A(n28937), .Z(n28939) );
  NOR U29265 ( .A(n28939), .B(n28938), .Z(n28944) );
  IV U29266 ( .A(n28940), .Z(n28941) );
  NOR U29267 ( .A(n28942), .B(n28941), .Z(n28943) );
  NOR U29268 ( .A(n28944), .B(n28943), .Z(n29131) );
  NOR U29269 ( .A(n128), .B(n159), .Z(n29129) );
  XOR U29270 ( .A(n29131), .B(n29129), .Z(n29133) );
  XOR U29271 ( .A(n29132), .B(n29133), .Z(n29099) );
  IV U29272 ( .A(n28945), .Z(n28946) );
  NOR U29273 ( .A(n28947), .B(n28946), .Z(n28951) );
  NOR U29274 ( .A(n28949), .B(n28948), .Z(n28950) );
  NOR U29275 ( .A(n28951), .B(n28950), .Z(n29098) );
  NOR U29276 ( .A(n131), .B(n157), .Z(n29096) );
  XOR U29277 ( .A(n29098), .B(n29096), .Z(n29101) );
  XOR U29278 ( .A(n29099), .B(n29101), .Z(n29089) );
  XOR U29279 ( .A(n29090), .B(n29089), .Z(n29091) );
  XOR U29280 ( .A(n29092), .B(n29091), .Z(n29136) );
  XOR U29281 ( .A(n28952), .B(n29136), .Z(n29140) );
  XOR U29282 ( .A(n29138), .B(n29140), .Z(n29143) );
  XOR U29283 ( .A(n29144), .B(n29143), .Z(n29145) );
  XOR U29284 ( .A(n29146), .B(n29145), .Z(n29085) );
  IV U29285 ( .A(n28953), .Z(n28954) );
  NOR U29286 ( .A(n28955), .B(n28954), .Z(n28959) );
  NOR U29287 ( .A(n28957), .B(n28956), .Z(n28958) );
  NOR U29288 ( .A(n28959), .B(n28958), .Z(n29084) );
  NOR U29289 ( .A(n139), .B(n149), .Z(n29082) );
  XOR U29290 ( .A(n29084), .B(n29082), .Z(n29086) );
  XOR U29291 ( .A(n29085), .B(n29086), .Z(n29153) );
  IV U29292 ( .A(n28960), .Z(n28962) );
  NOR U29293 ( .A(n28962), .B(n28961), .Z(n28967) );
  IV U29294 ( .A(n28963), .Z(n28964) );
  NOR U29295 ( .A(n28965), .B(n28964), .Z(n28966) );
  NOR U29296 ( .A(n28967), .B(n28966), .Z(n29152) );
  NOR U29297 ( .A(n141), .B(n146), .Z(n29150) );
  XOR U29298 ( .A(n29152), .B(n29150), .Z(n29155) );
  XOR U29299 ( .A(n29153), .B(n29155), .Z(n29075) );
  XOR U29300 ( .A(n29076), .B(n29075), .Z(n29077) );
  XOR U29301 ( .A(n29078), .B(n29077), .Z(n29161) );
  XOR U29302 ( .A(n29162), .B(n29161), .Z(n29070) );
  IV U29303 ( .A(n28968), .Z(n28969) );
  NOR U29304 ( .A(n28970), .B(n28969), .Z(n28974) );
  NOR U29305 ( .A(n28972), .B(n28971), .Z(n28973) );
  NOR U29306 ( .A(n28974), .B(n28973), .Z(n29069) );
  NOR U29307 ( .A(n147), .B(n140), .Z(n29067) );
  XOR U29308 ( .A(n29069), .B(n29067), .Z(n29072) );
  XOR U29309 ( .A(n29070), .B(n29072), .Z(n29168) );
  IV U29310 ( .A(n28975), .Z(n28976) );
  NOR U29311 ( .A(n28977), .B(n28976), .Z(n28982) );
  IV U29312 ( .A(n28978), .Z(n28979) );
  NOR U29313 ( .A(n28980), .B(n28979), .Z(n28981) );
  NOR U29314 ( .A(n28982), .B(n28981), .Z(n29167) );
  NOR U29315 ( .A(n148), .B(n138), .Z(n29165) );
  XOR U29316 ( .A(n29167), .B(n29165), .Z(n29169) );
  XOR U29317 ( .A(n29168), .B(n29169), .Z(n29059) );
  XOR U29318 ( .A(n29061), .B(n29059), .Z(n29064) );
  XOR U29319 ( .A(n29062), .B(n29064), .Z(n29175) );
  IV U29320 ( .A(n28983), .Z(n28984) );
  NOR U29321 ( .A(n28985), .B(n28984), .Z(n28990) );
  IV U29322 ( .A(n28986), .Z(n28987) );
  NOR U29323 ( .A(n28988), .B(n28987), .Z(n28989) );
  NOR U29324 ( .A(n28990), .B(n28989), .Z(n29174) );
  NOR U29325 ( .A(n153), .B(n134), .Z(n29172) );
  XOR U29326 ( .A(n29174), .B(n29172), .Z(n29176) );
  XOR U29327 ( .A(n29175), .B(n29176), .Z(n29054) );
  IV U29328 ( .A(n28991), .Z(n28992) );
  NOR U29329 ( .A(n28993), .B(n28992), .Z(n28997) );
  NOR U29330 ( .A(n28995), .B(n28994), .Z(n28996) );
  NOR U29331 ( .A(n28997), .B(n28996), .Z(n29053) );
  NOR U29332 ( .A(n155), .B(n132), .Z(n29051) );
  XOR U29333 ( .A(n29053), .B(n29051), .Z(n29056) );
  XOR U29334 ( .A(n29054), .B(n29056), .Z(n29182) );
  IV U29335 ( .A(n28998), .Z(n28999) );
  NOR U29336 ( .A(n29000), .B(n28999), .Z(n29005) );
  IV U29337 ( .A(n29001), .Z(n29002) );
  NOR U29338 ( .A(n29003), .B(n29002), .Z(n29004) );
  NOR U29339 ( .A(n29005), .B(n29004), .Z(n29181) );
  NOR U29340 ( .A(n156), .B(n130), .Z(n29179) );
  XOR U29341 ( .A(n29181), .B(n29179), .Z(n29183) );
  XOR U29342 ( .A(n29182), .B(n29183), .Z(n29186) );
  XOR U29343 ( .A(n29188), .B(n29186), .Z(n29191) );
  XOR U29344 ( .A(n29189), .B(n29191), .Z(n29194) );
  XOR U29345 ( .A(n29195), .B(n29194), .Z(n29196) );
  XOR U29346 ( .A(n29197), .B(n29196), .Z(n29047) );
  IV U29347 ( .A(n29006), .Z(n29007) );
  NOR U29348 ( .A(n29008), .B(n29007), .Z(n29012) );
  NOR U29349 ( .A(n29010), .B(n29009), .Z(n29011) );
  NOR U29350 ( .A(n29012), .B(n29011), .Z(n29046) );
  NOR U29351 ( .A(n163), .B(n124), .Z(n29044) );
  XOR U29352 ( .A(n29046), .B(n29044), .Z(n29048) );
  XOR U29353 ( .A(n29047), .B(n29048), .Z(n29039) );
  IV U29354 ( .A(n29013), .Z(n29014) );
  NOR U29355 ( .A(n29015), .B(n29014), .Z(n29020) );
  IV U29356 ( .A(n29016), .Z(n29017) );
  NOR U29357 ( .A(n29018), .B(n29017), .Z(n29019) );
  NOR U29358 ( .A(n29020), .B(n29019), .Z(n29038) );
  NOR U29359 ( .A(n165), .B(n122), .Z(n29036) );
  XOR U29360 ( .A(n29038), .B(n29036), .Z(n29041) );
  XOR U29361 ( .A(n29039), .B(n29041), .Z(n29029) );
  XOR U29362 ( .A(n29030), .B(n29029), .Z(n29031) );
  NOR U29363 ( .A(n167), .B(n121), .Z(n29021) );
  IV U29364 ( .A(n29021), .Z(n29032) );
  XOR U29365 ( .A(n29031), .B(n29032), .Z(n29201) );
  IV U29366 ( .A(n29201), .Z(n29391) );
  XOR U29367 ( .A(n29389), .B(n29391), .Z(n29405) );
  NOR U29368 ( .A(n29022), .B(n29392), .Z(n29408) );
  IV U29369 ( .A(n29409), .Z(n29024) );
  NOR U29370 ( .A(n29024), .B(n29023), .Z(n29025) );
  NOR U29371 ( .A(n29408), .B(n29025), .Z(n29026) );
  IV U29372 ( .A(n29026), .Z(n29202) );
  NOR U29373 ( .A(n29028), .B(n29027), .Z(n29407) );
  XOR U29374 ( .A(n29202), .B(n29407), .Z(n29206) );
  XOR U29375 ( .A(n29405), .B(n29206), .Z(c[103]) );
  NOR U29376 ( .A(n29030), .B(n29029), .Z(n29035) );
  IV U29377 ( .A(n29031), .Z(n29033) );
  NOR U29378 ( .A(n29033), .B(n29032), .Z(n29034) );
  NOR U29379 ( .A(n29035), .B(n29034), .Z(n29382) );
  IV U29380 ( .A(n29036), .Z(n29037) );
  NOR U29381 ( .A(n29038), .B(n29037), .Z(n29043) );
  IV U29382 ( .A(n29039), .Z(n29040) );
  NOR U29383 ( .A(n29041), .B(n29040), .Z(n29042) );
  NOR U29384 ( .A(n29043), .B(n29042), .Z(n29214) );
  NOR U29385 ( .A(n167), .B(n122), .Z(n29212) );
  XOR U29386 ( .A(n29214), .B(n29212), .Z(n29216) );
  NOR U29387 ( .A(n165), .B(n124), .Z(n29222) );
  IV U29388 ( .A(n29044), .Z(n29045) );
  NOR U29389 ( .A(n29046), .B(n29045), .Z(n29050) );
  NOR U29390 ( .A(n29048), .B(n29047), .Z(n29049) );
  NOR U29391 ( .A(n29050), .B(n29049), .Z(n29221) );
  NOR U29392 ( .A(n156), .B(n132), .Z(n29244) );
  IV U29393 ( .A(n29051), .Z(n29052) );
  NOR U29394 ( .A(n29053), .B(n29052), .Z(n29058) );
  IV U29395 ( .A(n29054), .Z(n29055) );
  NOR U29396 ( .A(n29056), .B(n29055), .Z(n29057) );
  NOR U29397 ( .A(n29058), .B(n29057), .Z(n29243) );
  NOR U29398 ( .A(n153), .B(n136), .Z(n29253) );
  IV U29399 ( .A(n29059), .Z(n29060) );
  NOR U29400 ( .A(n29061), .B(n29060), .Z(n29066) );
  IV U29401 ( .A(n29062), .Z(n29063) );
  NOR U29402 ( .A(n29064), .B(n29063), .Z(n29065) );
  NOR U29403 ( .A(n29066), .B(n29065), .Z(n29252) );
  NOR U29404 ( .A(n148), .B(n140), .Z(n29352) );
  IV U29405 ( .A(n29067), .Z(n29068) );
  NOR U29406 ( .A(n29069), .B(n29068), .Z(n29074) );
  IV U29407 ( .A(n29070), .Z(n29071) );
  NOR U29408 ( .A(n29072), .B(n29071), .Z(n29073) );
  NOR U29409 ( .A(n29074), .B(n29073), .Z(n29351) );
  NOR U29410 ( .A(n145), .B(n144), .Z(n29344) );
  NOR U29411 ( .A(n29076), .B(n29075), .Z(n29081) );
  IV U29412 ( .A(n29077), .Z(n29079) );
  NOR U29413 ( .A(n29079), .B(n29078), .Z(n29080) );
  NOR U29414 ( .A(n29081), .B(n29080), .Z(n29343) );
  NOR U29415 ( .A(n141), .B(n149), .Z(n29275) );
  IV U29416 ( .A(n29082), .Z(n29083) );
  NOR U29417 ( .A(n29084), .B(n29083), .Z(n29088) );
  NOR U29418 ( .A(n29086), .B(n29085), .Z(n29087) );
  NOR U29419 ( .A(n29088), .B(n29087), .Z(n29274) );
  NOR U29420 ( .A(n29090), .B(n29089), .Z(n29095) );
  IV U29421 ( .A(n29091), .Z(n29093) );
  NOR U29422 ( .A(n29093), .B(n29092), .Z(n29094) );
  NOR U29423 ( .A(n29095), .B(n29094), .Z(n29330) );
  NOR U29424 ( .A(n135), .B(n154), .Z(n29326) );
  NOR U29425 ( .A(n133), .B(n157), .Z(n29292) );
  IV U29426 ( .A(n29096), .Z(n29097) );
  NOR U29427 ( .A(n29098), .B(n29097), .Z(n29103) );
  IV U29428 ( .A(n29099), .Z(n29100) );
  NOR U29429 ( .A(n29101), .B(n29100), .Z(n29102) );
  NOR U29430 ( .A(n29103), .B(n29102), .Z(n29291) );
  NOR U29431 ( .A(n128), .B(n160), .Z(n29321) );
  IV U29432 ( .A(n29104), .Z(n29105) );
  NOR U29433 ( .A(n29106), .B(n29105), .Z(n29111) );
  IV U29434 ( .A(n29107), .Z(n29108) );
  NOR U29435 ( .A(n29109), .B(n29108), .Z(n29110) );
  NOR U29436 ( .A(n29111), .B(n29110), .Z(n29320) );
  NOR U29437 ( .A(n29113), .B(n29112), .Z(n29115) );
  NOR U29438 ( .A(n29115), .B(n29114), .Z(n29120) );
  NOR U29439 ( .A(n29116), .B(n29120), .Z(n29118) );
  NOR U29440 ( .A(n166), .B(n123), .Z(n29119) );
  IV U29441 ( .A(n29119), .Z(n29117) );
  NOR U29442 ( .A(n29118), .B(n29117), .Z(n29315) );
  NOR U29443 ( .A(n29120), .B(n29119), .Z(n29121) );
  NOR U29444 ( .A(n29315), .B(n29121), .Z(n29311) );
  NOR U29445 ( .A(n125), .B(n164), .Z(n29517) );
  IV U29446 ( .A(n29517), .Z(n29313) );
  XOR U29447 ( .A(n29311), .B(n29313), .Z(n29307) );
  IV U29448 ( .A(n29122), .Z(n29123) );
  NOR U29449 ( .A(n29124), .B(n29123), .Z(n29128) );
  NOR U29450 ( .A(n29126), .B(n29125), .Z(n29127) );
  NOR U29451 ( .A(n29128), .B(n29127), .Z(n29306) );
  NOR U29452 ( .A(n126), .B(n162), .Z(n29304) );
  XOR U29453 ( .A(n29306), .B(n29304), .Z(n29308) );
  XOR U29454 ( .A(n29307), .B(n29308), .Z(n29318) );
  XOR U29455 ( .A(n29320), .B(n29318), .Z(n29323) );
  XOR U29456 ( .A(n29321), .B(n29323), .Z(n29301) );
  IV U29457 ( .A(n29129), .Z(n29130) );
  NOR U29458 ( .A(n29131), .B(n29130), .Z(n29135) );
  NOR U29459 ( .A(n29133), .B(n29132), .Z(n29134) );
  NOR U29460 ( .A(n29135), .B(n29134), .Z(n29299) );
  NOR U29461 ( .A(n131), .B(n159), .Z(n29297) );
  XOR U29462 ( .A(n29299), .B(n29297), .Z(n29300) );
  XOR U29463 ( .A(n29301), .B(n29300), .Z(n29289) );
  XOR U29464 ( .A(n29291), .B(n29289), .Z(n29294) );
  XOR U29465 ( .A(n29292), .B(n29294), .Z(n29328) );
  XOR U29466 ( .A(n29326), .B(n29328), .Z(n29329) );
  XOR U29467 ( .A(n29330), .B(n29329), .Z(n29283) );
  NOR U29468 ( .A(n29137), .B(n29136), .Z(n29142) );
  IV U29469 ( .A(n29138), .Z(n29139) );
  NOR U29470 ( .A(n29140), .B(n29139), .Z(n29141) );
  NOR U29471 ( .A(n29142), .B(n29141), .Z(n29282) );
  NOR U29472 ( .A(n137), .B(n152), .Z(n29280) );
  XOR U29473 ( .A(n29282), .B(n29280), .Z(n29285) );
  XOR U29474 ( .A(n29283), .B(n29285), .Z(n29336) );
  NOR U29475 ( .A(n29144), .B(n29143), .Z(n29149) );
  IV U29476 ( .A(n29145), .Z(n29147) );
  NOR U29477 ( .A(n29147), .B(n29146), .Z(n29148) );
  NOR U29478 ( .A(n29149), .B(n29148), .Z(n29335) );
  NOR U29479 ( .A(n139), .B(n151), .Z(n29333) );
  XOR U29480 ( .A(n29335), .B(n29333), .Z(n29337) );
  XOR U29481 ( .A(n29336), .B(n29337), .Z(n29272) );
  XOR U29482 ( .A(n29274), .B(n29272), .Z(n29277) );
  XOR U29483 ( .A(n29275), .B(n29277), .Z(n29268) );
  IV U29484 ( .A(n29150), .Z(n29151) );
  NOR U29485 ( .A(n29152), .B(n29151), .Z(n29157) );
  IV U29486 ( .A(n29153), .Z(n29154) );
  NOR U29487 ( .A(n29155), .B(n29154), .Z(n29156) );
  NOR U29488 ( .A(n29157), .B(n29156), .Z(n29267) );
  NOR U29489 ( .A(n143), .B(n146), .Z(n29265) );
  XOR U29490 ( .A(n29267), .B(n29265), .Z(n29269) );
  XOR U29491 ( .A(n29268), .B(n29269), .Z(n29341) );
  XOR U29492 ( .A(n29343), .B(n29341), .Z(n29346) );
  XOR U29493 ( .A(n29344), .B(n29346), .Z(n29262) );
  IV U29494 ( .A(n29158), .Z(n29159) );
  NOR U29495 ( .A(n29160), .B(n29159), .Z(n29164) );
  NOR U29496 ( .A(n29162), .B(n29161), .Z(n29163) );
  NOR U29497 ( .A(n29164), .B(n29163), .Z(n29260) );
  NOR U29498 ( .A(n147), .B(n142), .Z(n29258) );
  XOR U29499 ( .A(n29260), .B(n29258), .Z(n29261) );
  XOR U29500 ( .A(n29262), .B(n29261), .Z(n29349) );
  XOR U29501 ( .A(n29351), .B(n29349), .Z(n29354) );
  XOR U29502 ( .A(n29352), .B(n29354), .Z(n29360) );
  IV U29503 ( .A(n29165), .Z(n29166) );
  NOR U29504 ( .A(n29167), .B(n29166), .Z(n29171) );
  NOR U29505 ( .A(n29169), .B(n29168), .Z(n29170) );
  NOR U29506 ( .A(n29171), .B(n29170), .Z(n29359) );
  NOR U29507 ( .A(n150), .B(n138), .Z(n29357) );
  XOR U29508 ( .A(n29359), .B(n29357), .Z(n29361) );
  XOR U29509 ( .A(n29360), .B(n29361), .Z(n29250) );
  XOR U29510 ( .A(n29252), .B(n29250), .Z(n29255) );
  XOR U29511 ( .A(n29253), .B(n29255), .Z(n29368) );
  IV U29512 ( .A(n29172), .Z(n29173) );
  NOR U29513 ( .A(n29174), .B(n29173), .Z(n29178) );
  NOR U29514 ( .A(n29176), .B(n29175), .Z(n29177) );
  NOR U29515 ( .A(n29178), .B(n29177), .Z(n29366) );
  NOR U29516 ( .A(n155), .B(n134), .Z(n29364) );
  XOR U29517 ( .A(n29366), .B(n29364), .Z(n29367) );
  XOR U29518 ( .A(n29368), .B(n29367), .Z(n29241) );
  XOR U29519 ( .A(n29243), .B(n29241), .Z(n29246) );
  XOR U29520 ( .A(n29244), .B(n29246), .Z(n29237) );
  IV U29521 ( .A(n29179), .Z(n29180) );
  NOR U29522 ( .A(n29181), .B(n29180), .Z(n29185) );
  NOR U29523 ( .A(n29183), .B(n29182), .Z(n29184) );
  NOR U29524 ( .A(n29185), .B(n29184), .Z(n29236) );
  NOR U29525 ( .A(n158), .B(n130), .Z(n29234) );
  XOR U29526 ( .A(n29236), .B(n29234), .Z(n29238) );
  XOR U29527 ( .A(n29237), .B(n29238), .Z(n29375) );
  IV U29528 ( .A(n29186), .Z(n29187) );
  NOR U29529 ( .A(n29188), .B(n29187), .Z(n29193) );
  IV U29530 ( .A(n29189), .Z(n29190) );
  NOR U29531 ( .A(n29191), .B(n29190), .Z(n29192) );
  NOR U29532 ( .A(n29193), .B(n29192), .Z(n29374) );
  NOR U29533 ( .A(n161), .B(n129), .Z(n29372) );
  XOR U29534 ( .A(n29374), .B(n29372), .Z(n29377) );
  XOR U29535 ( .A(n29375), .B(n29377), .Z(n29230) );
  NOR U29536 ( .A(n29195), .B(n29194), .Z(n29200) );
  IV U29537 ( .A(n29196), .Z(n29198) );
  NOR U29538 ( .A(n29198), .B(n29197), .Z(n29199) );
  NOR U29539 ( .A(n29200), .B(n29199), .Z(n29229) );
  NOR U29540 ( .A(n163), .B(n127), .Z(n29227) );
  XOR U29541 ( .A(n29229), .B(n29227), .Z(n29231) );
  XOR U29542 ( .A(n29230), .B(n29231), .Z(n29219) );
  XOR U29543 ( .A(n29221), .B(n29219), .Z(n29224) );
  XOR U29544 ( .A(n29222), .B(n29224), .Z(n29215) );
  XOR U29545 ( .A(n29216), .B(n29215), .Z(n29383) );
  IV U29546 ( .A(n29383), .Z(n29380) );
  XOR U29547 ( .A(n29382), .B(n29380), .Z(n29403) );
  NOR U29548 ( .A(n29389), .B(n29201), .Z(n29404) );
  IV U29549 ( .A(n29404), .Z(n29205) );
  IV U29550 ( .A(n29407), .Z(n29203) );
  NOR U29551 ( .A(n29203), .B(n29202), .Z(n29208) );
  IV U29552 ( .A(n29208), .Z(n29204) );
  NOR U29553 ( .A(n29205), .B(n29204), .Z(n29381) );
  NOR U29554 ( .A(n29405), .B(n29206), .Z(n29207) );
  NOR U29555 ( .A(n29208), .B(n29207), .Z(n29209) );
  IV U29556 ( .A(n29209), .Z(n29210) );
  NOR U29557 ( .A(n29404), .B(n29210), .Z(n29385) );
  NOR U29558 ( .A(n29381), .B(n29385), .Z(n29211) );
  XOR U29559 ( .A(n29403), .B(n29211), .Z(c[104]) );
  IV U29560 ( .A(n29212), .Z(n29213) );
  NOR U29561 ( .A(n29214), .B(n29213), .Z(n29218) );
  NOR U29562 ( .A(n29216), .B(n29215), .Z(n29217) );
  NOR U29563 ( .A(n29218), .B(n29217), .Z(n29428) );
  IV U29564 ( .A(n29219), .Z(n29220) );
  NOR U29565 ( .A(n29221), .B(n29220), .Z(n29226) );
  IV U29566 ( .A(n29222), .Z(n29223) );
  NOR U29567 ( .A(n29224), .B(n29223), .Z(n29225) );
  NOR U29568 ( .A(n29226), .B(n29225), .Z(n29433) );
  NOR U29569 ( .A(n167), .B(n124), .Z(n29429) );
  NOR U29570 ( .A(n165), .B(n127), .Z(n29588) );
  IV U29571 ( .A(n29227), .Z(n29228) );
  NOR U29572 ( .A(n29229), .B(n29228), .Z(n29233) );
  NOR U29573 ( .A(n29231), .B(n29230), .Z(n29232) );
  NOR U29574 ( .A(n29233), .B(n29232), .Z(n29587) );
  NOR U29575 ( .A(n161), .B(n130), .Z(n29579) );
  IV U29576 ( .A(n29234), .Z(n29235) );
  NOR U29577 ( .A(n29236), .B(n29235), .Z(n29240) );
  NOR U29578 ( .A(n29238), .B(n29237), .Z(n29239) );
  NOR U29579 ( .A(n29240), .B(n29239), .Z(n29578) );
  IV U29580 ( .A(n29241), .Z(n29242) );
  NOR U29581 ( .A(n29243), .B(n29242), .Z(n29248) );
  IV U29582 ( .A(n29244), .Z(n29245) );
  NOR U29583 ( .A(n29246), .B(n29245), .Z(n29247) );
  NOR U29584 ( .A(n29248), .B(n29247), .Z(n29447) );
  NOR U29585 ( .A(n158), .B(n132), .Z(n29443) );
  NOR U29586 ( .A(n155), .B(n136), .Z(n29249) );
  IV U29587 ( .A(n29249), .Z(n29565) );
  IV U29588 ( .A(n29250), .Z(n29251) );
  NOR U29589 ( .A(n29252), .B(n29251), .Z(n29257) );
  IV U29590 ( .A(n29253), .Z(n29254) );
  NOR U29591 ( .A(n29255), .B(n29254), .Z(n29256) );
  NOR U29592 ( .A(n29257), .B(n29256), .Z(n29563) );
  NOR U29593 ( .A(n148), .B(n142), .Z(n29550) );
  IV U29594 ( .A(n29258), .Z(n29259) );
  NOR U29595 ( .A(n29260), .B(n29259), .Z(n29264) );
  NOR U29596 ( .A(n29262), .B(n29261), .Z(n29263) );
  NOR U29597 ( .A(n29264), .B(n29263), .Z(n29549) );
  NOR U29598 ( .A(n145), .B(n146), .Z(n29470) );
  IV U29599 ( .A(n29265), .Z(n29266) );
  NOR U29600 ( .A(n29267), .B(n29266), .Z(n29271) );
  NOR U29601 ( .A(n29269), .B(n29268), .Z(n29270) );
  NOR U29602 ( .A(n29271), .B(n29270), .Z(n29469) );
  IV U29603 ( .A(n29272), .Z(n29273) );
  NOR U29604 ( .A(n29274), .B(n29273), .Z(n29279) );
  IV U29605 ( .A(n29275), .Z(n29276) );
  NOR U29606 ( .A(n29277), .B(n29276), .Z(n29278) );
  NOR U29607 ( .A(n29279), .B(n29278), .Z(n29479) );
  NOR U29608 ( .A(n143), .B(n149), .Z(n29475) );
  NOR U29609 ( .A(n139), .B(n152), .Z(n29485) );
  IV U29610 ( .A(n29280), .Z(n29281) );
  NOR U29611 ( .A(n29282), .B(n29281), .Z(n29287) );
  IV U29612 ( .A(n29283), .Z(n29284) );
  NOR U29613 ( .A(n29285), .B(n29284), .Z(n29286) );
  NOR U29614 ( .A(n29287), .B(n29286), .Z(n29484) );
  NOR U29615 ( .A(n135), .B(n157), .Z(n29288) );
  IV U29616 ( .A(n29288), .Z(n29536) );
  IV U29617 ( .A(n29289), .Z(n29290) );
  NOR U29618 ( .A(n29291), .B(n29290), .Z(n29296) );
  IV U29619 ( .A(n29292), .Z(n29293) );
  NOR U29620 ( .A(n29294), .B(n29293), .Z(n29295) );
  NOR U29621 ( .A(n29296), .B(n29295), .Z(n29534) );
  NOR U29622 ( .A(n133), .B(n159), .Z(n29528) );
  IV U29623 ( .A(n29297), .Z(n29298) );
  NOR U29624 ( .A(n29299), .B(n29298), .Z(n29303) );
  NOR U29625 ( .A(n29301), .B(n29300), .Z(n29302) );
  NOR U29626 ( .A(n29303), .B(n29302), .Z(n29527) );
  NOR U29627 ( .A(n128), .B(n162), .Z(n29508) );
  IV U29628 ( .A(n29304), .Z(n29305) );
  NOR U29629 ( .A(n29306), .B(n29305), .Z(n29310) );
  NOR U29630 ( .A(n29308), .B(n29307), .Z(n29309) );
  NOR U29631 ( .A(n29310), .B(n29309), .Z(n29507) );
  IV U29632 ( .A(n29507), .Z(n29317) );
  IV U29633 ( .A(n29311), .Z(n29312) );
  NOR U29634 ( .A(n29313), .B(n29312), .Z(n29314) );
  NOR U29635 ( .A(n29315), .B(n29314), .Z(n29515) );
  NOR U29636 ( .A(n164), .B(n126), .Z(n29514) );
  NOR U29637 ( .A(n125), .B(n166), .Z(n29513) );
  XOR U29638 ( .A(n29514), .B(n29513), .Z(n29316) );
  XOR U29639 ( .A(n29515), .B(n29316), .Z(n29506) );
  XOR U29640 ( .A(n29317), .B(n29506), .Z(n29510) );
  XOR U29641 ( .A(n29508), .B(n29510), .Z(n29502) );
  IV U29642 ( .A(n29318), .Z(n29319) );
  NOR U29643 ( .A(n29320), .B(n29319), .Z(n29325) );
  IV U29644 ( .A(n29321), .Z(n29322) );
  NOR U29645 ( .A(n29323), .B(n29322), .Z(n29324) );
  NOR U29646 ( .A(n29325), .B(n29324), .Z(n29501) );
  NOR U29647 ( .A(n131), .B(n160), .Z(n29499) );
  XOR U29648 ( .A(n29501), .B(n29499), .Z(n29503) );
  XOR U29649 ( .A(n29502), .B(n29503), .Z(n29525) );
  XOR U29650 ( .A(n29527), .B(n29525), .Z(n29530) );
  XOR U29651 ( .A(n29528), .B(n29530), .Z(n29533) );
  XOR U29652 ( .A(n29534), .B(n29533), .Z(n29535) );
  XOR U29653 ( .A(n29536), .B(n29535), .Z(n29495) );
  IV U29654 ( .A(n29326), .Z(n29327) );
  NOR U29655 ( .A(n29328), .B(n29327), .Z(n29332) );
  NOR U29656 ( .A(n29330), .B(n29329), .Z(n29331) );
  NOR U29657 ( .A(n29332), .B(n29331), .Z(n29493) );
  NOR U29658 ( .A(n137), .B(n154), .Z(n29491) );
  XOR U29659 ( .A(n29493), .B(n29491), .Z(n29494) );
  XOR U29660 ( .A(n29495), .B(n29494), .Z(n29482) );
  XOR U29661 ( .A(n29484), .B(n29482), .Z(n29487) );
  XOR U29662 ( .A(n29485), .B(n29487), .Z(n29543) );
  IV U29663 ( .A(n29543), .Z(n29340) );
  IV U29664 ( .A(n29333), .Z(n29334) );
  NOR U29665 ( .A(n29335), .B(n29334), .Z(n29339) );
  NOR U29666 ( .A(n29337), .B(n29336), .Z(n29338) );
  NOR U29667 ( .A(n29339), .B(n29338), .Z(n29542) );
  NOR U29668 ( .A(n141), .B(n151), .Z(n29540) );
  XOR U29669 ( .A(n29542), .B(n29540), .Z(n29544) );
  XOR U29670 ( .A(n29340), .B(n29544), .Z(n29477) );
  XOR U29671 ( .A(n29475), .B(n29477), .Z(n29478) );
  XOR U29672 ( .A(n29479), .B(n29478), .Z(n29467) );
  XOR U29673 ( .A(n29469), .B(n29467), .Z(n29472) );
  XOR U29674 ( .A(n29470), .B(n29472), .Z(n29463) );
  IV U29675 ( .A(n29341), .Z(n29342) );
  NOR U29676 ( .A(n29343), .B(n29342), .Z(n29348) );
  IV U29677 ( .A(n29344), .Z(n29345) );
  NOR U29678 ( .A(n29346), .B(n29345), .Z(n29347) );
  NOR U29679 ( .A(n29348), .B(n29347), .Z(n29462) );
  NOR U29680 ( .A(n147), .B(n144), .Z(n29460) );
  XOR U29681 ( .A(n29462), .B(n29460), .Z(n29464) );
  XOR U29682 ( .A(n29463), .B(n29464), .Z(n29547) );
  XOR U29683 ( .A(n29549), .B(n29547), .Z(n29552) );
  XOR U29684 ( .A(n29550), .B(n29552), .Z(n29559) );
  IV U29685 ( .A(n29349), .Z(n29350) );
  NOR U29686 ( .A(n29351), .B(n29350), .Z(n29356) );
  IV U29687 ( .A(n29352), .Z(n29353) );
  NOR U29688 ( .A(n29354), .B(n29353), .Z(n29355) );
  NOR U29689 ( .A(n29356), .B(n29355), .Z(n29557) );
  NOR U29690 ( .A(n150), .B(n140), .Z(n29555) );
  XOR U29691 ( .A(n29557), .B(n29555), .Z(n29558) );
  XOR U29692 ( .A(n29559), .B(n29558), .Z(n29454) );
  IV U29693 ( .A(n29357), .Z(n29358) );
  NOR U29694 ( .A(n29359), .B(n29358), .Z(n29363) );
  NOR U29695 ( .A(n29361), .B(n29360), .Z(n29362) );
  NOR U29696 ( .A(n29363), .B(n29362), .Z(n29453) );
  NOR U29697 ( .A(n153), .B(n138), .Z(n29451) );
  XOR U29698 ( .A(n29453), .B(n29451), .Z(n29456) );
  XOR U29699 ( .A(n29454), .B(n29456), .Z(n29562) );
  XOR U29700 ( .A(n29563), .B(n29562), .Z(n29564) );
  XOR U29701 ( .A(n29565), .B(n29564), .Z(n29572) );
  IV U29702 ( .A(n29572), .Z(n29371) );
  IV U29703 ( .A(n29364), .Z(n29365) );
  NOR U29704 ( .A(n29366), .B(n29365), .Z(n29370) );
  NOR U29705 ( .A(n29368), .B(n29367), .Z(n29369) );
  NOR U29706 ( .A(n29370), .B(n29369), .Z(n29571) );
  NOR U29707 ( .A(n156), .B(n134), .Z(n29569) );
  XOR U29708 ( .A(n29571), .B(n29569), .Z(n29573) );
  XOR U29709 ( .A(n29371), .B(n29573), .Z(n29445) );
  XOR U29710 ( .A(n29443), .B(n29445), .Z(n29446) );
  XOR U29711 ( .A(n29447), .B(n29446), .Z(n29576) );
  XOR U29712 ( .A(n29578), .B(n29576), .Z(n29581) );
  XOR U29713 ( .A(n29579), .B(n29581), .Z(n29439) );
  IV U29714 ( .A(n29372), .Z(n29373) );
  NOR U29715 ( .A(n29374), .B(n29373), .Z(n29379) );
  IV U29716 ( .A(n29375), .Z(n29376) );
  NOR U29717 ( .A(n29377), .B(n29376), .Z(n29378) );
  NOR U29718 ( .A(n29379), .B(n29378), .Z(n29438) );
  NOR U29719 ( .A(n163), .B(n129), .Z(n29436) );
  XOR U29720 ( .A(n29438), .B(n29436), .Z(n29440) );
  XOR U29721 ( .A(n29439), .B(n29440), .Z(n29585) );
  XOR U29722 ( .A(n29587), .B(n29585), .Z(n29590) );
  XOR U29723 ( .A(n29588), .B(n29590), .Z(n29431) );
  XOR U29724 ( .A(n29429), .B(n29431), .Z(n29432) );
  XOR U29725 ( .A(n29433), .B(n29432), .Z(n29426) );
  XOR U29726 ( .A(n29428), .B(n29426), .Z(n29423) );
  NOR U29727 ( .A(n29380), .B(n29382), .Z(n29421) );
  XOR U29728 ( .A(n29381), .B(n29421), .Z(n29387) );
  XOR U29729 ( .A(n29383), .B(n29382), .Z(n29384) );
  NOR U29730 ( .A(n29385), .B(n29384), .Z(n29386) );
  NOR U29731 ( .A(n29387), .B(n29386), .Z(n29388) );
  XOR U29732 ( .A(n29423), .B(n29388), .Z(c[105]) );
  IV U29733 ( .A(n29389), .Z(n29390) );
  NOR U29734 ( .A(n29391), .B(n29390), .Z(n29402) );
  IV U29735 ( .A(n29392), .Z(n29393) );
  NOR U29736 ( .A(n29394), .B(n29393), .Z(n29397) );
  NOR U29737 ( .A(n29407), .B(n29404), .Z(n29395) );
  IV U29738 ( .A(n29395), .Z(n29396) );
  NOR U29739 ( .A(n29397), .B(n29396), .Z(n29399) );
  IV U29740 ( .A(n29403), .Z(n29398) );
  NOR U29741 ( .A(n29399), .B(n29398), .Z(n29400) );
  IV U29742 ( .A(n29400), .Z(n29401) );
  NOR U29743 ( .A(n29402), .B(n29401), .Z(n29417) );
  NOR U29744 ( .A(n29404), .B(n29403), .Z(n29415) );
  IV U29745 ( .A(n29405), .Z(n29406) );
  NOR U29746 ( .A(n29407), .B(n29406), .Z(n29412) );
  NOR U29747 ( .A(n29409), .B(n29408), .Z(n29410) );
  IV U29748 ( .A(n29410), .Z(n29411) );
  NOR U29749 ( .A(n29412), .B(n29411), .Z(n29413) );
  IV U29750 ( .A(n29413), .Z(n29414) );
  NOR U29751 ( .A(n29415), .B(n29414), .Z(n29416) );
  NOR U29752 ( .A(n29417), .B(n29416), .Z(n29419) );
  IV U29753 ( .A(n29421), .Z(n29418) );
  NOR U29754 ( .A(n29419), .B(n29418), .Z(n29425) );
  IV U29755 ( .A(n29419), .Z(n29420) );
  NOR U29756 ( .A(n29421), .B(n29420), .Z(n29422) );
  NOR U29757 ( .A(n29423), .B(n29422), .Z(n29424) );
  NOR U29758 ( .A(n29425), .B(n29424), .Z(n29748) );
  IV U29759 ( .A(n29426), .Z(n29427) );
  NOR U29760 ( .A(n29428), .B(n29427), .Z(n29747) );
  IV U29761 ( .A(n29747), .Z(n29752) );
  IV U29762 ( .A(n29429), .Z(n29430) );
  NOR U29763 ( .A(n29431), .B(n29430), .Z(n29435) );
  NOR U29764 ( .A(n29433), .B(n29432), .Z(n29434) );
  NOR U29765 ( .A(n29435), .B(n29434), .Z(n29743) );
  NOR U29766 ( .A(n165), .B(n129), .Z(n29737) );
  IV U29767 ( .A(n29436), .Z(n29437) );
  NOR U29768 ( .A(n29438), .B(n29437), .Z(n29442) );
  NOR U29769 ( .A(n29440), .B(n29439), .Z(n29441) );
  NOR U29770 ( .A(n29442), .B(n29441), .Z(n29736) );
  IV U29771 ( .A(n29443), .Z(n29444) );
  NOR U29772 ( .A(n29445), .B(n29444), .Z(n29449) );
  NOR U29773 ( .A(n29447), .B(n29446), .Z(n29448) );
  NOR U29774 ( .A(n29449), .B(n29448), .Z(n29731) );
  NOR U29775 ( .A(n161), .B(n132), .Z(n29727) );
  NOR U29776 ( .A(n155), .B(n138), .Z(n29450) );
  IV U29777 ( .A(n29450), .Z(n29708) );
  IV U29778 ( .A(n29451), .Z(n29452) );
  NOR U29779 ( .A(n29453), .B(n29452), .Z(n29458) );
  IV U29780 ( .A(n29454), .Z(n29455) );
  NOR U29781 ( .A(n29456), .B(n29455), .Z(n29457) );
  NOR U29782 ( .A(n29458), .B(n29457), .Z(n29706) );
  NOR U29783 ( .A(n148), .B(n144), .Z(n29459) );
  IV U29784 ( .A(n29459), .Z(n29694) );
  IV U29785 ( .A(n29460), .Z(n29461) );
  NOR U29786 ( .A(n29462), .B(n29461), .Z(n29466) );
  NOR U29787 ( .A(n29464), .B(n29463), .Z(n29465) );
  NOR U29788 ( .A(n29466), .B(n29465), .Z(n29692) );
  NOR U29789 ( .A(n147), .B(n146), .Z(n29621) );
  IV U29790 ( .A(n29467), .Z(n29468) );
  NOR U29791 ( .A(n29469), .B(n29468), .Z(n29474) );
  IV U29792 ( .A(n29470), .Z(n29471) );
  NOR U29793 ( .A(n29472), .B(n29471), .Z(n29473) );
  NOR U29794 ( .A(n29474), .B(n29473), .Z(n29620) );
  IV U29795 ( .A(n29475), .Z(n29476) );
  NOR U29796 ( .A(n29477), .B(n29476), .Z(n29481) );
  NOR U29797 ( .A(n29479), .B(n29478), .Z(n29480) );
  NOR U29798 ( .A(n29481), .B(n29480), .Z(n29630) );
  NOR U29799 ( .A(n145), .B(n149), .Z(n29626) );
  IV U29800 ( .A(n29482), .Z(n29483) );
  NOR U29801 ( .A(n29484), .B(n29483), .Z(n29489) );
  IV U29802 ( .A(n29485), .Z(n29486) );
  NOR U29803 ( .A(n29487), .B(n29486), .Z(n29488) );
  NOR U29804 ( .A(n29489), .B(n29488), .Z(n29686) );
  NOR U29805 ( .A(n141), .B(n152), .Z(n29682) );
  NOR U29806 ( .A(n139), .B(n154), .Z(n29490) );
  IV U29807 ( .A(n29490), .Z(n29644) );
  IV U29808 ( .A(n29491), .Z(n29492) );
  NOR U29809 ( .A(n29493), .B(n29492), .Z(n29497) );
  NOR U29810 ( .A(n29495), .B(n29494), .Z(n29496) );
  NOR U29811 ( .A(n29497), .B(n29496), .Z(n29642) );
  NOR U29812 ( .A(n133), .B(n160), .Z(n29498) );
  IV U29813 ( .A(n29498), .Z(n29671) );
  IV U29814 ( .A(n29499), .Z(n29500) );
  NOR U29815 ( .A(n29501), .B(n29500), .Z(n29505) );
  NOR U29816 ( .A(n29503), .B(n29502), .Z(n29504) );
  NOR U29817 ( .A(n29505), .B(n29504), .Z(n29669) );
  NOR U29818 ( .A(n131), .B(n162), .Z(n29663) );
  NOR U29819 ( .A(n29507), .B(n29506), .Z(n29512) );
  IV U29820 ( .A(n29508), .Z(n29509) );
  NOR U29821 ( .A(n29510), .B(n29509), .Z(n29511) );
  NOR U29822 ( .A(n29512), .B(n29511), .Z(n29662) );
  IV U29823 ( .A(n29662), .Z(n29524) );
  NOR U29824 ( .A(n29514), .B(n29513), .Z(n29516) );
  NOR U29825 ( .A(n29516), .B(n29515), .Z(n29521) );
  NOR U29826 ( .A(n29517), .B(n29521), .Z(n29519) );
  NOR U29827 ( .A(n126), .B(n166), .Z(n29520) );
  IV U29828 ( .A(n29520), .Z(n29518) );
  NOR U29829 ( .A(n29519), .B(n29518), .Z(n29660) );
  NOR U29830 ( .A(n29521), .B(n29520), .Z(n29522) );
  NOR U29831 ( .A(n29660), .B(n29522), .Z(n29523) );
  IV U29832 ( .A(n29523), .Z(n29658) );
  NOR U29833 ( .A(n164), .B(n128), .Z(n29656) );
  XOR U29834 ( .A(n29658), .B(n29656), .Z(n29661) );
  XOR U29835 ( .A(n29524), .B(n29661), .Z(n29665) );
  XOR U29836 ( .A(n29663), .B(n29665), .Z(n29668) );
  XOR U29837 ( .A(n29669), .B(n29668), .Z(n29670) );
  XOR U29838 ( .A(n29671), .B(n29670), .Z(n29678) );
  IV U29839 ( .A(n29525), .Z(n29526) );
  NOR U29840 ( .A(n29527), .B(n29526), .Z(n29532) );
  IV U29841 ( .A(n29528), .Z(n29529) );
  NOR U29842 ( .A(n29530), .B(n29529), .Z(n29531) );
  NOR U29843 ( .A(n29532), .B(n29531), .Z(n29677) );
  NOR U29844 ( .A(n135), .B(n159), .Z(n29675) );
  XOR U29845 ( .A(n29677), .B(n29675), .Z(n29679) );
  XOR U29846 ( .A(n29678), .B(n29679), .Z(n29651) );
  NOR U29847 ( .A(n29534), .B(n29533), .Z(n29539) );
  IV U29848 ( .A(n29535), .Z(n29537) );
  NOR U29849 ( .A(n29537), .B(n29536), .Z(n29538) );
  NOR U29850 ( .A(n29539), .B(n29538), .Z(n29650) );
  NOR U29851 ( .A(n137), .B(n157), .Z(n29648) );
  XOR U29852 ( .A(n29650), .B(n29648), .Z(n29653) );
  XOR U29853 ( .A(n29651), .B(n29653), .Z(n29641) );
  XOR U29854 ( .A(n29642), .B(n29641), .Z(n29643) );
  XOR U29855 ( .A(n29644), .B(n29643), .Z(n29684) );
  XOR U29856 ( .A(n29682), .B(n29684), .Z(n29685) );
  XOR U29857 ( .A(n29686), .B(n29685), .Z(n29636) );
  IV U29858 ( .A(n29540), .Z(n29541) );
  NOR U29859 ( .A(n29542), .B(n29541), .Z(n29546) );
  NOR U29860 ( .A(n29544), .B(n29543), .Z(n29545) );
  NOR U29861 ( .A(n29546), .B(n29545), .Z(n29635) );
  NOR U29862 ( .A(n143), .B(n151), .Z(n29633) );
  XOR U29863 ( .A(n29635), .B(n29633), .Z(n29638) );
  XOR U29864 ( .A(n29636), .B(n29638), .Z(n29628) );
  XOR U29865 ( .A(n29626), .B(n29628), .Z(n29629) );
  XOR U29866 ( .A(n29630), .B(n29629), .Z(n29618) );
  XOR U29867 ( .A(n29620), .B(n29618), .Z(n29623) );
  XOR U29868 ( .A(n29621), .B(n29623), .Z(n29691) );
  XOR U29869 ( .A(n29692), .B(n29691), .Z(n29693) );
  XOR U29870 ( .A(n29694), .B(n29693), .Z(n29701) );
  IV U29871 ( .A(n29547), .Z(n29548) );
  NOR U29872 ( .A(n29549), .B(n29548), .Z(n29554) );
  IV U29873 ( .A(n29550), .Z(n29551) );
  NOR U29874 ( .A(n29552), .B(n29551), .Z(n29553) );
  NOR U29875 ( .A(n29554), .B(n29553), .Z(n29700) );
  NOR U29876 ( .A(n150), .B(n142), .Z(n29698) );
  XOR U29877 ( .A(n29700), .B(n29698), .Z(n29702) );
  XOR U29878 ( .A(n29701), .B(n29702), .Z(n29613) );
  IV U29879 ( .A(n29555), .Z(n29556) );
  NOR U29880 ( .A(n29557), .B(n29556), .Z(n29561) );
  NOR U29881 ( .A(n29559), .B(n29558), .Z(n29560) );
  NOR U29882 ( .A(n29561), .B(n29560), .Z(n29612) );
  NOR U29883 ( .A(n153), .B(n140), .Z(n29610) );
  XOR U29884 ( .A(n29612), .B(n29610), .Z(n29615) );
  XOR U29885 ( .A(n29613), .B(n29615), .Z(n29705) );
  XOR U29886 ( .A(n29706), .B(n29705), .Z(n29707) );
  XOR U29887 ( .A(n29708), .B(n29707), .Z(n29715) );
  NOR U29888 ( .A(n29563), .B(n29562), .Z(n29568) );
  IV U29889 ( .A(n29564), .Z(n29566) );
  NOR U29890 ( .A(n29566), .B(n29565), .Z(n29567) );
  NOR U29891 ( .A(n29568), .B(n29567), .Z(n29714) );
  NOR U29892 ( .A(n156), .B(n136), .Z(n29712) );
  XOR U29893 ( .A(n29714), .B(n29712), .Z(n29716) );
  XOR U29894 ( .A(n29715), .B(n29716), .Z(n29722) );
  IV U29895 ( .A(n29569), .Z(n29570) );
  NOR U29896 ( .A(n29571), .B(n29570), .Z(n29575) );
  NOR U29897 ( .A(n29573), .B(n29572), .Z(n29574) );
  NOR U29898 ( .A(n29575), .B(n29574), .Z(n29721) );
  NOR U29899 ( .A(n158), .B(n134), .Z(n29719) );
  XOR U29900 ( .A(n29721), .B(n29719), .Z(n29724) );
  XOR U29901 ( .A(n29722), .B(n29724), .Z(n29729) );
  XOR U29902 ( .A(n29727), .B(n29729), .Z(n29730) );
  XOR U29903 ( .A(n29731), .B(n29730), .Z(n29605) );
  IV U29904 ( .A(n29576), .Z(n29577) );
  NOR U29905 ( .A(n29578), .B(n29577), .Z(n29583) );
  IV U29906 ( .A(n29579), .Z(n29580) );
  NOR U29907 ( .A(n29581), .B(n29580), .Z(n29582) );
  NOR U29908 ( .A(n29583), .B(n29582), .Z(n29604) );
  NOR U29909 ( .A(n163), .B(n130), .Z(n29602) );
  XOR U29910 ( .A(n29604), .B(n29602), .Z(n29607) );
  XOR U29911 ( .A(n29605), .B(n29607), .Z(n29735) );
  XOR U29912 ( .A(n29736), .B(n29735), .Z(n29584) );
  IV U29913 ( .A(n29584), .Z(n29739) );
  XOR U29914 ( .A(n29737), .B(n29739), .Z(n29598) );
  IV U29915 ( .A(n29585), .Z(n29586) );
  NOR U29916 ( .A(n29587), .B(n29586), .Z(n29592) );
  IV U29917 ( .A(n29588), .Z(n29589) );
  NOR U29918 ( .A(n29590), .B(n29589), .Z(n29591) );
  NOR U29919 ( .A(n29592), .B(n29591), .Z(n29597) );
  NOR U29920 ( .A(n167), .B(n127), .Z(n29595) );
  XOR U29921 ( .A(n29597), .B(n29595), .Z(n29599) );
  XOR U29922 ( .A(n29598), .B(n29599), .Z(n29593) );
  IV U29923 ( .A(n29593), .Z(n29742) );
  XOR U29924 ( .A(n29743), .B(n29742), .Z(n29750) );
  XOR U29925 ( .A(n29752), .B(n29750), .Z(n29594) );
  XOR U29926 ( .A(n29748), .B(n29594), .Z(c[106]) );
  IV U29927 ( .A(n29595), .Z(n29596) );
  NOR U29928 ( .A(n29597), .B(n29596), .Z(n29601) );
  NOR U29929 ( .A(n29599), .B(n29598), .Z(n29600) );
  NOR U29930 ( .A(n29601), .B(n29600), .Z(n30074) );
  IV U29931 ( .A(n29602), .Z(n29603) );
  NOR U29932 ( .A(n29604), .B(n29603), .Z(n29609) );
  IV U29933 ( .A(n29605), .Z(n29606) );
  NOR U29934 ( .A(n29607), .B(n29606), .Z(n29608) );
  NOR U29935 ( .A(n29609), .B(n29608), .Z(n29769) );
  NOR U29936 ( .A(n165), .B(n130), .Z(n29765) );
  NOR U29937 ( .A(n155), .B(n140), .Z(n29878) );
  IV U29938 ( .A(n29610), .Z(n29611) );
  NOR U29939 ( .A(n29612), .B(n29611), .Z(n29617) );
  IV U29940 ( .A(n29613), .Z(n29614) );
  NOR U29941 ( .A(n29615), .B(n29614), .Z(n29616) );
  NOR U29942 ( .A(n29617), .B(n29616), .Z(n29877) );
  IV U29943 ( .A(n29618), .Z(n29619) );
  NOR U29944 ( .A(n29620), .B(n29619), .Z(n29625) );
  IV U29945 ( .A(n29621), .Z(n29622) );
  NOR U29946 ( .A(n29623), .B(n29622), .Z(n29624) );
  NOR U29947 ( .A(n29625), .B(n29624), .Z(n29793) );
  NOR U29948 ( .A(n148), .B(n146), .Z(n29789) );
  NOR U29949 ( .A(n147), .B(n149), .Z(n29862) );
  IV U29950 ( .A(n29626), .Z(n29627) );
  NOR U29951 ( .A(n29628), .B(n29627), .Z(n29632) );
  NOR U29952 ( .A(n29630), .B(n29629), .Z(n29631) );
  NOR U29953 ( .A(n29632), .B(n29631), .Z(n29861) );
  IV U29954 ( .A(n29861), .Z(n29690) );
  NOR U29955 ( .A(n145), .B(n151), .Z(n29855) );
  IV U29956 ( .A(n29633), .Z(n29634) );
  NOR U29957 ( .A(n29635), .B(n29634), .Z(n29640) );
  IV U29958 ( .A(n29636), .Z(n29637) );
  NOR U29959 ( .A(n29638), .B(n29637), .Z(n29639) );
  NOR U29960 ( .A(n29640), .B(n29639), .Z(n29854) );
  NOR U29961 ( .A(n29642), .B(n29641), .Z(n29647) );
  IV U29962 ( .A(n29643), .Z(n29645) );
  NOR U29963 ( .A(n29645), .B(n29644), .Z(n29646) );
  NOR U29964 ( .A(n29647), .B(n29646), .Z(n29849) );
  NOR U29965 ( .A(n141), .B(n154), .Z(n29845) );
  NOR U29966 ( .A(n139), .B(n157), .Z(n29840) );
  IV U29967 ( .A(n29648), .Z(n29649) );
  NOR U29968 ( .A(n29650), .B(n29649), .Z(n29655) );
  IV U29969 ( .A(n29651), .Z(n29652) );
  NOR U29970 ( .A(n29653), .B(n29652), .Z(n29654) );
  NOR U29971 ( .A(n29655), .B(n29654), .Z(n29839) );
  NOR U29972 ( .A(n164), .B(n131), .Z(n29823) );
  IV U29973 ( .A(n29656), .Z(n29657) );
  NOR U29974 ( .A(n29658), .B(n29657), .Z(n29659) );
  NOR U29975 ( .A(n29660), .B(n29659), .Z(n29822) );
  NOR U29976 ( .A(n166), .B(n128), .Z(n29820) );
  XOR U29977 ( .A(n29822), .B(n29820), .Z(n29825) );
  XOR U29978 ( .A(n29823), .B(n29825), .Z(n29816) );
  NOR U29979 ( .A(n29662), .B(n29661), .Z(n29667) );
  IV U29980 ( .A(n29663), .Z(n29664) );
  NOR U29981 ( .A(n29665), .B(n29664), .Z(n29666) );
  NOR U29982 ( .A(n29667), .B(n29666), .Z(n29815) );
  NOR U29983 ( .A(n133), .B(n162), .Z(n29813) );
  XOR U29984 ( .A(n29815), .B(n29813), .Z(n29817) );
  XOR U29985 ( .A(n29816), .B(n29817), .Z(n29807) );
  NOR U29986 ( .A(n29669), .B(n29668), .Z(n29674) );
  IV U29987 ( .A(n29670), .Z(n29672) );
  NOR U29988 ( .A(n29672), .B(n29671), .Z(n29673) );
  NOR U29989 ( .A(n29674), .B(n29673), .Z(n29806) );
  NOR U29990 ( .A(n135), .B(n160), .Z(n29804) );
  XOR U29991 ( .A(n29806), .B(n29804), .Z(n29809) );
  XOR U29992 ( .A(n29807), .B(n29809), .Z(n29833) );
  IV U29993 ( .A(n29675), .Z(n29676) );
  NOR U29994 ( .A(n29677), .B(n29676), .Z(n29681) );
  NOR U29995 ( .A(n29679), .B(n29678), .Z(n29680) );
  NOR U29996 ( .A(n29681), .B(n29680), .Z(n29832) );
  NOR U29997 ( .A(n137), .B(n159), .Z(n29830) );
  XOR U29998 ( .A(n29832), .B(n29830), .Z(n29834) );
  XOR U29999 ( .A(n29833), .B(n29834), .Z(n29837) );
  XOR U30000 ( .A(n29839), .B(n29837), .Z(n29842) );
  XOR U30001 ( .A(n29840), .B(n29842), .Z(n29847) );
  XOR U30002 ( .A(n29845), .B(n29847), .Z(n29848) );
  XOR U30003 ( .A(n29849), .B(n29848), .Z(n29799) );
  IV U30004 ( .A(n29682), .Z(n29683) );
  NOR U30005 ( .A(n29684), .B(n29683), .Z(n29688) );
  NOR U30006 ( .A(n29686), .B(n29685), .Z(n29687) );
  NOR U30007 ( .A(n29688), .B(n29687), .Z(n29798) );
  NOR U30008 ( .A(n143), .B(n152), .Z(n29796) );
  XOR U30009 ( .A(n29798), .B(n29796), .Z(n29800) );
  XOR U30010 ( .A(n29799), .B(n29800), .Z(n29853) );
  XOR U30011 ( .A(n29854), .B(n29853), .Z(n29689) );
  IV U30012 ( .A(n29689), .Z(n29857) );
  XOR U30013 ( .A(n29855), .B(n29857), .Z(n29860) );
  XOR U30014 ( .A(n29690), .B(n29860), .Z(n29864) );
  XOR U30015 ( .A(n29862), .B(n29864), .Z(n29791) );
  XOR U30016 ( .A(n29789), .B(n29791), .Z(n29792) );
  XOR U30017 ( .A(n29793), .B(n29792), .Z(n29870) );
  NOR U30018 ( .A(n29692), .B(n29691), .Z(n29697) );
  IV U30019 ( .A(n29693), .Z(n29695) );
  NOR U30020 ( .A(n29695), .B(n29694), .Z(n29696) );
  NOR U30021 ( .A(n29697), .B(n29696), .Z(n29869) );
  NOR U30022 ( .A(n150), .B(n144), .Z(n29867) );
  XOR U30023 ( .A(n29869), .B(n29867), .Z(n29872) );
  XOR U30024 ( .A(n29870), .B(n29872), .Z(n29784) );
  IV U30025 ( .A(n29698), .Z(n29699) );
  NOR U30026 ( .A(n29700), .B(n29699), .Z(n29704) );
  NOR U30027 ( .A(n29702), .B(n29701), .Z(n29703) );
  NOR U30028 ( .A(n29704), .B(n29703), .Z(n29783) );
  NOR U30029 ( .A(n153), .B(n142), .Z(n29781) );
  XOR U30030 ( .A(n29783), .B(n29781), .Z(n29785) );
  XOR U30031 ( .A(n29784), .B(n29785), .Z(n29875) );
  XOR U30032 ( .A(n29877), .B(n29875), .Z(n29880) );
  XOR U30033 ( .A(n29878), .B(n29880), .Z(n29886) );
  NOR U30034 ( .A(n29706), .B(n29705), .Z(n29711) );
  IV U30035 ( .A(n29707), .Z(n29709) );
  NOR U30036 ( .A(n29709), .B(n29708), .Z(n29710) );
  NOR U30037 ( .A(n29711), .B(n29710), .Z(n29885) );
  NOR U30038 ( .A(n156), .B(n138), .Z(n29883) );
  XOR U30039 ( .A(n29885), .B(n29883), .Z(n29887) );
  XOR U30040 ( .A(n29886), .B(n29887), .Z(n29776) );
  IV U30041 ( .A(n29712), .Z(n29713) );
  NOR U30042 ( .A(n29714), .B(n29713), .Z(n29718) );
  NOR U30043 ( .A(n29716), .B(n29715), .Z(n29717) );
  NOR U30044 ( .A(n29718), .B(n29717), .Z(n29775) );
  NOR U30045 ( .A(n158), .B(n136), .Z(n29773) );
  XOR U30046 ( .A(n29775), .B(n29773), .Z(n29778) );
  XOR U30047 ( .A(n29776), .B(n29778), .Z(n29893) );
  IV U30048 ( .A(n29719), .Z(n29720) );
  NOR U30049 ( .A(n29721), .B(n29720), .Z(n29726) );
  IV U30050 ( .A(n29722), .Z(n29723) );
  NOR U30051 ( .A(n29724), .B(n29723), .Z(n29725) );
  NOR U30052 ( .A(n29726), .B(n29725), .Z(n29892) );
  NOR U30053 ( .A(n161), .B(n134), .Z(n29890) );
  XOR U30054 ( .A(n29892), .B(n29890), .Z(n29894) );
  XOR U30055 ( .A(n29893), .B(n29894), .Z(n29900) );
  IV U30056 ( .A(n29727), .Z(n29728) );
  NOR U30057 ( .A(n29729), .B(n29728), .Z(n29733) );
  NOR U30058 ( .A(n29731), .B(n29730), .Z(n29732) );
  NOR U30059 ( .A(n29733), .B(n29732), .Z(n29899) );
  NOR U30060 ( .A(n163), .B(n132), .Z(n29897) );
  XOR U30061 ( .A(n29899), .B(n29897), .Z(n29902) );
  XOR U30062 ( .A(n29900), .B(n29902), .Z(n29767) );
  XOR U30063 ( .A(n29765), .B(n29767), .Z(n29768) );
  XOR U30064 ( .A(n29769), .B(n29768), .Z(n29734) );
  IV U30065 ( .A(n29734), .Z(n29760) );
  NOR U30066 ( .A(n29736), .B(n29735), .Z(n29741) );
  IV U30067 ( .A(n29737), .Z(n29738) );
  NOR U30068 ( .A(n29739), .B(n29738), .Z(n29740) );
  NOR U30069 ( .A(n29741), .B(n29740), .Z(n29759) );
  NOR U30070 ( .A(n167), .B(n129), .Z(n29757) );
  XOR U30071 ( .A(n29759), .B(n29757), .Z(n29761) );
  XOR U30072 ( .A(n29760), .B(n29761), .Z(n30076) );
  XOR U30073 ( .A(n30074), .B(n30076), .Z(n30065) );
  NOR U30074 ( .A(n29743), .B(n29742), .Z(n30067) );
  IV U30075 ( .A(n30067), .Z(n29744) );
  NOR U30076 ( .A(n29744), .B(n29748), .Z(n29745) );
  IV U30077 ( .A(n29745), .Z(n29746) );
  NOR U30078 ( .A(n29752), .B(n29746), .Z(n29914) );
  NOR U30079 ( .A(n29747), .B(n29750), .Z(n29749) );
  NOR U30080 ( .A(n29749), .B(n29748), .Z(n30068) );
  IV U30081 ( .A(n29750), .Z(n29751) );
  NOR U30082 ( .A(n29752), .B(n29751), .Z(n29753) );
  NOR U30083 ( .A(n30067), .B(n29753), .Z(n30077) );
  IV U30084 ( .A(n30077), .Z(n29754) );
  NOR U30085 ( .A(n30068), .B(n29754), .Z(n29755) );
  NOR U30086 ( .A(n29914), .B(n29755), .Z(n29756) );
  IV U30087 ( .A(n29756), .Z(n29906) );
  XOR U30088 ( .A(n30065), .B(n29906), .Z(c[107]) );
  IV U30089 ( .A(n29757), .Z(n29758) );
  NOR U30090 ( .A(n29759), .B(n29758), .Z(n29763) );
  NOR U30091 ( .A(n29761), .B(n29760), .Z(n29762) );
  NOR U30092 ( .A(n29763), .B(n29762), .Z(n30058) );
  NOR U30093 ( .A(n167), .B(n130), .Z(n29764) );
  IV U30094 ( .A(n29764), .Z(n29922) );
  IV U30095 ( .A(n29765), .Z(n29766) );
  NOR U30096 ( .A(n29767), .B(n29766), .Z(n29771) );
  NOR U30097 ( .A(n29769), .B(n29768), .Z(n29770) );
  NOR U30098 ( .A(n29771), .B(n29770), .Z(n29920) );
  NOR U30099 ( .A(n161), .B(n136), .Z(n29772) );
  IV U30100 ( .A(n29772), .Z(n29937) );
  IV U30101 ( .A(n29773), .Z(n29774) );
  NOR U30102 ( .A(n29775), .B(n29774), .Z(n29780) );
  IV U30103 ( .A(n29776), .Z(n29777) );
  NOR U30104 ( .A(n29778), .B(n29777), .Z(n29779) );
  NOR U30105 ( .A(n29780), .B(n29779), .Z(n29935) );
  NOR U30106 ( .A(n155), .B(n142), .Z(n29952) );
  IV U30107 ( .A(n29781), .Z(n29782) );
  NOR U30108 ( .A(n29783), .B(n29782), .Z(n29787) );
  NOR U30109 ( .A(n29785), .B(n29784), .Z(n29786) );
  NOR U30110 ( .A(n29787), .B(n29786), .Z(n29951) );
  NOR U30111 ( .A(n150), .B(n146), .Z(n29788) );
  IV U30112 ( .A(n29788), .Z(n29967) );
  IV U30113 ( .A(n29789), .Z(n29790) );
  NOR U30114 ( .A(n29791), .B(n29790), .Z(n29795) );
  NOR U30115 ( .A(n29793), .B(n29792), .Z(n29794) );
  NOR U30116 ( .A(n29795), .B(n29794), .Z(n29965) );
  NOR U30117 ( .A(n145), .B(n152), .Z(n29980) );
  IV U30118 ( .A(n29796), .Z(n29797) );
  NOR U30119 ( .A(n29798), .B(n29797), .Z(n29803) );
  IV U30120 ( .A(n29799), .Z(n29801) );
  NOR U30121 ( .A(n29801), .B(n29800), .Z(n29802) );
  NOR U30122 ( .A(n29803), .B(n29802), .Z(n29979) );
  NOR U30123 ( .A(n139), .B(n159), .Z(n29996) );
  IV U30124 ( .A(n29804), .Z(n29805) );
  NOR U30125 ( .A(n29806), .B(n29805), .Z(n29811) );
  IV U30126 ( .A(n29807), .Z(n29808) );
  NOR U30127 ( .A(n29809), .B(n29808), .Z(n29810) );
  NOR U30128 ( .A(n29811), .B(n29810), .Z(n30000) );
  NOR U30129 ( .A(n135), .B(n162), .Z(n29812) );
  IV U30130 ( .A(n29812), .Z(n30008) );
  IV U30131 ( .A(n29813), .Z(n29814) );
  NOR U30132 ( .A(n29815), .B(n29814), .Z(n29819) );
  NOR U30133 ( .A(n29817), .B(n29816), .Z(n29818) );
  NOR U30134 ( .A(n29819), .B(n29818), .Z(n30006) );
  NOR U30135 ( .A(n164), .B(n133), .Z(n30015) );
  IV U30136 ( .A(n29820), .Z(n29821) );
  NOR U30137 ( .A(n29822), .B(n29821), .Z(n29827) );
  IV U30138 ( .A(n29823), .Z(n29824) );
  NOR U30139 ( .A(n29825), .B(n29824), .Z(n29826) );
  NOR U30140 ( .A(n29827), .B(n29826), .Z(n30014) );
  NOR U30141 ( .A(n166), .B(n131), .Z(n30012) );
  XOR U30142 ( .A(n30014), .B(n30012), .Z(n30017) );
  XOR U30143 ( .A(n30015), .B(n30017), .Z(n30005) );
  XOR U30144 ( .A(n30006), .B(n30005), .Z(n30007) );
  XOR U30145 ( .A(n30008), .B(n30007), .Z(n29999) );
  XOR U30146 ( .A(n30000), .B(n29999), .Z(n29828) );
  IV U30147 ( .A(n29828), .Z(n30002) );
  NOR U30148 ( .A(n137), .B(n160), .Z(n29829) );
  IV U30149 ( .A(n29829), .Z(n30001) );
  XOR U30150 ( .A(n30002), .B(n30001), .Z(n29994) );
  IV U30151 ( .A(n29830), .Z(n29831) );
  NOR U30152 ( .A(n29832), .B(n29831), .Z(n29836) );
  NOR U30153 ( .A(n29834), .B(n29833), .Z(n29835) );
  NOR U30154 ( .A(n29836), .B(n29835), .Z(n29992) );
  XOR U30155 ( .A(n29994), .B(n29992), .Z(n29995) );
  XOR U30156 ( .A(n29996), .B(n29995), .Z(n29989) );
  IV U30157 ( .A(n29837), .Z(n29838) );
  NOR U30158 ( .A(n29839), .B(n29838), .Z(n29844) );
  IV U30159 ( .A(n29840), .Z(n29841) );
  NOR U30160 ( .A(n29842), .B(n29841), .Z(n29843) );
  NOR U30161 ( .A(n29844), .B(n29843), .Z(n29987) );
  NOR U30162 ( .A(n141), .B(n157), .Z(n29985) );
  XOR U30163 ( .A(n29987), .B(n29985), .Z(n29988) );
  XOR U30164 ( .A(n29989), .B(n29988), .Z(n30026) );
  IV U30165 ( .A(n29845), .Z(n29846) );
  NOR U30166 ( .A(n29847), .B(n29846), .Z(n29851) );
  NOR U30167 ( .A(n29849), .B(n29848), .Z(n29850) );
  NOR U30168 ( .A(n29851), .B(n29850), .Z(n30025) );
  NOR U30169 ( .A(n143), .B(n154), .Z(n30023) );
  XOR U30170 ( .A(n30025), .B(n30023), .Z(n30027) );
  XOR U30171 ( .A(n30026), .B(n30027), .Z(n29978) );
  XOR U30172 ( .A(n29979), .B(n29978), .Z(n29852) );
  IV U30173 ( .A(n29852), .Z(n29982) );
  XOR U30174 ( .A(n29980), .B(n29982), .Z(n29974) );
  NOR U30175 ( .A(n29854), .B(n29853), .Z(n29859) );
  IV U30176 ( .A(n29855), .Z(n29856) );
  NOR U30177 ( .A(n29857), .B(n29856), .Z(n29858) );
  NOR U30178 ( .A(n29859), .B(n29858), .Z(n29973) );
  NOR U30179 ( .A(n147), .B(n151), .Z(n29971) );
  XOR U30180 ( .A(n29973), .B(n29971), .Z(n29975) );
  XOR U30181 ( .A(n29974), .B(n29975), .Z(n30035) );
  NOR U30182 ( .A(n29861), .B(n29860), .Z(n29866) );
  IV U30183 ( .A(n29862), .Z(n29863) );
  NOR U30184 ( .A(n29864), .B(n29863), .Z(n29865) );
  NOR U30185 ( .A(n29866), .B(n29865), .Z(n30034) );
  NOR U30186 ( .A(n148), .B(n149), .Z(n30032) );
  XOR U30187 ( .A(n30034), .B(n30032), .Z(n30037) );
  XOR U30188 ( .A(n30035), .B(n30037), .Z(n29964) );
  XOR U30189 ( .A(n29965), .B(n29964), .Z(n29966) );
  XOR U30190 ( .A(n29967), .B(n29966), .Z(n29961) );
  IV U30191 ( .A(n29867), .Z(n29868) );
  NOR U30192 ( .A(n29869), .B(n29868), .Z(n29874) );
  IV U30193 ( .A(n29870), .Z(n29871) );
  NOR U30194 ( .A(n29872), .B(n29871), .Z(n29873) );
  NOR U30195 ( .A(n29874), .B(n29873), .Z(n29959) );
  NOR U30196 ( .A(n153), .B(n144), .Z(n29957) );
  XOR U30197 ( .A(n29959), .B(n29957), .Z(n29960) );
  XOR U30198 ( .A(n29961), .B(n29960), .Z(n29949) );
  XOR U30199 ( .A(n29951), .B(n29949), .Z(n29954) );
  XOR U30200 ( .A(n29952), .B(n29954), .Z(n30044) );
  IV U30201 ( .A(n29875), .Z(n29876) );
  NOR U30202 ( .A(n29877), .B(n29876), .Z(n29882) );
  IV U30203 ( .A(n29878), .Z(n29879) );
  NOR U30204 ( .A(n29880), .B(n29879), .Z(n29881) );
  NOR U30205 ( .A(n29882), .B(n29881), .Z(n30043) );
  NOR U30206 ( .A(n156), .B(n140), .Z(n30041) );
  XOR U30207 ( .A(n30043), .B(n30041), .Z(n30045) );
  XOR U30208 ( .A(n30044), .B(n30045), .Z(n29944) );
  IV U30209 ( .A(n29883), .Z(n29884) );
  NOR U30210 ( .A(n29885), .B(n29884), .Z(n29889) );
  NOR U30211 ( .A(n29887), .B(n29886), .Z(n29888) );
  NOR U30212 ( .A(n29889), .B(n29888), .Z(n29943) );
  NOR U30213 ( .A(n158), .B(n138), .Z(n29941) );
  XOR U30214 ( .A(n29943), .B(n29941), .Z(n29945) );
  XOR U30215 ( .A(n29944), .B(n29945), .Z(n29934) );
  XOR U30216 ( .A(n29935), .B(n29934), .Z(n29936) );
  XOR U30217 ( .A(n29937), .B(n29936), .Z(n30052) );
  IV U30218 ( .A(n29890), .Z(n29891) );
  NOR U30219 ( .A(n29892), .B(n29891), .Z(n29896) );
  NOR U30220 ( .A(n29894), .B(n29893), .Z(n29895) );
  NOR U30221 ( .A(n29896), .B(n29895), .Z(n30051) );
  NOR U30222 ( .A(n163), .B(n134), .Z(n30049) );
  XOR U30223 ( .A(n30051), .B(n30049), .Z(n30053) );
  XOR U30224 ( .A(n30052), .B(n30053), .Z(n29929) );
  IV U30225 ( .A(n29897), .Z(n29898) );
  NOR U30226 ( .A(n29899), .B(n29898), .Z(n29904) );
  IV U30227 ( .A(n29900), .Z(n29901) );
  NOR U30228 ( .A(n29902), .B(n29901), .Z(n29903) );
  NOR U30229 ( .A(n29904), .B(n29903), .Z(n29928) );
  NOR U30230 ( .A(n165), .B(n132), .Z(n29926) );
  XOR U30231 ( .A(n29928), .B(n29926), .Z(n29931) );
  XOR U30232 ( .A(n29929), .B(n29931), .Z(n29919) );
  XOR U30233 ( .A(n29920), .B(n29919), .Z(n29921) );
  XOR U30234 ( .A(n29922), .B(n29921), .Z(n30057) );
  XOR U30235 ( .A(n30058), .B(n30057), .Z(n29911) );
  IV U30236 ( .A(n29911), .Z(n30081) );
  IV U30237 ( .A(n30076), .Z(n29905) );
  NOR U30238 ( .A(n30074), .B(n29905), .Z(n30080) );
  XOR U30239 ( .A(n30080), .B(n29914), .Z(n29909) );
  NOR U30240 ( .A(n30065), .B(n29906), .Z(n29913) );
  IV U30241 ( .A(n29913), .Z(n29907) );
  NOR U30242 ( .A(n29914), .B(n29907), .Z(n29908) );
  NOR U30243 ( .A(n29909), .B(n29908), .Z(n29910) );
  XOR U30244 ( .A(n30081), .B(n29910), .Z(c[108]) );
  NOR U30245 ( .A(n30080), .B(n29911), .Z(n30070) );
  IV U30246 ( .A(n30080), .Z(n29912) );
  NOR U30247 ( .A(n30081), .B(n29912), .Z(n29917) );
  NOR U30248 ( .A(n29914), .B(n29913), .Z(n29915) );
  IV U30249 ( .A(n29915), .Z(n29916) );
  NOR U30250 ( .A(n29917), .B(n29916), .Z(n29918) );
  NOR U30251 ( .A(n30070), .B(n29918), .Z(n30060) );
  NOR U30252 ( .A(n29920), .B(n29919), .Z(n29925) );
  IV U30253 ( .A(n29921), .Z(n29923) );
  NOR U30254 ( .A(n29923), .B(n29922), .Z(n29924) );
  NOR U30255 ( .A(n29925), .B(n29924), .Z(n30090) );
  NOR U30256 ( .A(n167), .B(n132), .Z(n30093) );
  IV U30257 ( .A(n29926), .Z(n29927) );
  NOR U30258 ( .A(n29928), .B(n29927), .Z(n29933) );
  IV U30259 ( .A(n29929), .Z(n29930) );
  NOR U30260 ( .A(n29931), .B(n29930), .Z(n29932) );
  NOR U30261 ( .A(n29933), .B(n29932), .Z(n30092) );
  NOR U30262 ( .A(n29935), .B(n29934), .Z(n29940) );
  IV U30263 ( .A(n29936), .Z(n29938) );
  NOR U30264 ( .A(n29938), .B(n29937), .Z(n29939) );
  NOR U30265 ( .A(n29940), .B(n29939), .Z(n30218) );
  NOR U30266 ( .A(n163), .B(n136), .Z(n30214) );
  NOR U30267 ( .A(n161), .B(n138), .Z(n30209) );
  IV U30268 ( .A(n29941), .Z(n29942) );
  NOR U30269 ( .A(n29943), .B(n29942), .Z(n29948) );
  IV U30270 ( .A(n29944), .Z(n29946) );
  NOR U30271 ( .A(n29946), .B(n29945), .Z(n29947) );
  NOR U30272 ( .A(n29948), .B(n29947), .Z(n30208) );
  IV U30273 ( .A(n29949), .Z(n29950) );
  NOR U30274 ( .A(n29951), .B(n29950), .Z(n29956) );
  IV U30275 ( .A(n29952), .Z(n29953) );
  NOR U30276 ( .A(n29954), .B(n29953), .Z(n29955) );
  NOR U30277 ( .A(n29956), .B(n29955), .Z(n30204) );
  NOR U30278 ( .A(n156), .B(n142), .Z(n30200) );
  NOR U30279 ( .A(n155), .B(n144), .Z(n30195) );
  IV U30280 ( .A(n29957), .Z(n29958) );
  NOR U30281 ( .A(n29959), .B(n29958), .Z(n29963) );
  NOR U30282 ( .A(n29961), .B(n29960), .Z(n29962) );
  NOR U30283 ( .A(n29963), .B(n29962), .Z(n30194) );
  IV U30284 ( .A(n30194), .Z(n30040) );
  NOR U30285 ( .A(n153), .B(n146), .Z(n30118) );
  NOR U30286 ( .A(n29965), .B(n29964), .Z(n29970) );
  IV U30287 ( .A(n29966), .Z(n29968) );
  NOR U30288 ( .A(n29968), .B(n29967), .Z(n29969) );
  NOR U30289 ( .A(n29970), .B(n29969), .Z(n30117) );
  NOR U30290 ( .A(n148), .B(n151), .Z(n30133) );
  IV U30291 ( .A(n29971), .Z(n29972) );
  NOR U30292 ( .A(n29973), .B(n29972), .Z(n29977) );
  NOR U30293 ( .A(n29975), .B(n29974), .Z(n29976) );
  NOR U30294 ( .A(n29977), .B(n29976), .Z(n30132) );
  NOR U30295 ( .A(n29979), .B(n29978), .Z(n29984) );
  IV U30296 ( .A(n29980), .Z(n29981) );
  NOR U30297 ( .A(n29982), .B(n29981), .Z(n29983) );
  NOR U30298 ( .A(n29984), .B(n29983), .Z(n30142) );
  NOR U30299 ( .A(n147), .B(n152), .Z(n30138) );
  NOR U30300 ( .A(n143), .B(n157), .Z(n30179) );
  IV U30301 ( .A(n29985), .Z(n29986) );
  NOR U30302 ( .A(n29987), .B(n29986), .Z(n29991) );
  NOR U30303 ( .A(n29989), .B(n29988), .Z(n29990) );
  NOR U30304 ( .A(n29991), .B(n29990), .Z(n30178) );
  IV U30305 ( .A(n30178), .Z(n30022) );
  NOR U30306 ( .A(n141), .B(n159), .Z(n30148) );
  IV U30307 ( .A(n29992), .Z(n29993) );
  NOR U30308 ( .A(n29994), .B(n29993), .Z(n29998) );
  NOR U30309 ( .A(n29996), .B(n29995), .Z(n29997) );
  NOR U30310 ( .A(n29998), .B(n29997), .Z(n30145) );
  NOR U30311 ( .A(n139), .B(n160), .Z(n30171) );
  NOR U30312 ( .A(n30000), .B(n29999), .Z(n30004) );
  NOR U30313 ( .A(n30002), .B(n30001), .Z(n30003) );
  NOR U30314 ( .A(n30004), .B(n30003), .Z(n30170) );
  IV U30315 ( .A(n30170), .Z(n30021) );
  NOR U30316 ( .A(n137), .B(n162), .Z(n30155) );
  NOR U30317 ( .A(n30006), .B(n30005), .Z(n30011) );
  IV U30318 ( .A(n30007), .Z(n30009) );
  NOR U30319 ( .A(n30009), .B(n30008), .Z(n30010) );
  NOR U30320 ( .A(n30011), .B(n30010), .Z(n30154) );
  IV U30321 ( .A(n30154), .Z(n30020) );
  NOR U30322 ( .A(n164), .B(n135), .Z(n30163) );
  IV U30323 ( .A(n30012), .Z(n30013) );
  NOR U30324 ( .A(n30014), .B(n30013), .Z(n30019) );
  IV U30325 ( .A(n30015), .Z(n30016) );
  NOR U30326 ( .A(n30017), .B(n30016), .Z(n30018) );
  NOR U30327 ( .A(n30019), .B(n30018), .Z(n30162) );
  NOR U30328 ( .A(n166), .B(n133), .Z(n30160) );
  XOR U30329 ( .A(n30162), .B(n30160), .Z(n30165) );
  XOR U30330 ( .A(n30163), .B(n30165), .Z(n30153) );
  XOR U30331 ( .A(n30020), .B(n30153), .Z(n30157) );
  XOR U30332 ( .A(n30155), .B(n30157), .Z(n30169) );
  XOR U30333 ( .A(n30021), .B(n30169), .Z(n30173) );
  XOR U30334 ( .A(n30171), .B(n30173), .Z(n30147) );
  XOR U30335 ( .A(n30145), .B(n30147), .Z(n30150) );
  XOR U30336 ( .A(n30148), .B(n30150), .Z(n30177) );
  XOR U30337 ( .A(n30022), .B(n30177), .Z(n30181) );
  XOR U30338 ( .A(n30179), .B(n30181), .Z(n30187) );
  IV U30339 ( .A(n30187), .Z(n30031) );
  IV U30340 ( .A(n30023), .Z(n30024) );
  NOR U30341 ( .A(n30025), .B(n30024), .Z(n30030) );
  IV U30342 ( .A(n30026), .Z(n30028) );
  NOR U30343 ( .A(n30028), .B(n30027), .Z(n30029) );
  NOR U30344 ( .A(n30030), .B(n30029), .Z(n30186) );
  NOR U30345 ( .A(n145), .B(n154), .Z(n30184) );
  XOR U30346 ( .A(n30186), .B(n30184), .Z(n30188) );
  XOR U30347 ( .A(n30031), .B(n30188), .Z(n30140) );
  XOR U30348 ( .A(n30138), .B(n30140), .Z(n30141) );
  XOR U30349 ( .A(n30142), .B(n30141), .Z(n30130) );
  XOR U30350 ( .A(n30132), .B(n30130), .Z(n30135) );
  XOR U30351 ( .A(n30133), .B(n30135), .Z(n30126) );
  IV U30352 ( .A(n30032), .Z(n30033) );
  NOR U30353 ( .A(n30034), .B(n30033), .Z(n30039) );
  IV U30354 ( .A(n30035), .Z(n30036) );
  NOR U30355 ( .A(n30037), .B(n30036), .Z(n30038) );
  NOR U30356 ( .A(n30039), .B(n30038), .Z(n30125) );
  NOR U30357 ( .A(n150), .B(n149), .Z(n30123) );
  XOR U30358 ( .A(n30125), .B(n30123), .Z(n30127) );
  XOR U30359 ( .A(n30126), .B(n30127), .Z(n30115) );
  XOR U30360 ( .A(n30117), .B(n30115), .Z(n30120) );
  XOR U30361 ( .A(n30118), .B(n30120), .Z(n30193) );
  XOR U30362 ( .A(n30040), .B(n30193), .Z(n30197) );
  XOR U30363 ( .A(n30195), .B(n30197), .Z(n30202) );
  XOR U30364 ( .A(n30200), .B(n30202), .Z(n30203) );
  XOR U30365 ( .A(n30204), .B(n30203), .Z(n30110) );
  IV U30366 ( .A(n30041), .Z(n30042) );
  NOR U30367 ( .A(n30043), .B(n30042), .Z(n30047) );
  NOR U30368 ( .A(n30045), .B(n30044), .Z(n30046) );
  NOR U30369 ( .A(n30047), .B(n30046), .Z(n30109) );
  NOR U30370 ( .A(n158), .B(n140), .Z(n30107) );
  XOR U30371 ( .A(n30109), .B(n30107), .Z(n30111) );
  XOR U30372 ( .A(n30110), .B(n30111), .Z(n30207) );
  XOR U30373 ( .A(n30208), .B(n30207), .Z(n30048) );
  IV U30374 ( .A(n30048), .Z(n30211) );
  XOR U30375 ( .A(n30209), .B(n30211), .Z(n30216) );
  XOR U30376 ( .A(n30214), .B(n30216), .Z(n30217) );
  XOR U30377 ( .A(n30218), .B(n30217), .Z(n30102) );
  IV U30378 ( .A(n30049), .Z(n30050) );
  NOR U30379 ( .A(n30051), .B(n30050), .Z(n30055) );
  NOR U30380 ( .A(n30053), .B(n30052), .Z(n30054) );
  NOR U30381 ( .A(n30055), .B(n30054), .Z(n30101) );
  NOR U30382 ( .A(n165), .B(n134), .Z(n30099) );
  XOR U30383 ( .A(n30101), .B(n30099), .Z(n30104) );
  XOR U30384 ( .A(n30102), .B(n30104), .Z(n30091) );
  XOR U30385 ( .A(n30092), .B(n30091), .Z(n30056) );
  IV U30386 ( .A(n30056), .Z(n30095) );
  XOR U30387 ( .A(n30093), .B(n30095), .Z(n30089) );
  XOR U30388 ( .A(n30090), .B(n30089), .Z(n30063) );
  IV U30389 ( .A(n30063), .Z(n30061) );
  NOR U30390 ( .A(n30058), .B(n30057), .Z(n30064) );
  IV U30391 ( .A(n30064), .Z(n30062) );
  XOR U30392 ( .A(n30061), .B(n30062), .Z(n30059) );
  XOR U30393 ( .A(n30060), .B(n30059), .Z(c[109]) );
  NOR U30394 ( .A(n30062), .B(n30061), .Z(n30088) );
  NOR U30395 ( .A(n30064), .B(n30063), .Z(n30086) );
  IV U30396 ( .A(n30065), .Z(n30066) );
  NOR U30397 ( .A(n30067), .B(n30066), .Z(n30073) );
  IV U30398 ( .A(n30068), .Z(n30069) );
  NOR U30399 ( .A(n30070), .B(n30069), .Z(n30071) );
  IV U30400 ( .A(n30071), .Z(n30072) );
  NOR U30401 ( .A(n30073), .B(n30072), .Z(n30084) );
  IV U30402 ( .A(n30074), .Z(n30075) );
  NOR U30403 ( .A(n30076), .B(n30075), .Z(n30078) );
  NOR U30404 ( .A(n30078), .B(n30077), .Z(n30079) );
  NOR U30405 ( .A(n30080), .B(n30079), .Z(n30082) );
  NOR U30406 ( .A(n30082), .B(n30081), .Z(n30083) );
  NOR U30407 ( .A(n30084), .B(n30083), .Z(n30085) );
  NOR U30408 ( .A(n30086), .B(n30085), .Z(n30087) );
  NOR U30409 ( .A(n30088), .B(n30087), .Z(n30226) );
  NOR U30410 ( .A(n30090), .B(n30089), .Z(n30222) );
  NOR U30411 ( .A(n30092), .B(n30091), .Z(n30097) );
  IV U30412 ( .A(n30093), .Z(n30094) );
  NOR U30413 ( .A(n30095), .B(n30094), .Z(n30096) );
  NOR U30414 ( .A(n30097), .B(n30096), .Z(n30231) );
  IV U30415 ( .A(n30231), .Z(n30221) );
  NOR U30416 ( .A(n167), .B(n134), .Z(n30098) );
  IV U30417 ( .A(n30098), .Z(n30235) );
  IV U30418 ( .A(n30099), .Z(n30100) );
  NOR U30419 ( .A(n30101), .B(n30100), .Z(n30106) );
  IV U30420 ( .A(n30102), .Z(n30103) );
  NOR U30421 ( .A(n30104), .B(n30103), .Z(n30105) );
  NOR U30422 ( .A(n30106), .B(n30105), .Z(n30233) );
  NOR U30423 ( .A(n161), .B(n140), .Z(n30344) );
  IV U30424 ( .A(n30107), .Z(n30108) );
  NOR U30425 ( .A(n30109), .B(n30108), .Z(n30114) );
  IV U30426 ( .A(n30110), .Z(n30112) );
  NOR U30427 ( .A(n30112), .B(n30111), .Z(n30113) );
  NOR U30428 ( .A(n30114), .B(n30113), .Z(n30343) );
  IV U30429 ( .A(n30115), .Z(n30116) );
  NOR U30430 ( .A(n30117), .B(n30116), .Z(n30122) );
  IV U30431 ( .A(n30118), .Z(n30119) );
  NOR U30432 ( .A(n30120), .B(n30119), .Z(n30121) );
  NOR U30433 ( .A(n30122), .B(n30121), .Z(n30259) );
  NOR U30434 ( .A(n155), .B(n146), .Z(n30255) );
  NOR U30435 ( .A(n153), .B(n149), .Z(n30327) );
  IV U30436 ( .A(n30123), .Z(n30124) );
  NOR U30437 ( .A(n30125), .B(n30124), .Z(n30129) );
  NOR U30438 ( .A(n30127), .B(n30126), .Z(n30128) );
  NOR U30439 ( .A(n30129), .B(n30128), .Z(n30326) );
  IV U30440 ( .A(n30326), .Z(n30192) );
  NOR U30441 ( .A(n150), .B(n151), .Z(n30264) );
  IV U30442 ( .A(n30130), .Z(n30131) );
  NOR U30443 ( .A(n30132), .B(n30131), .Z(n30137) );
  IV U30444 ( .A(n30133), .Z(n30134) );
  NOR U30445 ( .A(n30135), .B(n30134), .Z(n30136) );
  NOR U30446 ( .A(n30137), .B(n30136), .Z(n30263) );
  IV U30447 ( .A(n30263), .Z(n30191) );
  NOR U30448 ( .A(n148), .B(n152), .Z(n30272) );
  IV U30449 ( .A(n30138), .Z(n30139) );
  NOR U30450 ( .A(n30140), .B(n30139), .Z(n30144) );
  NOR U30451 ( .A(n30142), .B(n30141), .Z(n30143) );
  NOR U30452 ( .A(n30144), .B(n30143), .Z(n30271) );
  IV U30453 ( .A(n30145), .Z(n30146) );
  NOR U30454 ( .A(n30147), .B(n30146), .Z(n30152) );
  IV U30455 ( .A(n30148), .Z(n30149) );
  NOR U30456 ( .A(n30150), .B(n30149), .Z(n30151) );
  NOR U30457 ( .A(n30152), .B(n30151), .Z(n30312) );
  NOR U30458 ( .A(n143), .B(n159), .Z(n30308) );
  NOR U30459 ( .A(n139), .B(n162), .Z(n30293) );
  NOR U30460 ( .A(n30154), .B(n30153), .Z(n30159) );
  IV U30461 ( .A(n30155), .Z(n30156) );
  NOR U30462 ( .A(n30157), .B(n30156), .Z(n30158) );
  NOR U30463 ( .A(n30159), .B(n30158), .Z(n30292) );
  IV U30464 ( .A(n30292), .Z(n30168) );
  NOR U30465 ( .A(n164), .B(n137), .Z(n30301) );
  IV U30466 ( .A(n30160), .Z(n30161) );
  NOR U30467 ( .A(n30162), .B(n30161), .Z(n30167) );
  IV U30468 ( .A(n30163), .Z(n30164) );
  NOR U30469 ( .A(n30165), .B(n30164), .Z(n30166) );
  NOR U30470 ( .A(n30167), .B(n30166), .Z(n30300) );
  NOR U30471 ( .A(n166), .B(n135), .Z(n30298) );
  XOR U30472 ( .A(n30300), .B(n30298), .Z(n30303) );
  XOR U30473 ( .A(n30301), .B(n30303), .Z(n30291) );
  XOR U30474 ( .A(n30168), .B(n30291), .Z(n30295) );
  XOR U30475 ( .A(n30293), .B(n30295), .Z(n30287) );
  NOR U30476 ( .A(n30170), .B(n30169), .Z(n30175) );
  IV U30477 ( .A(n30171), .Z(n30172) );
  NOR U30478 ( .A(n30173), .B(n30172), .Z(n30174) );
  NOR U30479 ( .A(n30175), .B(n30174), .Z(n30286) );
  NOR U30480 ( .A(n141), .B(n160), .Z(n30284) );
  XOR U30481 ( .A(n30286), .B(n30284), .Z(n30288) );
  XOR U30482 ( .A(n30287), .B(n30288), .Z(n30176) );
  IV U30483 ( .A(n30176), .Z(n30310) );
  XOR U30484 ( .A(n30308), .B(n30310), .Z(n30311) );
  XOR U30485 ( .A(n30312), .B(n30311), .Z(n30281) );
  NOR U30486 ( .A(n145), .B(n157), .Z(n30279) );
  NOR U30487 ( .A(n30178), .B(n30177), .Z(n30183) );
  IV U30488 ( .A(n30179), .Z(n30180) );
  NOR U30489 ( .A(n30181), .B(n30180), .Z(n30182) );
  NOR U30490 ( .A(n30183), .B(n30182), .Z(n30277) );
  XOR U30491 ( .A(n30279), .B(n30277), .Z(n30280) );
  XOR U30492 ( .A(n30281), .B(n30280), .Z(n30320) );
  IV U30493 ( .A(n30184), .Z(n30185) );
  NOR U30494 ( .A(n30186), .B(n30185), .Z(n30190) );
  NOR U30495 ( .A(n30188), .B(n30187), .Z(n30189) );
  NOR U30496 ( .A(n30190), .B(n30189), .Z(n30318) );
  NOR U30497 ( .A(n147), .B(n154), .Z(n30316) );
  XOR U30498 ( .A(n30318), .B(n30316), .Z(n30319) );
  XOR U30499 ( .A(n30320), .B(n30319), .Z(n30269) );
  XOR U30500 ( .A(n30271), .B(n30269), .Z(n30274) );
  XOR U30501 ( .A(n30272), .B(n30274), .Z(n30262) );
  XOR U30502 ( .A(n30191), .B(n30262), .Z(n30266) );
  XOR U30503 ( .A(n30264), .B(n30266), .Z(n30325) );
  XOR U30504 ( .A(n30192), .B(n30325), .Z(n30329) );
  XOR U30505 ( .A(n30327), .B(n30329), .Z(n30257) );
  XOR U30506 ( .A(n30255), .B(n30257), .Z(n30258) );
  XOR U30507 ( .A(n30259), .B(n30258), .Z(n30336) );
  NOR U30508 ( .A(n30194), .B(n30193), .Z(n30199) );
  IV U30509 ( .A(n30195), .Z(n30196) );
  NOR U30510 ( .A(n30197), .B(n30196), .Z(n30198) );
  NOR U30511 ( .A(n30199), .B(n30198), .Z(n30335) );
  NOR U30512 ( .A(n156), .B(n144), .Z(n30333) );
  XOR U30513 ( .A(n30335), .B(n30333), .Z(n30338) );
  XOR U30514 ( .A(n30336), .B(n30338), .Z(n30251) );
  IV U30515 ( .A(n30200), .Z(n30201) );
  NOR U30516 ( .A(n30202), .B(n30201), .Z(n30206) );
  NOR U30517 ( .A(n30204), .B(n30203), .Z(n30205) );
  NOR U30518 ( .A(n30206), .B(n30205), .Z(n30250) );
  NOR U30519 ( .A(n158), .B(n142), .Z(n30248) );
  XOR U30520 ( .A(n30250), .B(n30248), .Z(n30252) );
  XOR U30521 ( .A(n30251), .B(n30252), .Z(n30341) );
  XOR U30522 ( .A(n30343), .B(n30341), .Z(n30346) );
  XOR U30523 ( .A(n30344), .B(n30346), .Z(n30352) );
  NOR U30524 ( .A(n30208), .B(n30207), .Z(n30213) );
  IV U30525 ( .A(n30209), .Z(n30210) );
  NOR U30526 ( .A(n30211), .B(n30210), .Z(n30212) );
  NOR U30527 ( .A(n30213), .B(n30212), .Z(n30351) );
  NOR U30528 ( .A(n163), .B(n138), .Z(n30349) );
  XOR U30529 ( .A(n30351), .B(n30349), .Z(n30353) );
  XOR U30530 ( .A(n30352), .B(n30353), .Z(n30243) );
  IV U30531 ( .A(n30214), .Z(n30215) );
  NOR U30532 ( .A(n30216), .B(n30215), .Z(n30220) );
  NOR U30533 ( .A(n30218), .B(n30217), .Z(n30219) );
  NOR U30534 ( .A(n30220), .B(n30219), .Z(n30242) );
  NOR U30535 ( .A(n165), .B(n136), .Z(n30240) );
  XOR U30536 ( .A(n30242), .B(n30240), .Z(n30244) );
  XOR U30537 ( .A(n30243), .B(n30244), .Z(n30232) );
  XOR U30538 ( .A(n30233), .B(n30232), .Z(n30234) );
  XOR U30539 ( .A(n30235), .B(n30234), .Z(n30230) );
  XOR U30540 ( .A(n30221), .B(n30230), .Z(n30224) );
  XOR U30541 ( .A(n30222), .B(n30224), .Z(n30225) );
  XOR U30542 ( .A(n30226), .B(n30225), .Z(c[110]) );
  IV U30543 ( .A(n30222), .Z(n30223) );
  NOR U30544 ( .A(n30224), .B(n30223), .Z(n30228) );
  NOR U30545 ( .A(n30226), .B(n30225), .Z(n30227) );
  NOR U30546 ( .A(n30228), .B(n30227), .Z(n30229) );
  IV U30547 ( .A(n30229), .Z(n30359) );
  NOR U30548 ( .A(n30231), .B(n30230), .Z(n30357) );
  NOR U30549 ( .A(n30233), .B(n30232), .Z(n30238) );
  IV U30550 ( .A(n30234), .Z(n30236) );
  NOR U30551 ( .A(n30236), .B(n30235), .Z(n30237) );
  NOR U30552 ( .A(n30238), .B(n30237), .Z(n30364) );
  NOR U30553 ( .A(n167), .B(n136), .Z(n30239) );
  IV U30554 ( .A(n30239), .Z(n30368) );
  IV U30555 ( .A(n30240), .Z(n30241) );
  NOR U30556 ( .A(n30242), .B(n30241), .Z(n30247) );
  IV U30557 ( .A(n30243), .Z(n30245) );
  NOR U30558 ( .A(n30245), .B(n30244), .Z(n30246) );
  NOR U30559 ( .A(n30247), .B(n30246), .Z(n30366) );
  NOR U30560 ( .A(n161), .B(n142), .Z(n30384) );
  IV U30561 ( .A(n30248), .Z(n30249) );
  NOR U30562 ( .A(n30250), .B(n30249), .Z(n30254) );
  NOR U30563 ( .A(n30252), .B(n30251), .Z(n30253) );
  NOR U30564 ( .A(n30254), .B(n30253), .Z(n30383) );
  NOR U30565 ( .A(n156), .B(n146), .Z(n30398) );
  IV U30566 ( .A(n30255), .Z(n30256) );
  NOR U30567 ( .A(n30257), .B(n30256), .Z(n30261) );
  NOR U30568 ( .A(n30259), .B(n30258), .Z(n30260) );
  NOR U30569 ( .A(n30261), .B(n30260), .Z(n30396) );
  IV U30570 ( .A(n30396), .Z(n30332) );
  NOR U30571 ( .A(n155), .B(n149), .Z(n30407) );
  NOR U30572 ( .A(n30263), .B(n30262), .Z(n30268) );
  IV U30573 ( .A(n30264), .Z(n30265) );
  NOR U30574 ( .A(n30266), .B(n30265), .Z(n30267) );
  NOR U30575 ( .A(n30268), .B(n30267), .Z(n30411) );
  NOR U30576 ( .A(n150), .B(n152), .Z(n30419) );
  IV U30577 ( .A(n30269), .Z(n30270) );
  NOR U30578 ( .A(n30271), .B(n30270), .Z(n30276) );
  IV U30579 ( .A(n30272), .Z(n30273) );
  NOR U30580 ( .A(n30274), .B(n30273), .Z(n30275) );
  NOR U30581 ( .A(n30276), .B(n30275), .Z(n30418) );
  NOR U30582 ( .A(n147), .B(n157), .Z(n30460) );
  IV U30583 ( .A(n30277), .Z(n30278) );
  NOR U30584 ( .A(n30279), .B(n30278), .Z(n30283) );
  NOR U30585 ( .A(n30281), .B(n30280), .Z(n30282) );
  NOR U30586 ( .A(n30283), .B(n30282), .Z(n30457) );
  NOR U30587 ( .A(n143), .B(n160), .Z(n30450) );
  IV U30588 ( .A(n30284), .Z(n30285) );
  NOR U30589 ( .A(n30286), .B(n30285), .Z(n30290) );
  NOR U30590 ( .A(n30288), .B(n30287), .Z(n30289) );
  NOR U30591 ( .A(n30290), .B(n30289), .Z(n30449) );
  IV U30592 ( .A(n30449), .Z(n30307) );
  NOR U30593 ( .A(n141), .B(n162), .Z(n30433) );
  NOR U30594 ( .A(n30292), .B(n30291), .Z(n30297) );
  IV U30595 ( .A(n30293), .Z(n30294) );
  NOR U30596 ( .A(n30295), .B(n30294), .Z(n30296) );
  NOR U30597 ( .A(n30297), .B(n30296), .Z(n30432) );
  IV U30598 ( .A(n30432), .Z(n30306) );
  NOR U30599 ( .A(n164), .B(n139), .Z(n30441) );
  IV U30600 ( .A(n30298), .Z(n30299) );
  NOR U30601 ( .A(n30300), .B(n30299), .Z(n30305) );
  IV U30602 ( .A(n30301), .Z(n30302) );
  NOR U30603 ( .A(n30303), .B(n30302), .Z(n30304) );
  NOR U30604 ( .A(n30305), .B(n30304), .Z(n30440) );
  NOR U30605 ( .A(n166), .B(n137), .Z(n30438) );
  XOR U30606 ( .A(n30440), .B(n30438), .Z(n30443) );
  XOR U30607 ( .A(n30441), .B(n30443), .Z(n30431) );
  XOR U30608 ( .A(n30306), .B(n30431), .Z(n30435) );
  XOR U30609 ( .A(n30433), .B(n30435), .Z(n30448) );
  XOR U30610 ( .A(n30307), .B(n30448), .Z(n30452) );
  XOR U30611 ( .A(n30450), .B(n30452), .Z(n30427) );
  IV U30612 ( .A(n30308), .Z(n30309) );
  NOR U30613 ( .A(n30310), .B(n30309), .Z(n30314) );
  NOR U30614 ( .A(n30312), .B(n30311), .Z(n30313) );
  NOR U30615 ( .A(n30314), .B(n30313), .Z(n30426) );
  NOR U30616 ( .A(n145), .B(n159), .Z(n30424) );
  XOR U30617 ( .A(n30426), .B(n30424), .Z(n30428) );
  XOR U30618 ( .A(n30427), .B(n30428), .Z(n30315) );
  IV U30619 ( .A(n30315), .Z(n30458) );
  XOR U30620 ( .A(n30457), .B(n30458), .Z(n30462) );
  XOR U30621 ( .A(n30460), .B(n30462), .Z(n30468) );
  IV U30622 ( .A(n30316), .Z(n30317) );
  NOR U30623 ( .A(n30318), .B(n30317), .Z(n30322) );
  NOR U30624 ( .A(n30320), .B(n30319), .Z(n30321) );
  NOR U30625 ( .A(n30322), .B(n30321), .Z(n30467) );
  NOR U30626 ( .A(n148), .B(n154), .Z(n30465) );
  XOR U30627 ( .A(n30467), .B(n30465), .Z(n30469) );
  XOR U30628 ( .A(n30468), .B(n30469), .Z(n30416) );
  XOR U30629 ( .A(n30418), .B(n30416), .Z(n30421) );
  XOR U30630 ( .A(n30419), .B(n30421), .Z(n30410) );
  XOR U30631 ( .A(n30411), .B(n30410), .Z(n30323) );
  IV U30632 ( .A(n30323), .Z(n30413) );
  NOR U30633 ( .A(n153), .B(n151), .Z(n30324) );
  IV U30634 ( .A(n30324), .Z(n30412) );
  XOR U30635 ( .A(n30413), .B(n30412), .Z(n30405) );
  NOR U30636 ( .A(n30326), .B(n30325), .Z(n30331) );
  IV U30637 ( .A(n30327), .Z(n30328) );
  NOR U30638 ( .A(n30329), .B(n30328), .Z(n30330) );
  NOR U30639 ( .A(n30331), .B(n30330), .Z(n30403) );
  XOR U30640 ( .A(n30405), .B(n30403), .Z(n30406) );
  XOR U30641 ( .A(n30407), .B(n30406), .Z(n30397) );
  XOR U30642 ( .A(n30332), .B(n30397), .Z(n30400) );
  XOR U30643 ( .A(n30398), .B(n30400), .Z(n30392) );
  IV U30644 ( .A(n30333), .Z(n30334) );
  NOR U30645 ( .A(n30335), .B(n30334), .Z(n30340) );
  IV U30646 ( .A(n30336), .Z(n30337) );
  NOR U30647 ( .A(n30338), .B(n30337), .Z(n30339) );
  NOR U30648 ( .A(n30340), .B(n30339), .Z(n30391) );
  NOR U30649 ( .A(n158), .B(n144), .Z(n30389) );
  XOR U30650 ( .A(n30391), .B(n30389), .Z(n30393) );
  XOR U30651 ( .A(n30392), .B(n30393), .Z(n30381) );
  XOR U30652 ( .A(n30383), .B(n30381), .Z(n30386) );
  XOR U30653 ( .A(n30384), .B(n30386), .Z(n30478) );
  IV U30654 ( .A(n30341), .Z(n30342) );
  NOR U30655 ( .A(n30343), .B(n30342), .Z(n30348) );
  IV U30656 ( .A(n30344), .Z(n30345) );
  NOR U30657 ( .A(n30346), .B(n30345), .Z(n30347) );
  NOR U30658 ( .A(n30348), .B(n30347), .Z(n30477) );
  NOR U30659 ( .A(n163), .B(n140), .Z(n30475) );
  XOR U30660 ( .A(n30477), .B(n30475), .Z(n30479) );
  XOR U30661 ( .A(n30478), .B(n30479), .Z(n30375) );
  IV U30662 ( .A(n30349), .Z(n30350) );
  NOR U30663 ( .A(n30351), .B(n30350), .Z(n30355) );
  NOR U30664 ( .A(n30353), .B(n30352), .Z(n30354) );
  NOR U30665 ( .A(n30355), .B(n30354), .Z(n30374) );
  NOR U30666 ( .A(n165), .B(n138), .Z(n30372) );
  XOR U30667 ( .A(n30374), .B(n30372), .Z(n30377) );
  XOR U30668 ( .A(n30375), .B(n30377), .Z(n30365) );
  XOR U30669 ( .A(n30366), .B(n30365), .Z(n30367) );
  XOR U30670 ( .A(n30368), .B(n30367), .Z(n30363) );
  XOR U30671 ( .A(n30364), .B(n30363), .Z(n30356) );
  XOR U30672 ( .A(n30357), .B(n30356), .Z(n30358) );
  XOR U30673 ( .A(n30359), .B(n30358), .Z(c[111]) );
  NOR U30674 ( .A(n30357), .B(n30356), .Z(n30362) );
  IV U30675 ( .A(n30358), .Z(n30360) );
  NOR U30676 ( .A(n30360), .B(n30359), .Z(n30361) );
  NOR U30677 ( .A(n30362), .B(n30361), .Z(n30593) );
  NOR U30678 ( .A(n30364), .B(n30363), .Z(n30590) );
  NOR U30679 ( .A(n30366), .B(n30365), .Z(n30371) );
  IV U30680 ( .A(n30367), .Z(n30369) );
  NOR U30681 ( .A(n30369), .B(n30368), .Z(n30370) );
  NOR U30682 ( .A(n30371), .B(n30370), .Z(n30483) );
  NOR U30683 ( .A(n167), .B(n138), .Z(n30487) );
  IV U30684 ( .A(n30372), .Z(n30373) );
  NOR U30685 ( .A(n30374), .B(n30373), .Z(n30379) );
  IV U30686 ( .A(n30375), .Z(n30376) );
  NOR U30687 ( .A(n30377), .B(n30376), .Z(n30378) );
  NOR U30688 ( .A(n30379), .B(n30378), .Z(n30486) );
  NOR U30689 ( .A(n163), .B(n142), .Z(n30380) );
  IV U30690 ( .A(n30380), .Z(n30584) );
  IV U30691 ( .A(n30381), .Z(n30382) );
  NOR U30692 ( .A(n30383), .B(n30382), .Z(n30388) );
  IV U30693 ( .A(n30384), .Z(n30385) );
  NOR U30694 ( .A(n30386), .B(n30385), .Z(n30387) );
  NOR U30695 ( .A(n30388), .B(n30387), .Z(n30582) );
  NOR U30696 ( .A(n161), .B(n144), .Z(n30576) );
  IV U30697 ( .A(n30389), .Z(n30390) );
  NOR U30698 ( .A(n30391), .B(n30390), .Z(n30395) );
  NOR U30699 ( .A(n30393), .B(n30392), .Z(n30394) );
  NOR U30700 ( .A(n30395), .B(n30394), .Z(n30575) );
  IV U30701 ( .A(n30575), .Z(n30474) );
  NOR U30702 ( .A(n158), .B(n146), .Z(n30501) );
  NOR U30703 ( .A(n30397), .B(n30396), .Z(n30402) );
  IV U30704 ( .A(n30398), .Z(n30399) );
  NOR U30705 ( .A(n30400), .B(n30399), .Z(n30401) );
  NOR U30706 ( .A(n30402), .B(n30401), .Z(n30500) );
  IV U30707 ( .A(n30500), .Z(n30473) );
  NOR U30708 ( .A(n156), .B(n149), .Z(n30569) );
  IV U30709 ( .A(n30403), .Z(n30404) );
  NOR U30710 ( .A(n30405), .B(n30404), .Z(n30409) );
  NOR U30711 ( .A(n30407), .B(n30406), .Z(n30408) );
  NOR U30712 ( .A(n30409), .B(n30408), .Z(n30566) );
  NOR U30713 ( .A(n155), .B(n151), .Z(n30561) );
  NOR U30714 ( .A(n30411), .B(n30410), .Z(n30415) );
  NOR U30715 ( .A(n30413), .B(n30412), .Z(n30414) );
  NOR U30716 ( .A(n30415), .B(n30414), .Z(n30560) );
  IV U30717 ( .A(n30560), .Z(n30472) );
  NOR U30718 ( .A(n153), .B(n152), .Z(n30510) );
  IV U30719 ( .A(n30416), .Z(n30417) );
  NOR U30720 ( .A(n30418), .B(n30417), .Z(n30423) );
  IV U30721 ( .A(n30419), .Z(n30420) );
  NOR U30722 ( .A(n30421), .B(n30420), .Z(n30422) );
  NOR U30723 ( .A(n30423), .B(n30422), .Z(n30509) );
  IV U30724 ( .A(n30424), .Z(n30425) );
  NOR U30725 ( .A(n30426), .B(n30425), .Z(n30430) );
  NOR U30726 ( .A(n30428), .B(n30427), .Z(n30429) );
  NOR U30727 ( .A(n30430), .B(n30429), .Z(n30530) );
  NOR U30728 ( .A(n145), .B(n160), .Z(n30540) );
  NOR U30729 ( .A(n30432), .B(n30431), .Z(n30437) );
  IV U30730 ( .A(n30433), .Z(n30434) );
  NOR U30731 ( .A(n30435), .B(n30434), .Z(n30436) );
  NOR U30732 ( .A(n30437), .B(n30436), .Z(n30544) );
  NOR U30733 ( .A(n164), .B(n141), .Z(n30552) );
  IV U30734 ( .A(n30438), .Z(n30439) );
  NOR U30735 ( .A(n30440), .B(n30439), .Z(n30445) );
  IV U30736 ( .A(n30441), .Z(n30442) );
  NOR U30737 ( .A(n30443), .B(n30442), .Z(n30444) );
  NOR U30738 ( .A(n30445), .B(n30444), .Z(n30551) );
  NOR U30739 ( .A(n166), .B(n139), .Z(n30549) );
  XOR U30740 ( .A(n30551), .B(n30549), .Z(n30554) );
  XOR U30741 ( .A(n30552), .B(n30554), .Z(n30543) );
  XOR U30742 ( .A(n30544), .B(n30543), .Z(n30446) );
  IV U30743 ( .A(n30446), .Z(n30546) );
  NOR U30744 ( .A(n143), .B(n162), .Z(n30447) );
  IV U30745 ( .A(n30447), .Z(n30545) );
  XOR U30746 ( .A(n30546), .B(n30545), .Z(n30538) );
  NOR U30747 ( .A(n30449), .B(n30448), .Z(n30454) );
  IV U30748 ( .A(n30450), .Z(n30451) );
  NOR U30749 ( .A(n30452), .B(n30451), .Z(n30453) );
  NOR U30750 ( .A(n30454), .B(n30453), .Z(n30536) );
  XOR U30751 ( .A(n30538), .B(n30536), .Z(n30539) );
  XOR U30752 ( .A(n30540), .B(n30539), .Z(n30531) );
  XOR U30753 ( .A(n30530), .B(n30531), .Z(n30455) );
  IV U30754 ( .A(n30455), .Z(n30533) );
  NOR U30755 ( .A(n147), .B(n159), .Z(n30456) );
  IV U30756 ( .A(n30456), .Z(n30532) );
  XOR U30757 ( .A(n30533), .B(n30532), .Z(n30526) );
  NOR U30758 ( .A(n148), .B(n157), .Z(n30524) );
  IV U30759 ( .A(n30457), .Z(n30459) );
  NOR U30760 ( .A(n30459), .B(n30458), .Z(n30464) );
  IV U30761 ( .A(n30460), .Z(n30461) );
  NOR U30762 ( .A(n30462), .B(n30461), .Z(n30463) );
  NOR U30763 ( .A(n30464), .B(n30463), .Z(n30522) );
  XOR U30764 ( .A(n30524), .B(n30522), .Z(n30525) );
  XOR U30765 ( .A(n30526), .B(n30525), .Z(n30519) );
  IV U30766 ( .A(n30465), .Z(n30466) );
  NOR U30767 ( .A(n30467), .B(n30466), .Z(n30471) );
  NOR U30768 ( .A(n30469), .B(n30468), .Z(n30470) );
  NOR U30769 ( .A(n30471), .B(n30470), .Z(n30517) );
  NOR U30770 ( .A(n150), .B(n154), .Z(n30515) );
  XOR U30771 ( .A(n30517), .B(n30515), .Z(n30518) );
  XOR U30772 ( .A(n30519), .B(n30518), .Z(n30507) );
  XOR U30773 ( .A(n30509), .B(n30507), .Z(n30512) );
  XOR U30774 ( .A(n30510), .B(n30512), .Z(n30559) );
  XOR U30775 ( .A(n30472), .B(n30559), .Z(n30563) );
  XOR U30776 ( .A(n30561), .B(n30563), .Z(n30567) );
  XOR U30777 ( .A(n30566), .B(n30567), .Z(n30571) );
  XOR U30778 ( .A(n30569), .B(n30571), .Z(n30499) );
  XOR U30779 ( .A(n30473), .B(n30499), .Z(n30503) );
  XOR U30780 ( .A(n30501), .B(n30503), .Z(n30574) );
  XOR U30781 ( .A(n30474), .B(n30574), .Z(n30578) );
  XOR U30782 ( .A(n30576), .B(n30578), .Z(n30581) );
  XOR U30783 ( .A(n30582), .B(n30581), .Z(n30583) );
  XOR U30784 ( .A(n30584), .B(n30583), .Z(n30495) );
  IV U30785 ( .A(n30475), .Z(n30476) );
  NOR U30786 ( .A(n30477), .B(n30476), .Z(n30481) );
  NOR U30787 ( .A(n30479), .B(n30478), .Z(n30480) );
  NOR U30788 ( .A(n30481), .B(n30480), .Z(n30494) );
  NOR U30789 ( .A(n165), .B(n140), .Z(n30492) );
  XOR U30790 ( .A(n30494), .B(n30492), .Z(n30496) );
  XOR U30791 ( .A(n30495), .B(n30496), .Z(n30484) );
  XOR U30792 ( .A(n30486), .B(n30484), .Z(n30489) );
  XOR U30793 ( .A(n30487), .B(n30489), .Z(n30482) );
  XOR U30794 ( .A(n30483), .B(n30482), .Z(n30589) );
  XOR U30795 ( .A(n30590), .B(n30589), .Z(n30591) );
  XOR U30796 ( .A(n30593), .B(n30591), .Z(c[112]) );
  NOR U30797 ( .A(n30483), .B(n30482), .Z(n30597) );
  IV U30798 ( .A(n30484), .Z(n30485) );
  NOR U30799 ( .A(n30486), .B(n30485), .Z(n30491) );
  IV U30800 ( .A(n30487), .Z(n30488) );
  NOR U30801 ( .A(n30489), .B(n30488), .Z(n30490) );
  NOR U30802 ( .A(n30491), .B(n30490), .Z(n30605) );
  IV U30803 ( .A(n30605), .Z(n30588) );
  NOR U30804 ( .A(n167), .B(n140), .Z(n30609) );
  IV U30805 ( .A(n30492), .Z(n30493) );
  NOR U30806 ( .A(n30494), .B(n30493), .Z(n30498) );
  NOR U30807 ( .A(n30496), .B(n30495), .Z(n30497) );
  NOR U30808 ( .A(n30498), .B(n30497), .Z(n30608) );
  NOR U30809 ( .A(n30500), .B(n30499), .Z(n30505) );
  IV U30810 ( .A(n30501), .Z(n30502) );
  NOR U30811 ( .A(n30503), .B(n30502), .Z(n30504) );
  NOR U30812 ( .A(n30505), .B(n30504), .Z(n30625) );
  NOR U30813 ( .A(n161), .B(n146), .Z(n30621) );
  NOR U30814 ( .A(n155), .B(n152), .Z(n30506) );
  IV U30815 ( .A(n30506), .Z(n30686) );
  IV U30816 ( .A(n30507), .Z(n30508) );
  NOR U30817 ( .A(n30509), .B(n30508), .Z(n30514) );
  IV U30818 ( .A(n30510), .Z(n30511) );
  NOR U30819 ( .A(n30512), .B(n30511), .Z(n30513) );
  NOR U30820 ( .A(n30514), .B(n30513), .Z(n30684) );
  NOR U30821 ( .A(n153), .B(n154), .Z(n30678) );
  IV U30822 ( .A(n30515), .Z(n30516) );
  NOR U30823 ( .A(n30517), .B(n30516), .Z(n30521) );
  NOR U30824 ( .A(n30519), .B(n30518), .Z(n30520) );
  NOR U30825 ( .A(n30521), .B(n30520), .Z(n30677) );
  IV U30826 ( .A(n30677), .Z(n30558) );
  IV U30827 ( .A(n30522), .Z(n30523) );
  NOR U30828 ( .A(n30524), .B(n30523), .Z(n30528) );
  NOR U30829 ( .A(n30526), .B(n30525), .Z(n30527) );
  NOR U30830 ( .A(n30528), .B(n30527), .Z(n30636) );
  NOR U30831 ( .A(n150), .B(n157), .Z(n30529) );
  IV U30832 ( .A(n30529), .Z(n30637) );
  XOR U30833 ( .A(n30636), .B(n30637), .Z(n30640) );
  NOR U30834 ( .A(n30531), .B(n30530), .Z(n30535) );
  NOR U30835 ( .A(n30533), .B(n30532), .Z(n30534) );
  NOR U30836 ( .A(n30535), .B(n30534), .Z(n30673) );
  NOR U30837 ( .A(n148), .B(n159), .Z(n30669) );
  IV U30838 ( .A(n30536), .Z(n30537) );
  NOR U30839 ( .A(n30538), .B(n30537), .Z(n30542) );
  NOR U30840 ( .A(n30540), .B(n30539), .Z(n30541) );
  NOR U30841 ( .A(n30542), .B(n30541), .Z(n30648) );
  NOR U30842 ( .A(n147), .B(n160), .Z(n30645) );
  NOR U30843 ( .A(n145), .B(n162), .Z(n30655) );
  NOR U30844 ( .A(n30544), .B(n30543), .Z(n30548) );
  NOR U30845 ( .A(n30546), .B(n30545), .Z(n30547) );
  NOR U30846 ( .A(n30548), .B(n30547), .Z(n30654) );
  IV U30847 ( .A(n30654), .Z(n30557) );
  NOR U30848 ( .A(n164), .B(n143), .Z(n30663) );
  IV U30849 ( .A(n30549), .Z(n30550) );
  NOR U30850 ( .A(n30551), .B(n30550), .Z(n30556) );
  IV U30851 ( .A(n30552), .Z(n30553) );
  NOR U30852 ( .A(n30554), .B(n30553), .Z(n30555) );
  NOR U30853 ( .A(n30556), .B(n30555), .Z(n30662) );
  NOR U30854 ( .A(n166), .B(n141), .Z(n30660) );
  XOR U30855 ( .A(n30662), .B(n30660), .Z(n30665) );
  XOR U30856 ( .A(n30663), .B(n30665), .Z(n30653) );
  XOR U30857 ( .A(n30557), .B(n30653), .Z(n30657) );
  XOR U30858 ( .A(n30655), .B(n30657), .Z(n30647) );
  XOR U30859 ( .A(n30645), .B(n30647), .Z(n30650) );
  XOR U30860 ( .A(n30648), .B(n30650), .Z(n30671) );
  XOR U30861 ( .A(n30669), .B(n30671), .Z(n30672) );
  XOR U30862 ( .A(n30673), .B(n30672), .Z(n30639) );
  XOR U30863 ( .A(n30640), .B(n30639), .Z(n30676) );
  XOR U30864 ( .A(n30558), .B(n30676), .Z(n30680) );
  XOR U30865 ( .A(n30678), .B(n30680), .Z(n30683) );
  XOR U30866 ( .A(n30684), .B(n30683), .Z(n30685) );
  XOR U30867 ( .A(n30686), .B(n30685), .Z(n30633) );
  NOR U30868 ( .A(n30560), .B(n30559), .Z(n30565) );
  IV U30869 ( .A(n30561), .Z(n30562) );
  NOR U30870 ( .A(n30563), .B(n30562), .Z(n30564) );
  NOR U30871 ( .A(n30565), .B(n30564), .Z(n30631) );
  NOR U30872 ( .A(n156), .B(n151), .Z(n30629) );
  XOR U30873 ( .A(n30631), .B(n30629), .Z(n30632) );
  XOR U30874 ( .A(n30633), .B(n30632), .Z(n30693) );
  IV U30875 ( .A(n30566), .Z(n30568) );
  NOR U30876 ( .A(n30568), .B(n30567), .Z(n30573) );
  IV U30877 ( .A(n30569), .Z(n30570) );
  NOR U30878 ( .A(n30571), .B(n30570), .Z(n30572) );
  NOR U30879 ( .A(n30573), .B(n30572), .Z(n30692) );
  NOR U30880 ( .A(n158), .B(n149), .Z(n30690) );
  XOR U30881 ( .A(n30692), .B(n30690), .Z(n30695) );
  XOR U30882 ( .A(n30693), .B(n30695), .Z(n30623) );
  XOR U30883 ( .A(n30621), .B(n30623), .Z(n30624) );
  XOR U30884 ( .A(n30625), .B(n30624), .Z(n30701) );
  NOR U30885 ( .A(n30575), .B(n30574), .Z(n30580) );
  IV U30886 ( .A(n30576), .Z(n30577) );
  NOR U30887 ( .A(n30578), .B(n30577), .Z(n30579) );
  NOR U30888 ( .A(n30580), .B(n30579), .Z(n30700) );
  NOR U30889 ( .A(n163), .B(n144), .Z(n30698) );
  XOR U30890 ( .A(n30700), .B(n30698), .Z(n30703) );
  XOR U30891 ( .A(n30701), .B(n30703), .Z(n30617) );
  NOR U30892 ( .A(n30582), .B(n30581), .Z(n30587) );
  IV U30893 ( .A(n30583), .Z(n30585) );
  NOR U30894 ( .A(n30585), .B(n30584), .Z(n30586) );
  NOR U30895 ( .A(n30587), .B(n30586), .Z(n30616) );
  NOR U30896 ( .A(n165), .B(n142), .Z(n30614) );
  XOR U30897 ( .A(n30616), .B(n30614), .Z(n30618) );
  XOR U30898 ( .A(n30617), .B(n30618), .Z(n30606) );
  XOR U30899 ( .A(n30608), .B(n30606), .Z(n30611) );
  XOR U30900 ( .A(n30609), .B(n30611), .Z(n30604) );
  XOR U30901 ( .A(n30588), .B(n30604), .Z(n30599) );
  XOR U30902 ( .A(n30597), .B(n30599), .Z(n30601) );
  NOR U30903 ( .A(n30590), .B(n30589), .Z(n30595) );
  IV U30904 ( .A(n30591), .Z(n30592) );
  NOR U30905 ( .A(n30593), .B(n30592), .Z(n30594) );
  NOR U30906 ( .A(n30595), .B(n30594), .Z(n30596) );
  IV U30907 ( .A(n30596), .Z(n30600) );
  XOR U30908 ( .A(n30601), .B(n30600), .Z(c[113]) );
  IV U30909 ( .A(n30597), .Z(n30598) );
  NOR U30910 ( .A(n30599), .B(n30598), .Z(n30603) );
  NOR U30911 ( .A(n30601), .B(n30600), .Z(n30602) );
  NOR U30912 ( .A(n30603), .B(n30602), .Z(n30711) );
  NOR U30913 ( .A(n30605), .B(n30604), .Z(n30707) );
  IV U30914 ( .A(n30606), .Z(n30607) );
  NOR U30915 ( .A(n30608), .B(n30607), .Z(n30613) );
  IV U30916 ( .A(n30609), .Z(n30610) );
  NOR U30917 ( .A(n30611), .B(n30610), .Z(n30612) );
  NOR U30918 ( .A(n30613), .B(n30612), .Z(n30714) );
  IV U30919 ( .A(n30714), .Z(n30706) );
  NOR U30920 ( .A(n167), .B(n142), .Z(n30718) );
  IV U30921 ( .A(n30614), .Z(n30615) );
  NOR U30922 ( .A(n30616), .B(n30615), .Z(n30620) );
  NOR U30923 ( .A(n30618), .B(n30617), .Z(n30619) );
  NOR U30924 ( .A(n30620), .B(n30619), .Z(n30717) );
  NOR U30925 ( .A(n163), .B(n146), .Z(n30733) );
  IV U30926 ( .A(n30621), .Z(n30622) );
  NOR U30927 ( .A(n30623), .B(n30622), .Z(n30627) );
  NOR U30928 ( .A(n30625), .B(n30624), .Z(n30626) );
  NOR U30929 ( .A(n30627), .B(n30626), .Z(n30732) );
  NOR U30930 ( .A(n158), .B(n151), .Z(n30628) );
  IV U30931 ( .A(n30628), .Z(n30741) );
  IV U30932 ( .A(n30629), .Z(n30630) );
  NOR U30933 ( .A(n30631), .B(n30630), .Z(n30635) );
  NOR U30934 ( .A(n30633), .B(n30632), .Z(n30634) );
  NOR U30935 ( .A(n30635), .B(n30634), .Z(n30739) );
  NOR U30936 ( .A(n153), .B(n157), .Z(n30789) );
  IV U30937 ( .A(n30636), .Z(n30638) );
  NOR U30938 ( .A(n30638), .B(n30637), .Z(n30643) );
  IV U30939 ( .A(n30639), .Z(n30641) );
  NOR U30940 ( .A(n30641), .B(n30640), .Z(n30642) );
  NOR U30941 ( .A(n30643), .B(n30642), .Z(n30788) );
  NOR U30942 ( .A(n148), .B(n160), .Z(n30644) );
  IV U30943 ( .A(n30644), .Z(n30781) );
  IV U30944 ( .A(n30645), .Z(n30646) );
  NOR U30945 ( .A(n30647), .B(n30646), .Z(n30652) );
  IV U30946 ( .A(n30648), .Z(n30649) );
  NOR U30947 ( .A(n30650), .B(n30649), .Z(n30651) );
  NOR U30948 ( .A(n30652), .B(n30651), .Z(n30779) );
  NOR U30949 ( .A(n147), .B(n162), .Z(n30763) );
  NOR U30950 ( .A(n30654), .B(n30653), .Z(n30659) );
  IV U30951 ( .A(n30655), .Z(n30656) );
  NOR U30952 ( .A(n30657), .B(n30656), .Z(n30658) );
  NOR U30953 ( .A(n30659), .B(n30658), .Z(n30762) );
  IV U30954 ( .A(n30762), .Z(n30668) );
  NOR U30955 ( .A(n164), .B(n145), .Z(n30771) );
  IV U30956 ( .A(n30660), .Z(n30661) );
  NOR U30957 ( .A(n30662), .B(n30661), .Z(n30667) );
  IV U30958 ( .A(n30663), .Z(n30664) );
  NOR U30959 ( .A(n30665), .B(n30664), .Z(n30666) );
  NOR U30960 ( .A(n30667), .B(n30666), .Z(n30770) );
  NOR U30961 ( .A(n166), .B(n143), .Z(n30768) );
  XOR U30962 ( .A(n30770), .B(n30768), .Z(n30773) );
  XOR U30963 ( .A(n30771), .B(n30773), .Z(n30761) );
  XOR U30964 ( .A(n30668), .B(n30761), .Z(n30765) );
  XOR U30965 ( .A(n30763), .B(n30765), .Z(n30778) );
  XOR U30966 ( .A(n30779), .B(n30778), .Z(n30780) );
  XOR U30967 ( .A(n30781), .B(n30780), .Z(n30757) );
  IV U30968 ( .A(n30669), .Z(n30670) );
  NOR U30969 ( .A(n30671), .B(n30670), .Z(n30675) );
  NOR U30970 ( .A(n30673), .B(n30672), .Z(n30674) );
  NOR U30971 ( .A(n30675), .B(n30674), .Z(n30756) );
  NOR U30972 ( .A(n150), .B(n159), .Z(n30754) );
  XOR U30973 ( .A(n30756), .B(n30754), .Z(n30758) );
  XOR U30974 ( .A(n30757), .B(n30758), .Z(n30786) );
  XOR U30975 ( .A(n30788), .B(n30786), .Z(n30791) );
  XOR U30976 ( .A(n30789), .B(n30791), .Z(n30797) );
  NOR U30977 ( .A(n30677), .B(n30676), .Z(n30682) );
  IV U30978 ( .A(n30678), .Z(n30679) );
  NOR U30979 ( .A(n30680), .B(n30679), .Z(n30681) );
  NOR U30980 ( .A(n30682), .B(n30681), .Z(n30796) );
  NOR U30981 ( .A(n155), .B(n154), .Z(n30794) );
  XOR U30982 ( .A(n30796), .B(n30794), .Z(n30798) );
  XOR U30983 ( .A(n30797), .B(n30798), .Z(n30749) );
  NOR U30984 ( .A(n30684), .B(n30683), .Z(n30689) );
  IV U30985 ( .A(n30685), .Z(n30687) );
  NOR U30986 ( .A(n30687), .B(n30686), .Z(n30688) );
  NOR U30987 ( .A(n30689), .B(n30688), .Z(n30748) );
  NOR U30988 ( .A(n156), .B(n152), .Z(n30746) );
  XOR U30989 ( .A(n30748), .B(n30746), .Z(n30751) );
  XOR U30990 ( .A(n30749), .B(n30751), .Z(n30738) );
  XOR U30991 ( .A(n30739), .B(n30738), .Z(n30740) );
  XOR U30992 ( .A(n30741), .B(n30740), .Z(n30804) );
  IV U30993 ( .A(n30690), .Z(n30691) );
  NOR U30994 ( .A(n30692), .B(n30691), .Z(n30697) );
  IV U30995 ( .A(n30693), .Z(n30694) );
  NOR U30996 ( .A(n30695), .B(n30694), .Z(n30696) );
  NOR U30997 ( .A(n30697), .B(n30696), .Z(n30803) );
  NOR U30998 ( .A(n161), .B(n149), .Z(n30801) );
  XOR U30999 ( .A(n30803), .B(n30801), .Z(n30805) );
  XOR U31000 ( .A(n30804), .B(n30805), .Z(n30730) );
  XOR U31001 ( .A(n30732), .B(n30730), .Z(n30735) );
  XOR U31002 ( .A(n30733), .B(n30735), .Z(n30726) );
  IV U31003 ( .A(n30698), .Z(n30699) );
  NOR U31004 ( .A(n30700), .B(n30699), .Z(n30705) );
  IV U31005 ( .A(n30701), .Z(n30702) );
  NOR U31006 ( .A(n30703), .B(n30702), .Z(n30704) );
  NOR U31007 ( .A(n30705), .B(n30704), .Z(n30725) );
  NOR U31008 ( .A(n165), .B(n144), .Z(n30723) );
  XOR U31009 ( .A(n30725), .B(n30723), .Z(n30727) );
  XOR U31010 ( .A(n30726), .B(n30727), .Z(n30715) );
  XOR U31011 ( .A(n30717), .B(n30715), .Z(n30720) );
  XOR U31012 ( .A(n30718), .B(n30720), .Z(n30713) );
  XOR U31013 ( .A(n30706), .B(n30713), .Z(n30709) );
  XOR U31014 ( .A(n30707), .B(n30709), .Z(n30710) );
  XOR U31015 ( .A(n30711), .B(n30710), .Z(c[114]) );
  IV U31016 ( .A(n30707), .Z(n30708) );
  NOR U31017 ( .A(n30709), .B(n30708), .Z(n30712) );
  NOR U31018 ( .A(n30711), .B(n30710), .Z(n30901) );
  NOR U31019 ( .A(n30712), .B(n30901), .Z(n30910) );
  NOR U31020 ( .A(n30714), .B(n30713), .Z(n30895) );
  IV U31021 ( .A(n30895), .Z(n30904) );
  IV U31022 ( .A(n30715), .Z(n30716) );
  NOR U31023 ( .A(n30717), .B(n30716), .Z(n30722) );
  IV U31024 ( .A(n30718), .Z(n30719) );
  NOR U31025 ( .A(n30720), .B(n30719), .Z(n30721) );
  NOR U31026 ( .A(n30722), .B(n30721), .Z(n30893) );
  NOR U31027 ( .A(n167), .B(n144), .Z(n30812) );
  IV U31028 ( .A(n30723), .Z(n30724) );
  NOR U31029 ( .A(n30725), .B(n30724), .Z(n30729) );
  NOR U31030 ( .A(n30727), .B(n30726), .Z(n30728) );
  NOR U31031 ( .A(n30729), .B(n30728), .Z(n30811) );
  IV U31032 ( .A(n30811), .Z(n30809) );
  NOR U31033 ( .A(n165), .B(n146), .Z(n30819) );
  IV U31034 ( .A(n30730), .Z(n30731) );
  NOR U31035 ( .A(n30732), .B(n30731), .Z(n30737) );
  IV U31036 ( .A(n30733), .Z(n30734) );
  NOR U31037 ( .A(n30735), .B(n30734), .Z(n30736) );
  NOR U31038 ( .A(n30737), .B(n30736), .Z(n30818) );
  NOR U31039 ( .A(n30739), .B(n30738), .Z(n30744) );
  IV U31040 ( .A(n30740), .Z(n30742) );
  NOR U31041 ( .A(n30742), .B(n30741), .Z(n30743) );
  NOR U31042 ( .A(n30744), .B(n30743), .Z(n30889) );
  NOR U31043 ( .A(n161), .B(n151), .Z(n30885) );
  NOR U31044 ( .A(n158), .B(n152), .Z(n30745) );
  IV U31045 ( .A(n30745), .Z(n30835) );
  IV U31046 ( .A(n30746), .Z(n30747) );
  NOR U31047 ( .A(n30748), .B(n30747), .Z(n30753) );
  IV U31048 ( .A(n30749), .Z(n30750) );
  NOR U31049 ( .A(n30751), .B(n30750), .Z(n30752) );
  NOR U31050 ( .A(n30753), .B(n30752), .Z(n30833) );
  NOR U31051 ( .A(n153), .B(n159), .Z(n30872) );
  IV U31052 ( .A(n30754), .Z(n30755) );
  NOR U31053 ( .A(n30756), .B(n30755), .Z(n30760) );
  NOR U31054 ( .A(n30758), .B(n30757), .Z(n30759) );
  NOR U31055 ( .A(n30760), .B(n30759), .Z(n30870) );
  IV U31056 ( .A(n30870), .Z(n30785) );
  NOR U31057 ( .A(n150), .B(n160), .Z(n30852) );
  NOR U31058 ( .A(n30762), .B(n30761), .Z(n30767) );
  IV U31059 ( .A(n30763), .Z(n30764) );
  NOR U31060 ( .A(n30765), .B(n30764), .Z(n30766) );
  NOR U31061 ( .A(n30767), .B(n30766), .Z(n30856) );
  NOR U31062 ( .A(n164), .B(n147), .Z(n30864) );
  IV U31063 ( .A(n30768), .Z(n30769) );
  NOR U31064 ( .A(n30770), .B(n30769), .Z(n30775) );
  IV U31065 ( .A(n30771), .Z(n30772) );
  NOR U31066 ( .A(n30773), .B(n30772), .Z(n30774) );
  NOR U31067 ( .A(n30775), .B(n30774), .Z(n30863) );
  NOR U31068 ( .A(n166), .B(n145), .Z(n30861) );
  XOR U31069 ( .A(n30863), .B(n30861), .Z(n30866) );
  XOR U31070 ( .A(n30864), .B(n30866), .Z(n30855) );
  XOR U31071 ( .A(n30856), .B(n30855), .Z(n30776) );
  IV U31072 ( .A(n30776), .Z(n30858) );
  NOR U31073 ( .A(n148), .B(n162), .Z(n30777) );
  IV U31074 ( .A(n30777), .Z(n30857) );
  XOR U31075 ( .A(n30858), .B(n30857), .Z(n30850) );
  NOR U31076 ( .A(n30779), .B(n30778), .Z(n30784) );
  IV U31077 ( .A(n30780), .Z(n30782) );
  NOR U31078 ( .A(n30782), .B(n30781), .Z(n30783) );
  NOR U31079 ( .A(n30784), .B(n30783), .Z(n30848) );
  XOR U31080 ( .A(n30850), .B(n30848), .Z(n30851) );
  XOR U31081 ( .A(n30852), .B(n30851), .Z(n30871) );
  XOR U31082 ( .A(n30785), .B(n30871), .Z(n30874) );
  XOR U31083 ( .A(n30872), .B(n30874), .Z(n30880) );
  IV U31084 ( .A(n30786), .Z(n30787) );
  NOR U31085 ( .A(n30788), .B(n30787), .Z(n30793) );
  IV U31086 ( .A(n30789), .Z(n30790) );
  NOR U31087 ( .A(n30791), .B(n30790), .Z(n30792) );
  NOR U31088 ( .A(n30793), .B(n30792), .Z(n30879) );
  NOR U31089 ( .A(n155), .B(n157), .Z(n30877) );
  XOR U31090 ( .A(n30879), .B(n30877), .Z(n30881) );
  XOR U31091 ( .A(n30880), .B(n30881), .Z(n30843) );
  IV U31092 ( .A(n30794), .Z(n30795) );
  NOR U31093 ( .A(n30796), .B(n30795), .Z(n30800) );
  NOR U31094 ( .A(n30798), .B(n30797), .Z(n30799) );
  NOR U31095 ( .A(n30800), .B(n30799), .Z(n30842) );
  NOR U31096 ( .A(n156), .B(n154), .Z(n30840) );
  XOR U31097 ( .A(n30842), .B(n30840), .Z(n30844) );
  XOR U31098 ( .A(n30843), .B(n30844), .Z(n30832) );
  XOR U31099 ( .A(n30833), .B(n30832), .Z(n30834) );
  XOR U31100 ( .A(n30835), .B(n30834), .Z(n30887) );
  XOR U31101 ( .A(n30885), .B(n30887), .Z(n30888) );
  XOR U31102 ( .A(n30889), .B(n30888), .Z(n30827) );
  IV U31103 ( .A(n30801), .Z(n30802) );
  NOR U31104 ( .A(n30803), .B(n30802), .Z(n30807) );
  NOR U31105 ( .A(n30805), .B(n30804), .Z(n30806) );
  NOR U31106 ( .A(n30807), .B(n30806), .Z(n30826) );
  NOR U31107 ( .A(n163), .B(n149), .Z(n30824) );
  XOR U31108 ( .A(n30826), .B(n30824), .Z(n30828) );
  XOR U31109 ( .A(n30827), .B(n30828), .Z(n30817) );
  XOR U31110 ( .A(n30818), .B(n30817), .Z(n30808) );
  IV U31111 ( .A(n30808), .Z(n30821) );
  XOR U31112 ( .A(n30819), .B(n30821), .Z(n30810) );
  XOR U31113 ( .A(n30809), .B(n30810), .Z(n30814) );
  XOR U31114 ( .A(n30812), .B(n30814), .Z(n30892) );
  XOR U31115 ( .A(n30893), .B(n30892), .Z(n30894) );
  XOR U31116 ( .A(n30904), .B(n30894), .Z(n30896) );
  XOR U31117 ( .A(n30910), .B(n30896), .Z(c[115]) );
  NOR U31118 ( .A(n30811), .B(n30810), .Z(n30816) );
  IV U31119 ( .A(n30812), .Z(n30813) );
  NOR U31120 ( .A(n30814), .B(n30813), .Z(n30815) );
  NOR U31121 ( .A(n30816), .B(n30815), .Z(n30918) );
  NOR U31122 ( .A(n30818), .B(n30817), .Z(n30823) );
  IV U31123 ( .A(n30819), .Z(n30820) );
  NOR U31124 ( .A(n30821), .B(n30820), .Z(n30822) );
  NOR U31125 ( .A(n30823), .B(n30822), .Z(n30923) );
  NOR U31126 ( .A(n167), .B(n146), .Z(n30919) );
  NOR U31127 ( .A(n165), .B(n149), .Z(n30991) );
  IV U31128 ( .A(n30824), .Z(n30825) );
  NOR U31129 ( .A(n30826), .B(n30825), .Z(n30831) );
  IV U31130 ( .A(n30827), .Z(n30829) );
  NOR U31131 ( .A(n30829), .B(n30828), .Z(n30830) );
  NOR U31132 ( .A(n30831), .B(n30830), .Z(n30990) );
  NOR U31133 ( .A(n161), .B(n152), .Z(n30982) );
  NOR U31134 ( .A(n30833), .B(n30832), .Z(n30838) );
  IV U31135 ( .A(n30834), .Z(n30836) );
  NOR U31136 ( .A(n30836), .B(n30835), .Z(n30837) );
  NOR U31137 ( .A(n30838), .B(n30837), .Z(n30981) );
  IV U31138 ( .A(n30981), .Z(n30884) );
  NOR U31139 ( .A(n158), .B(n154), .Z(n30839) );
  IV U31140 ( .A(n30839), .Z(n30936) );
  IV U31141 ( .A(n30840), .Z(n30841) );
  NOR U31142 ( .A(n30842), .B(n30841), .Z(n30847) );
  IV U31143 ( .A(n30843), .Z(n30845) );
  NOR U31144 ( .A(n30845), .B(n30844), .Z(n30846) );
  NOR U31145 ( .A(n30847), .B(n30846), .Z(n30934) );
  IV U31146 ( .A(n30848), .Z(n30849) );
  NOR U31147 ( .A(n30850), .B(n30849), .Z(n30854) );
  NOR U31148 ( .A(n30852), .B(n30851), .Z(n30853) );
  NOR U31149 ( .A(n30854), .B(n30853), .Z(n30952) );
  NOR U31150 ( .A(n153), .B(n160), .Z(n30949) );
  NOR U31151 ( .A(n150), .B(n162), .Z(n30959) );
  NOR U31152 ( .A(n30856), .B(n30855), .Z(n30860) );
  NOR U31153 ( .A(n30858), .B(n30857), .Z(n30859) );
  NOR U31154 ( .A(n30860), .B(n30859), .Z(n30958) );
  IV U31155 ( .A(n30958), .Z(n30869) );
  NOR U31156 ( .A(n164), .B(n148), .Z(n30967) );
  IV U31157 ( .A(n30861), .Z(n30862) );
  NOR U31158 ( .A(n30863), .B(n30862), .Z(n30868) );
  IV U31159 ( .A(n30864), .Z(n30865) );
  NOR U31160 ( .A(n30866), .B(n30865), .Z(n30867) );
  NOR U31161 ( .A(n30868), .B(n30867), .Z(n30966) );
  NOR U31162 ( .A(n166), .B(n147), .Z(n30964) );
  XOR U31163 ( .A(n30966), .B(n30964), .Z(n30969) );
  XOR U31164 ( .A(n30967), .B(n30969), .Z(n30957) );
  XOR U31165 ( .A(n30869), .B(n30957), .Z(n30961) );
  XOR U31166 ( .A(n30959), .B(n30961), .Z(n30951) );
  XOR U31167 ( .A(n30949), .B(n30951), .Z(n30954) );
  XOR U31168 ( .A(n30952), .B(n30954), .Z(n30976) );
  NOR U31169 ( .A(n30871), .B(n30870), .Z(n30876) );
  IV U31170 ( .A(n30872), .Z(n30873) );
  NOR U31171 ( .A(n30874), .B(n30873), .Z(n30875) );
  NOR U31172 ( .A(n30876), .B(n30875), .Z(n30975) );
  NOR U31173 ( .A(n155), .B(n159), .Z(n30973) );
  XOR U31174 ( .A(n30975), .B(n30973), .Z(n30977) );
  XOR U31175 ( .A(n30976), .B(n30977), .Z(n30943) );
  IV U31176 ( .A(n30877), .Z(n30878) );
  NOR U31177 ( .A(n30879), .B(n30878), .Z(n30883) );
  NOR U31178 ( .A(n30881), .B(n30880), .Z(n30882) );
  NOR U31179 ( .A(n30883), .B(n30882), .Z(n30942) );
  NOR U31180 ( .A(n156), .B(n157), .Z(n30940) );
  XOR U31181 ( .A(n30942), .B(n30940), .Z(n30944) );
  XOR U31182 ( .A(n30943), .B(n30944), .Z(n30933) );
  XOR U31183 ( .A(n30934), .B(n30933), .Z(n30935) );
  XOR U31184 ( .A(n30936), .B(n30935), .Z(n30980) );
  XOR U31185 ( .A(n30884), .B(n30980), .Z(n30984) );
  XOR U31186 ( .A(n30982), .B(n30984), .Z(n30930) );
  IV U31187 ( .A(n30885), .Z(n30886) );
  NOR U31188 ( .A(n30887), .B(n30886), .Z(n30891) );
  NOR U31189 ( .A(n30889), .B(n30888), .Z(n30890) );
  NOR U31190 ( .A(n30891), .B(n30890), .Z(n30928) );
  NOR U31191 ( .A(n163), .B(n151), .Z(n30926) );
  XOR U31192 ( .A(n30928), .B(n30926), .Z(n30929) );
  XOR U31193 ( .A(n30930), .B(n30929), .Z(n30988) );
  XOR U31194 ( .A(n30990), .B(n30988), .Z(n30993) );
  XOR U31195 ( .A(n30991), .B(n30993), .Z(n30921) );
  XOR U31196 ( .A(n30919), .B(n30921), .Z(n30922) );
  XOR U31197 ( .A(n30923), .B(n30922), .Z(n30916) );
  XOR U31198 ( .A(n30918), .B(n30916), .Z(n30912) );
  NOR U31199 ( .A(n30893), .B(n30892), .Z(n30902) );
  NOR U31200 ( .A(n30895), .B(n30894), .Z(n30899) );
  IV U31201 ( .A(n30910), .Z(n30897) );
  NOR U31202 ( .A(n30897), .B(n30896), .Z(n30898) );
  NOR U31203 ( .A(n30899), .B(n30898), .Z(n30900) );
  NOR U31204 ( .A(n30902), .B(n30900), .Z(n30913) );
  IV U31205 ( .A(n30901), .Z(n30906) );
  IV U31206 ( .A(n30902), .Z(n30903) );
  NOR U31207 ( .A(n30904), .B(n30903), .Z(n30905) );
  IV U31208 ( .A(n30905), .Z(n30911) );
  NOR U31209 ( .A(n30906), .B(n30911), .Z(n30907) );
  NOR U31210 ( .A(n30913), .B(n30907), .Z(n30908) );
  XOR U31211 ( .A(n30912), .B(n30908), .Z(n30909) );
  IV U31212 ( .A(n30909), .Z(c[116]) );
  NOR U31213 ( .A(n30911), .B(n30910), .Z(n30915) );
  NOR U31214 ( .A(n30913), .B(n30912), .Z(n30914) );
  NOR U31215 ( .A(n30915), .B(n30914), .Z(n31069) );
  IV U31216 ( .A(n30916), .Z(n30917) );
  NOR U31217 ( .A(n30918), .B(n30917), .Z(n31072) );
  IV U31218 ( .A(n30919), .Z(n30920) );
  NOR U31219 ( .A(n30921), .B(n30920), .Z(n30925) );
  NOR U31220 ( .A(n30923), .B(n30922), .Z(n30924) );
  NOR U31221 ( .A(n30925), .B(n30924), .Z(n31067) );
  IV U31222 ( .A(n30926), .Z(n30927) );
  NOR U31223 ( .A(n30928), .B(n30927), .Z(n30932) );
  NOR U31224 ( .A(n30930), .B(n30929), .Z(n30931) );
  NOR U31225 ( .A(n30932), .B(n30931), .Z(n31059) );
  NOR U31226 ( .A(n30934), .B(n30933), .Z(n30939) );
  IV U31227 ( .A(n30935), .Z(n30937) );
  NOR U31228 ( .A(n30937), .B(n30936), .Z(n30938) );
  NOR U31229 ( .A(n30939), .B(n30938), .Z(n31055) );
  NOR U31230 ( .A(n161), .B(n154), .Z(n31051) );
  NOR U31231 ( .A(n158), .B(n157), .Z(n31046) );
  IV U31232 ( .A(n30940), .Z(n30941) );
  NOR U31233 ( .A(n30942), .B(n30941), .Z(n30947) );
  IV U31234 ( .A(n30943), .Z(n30945) );
  NOR U31235 ( .A(n30945), .B(n30944), .Z(n30946) );
  NOR U31236 ( .A(n30947), .B(n30946), .Z(n31045) );
  NOR U31237 ( .A(n155), .B(n160), .Z(n30948) );
  IV U31238 ( .A(n30948), .Z(n31038) );
  IV U31239 ( .A(n30949), .Z(n30950) );
  NOR U31240 ( .A(n30951), .B(n30950), .Z(n30956) );
  IV U31241 ( .A(n30952), .Z(n30953) );
  NOR U31242 ( .A(n30954), .B(n30953), .Z(n30955) );
  NOR U31243 ( .A(n30956), .B(n30955), .Z(n31036) );
  NOR U31244 ( .A(n153), .B(n162), .Z(n31020) );
  NOR U31245 ( .A(n30958), .B(n30957), .Z(n30963) );
  IV U31246 ( .A(n30959), .Z(n30960) );
  NOR U31247 ( .A(n30961), .B(n30960), .Z(n30962) );
  NOR U31248 ( .A(n30963), .B(n30962), .Z(n31019) );
  IV U31249 ( .A(n31019), .Z(n30972) );
  NOR U31250 ( .A(n164), .B(n150), .Z(n31028) );
  IV U31251 ( .A(n30964), .Z(n30965) );
  NOR U31252 ( .A(n30966), .B(n30965), .Z(n30971) );
  IV U31253 ( .A(n30967), .Z(n30968) );
  NOR U31254 ( .A(n30969), .B(n30968), .Z(n30970) );
  NOR U31255 ( .A(n30971), .B(n30970), .Z(n31027) );
  NOR U31256 ( .A(n166), .B(n148), .Z(n31025) );
  XOR U31257 ( .A(n31027), .B(n31025), .Z(n31030) );
  XOR U31258 ( .A(n31028), .B(n31030), .Z(n31018) );
  XOR U31259 ( .A(n30972), .B(n31018), .Z(n31022) );
  XOR U31260 ( .A(n31020), .B(n31022), .Z(n31035) );
  XOR U31261 ( .A(n31036), .B(n31035), .Z(n31037) );
  XOR U31262 ( .A(n31038), .B(n31037), .Z(n31014) );
  IV U31263 ( .A(n30973), .Z(n30974) );
  NOR U31264 ( .A(n30975), .B(n30974), .Z(n30979) );
  NOR U31265 ( .A(n30977), .B(n30976), .Z(n30978) );
  NOR U31266 ( .A(n30979), .B(n30978), .Z(n31013) );
  NOR U31267 ( .A(n156), .B(n159), .Z(n31011) );
  XOR U31268 ( .A(n31013), .B(n31011), .Z(n31015) );
  XOR U31269 ( .A(n31014), .B(n31015), .Z(n31043) );
  XOR U31270 ( .A(n31045), .B(n31043), .Z(n31048) );
  XOR U31271 ( .A(n31046), .B(n31048), .Z(n31053) );
  XOR U31272 ( .A(n31051), .B(n31053), .Z(n31054) );
  XOR U31273 ( .A(n31055), .B(n31054), .Z(n31006) );
  NOR U31274 ( .A(n30981), .B(n30980), .Z(n30986) );
  IV U31275 ( .A(n30982), .Z(n30983) );
  NOR U31276 ( .A(n30984), .B(n30983), .Z(n30985) );
  NOR U31277 ( .A(n30986), .B(n30985), .Z(n31005) );
  NOR U31278 ( .A(n163), .B(n152), .Z(n31003) );
  XOR U31279 ( .A(n31005), .B(n31003), .Z(n31007) );
  XOR U31280 ( .A(n31006), .B(n31007), .Z(n31058) );
  XOR U31281 ( .A(n31059), .B(n31058), .Z(n31060) );
  NOR U31282 ( .A(n165), .B(n151), .Z(n30987) );
  IV U31283 ( .A(n30987), .Z(n31061) );
  XOR U31284 ( .A(n31060), .B(n31061), .Z(n30999) );
  IV U31285 ( .A(n30988), .Z(n30989) );
  NOR U31286 ( .A(n30990), .B(n30989), .Z(n30995) );
  IV U31287 ( .A(n30991), .Z(n30992) );
  NOR U31288 ( .A(n30993), .B(n30992), .Z(n30994) );
  NOR U31289 ( .A(n30995), .B(n30994), .Z(n30998) );
  NOR U31290 ( .A(n167), .B(n149), .Z(n30996) );
  XOR U31291 ( .A(n30998), .B(n30996), .Z(n31000) );
  XOR U31292 ( .A(n30999), .B(n31000), .Z(n31065) );
  XOR U31293 ( .A(n31067), .B(n31065), .Z(n31073) );
  XOR U31294 ( .A(n31072), .B(n31073), .Z(n31068) );
  XOR U31295 ( .A(n31069), .B(n31068), .Z(c[117]) );
  IV U31296 ( .A(n30996), .Z(n30997) );
  NOR U31297 ( .A(n30998), .B(n30997), .Z(n31002) );
  NOR U31298 ( .A(n31000), .B(n30999), .Z(n31001) );
  NOR U31299 ( .A(n31002), .B(n31001), .Z(n31082) );
  IV U31300 ( .A(n31003), .Z(n31004) );
  NOR U31301 ( .A(n31005), .B(n31004), .Z(n31010) );
  IV U31302 ( .A(n31006), .Z(n31008) );
  NOR U31303 ( .A(n31008), .B(n31007), .Z(n31009) );
  NOR U31304 ( .A(n31010), .B(n31009), .Z(n31144) );
  NOR U31305 ( .A(n158), .B(n159), .Z(n31129) );
  IV U31306 ( .A(n31011), .Z(n31012) );
  NOR U31307 ( .A(n31013), .B(n31012), .Z(n31017) );
  NOR U31308 ( .A(n31015), .B(n31014), .Z(n31016) );
  NOR U31309 ( .A(n31017), .B(n31016), .Z(n31127) );
  IV U31310 ( .A(n31127), .Z(n31042) );
  NOR U31311 ( .A(n156), .B(n160), .Z(n31109) );
  NOR U31312 ( .A(n31019), .B(n31018), .Z(n31024) );
  IV U31313 ( .A(n31020), .Z(n31021) );
  NOR U31314 ( .A(n31022), .B(n31021), .Z(n31023) );
  NOR U31315 ( .A(n31024), .B(n31023), .Z(n31113) );
  NOR U31316 ( .A(n164), .B(n153), .Z(n31121) );
  IV U31317 ( .A(n31025), .Z(n31026) );
  NOR U31318 ( .A(n31027), .B(n31026), .Z(n31032) );
  IV U31319 ( .A(n31028), .Z(n31029) );
  NOR U31320 ( .A(n31030), .B(n31029), .Z(n31031) );
  NOR U31321 ( .A(n31032), .B(n31031), .Z(n31120) );
  NOR U31322 ( .A(n166), .B(n150), .Z(n31118) );
  XOR U31323 ( .A(n31120), .B(n31118), .Z(n31123) );
  XOR U31324 ( .A(n31121), .B(n31123), .Z(n31112) );
  XOR U31325 ( .A(n31113), .B(n31112), .Z(n31033) );
  IV U31326 ( .A(n31033), .Z(n31115) );
  NOR U31327 ( .A(n155), .B(n162), .Z(n31034) );
  IV U31328 ( .A(n31034), .Z(n31114) );
  XOR U31329 ( .A(n31115), .B(n31114), .Z(n31107) );
  NOR U31330 ( .A(n31036), .B(n31035), .Z(n31041) );
  IV U31331 ( .A(n31037), .Z(n31039) );
  NOR U31332 ( .A(n31039), .B(n31038), .Z(n31040) );
  NOR U31333 ( .A(n31041), .B(n31040), .Z(n31105) );
  XOR U31334 ( .A(n31107), .B(n31105), .Z(n31108) );
  XOR U31335 ( .A(n31109), .B(n31108), .Z(n31128) );
  XOR U31336 ( .A(n31042), .B(n31128), .Z(n31131) );
  XOR U31337 ( .A(n31129), .B(n31131), .Z(n31137) );
  IV U31338 ( .A(n31043), .Z(n31044) );
  NOR U31339 ( .A(n31045), .B(n31044), .Z(n31050) );
  IV U31340 ( .A(n31046), .Z(n31047) );
  NOR U31341 ( .A(n31048), .B(n31047), .Z(n31049) );
  NOR U31342 ( .A(n31050), .B(n31049), .Z(n31136) );
  NOR U31343 ( .A(n161), .B(n157), .Z(n31134) );
  XOR U31344 ( .A(n31136), .B(n31134), .Z(n31138) );
  XOR U31345 ( .A(n31137), .B(n31138), .Z(n31100) );
  IV U31346 ( .A(n31051), .Z(n31052) );
  NOR U31347 ( .A(n31053), .B(n31052), .Z(n31057) );
  NOR U31348 ( .A(n31055), .B(n31054), .Z(n31056) );
  NOR U31349 ( .A(n31057), .B(n31056), .Z(n31099) );
  NOR U31350 ( .A(n163), .B(n154), .Z(n31097) );
  XOR U31351 ( .A(n31099), .B(n31097), .Z(n31102) );
  XOR U31352 ( .A(n31100), .B(n31102), .Z(n31143) );
  XOR U31353 ( .A(n31144), .B(n31143), .Z(n31145) );
  NOR U31354 ( .A(n165), .B(n152), .Z(n31146) );
  XOR U31355 ( .A(n31145), .B(n31146), .Z(n31094) );
  NOR U31356 ( .A(n167), .B(n151), .Z(n31092) );
  NOR U31357 ( .A(n31059), .B(n31058), .Z(n31064) );
  IV U31358 ( .A(n31060), .Z(n31062) );
  NOR U31359 ( .A(n31062), .B(n31061), .Z(n31063) );
  NOR U31360 ( .A(n31064), .B(n31063), .Z(n31090) );
  XOR U31361 ( .A(n31092), .B(n31090), .Z(n31093) );
  XOR U31362 ( .A(n31094), .B(n31093), .Z(n31081) );
  XOR U31363 ( .A(n31082), .B(n31081), .Z(n31083) );
  IV U31364 ( .A(n31065), .Z(n31066) );
  NOR U31365 ( .A(n31067), .B(n31066), .Z(n31079) );
  IV U31366 ( .A(n31079), .Z(n31071) );
  NOR U31367 ( .A(n31069), .B(n31068), .Z(n31075) );
  IV U31368 ( .A(n31075), .Z(n31070) );
  NOR U31369 ( .A(n31071), .B(n31070), .Z(n31087) );
  IV U31370 ( .A(n31072), .Z(n31074) );
  NOR U31371 ( .A(n31074), .B(n31073), .Z(n31076) );
  NOR U31372 ( .A(n31076), .B(n31075), .Z(n31077) );
  IV U31373 ( .A(n31077), .Z(n31078) );
  NOR U31374 ( .A(n31079), .B(n31078), .Z(n31085) );
  NOR U31375 ( .A(n31087), .B(n31085), .Z(n31080) );
  XOR U31376 ( .A(n31083), .B(n31080), .Z(c[118]) );
  NOR U31377 ( .A(n31082), .B(n31081), .Z(n31212) );
  IV U31378 ( .A(n31212), .Z(n31209) );
  NOR U31379 ( .A(n31087), .B(n31209), .Z(n31089) );
  IV U31380 ( .A(n31083), .Z(n31084) );
  NOR U31381 ( .A(n31085), .B(n31084), .Z(n31086) );
  NOR U31382 ( .A(n31087), .B(n31086), .Z(n31214) );
  NOR U31383 ( .A(n31212), .B(n31214), .Z(n31088) );
  NOR U31384 ( .A(n31089), .B(n31088), .Z(n31151) );
  IV U31385 ( .A(n31090), .Z(n31091) );
  NOR U31386 ( .A(n31092), .B(n31091), .Z(n31096) );
  NOR U31387 ( .A(n31094), .B(n31093), .Z(n31095) );
  NOR U31388 ( .A(n31096), .B(n31095), .Z(n31206) );
  NOR U31389 ( .A(n167), .B(n152), .Z(n31156) );
  IV U31390 ( .A(n31097), .Z(n31098) );
  NOR U31391 ( .A(n31099), .B(n31098), .Z(n31104) );
  IV U31392 ( .A(n31100), .Z(n31101) );
  NOR U31393 ( .A(n31102), .B(n31101), .Z(n31103) );
  NOR U31394 ( .A(n31104), .B(n31103), .Z(n31160) );
  IV U31395 ( .A(n31105), .Z(n31106) );
  NOR U31396 ( .A(n31107), .B(n31106), .Z(n31111) );
  NOR U31397 ( .A(n31109), .B(n31108), .Z(n31110) );
  NOR U31398 ( .A(n31111), .B(n31110), .Z(n31177) );
  NOR U31399 ( .A(n158), .B(n160), .Z(n31174) );
  NOR U31400 ( .A(n156), .B(n162), .Z(n31184) );
  NOR U31401 ( .A(n31113), .B(n31112), .Z(n31117) );
  NOR U31402 ( .A(n31115), .B(n31114), .Z(n31116) );
  NOR U31403 ( .A(n31117), .B(n31116), .Z(n31183) );
  IV U31404 ( .A(n31183), .Z(n31126) );
  NOR U31405 ( .A(n164), .B(n155), .Z(n31192) );
  IV U31406 ( .A(n31118), .Z(n31119) );
  NOR U31407 ( .A(n31120), .B(n31119), .Z(n31125) );
  IV U31408 ( .A(n31121), .Z(n31122) );
  NOR U31409 ( .A(n31123), .B(n31122), .Z(n31124) );
  NOR U31410 ( .A(n31125), .B(n31124), .Z(n31191) );
  NOR U31411 ( .A(n166), .B(n153), .Z(n31189) );
  XOR U31412 ( .A(n31191), .B(n31189), .Z(n31194) );
  XOR U31413 ( .A(n31192), .B(n31194), .Z(n31182) );
  XOR U31414 ( .A(n31126), .B(n31182), .Z(n31186) );
  XOR U31415 ( .A(n31184), .B(n31186), .Z(n31176) );
  XOR U31416 ( .A(n31174), .B(n31176), .Z(n31179) );
  XOR U31417 ( .A(n31177), .B(n31179), .Z(n31202) );
  NOR U31418 ( .A(n31128), .B(n31127), .Z(n31133) );
  IV U31419 ( .A(n31129), .Z(n31130) );
  NOR U31420 ( .A(n31131), .B(n31130), .Z(n31132) );
  NOR U31421 ( .A(n31133), .B(n31132), .Z(n31200) );
  NOR U31422 ( .A(n161), .B(n159), .Z(n31198) );
  XOR U31423 ( .A(n31200), .B(n31198), .Z(n31201) );
  XOR U31424 ( .A(n31202), .B(n31201), .Z(n31168) );
  IV U31425 ( .A(n31134), .Z(n31135) );
  NOR U31426 ( .A(n31136), .B(n31135), .Z(n31140) );
  NOR U31427 ( .A(n31138), .B(n31137), .Z(n31139) );
  NOR U31428 ( .A(n31140), .B(n31139), .Z(n31167) );
  NOR U31429 ( .A(n163), .B(n157), .Z(n31165) );
  XOR U31430 ( .A(n31167), .B(n31165), .Z(n31169) );
  XOR U31431 ( .A(n31168), .B(n31169), .Z(n31159) );
  XOR U31432 ( .A(n31160), .B(n31159), .Z(n31141) );
  IV U31433 ( .A(n31141), .Z(n31162) );
  NOR U31434 ( .A(n165), .B(n154), .Z(n31142) );
  IV U31435 ( .A(n31142), .Z(n31161) );
  XOR U31436 ( .A(n31162), .B(n31161), .Z(n31154) );
  NOR U31437 ( .A(n31144), .B(n31143), .Z(n31150) );
  IV U31438 ( .A(n31145), .Z(n31148) );
  IV U31439 ( .A(n31146), .Z(n31147) );
  NOR U31440 ( .A(n31148), .B(n31147), .Z(n31149) );
  NOR U31441 ( .A(n31150), .B(n31149), .Z(n31152) );
  XOR U31442 ( .A(n31154), .B(n31152), .Z(n31155) );
  XOR U31443 ( .A(n31156), .B(n31155), .Z(n31208) );
  XOR U31444 ( .A(n31206), .B(n31208), .Z(n31210) );
  XOR U31445 ( .A(n31151), .B(n31210), .Z(c[119]) );
  IV U31446 ( .A(n31152), .Z(n31153) );
  NOR U31447 ( .A(n31154), .B(n31153), .Z(n31158) );
  NOR U31448 ( .A(n31156), .B(n31155), .Z(n31157) );
  NOR U31449 ( .A(n31158), .B(n31157), .Z(n31268) );
  NOR U31450 ( .A(n167), .B(n154), .Z(n31220) );
  NOR U31451 ( .A(n31160), .B(n31159), .Z(n31164) );
  NOR U31452 ( .A(n31162), .B(n31161), .Z(n31163) );
  NOR U31453 ( .A(n31164), .B(n31163), .Z(n31219) );
  IV U31454 ( .A(n31219), .Z(n31205) );
  NOR U31455 ( .A(n165), .B(n157), .Z(n31260) );
  IV U31456 ( .A(n31165), .Z(n31166) );
  NOR U31457 ( .A(n31167), .B(n31166), .Z(n31172) );
  IV U31458 ( .A(n31168), .Z(n31170) );
  NOR U31459 ( .A(n31170), .B(n31169), .Z(n31171) );
  NOR U31460 ( .A(n31172), .B(n31171), .Z(n31259) );
  NOR U31461 ( .A(n161), .B(n160), .Z(n31173) );
  IV U31462 ( .A(n31173), .Z(n31252) );
  IV U31463 ( .A(n31174), .Z(n31175) );
  NOR U31464 ( .A(n31176), .B(n31175), .Z(n31181) );
  IV U31465 ( .A(n31177), .Z(n31178) );
  NOR U31466 ( .A(n31179), .B(n31178), .Z(n31180) );
  NOR U31467 ( .A(n31181), .B(n31180), .Z(n31250) );
  NOR U31468 ( .A(n158), .B(n162), .Z(n31234) );
  NOR U31469 ( .A(n31183), .B(n31182), .Z(n31188) );
  IV U31470 ( .A(n31184), .Z(n31185) );
  NOR U31471 ( .A(n31186), .B(n31185), .Z(n31187) );
  NOR U31472 ( .A(n31188), .B(n31187), .Z(n31233) );
  IV U31473 ( .A(n31233), .Z(n31197) );
  NOR U31474 ( .A(n164), .B(n156), .Z(n31242) );
  IV U31475 ( .A(n31189), .Z(n31190) );
  NOR U31476 ( .A(n31191), .B(n31190), .Z(n31196) );
  IV U31477 ( .A(n31192), .Z(n31193) );
  NOR U31478 ( .A(n31194), .B(n31193), .Z(n31195) );
  NOR U31479 ( .A(n31196), .B(n31195), .Z(n31241) );
  NOR U31480 ( .A(n166), .B(n155), .Z(n31239) );
  XOR U31481 ( .A(n31241), .B(n31239), .Z(n31244) );
  XOR U31482 ( .A(n31242), .B(n31244), .Z(n31232) );
  XOR U31483 ( .A(n31197), .B(n31232), .Z(n31236) );
  XOR U31484 ( .A(n31234), .B(n31236), .Z(n31249) );
  XOR U31485 ( .A(n31250), .B(n31249), .Z(n31251) );
  XOR U31486 ( .A(n31252), .B(n31251), .Z(n31228) );
  IV U31487 ( .A(n31198), .Z(n31199) );
  NOR U31488 ( .A(n31200), .B(n31199), .Z(n31204) );
  NOR U31489 ( .A(n31202), .B(n31201), .Z(n31203) );
  NOR U31490 ( .A(n31204), .B(n31203), .Z(n31227) );
  NOR U31491 ( .A(n163), .B(n159), .Z(n31225) );
  XOR U31492 ( .A(n31227), .B(n31225), .Z(n31229) );
  XOR U31493 ( .A(n31228), .B(n31229), .Z(n31257) );
  XOR U31494 ( .A(n31259), .B(n31257), .Z(n31262) );
  XOR U31495 ( .A(n31260), .B(n31262), .Z(n31218) );
  XOR U31496 ( .A(n31205), .B(n31218), .Z(n31222) );
  XOR U31497 ( .A(n31220), .B(n31222), .Z(n31269) );
  XOR U31498 ( .A(n31268), .B(n31269), .Z(n31276) );
  IV U31499 ( .A(n31206), .Z(n31207) );
  NOR U31500 ( .A(n31208), .B(n31207), .Z(n31274) );
  IV U31501 ( .A(n31274), .Z(n31267) );
  NOR U31502 ( .A(n31209), .B(n31210), .Z(n31216) );
  IV U31503 ( .A(n31210), .Z(n31211) );
  NOR U31504 ( .A(n31212), .B(n31211), .Z(n31213) );
  NOR U31505 ( .A(n31214), .B(n31213), .Z(n31215) );
  NOR U31506 ( .A(n31216), .B(n31215), .Z(n31266) );
  IV U31507 ( .A(n31266), .Z(n31273) );
  XOR U31508 ( .A(n31267), .B(n31273), .Z(n31217) );
  XOR U31509 ( .A(n31276), .B(n31217), .Z(c[120]) );
  NOR U31510 ( .A(n31219), .B(n31218), .Z(n31224) );
  IV U31511 ( .A(n31220), .Z(n31221) );
  NOR U31512 ( .A(n31222), .B(n31221), .Z(n31223) );
  NOR U31513 ( .A(n31224), .B(n31223), .Z(n31284) );
  NOR U31514 ( .A(n165), .B(n159), .Z(n31324) );
  IV U31515 ( .A(n31225), .Z(n31226) );
  NOR U31516 ( .A(n31227), .B(n31226), .Z(n31231) );
  NOR U31517 ( .A(n31229), .B(n31228), .Z(n31230) );
  NOR U31518 ( .A(n31231), .B(n31230), .Z(n31322) );
  IV U31519 ( .A(n31322), .Z(n31256) );
  NOR U31520 ( .A(n163), .B(n160), .Z(n31303) );
  NOR U31521 ( .A(n31233), .B(n31232), .Z(n31238) );
  IV U31522 ( .A(n31234), .Z(n31235) );
  NOR U31523 ( .A(n31236), .B(n31235), .Z(n31237) );
  NOR U31524 ( .A(n31238), .B(n31237), .Z(n31308) );
  NOR U31525 ( .A(n164), .B(n158), .Z(n31316) );
  IV U31526 ( .A(n31239), .Z(n31240) );
  NOR U31527 ( .A(n31241), .B(n31240), .Z(n31246) );
  IV U31528 ( .A(n31242), .Z(n31243) );
  NOR U31529 ( .A(n31244), .B(n31243), .Z(n31245) );
  NOR U31530 ( .A(n31246), .B(n31245), .Z(n31315) );
  NOR U31531 ( .A(n166), .B(n156), .Z(n31313) );
  XOR U31532 ( .A(n31315), .B(n31313), .Z(n31318) );
  XOR U31533 ( .A(n31316), .B(n31318), .Z(n31307) );
  XOR U31534 ( .A(n31308), .B(n31307), .Z(n31247) );
  IV U31535 ( .A(n31247), .Z(n31310) );
  NOR U31536 ( .A(n161), .B(n162), .Z(n31248) );
  IV U31537 ( .A(n31248), .Z(n31309) );
  XOR U31538 ( .A(n31310), .B(n31309), .Z(n31301) );
  NOR U31539 ( .A(n31250), .B(n31249), .Z(n31255) );
  IV U31540 ( .A(n31251), .Z(n31253) );
  NOR U31541 ( .A(n31253), .B(n31252), .Z(n31254) );
  NOR U31542 ( .A(n31255), .B(n31254), .Z(n31299) );
  XOR U31543 ( .A(n31301), .B(n31299), .Z(n31302) );
  XOR U31544 ( .A(n31303), .B(n31302), .Z(n31323) );
  XOR U31545 ( .A(n31256), .B(n31323), .Z(n31326) );
  XOR U31546 ( .A(n31324), .B(n31326), .Z(n31295) );
  IV U31547 ( .A(n31295), .Z(n31265) );
  IV U31548 ( .A(n31257), .Z(n31258) );
  NOR U31549 ( .A(n31259), .B(n31258), .Z(n31264) );
  IV U31550 ( .A(n31260), .Z(n31261) );
  NOR U31551 ( .A(n31262), .B(n31261), .Z(n31263) );
  NOR U31552 ( .A(n31264), .B(n31263), .Z(n31294) );
  NOR U31553 ( .A(n167), .B(n157), .Z(n31292) );
  XOR U31554 ( .A(n31294), .B(n31292), .Z(n31296) );
  XOR U31555 ( .A(n31265), .B(n31296), .Z(n31283) );
  XOR U31556 ( .A(n31284), .B(n31283), .Z(n31285) );
  NOR U31557 ( .A(n31267), .B(n31266), .Z(n31278) );
  IV U31558 ( .A(n31278), .Z(n31272) );
  IV U31559 ( .A(n31268), .Z(n31270) );
  NOR U31560 ( .A(n31270), .B(n31269), .Z(n31277) );
  IV U31561 ( .A(n31277), .Z(n31271) );
  NOR U31562 ( .A(n31272), .B(n31271), .Z(n31289) );
  NOR U31563 ( .A(n31274), .B(n31273), .Z(n31275) );
  NOR U31564 ( .A(n31276), .B(n31275), .Z(n31281) );
  NOR U31565 ( .A(n31278), .B(n31277), .Z(n31279) );
  IV U31566 ( .A(n31279), .Z(n31280) );
  NOR U31567 ( .A(n31281), .B(n31280), .Z(n31286) );
  NOR U31568 ( .A(n31289), .B(n31286), .Z(n31282) );
  XOR U31569 ( .A(n31285), .B(n31282), .Z(c[121]) );
  NOR U31570 ( .A(n31284), .B(n31283), .Z(n31332) );
  IV U31571 ( .A(n31332), .Z(n31330) );
  NOR U31572 ( .A(n31289), .B(n31330), .Z(n31291) );
  IV U31573 ( .A(n31285), .Z(n31287) );
  NOR U31574 ( .A(n31287), .B(n31286), .Z(n31288) );
  NOR U31575 ( .A(n31289), .B(n31288), .Z(n31335) );
  NOR U31576 ( .A(n31332), .B(n31335), .Z(n31290) );
  NOR U31577 ( .A(n31291), .B(n31290), .Z(n31329) );
  IV U31578 ( .A(n31292), .Z(n31293) );
  NOR U31579 ( .A(n31294), .B(n31293), .Z(n31298) );
  NOR U31580 ( .A(n31296), .B(n31295), .Z(n31297) );
  NOR U31581 ( .A(n31298), .B(n31297), .Z(n31338) );
  IV U31582 ( .A(n31299), .Z(n31300) );
  NOR U31583 ( .A(n31301), .B(n31300), .Z(n31305) );
  NOR U31584 ( .A(n31303), .B(n31302), .Z(n31304) );
  NOR U31585 ( .A(n31305), .B(n31304), .Z(n31306) );
  IV U31586 ( .A(n31306), .Z(n31351) );
  NOR U31587 ( .A(n165), .B(n160), .Z(n31348) );
  NOR U31588 ( .A(n163), .B(n162), .Z(n31357) );
  NOR U31589 ( .A(n31308), .B(n31307), .Z(n31312) );
  NOR U31590 ( .A(n31310), .B(n31309), .Z(n31311) );
  NOR U31591 ( .A(n31312), .B(n31311), .Z(n31356) );
  IV U31592 ( .A(n31356), .Z(n31321) );
  NOR U31593 ( .A(n164), .B(n161), .Z(n31365) );
  IV U31594 ( .A(n31313), .Z(n31314) );
  NOR U31595 ( .A(n31315), .B(n31314), .Z(n31320) );
  IV U31596 ( .A(n31316), .Z(n31317) );
  NOR U31597 ( .A(n31318), .B(n31317), .Z(n31319) );
  NOR U31598 ( .A(n31320), .B(n31319), .Z(n31364) );
  NOR U31599 ( .A(n166), .B(n158), .Z(n31362) );
  XOR U31600 ( .A(n31364), .B(n31362), .Z(n31367) );
  XOR U31601 ( .A(n31365), .B(n31367), .Z(n31355) );
  XOR U31602 ( .A(n31321), .B(n31355), .Z(n31359) );
  XOR U31603 ( .A(n31357), .B(n31359), .Z(n31350) );
  XOR U31604 ( .A(n31348), .B(n31350), .Z(n31352) );
  XOR U31605 ( .A(n31351), .B(n31352), .Z(n31342) );
  NOR U31606 ( .A(n31323), .B(n31322), .Z(n31328) );
  IV U31607 ( .A(n31324), .Z(n31325) );
  NOR U31608 ( .A(n31326), .B(n31325), .Z(n31327) );
  NOR U31609 ( .A(n31328), .B(n31327), .Z(n31341) );
  NOR U31610 ( .A(n167), .B(n159), .Z(n31339) );
  XOR U31611 ( .A(n31341), .B(n31339), .Z(n31343) );
  XOR U31612 ( .A(n31342), .B(n31343), .Z(n31337) );
  XOR U31613 ( .A(n31338), .B(n31337), .Z(n31333) );
  IV U31614 ( .A(n31333), .Z(n31331) );
  XOR U31615 ( .A(n31329), .B(n31331), .Z(c[122]) );
  NOR U31616 ( .A(n31331), .B(n31330), .Z(n31336) );
  NOR U31617 ( .A(n31333), .B(n31332), .Z(n31334) );
  NOR U31618 ( .A(n31335), .B(n31334), .Z(n31381) );
  NOR U31619 ( .A(n31336), .B(n31381), .Z(n31375) );
  NOR U31620 ( .A(n31338), .B(n31337), .Z(n31374) );
  IV U31621 ( .A(n31374), .Z(n31383) );
  IV U31622 ( .A(n31339), .Z(n31340) );
  NOR U31623 ( .A(n31341), .B(n31340), .Z(n31346) );
  IV U31624 ( .A(n31342), .Z(n31344) );
  NOR U31625 ( .A(n31344), .B(n31343), .Z(n31345) );
  NOR U31626 ( .A(n31346), .B(n31345), .Z(n31372) );
  NOR U31627 ( .A(n167), .B(n160), .Z(n31347) );
  IV U31628 ( .A(n31347), .Z(n31390) );
  IV U31629 ( .A(n31348), .Z(n31349) );
  NOR U31630 ( .A(n31350), .B(n31349), .Z(n31354) );
  NOR U31631 ( .A(n31352), .B(n31351), .Z(n31353) );
  NOR U31632 ( .A(n31354), .B(n31353), .Z(n31388) );
  NOR U31633 ( .A(n31356), .B(n31355), .Z(n31361) );
  IV U31634 ( .A(n31357), .Z(n31358) );
  NOR U31635 ( .A(n31359), .B(n31358), .Z(n31360) );
  NOR U31636 ( .A(n31361), .B(n31360), .Z(n31395) );
  NOR U31637 ( .A(n164), .B(n163), .Z(n31404) );
  IV U31638 ( .A(n31362), .Z(n31363) );
  NOR U31639 ( .A(n31364), .B(n31363), .Z(n31369) );
  IV U31640 ( .A(n31365), .Z(n31366) );
  NOR U31641 ( .A(n31367), .B(n31366), .Z(n31368) );
  NOR U31642 ( .A(n31369), .B(n31368), .Z(n31403) );
  NOR U31643 ( .A(n166), .B(n161), .Z(n31401) );
  XOR U31644 ( .A(n31403), .B(n31401), .Z(n31406) );
  XOR U31645 ( .A(n31404), .B(n31406), .Z(n31394) );
  XOR U31646 ( .A(n31395), .B(n31394), .Z(n31396) );
  NOR U31647 ( .A(n165), .B(n162), .Z(n31370) );
  IV U31648 ( .A(n31370), .Z(n31397) );
  XOR U31649 ( .A(n31396), .B(n31397), .Z(n31387) );
  XOR U31650 ( .A(n31388), .B(n31387), .Z(n31389) );
  XOR U31651 ( .A(n31390), .B(n31389), .Z(n31371) );
  XOR U31652 ( .A(n31372), .B(n31371), .Z(n31373) );
  XOR U31653 ( .A(n31383), .B(n31373), .Z(n31377) );
  XOR U31654 ( .A(n31375), .B(n31377), .Z(c[123]) );
  NOR U31655 ( .A(n31372), .B(n31371), .Z(n31410) );
  NOR U31656 ( .A(n31374), .B(n31373), .Z(n31379) );
  IV U31657 ( .A(n31375), .Z(n31376) );
  NOR U31658 ( .A(n31377), .B(n31376), .Z(n31378) );
  NOR U31659 ( .A(n31379), .B(n31378), .Z(n31380) );
  IV U31660 ( .A(n31380), .Z(n31411) );
  NOR U31661 ( .A(n31410), .B(n31411), .Z(n31386) );
  IV U31662 ( .A(n31381), .Z(n31382) );
  NOR U31663 ( .A(n31383), .B(n31382), .Z(n31384) );
  IV U31664 ( .A(n31410), .Z(n31414) );
  NOR U31665 ( .A(n31384), .B(n31414), .Z(n31385) );
  NOR U31666 ( .A(n31386), .B(n31385), .Z(n31409) );
  NOR U31667 ( .A(n31388), .B(n31387), .Z(n31393) );
  IV U31668 ( .A(n31389), .Z(n31391) );
  NOR U31669 ( .A(n31391), .B(n31390), .Z(n31392) );
  NOR U31670 ( .A(n31393), .B(n31392), .Z(n31419) );
  NOR U31671 ( .A(n31395), .B(n31394), .Z(n31400) );
  IV U31672 ( .A(n31396), .Z(n31398) );
  NOR U31673 ( .A(n31398), .B(n31397), .Z(n31399) );
  NOR U31674 ( .A(n31400), .B(n31399), .Z(n31422) );
  NOR U31675 ( .A(n167), .B(n162), .Z(n31420) );
  XOR U31676 ( .A(n31422), .B(n31420), .Z(n31424) );
  NOR U31677 ( .A(n164), .B(n165), .Z(n31430) );
  IV U31678 ( .A(n31401), .Z(n31402) );
  NOR U31679 ( .A(n31403), .B(n31402), .Z(n31408) );
  IV U31680 ( .A(n31404), .Z(n31405) );
  NOR U31681 ( .A(n31406), .B(n31405), .Z(n31407) );
  NOR U31682 ( .A(n31408), .B(n31407), .Z(n31429) );
  NOR U31683 ( .A(n166), .B(n163), .Z(n31427) );
  XOR U31684 ( .A(n31429), .B(n31427), .Z(n31432) );
  XOR U31685 ( .A(n31430), .B(n31432), .Z(n31423) );
  XOR U31686 ( .A(n31424), .B(n31423), .Z(n31417) );
  XOR U31687 ( .A(n31419), .B(n31417), .Z(n31413) );
  XOR U31688 ( .A(n31409), .B(n31413), .Z(c[124]) );
  XOR U31689 ( .A(n31410), .B(n31413), .Z(n31412) );
  NOR U31690 ( .A(n31412), .B(n31411), .Z(n31416) );
  NOR U31691 ( .A(n31414), .B(n31413), .Z(n31415) );
  NOR U31692 ( .A(n31416), .B(n31415), .Z(n31439) );
  IV U31693 ( .A(n31417), .Z(n31418) );
  NOR U31694 ( .A(n31419), .B(n31418), .Z(n31442) );
  IV U31695 ( .A(n31420), .Z(n31421) );
  NOR U31696 ( .A(n31422), .B(n31421), .Z(n31426) );
  NOR U31697 ( .A(n31424), .B(n31423), .Z(n31425) );
  NOR U31698 ( .A(n31426), .B(n31425), .Z(n31437) );
  IV U31699 ( .A(n31437), .Z(n31435) );
  NOR U31700 ( .A(n167), .B(n164), .Z(n31453) );
  IV U31701 ( .A(n31427), .Z(n31428) );
  NOR U31702 ( .A(n31429), .B(n31428), .Z(n31434) );
  IV U31703 ( .A(n31430), .Z(n31431) );
  NOR U31704 ( .A(n31432), .B(n31431), .Z(n31433) );
  NOR U31705 ( .A(n31434), .B(n31433), .Z(n31452) );
  NOR U31706 ( .A(n166), .B(n165), .Z(n31450) );
  XOR U31707 ( .A(n31452), .B(n31450), .Z(n31455) );
  XOR U31708 ( .A(n31453), .B(n31455), .Z(n31436) );
  XOR U31709 ( .A(n31435), .B(n31436), .Z(n31443) );
  XOR U31710 ( .A(n31442), .B(n31443), .Z(n31438) );
  XOR U31711 ( .A(n31439), .B(n31438), .Z(c[125]) );
  NOR U31712 ( .A(n31437), .B(n31436), .Z(n31449) );
  IV U31713 ( .A(n31449), .Z(n31441) );
  NOR U31714 ( .A(n31439), .B(n31438), .Z(n31445) );
  IV U31715 ( .A(n31445), .Z(n31440) );
  NOR U31716 ( .A(n31441), .B(n31440), .Z(n31692) );
  IV U31717 ( .A(n31442), .Z(n31444) );
  NOR U31718 ( .A(n31444), .B(n31443), .Z(n31446) );
  NOR U31719 ( .A(n31446), .B(n31445), .Z(n31447) );
  IV U31720 ( .A(n31447), .Z(n31448) );
  NOR U31721 ( .A(n31449), .B(n31448), .Z(n31690) );
  NOR U31722 ( .A(n31692), .B(n31690), .Z(n31459) );
  IV U31723 ( .A(n31450), .Z(n31451) );
  NOR U31724 ( .A(n31452), .B(n31451), .Z(n31457) );
  IV U31725 ( .A(n31453), .Z(n31454) );
  NOR U31726 ( .A(n31455), .B(n31454), .Z(n31456) );
  NOR U31727 ( .A(n31457), .B(n31456), .Z(n31694) );
  NOR U31728 ( .A(n166), .B(n167), .Z(n31458) );
  XOR U31729 ( .A(n31694), .B(n31458), .Z(n31689) );
  XOR U31730 ( .A(n31459), .B(n31689), .Z(n31460) );
  IV U31731 ( .A(n31460), .Z(c[126]) );
  XOR U31732 ( .A(n31462), .B(n31461), .Z(c[65]) );
  NOR U31733 ( .A(n31464), .B(n31463), .Z(n31466) );
  XOR U31734 ( .A(n31466), .B(n31465), .Z(c[66]) );
  NOR U31735 ( .A(n31466), .B(n31465), .Z(n31467) );
  NOR U31736 ( .A(n31468), .B(n31467), .Z(n31470) );
  XOR U31737 ( .A(n31470), .B(n31469), .Z(c[67]) );
  NOR U31738 ( .A(n31470), .B(n31469), .Z(n31471) );
  IV U31739 ( .A(n31471), .Z(n31475) );
  XOR U31740 ( .A(n31473), .B(n31472), .Z(n31474) );
  XOR U31741 ( .A(n31475), .B(n31474), .Z(c[68]) );
  NOR U31742 ( .A(n31475), .B(n31474), .Z(n31480) );
  NOR U31743 ( .A(n31477), .B(n31476), .Z(n31478) );
  IV U31744 ( .A(n31478), .Z(n31479) );
  NOR U31745 ( .A(n31480), .B(n31479), .Z(n31482) );
  XOR U31746 ( .A(n31482), .B(n31481), .Z(c[69]) );
  XOR U31747 ( .A(n31484), .B(n31483), .Z(n31485) );
  XOR U31748 ( .A(n31486), .B(n31485), .Z(c[70]) );
  NOR U31749 ( .A(n31486), .B(n31485), .Z(n31489) );
  NOR U31750 ( .A(n31487), .B(n31489), .Z(n31496) );
  XOR U31751 ( .A(n31494), .B(n31488), .Z(n31495) );
  XOR U31752 ( .A(n31496), .B(n31495), .Z(c[71]) );
  IV U31753 ( .A(n31489), .Z(n31490) );
  NOR U31754 ( .A(n31491), .B(n31490), .Z(n31492) );
  IV U31755 ( .A(n31492), .Z(n31493) );
  NOR U31756 ( .A(n31494), .B(n31493), .Z(n31505) );
  NOR U31757 ( .A(n31496), .B(n31495), .Z(n31497) );
  NOR U31758 ( .A(n31498), .B(n31497), .Z(n31499) );
  IV U31759 ( .A(n31499), .Z(n31500) );
  NOR U31760 ( .A(n31501), .B(n31500), .Z(n31509) );
  NOR U31761 ( .A(n31505), .B(n31509), .Z(n31502) );
  XOR U31762 ( .A(n31503), .B(n31502), .Z(c[72]) );
  XOR U31763 ( .A(n31505), .B(n31504), .Z(n31511) );
  XOR U31764 ( .A(n31507), .B(n31506), .Z(n31508) );
  NOR U31765 ( .A(n31509), .B(n31508), .Z(n31510) );
  NOR U31766 ( .A(n31511), .B(n31510), .Z(n31512) );
  XOR U31767 ( .A(n31513), .B(n31512), .Z(c[73]) );
  XOR U31768 ( .A(n31515), .B(n31514), .Z(n31516) );
  XOR U31769 ( .A(n31517), .B(n31516), .Z(c[74]) );
  NOR U31770 ( .A(n31517), .B(n31516), .Z(n31518) );
  NOR U31771 ( .A(n31519), .B(n31518), .Z(n31522) );
  XOR U31772 ( .A(n31524), .B(n31523), .Z(n31521) );
  XOR U31773 ( .A(n31522), .B(n31521), .Z(c[75]) );
  IV U31774 ( .A(n31520), .Z(n31532) );
  NOR U31775 ( .A(n31522), .B(n31521), .Z(n31528) );
  IV U31776 ( .A(n31528), .Z(n31531) );
  XOR U31777 ( .A(n31532), .B(n31531), .Z(n31530) );
  IV U31778 ( .A(n31523), .Z(n31525) );
  NOR U31779 ( .A(n31525), .B(n31524), .Z(n31526) );
  IV U31780 ( .A(n31526), .Z(n31527) );
  NOR U31781 ( .A(n31528), .B(n31527), .Z(n31529) );
  NOR U31782 ( .A(n31530), .B(n31529), .Z(n31533) );
  XOR U31783 ( .A(n31534), .B(n31533), .Z(c[76]) );
  NOR U31784 ( .A(n31532), .B(n31531), .Z(n31536) );
  NOR U31785 ( .A(n31534), .B(n31533), .Z(n31535) );
  NOR U31786 ( .A(n31536), .B(n31535), .Z(n31540) );
  XOR U31787 ( .A(n31538), .B(n31537), .Z(n31539) );
  XOR U31788 ( .A(n31540), .B(n31539), .Z(c[77]) );
  XOR U31789 ( .A(n31542), .B(n31541), .Z(c[78]) );
  XOR U31790 ( .A(n31544), .B(n31543), .Z(c[79]) );
  IV U31791 ( .A(n31545), .Z(n31550) );
  XOR U31792 ( .A(n31550), .B(n31546), .Z(c[80]) );
  NOR U31793 ( .A(n31548), .B(n31547), .Z(n31554) );
  NOR U31794 ( .A(n31550), .B(n31549), .Z(n31551) );
  NOR U31795 ( .A(n31552), .B(n31551), .Z(n31553) );
  NOR U31796 ( .A(n31554), .B(n31553), .Z(n31556) );
  XOR U31797 ( .A(n31556), .B(n31555), .Z(c[81]) );
  XOR U31798 ( .A(n31558), .B(n31557), .Z(n31559) );
  XOR U31799 ( .A(n31560), .B(n31559), .Z(c[82]) );
  NOR U31800 ( .A(n31562), .B(n31561), .Z(n31565) );
  XOR U31801 ( .A(n31575), .B(n31563), .Z(n31564) );
  XOR U31802 ( .A(n31565), .B(n31564), .Z(c[83]) );
  NOR U31803 ( .A(n31565), .B(n31564), .Z(n31566) );
  NOR U31804 ( .A(n31567), .B(n31566), .Z(n31568) );
  IV U31805 ( .A(n31568), .Z(n31569) );
  NOR U31806 ( .A(n31570), .B(n31569), .Z(n31583) );
  NOR U31807 ( .A(n31572), .B(n31571), .Z(n31573) );
  IV U31808 ( .A(n31573), .Z(n31574) );
  NOR U31809 ( .A(n31575), .B(n31574), .Z(n31579) );
  NOR U31810 ( .A(n31583), .B(n31579), .Z(n31576) );
  XOR U31811 ( .A(n31577), .B(n31576), .Z(c[84]) );
  XOR U31812 ( .A(n31579), .B(n31578), .Z(n31585) );
  XOR U31813 ( .A(n31581), .B(n31580), .Z(n31582) );
  NOR U31814 ( .A(n31583), .B(n31582), .Z(n31584) );
  NOR U31815 ( .A(n31585), .B(n31584), .Z(n31586) );
  XOR U31816 ( .A(n31587), .B(n31586), .Z(c[85]) );
  XOR U31817 ( .A(n31589), .B(n31588), .Z(n31590) );
  XOR U31818 ( .A(n31591), .B(n31590), .Z(c[86]) );
  NOR U31819 ( .A(n31591), .B(n31590), .Z(n31592) );
  NOR U31820 ( .A(n31593), .B(n31592), .Z(n31597) );
  IV U31821 ( .A(n31594), .Z(n31596) );
  XOR U31822 ( .A(n31596), .B(n31595), .Z(n31598) );
  XOR U31823 ( .A(n31597), .B(n31598), .Z(c[87]) );
  IV U31824 ( .A(n31597), .Z(n31599) );
  NOR U31825 ( .A(n31599), .B(n31598), .Z(n31600) );
  NOR U31826 ( .A(n31601), .B(n31600), .Z(n31609) );
  XOR U31827 ( .A(n31610), .B(n31602), .Z(n31603) );
  XOR U31828 ( .A(n31609), .B(n31603), .Z(c[88]) );
  IV U31829 ( .A(n31610), .Z(n31605) );
  IV U31830 ( .A(n31609), .Z(n31604) );
  NOR U31831 ( .A(n31605), .B(n31604), .Z(n31608) );
  IV U31832 ( .A(n31606), .Z(n31607) );
  NOR U31833 ( .A(n31608), .B(n31607), .Z(n31615) );
  XOR U31834 ( .A(n31609), .B(n31611), .Z(n31613) );
  XOR U31835 ( .A(n31611), .B(n31610), .Z(n31612) );
  NOR U31836 ( .A(n31613), .B(n31612), .Z(n31614) );
  NOR U31837 ( .A(n31615), .B(n31614), .Z(n31616) );
  XOR U31838 ( .A(n31617), .B(n31616), .Z(c[89]) );
  XOR U31839 ( .A(n31631), .B(n31618), .Z(n31619) );
  XOR U31840 ( .A(n31622), .B(n31619), .Z(c[90]) );
  NOR U31841 ( .A(n31631), .B(n31628), .Z(n31620) );
  XOR U31842 ( .A(n31626), .B(n31620), .Z(n31625) );
  XOR U31843 ( .A(n31621), .B(n31628), .Z(n31623) );
  NOR U31844 ( .A(n31623), .B(n31622), .Z(n31624) );
  NOR U31845 ( .A(n31625), .B(n31624), .Z(n31632) );
  XOR U31846 ( .A(n31633), .B(n31632), .Z(c[91]) );
  IV U31847 ( .A(n31626), .Z(n31627) );
  NOR U31848 ( .A(n31628), .B(n31627), .Z(n31629) );
  IV U31849 ( .A(n31629), .Z(n31630) );
  NOR U31850 ( .A(n31631), .B(n31630), .Z(n31635) );
  NOR U31851 ( .A(n31633), .B(n31632), .Z(n31634) );
  NOR U31852 ( .A(n31635), .B(n31634), .Z(n31639) );
  XOR U31853 ( .A(n31637), .B(n31636), .Z(n31638) );
  XOR U31854 ( .A(n31639), .B(n31638), .Z(c[92]) );
  NOR U31855 ( .A(n31639), .B(n31638), .Z(n31640) );
  NOR U31856 ( .A(n31641), .B(n31640), .Z(n31642) );
  XOR U31857 ( .A(n31643), .B(n31642), .Z(n31644) );
  XOR U31858 ( .A(n31645), .B(n31644), .Z(c[93]) );
  XOR U31859 ( .A(n31650), .B(n31646), .Z(c[94]) );
  NOR U31860 ( .A(n31648), .B(n31647), .Z(n31654) );
  NOR U31861 ( .A(n31650), .B(n31649), .Z(n31651) );
  NOR U31862 ( .A(n31652), .B(n31651), .Z(n31653) );
  NOR U31863 ( .A(n31654), .B(n31653), .Z(n31656) );
  XOR U31864 ( .A(n31656), .B(n31655), .Z(c[95]) );
  XOR U31865 ( .A(n31658), .B(n31657), .Z(c[96]) );
  XOR U31866 ( .A(n31660), .B(n31659), .Z(c[97]) );
  XOR U31867 ( .A(n31669), .B(n31661), .Z(n31662) );
  XOR U31868 ( .A(n31663), .B(n31662), .Z(c[98]) );
  IV U31869 ( .A(n31664), .Z(n31666) );
  NOR U31870 ( .A(n31666), .B(n31665), .Z(n31667) );
  IV U31871 ( .A(n31667), .Z(n31668) );
  NOR U31872 ( .A(n31669), .B(n31668), .Z(n31678) );
  IV U31873 ( .A(n31670), .Z(n31671) );
  NOR U31874 ( .A(n31672), .B(n31671), .Z(n31673) );
  NOR U31875 ( .A(n31678), .B(n31673), .Z(n31674) );
  IV U31876 ( .A(n31674), .Z(n31675) );
  XOR U31877 ( .A(n31676), .B(n31675), .Z(c[99]) );
  NOR U31878 ( .A(n31676), .B(n31675), .Z(n31677) );
  NOR U31879 ( .A(n31678), .B(n31677), .Z(n31682) );
  XOR U31880 ( .A(n31680), .B(n31679), .Z(n31681) );
  XOR U31881 ( .A(n31682), .B(n31681), .Z(c[100]) );
  NOR U31882 ( .A(n31682), .B(n31681), .Z(n31683) );
  NOR U31883 ( .A(n31684), .B(n31683), .Z(n31688) );
  XOR U31884 ( .A(n31686), .B(n31685), .Z(n31687) );
  XOR U31885 ( .A(n31688), .B(n31687), .Z(c[101]) );
  NOR U31886 ( .A(n31690), .B(n31689), .Z(n31691) );
  NOR U31887 ( .A(n31692), .B(n31691), .Z(n31693) );
  IV U31888 ( .A(n31693), .Z(n31696) );
  NOR U31889 ( .A(n31694), .B(n167), .Z(n31695) );
  XOR U31890 ( .A(n31696), .B(n31695), .Z(c[127]) );
  XOR U31891 ( .A(n31698), .B(n31697), .Z(c[2]) );
  XOR U31892 ( .A(n31700), .B(n31699), .Z(c[12]) );
  XOR U31893 ( .A(n31702), .B(n31701), .Z(c[13]) );
  XOR U31894 ( .A(n31704), .B(n31703), .Z(c[14]) );
  XOR U31895 ( .A(n31706), .B(n31705), .Z(c[15]) );
  XOR U31896 ( .A(n31708), .B(n31707), .Z(c[16]) );
  XOR U31897 ( .A(n31710), .B(n31709), .Z(c[17]) );
  XOR U31898 ( .A(n31712), .B(n31711), .Z(c[18]) );
  XOR U31899 ( .A(n31714), .B(n31713), .Z(c[19]) );
  XOR U31900 ( .A(n31716), .B(n31715), .Z(c[20]) );
  XOR U31901 ( .A(n31718), .B(n31717), .Z(c[21]) );
  XOR U31902 ( .A(n31720), .B(n31719), .Z(c[3]) );
  XOR U31903 ( .A(n31722), .B(n31721), .Z(c[22]) );
  XOR U31904 ( .A(n31724), .B(n31723), .Z(c[23]) );
  XOR U31905 ( .A(n31726), .B(n31725), .Z(c[24]) );
  XOR U31906 ( .A(n31728), .B(n31727), .Z(c[25]) );
  XOR U31907 ( .A(n31730), .B(n31729), .Z(c[26]) );
  XOR U31908 ( .A(n31732), .B(n31731), .Z(c[27]) );
  XOR U31909 ( .A(n31734), .B(n31733), .Z(c[28]) );
  XOR U31910 ( .A(n31736), .B(n31735), .Z(c[29]) );
  XOR U31911 ( .A(n31738), .B(n31737), .Z(c[30]) );
  XOR U31912 ( .A(n31740), .B(n31739), .Z(c[31]) );
  XOR U31913 ( .A(n31742), .B(n31741), .Z(c[4]) );
  XOR U31914 ( .A(n31744), .B(n31743), .Z(c[32]) );
  XOR U31915 ( .A(n31746), .B(n31745), .Z(c[33]) );
  XOR U31916 ( .A(n31748), .B(n31747), .Z(c[34]) );
  XOR U31917 ( .A(n31750), .B(n31749), .Z(c[35]) );
  XOR U31918 ( .A(n31752), .B(n31751), .Z(c[36]) );
  XOR U31919 ( .A(n31754), .B(n31753), .Z(c[37]) );
  XOR U31920 ( .A(n31756), .B(n31755), .Z(c[38]) );
  XOR U31921 ( .A(n31758), .B(n31757), .Z(c[39]) );
  XOR U31922 ( .A(n31760), .B(n31759), .Z(c[40]) );
  XOR U31923 ( .A(n31762), .B(n31761), .Z(c[41]) );
  XOR U31924 ( .A(n31764), .B(n31763), .Z(c[5]) );
  XOR U31925 ( .A(n31766), .B(n31765), .Z(c[42]) );
  XOR U31926 ( .A(n31768), .B(n31767), .Z(c[43]) );
  XOR U31927 ( .A(n31770), .B(n31769), .Z(c[44]) );
  XOR U31928 ( .A(n31772), .B(n31771), .Z(c[45]) );
  IV U31929 ( .A(n31773), .Z(n31775) );
  XOR U31930 ( .A(n31775), .B(n31774), .Z(c[46]) );
  XOR U31931 ( .A(n31777), .B(n31776), .Z(c[47]) );
  XOR U31932 ( .A(n31779), .B(n31778), .Z(c[48]) );
  XOR U31933 ( .A(n31781), .B(n31780), .Z(c[49]) );
  XOR U31934 ( .A(n31783), .B(n31782), .Z(c[50]) );
  XOR U31935 ( .A(n31785), .B(n31784), .Z(c[51]) );
  XOR U31936 ( .A(n31787), .B(n31786), .Z(c[6]) );
  XOR U31937 ( .A(n31789), .B(n31788), .Z(c[52]) );
  XOR U31938 ( .A(n31791), .B(n31790), .Z(c[53]) );
  XOR U31939 ( .A(n31793), .B(n31792), .Z(c[54]) );
  XOR U31940 ( .A(n31795), .B(n31794), .Z(c[55]) );
  XOR U31941 ( .A(n31797), .B(n31796), .Z(c[56]) );
  XOR U31942 ( .A(n31799), .B(n31798), .Z(n31800) );
  XOR U31943 ( .A(n31801), .B(n31800), .Z(c[57]) );
  XOR U31944 ( .A(n31803), .B(n31802), .Z(c[58]) );
  XOR U31945 ( .A(n31805), .B(n31804), .Z(n31806) );
  XOR U31946 ( .A(n31807), .B(n31806), .Z(c[59]) );
  XOR U31947 ( .A(n31809), .B(n31808), .Z(c[60]) );
  XOR U31948 ( .A(n31811), .B(n31810), .Z(c[61]) );
  XOR U31949 ( .A(n31813), .B(n31812), .Z(c[7]) );
  XOR U31950 ( .A(n31815), .B(n31814), .Z(n31816) );
  XOR U31951 ( .A(n31817), .B(n31816), .Z(c[62]) );
  XOR U31952 ( .A(n31819), .B(n31818), .Z(c[63]) );
  XOR U31953 ( .A(n31821), .B(n31820), .Z(c[64]) );
  XOR U31954 ( .A(n31823), .B(n31822), .Z(c[8]) );
  XOR U31955 ( .A(n31825), .B(n31824), .Z(c[9]) );
  XOR U31956 ( .A(n31827), .B(n31826), .Z(c[10]) );
  XOR U31957 ( .A(n31829), .B(n31828), .Z(c[11]) );
  NOR U31958 ( .A(n169), .B(n168), .Z(n31830) );
  XOR U31959 ( .A(n31831), .B(n31830), .Z(c[1]) );
endmodule

