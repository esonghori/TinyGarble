
module modexp_2N_NN_N1024_CC2097152 ( clk, rst, g_init, e_init, g_input, 
        e_input, o );
  input [1023:0] g_init;
  input [1023:0] e_init;
  input [1023:0] g_input;
  input [1023:0] e_input;
  output [1023:0] o;
  input clk, rst;
  wire   first_one, mul_pow, n6, n8, \modmult_1/xin[1023] ,
         \modmult_1/xin[1022] , \modmult_1/xin[1021] , \modmult_1/xin[1020] ,
         \modmult_1/xin[1019] , \modmult_1/xin[1018] , \modmult_1/xin[1017] ,
         \modmult_1/xin[1016] , \modmult_1/xin[1015] , \modmult_1/xin[1014] ,
         \modmult_1/xin[1013] , \modmult_1/xin[1012] , \modmult_1/xin[1011] ,
         \modmult_1/xin[1010] , \modmult_1/xin[1009] , \modmult_1/xin[1008] ,
         \modmult_1/xin[1007] , \modmult_1/xin[1006] , \modmult_1/xin[1005] ,
         \modmult_1/xin[1004] , \modmult_1/xin[1003] , \modmult_1/xin[1002] ,
         \modmult_1/xin[1001] , \modmult_1/xin[1000] , \modmult_1/xin[999] ,
         \modmult_1/xin[998] , \modmult_1/xin[997] , \modmult_1/xin[996] ,
         \modmult_1/xin[995] , \modmult_1/xin[994] , \modmult_1/xin[993] ,
         \modmult_1/xin[992] , \modmult_1/xin[991] , \modmult_1/xin[990] ,
         \modmult_1/xin[989] , \modmult_1/xin[988] , \modmult_1/xin[987] ,
         \modmult_1/xin[986] , \modmult_1/xin[985] , \modmult_1/xin[984] ,
         \modmult_1/xin[983] , \modmult_1/xin[982] , \modmult_1/xin[981] ,
         \modmult_1/xin[980] , \modmult_1/xin[979] , \modmult_1/xin[978] ,
         \modmult_1/xin[977] , \modmult_1/xin[976] , \modmult_1/xin[975] ,
         \modmult_1/xin[974] , \modmult_1/xin[973] , \modmult_1/xin[972] ,
         \modmult_1/xin[971] , \modmult_1/xin[970] , \modmult_1/xin[969] ,
         \modmult_1/xin[968] , \modmult_1/xin[967] , \modmult_1/xin[966] ,
         \modmult_1/xin[965] , \modmult_1/xin[964] , \modmult_1/xin[963] ,
         \modmult_1/xin[962] , \modmult_1/xin[961] , \modmult_1/xin[960] ,
         \modmult_1/xin[959] , \modmult_1/xin[958] , \modmult_1/xin[957] ,
         \modmult_1/xin[956] , \modmult_1/xin[955] , \modmult_1/xin[954] ,
         \modmult_1/xin[953] , \modmult_1/xin[952] , \modmult_1/xin[951] ,
         \modmult_1/xin[950] , \modmult_1/xin[949] , \modmult_1/xin[948] ,
         \modmult_1/xin[947] , \modmult_1/xin[946] , \modmult_1/xin[945] ,
         \modmult_1/xin[944] , \modmult_1/xin[943] , \modmult_1/xin[942] ,
         \modmult_1/xin[941] , \modmult_1/xin[940] , \modmult_1/xin[939] ,
         \modmult_1/xin[938] , \modmult_1/xin[937] , \modmult_1/xin[936] ,
         \modmult_1/xin[935] , \modmult_1/xin[934] , \modmult_1/xin[933] ,
         \modmult_1/xin[932] , \modmult_1/xin[931] , \modmult_1/xin[930] ,
         \modmult_1/xin[929] , \modmult_1/xin[928] , \modmult_1/xin[927] ,
         \modmult_1/xin[926] , \modmult_1/xin[925] , \modmult_1/xin[924] ,
         \modmult_1/xin[923] , \modmult_1/xin[922] , \modmult_1/xin[921] ,
         \modmult_1/xin[920] , \modmult_1/xin[919] , \modmult_1/xin[918] ,
         \modmult_1/xin[917] , \modmult_1/xin[916] , \modmult_1/xin[915] ,
         \modmult_1/xin[914] , \modmult_1/xin[913] , \modmult_1/xin[912] ,
         \modmult_1/xin[911] , \modmult_1/xin[910] , \modmult_1/xin[909] ,
         \modmult_1/xin[908] , \modmult_1/xin[907] , \modmult_1/xin[906] ,
         \modmult_1/xin[905] , \modmult_1/xin[904] , \modmult_1/xin[903] ,
         \modmult_1/xin[902] , \modmult_1/xin[901] , \modmult_1/xin[900] ,
         \modmult_1/xin[899] , \modmult_1/xin[898] , \modmult_1/xin[897] ,
         \modmult_1/xin[896] , \modmult_1/xin[895] , \modmult_1/xin[894] ,
         \modmult_1/xin[893] , \modmult_1/xin[892] , \modmult_1/xin[891] ,
         \modmult_1/xin[890] , \modmult_1/xin[889] , \modmult_1/xin[888] ,
         \modmult_1/xin[887] , \modmult_1/xin[886] , \modmult_1/xin[885] ,
         \modmult_1/xin[884] , \modmult_1/xin[883] , \modmult_1/xin[882] ,
         \modmult_1/xin[881] , \modmult_1/xin[880] , \modmult_1/xin[879] ,
         \modmult_1/xin[878] , \modmult_1/xin[877] , \modmult_1/xin[876] ,
         \modmult_1/xin[875] , \modmult_1/xin[874] , \modmult_1/xin[873] ,
         \modmult_1/xin[872] , \modmult_1/xin[871] , \modmult_1/xin[870] ,
         \modmult_1/xin[869] , \modmult_1/xin[868] , \modmult_1/xin[867] ,
         \modmult_1/xin[866] , \modmult_1/xin[865] , \modmult_1/xin[864] ,
         \modmult_1/xin[863] , \modmult_1/xin[862] , \modmult_1/xin[861] ,
         \modmult_1/xin[860] , \modmult_1/xin[859] , \modmult_1/xin[858] ,
         \modmult_1/xin[857] , \modmult_1/xin[856] , \modmult_1/xin[855] ,
         \modmult_1/xin[854] , \modmult_1/xin[853] , \modmult_1/xin[852] ,
         \modmult_1/xin[851] , \modmult_1/xin[850] , \modmult_1/xin[849] ,
         \modmult_1/xin[848] , \modmult_1/xin[847] , \modmult_1/xin[846] ,
         \modmult_1/xin[845] , \modmult_1/xin[844] , \modmult_1/xin[843] ,
         \modmult_1/xin[842] , \modmult_1/xin[841] , \modmult_1/xin[840] ,
         \modmult_1/xin[839] , \modmult_1/xin[838] , \modmult_1/xin[837] ,
         \modmult_1/xin[836] , \modmult_1/xin[835] , \modmult_1/xin[834] ,
         \modmult_1/xin[833] , \modmult_1/xin[832] , \modmult_1/xin[831] ,
         \modmult_1/xin[830] , \modmult_1/xin[829] , \modmult_1/xin[828] ,
         \modmult_1/xin[827] , \modmult_1/xin[826] , \modmult_1/xin[825] ,
         \modmult_1/xin[824] , \modmult_1/xin[823] , \modmult_1/xin[822] ,
         \modmult_1/xin[821] , \modmult_1/xin[820] , \modmult_1/xin[819] ,
         \modmult_1/xin[818] , \modmult_1/xin[817] , \modmult_1/xin[816] ,
         \modmult_1/xin[815] , \modmult_1/xin[814] , \modmult_1/xin[813] ,
         \modmult_1/xin[812] , \modmult_1/xin[811] , \modmult_1/xin[810] ,
         \modmult_1/xin[809] , \modmult_1/xin[808] , \modmult_1/xin[807] ,
         \modmult_1/xin[806] , \modmult_1/xin[805] , \modmult_1/xin[804] ,
         \modmult_1/xin[803] , \modmult_1/xin[802] , \modmult_1/xin[801] ,
         \modmult_1/xin[800] , \modmult_1/xin[799] , \modmult_1/xin[798] ,
         \modmult_1/xin[797] , \modmult_1/xin[796] , \modmult_1/xin[795] ,
         \modmult_1/xin[794] , \modmult_1/xin[793] , \modmult_1/xin[792] ,
         \modmult_1/xin[791] , \modmult_1/xin[790] , \modmult_1/xin[789] ,
         \modmult_1/xin[788] , \modmult_1/xin[787] , \modmult_1/xin[786] ,
         \modmult_1/xin[785] , \modmult_1/xin[784] , \modmult_1/xin[783] ,
         \modmult_1/xin[782] , \modmult_1/xin[781] , \modmult_1/xin[780] ,
         \modmult_1/xin[779] , \modmult_1/xin[778] , \modmult_1/xin[777] ,
         \modmult_1/xin[776] , \modmult_1/xin[775] , \modmult_1/xin[774] ,
         \modmult_1/xin[773] , \modmult_1/xin[772] , \modmult_1/xin[771] ,
         \modmult_1/xin[770] , \modmult_1/xin[769] , \modmult_1/xin[768] ,
         \modmult_1/xin[767] , \modmult_1/xin[766] , \modmult_1/xin[765] ,
         \modmult_1/xin[764] , \modmult_1/xin[763] , \modmult_1/xin[762] ,
         \modmult_1/xin[761] , \modmult_1/xin[760] , \modmult_1/xin[759] ,
         \modmult_1/xin[758] , \modmult_1/xin[757] , \modmult_1/xin[756] ,
         \modmult_1/xin[755] , \modmult_1/xin[754] , \modmult_1/xin[753] ,
         \modmult_1/xin[752] , \modmult_1/xin[751] , \modmult_1/xin[750] ,
         \modmult_1/xin[749] , \modmult_1/xin[748] , \modmult_1/xin[747] ,
         \modmult_1/xin[746] , \modmult_1/xin[745] , \modmult_1/xin[744] ,
         \modmult_1/xin[743] , \modmult_1/xin[742] , \modmult_1/xin[741] ,
         \modmult_1/xin[740] , \modmult_1/xin[739] , \modmult_1/xin[738] ,
         \modmult_1/xin[737] , \modmult_1/xin[736] , \modmult_1/xin[735] ,
         \modmult_1/xin[734] , \modmult_1/xin[733] , \modmult_1/xin[732] ,
         \modmult_1/xin[731] , \modmult_1/xin[730] , \modmult_1/xin[729] ,
         \modmult_1/xin[728] , \modmult_1/xin[727] , \modmult_1/xin[726] ,
         \modmult_1/xin[725] , \modmult_1/xin[724] , \modmult_1/xin[723] ,
         \modmult_1/xin[722] , \modmult_1/xin[721] , \modmult_1/xin[720] ,
         \modmult_1/xin[719] , \modmult_1/xin[718] , \modmult_1/xin[717] ,
         \modmult_1/xin[716] , \modmult_1/xin[715] , \modmult_1/xin[714] ,
         \modmult_1/xin[713] , \modmult_1/xin[712] , \modmult_1/xin[711] ,
         \modmult_1/xin[710] , \modmult_1/xin[709] , \modmult_1/xin[708] ,
         \modmult_1/xin[707] , \modmult_1/xin[706] , \modmult_1/xin[705] ,
         \modmult_1/xin[704] , \modmult_1/xin[703] , \modmult_1/xin[702] ,
         \modmult_1/xin[701] , \modmult_1/xin[700] , \modmult_1/xin[699] ,
         \modmult_1/xin[698] , \modmult_1/xin[697] , \modmult_1/xin[696] ,
         \modmult_1/xin[695] , \modmult_1/xin[694] , \modmult_1/xin[693] ,
         \modmult_1/xin[692] , \modmult_1/xin[691] , \modmult_1/xin[690] ,
         \modmult_1/xin[689] , \modmult_1/xin[688] , \modmult_1/xin[687] ,
         \modmult_1/xin[686] , \modmult_1/xin[685] , \modmult_1/xin[684] ,
         \modmult_1/xin[683] , \modmult_1/xin[682] , \modmult_1/xin[681] ,
         \modmult_1/xin[680] , \modmult_1/xin[679] , \modmult_1/xin[678] ,
         \modmult_1/xin[677] , \modmult_1/xin[676] , \modmult_1/xin[675] ,
         \modmult_1/xin[674] , \modmult_1/xin[673] , \modmult_1/xin[672] ,
         \modmult_1/xin[671] , \modmult_1/xin[670] , \modmult_1/xin[669] ,
         \modmult_1/xin[668] , \modmult_1/xin[667] , \modmult_1/xin[666] ,
         \modmult_1/xin[665] , \modmult_1/xin[664] , \modmult_1/xin[663] ,
         \modmult_1/xin[662] , \modmult_1/xin[661] , \modmult_1/xin[660] ,
         \modmult_1/xin[659] , \modmult_1/xin[658] , \modmult_1/xin[657] ,
         \modmult_1/xin[656] , \modmult_1/xin[655] , \modmult_1/xin[654] ,
         \modmult_1/xin[653] , \modmult_1/xin[652] , \modmult_1/xin[651] ,
         \modmult_1/xin[650] , \modmult_1/xin[649] , \modmult_1/xin[648] ,
         \modmult_1/xin[647] , \modmult_1/xin[646] , \modmult_1/xin[645] ,
         \modmult_1/xin[644] , \modmult_1/xin[643] , \modmult_1/xin[642] ,
         \modmult_1/xin[641] , \modmult_1/xin[640] , \modmult_1/xin[639] ,
         \modmult_1/xin[638] , \modmult_1/xin[637] , \modmult_1/xin[636] ,
         \modmult_1/xin[635] , \modmult_1/xin[634] , \modmult_1/xin[633] ,
         \modmult_1/xin[632] , \modmult_1/xin[631] , \modmult_1/xin[630] ,
         \modmult_1/xin[629] , \modmult_1/xin[628] , \modmult_1/xin[627] ,
         \modmult_1/xin[626] , \modmult_1/xin[625] , \modmult_1/xin[624] ,
         \modmult_1/xin[623] , \modmult_1/xin[622] , \modmult_1/xin[621] ,
         \modmult_1/xin[620] , \modmult_1/xin[619] , \modmult_1/xin[618] ,
         \modmult_1/xin[617] , \modmult_1/xin[616] , \modmult_1/xin[615] ,
         \modmult_1/xin[614] , \modmult_1/xin[613] , \modmult_1/xin[612] ,
         \modmult_1/xin[611] , \modmult_1/xin[610] , \modmult_1/xin[609] ,
         \modmult_1/xin[608] , \modmult_1/xin[607] , \modmult_1/xin[606] ,
         \modmult_1/xin[605] , \modmult_1/xin[604] , \modmult_1/xin[603] ,
         \modmult_1/xin[602] , \modmult_1/xin[601] , \modmult_1/xin[600] ,
         \modmult_1/xin[599] , \modmult_1/xin[598] , \modmult_1/xin[597] ,
         \modmult_1/xin[596] , \modmult_1/xin[595] , \modmult_1/xin[594] ,
         \modmult_1/xin[593] , \modmult_1/xin[592] , \modmult_1/xin[591] ,
         \modmult_1/xin[590] , \modmult_1/xin[589] , \modmult_1/xin[588] ,
         \modmult_1/xin[587] , \modmult_1/xin[586] , \modmult_1/xin[585] ,
         \modmult_1/xin[584] , \modmult_1/xin[583] , \modmult_1/xin[582] ,
         \modmult_1/xin[581] , \modmult_1/xin[580] , \modmult_1/xin[579] ,
         \modmult_1/xin[578] , \modmult_1/xin[577] , \modmult_1/xin[576] ,
         \modmult_1/xin[575] , \modmult_1/xin[574] , \modmult_1/xin[573] ,
         \modmult_1/xin[572] , \modmult_1/xin[571] , \modmult_1/xin[570] ,
         \modmult_1/xin[569] , \modmult_1/xin[568] , \modmult_1/xin[567] ,
         \modmult_1/xin[566] , \modmult_1/xin[565] , \modmult_1/xin[564] ,
         \modmult_1/xin[563] , \modmult_1/xin[562] , \modmult_1/xin[561] ,
         \modmult_1/xin[560] , \modmult_1/xin[559] , \modmult_1/xin[558] ,
         \modmult_1/xin[557] , \modmult_1/xin[556] , \modmult_1/xin[555] ,
         \modmult_1/xin[554] , \modmult_1/xin[553] , \modmult_1/xin[552] ,
         \modmult_1/xin[551] , \modmult_1/xin[550] , \modmult_1/xin[549] ,
         \modmult_1/xin[548] , \modmult_1/xin[547] , \modmult_1/xin[546] ,
         \modmult_1/xin[545] , \modmult_1/xin[544] , \modmult_1/xin[543] ,
         \modmult_1/xin[542] , \modmult_1/xin[541] , \modmult_1/xin[540] ,
         \modmult_1/xin[539] , \modmult_1/xin[538] , \modmult_1/xin[537] ,
         \modmult_1/xin[536] , \modmult_1/xin[535] , \modmult_1/xin[534] ,
         \modmult_1/xin[533] , \modmult_1/xin[532] , \modmult_1/xin[531] ,
         \modmult_1/xin[530] , \modmult_1/xin[529] , \modmult_1/xin[528] ,
         \modmult_1/xin[527] , \modmult_1/xin[526] , \modmult_1/xin[525] ,
         \modmult_1/xin[524] , \modmult_1/xin[523] , \modmult_1/xin[522] ,
         \modmult_1/xin[521] , \modmult_1/xin[520] , \modmult_1/xin[519] ,
         \modmult_1/xin[518] , \modmult_1/xin[517] , \modmult_1/xin[516] ,
         \modmult_1/xin[515] , \modmult_1/xin[514] , \modmult_1/xin[513] ,
         \modmult_1/xin[512] , \modmult_1/xin[511] , \modmult_1/xin[510] ,
         \modmult_1/xin[509] , \modmult_1/xin[508] , \modmult_1/xin[507] ,
         \modmult_1/xin[506] , \modmult_1/xin[505] , \modmult_1/xin[504] ,
         \modmult_1/xin[503] , \modmult_1/xin[502] , \modmult_1/xin[501] ,
         \modmult_1/xin[500] , \modmult_1/xin[499] , \modmult_1/xin[498] ,
         \modmult_1/xin[497] , \modmult_1/xin[496] , \modmult_1/xin[495] ,
         \modmult_1/xin[494] , \modmult_1/xin[493] , \modmult_1/xin[492] ,
         \modmult_1/xin[491] , \modmult_1/xin[490] , \modmult_1/xin[489] ,
         \modmult_1/xin[488] , \modmult_1/xin[487] , \modmult_1/xin[486] ,
         \modmult_1/xin[485] , \modmult_1/xin[484] , \modmult_1/xin[483] ,
         \modmult_1/xin[482] , \modmult_1/xin[481] , \modmult_1/xin[480] ,
         \modmult_1/xin[479] , \modmult_1/xin[478] , \modmult_1/xin[477] ,
         \modmult_1/xin[476] , \modmult_1/xin[475] , \modmult_1/xin[474] ,
         \modmult_1/xin[473] , \modmult_1/xin[472] , \modmult_1/xin[471] ,
         \modmult_1/xin[470] , \modmult_1/xin[469] , \modmult_1/xin[468] ,
         \modmult_1/xin[467] , \modmult_1/xin[466] , \modmult_1/xin[465] ,
         \modmult_1/xin[464] , \modmult_1/xin[463] , \modmult_1/xin[462] ,
         \modmult_1/xin[461] , \modmult_1/xin[460] , \modmult_1/xin[459] ,
         \modmult_1/xin[458] , \modmult_1/xin[457] , \modmult_1/xin[456] ,
         \modmult_1/xin[455] , \modmult_1/xin[454] , \modmult_1/xin[453] ,
         \modmult_1/xin[452] , \modmult_1/xin[451] , \modmult_1/xin[450] ,
         \modmult_1/xin[449] , \modmult_1/xin[448] , \modmult_1/xin[447] ,
         \modmult_1/xin[446] , \modmult_1/xin[445] , \modmult_1/xin[444] ,
         \modmult_1/xin[443] , \modmult_1/xin[442] , \modmult_1/xin[441] ,
         \modmult_1/xin[440] , \modmult_1/xin[439] , \modmult_1/xin[438] ,
         \modmult_1/xin[437] , \modmult_1/xin[436] , \modmult_1/xin[435] ,
         \modmult_1/xin[434] , \modmult_1/xin[433] , \modmult_1/xin[432] ,
         \modmult_1/xin[431] , \modmult_1/xin[430] , \modmult_1/xin[429] ,
         \modmult_1/xin[428] , \modmult_1/xin[427] , \modmult_1/xin[426] ,
         \modmult_1/xin[425] , \modmult_1/xin[424] , \modmult_1/xin[423] ,
         \modmult_1/xin[422] , \modmult_1/xin[421] , \modmult_1/xin[420] ,
         \modmult_1/xin[419] , \modmult_1/xin[418] , \modmult_1/xin[417] ,
         \modmult_1/xin[416] , \modmult_1/xin[415] , \modmult_1/xin[414] ,
         \modmult_1/xin[413] , \modmult_1/xin[412] , \modmult_1/xin[411] ,
         \modmult_1/xin[410] , \modmult_1/xin[409] , \modmult_1/xin[408] ,
         \modmult_1/xin[407] , \modmult_1/xin[406] , \modmult_1/xin[405] ,
         \modmult_1/xin[404] , \modmult_1/xin[403] , \modmult_1/xin[402] ,
         \modmult_1/xin[401] , \modmult_1/xin[400] , \modmult_1/xin[399] ,
         \modmult_1/xin[398] , \modmult_1/xin[397] , \modmult_1/xin[396] ,
         \modmult_1/xin[395] , \modmult_1/xin[394] , \modmult_1/xin[393] ,
         \modmult_1/xin[392] , \modmult_1/xin[391] , \modmult_1/xin[390] ,
         \modmult_1/xin[389] , \modmult_1/xin[388] , \modmult_1/xin[387] ,
         \modmult_1/xin[386] , \modmult_1/xin[385] , \modmult_1/xin[384] ,
         \modmult_1/xin[383] , \modmult_1/xin[382] , \modmult_1/xin[381] ,
         \modmult_1/xin[380] , \modmult_1/xin[379] , \modmult_1/xin[378] ,
         \modmult_1/xin[377] , \modmult_1/xin[376] , \modmult_1/xin[375] ,
         \modmult_1/xin[374] , \modmult_1/xin[373] , \modmult_1/xin[372] ,
         \modmult_1/xin[371] , \modmult_1/xin[370] , \modmult_1/xin[369] ,
         \modmult_1/xin[368] , \modmult_1/xin[367] , \modmult_1/xin[366] ,
         \modmult_1/xin[365] , \modmult_1/xin[364] , \modmult_1/xin[363] ,
         \modmult_1/xin[362] , \modmult_1/xin[361] , \modmult_1/xin[360] ,
         \modmult_1/xin[359] , \modmult_1/xin[358] , \modmult_1/xin[357] ,
         \modmult_1/xin[356] , \modmult_1/xin[355] , \modmult_1/xin[354] ,
         \modmult_1/xin[353] , \modmult_1/xin[352] , \modmult_1/xin[351] ,
         \modmult_1/xin[350] , \modmult_1/xin[349] , \modmult_1/xin[348] ,
         \modmult_1/xin[347] , \modmult_1/xin[346] , \modmult_1/xin[345] ,
         \modmult_1/xin[344] , \modmult_1/xin[343] , \modmult_1/xin[342] ,
         \modmult_1/xin[341] , \modmult_1/xin[340] , \modmult_1/xin[339] ,
         \modmult_1/xin[338] , \modmult_1/xin[337] , \modmult_1/xin[336] ,
         \modmult_1/xin[335] , \modmult_1/xin[334] , \modmult_1/xin[333] ,
         \modmult_1/xin[332] , \modmult_1/xin[331] , \modmult_1/xin[330] ,
         \modmult_1/xin[329] , \modmult_1/xin[328] , \modmult_1/xin[327] ,
         \modmult_1/xin[326] , \modmult_1/xin[325] , \modmult_1/xin[324] ,
         \modmult_1/xin[323] , \modmult_1/xin[322] , \modmult_1/xin[321] ,
         \modmult_1/xin[320] , \modmult_1/xin[319] , \modmult_1/xin[318] ,
         \modmult_1/xin[317] , \modmult_1/xin[316] , \modmult_1/xin[315] ,
         \modmult_1/xin[314] , \modmult_1/xin[313] , \modmult_1/xin[312] ,
         \modmult_1/xin[311] , \modmult_1/xin[310] , \modmult_1/xin[309] ,
         \modmult_1/xin[308] , \modmult_1/xin[307] , \modmult_1/xin[306] ,
         \modmult_1/xin[305] , \modmult_1/xin[304] , \modmult_1/xin[303] ,
         \modmult_1/xin[302] , \modmult_1/xin[301] , \modmult_1/xin[300] ,
         \modmult_1/xin[299] , \modmult_1/xin[298] , \modmult_1/xin[297] ,
         \modmult_1/xin[296] , \modmult_1/xin[295] , \modmult_1/xin[294] ,
         \modmult_1/xin[293] , \modmult_1/xin[292] , \modmult_1/xin[291] ,
         \modmult_1/xin[290] , \modmult_1/xin[289] , \modmult_1/xin[288] ,
         \modmult_1/xin[287] , \modmult_1/xin[286] , \modmult_1/xin[285] ,
         \modmult_1/xin[284] , \modmult_1/xin[283] , \modmult_1/xin[282] ,
         \modmult_1/xin[281] , \modmult_1/xin[280] , \modmult_1/xin[279] ,
         \modmult_1/xin[278] , \modmult_1/xin[277] , \modmult_1/xin[276] ,
         \modmult_1/xin[275] , \modmult_1/xin[274] , \modmult_1/xin[273] ,
         \modmult_1/xin[272] , \modmult_1/xin[271] , \modmult_1/xin[270] ,
         \modmult_1/xin[269] , \modmult_1/xin[268] , \modmult_1/xin[267] ,
         \modmult_1/xin[266] , \modmult_1/xin[265] , \modmult_1/xin[264] ,
         \modmult_1/xin[263] , \modmult_1/xin[262] , \modmult_1/xin[261] ,
         \modmult_1/xin[260] , \modmult_1/xin[259] , \modmult_1/xin[258] ,
         \modmult_1/xin[257] , \modmult_1/xin[256] , \modmult_1/xin[255] ,
         \modmult_1/xin[254] , \modmult_1/xin[253] , \modmult_1/xin[252] ,
         \modmult_1/xin[251] , \modmult_1/xin[250] , \modmult_1/xin[249] ,
         \modmult_1/xin[248] , \modmult_1/xin[247] , \modmult_1/xin[246] ,
         \modmult_1/xin[245] , \modmult_1/xin[244] , \modmult_1/xin[243] ,
         \modmult_1/xin[242] , \modmult_1/xin[241] , \modmult_1/xin[240] ,
         \modmult_1/xin[239] , \modmult_1/xin[238] , \modmult_1/xin[237] ,
         \modmult_1/xin[236] , \modmult_1/xin[235] , \modmult_1/xin[234] ,
         \modmult_1/xin[233] , \modmult_1/xin[232] , \modmult_1/xin[231] ,
         \modmult_1/xin[230] , \modmult_1/xin[229] , \modmult_1/xin[228] ,
         \modmult_1/xin[227] , \modmult_1/xin[226] , \modmult_1/xin[225] ,
         \modmult_1/xin[224] , \modmult_1/xin[223] , \modmult_1/xin[222] ,
         \modmult_1/xin[221] , \modmult_1/xin[220] , \modmult_1/xin[219] ,
         \modmult_1/xin[218] , \modmult_1/xin[217] , \modmult_1/xin[216] ,
         \modmult_1/xin[215] , \modmult_1/xin[214] , \modmult_1/xin[213] ,
         \modmult_1/xin[212] , \modmult_1/xin[211] , \modmult_1/xin[210] ,
         \modmult_1/xin[209] , \modmult_1/xin[208] , \modmult_1/xin[207] ,
         \modmult_1/xin[206] , \modmult_1/xin[205] , \modmult_1/xin[204] ,
         \modmult_1/xin[203] , \modmult_1/xin[202] , \modmult_1/xin[201] ,
         \modmult_1/xin[200] , \modmult_1/xin[199] , \modmult_1/xin[198] ,
         \modmult_1/xin[197] , \modmult_1/xin[196] , \modmult_1/xin[195] ,
         \modmult_1/xin[194] , \modmult_1/xin[193] , \modmult_1/xin[192] ,
         \modmult_1/xin[191] , \modmult_1/xin[190] , \modmult_1/xin[189] ,
         \modmult_1/xin[188] , \modmult_1/xin[187] , \modmult_1/xin[186] ,
         \modmult_1/xin[185] , \modmult_1/xin[184] , \modmult_1/xin[183] ,
         \modmult_1/xin[182] , \modmult_1/xin[181] , \modmult_1/xin[180] ,
         \modmult_1/xin[179] , \modmult_1/xin[178] , \modmult_1/xin[177] ,
         \modmult_1/xin[176] , \modmult_1/xin[175] , \modmult_1/xin[174] ,
         \modmult_1/xin[173] , \modmult_1/xin[172] , \modmult_1/xin[171] ,
         \modmult_1/xin[170] , \modmult_1/xin[169] , \modmult_1/xin[168] ,
         \modmult_1/xin[167] , \modmult_1/xin[166] , \modmult_1/xin[165] ,
         \modmult_1/xin[164] , \modmult_1/xin[163] , \modmult_1/xin[162] ,
         \modmult_1/xin[161] , \modmult_1/xin[160] , \modmult_1/xin[159] ,
         \modmult_1/xin[158] , \modmult_1/xin[157] , \modmult_1/xin[156] ,
         \modmult_1/xin[155] , \modmult_1/xin[154] , \modmult_1/xin[153] ,
         \modmult_1/xin[152] , \modmult_1/xin[151] , \modmult_1/xin[150] ,
         \modmult_1/xin[149] , \modmult_1/xin[148] , \modmult_1/xin[147] ,
         \modmult_1/xin[146] , \modmult_1/xin[145] , \modmult_1/xin[144] ,
         \modmult_1/xin[143] , \modmult_1/xin[142] , \modmult_1/xin[141] ,
         \modmult_1/xin[140] , \modmult_1/xin[139] , \modmult_1/xin[138] ,
         \modmult_1/xin[137] , \modmult_1/xin[136] , \modmult_1/xin[135] ,
         \modmult_1/xin[134] , \modmult_1/xin[133] , \modmult_1/xin[132] ,
         \modmult_1/xin[131] , \modmult_1/xin[130] , \modmult_1/xin[129] ,
         \modmult_1/xin[128] , \modmult_1/xin[127] , \modmult_1/xin[126] ,
         \modmult_1/xin[125] , \modmult_1/xin[124] , \modmult_1/xin[123] ,
         \modmult_1/xin[122] , \modmult_1/xin[121] , \modmult_1/xin[120] ,
         \modmult_1/xin[119] , \modmult_1/xin[118] , \modmult_1/xin[117] ,
         \modmult_1/xin[116] , \modmult_1/xin[115] , \modmult_1/xin[114] ,
         \modmult_1/xin[113] , \modmult_1/xin[112] , \modmult_1/xin[111] ,
         \modmult_1/xin[110] , \modmult_1/xin[109] , \modmult_1/xin[108] ,
         \modmult_1/xin[107] , \modmult_1/xin[106] , \modmult_1/xin[105] ,
         \modmult_1/xin[104] , \modmult_1/xin[103] , \modmult_1/xin[102] ,
         \modmult_1/xin[101] , \modmult_1/xin[100] , \modmult_1/xin[99] ,
         \modmult_1/xin[98] , \modmult_1/xin[97] , \modmult_1/xin[96] ,
         \modmult_1/xin[95] , \modmult_1/xin[94] , \modmult_1/xin[93] ,
         \modmult_1/xin[92] , \modmult_1/xin[91] , \modmult_1/xin[90] ,
         \modmult_1/xin[89] , \modmult_1/xin[88] , \modmult_1/xin[87] ,
         \modmult_1/xin[86] , \modmult_1/xin[85] , \modmult_1/xin[84] ,
         \modmult_1/xin[83] , \modmult_1/xin[82] , \modmult_1/xin[81] ,
         \modmult_1/xin[80] , \modmult_1/xin[79] , \modmult_1/xin[78] ,
         \modmult_1/xin[77] , \modmult_1/xin[76] , \modmult_1/xin[75] ,
         \modmult_1/xin[74] , \modmult_1/xin[73] , \modmult_1/xin[72] ,
         \modmult_1/xin[71] , \modmult_1/xin[70] , \modmult_1/xin[69] ,
         \modmult_1/xin[68] , \modmult_1/xin[67] , \modmult_1/xin[66] ,
         \modmult_1/xin[65] , \modmult_1/xin[64] , \modmult_1/xin[63] ,
         \modmult_1/xin[62] , \modmult_1/xin[61] , \modmult_1/xin[60] ,
         \modmult_1/xin[59] , \modmult_1/xin[58] , \modmult_1/xin[57] ,
         \modmult_1/xin[56] , \modmult_1/xin[55] , \modmult_1/xin[54] ,
         \modmult_1/xin[53] , \modmult_1/xin[52] , \modmult_1/xin[51] ,
         \modmult_1/xin[50] , \modmult_1/xin[49] , \modmult_1/xin[48] ,
         \modmult_1/xin[47] , \modmult_1/xin[46] , \modmult_1/xin[45] ,
         \modmult_1/xin[44] , \modmult_1/xin[43] , \modmult_1/xin[42] ,
         \modmult_1/xin[41] , \modmult_1/xin[40] , \modmult_1/xin[39] ,
         \modmult_1/xin[38] , \modmult_1/xin[37] , \modmult_1/xin[36] ,
         \modmult_1/xin[35] , \modmult_1/xin[34] , \modmult_1/xin[33] ,
         \modmult_1/xin[32] , \modmult_1/xin[31] , \modmult_1/xin[30] ,
         \modmult_1/xin[29] , \modmult_1/xin[28] , \modmult_1/xin[27] ,
         \modmult_1/xin[26] , \modmult_1/xin[25] , \modmult_1/xin[24] ,
         \modmult_1/xin[23] , \modmult_1/xin[22] , \modmult_1/xin[21] ,
         \modmult_1/xin[20] , \modmult_1/xin[19] , \modmult_1/xin[18] ,
         \modmult_1/xin[17] , \modmult_1/xin[16] , \modmult_1/xin[15] ,
         \modmult_1/xin[14] , \modmult_1/xin[13] , \modmult_1/xin[12] ,
         \modmult_1/xin[11] , \modmult_1/xin[10] , \modmult_1/xin[9] ,
         \modmult_1/xin[8] , \modmult_1/xin[7] , \modmult_1/xin[6] ,
         \modmult_1/xin[5] , \modmult_1/xin[4] , \modmult_1/xin[3] ,
         \modmult_1/xin[2] , \modmult_1/xin[1] , \modmult_1/xin[0] ,
         \modmult_1/zin[0][1024] , \modmult_1/zin[0][1023] ,
         \modmult_1/zin[0][1022] , \modmult_1/zin[0][1021] ,
         \modmult_1/zin[0][1020] , \modmult_1/zin[0][1019] ,
         \modmult_1/zin[0][1018] , \modmult_1/zin[0][1017] ,
         \modmult_1/zin[0][1016] , \modmult_1/zin[0][1015] ,
         \modmult_1/zin[0][1014] , \modmult_1/zin[0][1013] ,
         \modmult_1/zin[0][1012] , \modmult_1/zin[0][1011] ,
         \modmult_1/zin[0][1010] , \modmult_1/zin[0][1009] ,
         \modmult_1/zin[0][1008] , \modmult_1/zin[0][1007] ,
         \modmult_1/zin[0][1006] , \modmult_1/zin[0][1005] ,
         \modmult_1/zin[0][1004] , \modmult_1/zin[0][1003] ,
         \modmult_1/zin[0][1002] , \modmult_1/zin[0][1001] ,
         \modmult_1/zin[0][1000] , \modmult_1/zin[0][999] ,
         \modmult_1/zin[0][998] , \modmult_1/zin[0][997] ,
         \modmult_1/zin[0][996] , \modmult_1/zin[0][995] ,
         \modmult_1/zin[0][994] , \modmult_1/zin[0][993] ,
         \modmult_1/zin[0][992] , \modmult_1/zin[0][991] ,
         \modmult_1/zin[0][990] , \modmult_1/zin[0][989] ,
         \modmult_1/zin[0][988] , \modmult_1/zin[0][987] ,
         \modmult_1/zin[0][986] , \modmult_1/zin[0][985] ,
         \modmult_1/zin[0][984] , \modmult_1/zin[0][983] ,
         \modmult_1/zin[0][982] , \modmult_1/zin[0][981] ,
         \modmult_1/zin[0][980] , \modmult_1/zin[0][979] ,
         \modmult_1/zin[0][978] , \modmult_1/zin[0][977] ,
         \modmult_1/zin[0][976] , \modmult_1/zin[0][975] ,
         \modmult_1/zin[0][974] , \modmult_1/zin[0][973] ,
         \modmult_1/zin[0][972] , \modmult_1/zin[0][971] ,
         \modmult_1/zin[0][970] , \modmult_1/zin[0][969] ,
         \modmult_1/zin[0][968] , \modmult_1/zin[0][967] ,
         \modmult_1/zin[0][966] , \modmult_1/zin[0][965] ,
         \modmult_1/zin[0][964] , \modmult_1/zin[0][963] ,
         \modmult_1/zin[0][962] , \modmult_1/zin[0][961] ,
         \modmult_1/zin[0][960] , \modmult_1/zin[0][959] ,
         \modmult_1/zin[0][958] , \modmult_1/zin[0][957] ,
         \modmult_1/zin[0][956] , \modmult_1/zin[0][955] ,
         \modmult_1/zin[0][954] , \modmult_1/zin[0][953] ,
         \modmult_1/zin[0][952] , \modmult_1/zin[0][951] ,
         \modmult_1/zin[0][950] , \modmult_1/zin[0][949] ,
         \modmult_1/zin[0][948] , \modmult_1/zin[0][947] ,
         \modmult_1/zin[0][946] , \modmult_1/zin[0][945] ,
         \modmult_1/zin[0][944] , \modmult_1/zin[0][943] ,
         \modmult_1/zin[0][942] , \modmult_1/zin[0][941] ,
         \modmult_1/zin[0][940] , \modmult_1/zin[0][939] ,
         \modmult_1/zin[0][938] , \modmult_1/zin[0][937] ,
         \modmult_1/zin[0][936] , \modmult_1/zin[0][935] ,
         \modmult_1/zin[0][934] , \modmult_1/zin[0][933] ,
         \modmult_1/zin[0][932] , \modmult_1/zin[0][931] ,
         \modmult_1/zin[0][930] , \modmult_1/zin[0][929] ,
         \modmult_1/zin[0][928] , \modmult_1/zin[0][927] ,
         \modmult_1/zin[0][926] , \modmult_1/zin[0][925] ,
         \modmult_1/zin[0][924] , \modmult_1/zin[0][923] ,
         \modmult_1/zin[0][922] , \modmult_1/zin[0][921] ,
         \modmult_1/zin[0][920] , \modmult_1/zin[0][919] ,
         \modmult_1/zin[0][918] , \modmult_1/zin[0][917] ,
         \modmult_1/zin[0][916] , \modmult_1/zin[0][915] ,
         \modmult_1/zin[0][914] , \modmult_1/zin[0][913] ,
         \modmult_1/zin[0][912] , \modmult_1/zin[0][911] ,
         \modmult_1/zin[0][910] , \modmult_1/zin[0][909] ,
         \modmult_1/zin[0][908] , \modmult_1/zin[0][907] ,
         \modmult_1/zin[0][906] , \modmult_1/zin[0][905] ,
         \modmult_1/zin[0][904] , \modmult_1/zin[0][903] ,
         \modmult_1/zin[0][902] , \modmult_1/zin[0][901] ,
         \modmult_1/zin[0][900] , \modmult_1/zin[0][899] ,
         \modmult_1/zin[0][898] , \modmult_1/zin[0][897] ,
         \modmult_1/zin[0][896] , \modmult_1/zin[0][895] ,
         \modmult_1/zin[0][894] , \modmult_1/zin[0][893] ,
         \modmult_1/zin[0][892] , \modmult_1/zin[0][891] ,
         \modmult_1/zin[0][890] , \modmult_1/zin[0][889] ,
         \modmult_1/zin[0][888] , \modmult_1/zin[0][887] ,
         \modmult_1/zin[0][886] , \modmult_1/zin[0][885] ,
         \modmult_1/zin[0][884] , \modmult_1/zin[0][883] ,
         \modmult_1/zin[0][882] , \modmult_1/zin[0][881] ,
         \modmult_1/zin[0][880] , \modmult_1/zin[0][879] ,
         \modmult_1/zin[0][878] , \modmult_1/zin[0][877] ,
         \modmult_1/zin[0][876] , \modmult_1/zin[0][875] ,
         \modmult_1/zin[0][874] , \modmult_1/zin[0][873] ,
         \modmult_1/zin[0][872] , \modmult_1/zin[0][871] ,
         \modmult_1/zin[0][870] , \modmult_1/zin[0][869] ,
         \modmult_1/zin[0][868] , \modmult_1/zin[0][867] ,
         \modmult_1/zin[0][866] , \modmult_1/zin[0][865] ,
         \modmult_1/zin[0][864] , \modmult_1/zin[0][863] ,
         \modmult_1/zin[0][862] , \modmult_1/zin[0][861] ,
         \modmult_1/zin[0][860] , \modmult_1/zin[0][859] ,
         \modmult_1/zin[0][858] , \modmult_1/zin[0][857] ,
         \modmult_1/zin[0][856] , \modmult_1/zin[0][855] ,
         \modmult_1/zin[0][854] , \modmult_1/zin[0][853] ,
         \modmult_1/zin[0][852] , \modmult_1/zin[0][851] ,
         \modmult_1/zin[0][850] , \modmult_1/zin[0][849] ,
         \modmult_1/zin[0][848] , \modmult_1/zin[0][847] ,
         \modmult_1/zin[0][846] , \modmult_1/zin[0][845] ,
         \modmult_1/zin[0][844] , \modmult_1/zin[0][843] ,
         \modmult_1/zin[0][842] , \modmult_1/zin[0][841] ,
         \modmult_1/zin[0][840] , \modmult_1/zin[0][839] ,
         \modmult_1/zin[0][838] , \modmult_1/zin[0][837] ,
         \modmult_1/zin[0][836] , \modmult_1/zin[0][835] ,
         \modmult_1/zin[0][834] , \modmult_1/zin[0][833] ,
         \modmult_1/zin[0][832] , \modmult_1/zin[0][831] ,
         \modmult_1/zin[0][830] , \modmult_1/zin[0][829] ,
         \modmult_1/zin[0][828] , \modmult_1/zin[0][827] ,
         \modmult_1/zin[0][826] , \modmult_1/zin[0][825] ,
         \modmult_1/zin[0][824] , \modmult_1/zin[0][823] ,
         \modmult_1/zin[0][822] , \modmult_1/zin[0][821] ,
         \modmult_1/zin[0][820] , \modmult_1/zin[0][819] ,
         \modmult_1/zin[0][818] , \modmult_1/zin[0][817] ,
         \modmult_1/zin[0][816] , \modmult_1/zin[0][815] ,
         \modmult_1/zin[0][814] , \modmult_1/zin[0][813] ,
         \modmult_1/zin[0][812] , \modmult_1/zin[0][811] ,
         \modmult_1/zin[0][810] , \modmult_1/zin[0][809] ,
         \modmult_1/zin[0][808] , \modmult_1/zin[0][807] ,
         \modmult_1/zin[0][806] , \modmult_1/zin[0][805] ,
         \modmult_1/zin[0][804] , \modmult_1/zin[0][803] ,
         \modmult_1/zin[0][802] , \modmult_1/zin[0][801] ,
         \modmult_1/zin[0][800] , \modmult_1/zin[0][799] ,
         \modmult_1/zin[0][798] , \modmult_1/zin[0][797] ,
         \modmult_1/zin[0][796] , \modmult_1/zin[0][795] ,
         \modmult_1/zin[0][794] , \modmult_1/zin[0][793] ,
         \modmult_1/zin[0][792] , \modmult_1/zin[0][791] ,
         \modmult_1/zin[0][790] , \modmult_1/zin[0][789] ,
         \modmult_1/zin[0][788] , \modmult_1/zin[0][787] ,
         \modmult_1/zin[0][786] , \modmult_1/zin[0][785] ,
         \modmult_1/zin[0][784] , \modmult_1/zin[0][783] ,
         \modmult_1/zin[0][782] , \modmult_1/zin[0][781] ,
         \modmult_1/zin[0][780] , \modmult_1/zin[0][779] ,
         \modmult_1/zin[0][778] , \modmult_1/zin[0][777] ,
         \modmult_1/zin[0][776] , \modmult_1/zin[0][775] ,
         \modmult_1/zin[0][774] , \modmult_1/zin[0][773] ,
         \modmult_1/zin[0][772] , \modmult_1/zin[0][771] ,
         \modmult_1/zin[0][770] , \modmult_1/zin[0][769] ,
         \modmult_1/zin[0][768] , \modmult_1/zin[0][767] ,
         \modmult_1/zin[0][766] , \modmult_1/zin[0][765] ,
         \modmult_1/zin[0][764] , \modmult_1/zin[0][763] ,
         \modmult_1/zin[0][762] , \modmult_1/zin[0][761] ,
         \modmult_1/zin[0][760] , \modmult_1/zin[0][759] ,
         \modmult_1/zin[0][758] , \modmult_1/zin[0][757] ,
         \modmult_1/zin[0][756] , \modmult_1/zin[0][755] ,
         \modmult_1/zin[0][754] , \modmult_1/zin[0][753] ,
         \modmult_1/zin[0][752] , \modmult_1/zin[0][751] ,
         \modmult_1/zin[0][750] , \modmult_1/zin[0][749] ,
         \modmult_1/zin[0][748] , \modmult_1/zin[0][747] ,
         \modmult_1/zin[0][746] , \modmult_1/zin[0][745] ,
         \modmult_1/zin[0][744] , \modmult_1/zin[0][743] ,
         \modmult_1/zin[0][742] , \modmult_1/zin[0][741] ,
         \modmult_1/zin[0][740] , \modmult_1/zin[0][739] ,
         \modmult_1/zin[0][738] , \modmult_1/zin[0][737] ,
         \modmult_1/zin[0][736] , \modmult_1/zin[0][735] ,
         \modmult_1/zin[0][734] , \modmult_1/zin[0][733] ,
         \modmult_1/zin[0][732] , \modmult_1/zin[0][731] ,
         \modmult_1/zin[0][730] , \modmult_1/zin[0][729] ,
         \modmult_1/zin[0][728] , \modmult_1/zin[0][727] ,
         \modmult_1/zin[0][726] , \modmult_1/zin[0][725] ,
         \modmult_1/zin[0][724] , \modmult_1/zin[0][723] ,
         \modmult_1/zin[0][722] , \modmult_1/zin[0][721] ,
         \modmult_1/zin[0][720] , \modmult_1/zin[0][719] ,
         \modmult_1/zin[0][718] , \modmult_1/zin[0][717] ,
         \modmult_1/zin[0][716] , \modmult_1/zin[0][715] ,
         \modmult_1/zin[0][714] , \modmult_1/zin[0][713] ,
         \modmult_1/zin[0][712] , \modmult_1/zin[0][711] ,
         \modmult_1/zin[0][710] , \modmult_1/zin[0][709] ,
         \modmult_1/zin[0][708] , \modmult_1/zin[0][707] ,
         \modmult_1/zin[0][706] , \modmult_1/zin[0][705] ,
         \modmult_1/zin[0][704] , \modmult_1/zin[0][703] ,
         \modmult_1/zin[0][702] , \modmult_1/zin[0][701] ,
         \modmult_1/zin[0][700] , \modmult_1/zin[0][699] ,
         \modmult_1/zin[0][698] , \modmult_1/zin[0][697] ,
         \modmult_1/zin[0][696] , \modmult_1/zin[0][695] ,
         \modmult_1/zin[0][694] , \modmult_1/zin[0][693] ,
         \modmult_1/zin[0][692] , \modmult_1/zin[0][691] ,
         \modmult_1/zin[0][690] , \modmult_1/zin[0][689] ,
         \modmult_1/zin[0][688] , \modmult_1/zin[0][687] ,
         \modmult_1/zin[0][686] , \modmult_1/zin[0][685] ,
         \modmult_1/zin[0][684] , \modmult_1/zin[0][683] ,
         \modmult_1/zin[0][682] , \modmult_1/zin[0][681] ,
         \modmult_1/zin[0][680] , \modmult_1/zin[0][679] ,
         \modmult_1/zin[0][678] , \modmult_1/zin[0][677] ,
         \modmult_1/zin[0][676] , \modmult_1/zin[0][675] ,
         \modmult_1/zin[0][674] , \modmult_1/zin[0][673] ,
         \modmult_1/zin[0][672] , \modmult_1/zin[0][671] ,
         \modmult_1/zin[0][670] , \modmult_1/zin[0][669] ,
         \modmult_1/zin[0][668] , \modmult_1/zin[0][667] ,
         \modmult_1/zin[0][666] , \modmult_1/zin[0][665] ,
         \modmult_1/zin[0][664] , \modmult_1/zin[0][663] ,
         \modmult_1/zin[0][662] , \modmult_1/zin[0][661] ,
         \modmult_1/zin[0][660] , \modmult_1/zin[0][659] ,
         \modmult_1/zin[0][658] , \modmult_1/zin[0][657] ,
         \modmult_1/zin[0][656] , \modmult_1/zin[0][655] ,
         \modmult_1/zin[0][654] , \modmult_1/zin[0][653] ,
         \modmult_1/zin[0][652] , \modmult_1/zin[0][651] ,
         \modmult_1/zin[0][650] , \modmult_1/zin[0][649] ,
         \modmult_1/zin[0][648] , \modmult_1/zin[0][647] ,
         \modmult_1/zin[0][646] , \modmult_1/zin[0][645] ,
         \modmult_1/zin[0][644] , \modmult_1/zin[0][643] ,
         \modmult_1/zin[0][642] , \modmult_1/zin[0][641] ,
         \modmult_1/zin[0][640] , \modmult_1/zin[0][639] ,
         \modmult_1/zin[0][638] , \modmult_1/zin[0][637] ,
         \modmult_1/zin[0][636] , \modmult_1/zin[0][635] ,
         \modmult_1/zin[0][634] , \modmult_1/zin[0][633] ,
         \modmult_1/zin[0][632] , \modmult_1/zin[0][631] ,
         \modmult_1/zin[0][630] , \modmult_1/zin[0][629] ,
         \modmult_1/zin[0][628] , \modmult_1/zin[0][627] ,
         \modmult_1/zin[0][626] , \modmult_1/zin[0][625] ,
         \modmult_1/zin[0][624] , \modmult_1/zin[0][623] ,
         \modmult_1/zin[0][622] , \modmult_1/zin[0][621] ,
         \modmult_1/zin[0][620] , \modmult_1/zin[0][619] ,
         \modmult_1/zin[0][618] , \modmult_1/zin[0][617] ,
         \modmult_1/zin[0][616] , \modmult_1/zin[0][615] ,
         \modmult_1/zin[0][614] , \modmult_1/zin[0][613] ,
         \modmult_1/zin[0][612] , \modmult_1/zin[0][611] ,
         \modmult_1/zin[0][610] , \modmult_1/zin[0][609] ,
         \modmult_1/zin[0][608] , \modmult_1/zin[0][607] ,
         \modmult_1/zin[0][606] , \modmult_1/zin[0][605] ,
         \modmult_1/zin[0][604] , \modmult_1/zin[0][603] ,
         \modmult_1/zin[0][602] , \modmult_1/zin[0][601] ,
         \modmult_1/zin[0][600] , \modmult_1/zin[0][599] ,
         \modmult_1/zin[0][598] , \modmult_1/zin[0][597] ,
         \modmult_1/zin[0][596] , \modmult_1/zin[0][595] ,
         \modmult_1/zin[0][594] , \modmult_1/zin[0][593] ,
         \modmult_1/zin[0][592] , \modmult_1/zin[0][591] ,
         \modmult_1/zin[0][590] , \modmult_1/zin[0][589] ,
         \modmult_1/zin[0][588] , \modmult_1/zin[0][587] ,
         \modmult_1/zin[0][586] , \modmult_1/zin[0][585] ,
         \modmult_1/zin[0][584] , \modmult_1/zin[0][583] ,
         \modmult_1/zin[0][582] , \modmult_1/zin[0][581] ,
         \modmult_1/zin[0][580] , \modmult_1/zin[0][579] ,
         \modmult_1/zin[0][578] , \modmult_1/zin[0][577] ,
         \modmult_1/zin[0][576] , \modmult_1/zin[0][575] ,
         \modmult_1/zin[0][574] , \modmult_1/zin[0][573] ,
         \modmult_1/zin[0][572] , \modmult_1/zin[0][571] ,
         \modmult_1/zin[0][570] , \modmult_1/zin[0][569] ,
         \modmult_1/zin[0][568] , \modmult_1/zin[0][567] ,
         \modmult_1/zin[0][566] , \modmult_1/zin[0][565] ,
         \modmult_1/zin[0][564] , \modmult_1/zin[0][563] ,
         \modmult_1/zin[0][562] , \modmult_1/zin[0][561] ,
         \modmult_1/zin[0][560] , \modmult_1/zin[0][559] ,
         \modmult_1/zin[0][558] , \modmult_1/zin[0][557] ,
         \modmult_1/zin[0][556] , \modmult_1/zin[0][555] ,
         \modmult_1/zin[0][554] , \modmult_1/zin[0][553] ,
         \modmult_1/zin[0][552] , \modmult_1/zin[0][551] ,
         \modmult_1/zin[0][550] , \modmult_1/zin[0][549] ,
         \modmult_1/zin[0][548] , \modmult_1/zin[0][547] ,
         \modmult_1/zin[0][546] , \modmult_1/zin[0][545] ,
         \modmult_1/zin[0][544] , \modmult_1/zin[0][543] ,
         \modmult_1/zin[0][542] , \modmult_1/zin[0][541] ,
         \modmult_1/zin[0][540] , \modmult_1/zin[0][539] ,
         \modmult_1/zin[0][538] , \modmult_1/zin[0][537] ,
         \modmult_1/zin[0][536] , \modmult_1/zin[0][535] ,
         \modmult_1/zin[0][534] , \modmult_1/zin[0][533] ,
         \modmult_1/zin[0][532] , \modmult_1/zin[0][531] ,
         \modmult_1/zin[0][530] , \modmult_1/zin[0][529] ,
         \modmult_1/zin[0][528] , \modmult_1/zin[0][527] ,
         \modmult_1/zin[0][526] , \modmult_1/zin[0][525] ,
         \modmult_1/zin[0][524] , \modmult_1/zin[0][523] ,
         \modmult_1/zin[0][522] , \modmult_1/zin[0][521] ,
         \modmult_1/zin[0][520] , \modmult_1/zin[0][519] ,
         \modmult_1/zin[0][518] , \modmult_1/zin[0][517] ,
         \modmult_1/zin[0][516] , \modmult_1/zin[0][515] ,
         \modmult_1/zin[0][514] , \modmult_1/zin[0][513] ,
         \modmult_1/zin[0][512] , \modmult_1/zin[0][511] ,
         \modmult_1/zin[0][510] , \modmult_1/zin[0][509] ,
         \modmult_1/zin[0][508] , \modmult_1/zin[0][507] ,
         \modmult_1/zin[0][506] , \modmult_1/zin[0][505] ,
         \modmult_1/zin[0][504] , \modmult_1/zin[0][503] ,
         \modmult_1/zin[0][502] , \modmult_1/zin[0][501] ,
         \modmult_1/zin[0][500] , \modmult_1/zin[0][499] ,
         \modmult_1/zin[0][498] , \modmult_1/zin[0][497] ,
         \modmult_1/zin[0][496] , \modmult_1/zin[0][495] ,
         \modmult_1/zin[0][494] , \modmult_1/zin[0][493] ,
         \modmult_1/zin[0][492] , \modmult_1/zin[0][491] ,
         \modmult_1/zin[0][490] , \modmult_1/zin[0][489] ,
         \modmult_1/zin[0][488] , \modmult_1/zin[0][487] ,
         \modmult_1/zin[0][486] , \modmult_1/zin[0][485] ,
         \modmult_1/zin[0][484] , \modmult_1/zin[0][483] ,
         \modmult_1/zin[0][482] , \modmult_1/zin[0][481] ,
         \modmult_1/zin[0][480] , \modmult_1/zin[0][479] ,
         \modmult_1/zin[0][478] , \modmult_1/zin[0][477] ,
         \modmult_1/zin[0][476] , \modmult_1/zin[0][475] ,
         \modmult_1/zin[0][474] , \modmult_1/zin[0][473] ,
         \modmult_1/zin[0][472] , \modmult_1/zin[0][471] ,
         \modmult_1/zin[0][470] , \modmult_1/zin[0][469] ,
         \modmult_1/zin[0][468] , \modmult_1/zin[0][467] ,
         \modmult_1/zin[0][466] , \modmult_1/zin[0][465] ,
         \modmult_1/zin[0][464] , \modmult_1/zin[0][463] ,
         \modmult_1/zin[0][462] , \modmult_1/zin[0][461] ,
         \modmult_1/zin[0][460] , \modmult_1/zin[0][459] ,
         \modmult_1/zin[0][458] , \modmult_1/zin[0][457] ,
         \modmult_1/zin[0][456] , \modmult_1/zin[0][455] ,
         \modmult_1/zin[0][454] , \modmult_1/zin[0][453] ,
         \modmult_1/zin[0][452] , \modmult_1/zin[0][451] ,
         \modmult_1/zin[0][450] , \modmult_1/zin[0][449] ,
         \modmult_1/zin[0][448] , \modmult_1/zin[0][447] ,
         \modmult_1/zin[0][446] , \modmult_1/zin[0][445] ,
         \modmult_1/zin[0][444] , \modmult_1/zin[0][443] ,
         \modmult_1/zin[0][442] , \modmult_1/zin[0][441] ,
         \modmult_1/zin[0][440] , \modmult_1/zin[0][439] ,
         \modmult_1/zin[0][438] , \modmult_1/zin[0][437] ,
         \modmult_1/zin[0][436] , \modmult_1/zin[0][435] ,
         \modmult_1/zin[0][434] , \modmult_1/zin[0][433] ,
         \modmult_1/zin[0][432] , \modmult_1/zin[0][431] ,
         \modmult_1/zin[0][430] , \modmult_1/zin[0][429] ,
         \modmult_1/zin[0][428] , \modmult_1/zin[0][427] ,
         \modmult_1/zin[0][426] , \modmult_1/zin[0][425] ,
         \modmult_1/zin[0][424] , \modmult_1/zin[0][423] ,
         \modmult_1/zin[0][422] , \modmult_1/zin[0][421] ,
         \modmult_1/zin[0][420] , \modmult_1/zin[0][419] ,
         \modmult_1/zin[0][418] , \modmult_1/zin[0][417] ,
         \modmult_1/zin[0][416] , \modmult_1/zin[0][415] ,
         \modmult_1/zin[0][414] , \modmult_1/zin[0][413] ,
         \modmult_1/zin[0][412] , \modmult_1/zin[0][411] ,
         \modmult_1/zin[0][410] , \modmult_1/zin[0][409] ,
         \modmult_1/zin[0][408] , \modmult_1/zin[0][407] ,
         \modmult_1/zin[0][406] , \modmult_1/zin[0][405] ,
         \modmult_1/zin[0][404] , \modmult_1/zin[0][403] ,
         \modmult_1/zin[0][402] , \modmult_1/zin[0][401] ,
         \modmult_1/zin[0][400] , \modmult_1/zin[0][399] ,
         \modmult_1/zin[0][398] , \modmult_1/zin[0][397] ,
         \modmult_1/zin[0][396] , \modmult_1/zin[0][395] ,
         \modmult_1/zin[0][394] , \modmult_1/zin[0][393] ,
         \modmult_1/zin[0][392] , \modmult_1/zin[0][391] ,
         \modmult_1/zin[0][390] , \modmult_1/zin[0][389] ,
         \modmult_1/zin[0][388] , \modmult_1/zin[0][387] ,
         \modmult_1/zin[0][386] , \modmult_1/zin[0][385] ,
         \modmult_1/zin[0][384] , \modmult_1/zin[0][383] ,
         \modmult_1/zin[0][382] , \modmult_1/zin[0][381] ,
         \modmult_1/zin[0][380] , \modmult_1/zin[0][379] ,
         \modmult_1/zin[0][378] , \modmult_1/zin[0][377] ,
         \modmult_1/zin[0][376] , \modmult_1/zin[0][375] ,
         \modmult_1/zin[0][374] , \modmult_1/zin[0][373] ,
         \modmult_1/zin[0][372] , \modmult_1/zin[0][371] ,
         \modmult_1/zin[0][370] , \modmult_1/zin[0][369] ,
         \modmult_1/zin[0][368] , \modmult_1/zin[0][367] ,
         \modmult_1/zin[0][366] , \modmult_1/zin[0][365] ,
         \modmult_1/zin[0][364] , \modmult_1/zin[0][363] ,
         \modmult_1/zin[0][362] , \modmult_1/zin[0][361] ,
         \modmult_1/zin[0][360] , \modmult_1/zin[0][359] ,
         \modmult_1/zin[0][358] , \modmult_1/zin[0][357] ,
         \modmult_1/zin[0][356] , \modmult_1/zin[0][355] ,
         \modmult_1/zin[0][354] , \modmult_1/zin[0][353] ,
         \modmult_1/zin[0][352] , \modmult_1/zin[0][351] ,
         \modmult_1/zin[0][350] , \modmult_1/zin[0][349] ,
         \modmult_1/zin[0][348] , \modmult_1/zin[0][347] ,
         \modmult_1/zin[0][346] , \modmult_1/zin[0][345] ,
         \modmult_1/zin[0][344] , \modmult_1/zin[0][343] ,
         \modmult_1/zin[0][342] , \modmult_1/zin[0][341] ,
         \modmult_1/zin[0][340] , \modmult_1/zin[0][339] ,
         \modmult_1/zin[0][338] , \modmult_1/zin[0][337] ,
         \modmult_1/zin[0][336] , \modmult_1/zin[0][335] ,
         \modmult_1/zin[0][334] , \modmult_1/zin[0][333] ,
         \modmult_1/zin[0][332] , \modmult_1/zin[0][331] ,
         \modmult_1/zin[0][330] , \modmult_1/zin[0][329] ,
         \modmult_1/zin[0][328] , \modmult_1/zin[0][327] ,
         \modmult_1/zin[0][326] , \modmult_1/zin[0][325] ,
         \modmult_1/zin[0][324] , \modmult_1/zin[0][323] ,
         \modmult_1/zin[0][322] , \modmult_1/zin[0][321] ,
         \modmult_1/zin[0][320] , \modmult_1/zin[0][319] ,
         \modmult_1/zin[0][318] , \modmult_1/zin[0][317] ,
         \modmult_1/zin[0][316] , \modmult_1/zin[0][315] ,
         \modmult_1/zin[0][314] , \modmult_1/zin[0][313] ,
         \modmult_1/zin[0][312] , \modmult_1/zin[0][311] ,
         \modmult_1/zin[0][310] , \modmult_1/zin[0][309] ,
         \modmult_1/zin[0][308] , \modmult_1/zin[0][307] ,
         \modmult_1/zin[0][306] , \modmult_1/zin[0][305] ,
         \modmult_1/zin[0][304] , \modmult_1/zin[0][303] ,
         \modmult_1/zin[0][302] , \modmult_1/zin[0][301] ,
         \modmult_1/zin[0][300] , \modmult_1/zin[0][299] ,
         \modmult_1/zin[0][298] , \modmult_1/zin[0][297] ,
         \modmult_1/zin[0][296] , \modmult_1/zin[0][295] ,
         \modmult_1/zin[0][294] , \modmult_1/zin[0][293] ,
         \modmult_1/zin[0][292] , \modmult_1/zin[0][291] ,
         \modmult_1/zin[0][290] , \modmult_1/zin[0][289] ,
         \modmult_1/zin[0][288] , \modmult_1/zin[0][287] ,
         \modmult_1/zin[0][286] , \modmult_1/zin[0][285] ,
         \modmult_1/zin[0][284] , \modmult_1/zin[0][283] ,
         \modmult_1/zin[0][282] , \modmult_1/zin[0][281] ,
         \modmult_1/zin[0][280] , \modmult_1/zin[0][279] ,
         \modmult_1/zin[0][278] , \modmult_1/zin[0][277] ,
         \modmult_1/zin[0][276] , \modmult_1/zin[0][275] ,
         \modmult_1/zin[0][274] , \modmult_1/zin[0][273] ,
         \modmult_1/zin[0][272] , \modmult_1/zin[0][271] ,
         \modmult_1/zin[0][270] , \modmult_1/zin[0][269] ,
         \modmult_1/zin[0][268] , \modmult_1/zin[0][267] ,
         \modmult_1/zin[0][266] , \modmult_1/zin[0][265] ,
         \modmult_1/zin[0][264] , \modmult_1/zin[0][263] ,
         \modmult_1/zin[0][262] , \modmult_1/zin[0][261] ,
         \modmult_1/zin[0][260] , \modmult_1/zin[0][259] ,
         \modmult_1/zin[0][258] , \modmult_1/zin[0][257] ,
         \modmult_1/zin[0][256] , \modmult_1/zin[0][255] ,
         \modmult_1/zin[0][254] , \modmult_1/zin[0][253] ,
         \modmult_1/zin[0][252] , \modmult_1/zin[0][251] ,
         \modmult_1/zin[0][250] , \modmult_1/zin[0][249] ,
         \modmult_1/zin[0][248] , \modmult_1/zin[0][247] ,
         \modmult_1/zin[0][246] , \modmult_1/zin[0][245] ,
         \modmult_1/zin[0][244] , \modmult_1/zin[0][243] ,
         \modmult_1/zin[0][242] , \modmult_1/zin[0][241] ,
         \modmult_1/zin[0][240] , \modmult_1/zin[0][239] ,
         \modmult_1/zin[0][238] , \modmult_1/zin[0][237] ,
         \modmult_1/zin[0][236] , \modmult_1/zin[0][235] ,
         \modmult_1/zin[0][234] , \modmult_1/zin[0][233] ,
         \modmult_1/zin[0][232] , \modmult_1/zin[0][231] ,
         \modmult_1/zin[0][230] , \modmult_1/zin[0][229] ,
         \modmult_1/zin[0][228] , \modmult_1/zin[0][227] ,
         \modmult_1/zin[0][226] , \modmult_1/zin[0][225] ,
         \modmult_1/zin[0][224] , \modmult_1/zin[0][223] ,
         \modmult_1/zin[0][222] , \modmult_1/zin[0][221] ,
         \modmult_1/zin[0][220] , \modmult_1/zin[0][219] ,
         \modmult_1/zin[0][218] , \modmult_1/zin[0][217] ,
         \modmult_1/zin[0][216] , \modmult_1/zin[0][215] ,
         \modmult_1/zin[0][214] , \modmult_1/zin[0][213] ,
         \modmult_1/zin[0][212] , \modmult_1/zin[0][211] ,
         \modmult_1/zin[0][210] , \modmult_1/zin[0][209] ,
         \modmult_1/zin[0][208] , \modmult_1/zin[0][207] ,
         \modmult_1/zin[0][206] , \modmult_1/zin[0][205] ,
         \modmult_1/zin[0][204] , \modmult_1/zin[0][203] ,
         \modmult_1/zin[0][202] , \modmult_1/zin[0][201] ,
         \modmult_1/zin[0][200] , \modmult_1/zin[0][199] ,
         \modmult_1/zin[0][198] , \modmult_1/zin[0][197] ,
         \modmult_1/zin[0][196] , \modmult_1/zin[0][195] ,
         \modmult_1/zin[0][194] , \modmult_1/zin[0][193] ,
         \modmult_1/zin[0][192] , \modmult_1/zin[0][191] ,
         \modmult_1/zin[0][190] , \modmult_1/zin[0][189] ,
         \modmult_1/zin[0][188] , \modmult_1/zin[0][187] ,
         \modmult_1/zin[0][186] , \modmult_1/zin[0][185] ,
         \modmult_1/zin[0][184] , \modmult_1/zin[0][183] ,
         \modmult_1/zin[0][182] , \modmult_1/zin[0][181] ,
         \modmult_1/zin[0][180] , \modmult_1/zin[0][179] ,
         \modmult_1/zin[0][178] , \modmult_1/zin[0][177] ,
         \modmult_1/zin[0][176] , \modmult_1/zin[0][175] ,
         \modmult_1/zin[0][174] , \modmult_1/zin[0][173] ,
         \modmult_1/zin[0][172] , \modmult_1/zin[0][171] ,
         \modmult_1/zin[0][170] , \modmult_1/zin[0][169] ,
         \modmult_1/zin[0][168] , \modmult_1/zin[0][167] ,
         \modmult_1/zin[0][166] , \modmult_1/zin[0][165] ,
         \modmult_1/zin[0][164] , \modmult_1/zin[0][163] ,
         \modmult_1/zin[0][162] , \modmult_1/zin[0][161] ,
         \modmult_1/zin[0][160] , \modmult_1/zin[0][159] ,
         \modmult_1/zin[0][158] , \modmult_1/zin[0][157] ,
         \modmult_1/zin[0][156] , \modmult_1/zin[0][155] ,
         \modmult_1/zin[0][154] , \modmult_1/zin[0][153] ,
         \modmult_1/zin[0][152] , \modmult_1/zin[0][151] ,
         \modmult_1/zin[0][150] , \modmult_1/zin[0][149] ,
         \modmult_1/zin[0][148] , \modmult_1/zin[0][147] ,
         \modmult_1/zin[0][146] , \modmult_1/zin[0][145] ,
         \modmult_1/zin[0][144] , \modmult_1/zin[0][143] ,
         \modmult_1/zin[0][142] , \modmult_1/zin[0][141] ,
         \modmult_1/zin[0][140] , \modmult_1/zin[0][139] ,
         \modmult_1/zin[0][138] , \modmult_1/zin[0][137] ,
         \modmult_1/zin[0][136] , \modmult_1/zin[0][135] ,
         \modmult_1/zin[0][134] , \modmult_1/zin[0][133] ,
         \modmult_1/zin[0][132] , \modmult_1/zin[0][131] ,
         \modmult_1/zin[0][130] , \modmult_1/zin[0][129] ,
         \modmult_1/zin[0][128] , \modmult_1/zin[0][127] ,
         \modmult_1/zin[0][126] , \modmult_1/zin[0][125] ,
         \modmult_1/zin[0][124] , \modmult_1/zin[0][123] ,
         \modmult_1/zin[0][122] , \modmult_1/zin[0][121] ,
         \modmult_1/zin[0][120] , \modmult_1/zin[0][119] ,
         \modmult_1/zin[0][118] , \modmult_1/zin[0][117] ,
         \modmult_1/zin[0][116] , \modmult_1/zin[0][115] ,
         \modmult_1/zin[0][114] , \modmult_1/zin[0][113] ,
         \modmult_1/zin[0][112] , \modmult_1/zin[0][111] ,
         \modmult_1/zin[0][110] , \modmult_1/zin[0][109] ,
         \modmult_1/zin[0][108] , \modmult_1/zin[0][107] ,
         \modmult_1/zin[0][106] , \modmult_1/zin[0][105] ,
         \modmult_1/zin[0][104] , \modmult_1/zin[0][103] ,
         \modmult_1/zin[0][102] , \modmult_1/zin[0][101] ,
         \modmult_1/zin[0][100] , \modmult_1/zin[0][99] ,
         \modmult_1/zin[0][98] , \modmult_1/zin[0][97] ,
         \modmult_1/zin[0][96] , \modmult_1/zin[0][95] ,
         \modmult_1/zin[0][94] , \modmult_1/zin[0][93] ,
         \modmult_1/zin[0][92] , \modmult_1/zin[0][91] ,
         \modmult_1/zin[0][90] , \modmult_1/zin[0][89] ,
         \modmult_1/zin[0][88] , \modmult_1/zin[0][87] ,
         \modmult_1/zin[0][86] , \modmult_1/zin[0][85] ,
         \modmult_1/zin[0][84] , \modmult_1/zin[0][83] ,
         \modmult_1/zin[0][82] , \modmult_1/zin[0][81] ,
         \modmult_1/zin[0][80] , \modmult_1/zin[0][79] ,
         \modmult_1/zin[0][78] , \modmult_1/zin[0][77] ,
         \modmult_1/zin[0][76] , \modmult_1/zin[0][75] ,
         \modmult_1/zin[0][74] , \modmult_1/zin[0][73] ,
         \modmult_1/zin[0][72] , \modmult_1/zin[0][71] ,
         \modmult_1/zin[0][70] , \modmult_1/zin[0][69] ,
         \modmult_1/zin[0][68] , \modmult_1/zin[0][67] ,
         \modmult_1/zin[0][66] , \modmult_1/zin[0][65] ,
         \modmult_1/zin[0][64] , \modmult_1/zin[0][63] ,
         \modmult_1/zin[0][62] , \modmult_1/zin[0][61] ,
         \modmult_1/zin[0][60] , \modmult_1/zin[0][59] ,
         \modmult_1/zin[0][58] , \modmult_1/zin[0][57] ,
         \modmult_1/zin[0][56] , \modmult_1/zin[0][55] ,
         \modmult_1/zin[0][54] , \modmult_1/zin[0][53] ,
         \modmult_1/zin[0][52] , \modmult_1/zin[0][51] ,
         \modmult_1/zin[0][50] , \modmult_1/zin[0][49] ,
         \modmult_1/zin[0][48] , \modmult_1/zin[0][47] ,
         \modmult_1/zin[0][46] , \modmult_1/zin[0][45] ,
         \modmult_1/zin[0][44] , \modmult_1/zin[0][43] ,
         \modmult_1/zin[0][42] , \modmult_1/zin[0][41] ,
         \modmult_1/zin[0][40] , \modmult_1/zin[0][39] ,
         \modmult_1/zin[0][38] , \modmult_1/zin[0][37] ,
         \modmult_1/zin[0][36] , \modmult_1/zin[0][35] ,
         \modmult_1/zin[0][34] , \modmult_1/zin[0][33] ,
         \modmult_1/zin[0][32] , \modmult_1/zin[0][31] ,
         \modmult_1/zin[0][30] , \modmult_1/zin[0][29] ,
         \modmult_1/zin[0][28] , \modmult_1/zin[0][27] ,
         \modmult_1/zin[0][26] , \modmult_1/zin[0][25] ,
         \modmult_1/zin[0][24] , \modmult_1/zin[0][23] ,
         \modmult_1/zin[0][22] , \modmult_1/zin[0][21] ,
         \modmult_1/zin[0][20] , \modmult_1/zin[0][19] ,
         \modmult_1/zin[0][18] , \modmult_1/zin[0][17] ,
         \modmult_1/zin[0][16] , \modmult_1/zin[0][15] ,
         \modmult_1/zin[0][14] , \modmult_1/zin[0][13] ,
         \modmult_1/zin[0][12] , \modmult_1/zin[0][11] ,
         \modmult_1/zin[0][10] , \modmult_1/zin[0][9] , \modmult_1/zin[0][8] ,
         \modmult_1/zin[0][7] , \modmult_1/zin[0][6] , \modmult_1/zin[0][5] ,
         \modmult_1/zin[0][4] , \modmult_1/zin[0][3] , \modmult_1/zin[0][2] ,
         \modmult_1/zin[0][1] , \modmult_1/zin[0][0] ,
         \modmult_1/zout[0][1024] , n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
         n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
         n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
         n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
         n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
         n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
         n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
         n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511,
         n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
         n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
         n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
         n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
         n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
         n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
         n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575,
         n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
         n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
         n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
         n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
         n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711,
         n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719,
         n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727,
         n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735,
         n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
         n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751,
         n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
         n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
         n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775,
         n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
         n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791,
         n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799,
         n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807,
         n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
         n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823,
         n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
         n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839,
         n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847,
         n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855,
         n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863,
         n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871,
         n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879,
         n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887,
         n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895,
         n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
         n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911,
         n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919,
         n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927,
         n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935,
         n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943,
         n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951,
         n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959,
         n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967,
         n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975,
         n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983,
         n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991,
         n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999,
         n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007,
         n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015,
         n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023,
         n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
         n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039,
         n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047,
         n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055,
         n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063,
         n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071,
         n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079,
         n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087,
         n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095,
         n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103,
         n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111,
         n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
         n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127,
         n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135,
         n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143,
         n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151,
         n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159,
         n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167,
         n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175,
         n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183,
         n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191,
         n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199,
         n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207,
         n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215,
         n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223,
         n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231,
         n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239,
         n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247,
         n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255,
         n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263,
         n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271,
         n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279,
         n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287,
         n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295,
         n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303,
         n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311,
         n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319,
         n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327,
         n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335,
         n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343,
         n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351,
         n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359,
         n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367,
         n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375,
         n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383,
         n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391,
         n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399,
         n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407,
         n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415,
         n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423,
         n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431,
         n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439,
         n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
         n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455,
         n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
         n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471,
         n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
         n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487,
         n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495,
         n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503,
         n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511,
         n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519,
         n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527,
         n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
         n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543,
         n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
         n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559,
         n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567,
         n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575,
         n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583,
         n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591,
         n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599,
         n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
         n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615,
         n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
         n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631,
         n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639,
         n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647,
         n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655,
         n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663,
         n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671,
         n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
         n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687,
         n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
         n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703,
         n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711,
         n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
         n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727,
         n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735,
         n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743,
         n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751,
         n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759,
         n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767,
         n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775,
         n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783,
         n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791,
         n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799,
         n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807,
         n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815,
         n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823,
         n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831,
         n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839,
         n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847,
         n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855,
         n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863,
         n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871,
         n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879,
         n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887,
         n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895,
         n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903,
         n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911,
         n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919,
         n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927,
         n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935,
         n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943,
         n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951,
         n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959,
         n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967,
         n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975,
         n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983,
         n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991,
         n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999,
         n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007,
         n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015,
         n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023,
         n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031,
         n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039,
         n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047,
         n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055,
         n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063,
         n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071,
         n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079,
         n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087,
         n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095,
         n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103,
         n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111,
         n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119,
         n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127,
         n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135,
         n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143,
         n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151,
         n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159,
         n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167,
         n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175,
         n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183,
         n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191,
         n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199,
         n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207,
         n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215,
         n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223,
         n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231,
         n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239,
         n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247,
         n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255,
         n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263,
         n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271,
         n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279,
         n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287,
         n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295,
         n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303,
         n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311,
         n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319,
         n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327,
         n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335,
         n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343,
         n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351,
         n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359,
         n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367,
         n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375,
         n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383,
         n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391,
         n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399,
         n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407,
         n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415,
         n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423,
         n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431,
         n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439,
         n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447,
         n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455,
         n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463,
         n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471,
         n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479,
         n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487,
         n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495,
         n16496, n16497, n16498, n16499, n16500, n16501, n16502, n16503,
         n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511,
         n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519,
         n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527,
         n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535,
         n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543,
         n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551,
         n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559,
         n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567,
         n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575,
         n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583,
         n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591,
         n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599,
         n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607,
         n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615,
         n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623,
         n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631,
         n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639,
         n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647,
         n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655,
         n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663,
         n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671,
         n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679,
         n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687,
         n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695,
         n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703,
         n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711,
         n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719,
         n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727,
         n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735,
         n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743,
         n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751,
         n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759,
         n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767,
         n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775,
         n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783,
         n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791,
         n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799,
         n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807,
         n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815,
         n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823,
         n16824, n16825, n16826, n16827, n16828, n16829, n16830, n16831,
         n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839,
         n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847,
         n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16855,
         n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863,
         n16864, n16865, n16866, n16867, n16868, n16869, n16870, n16871,
         n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879,
         n16880, n16881, n16882, n16883, n16884, n16885, n16886, n16887,
         n16888, n16889, n16890, n16891, n16892, n16893, n16894, n16895,
         n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903,
         n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911,
         n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919,
         n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927,
         n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935,
         n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943,
         n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951,
         n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959,
         n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967,
         n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975,
         n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983,
         n16984, n16985, n16986, n16987, n16988, n16989, n16990, n16991,
         n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999,
         n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007,
         n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015,
         n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023,
         n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031,
         n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039,
         n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047,
         n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055,
         n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063,
         n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071,
         n17072, n17073, n17074, n17075, n17076, n17077, n17078, n17079,
         n17080, n17081, n17082, n17083, n17084, n17085, n17086, n17087,
         n17088, n17089, n17090, n17091, n17092, n17093, n17094, n17095,
         n17096, n17097, n17098, n17099, n17100, n17101, n17102, n17103,
         n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111,
         n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119,
         n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127,
         n17128, n17129, n17130, n17131, n17132, n17133, n17134, n17135,
         n17136, n17137, n17138, n17139, n17140, n17141, n17142, n17143,
         n17144, n17145, n17146, n17147, n17148, n17149, n17150, n17151,
         n17152, n17153, n17154, n17155, n17156, n17157, n17158, n17159,
         n17160, n17161, n17162, n17163, n17164, n17165, n17166, n17167,
         n17168, n17169, n17170, n17171, n17172, n17173, n17174, n17175,
         n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183,
         n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191,
         n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199,
         n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207,
         n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215,
         n17216, n17217, n17218, n17219, n17220, n17221, n17222, n17223,
         n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231,
         n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239,
         n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247,
         n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255,
         n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17263,
         n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271,
         n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279,
         n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287,
         n17288, n17289, n17290, n17291, n17292, n17293, n17294, n17295,
         n17296, n17297, n17298, n17299, n17300, n17301, n17302, n17303,
         n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311,
         n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319,
         n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327,
         n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17335,
         n17336, n17337, n17338, n17339, n17340, n17341, n17342, n17343,
         n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351,
         n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359,
         n17360, n17361, n17362, n17363, n17364, n17365, n17366, n17367,
         n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375,
         n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383,
         n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391,
         n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399,
         n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407,
         n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415,
         n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423,
         n17424, n17425, n17426, n17427, n17428, n17429, n17430, n17431,
         n17432, n17433, n17434, n17435, n17436, n17437, n17438, n17439,
         n17440, n17441, n17442, n17443, n17444, n17445, n17446, n17447,
         n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455,
         n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463,
         n17464, n17465, n17466, n17467, n17468, n17469, n17470, n17471,
         n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479,
         n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487,
         n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495,
         n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503,
         n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511,
         n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519,
         n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527,
         n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535,
         n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543,
         n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17551,
         n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559,
         n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567,
         n17568, n17569, n17570, n17571, n17572, n17573, n17574, n17575,
         n17576, n17577, n17578, n17579, n17580, n17581, n17582, n17583,
         n17584, n17585, n17586, n17587, n17588, n17589, n17590, n17591,
         n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599,
         n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607,
         n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615,
         n17616, n17617, n17618, n17619, n17620, n17621, n17622, n17623,
         n17624, n17625, n17626, n17627, n17628, n17629, n17630, n17631,
         n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17639,
         n17640, n17641, n17642, n17643, n17644, n17645, n17646, n17647,
         n17648, n17649, n17650, n17651, n17652, n17653, n17654, n17655,
         n17656, n17657, n17658, n17659, n17660, n17661, n17662, n17663,
         n17664, n17665, n17666, n17667, n17668, n17669, n17670, n17671,
         n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679,
         n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687,
         n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695,
         n17696, n17697, n17698, n17699, n17700, n17701, n17702, n17703,
         n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711,
         n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719,
         n17720, n17721, n17722, n17723, n17724, n17725, n17726, n17727,
         n17728, n17729, n17730, n17731, n17732, n17733, n17734, n17735,
         n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743,
         n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751,
         n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759,
         n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767,
         n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775,
         n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783,
         n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791,
         n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799,
         n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807,
         n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815,
         n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823,
         n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831,
         n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839,
         n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847,
         n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855,
         n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863,
         n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871,
         n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879,
         n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887,
         n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895,
         n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903,
         n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17911,
         n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919,
         n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17927,
         n17928, n17929, n17930, n17931, n17932, n17933, n17934, n17935,
         n17936, n17937, n17938, n17939, n17940, n17941, n17942, n17943,
         n17944, n17945, n17946, n17947, n17948, n17949, n17950, n17951,
         n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959,
         n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967,
         n17968, n17969, n17970, n17971, n17972, n17973, n17974, n17975,
         n17976, n17977, n17978, n17979, n17980, n17981, n17982, n17983,
         n17984, n17985, n17986, n17987, n17988, n17989, n17990, n17991,
         n17992, n17993, n17994, n17995, n17996, n17997, n17998, n17999,
         n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007,
         n18008, n18009, n18010, n18011, n18012, n18013, n18014, n18015,
         n18016, n18017, n18018, n18019, n18020, n18021, n18022, n18023,
         n18024, n18025, n18026, n18027, n18028, n18029, n18030, n18031,
         n18032, n18033, n18034, n18035, n18036, n18037, n18038, n18039,
         n18040, n18041, n18042, n18043, n18044, n18045, n18046, n18047,
         n18048, n18049, n18050, n18051, n18052, n18053, n18054, n18055,
         n18056, n18057, n18058, n18059, n18060, n18061, n18062, n18063,
         n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071,
         n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18079,
         n18080, n18081, n18082, n18083, n18084, n18085, n18086, n18087,
         n18088, n18089, n18090, n18091, n18092, n18093, n18094, n18095,
         n18096, n18097, n18098, n18099, n18100, n18101, n18102, n18103,
         n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111,
         n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119,
         n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127,
         n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135,
         n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143,
         n18144, n18145, n18146, n18147, n18148, n18149, n18150, n18151,
         n18152, n18153, n18154, n18155, n18156, n18157, n18158, n18159,
         n18160, n18161, n18162, n18163, n18164, n18165, n18166, n18167,
         n18168, n18169, n18170, n18171, n18172, n18173, n18174, n18175,
         n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183,
         n18184, n18185, n18186, n18187, n18188, n18189, n18190, n18191,
         n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199,
         n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207,
         n18208, n18209, n18210, n18211, n18212, n18213, n18214, n18215,
         n18216, n18217, n18218, n18219, n18220, n18221, n18222, n18223,
         n18224, n18225, n18226, n18227, n18228, n18229, n18230, n18231,
         n18232, n18233, n18234, n18235, n18236, n18237, n18238, n18239,
         n18240, n18241, n18242, n18243, n18244, n18245, n18246, n18247,
         n18248, n18249, n18250, n18251, n18252, n18253, n18254, n18255,
         n18256, n18257, n18258, n18259, n18260, n18261, n18262, n18263,
         n18264, n18265, n18266, n18267, n18268, n18269, n18270, n18271,
         n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279,
         n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287,
         n18288, n18289, n18290, n18291, n18292, n18293, n18294, n18295,
         n18296, n18297, n18298, n18299, n18300, n18301, n18302, n18303,
         n18304, n18305, n18306, n18307, n18308, n18309, n18310, n18311,
         n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319,
         n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327,
         n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335,
         n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343,
         n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351,
         n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359,
         n18360, n18361, n18362, n18363, n18364, n18365, n18366, n18367,
         n18368, n18369, n18370, n18371, n18372, n18373, n18374, n18375,
         n18376, n18377, n18378, n18379, n18380, n18381, n18382, n18383,
         n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391,
         n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399,
         n18400, n18401, n18402, n18403, n18404, n18405, n18406, n18407,
         n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415,
         n18416, n18417, n18418, n18419, n18420, n18421, n18422, n18423,
         n18424, n18425, n18426, n18427, n18428, n18429, n18430, n18431,
         n18432, n18433, n18434, n18435, n18436, n18437, n18438, n18439,
         n18440, n18441, n18442, n18443, n18444, n18445, n18446, n18447,
         n18448, n18449, n18450, n18451, n18452, n18453, n18454, n18455,
         n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463,
         n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471,
         n18472, n18473, n18474, n18475, n18476, n18477, n18478, n18479,
         n18480, n18481, n18482, n18483, n18484, n18485, n18486, n18487,
         n18488, n18489, n18490, n18491, n18492, n18493, n18494, n18495,
         n18496, n18497, n18498, n18499, n18500, n18501, n18502, n18503,
         n18504, n18505, n18506, n18507, n18508, n18509, n18510, n18511,
         n18512, n18513, n18514, n18515, n18516, n18517, n18518, n18519,
         n18520, n18521, n18522, n18523, n18524, n18525, n18526, n18527,
         n18528, n18529, n18530, n18531, n18532, n18533, n18534, n18535,
         n18536, n18537, n18538, n18539, n18540, n18541, n18542, n18543,
         n18544, n18545, n18546, n18547, n18548, n18549, n18550, n18551,
         n18552, n18553, n18554, n18555, n18556, n18557, n18558, n18559,
         n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567,
         n18568, n18569, n18570, n18571, n18572, n18573, n18574, n18575,
         n18576, n18577, n18578, n18579, n18580, n18581, n18582, n18583,
         n18584, n18585, n18586, n18587, n18588, n18589, n18590, n18591,
         n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599,
         n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607,
         n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615,
         n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623,
         n18624, n18625, n18626, n18627, n18628, n18629, n18630, n18631,
         n18632, n18633, n18634, n18635, n18636, n18637, n18638, n18639,
         n18640, n18641, n18642, n18643, n18644, n18645, n18646, n18647,
         n18648, n18649, n18650, n18651, n18652, n18653, n18654, n18655,
         n18656, n18657, n18658, n18659, n18660, n18661, n18662, n18663,
         n18664, n18665, n18666, n18667, n18668, n18669, n18670, n18671,
         n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18679,
         n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687,
         n18688, n18689, n18690, n18691, n18692, n18693, n18694, n18695,
         n18696, n18697, n18698, n18699, n18700, n18701, n18702, n18703,
         n18704, n18705, n18706, n18707, n18708, n18709, n18710, n18711,
         n18712, n18713, n18714, n18715, n18716, n18717, n18718, n18719,
         n18720, n18721, n18722, n18723, n18724, n18725, n18726, n18727,
         n18728, n18729, n18730, n18731, n18732, n18733, n18734, n18735,
         n18736, n18737, n18738, n18739, n18740, n18741, n18742, n18743,
         n18744, n18745, n18746, n18747, n18748, n18749, n18750, n18751,
         n18752, n18753, n18754, n18755, n18756, n18757, n18758, n18759,
         n18760, n18761, n18762, n18763, n18764, n18765, n18766, n18767,
         n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18775,
         n18776, n18777, n18778, n18779, n18780, n18781, n18782, n18783,
         n18784, n18785, n18786, n18787, n18788, n18789, n18790, n18791,
         n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18799,
         n18800, n18801, n18802, n18803, n18804, n18805, n18806, n18807,
         n18808, n18809, n18810, n18811, n18812, n18813, n18814, n18815,
         n18816, n18817, n18818, n18819, n18820, n18821, n18822, n18823,
         n18824, n18825, n18826, n18827, n18828, n18829, n18830, n18831,
         n18832, n18833, n18834, n18835, n18836, n18837, n18838, n18839,
         n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847,
         n18848, n18849, n18850, n18851, n18852, n18853, n18854, n18855,
         n18856, n18857, n18858, n18859, n18860, n18861, n18862, n18863,
         n18864, n18865, n18866, n18867, n18868, n18869, n18870, n18871,
         n18872, n18873, n18874, n18875, n18876, n18877, n18878, n18879,
         n18880, n18881, n18882, n18883, n18884, n18885, n18886, n18887,
         n18888, n18889, n18890, n18891, n18892, n18893, n18894, n18895,
         n18896, n18897, n18898, n18899, n18900, n18901, n18902, n18903,
         n18904, n18905, n18906, n18907, n18908, n18909, n18910, n18911,
         n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18919,
         n18920, n18921, n18922, n18923, n18924, n18925, n18926, n18927,
         n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935,
         n18936, n18937, n18938, n18939, n18940, n18941, n18942, n18943,
         n18944, n18945, n18946, n18947, n18948, n18949, n18950, n18951,
         n18952, n18953, n18954, n18955, n18956, n18957, n18958, n18959,
         n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967,
         n18968, n18969, n18970, n18971, n18972, n18973, n18974, n18975,
         n18976, n18977, n18978, n18979, n18980, n18981, n18982, n18983,
         n18984, n18985, n18986, n18987, n18988, n18989, n18990, n18991,
         n18992, n18993, n18994, n18995, n18996, n18997, n18998, n18999,
         n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19007,
         n19008, n19009, n19010, n19011, n19012, n19013, n19014, n19015,
         n19016, n19017, n19018, n19019, n19020, n19021, n19022, n19023,
         n19024, n19025, n19026, n19027, n19028, n19029, n19030, n19031,
         n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039,
         n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047,
         n19048, n19049, n19050, n19051, n19052, n19053, n19054, n19055,
         n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19063,
         n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071,
         n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079,
         n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087,
         n19088, n19089, n19090, n19091, n19092, n19093, n19094, n19095,
         n19096, n19097, n19098, n19099, n19100, n19101, n19102, n19103,
         n19104, n19105, n19106, n19107, n19108, n19109, n19110, n19111,
         n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119,
         n19120, n19121, n19122, n19123, n19124, n19125, n19126, n19127,
         n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135,
         n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143,
         n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151,
         n19152, n19153, n19154, n19155, n19156, n19157, n19158, n19159,
         n19160, n19161, n19162, n19163, n19164, n19165, n19166, n19167,
         n19168, n19169, n19170, n19171, n19172, n19173, n19174, n19175,
         n19176, n19177, n19178, n19179, n19180, n19181, n19182, n19183,
         n19184, n19185, n19186, n19187, n19188, n19189, n19190, n19191,
         n19192, n19193, n19194, n19195, n19196, n19197, n19198, n19199,
         n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19207,
         n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215,
         n19216, n19217, n19218, n19219, n19220, n19221, n19222, n19223,
         n19224, n19225, n19226, n19227, n19228, n19229, n19230, n19231,
         n19232, n19233, n19234, n19235, n19236, n19237, n19238, n19239,
         n19240, n19241, n19242, n19243, n19244, n19245, n19246, n19247,
         n19248, n19249, n19250, n19251, n19252, n19253, n19254, n19255,
         n19256, n19257, n19258, n19259, n19260, n19261, n19262, n19263,
         n19264, n19265, n19266, n19267, n19268, n19269, n19270, n19271,
         n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279,
         n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287,
         n19288, n19289, n19290, n19291, n19292, n19293, n19294, n19295,
         n19296, n19297, n19298, n19299, n19300, n19301, n19302, n19303,
         n19304, n19305, n19306, n19307, n19308, n19309, n19310, n19311,
         n19312, n19313, n19314, n19315, n19316, n19317, n19318, n19319,
         n19320, n19321, n19322, n19323, n19324, n19325, n19326, n19327,
         n19328, n19329, n19330, n19331, n19332, n19333, n19334, n19335,
         n19336, n19337, n19338, n19339, n19340, n19341, n19342, n19343,
         n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351,
         n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359,
         n19360, n19361, n19362, n19363, n19364, n19365, n19366, n19367,
         n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19375,
         n19376, n19377, n19378, n19379, n19380, n19381, n19382, n19383,
         n19384, n19385, n19386, n19387, n19388, n19389, n19390, n19391,
         n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399,
         n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407,
         n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415,
         n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423,
         n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19431,
         n19432, n19433, n19434, n19435, n19436, n19437, n19438, n19439,
         n19440, n19441, n19442, n19443, n19444, n19445, n19446, n19447,
         n19448, n19449, n19450, n19451, n19452, n19453, n19454, n19455,
         n19456, n19457, n19458, n19459, n19460, n19461, n19462, n19463,
         n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471,
         n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479,
         n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487,
         n19488, n19489, n19490, n19491, n19492, n19493, n19494, n19495,
         n19496, n19497, n19498, n19499, n19500, n19501, n19502, n19503,
         n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511,
         n19512, n19513, n19514, n19515, n19516, n19517, n19518, n19519,
         n19520, n19521, n19522, n19523, n19524, n19525, n19526, n19527,
         n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535,
         n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543,
         n19544, n19545, n19546, n19547, n19548, n19549, n19550, n19551,
         n19552, n19553, n19554, n19555, n19556, n19557, n19558, n19559,
         n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567,
         n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575,
         n19576, n19577, n19578, n19579, n19580, n19581, n19582, n19583,
         n19584, n19585, n19586, n19587, n19588, n19589, n19590, n19591,
         n19592, n19593, n19594, n19595, n19596, n19597, n19598, n19599,
         n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607,
         n19608, n19609, n19610, n19611, n19612, n19613, n19614, n19615,
         n19616, n19617, n19618, n19619, n19620, n19621, n19622, n19623,
         n19624, n19625, n19626, n19627, n19628, n19629, n19630, n19631,
         n19632, n19633, n19634, n19635, n19636, n19637, n19638, n19639,
         n19640, n19641, n19642, n19643, n19644, n19645, n19646, n19647,
         n19648, n19649, n19650, n19651, n19652, n19653, n19654, n19655,
         n19656, n19657, n19658, n19659, n19660, n19661, n19662, n19663,
         n19664, n19665, n19666, n19667, n19668, n19669, n19670, n19671,
         n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679,
         n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687,
         n19688, n19689, n19690, n19691, n19692, n19693, n19694, n19695,
         n19696, n19697, n19698, n19699, n19700, n19701, n19702, n19703,
         n19704, n19705, n19706, n19707, n19708, n19709, n19710, n19711,
         n19712, n19713, n19714, n19715, n19716, n19717, n19718, n19719,
         n19720, n19721, n19722, n19723, n19724, n19725, n19726, n19727,
         n19728, n19729, n19730, n19731, n19732, n19733, n19734, n19735,
         n19736, n19737, n19738, n19739, n19740, n19741, n19742, n19743,
         n19744, n19745, n19746, n19747, n19748, n19749, n19750, n19751,
         n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759,
         n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19767,
         n19768, n19769, n19770, n19771, n19772, n19773, n19774, n19775,
         n19776, n19777, n19778, n19779, n19780, n19781, n19782, n19783,
         n19784, n19785, n19786, n19787, n19788, n19789, n19790, n19791,
         n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19799,
         n19800, n19801, n19802, n19803, n19804, n19805, n19806, n19807,
         n19808, n19809, n19810, n19811, n19812, n19813, n19814, n19815,
         n19816, n19817, n19818, n19819, n19820, n19821, n19822, n19823,
         n19824, n19825, n19826, n19827, n19828, n19829, n19830, n19831,
         n19832, n19833, n19834, n19835, n19836, n19837, n19838, n19839,
         n19840, n19841, n19842, n19843, n19844, n19845, n19846, n19847,
         n19848, n19849, n19850, n19851, n19852, n19853, n19854, n19855,
         n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19863,
         n19864, n19865, n19866, n19867, n19868, n19869, n19870, n19871,
         n19872, n19873, n19874, n19875, n19876, n19877, n19878, n19879,
         n19880, n19881, n19882, n19883, n19884, n19885, n19886, n19887,
         n19888, n19889, n19890, n19891, n19892, n19893, n19894, n19895,
         n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903,
         n19904, n19905, n19906, n19907, n19908, n19909, n19910, n19911,
         n19912, n19913, n19914, n19915, n19916, n19917, n19918, n19919,
         n19920, n19921, n19922, n19923, n19924, n19925, n19926, n19927,
         n19928, n19929, n19930, n19931, n19932, n19933, n19934, n19935,
         n19936, n19937, n19938, n19939, n19940, n19941, n19942, n19943,
         n19944, n19945, n19946, n19947, n19948, n19949, n19950, n19951,
         n19952, n19953, n19954, n19955, n19956, n19957, n19958, n19959,
         n19960, n19961, n19962, n19963, n19964, n19965, n19966, n19967,
         n19968, n19969, n19970, n19971, n19972, n19973, n19974, n19975,
         n19976, n19977, n19978, n19979, n19980, n19981, n19982, n19983,
         n19984, n19985, n19986, n19987, n19988, n19989, n19990, n19991,
         n19992, n19993, n19994, n19995, n19996, n19997, n19998, n19999,
         n20000, n20001, n20002, n20003, n20004, n20005, n20006, n20007,
         n20008, n20009, n20010, n20011, n20012, n20013, n20014, n20015,
         n20016, n20017, n20018, n20019, n20020, n20021, n20022, n20023,
         n20024, n20025, n20026, n20027, n20028, n20029, n20030, n20031,
         n20032, n20033, n20034, n20035, n20036, n20037, n20038, n20039,
         n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047,
         n20048, n20049, n20050, n20051, n20052, n20053, n20054, n20055,
         n20056, n20057, n20058, n20059, n20060, n20061, n20062, n20063,
         n20064, n20065, n20066, n20067, n20068, n20069, n20070, n20071,
         n20072, n20073, n20074, n20075, n20076, n20077, n20078, n20079,
         n20080, n20081, n20082, n20083, n20084, n20085, n20086, n20087,
         n20088, n20089, n20090, n20091, n20092, n20093, n20094, n20095,
         n20096, n20097, n20098, n20099, n20100, n20101, n20102, n20103,
         n20104, n20105, n20106, n20107, n20108, n20109, n20110, n20111,
         n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119,
         n20120, n20121, n20122, n20123, n20124, n20125, n20126, n20127,
         n20128, n20129, n20130, n20131, n20132, n20133, n20134, n20135,
         n20136, n20137, n20138, n20139, n20140, n20141, n20142, n20143,
         n20144, n20145, n20146, n20147, n20148, n20149, n20150, n20151,
         n20152, n20153, n20154, n20155, n20156, n20157, n20158, n20159,
         n20160, n20161, n20162, n20163, n20164, n20165, n20166, n20167,
         n20168, n20169, n20170, n20171, n20172, n20173, n20174, n20175,
         n20176, n20177, n20178, n20179, n20180, n20181, n20182, n20183,
         n20184, n20185, n20186, n20187, n20188, n20189, n20190, n20191,
         n20192, n20193, n20194, n20195, n20196, n20197, n20198, n20199,
         n20200, n20201, n20202, n20203, n20204, n20205, n20206, n20207,
         n20208, n20209, n20210, n20211, n20212, n20213, n20214, n20215,
         n20216, n20217, n20218, n20219, n20220, n20221, n20222, n20223,
         n20224, n20225, n20226, n20227, n20228, n20229, n20230, n20231,
         n20232, n20233, n20234, n20235, n20236, n20237, n20238, n20239,
         n20240, n20241, n20242, n20243, n20244, n20245, n20246, n20247,
         n20248, n20249, n20250, n20251, n20252, n20253, n20254, n20255,
         n20256, n20257, n20258, n20259, n20260, n20261, n20262, n20263,
         n20264, n20265, n20266, n20267, n20268, n20269, n20270, n20271,
         n20272, n20273, n20274, n20275, n20276, n20277, n20278, n20279,
         n20280, n20281, n20282, n20283, n20284, n20285, n20286, n20287,
         n20288, n20289, n20290, n20291, n20292, n20293, n20294, n20295,
         n20296, n20297, n20298, n20299, n20300, n20301, n20302, n20303,
         n20304, n20305, n20306, n20307, n20308, n20309, n20310, n20311,
         n20312, n20313, n20314, n20315, n20316, n20317, n20318, n20319,
         n20320, n20321, n20322, n20323, n20324, n20325, n20326, n20327,
         n20328, n20329, n20330, n20331, n20332, n20333, n20334, n20335,
         n20336, n20337, n20338, n20339, n20340, n20341, n20342, n20343,
         n20344, n20345, n20346, n20347, n20348, n20349, n20350, n20351,
         n20352, n20353, n20354, n20355, n20356, n20357, n20358, n20359,
         n20360, n20361, n20362, n20363, n20364, n20365, n20366, n20367,
         n20368, n20369, n20370, n20371, n20372, n20373, n20374, n20375,
         n20376, n20377, n20378, n20379, n20380, n20381, n20382, n20383,
         n20384, n20385, n20386, n20387, n20388, n20389, n20390, n20391,
         n20392, n20393, n20394, n20395, n20396, n20397, n20398, n20399,
         n20400, n20401, n20402, n20403, n20404, n20405, n20406, n20407,
         n20408, n20409, n20410, n20411, n20412, n20413, n20414, n20415,
         n20416, n20417, n20418, n20419, n20420, n20421, n20422, n20423,
         n20424, n20425, n20426, n20427, n20428, n20429, n20430, n20431,
         n20432, n20433, n20434, n20435, n20436, n20437, n20438, n20439,
         n20440, n20441, n20442, n20443, n20444, n20445, n20446, n20447,
         n20448, n20449, n20450, n20451, n20452, n20453, n20454, n20455,
         n20456, n20457, n20458, n20459, n20460, n20461, n20462, n20463,
         n20464, n20465, n20466, n20467, n20468, n20469, n20470, n20471,
         n20472, n20473, n20474, n20475, n20476, n20477, n20478, n20479,
         n20480, n20481, n20482, n20483, n20484, n20485, n20486, n20487,
         n20488, n20489, n20490, n20491, n20492, n20493, n20494, n20495,
         n20496, n20497, n20498, n20499, n20500, n20501, n20502, n20503,
         n20504, n20505, n20506, n20507, n20508, n20509, n20510, n20511,
         n20512, n20513, n20514, n20515, n20516, n20517, n20518, n20519,
         n20520, n20521, n20522, n20523, n20524, n20525, n20526, n20527,
         n20528, n20529, n20530, n20531, n20532, n20533, n20534, n20535,
         n20536, n20537, n20538, n20539, n20540, n20541, n20542, n20543,
         n20544, n20545, n20546, n20547, n20548, n20549, n20550, n20551,
         n20552, n20553, n20554, n20555, n20556, n20557, n20558, n20559,
         n20560, n20561, n20562, n20563, n20564, n20565, n20566, n20567,
         n20568, n20569, n20570, n20571, n20572, n20573, n20574, n20575,
         n20576, n20577, n20578, n20579, n20580, n20581, n20582, n20583,
         n20584, n20585, n20586, n20587, n20588, n20589, n20590, n20591,
         n20592, n20593, n20594, n20595, n20596, n20597, n20598, n20599,
         n20600, n20601, n20602, n20603, n20604, n20605, n20606, n20607,
         n20608, n20609, n20610, n20611, n20612, n20613, n20614, n20615,
         n20616, n20617, n20618, n20619, n20620, n20621, n20622, n20623,
         n20624, n20625, n20626, n20627, n20628, n20629, n20630, n20631,
         n20632, n20633, n20634, n20635, n20636, n20637, n20638, n20639,
         n20640, n20641, n20642, n20643, n20644, n20645, n20646, n20647,
         n20648, n20649, n20650, n20651, n20652, n20653, n20654, n20655,
         n20656, n20657, n20658, n20659, n20660, n20661, n20662, n20663,
         n20664, n20665, n20666, n20667, n20668, n20669, n20670, n20671,
         n20672, n20673, n20674, n20675, n20676, n20677, n20678, n20679,
         n20680, n20681, n20682, n20683, n20684, n20685, n20686, n20687,
         n20688, n20689, n20690, n20691, n20692, n20693, n20694, n20695,
         n20696, n20697, n20698, n20699, n20700, n20701, n20702, n20703,
         n20704, n20705, n20706, n20707, n20708, n20709, n20710, n20711,
         n20712, n20713, n20714, n20715, n20716, n20717, n20718, n20719,
         n20720, n20721, n20722, n20723, n20724, n20725, n20726, n20727,
         n20728, n20729, n20730, n20731, n20732, n20733, n20734, n20735,
         n20736, n20737, n20738, n20739, n20740, n20741, n20742, n20743,
         n20744, n20745, n20746, n20747, n20748, n20749, n20750, n20751,
         n20752, n20753, n20754, n20755, n20756, n20757, n20758, n20759,
         n20760, n20761, n20762, n20763, n20764, n20765, n20766, n20767,
         n20768, n20769, n20770, n20771, n20772, n20773, n20774, n20775,
         n20776, n20777, n20778, n20779, n20780, n20781, n20782, n20783,
         n20784, n20785, n20786, n20787, n20788, n20789, n20790, n20791,
         n20792, n20793, n20794, n20795, n20796, n20797, n20798, n20799,
         n20800, n20801, n20802, n20803, n20804, n20805, n20806, n20807,
         n20808, n20809, n20810, n20811, n20812, n20813, n20814, n20815,
         n20816, n20817, n20818, n20819, n20820, n20821, n20822, n20823,
         n20824, n20825, n20826, n20827, n20828, n20829, n20830, n20831,
         n20832, n20833, n20834, n20835, n20836, n20837, n20838, n20839,
         n20840, n20841, n20842, n20843, n20844, n20845, n20846, n20847,
         n20848, n20849, n20850, n20851, n20852, n20853, n20854, n20855,
         n20856, n20857, n20858, n20859, n20860, n20861, n20862, n20863,
         n20864, n20865, n20866, n20867, n20868, n20869, n20870, n20871,
         n20872, n20873, n20874, n20875, n20876, n20877, n20878, n20879,
         n20880, n20881, n20882, n20883, n20884, n20885, n20886, n20887,
         n20888, n20889, n20890, n20891, n20892, n20893, n20894, n20895,
         n20896, n20897, n20898, n20899, n20900, n20901, n20902, n20903,
         n20904, n20905, n20906, n20907, n20908, n20909, n20910, n20911,
         n20912, n20913, n20914, n20915, n20916, n20917, n20918, n20919,
         n20920, n20921, n20922, n20923, n20924, n20925, n20926, n20927,
         n20928, n20929, n20930, n20931, n20932, n20933, n20934, n20935,
         n20936, n20937, n20938, n20939, n20940, n20941, n20942, n20943,
         n20944, n20945, n20946, n20947, n20948, n20949, n20950, n20951,
         n20952, n20953, n20954, n20955, n20956, n20957, n20958, n20959,
         n20960, n20961, n20962, n20963, n20964, n20965, n20966, n20967,
         n20968, n20969, n20970, n20971, n20972, n20973, n20974, n20975,
         n20976, n20977, n20978, n20979, n20980, n20981, n20982, n20983,
         n20984, n20985, n20986, n20987, n20988, n20989, n20990, n20991,
         n20992, n20993, n20994, n20995, n20996, n20997, n20998, n20999,
         n21000, n21001, n21002, n21003, n21004, n21005, n21006, n21007,
         n21008, n21009, n21010, n21011, n21012, n21013, n21014, n21015,
         n21016, n21017, n21018, n21019, n21020, n21021, n21022, n21023,
         n21024, n21025, n21026, n21027, n21028, n21029, n21030, n21031,
         n21032, n21033, n21034, n21035, n21036, n21037, n21038, n21039,
         n21040, n21041, n21042, n21043, n21044, n21045, n21046, n21047,
         n21048, n21049, n21050, n21051, n21052, n21053, n21054, n21055,
         n21056, n21057, n21058, n21059, n21060, n21061, n21062, n21063,
         n21064, n21065, n21066, n21067, n21068, n21069, n21070, n21071,
         n21072, n21073, n21074, n21075, n21076, n21077, n21078, n21079,
         n21080, n21081, n21082, n21083, n21084, n21085, n21086, n21087,
         n21088, n21089, n21090, n21091, n21092, n21093, n21094, n21095,
         n21096, n21097, n21098, n21099, n21100, n21101, n21102, n21103,
         n21104, n21105, n21106, n21107, n21108, n21109, n21110, n21111,
         n21112, n21113, n21114, n21115, n21116, n21117, n21118, n21119,
         n21120, n21121, n21122, n21123, n21124, n21125, n21126, n21127,
         n21128, n21129, n21130, n21131, n21132, n21133, n21134, n21135,
         n21136, n21137, n21138, n21139, n21140, n21141, n21142, n21143,
         n21144, n21145, n21146, n21147, n21148, n21149, n21150, n21151,
         n21152, n21153, n21154, n21155, n21156, n21157, n21158, n21159,
         n21160, n21161, n21162, n21163, n21164, n21165, n21166, n21167,
         n21168, n21169, n21170, n21171, n21172, n21173, n21174, n21175,
         n21176, n21177, n21178, n21179, n21180, n21181, n21182, n21183,
         n21184, n21185, n21186, n21187, n21188, n21189, n21190, n21191,
         n21192, n21193, n21194, n21195, n21196, n21197, n21198, n21199,
         n21200, n21201, n21202, n21203, n21204, n21205, n21206, n21207,
         n21208, n21209, n21210, n21211, n21212, n21213, n21214, n21215,
         n21216, n21217, n21218, n21219, n21220, n21221, n21222, n21223,
         n21224, n21225, n21226, n21227, n21228, n21229, n21230, n21231,
         n21232, n21233, n21234, n21235, n21236, n21237, n21238, n21239,
         n21240, n21241, n21242, n21243, n21244, n21245, n21246, n21247,
         n21248, n21249, n21250, n21251, n21252, n21253, n21254, n21255,
         n21256, n21257, n21258, n21259, n21260, n21261, n21262, n21263,
         n21264, n21265, n21266, n21267, n21268, n21269, n21270, n21271,
         n21272, n21273, n21274, n21275, n21276, n21277, n21278, n21279,
         n21280, n21281, n21282, n21283, n21284, n21285, n21286, n21287,
         n21288, n21289, n21290, n21291, n21292, n21293, n21294, n21295,
         n21296, n21297, n21298, n21299, n21300, n21301, n21302, n21303,
         n21304, n21305, n21306, n21307, n21308, n21309, n21310, n21311,
         n21312, n21313, n21314, n21315, n21316, n21317, n21318, n21319,
         n21320, n21321, n21322, n21323, n21324, n21325, n21326, n21327,
         n21328, n21329, n21330, n21331, n21332, n21333, n21334, n21335,
         n21336, n21337, n21338, n21339, n21340, n21341, n21342, n21343,
         n21344, n21345, n21346, n21347, n21348, n21349, n21350, n21351,
         n21352, n21353, n21354, n21355, n21356, n21357, n21358, n21359,
         n21360, n21361, n21362, n21363, n21364, n21365, n21366, n21367,
         n21368, n21369, n21370, n21371, n21372, n21373, n21374, n21375,
         n21376, n21377, n21378, n21379, n21380, n21381, n21382, n21383,
         n21384, n21385, n21386, n21387, n21388, n21389, n21390, n21391,
         n21392, n21393, n21394, n21395, n21396, n21397, n21398, n21399,
         n21400, n21401, n21402, n21403, n21404, n21405, n21406, n21407,
         n21408, n21409, n21410, n21411, n21412, n21413, n21414, n21415,
         n21416, n21417, n21418, n21419, n21420, n21421, n21422, n21423,
         n21424, n21425, n21426, n21427, n21428, n21429, n21430, n21431,
         n21432, n21433, n21434, n21435, n21436, n21437, n21438, n21439,
         n21440, n21441, n21442, n21443, n21444, n21445, n21446, n21447,
         n21448, n21449, n21450, n21451, n21452, n21453, n21454, n21455,
         n21456, n21457, n21458, n21459, n21460, n21461, n21462, n21463,
         n21464, n21465, n21466, n21467, n21468, n21469, n21470, n21471,
         n21472, n21473, n21474, n21475, n21476, n21477, n21478, n21479,
         n21480, n21481, n21482, n21483, n21484, n21485, n21486, n21487,
         n21488, n21489, n21490, n21491, n21492, n21493, n21494, n21495,
         n21496, n21497, n21498, n21499, n21500, n21501, n21502, n21503,
         n21504, n21505, n21506, n21507, n21508, n21509, n21510, n21511,
         n21512, n21513, n21514, n21515, n21516, n21517, n21518, n21519,
         n21520, n21521, n21522, n21523, n21524, n21525, n21526, n21527,
         n21528, n21529, n21530, n21531, n21532, n21533, n21534, n21535,
         n21536, n21537, n21538, n21539, n21540, n21541, n21542, n21543,
         n21544, n21545, n21546, n21547, n21548, n21549, n21550, n21551,
         n21552, n21553, n21554, n21555, n21556, n21557, n21558, n21559,
         n21560, n21561, n21562, n21563, n21564, n21565, n21566, n21567,
         n21568, n21569, n21570, n21571, n21572, n21573, n21574, n21575,
         n21576, n21577, n21578, n21579, n21580, n21581, n21582, n21583,
         n21584, n21585, n21586, n21587, n21588, n21589, n21590, n21591,
         n21592, n21593, n21594, n21595, n21596, n21597, n21598, n21599,
         n21600, n21601, n21602, n21603, n21604, n21605, n21606, n21607,
         n21608, n21609, n21610, n21611, n21612, n21613, n21614, n21615,
         n21616, n21617, n21618, n21619, n21620, n21621, n21622, n21623,
         n21624, n21625, n21626, n21627, n21628, n21629, n21630, n21631,
         n21632, n21633, n21634, n21635, n21636, n21637, n21638, n21639,
         n21640, n21641, n21642, n21643, n21644, n21645, n21646, n21647,
         n21648, n21649, n21650, n21651, n21652, n21653, n21654, n21655,
         n21656, n21657, n21658, n21659, n21660, n21661, n21662, n21663,
         n21664, n21665, n21666, n21667, n21668, n21669, n21670, n21671,
         n21672, n21673, n21674, n21675, n21676, n21677, n21678, n21679,
         n21680, n21681, n21682, n21683, n21684, n21685, n21686, n21687,
         n21688, n21689, n21690, n21691, n21692, n21693, n21694, n21695,
         n21696, n21697, n21698, n21699, n21700, n21701, n21702, n21703,
         n21704, n21705, n21706, n21707, n21708, n21709, n21710, n21711,
         n21712, n21713, n21714, n21715, n21716, n21717, n21718, n21719,
         n21720, n21721, n21722, n21723, n21724, n21725, n21726, n21727,
         n21728, n21729, n21730, n21731, n21732, n21733, n21734, n21735,
         n21736, n21737, n21738, n21739, n21740, n21741, n21742, n21743,
         n21744, n21745, n21746, n21747, n21748, n21749, n21750, n21751,
         n21752, n21753, n21754, n21755, n21756, n21757, n21758, n21759,
         n21760, n21761, n21762, n21763, n21764, n21765, n21766, n21767,
         n21768, n21769, n21770, n21771, n21772, n21773, n21774, n21775,
         n21776, n21777, n21778, n21779, n21780, n21781, n21782, n21783,
         n21784, n21785, n21786, n21787, n21788, n21789, n21790, n21791,
         n21792, n21793, n21794, n21795, n21796, n21797, n21798, n21799,
         n21800, n21801, n21802, n21803, n21804, n21805, n21806, n21807,
         n21808, n21809, n21810, n21811, n21812, n21813, n21814, n21815,
         n21816, n21817, n21818, n21819, n21820, n21821, n21822, n21823,
         n21824, n21825, n21826, n21827, n21828, n21829, n21830, n21831,
         n21832, n21833, n21834, n21835, n21836, n21837, n21838, n21839,
         n21840, n21841, n21842, n21843, n21844, n21845, n21846, n21847,
         n21848, n21849, n21850, n21851, n21852, n21853, n21854, n21855,
         n21856, n21857, n21858, n21859, n21860, n21861, n21862, n21863,
         n21864, n21865, n21866, n21867, n21868, n21869, n21870, n21871,
         n21872, n21873, n21874, n21875, n21876, n21877, n21878, n21879,
         n21880, n21881, n21882, n21883, n21884, n21885, n21886, n21887,
         n21888, n21889, n21890, n21891, n21892, n21893, n21894, n21895,
         n21896, n21897, n21898, n21899, n21900, n21901, n21902, n21903,
         n21904, n21905, n21906, n21907, n21908, n21909, n21910, n21911,
         n21912, n21913, n21914, n21915, n21916, n21917, n21918, n21919,
         n21920, n21921, n21922, n21923, n21924, n21925, n21926, n21927,
         n21928, n21929, n21930, n21931, n21932, n21933, n21934, n21935,
         n21936, n21937, n21938, n21939, n21940, n21941, n21942, n21943,
         n21944, n21945, n21946, n21947, n21948, n21949, n21950, n21951,
         n21952, n21953, n21954, n21955, n21956, n21957, n21958, n21959,
         n21960, n21961, n21962, n21963, n21964, n21965, n21966, n21967,
         n21968, n21969, n21970, n21971, n21972, n21973, n21974, n21975,
         n21976, n21977, n21978, n21979, n21980, n21981, n21982, n21983,
         n21984, n21985, n21986, n21987, n21988, n21989, n21990, n21991,
         n21992, n21993, n21994, n21995, n21996, n21997, n21998, n21999,
         n22000, n22001, n22002, n22003, n22004, n22005, n22006, n22007,
         n22008, n22009, n22010, n22011, n22012, n22013, n22014, n22015,
         n22016, n22017, n22018, n22019, n22020, n22021, n22022, n22023,
         n22024, n22025, n22026, n22027, n22028, n22029, n22030, n22031,
         n22032, n22033, n22034, n22035, n22036, n22037, n22038, n22039,
         n22040, n22041, n22042, n22043, n22044, n22045, n22046, n22047,
         n22048, n22049, n22050, n22051, n22052, n22053, n22054, n22055,
         n22056, n22057, n22058, n22059, n22060, n22061, n22062, n22063,
         n22064, n22065, n22066, n22067, n22068, n22069, n22070, n22071,
         n22072, n22073, n22074, n22075, n22076, n22077, n22078, n22079,
         n22080, n22081, n22082, n22083, n22084, n22085, n22086, n22087,
         n22088, n22089, n22090, n22091, n22092, n22093, n22094, n22095,
         n22096, n22097, n22098, n22099, n22100, n22101, n22102, n22103,
         n22104, n22105, n22106, n22107, n22108, n22109, n22110, n22111,
         n22112, n22113, n22114, n22115, n22116, n22117, n22118, n22119,
         n22120, n22121, n22122, n22123, n22124, n22125, n22126, n22127,
         n22128, n22129, n22130, n22131, n22132, n22133, n22134, n22135,
         n22136, n22137, n22138, n22139, n22140, n22141, n22142, n22143,
         n22144, n22145, n22146, n22147, n22148, n22149, n22150, n22151,
         n22152, n22153, n22154, n22155, n22156, n22157, n22158, n22159,
         n22160, n22161, n22162, n22163, n22164, n22165, n22166, n22167,
         n22168, n22169, n22170, n22171, n22172, n22173, n22174, n22175,
         n22176, n22177, n22178, n22179, n22180, n22181, n22182, n22183,
         n22184, n22185, n22186, n22187, n22188, n22189, n22190, n22191,
         n22192, n22193, n22194, n22195, n22196, n22197, n22198, n22199,
         n22200, n22201, n22202, n22203, n22204, n22205, n22206, n22207,
         n22208, n22209, n22210, n22211, n22212, n22213, n22214, n22215,
         n22216, n22217, n22218, n22219, n22220, n22221, n22222, n22223,
         n22224, n22225, n22226, n22227, n22228, n22229, n22230, n22231,
         n22232, n22233, n22234, n22235, n22236, n22237, n22238, n22239,
         n22240, n22241, n22242, n22243, n22244, n22245, n22246, n22247,
         n22248, n22249, n22250, n22251, n22252, n22253, n22254, n22255,
         n22256, n22257, n22258, n22259, n22260, n22261, n22262, n22263,
         n22264, n22265, n22266, n22267, n22268, n22269, n22270, n22271,
         n22272, n22273, n22274, n22275, n22276, n22277, n22278, n22279,
         n22280, n22281, n22282, n22283, n22284, n22285, n22286, n22287,
         n22288, n22289, n22290, n22291, n22292, n22293, n22294, n22295,
         n22296, n22297, n22298, n22299, n22300, n22301, n22302, n22303,
         n22304, n22305, n22306, n22307, n22308, n22309, n22310, n22311,
         n22312, n22313, n22314, n22315, n22316, n22317, n22318, n22319,
         n22320, n22321, n22322, n22323, n22324, n22325, n22326, n22327,
         n22328, n22329, n22330, n22331, n22332, n22333, n22334, n22335,
         n22336, n22337, n22338, n22339, n22340, n22341, n22342, n22343,
         n22344, n22345, n22346, n22347, n22348, n22349, n22350, n22351,
         n22352, n22353, n22354, n22355, n22356, n22357, n22358, n22359,
         n22360, n22361, n22362, n22363, n22364, n22365, n22366, n22367,
         n22368, n22369, n22370, n22371, n22372, n22373, n22374, n22375,
         n22376, n22377, n22378, n22379, n22380, n22381, n22382, n22383,
         n22384, n22385, n22386, n22387, n22388, n22389, n22390, n22391,
         n22392, n22393, n22394, n22395, n22396, n22397, n22398, n22399,
         n22400, n22401, n22402, n22403, n22404, n22405, n22406, n22407,
         n22408, n22409, n22410, n22411, n22412, n22413, n22414, n22415,
         n22416, n22417, n22418, n22419, n22420, n22421, n22422, n22423,
         n22424, n22425, n22426, n22427, n22428, n22429, n22430, n22431,
         n22432, n22433, n22434, n22435, n22436, n22437, n22438, n22439,
         n22440, n22441, n22442, n22443, n22444, n22445, n22446, n22447,
         n22448, n22449, n22450, n22451, n22452, n22453, n22454, n22455,
         n22456, n22457, n22458, n22459, n22460, n22461, n22462, n22463,
         n22464, n22465, n22466, n22467, n22468, n22469, n22470, n22471,
         n22472, n22473, n22474, n22475, n22476, n22477, n22478, n22479,
         n22480, n22481, n22482, n22483, n22484, n22485, n22486, n22487,
         n22488, n22489, n22490, n22491, n22492, n22493, n22494, n22495,
         n22496, n22497, n22498, n22499, n22500, n22501, n22502, n22503,
         n22504, n22505, n22506, n22507, n22508, n22509, n22510, n22511,
         n22512, n22513, n22514, n22515, n22516, n22517, n22518, n22519,
         n22520, n22521, n22522, n22523, n22524, n22525, n22526, n22527,
         n22528, n22529, n22530, n22531, n22532, n22533, n22534, n22535,
         n22536, n22537, n22538, n22539, n22540, n22541, n22542, n22543,
         n22544, n22545, n22546, n22547, n22548, n22549, n22550, n22551,
         n22552, n22553, n22554, n22555, n22556, n22557, n22558, n22559,
         n22560, n22561, n22562, n22563, n22564, n22565, n22566, n22567,
         n22568, n22569, n22570, n22571, n22572, n22573, n22574, n22575,
         n22576, n22577, n22578, n22579, n22580, n22581, n22582, n22583,
         n22584, n22585, n22586, n22587, n22588, n22589, n22590, n22591,
         n22592, n22593, n22594, n22595, n22596, n22597, n22598, n22599,
         n22600, n22601, n22602, n22603, n22604, n22605, n22606, n22607,
         n22608, n22609, n22610, n22611, n22612, n22613, n22614, n22615,
         n22616, n22617, n22618, n22619, n22620, n22621, n22622, n22623,
         n22624, n22625, n22626, n22627, n22628, n22629, n22630, n22631,
         n22632, n22633, n22634, n22635, n22636, n22637, n22638, n22639,
         n22640, n22641, n22642, n22643, n22644, n22645, n22646, n22647,
         n22648, n22649, n22650, n22651, n22652, n22653, n22654, n22655,
         n22656, n22657, n22658, n22659, n22660, n22661, n22662, n22663,
         n22664, n22665, n22666, n22667, n22668, n22669, n22670, n22671,
         n22672, n22673, n22674, n22675, n22676, n22677, n22678, n22679,
         n22680, n22681, n22682, n22683, n22684, n22685, n22686, n22687,
         n22688, n22689, n22690, n22691, n22692, n22693, n22694, n22695,
         n22696, n22697, n22698, n22699, n22700, n22701, n22702, n22703,
         n22704, n22705, n22706, n22707, n22708, n22709, n22710, n22711,
         n22712, n22713, n22714, n22715, n22716, n22717, n22718, n22719,
         n22720, n22721, n22722, n22723, n22724, n22725, n22726, n22727,
         n22728, n22729, n22730, n22731, n22732, n22733, n22734, n22735,
         n22736, n22737, n22738, n22739, n22740, n22741, n22742, n22743,
         n22744, n22745, n22746, n22747, n22748, n22749, n22750, n22751,
         n22752, n22753, n22754, n22755, n22756, n22757, n22758, n22759,
         n22760, n22761, n22762, n22763, n22764, n22765, n22766, n22767,
         n22768, n22769, n22770, n22771, n22772, n22773, n22774, n22775,
         n22776, n22777, n22778, n22779, n22780, n22781, n22782, n22783,
         n22784, n22785, n22786, n22787, n22788, n22789, n22790, n22791,
         n22792, n22793, n22794, n22795, n22796, n22797, n22798, n22799,
         n22800, n22801, n22802, n22803, n22804, n22805, n22806, n22807,
         n22808, n22809, n22810, n22811, n22812, n22813, n22814, n22815,
         n22816, n22817, n22818, n22819, n22820, n22821, n22822, n22823,
         n22824, n22825, n22826, n22827, n22828, n22829, n22830, n22831,
         n22832, n22833, n22834, n22835, n22836, n22837, n22838, n22839,
         n22840, n22841, n22842, n22843, n22844, n22845, n22846, n22847,
         n22848, n22849, n22850, n22851, n22852, n22853, n22854, n22855,
         n22856, n22857, n22858, n22859, n22860, n22861, n22862, n22863,
         n22864, n22865, n22866, n22867, n22868, n22869, n22870, n22871,
         n22872, n22873, n22874, n22875, n22876, n22877, n22878, n22879,
         n22880, n22881, n22882, n22883, n22884, n22885, n22886, n22887,
         n22888, n22889, n22890, n22891, n22892, n22893, n22894, n22895,
         n22896, n22897, n22898, n22899, n22900, n22901, n22902, n22903,
         n22904, n22905, n22906, n22907, n22908, n22909, n22910, n22911,
         n22912, n22913, n22914, n22915, n22916, n22917, n22918, n22919,
         n22920, n22921, n22922, n22923, n22924, n22925, n22926, n22927,
         n22928, n22929, n22930, n22931, n22932, n22933, n22934, n22935,
         n22936, n22937, n22938, n22939, n22940, n22941, n22942, n22943,
         n22944, n22945, n22946, n22947, n22948, n22949, n22950, n22951,
         n22952, n22953, n22954, n22955, n22956, n22957, n22958, n22959,
         n22960, n22961, n22962, n22963, n22964, n22965, n22966, n22967,
         n22968, n22969, n22970, n22971, n22972, n22973, n22974, n22975,
         n22976, n22977, n22978, n22979, n22980, n22981, n22982, n22983,
         n22984, n22985, n22986, n22987, n22988, n22989, n22990, n22991,
         n22992, n22993, n22994, n22995, n22996, n22997, n22998, n22999,
         n23000, n23001, n23002, n23003, n23004, n23005, n23006, n23007,
         n23008, n23009, n23010, n23011, n23012, n23013, n23014, n23015,
         n23016, n23017, n23018, n23019, n23020, n23021, n23022, n23023,
         n23024, n23025, n23026, n23027, n23028, n23029, n23030, n23031,
         n23032, n23033, n23034, n23035, n23036, n23037, n23038, n23039,
         n23040, n23041, n23042, n23043, n23044, n23045, n23046, n23047,
         n23048, n23049, n23050, n23051, n23052, n23053, n23054, n23055,
         n23056, n23057, n23058, n23059, n23060, n23061, n23062, n23063,
         n23064, n23065, n23066, n23067, n23068, n23069, n23070, n23071,
         n23072, n23073, n23074, n23075, n23076, n23077, n23078, n23079,
         n23080, n23081, n23082, n23083, n23084, n23085, n23086, n23087,
         n23088, n23089, n23090, n23091, n23092, n23093, n23094, n23095,
         n23096, n23097, n23098, n23099, n23100, n23101, n23102, n23103,
         n23104, n23105, n23106, n23107, n23108, n23109, n23110, n23111,
         n23112, n23113, n23114, n23115, n23116, n23117, n23118, n23119,
         n23120, n23121, n23122, n23123, n23124, n23125, n23126, n23127,
         n23128, n23129, n23130, n23131, n23132, n23133, n23134, n23135,
         n23136, n23137, n23138, n23139, n23140, n23141, n23142, n23143,
         n23144, n23145, n23146, n23147, n23148, n23149, n23150, n23151,
         n23152, n23153, n23154, n23155, n23156, n23157, n23158, n23159,
         n23160, n23161, n23162, n23163, n23164, n23165, n23166, n23167,
         n23168, n23169, n23170, n23171, n23172, n23173, n23174, n23175,
         n23176, n23177, n23178, n23179, n23180, n23181, n23182, n23183,
         n23184, n23185, n23186, n23187, n23188, n23189, n23190, n23191,
         n23192, n23193, n23194, n23195, n23196, n23197, n23198, n23199,
         n23200, n23201, n23202, n23203, n23204, n23205, n23206, n23207,
         n23208, n23209, n23210, n23211, n23212, n23213, n23214, n23215,
         n23216, n23217, n23218, n23219, n23220, n23221, n23222, n23223,
         n23224, n23225, n23226, n23227, n23228, n23229, n23230, n23231,
         n23232, n23233, n23234, n23235, n23236, n23237, n23238, n23239,
         n23240, n23241, n23242, n23243, n23244, n23245, n23246, n23247,
         n23248, n23249, n23250, n23251, n23252, n23253, n23254, n23255,
         n23256, n23257, n23258, n23259, n23260, n23261, n23262, n23263,
         n23264, n23265, n23266, n23267, n23268, n23269, n23270, n23271,
         n23272, n23273, n23274, n23275, n23276, n23277, n23278, n23279,
         n23280, n23281, n23282, n23283, n23284, n23285, n23286, n23287,
         n23288, n23289, n23290, n23291, n23292, n23293, n23294, n23295,
         n23296, n23297, n23298, n23299, n23300, n23301, n23302, n23303,
         n23304, n23305, n23306, n23307, n23308, n23309, n23310, n23311,
         n23312, n23313, n23314, n23315, n23316, n23317, n23318, n23319,
         n23320, n23321, n23322, n23323, n23324, n23325, n23326, n23327,
         n23328, n23329, n23330, n23331, n23332, n23333, n23334, n23335,
         n23336, n23337, n23338, n23339, n23340, n23341, n23342, n23343,
         n23344, n23345, n23346, n23347, n23348, n23349, n23350, n23351,
         n23352, n23353, n23354, n23355, n23356, n23357, n23358, n23359,
         n23360, n23361, n23362, n23363, n23364, n23365, n23366, n23367,
         n23368, n23369, n23370, n23371, n23372, n23373, n23374, n23375,
         n23376, n23377, n23378, n23379, n23380, n23381, n23382, n23383,
         n23384, n23385, n23386, n23387, n23388, n23389, n23390, n23391,
         n23392, n23393, n23394, n23395, n23396, n23397, n23398, n23399,
         n23400, n23401, n23402, n23403, n23404, n23405, n23406, n23407,
         n23408, n23409, n23410, n23411, n23412, n23413, n23414, n23415,
         n23416, n23417, n23418, n23419, n23420, n23421, n23422, n23423,
         n23424, n23425, n23426, n23427, n23428, n23429, n23430, n23431,
         n23432, n23433, n23434, n23435, n23436, n23437, n23438, n23439,
         n23440, n23441, n23442, n23443, n23444, n23445, n23446, n23447,
         n23448, n23449, n23450, n23451, n23452, n23453, n23454, n23455,
         n23456, n23457, n23458, n23459, n23460, n23461, n23462, n23463,
         n23464, n23465, n23466, n23467, n23468, n23469, n23470, n23471,
         n23472, n23473, n23474, n23475, n23476, n23477, n23478, n23479,
         n23480, n23481, n23482, n23483, n23484, n23485, n23486, n23487,
         n23488, n23489, n23490, n23491, n23492, n23493, n23494, n23495,
         n23496, n23497, n23498, n23499, n23500, n23501, n23502, n23503,
         n23504, n23505, n23506, n23507, n23508, n23509, n23510, n23511,
         n23512, n23513, n23514, n23515, n23516, n23517, n23518, n23519,
         n23520, n23521, n23522, n23523, n23524, n23525, n23526, n23527,
         n23528, n23529, n23530, n23531, n23532, n23533, n23534, n23535,
         n23536, n23537, n23538, n23539, n23540, n23541, n23542, n23543,
         n23544, n23545, n23546, n23547, n23548, n23549, n23550, n23551,
         n23552, n23553, n23554, n23555, n23556, n23557, n23558, n23559,
         n23560, n23561, n23562, n23563, n23564, n23565, n23566, n23567,
         n23568, n23569, n23570, n23571, n23572, n23573, n23574, n23575,
         n23576, n23577, n23578, n23579, n23580, n23581, n23582, n23583,
         n23584, n23585, n23586, n23587, n23588, n23589, n23590, n23591,
         n23592, n23593, n23594, n23595, n23596, n23597, n23598, n23599,
         n23600, n23601, n23602, n23603, n23604, n23605, n23606, n23607,
         n23608, n23609, n23610, n23611, n23612, n23613, n23614, n23615,
         n23616, n23617, n23618, n23619, n23620, n23621, n23622, n23623,
         n23624, n23625, n23626, n23627, n23628, n23629, n23630, n23631,
         n23632, n23633, n23634, n23635, n23636, n23637, n23638, n23639,
         n23640, n23641, n23642, n23643, n23644, n23645, n23646, n23647,
         n23648, n23649, n23650, n23651, n23652, n23653, n23654, n23655,
         n23656, n23657, n23658, n23659, n23660, n23661, n23662, n23663,
         n23664, n23665, n23666, n23667, n23668, n23669, n23670, n23671,
         n23672, n23673, n23674, n23675, n23676, n23677, n23678, n23679,
         n23680, n23681, n23682, n23683, n23684, n23685, n23686, n23687,
         n23688, n23689, n23690, n23691, n23692, n23693, n23694, n23695,
         n23696, n23697, n23698, n23699, n23700, n23701, n23702, n23703,
         n23704, n23705, n23706, n23707, n23708, n23709, n23710, n23711,
         n23712, n23713, n23714, n23715, n23716, n23717, n23718, n23719,
         n23720, n23721, n23722, n23723, n23724, n23725, n23726, n23727,
         n23728, n23729, n23730, n23731, n23732, n23733, n23734, n23735,
         n23736, n23737, n23738, n23739, n23740, n23741, n23742, n23743,
         n23744, n23745, n23746, n23747, n23748, n23749, n23750, n23751,
         n23752, n23753, n23754, n23755, n23756, n23757, n23758, n23759,
         n23760, n23761, n23762, n23763, n23764, n23765, n23766, n23767,
         n23768, n23769, n23770, n23771, n23772, n23773, n23774, n23775,
         n23776, n23777, n23778, n23779, n23780, n23781, n23782, n23783,
         n23784, n23785, n23786, n23787, n23788, n23789, n23790, n23791,
         n23792, n23793, n23794, n23795, n23796, n23797, n23798, n23799,
         n23800, n23801, n23802, n23803, n23804, n23805, n23806, n23807,
         n23808, n23809, n23810, n23811, n23812, n23813, n23814, n23815,
         n23816, n23817, n23818, n23819, n23820, n23821, n23822, n23823,
         n23824, n23825, n23826, n23827, n23828, n23829, n23830, n23831,
         n23832, n23833, n23834, n23835, n23836, n23837, n23838, n23839,
         n23840, n23841, n23842, n23843, n23844, n23845, n23846, n23847,
         n23848, n23849, n23850, n23851, n23852, n23853, n23854, n23855,
         n23856, n23857, n23858, n23859, n23860, n23861, n23862, n23863,
         n23864, n23865, n23866, n23867, n23868, n23869, n23870, n23871,
         n23872, n23873, n23874, n23875, n23876, n23877, n23878, n23879,
         n23880, n23881, n23882, n23883, n23884, n23885, n23886, n23887,
         n23888, n23889, n23890, n23891, n23892, n23893, n23894, n23895,
         n23896, n23897, n23898, n23899, n23900, n23901, n23902, n23903,
         n23904, n23905, n23906, n23907, n23908, n23909, n23910, n23911,
         n23912, n23913, n23914, n23915, n23916, n23917, n23918, n23919,
         n23920, n23921, n23922, n23923, n23924, n23925, n23926, n23927,
         n23928, n23929, n23930, n23931, n23932, n23933, n23934, n23935,
         n23936, n23937, n23938, n23939, n23940, n23941, n23942, n23943,
         n23944, n23945, n23946, n23947, n23948, n23949, n23950, n23951,
         n23952, n23953, n23954, n23955, n23956, n23957, n23958, n23959,
         n23960, n23961, n23962, n23963, n23964, n23965, n23966, n23967,
         n23968, n23969, n23970, n23971, n23972, n23973, n23974, n23975,
         n23976, n23977, n23978, n23979, n23980, n23981, n23982, n23983,
         n23984, n23985, n23986, n23987, n23988, n23989, n23990, n23991,
         n23992, n23993, n23994, n23995, n23996, n23997, n23998, n23999,
         n24000, n24001, n24002, n24003, n24004, n24005, n24006, n24007,
         n24008, n24009, n24010, n24011, n24012, n24013, n24014, n24015,
         n24016, n24017, n24018, n24019, n24020, n24021, n24022, n24023,
         n24024, n24025, n24026, n24027, n24028, n24029, n24030, n24031,
         n24032, n24033, n24034, n24035, n24036, n24037, n24038, n24039,
         n24040, n24041, n24042, n24043, n24044, n24045, n24046, n24047,
         n24048, n24049, n24050, n24051, n24052, n24053, n24054, n24055,
         n24056, n24057, n24058, n24059, n24060, n24061, n24062, n24063,
         n24064, n24065, n24066, n24067, n24068, n24069, n24070, n24071,
         n24072, n24073, n24074, n24075, n24076, n24077, n24078, n24079,
         n24080, n24081, n24082, n24083, n24084, n24085, n24086, n24087,
         n24088, n24089, n24090, n24091, n24092, n24093, n24094, n24095,
         n24096, n24097, n24098, n24099, n24100, n24101, n24102, n24103,
         n24104, n24105, n24106, n24107, n24108, n24109, n24110, n24111,
         n24112, n24113, n24114, n24115, n24116, n24117, n24118, n24119,
         n24120, n24121, n24122, n24123, n24124, n24125, n24126, n24127,
         n24128, n24129, n24130, n24131, n24132, n24133, n24134, n24135,
         n24136, n24137, n24138, n24139, n24140, n24141, n24142, n24143,
         n24144, n24145, n24146, n24147, n24148, n24149, n24150, n24151,
         n24152, n24153, n24154, n24155, n24156, n24157, n24158, n24159,
         n24160, n24161, n24162, n24163, n24164, n24165, n24166, n24167,
         n24168, n24169, n24170, n24171, n24172, n24173, n24174, n24175,
         n24176, n24177, n24178, n24179, n24180, n24181, n24182, n24183,
         n24184, n24185, n24186, n24187, n24188, n24189, n24190, n24191,
         n24192, n24193, n24194, n24195, n24196, n24197, n24198, n24199,
         n24200, n24201, n24202, n24203, n24204, n24205, n24206, n24207,
         n24208, n24209, n24210, n24211, n24212, n24213, n24214, n24215,
         n24216, n24217, n24218, n24219, n24220, n24221, n24222, n24223,
         n24224, n24225, n24226, n24227, n24228, n24229, n24230, n24231,
         n24232, n24233, n24234, n24235, n24236, n24237, n24238, n24239,
         n24240, n24241, n24242, n24243, n24244, n24245, n24246, n24247,
         n24248, n24249, n24250, n24251, n24252, n24253, n24254, n24255,
         n24256, n24257, n24258, n24259, n24260, n24261, n24262, n24263,
         n24264, n24265, n24266, n24267, n24268, n24269, n24270, n24271,
         n24272, n24273, n24274, n24275, n24276, n24277, n24278, n24279,
         n24280, n24281, n24282, n24283, n24284, n24285, n24286, n24287,
         n24288, n24289, n24290, n24291, n24292, n24293, n24294, n24295,
         n24296, n24297, n24298, n24299, n24300, n24301, n24302, n24303,
         n24304, n24305, n24306, n24307, n24308, n24309, n24310, n24311,
         n24312, n24313, n24314, n24315, n24316, n24317, n24318, n24319,
         n24320, n24321, n24322, n24323, n24324, n24325, n24326, n24327,
         n24328, n24329, n24330, n24331, n24332, n24333, n24334, n24335,
         n24336, n24337, n24338, n24339, n24340, n24341, n24342, n24343,
         n24344, n24345, n24346, n24347, n24348, n24349, n24350, n24351,
         n24352, n24353, n24354, n24355, n24356, n24357, n24358, n24359,
         n24360, n24361, n24362, n24363, n24364, n24365, n24366, n24367,
         n24368, n24369, n24370, n24371, n24372, n24373, n24374, n24375,
         n24376, n24377, n24378, n24379, n24380, n24381, n24382, n24383,
         n24384, n24385, n24386, n24387, n24388, n24389, n24390, n24391,
         n24392, n24393, n24394, n24395, n24396, n24397, n24398, n24399,
         n24400, n24401, n24402, n24403, n24404, n24405, n24406, n24407,
         n24408, n24409, n24410, n24411, n24412, n24413, n24414, n24415,
         n24416, n24417, n24418, n24419, n24420, n24421, n24422, n24423,
         n24424, n24425, n24426, n24427, n24428, n24429, n24430, n24431,
         n24432, n24433, n24434, n24435, n24436, n24437, n24438, n24439,
         n24440, n24441, n24442, n24443, n24444, n24445, n24446, n24447,
         n24448, n24449, n24450, n24451, n24452, n24453, n24454, n24455,
         n24456, n24457, n24458, n24459, n24460, n24461, n24462, n24463,
         n24464, n24465, n24466, n24467, n24468, n24469, n24470, n24471,
         n24472, n24473, n24474, n24475, n24476, n24477, n24478, n24479,
         n24480, n24481, n24482, n24483, n24484, n24485, n24486, n24487,
         n24488, n24489, n24490, n24491, n24492, n24493, n24494, n24495,
         n24496, n24497, n24498, n24499, n24500, n24501, n24502, n24503,
         n24504, n24505, n24506, n24507, n24508, n24509, n24510, n24511,
         n24512, n24513, n24514, n24515, n24516, n24517, n24518, n24519,
         n24520, n24521, n24522, n24523, n24524, n24525, n24526, n24527,
         n24528, n24529, n24530, n24531, n24532, n24533, n24534, n24535,
         n24536, n24537, n24538, n24539, n24540, n24541, n24542, n24543,
         n24544, n24545, n24546, n24547, n24548, n24549, n24550, n24551,
         n24552, n24553, n24554, n24555, n24556, n24557, n24558, n24559,
         n24560, n24561, n24562, n24563, n24564, n24565, n24566, n24567,
         n24568, n24569, n24570, n24571, n24572, n24573, n24574, n24575,
         n24576, n24577, n24578, n24579, n24580, n24581, n24582, n24583,
         n24584, n24585, n24586, n24587, n24588, n24589, n24590, n24591,
         n24592, n24593, n24594, n24595, n24596, n24597, n24598, n24599,
         n24600, n24601, n24602, n24603, n24604, n24605, n24606, n24607,
         n24608, n24609, n24610, n24611, n24612, n24613, n24614, n24615,
         n24616, n24617, n24618, n24619, n24620, n24621, n24622, n24623,
         n24624, n24625, n24626, n24627, n24628, n24629, n24630, n24631,
         n24632, n24633, n24634, n24635, n24636, n24637, n24638, n24639,
         n24640, n24641, n24642, n24643, n24644, n24645, n24646, n24647,
         n24648, n24649, n24650, n24651, n24652, n24653, n24654, n24655,
         n24656, n24657, n24658, n24659, n24660, n24661, n24662, n24663,
         n24664, n24665, n24666, n24667, n24668, n24669, n24670, n24671,
         n24672, n24673, n24674, n24675, n24676, n24677, n24678, n24679,
         n24680, n24681, n24682, n24683, n24684, n24685, n24686, n24687,
         n24688, n24689, n24690, n24691, n24692, n24693, n24694, n24695,
         n24696, n24697, n24698, n24699, n24700, n24701, n24702, n24703,
         n24704, n24705, n24706, n24707, n24708, n24709, n24710, n24711,
         n24712, n24713, n24714, n24715, n24716, n24717, n24718, n24719,
         n24720, n24721, n24722, n24723, n24724, n24725, n24726, n24727,
         n24728, n24729, n24730, n24731, n24732, n24733, n24734, n24735,
         n24736, n24737, n24738, n24739, n24740, n24741, n24742, n24743,
         n24744, n24745, n24746, n24747, n24748, n24749, n24750, n24751,
         n24752, n24753, n24754, n24755, n24756, n24757, n24758, n24759,
         n24760, n24761, n24762, n24763, n24764, n24765, n24766, n24767,
         n24768, n24769, n24770, n24771, n24772, n24773, n24774, n24775,
         n24776, n24777, n24778, n24779, n24780, n24781, n24782, n24783,
         n24784, n24785, n24786, n24787, n24788, n24789, n24790, n24791,
         n24792, n24793, n24794, n24795, n24796, n24797, n24798, n24799,
         n24800, n24801, n24802, n24803, n24804, n24805, n24806, n24807,
         n24808, n24809, n24810, n24811, n24812, n24813, n24814, n24815,
         n24816, n24817, n24818, n24819, n24820, n24821, n24822, n24823,
         n24824, n24825, n24826, n24827, n24828, n24829, n24830, n24831,
         n24832, n24833, n24834, n24835, n24836, n24837, n24838, n24839,
         n24840, n24841, n24842, n24843, n24844, n24845, n24846, n24847,
         n24848, n24849, n24850, n24851, n24852, n24853, n24854, n24855,
         n24856, n24857, n24858, n24859, n24860, n24861, n24862, n24863,
         n24864, n24865, n24866, n24867, n24868, n24869, n24870, n24871,
         n24872, n24873, n24874, n24875, n24876, n24877, n24878, n24879,
         n24880, n24881, n24882, n24883, n24884, n24885, n24886, n24887,
         n24888, n24889, n24890, n24891, n24892, n24893, n24894, n24895,
         n24896, n24897, n24898, n24899, n24900, n24901, n24902, n24903,
         n24904, n24905, n24906, n24907, n24908, n24909, n24910, n24911,
         n24912, n24913, n24914, n24915, n24916, n24917, n24918, n24919,
         n24920, n24921, n24922, n24923, n24924, n24925, n24926, n24927,
         n24928, n24929, n24930, n24931, n24932, n24933, n24934, n24935,
         n24936, n24937, n24938, n24939, n24940, n24941, n24942, n24943,
         n24944, n24945, n24946, n24947, n24948, n24949, n24950, n24951,
         n24952, n24953, n24954, n24955, n24956, n24957, n24958, n24959,
         n24960, n24961, n24962, n24963, n24964, n24965, n24966, n24967,
         n24968, n24969, n24970, n24971, n24972, n24973, n24974, n24975,
         n24976, n24977, n24978, n24979, n24980, n24981, n24982, n24983,
         n24984, n24985, n24986, n24987, n24988, n24989, n24990, n24991,
         n24992, n24993, n24994, n24995, n24996, n24997, n24998, n24999,
         n25000, n25001, n25002, n25003, n25004, n25005, n25006, n25007,
         n25008, n25009, n25010, n25011, n25012, n25013, n25014, n25015,
         n25016, n25017, n25018, n25019, n25020, n25021, n25022, n25023,
         n25024, n25025, n25026, n25027, n25028, n25029, n25030, n25031,
         n25032, n25033, n25034, n25035, n25036, n25037, n25038, n25039,
         n25040, n25041, n25042, n25043, n25044, n25045, n25046, n25047,
         n25048, n25049, n25050, n25051, n25052, n25053, n25054, n25055,
         n25056, n25057, n25058, n25059, n25060, n25061, n25062, n25063,
         n25064, n25065, n25066, n25067, n25068, n25069, n25070, n25071,
         n25072, n25073, n25074, n25075, n25076, n25077, n25078, n25079,
         n25080, n25081, n25082, n25083, n25084, n25085, n25086, n25087,
         n25088, n25089, n25090, n25091, n25092, n25093, n25094, n25095,
         n25096, n25097, n25098, n25099, n25100, n25101, n25102, n25103,
         n25104, n25105, n25106, n25107, n25108, n25109, n25110, n25111,
         n25112, n25113, n25114, n25115, n25116, n25117, n25118, n25119,
         n25120, n25121, n25122, n25123, n25124, n25125, n25126, n25127,
         n25128, n25129, n25130, n25131, n25132, n25133, n25134, n25135,
         n25136, n25137, n25138, n25139, n25140, n25141, n25142, n25143,
         n25144, n25145, n25146, n25147, n25148, n25149, n25150, n25151,
         n25152, n25153, n25154, n25155, n25156, n25157, n25158, n25159,
         n25160, n25161, n25162, n25163, n25164, n25165, n25166, n25167,
         n25168, n25169, n25170, n25171, n25172, n25173, n25174, n25175,
         n25176, n25177, n25178, n25179, n25180, n25181, n25182, n25183,
         n25184, n25185, n25186, n25187, n25188, n25189, n25190, n25191,
         n25192, n25193, n25194, n25195, n25196, n25197, n25198, n25199,
         n25200, n25201, n25202, n25203, n25204, n25205, n25206, n25207,
         n25208, n25209, n25210, n25211, n25212, n25213, n25214, n25215,
         n25216, n25217, n25218, n25219, n25220, n25221, n25222, n25223,
         n25224, n25225, n25226, n25227, n25228, n25229, n25230, n25231,
         n25232, n25233, n25234, n25235, n25236, n25237, n25238, n25239,
         n25240, n25241, n25242, n25243, n25244, n25245, n25246, n25247,
         n25248, n25249, n25250, n25251, n25252, n25253, n25254, n25255,
         n25256, n25257, n25258, n25259, n25260, n25261, n25262, n25263,
         n25264, n25265, n25266, n25267, n25268, n25269, n25270, n25271,
         n25272, n25273, n25274, n25275, n25276, n25277, n25278, n25279,
         n25280, n25281, n25282, n25283, n25284, n25285, n25286, n25287,
         n25288, n25289, n25290, n25291, n25292, n25293, n25294, n25295,
         n25296, n25297, n25298, n25299, n25300, n25301, n25302, n25303,
         n25304, n25305, n25306, n25307, n25308, n25309, n25310, n25311,
         n25312, n25313, n25314, n25315, n25316, n25317, n25318, n25319,
         n25320, n25321, n25322, n25323, n25324, n25325, n25326, n25327,
         n25328, n25329, n25330, n25331, n25332, n25333, n25334, n25335,
         n25336, n25337, n25338, n25339, n25340, n25341, n25342, n25343,
         n25344, n25345, n25346, n25347, n25348, n25349, n25350, n25351,
         n25352, n25353, n25354, n25355, n25356, n25357, n25358, n25359,
         n25360, n25361, n25362, n25363, n25364, n25365, n25366, n25367,
         n25368, n25369, n25370, n25371, n25372, n25373, n25374, n25375,
         n25376, n25377, n25378, n25379, n25380, n25381, n25382, n25383,
         n25384, n25385, n25386, n25387, n25388, n25389, n25390, n25391,
         n25392, n25393, n25394, n25395, n25396, n25397, n25398, n25399,
         n25400, n25401, n25402, n25403, n25404, n25405, n25406, n25407,
         n25408, n25409, n25410, n25411, n25412, n25413, n25414, n25415,
         n25416, n25417, n25418, n25419, n25420, n25421, n25422, n25423,
         n25424, n25425, n25426, n25427, n25428, n25429, n25430, n25431,
         n25432, n25433, n25434, n25435, n25436, n25437, n25438, n25439,
         n25440, n25441, n25442, n25443, n25444, n25445, n25446, n25447,
         n25448, n25449, n25450, n25451, n25452, n25453, n25454, n25455,
         n25456, n25457, n25458, n25459, n25460, n25461, n25462, n25463,
         n25464, n25465, n25466, n25467, n25468, n25469, n25470, n25471,
         n25472, n25473, n25474, n25475, n25476, n25477, n25478, n25479,
         n25480, n25481, n25482, n25483, n25484, n25485, n25486, n25487,
         n25488, n25489, n25490, n25491, n25492, n25493, n25494, n25495,
         n25496, n25497, n25498, n25499, n25500, n25501, n25502, n25503,
         n25504, n25505, n25506, n25507, n25508, n25509, n25510, n25511,
         n25512, n25513, n25514, n25515, n25516, n25517, n25518, n25519,
         n25520, n25521, n25522, n25523, n25524, n25525, n25526, n25527,
         n25528, n25529, n25530, n25531, n25532, n25533, n25534, n25535,
         n25536, n25537, n25538, n25539, n25540, n25541, n25542, n25543,
         n25544, n25545, n25546, n25547, n25548, n25549, n25550, n25551,
         n25552, n25553, n25554, n25555, n25556, n25557, n25558, n25559,
         n25560, n25561, n25562, n25563, n25564, n25565, n25566, n25567,
         n25568, n25569, n25570, n25571, n25572, n25573, n25574, n25575,
         n25576, n25577, n25578, n25579, n25580, n25581, n25582, n25583,
         n25584, n25585, n25586, n25587, n25588, n25589, n25590, n25591,
         n25592, n25593, n25594, n25595, n25596, n25597, n25598, n25599,
         n25600, n25601, n25602, n25603, n25604, n25605, n25606, n25607,
         n25608, n25609, n25610, n25611, n25612, n25613, n25614, n25615,
         n25616, n25617, n25618, n25619, n25620, n25621, n25622, n25623,
         n25624, n25625, n25626, n25627, n25628, n25629, n25630, n25631,
         n25632, n25633, n25634, n25635, n25636, n25637, n25638, n25639,
         n25640, n25641, n25642, n25643, n25644, n25645, n25646, n25647,
         n25648, n25649, n25650, n25651, n25652, n25653, n25654, n25655,
         n25656, n25657, n25658, n25659, n25660, n25661, n25662, n25663,
         n25664, n25665, n25666, n25667, n25668, n25669, n25670, n25671,
         n25672, n25673, n25674, n25675, n25676, n25677, n25678, n25679,
         n25680, n25681, n25682, n25683, n25684, n25685, n25686, n25687,
         n25688, n25689, n25690, n25691, n25692, n25693, n25694, n25695,
         n25696, n25697, n25698, n25699, n25700, n25701, n25702, n25703,
         n25704, n25705, n25706, n25707, n25708, n25709, n25710, n25711,
         n25712, n25713, n25714, n25715, n25716, n25717, n25718, n25719,
         n25720, n25721, n25722, n25723, n25724, n25725, n25726, n25727,
         n25728, n25729, n25730, n25731, n25732, n25733, n25734, n25735,
         n25736, n25737, n25738, n25739, n25740, n25741, n25742, n25743,
         n25744, n25745, n25746, n25747, n25748, n25749, n25750, n25751,
         n25752, n25753, n25754, n25755, n25756, n25757, n25758, n25759,
         n25760, n25761, n25762, n25763, n25764, n25765, n25766, n25767,
         n25768, n25769, n25770, n25771, n25772, n25773, n25774, n25775,
         n25776, n25777, n25778, n25779, n25780, n25781, n25782, n25783,
         n25784, n25785, n25786, n25787, n25788, n25789, n25790, n25791,
         n25792, n25793, n25794, n25795, n25796, n25797, n25798, n25799,
         n25800, n25801, n25802, n25803, n25804, n25805, n25806, n25807,
         n25808, n25809, n25810, n25811, n25812, n25813, n25814, n25815,
         n25816, n25817, n25818, n25819, n25820, n25821, n25822, n25823,
         n25824, n25825, n25826, n25827, n25828, n25829, n25830, n25831,
         n25832, n25833, n25834, n25835, n25836, n25837, n25838, n25839,
         n25840, n25841, n25842, n25843, n25844, n25845, n25846, n25847,
         n25848, n25849, n25850, n25851, n25852, n25853, n25854, n25855,
         n25856, n25857, n25858, n25859, n25860, n25861, n25862, n25863,
         n25864, n25865, n25866, n25867, n25868, n25869, n25870, n25871,
         n25872, n25873, n25874, n25875, n25876, n25877, n25878, n25879,
         n25880, n25881, n25882, n25883, n25884, n25885, n25886, n25887,
         n25888, n25889, n25890, n25891, n25892, n25893, n25894, n25895,
         n25896, n25897, n25898, n25899, n25900, n25901, n25902, n25903,
         n25904, n25905, n25906, n25907, n25908, n25909, n25910, n25911,
         n25912, n25913, n25914, n25915, n25916, n25917, n25918, n25919,
         n25920, n25921, n25922, n25923, n25924, n25925, n25926, n25927,
         n25928, n25929, n25930, n25931, n25932, n25933, n25934, n25935,
         n25936, n25937, n25938, n25939, n25940, n25941, n25942, n25943,
         n25944, n25945, n25946, n25947, n25948, n25949, n25950, n25951,
         n25952, n25953, n25954, n25955, n25956, n25957, n25958, n25959,
         n25960, n25961, n25962, n25963, n25964, n25965, n25966, n25967,
         n25968, n25969, n25970, n25971, n25972, n25973, n25974, n25975,
         n25976, n25977, n25978, n25979, n25980, n25981, n25982, n25983,
         n25984, n25985, n25986, n25987, n25988, n25989, n25990, n25991,
         n25992, n25993, n25994, n25995, n25996, n25997, n25998, n25999,
         n26000, n26001, n26002, n26003, n26004, n26005, n26006, n26007,
         n26008, n26009, n26010, n26011, n26012, n26013, n26014, n26015,
         n26016, n26017, n26018, n26019, n26020, n26021, n26022, n26023,
         n26024, n26025, n26026, n26027, n26028, n26029, n26030, n26031,
         n26032, n26033, n26034, n26035, n26036, n26037, n26038, n26039,
         n26040, n26041, n26042, n26043, n26044, n26045, n26046, n26047,
         n26048, n26049, n26050, n26051, n26052, n26053, n26054, n26055,
         n26056, n26057, n26058, n26059, n26060, n26061, n26062, n26063,
         n26064, n26065, n26066, n26067, n26068, n26069, n26070, n26071,
         n26072, n26073, n26074, n26075, n26076, n26077, n26078, n26079,
         n26080, n26081, n26082, n26083, n26084, n26085, n26086, n26087,
         n26088, n26089, n26090, n26091, n26092, n26093, n26094, n26095,
         n26096, n26097, n26098, n26099, n26100, n26101, n26102, n26103,
         n26104, n26105, n26106, n26107, n26108, n26109, n26110, n26111,
         n26112, n26113, n26114, n26115, n26116, n26117, n26118, n26119,
         n26120, n26121, n26122, n26123, n26124, n26125, n26126, n26127,
         n26128, n26129, n26130, n26131, n26132, n26133, n26134, n26135,
         n26136, n26137, n26138, n26139, n26140, n26141, n26142, n26143,
         n26144, n26145, n26146, n26147, n26148, n26149, n26150, n26151,
         n26152, n26153, n26154, n26155, n26156, n26157, n26158, n26159,
         n26160, n26161, n26162, n26163, n26164, n26165, n26166, n26167,
         n26168, n26169, n26170, n26171, n26172, n26173, n26174, n26175,
         n26176, n26177, n26178, n26179, n26180, n26181, n26182, n26183,
         n26184, n26185, n26186, n26187, n26188, n26189, n26190, n26191,
         n26192, n26193, n26194, n26195, n26196, n26197, n26198, n26199,
         n26200, n26201, n26202, n26203, n26204, n26205, n26206, n26207,
         n26208, n26209, n26210, n26211, n26212, n26213, n26214, n26215,
         n26216, n26217, n26218, n26219, n26220, n26221, n26222, n26223,
         n26224, n26225, n26226, n26227, n26228, n26229, n26230, n26231,
         n26232, n26233, n26234, n26235, n26236, n26237, n26238, n26239,
         n26240, n26241, n26242, n26243, n26244, n26245, n26246, n26247,
         n26248, n26249, n26250, n26251, n26252, n26253, n26254, n26255,
         n26256, n26257, n26258, n26259, n26260, n26261, n26262, n26263,
         n26264, n26265, n26266, n26267, n26268, n26269, n26270, n26271,
         n26272, n26273, n26274, n26275, n26276, n26277, n26278, n26279,
         n26280, n26281, n26282, n26283, n26284, n26285, n26286, n26287,
         n26288, n26289, n26290, n26291, n26292, n26293, n26294, n26295,
         n26296, n26297, n26298, n26299, n26300, n26301, n26302, n26303,
         n26304, n26305, n26306, n26307, n26308, n26309, n26310, n26311,
         n26312, n26313, n26314, n26315, n26316, n26317, n26318, n26319,
         n26320, n26321, n26322, n26323, n26324, n26325, n26326, n26327,
         n26328, n26329, n26330, n26331, n26332, n26333, n26334, n26335,
         n26336, n26337, n26338, n26339, n26340, n26341, n26342, n26343,
         n26344, n26345, n26346, n26347, n26348, n26349, n26350, n26351,
         n26352, n26353, n26354, n26355, n26356, n26357, n26358, n26359,
         n26360, n26361, n26362, n26363, n26364, n26365, n26366, n26367,
         n26368, n26369, n26370, n26371, n26372, n26373, n26374, n26375,
         n26376, n26377, n26378, n26379, n26380, n26381, n26382, n26383,
         n26384, n26385, n26386, n26387, n26388, n26389, n26390, n26391,
         n26392, n26393, n26394, n26395, n26396, n26397, n26398, n26399,
         n26400, n26401, n26402, n26403, n26404, n26405, n26406, n26407,
         n26408, n26409, n26410, n26411, n26412, n26413, n26414, n26415,
         n26416, n26417, n26418, n26419, n26420, n26421, n26422, n26423,
         n26424, n26425, n26426, n26427, n26428, n26429, n26430, n26431,
         n26432, n26433, n26434, n26435, n26436, n26437, n26438, n26439,
         n26440, n26441, n26442, n26443, n26444, n26445, n26446, n26447,
         n26448, n26449, n26450, n26451, n26452, n26453, n26454, n26455,
         n26456, n26457, n26458, n26459, n26460, n26461, n26462, n26463,
         n26464, n26465, n26466, n26467, n26468, n26469, n26470, n26471,
         n26472, n26473, n26474, n26475, n26476, n26477, n26478, n26479,
         n26480, n26481, n26482, n26483, n26484, n26485, n26486, n26487,
         n26488, n26489, n26490, n26491, n26492, n26493, n26494, n26495,
         n26496, n26497, n26498, n26499, n26500, n26501, n26502, n26503,
         n26504, n26505, n26506, n26507, n26508, n26509, n26510, n26511,
         n26512, n26513, n26514, n26515, n26516, n26517, n26518, n26519,
         n26520, n26521, n26522, n26523, n26524, n26525, n26526, n26527,
         n26528, n26529, n26530, n26531, n26532, n26533, n26534, n26535,
         n26536, n26537, n26538, n26539, n26540, n26541, n26542, n26543,
         n26544, n26545, n26546, n26547, n26548, n26549, n26550, n26551,
         n26552, n26553, n26554, n26555, n26556, n26557, n26558, n26559,
         n26560, n26561, n26562, n26563, n26564, n26565, n26566, n26567,
         n26568, n26569, n26570, n26571, n26572, n26573, n26574, n26575,
         n26576, n26577, n26578, n26579, n26580, n26581, n26582, n26583,
         n26584, n26585, n26586, n26587, n26588, n26589, n26590, n26591,
         n26592, n26593, n26594, n26595, n26596, n26597, n26598, n26599,
         n26600, n26601, n26602, n26603, n26604, n26605, n26606, n26607,
         n26608, n26609, n26610, n26611, n26612, n26613, n26614, n26615,
         n26616, n26617, n26618, n26619, n26620, n26621, n26622, n26623,
         n26624, n26625, n26626, n26627, n26628, n26629, n26630, n26631,
         n26632, n26633, n26634, n26635, n26636, n26637, n26638, n26639,
         n26640, n26641, n26642, n26643, n26644, n26645, n26646, n26647,
         n26648, n26649, n26650, n26651, n26652, n26653, n26654, n26655,
         n26656, n26657, n26658, n26659, n26660, n26661, n26662, n26663,
         n26664, n26665, n26666, n26667, n26668, n26669, n26670, n26671,
         n26672, n26673, n26674, n26675, n26676, n26677, n26678, n26679,
         n26680, n26681, n26682, n26683, n26684, n26685, n26686, n26687,
         n26688, n26689, n26690, n26691, n26692, n26693, n26694, n26695,
         n26696, n26697, n26698, n26699, n26700, n26701, n26702, n26703,
         n26704, n26705, n26706, n26707, n26708, n26709, n26710, n26711,
         n26712, n26713, n26714, n26715, n26716, n26717, n26718, n26719,
         n26720, n26721, n26722, n26723, n26724, n26725, n26726, n26727,
         n26728, n26729, n26730, n26731, n26732, n26733, n26734, n26735,
         n26736, n26737, n26738, n26739, n26740, n26741, n26742, n26743,
         n26744, n26745, n26746, n26747, n26748, n26749, n26750, n26751,
         n26752, n26753, n26754, n26755, n26756, n26757, n26758, n26759,
         n26760, n26761, n26762, n26763, n26764, n26765, n26766, n26767,
         n26768, n26769, n26770, n26771, n26772, n26773, n26774, n26775,
         n26776, n26777, n26778, n26779, n26780, n26781, n26782, n26783,
         n26784, n26785, n26786, n26787, n26788, n26789, n26790, n26791,
         n26792, n26793, n26794, n26795, n26796, n26797, n26798, n26799,
         n26800, n26801, n26802, n26803, n26804, n26805, n26806, n26807,
         n26808, n26809, n26810, n26811, n26812, n26813, n26814, n26815,
         n26816, n26817, n26818, n26819, n26820, n26821, n26822, n26823,
         n26824, n26825, n26826, n26827, n26828, n26829, n26830, n26831,
         n26832, n26833, n26834, n26835, n26836, n26837, n26838, n26839,
         n26840, n26841, n26842, n26843, n26844, n26845, n26846, n26847,
         n26848, n26849, n26850, n26851, n26852, n26853, n26854, n26855,
         n26856, n26857, n26858, n26859, n26860, n26861, n26862, n26863,
         n26864, n26865, n26866, n26867, n26868, n26869, n26870, n26871,
         n26872, n26873, n26874, n26875, n26876, n26877, n26878, n26879,
         n26880, n26881, n26882, n26883, n26884, n26885, n26886, n26887,
         n26888, n26889, n26890, n26891, n26892, n26893, n26894, n26895,
         n26896, n26897, n26898, n26899, n26900, n26901, n26902, n26903,
         n26904, n26905, n26906, n26907, n26908, n26909, n26910, n26911,
         n26912, n26913, n26914, n26915, n26916, n26917, n26918, n26919,
         n26920, n26921, n26922, n26923, n26924, n26925, n26926, n26927,
         n26928, n26929, n26930, n26931, n26932, n26933, n26934, n26935,
         n26936, n26937, n26938, n26939, n26940, n26941, n26942, n26943,
         n26944, n26945, n26946, n26947, n26948, n26949, n26950, n26951,
         n26952, n26953, n26954, n26955, n26956, n26957, n26958, n26959,
         n26960, n26961, n26962, n26963, n26964, n26965, n26966, n26967,
         n26968, n26969, n26970, n26971, n26972, n26973, n26974, n26975,
         n26976, n26977, n26978, n26979, n26980, n26981, n26982, n26983,
         n26984, n26985, n26986, n26987, n26988, n26989, n26990, n26991,
         n26992, n26993, n26994, n26995, n26996, n26997, n26998, n26999,
         n27000, n27001, n27002, n27003, n27004, n27005, n27006, n27007,
         n27008, n27009, n27010, n27011, n27012, n27013, n27014, n27015,
         n27016, n27017, n27018, n27019, n27020, n27021, n27022, n27023,
         n27024, n27025, n27026, n27027, n27028, n27029, n27030, n27031,
         n27032, n27033, n27034, n27035, n27036, n27037, n27038, n27039,
         n27040, n27041, n27042, n27043, n27044, n27045, n27046, n27047,
         n27048, n27049, n27050, n27051, n27052, n27053, n27054, n27055,
         n27056, n27057, n27058, n27059, n27060, n27061, n27062, n27063,
         n27064, n27065, n27066, n27067, n27068, n27069, n27070, n27071,
         n27072, n27073, n27074, n27075, n27076, n27077, n27078, n27079,
         n27080, n27081, n27082, n27083, n27084, n27085, n27086, n27087,
         n27088, n27089, n27090, n27091, n27092, n27093, n27094, n27095,
         n27096, n27097, n27098, n27099, n27100, n27101, n27102, n27103,
         n27104, n27105, n27106, n27107, n27108, n27109, n27110, n27111,
         n27112, n27113, n27114, n27115, n27116, n27117, n27118, n27119,
         n27120, n27121, n27122, n27123, n27124, n27125, n27126, n27127,
         n27128, n27129, n27130, n27131, n27132, n27133, n27134, n27135,
         n27136, n27137, n27138, n27139, n27140, n27141, n27142, n27143,
         n27144, n27145, n27146, n27147, n27148, n27149, n27150, n27151,
         n27152, n27153, n27154, n27155, n27156, n27157, n27158, n27159,
         n27160, n27161, n27162, n27163, n27164, n27165, n27166, n27167,
         n27168, n27169, n27170, n27171, n27172, n27173, n27174, n27175,
         n27176, n27177, n27178, n27179, n27180, n27181, n27182, n27183,
         n27184, n27185, n27186, n27187, n27188, n27189, n27190, n27191,
         n27192, n27193, n27194, n27195, n27196, n27197, n27198, n27199,
         n27200, n27201, n27202, n27203, n27204, n27205, n27206, n27207,
         n27208, n27209, n27210, n27211, n27212, n27213, n27214, n27215,
         n27216, n27217, n27218, n27219, n27220, n27221, n27222, n27223,
         n27224, n27225, n27226, n27227, n27228, n27229, n27230, n27231,
         n27232, n27233, n27234, n27235, n27236, n27237, n27238, n27239,
         n27240, n27241, n27242, n27243, n27244, n27245, n27246, n27247,
         n27248, n27249, n27250, n27251, n27252, n27253, n27254, n27255,
         n27256, n27257, n27258, n27259, n27260, n27261, n27262, n27263,
         n27264, n27265, n27266, n27267, n27268, n27269, n27270, n27271,
         n27272, n27273, n27274, n27275, n27276, n27277, n27278, n27279,
         n27280, n27281, n27282, n27283, n27284, n27285, n27286, n27287,
         n27288, n27289, n27290, n27291, n27292, n27293, n27294, n27295,
         n27296, n27297, n27298, n27299, n27300, n27301, n27302, n27303,
         n27304, n27305, n27306, n27307, n27308, n27309, n27310, n27311,
         n27312, n27313, n27314, n27315, n27316, n27317, n27318, n27319,
         n27320, n27321, n27322, n27323, n27324, n27325, n27326, n27327,
         n27328, n27329, n27330, n27331, n27332, n27333, n27334, n27335,
         n27336, n27337, n27338, n27339, n27340, n27341, n27342, n27343,
         n27344, n27345, n27346, n27347, n27348, n27349, n27350, n27351,
         n27352, n27353, n27354, n27355, n27356, n27357, n27358, n27359,
         n27360, n27361, n27362, n27363, n27364, n27365, n27366, n27367,
         n27368, n27369, n27370, n27371, n27372, n27373, n27374, n27375,
         n27376, n27377, n27378, n27379, n27380, n27381, n27382, n27383,
         n27384, n27385, n27386, n27387, n27388, n27389, n27390, n27391,
         n27392, n27393, n27394, n27395, n27396, n27397, n27398, n27399,
         n27400, n27401, n27402, n27403, n27404, n27405, n27406, n27407,
         n27408, n27409, n27410, n27411, n27412, n27413, n27414, n27415,
         n27416, n27417, n27418, n27419, n27420, n27421, n27422, n27423,
         n27424, n27425, n27426, n27427, n27428, n27429, n27430, n27431,
         n27432, n27433, n27434, n27435, n27436, n27437, n27438, n27439,
         n27440, n27441, n27442, n27443, n27444, n27445, n27446, n27447,
         n27448, n27449, n27450, n27451, n27452, n27453, n27454, n27455,
         n27456, n27457, n27458, n27459, n27460, n27461, n27462, n27463,
         n27464, n27465, n27466, n27467, n27468, n27469, n27470, n27471,
         n27472, n27473, n27474, n27475, n27476, n27477, n27478, n27479,
         n27480, n27481, n27482, n27483, n27484, n27485, n27486, n27487,
         n27488, n27489, n27490, n27491, n27492, n27493, n27494, n27495,
         n27496, n27497, n27498, n27499, n27500, n27501, n27502, n27503,
         n27504, n27505, n27506, n27507, n27508, n27509, n27510, n27511,
         n27512, n27513, n27514, n27515, n27516, n27517, n27518, n27519,
         n27520, n27521, n27522, n27523, n27524, n27525, n27526, n27527,
         n27528, n27529, n27530, n27531, n27532, n27533, n27534, n27535,
         n27536, n27537, n27538, n27539, n27540, n27541, n27542, n27543,
         n27544, n27545, n27546, n27547, n27548, n27549, n27550, n27551,
         n27552, n27553, n27554, n27555, n27556, n27557, n27558, n27559,
         n27560, n27561, n27562, n27563, n27564, n27565, n27566, n27567,
         n27568, n27569, n27570, n27571, n27572, n27573, n27574, n27575,
         n27576, n27577, n27578, n27579, n27580, n27581, n27582, n27583,
         n27584, n27585, n27586, n27587, n27588, n27589, n27590, n27591,
         n27592, n27593, n27594, n27595, n27596, n27597, n27598, n27599,
         n27600, n27601, n27602, n27603, n27604, n27605, n27606, n27607,
         n27608, n27609, n27610, n27611, n27612, n27613, n27614, n27615,
         n27616, n27617, n27618, n27619, n27620, n27621, n27622, n27623,
         n27624, n27625, n27626, n27627, n27628, n27629, n27630, n27631,
         n27632, n27633, n27634, n27635, n27636, n27637, n27638, n27639,
         n27640, n27641, n27642, n27643, n27644, n27645, n27646, n27647,
         n27648, n27649, n27650, n27651, n27652, n27653, n27654, n27655,
         n27656, n27657, n27658, n27659, n27660, n27661, n27662, n27663,
         n27664, n27665, n27666, n27667, n27668, n27669, n27670, n27671,
         n27672, n27673, n27674, n27675, n27676, n27677, n27678, n27679,
         n27680, n27681, n27682, n27683, n27684, n27685, n27686, n27687,
         n27688, n27689, n27690, n27691, n27692, n27693, n27694, n27695,
         n27696, n27697, n27698, n27699, n27700, n27701, n27702, n27703,
         n27704, n27705, n27706, n27707, n27708, n27709, n27710, n27711,
         n27712, n27713, n27714, n27715, n27716, n27717, n27718, n27719,
         n27720, n27721, n27722, n27723, n27724, n27725, n27726, n27727,
         n27728, n27729, n27730, n27731, n27732, n27733, n27734, n27735,
         n27736, n27737, n27738, n27739, n27740, n27741, n27742, n27743,
         n27744, n27745, n27746, n27747, n27748, n27749, n27750, n27751,
         n27752, n27753, n27754, n27755, n27756, n27757, n27758, n27759,
         n27760, n27761, n27762, n27763, n27764, n27765, n27766, n27767,
         n27768, n27769, n27770, n27771, n27772, n27773, n27774, n27775,
         n27776, n27777, n27778, n27779, n27780, n27781, n27782, n27783,
         n27784, n27785, n27786, n27787, n27788, n27789, n27790, n27791,
         n27792, n27793, n27794, n27795, n27796, n27797, n27798, n27799,
         n27800, n27801, n27802, n27803, n27804, n27805, n27806, n27807,
         n27808, n27809, n27810, n27811, n27812, n27813, n27814, n27815,
         n27816, n27817, n27818, n27819, n27820, n27821, n27822, n27823,
         n27824, n27825, n27826, n27827, n27828, n27829, n27830, n27831,
         n27832, n27833, n27834, n27835, n27836, n27837, n27838, n27839,
         n27840, n27841, n27842, n27843, n27844, n27845, n27846, n27847,
         n27848, n27849, n27850, n27851, n27852, n27853, n27854, n27855,
         n27856, n27857, n27858, n27859, n27860, n27861, n27862, n27863,
         n27864, n27865, n27866, n27867, n27868, n27869, n27870, n27871,
         n27872, n27873, n27874, n27875, n27876, n27877, n27878, n27879,
         n27880, n27881, n27882, n27883, n27884, n27885, n27886, n27887,
         n27888, n27889, n27890, n27891, n27892, n27893, n27894, n27895,
         n27896, n27897, n27898, n27899, n27900, n27901, n27902, n27903,
         n27904, n27905, n27906, n27907, n27908, n27909, n27910, n27911,
         n27912, n27913, n27914, n27915, n27916, n27917, n27918, n27919,
         n27920, n27921, n27922, n27923, n27924, n27925, n27926, n27927,
         n27928, n27929, n27930, n27931, n27932, n27933, n27934, n27935,
         n27936, n27937, n27938, n27939, n27940, n27941, n27942, n27943,
         n27944, n27945, n27946, n27947, n27948, n27949, n27950, n27951,
         n27952, n27953, n27954, n27955, n27956, n27957, n27958, n27959,
         n27960, n27961, n27962, n27963, n27964, n27965, n27966, n27967,
         n27968, n27969, n27970, n27971, n27972, n27973, n27974, n27975,
         n27976, n27977, n27978, n27979, n27980, n27981, n27982, n27983,
         n27984, n27985, n27986, n27987, n27988, n27989, n27990, n27991,
         n27992, n27993, n27994, n27995, n27996, n27997, n27998, n27999,
         n28000, n28001, n28002, n28003, n28004, n28005, n28006, n28007,
         n28008, n28009, n28010, n28011, n28012, n28013, n28014, n28015,
         n28016, n28017, n28018, n28019, n28020, n28021, n28022, n28023,
         n28024, n28025, n28026, n28027, n28028, n28029, n28030, n28031,
         n28032, n28033, n28034, n28035, n28036, n28037, n28038, n28039,
         n28040, n28041, n28042, n28043, n28044, n28045, n28046, n28047,
         n28048, n28049, n28050, n28051, n28052, n28053, n28054, n28055,
         n28056, n28057, n28058, n28059, n28060, n28061, n28062, n28063,
         n28064, n28065, n28066, n28067, n28068, n28069, n28070, n28071,
         n28072, n28073, n28074, n28075, n28076, n28077, n28078, n28079,
         n28080, n28081, n28082, n28083, n28084, n28085, n28086, n28087,
         n28088, n28089, n28090, n28091, n28092, n28093, n28094, n28095,
         n28096, n28097, n28098, n28099, n28100, n28101, n28102, n28103,
         n28104, n28105, n28106, n28107, n28108, n28109, n28110, n28111,
         n28112, n28113, n28114, n28115, n28116, n28117, n28118, n28119,
         n28120, n28121, n28122, n28123, n28124, n28125, n28126, n28127,
         n28128, n28129, n28130, n28131, n28132, n28133, n28134, n28135,
         n28136, n28137, n28138, n28139, n28140, n28141, n28142, n28143,
         n28144, n28145, n28146, n28147, n28148, n28149, n28150, n28151,
         n28152, n28153, n28154, n28155, n28156, n28157, n28158, n28159,
         n28160, n28161, n28162, n28163, n28164, n28165, n28166, n28167,
         n28168, n28169, n28170, n28171, n28172, n28173, n28174, n28175,
         n28176, n28177, n28178, n28179, n28180, n28181, n28182, n28183,
         n28184, n28185, n28186, n28187, n28188, n28189, n28190, n28191,
         n28192, n28193, n28194, n28195, n28196, n28197, n28198, n28199,
         n28200, n28201, n28202, n28203, n28204, n28205, n28206, n28207,
         n28208, n28209, n28210, n28211, n28212, n28213, n28214, n28215,
         n28216, n28217, n28218, n28219, n28220, n28221, n28222, n28223,
         n28224, n28225, n28226, n28227, n28228, n28229, n28230, n28231,
         n28232, n28233, n28234, n28235, n28236, n28237, n28238, n28239,
         n28240, n28241, n28242, n28243, n28244, n28245, n28246, n28247,
         n28248, n28249, n28250, n28251, n28252, n28253, n28254, n28255,
         n28256, n28257, n28258, n28259, n28260, n28261, n28262, n28263,
         n28264, n28265, n28266, n28267, n28268, n28269, n28270, n28271,
         n28272, n28273, n28274, n28275, n28276, n28277, n28278, n28279,
         n28280, n28281, n28282, n28283, n28284, n28285, n28286, n28287,
         n28288, n28289, n28290, n28291, n28292, n28293, n28294, n28295,
         n28296, n28297, n28298, n28299, n28300, n28301, n28302, n28303,
         n28304, n28305, n28306, n28307, n28308, n28309, n28310, n28311,
         n28312, n28313, n28314, n28315, n28316, n28317, n28318, n28319,
         n28320, n28321, n28322, n28323, n28324, n28325, n28326, n28327,
         n28328, n28329, n28330, n28331, n28332, n28333, n28334, n28335,
         n28336, n28337, n28338, n28339, n28340, n28341, n28342, n28343,
         n28344, n28345, n28346, n28347, n28348, n28349, n28350, n28351,
         n28352, n28353, n28354, n28355, n28356, n28357, n28358, n28359,
         n28360, n28361, n28362, n28363, n28364, n28365, n28366, n28367,
         n28368, n28369, n28370, n28371, n28372, n28373, n28374, n28375,
         n28376, n28377, n28378, n28379, n28380, n28381, n28382, n28383,
         n28384, n28385, n28386, n28387, n28388, n28389, n28390, n28391,
         n28392, n28393, n28394, n28395, n28396, n28397, n28398, n28399,
         n28400, n28401, n28402, n28403, n28404, n28405, n28406, n28407,
         n28408, n28409, n28410, n28411, n28412, n28413, n28414, n28415,
         n28416, n28417, n28418, n28419, n28420, n28421, n28422, n28423,
         n28424, n28425, n28426, n28427, n28428, n28429, n28430, n28431,
         n28432, n28433, n28434, n28435, n28436, n28437, n28438, n28439,
         n28440, n28441, n28442, n28443, n28444, n28445, n28446, n28447,
         n28448, n28449, n28450, n28451, n28452, n28453, n28454, n28455,
         n28456, n28457, n28458, n28459, n28460, n28461, n28462, n28463,
         n28464, n28465, n28466, n28467, n28468, n28469, n28470, n28471,
         n28472, n28473, n28474, n28475, n28476, n28477, n28478, n28479,
         n28480, n28481, n28482, n28483, n28484, n28485, n28486, n28487,
         n28488, n28489, n28490, n28491, n28492, n28493, n28494, n28495,
         n28496, n28497, n28498, n28499, n28500, n28501, n28502, n28503,
         n28504, n28505, n28506, n28507, n28508, n28509, n28510, n28511,
         n28512, n28513, n28514, n28515, n28516, n28517, n28518, n28519,
         n28520, n28521, n28522, n28523, n28524, n28525, n28526, n28527,
         n28528, n28529, n28530, n28531, n28532, n28533, n28534, n28535,
         n28536, n28537, n28538, n28539, n28540, n28541, n28542, n28543,
         n28544, n28545, n28546, n28547, n28548, n28549, n28550, n28551,
         n28552, n28553, n28554, n28555, n28556, n28557, n28558, n28559,
         n28560, n28561, n28562, n28563, n28564, n28565, n28566, n28567,
         n28568, n28569, n28570, n28571, n28572, n28573, n28574, n28575,
         n28576, n28577, n28578, n28579, n28580, n28581, n28582, n28583,
         n28584, n28585, n28586, n28587, n28588, n28589, n28590, n28591,
         n28592, n28593, n28594, n28595, n28596, n28597, n28598, n28599,
         n28600, n28601, n28602, n28603, n28604, n28605, n28606, n28607,
         n28608, n28609, n28610, n28611, n28612, n28613, n28614, n28615,
         n28616, n28617, n28618, n28619, n28620, n28621, n28622, n28623,
         n28624, n28625, n28626, n28627, n28628, n28629, n28630, n28631,
         n28632, n28633, n28634, n28635, n28636, n28637, n28638, n28639,
         n28640, n28641, n28642, n28643, n28644, n28645, n28646, n28647,
         n28648, n28649, n28650, n28651, n28652, n28653, n28654, n28655,
         n28656, n28657, n28658, n28659, n28660, n28661, n28662, n28663,
         n28664, n28665, n28666, n28667, n28668, n28669, n28670, n28671,
         n28672, n28673, n28674, n28675, n28676, n28677, n28678, n28679,
         n28680, n28681, n28682, n28683, n28684, n28685, n28686, n28687,
         n28688, n28689, n28690, n28691, n28692, n28693, n28694, n28695,
         n28696, n28697, n28698, n28699, n28700, n28701, n28702, n28703,
         n28704, n28705, n28706, n28707, n28708, n28709, n28710, n28711,
         n28712, n28713, n28714, n28715, n28716, n28717, n28718, n28719,
         n28720, n28721, n28722, n28723, n28724, n28725, n28726, n28727,
         n28728, n28729, n28730, n28731, n28732, n28733, n28734, n28735,
         n28736, n28737, n28738, n28739, n28740, n28741, n28742, n28743,
         n28744, n28745, n28746, n28747, n28748, n28749, n28750, n28751,
         n28752, n28753, n28754, n28755, n28756, n28757, n28758, n28759,
         n28760, n28761, n28762, n28763, n28764, n28765, n28766, n28767,
         n28768, n28769, n28770, n28771, n28772, n28773, n28774, n28775,
         n28776, n28777, n28778, n28779, n28780, n28781, n28782, n28783,
         n28784, n28785, n28786, n28787, n28788, n28789, n28790, n28791,
         n28792, n28793, n28794, n28795, n28796, n28797, n28798, n28799,
         n28800, n28801, n28802, n28803, n28804, n28805, n28806, n28807,
         n28808, n28809, n28810, n28811, n28812, n28813, n28814, n28815,
         n28816, n28817, n28818, n28819, n28820, n28821, n28822, n28823,
         n28824, n28825, n28826, n28827, n28828, n28829, n28830, n28831,
         n28832, n28833, n28834, n28835, n28836, n28837, n28838, n28839,
         n28840, n28841, n28842, n28843, n28844, n28845, n28846, n28847,
         n28848, n28849, n28850, n28851, n28852, n28853, n28854, n28855,
         n28856, n28857, n28858, n28859, n28860, n28861, n28862, n28863,
         n28864, n28865, n28866, n28867, n28868, n28869, n28870, n28871,
         n28872, n28873, n28874, n28875, n28876, n28877, n28878, n28879,
         n28880, n28881, n28882, n28883, n28884, n28885, n28886, n28887,
         n28888, n28889, n28890, n28891, n28892, n28893, n28894, n28895,
         n28896, n28897, n28898, n28899, n28900, n28901, n28902, n28903,
         n28904, n28905, n28906, n28907, n28908, n28909, n28910, n28911,
         n28912, n28913, n28914, n28915, n28916, n28917, n28918, n28919,
         n28920, n28921, n28922, n28923, n28924, n28925, n28926, n28927,
         n28928, n28929, n28930, n28931, n28932, n28933, n28934, n28935,
         n28936, n28937, n28938, n28939, n28940, n28941, n28942, n28943,
         n28944, n28945, n28946, n28947, n28948, n28949, n28950, n28951,
         n28952, n28953, n28954, n28955, n28956, n28957, n28958, n28959,
         n28960, n28961, n28962, n28963, n28964, n28965, n28966, n28967,
         n28968, n28969, n28970, n28971, n28972, n28973, n28974, n28975,
         n28976, n28977, n28978, n28979, n28980, n28981, n28982, n28983,
         n28984, n28985, n28986, n28987, n28988, n28989, n28990, n28991,
         n28992, n28993, n28994, n28995, n28996, n28997, n28998, n28999,
         n29000, n29001, n29002, n29003, n29004, n29005, n29006, n29007,
         n29008, n29009, n29010, n29011, n29012, n29013, n29014, n29015,
         n29016, n29017, n29018, n29019, n29020, n29021, n29022, n29023,
         n29024, n29025, n29026, n29027, n29028, n29029, n29030, n29031,
         n29032, n29033, n29034, n29035, n29036, n29037, n29038, n29039,
         n29040, n29041, n29042, n29043, n29044, n29045, n29046, n29047,
         n29048, n29049, n29050, n29051, n29052, n29053, n29054, n29055,
         n29056, n29057, n29058, n29059, n29060, n29061, n29062, n29063,
         n29064, n29065, n29066, n29067, n29068, n29069, n29070, n29071,
         n29072, n29073, n29074, n29075, n29076, n29077, n29078, n29079,
         n29080, n29081, n29082, n29083, n29084, n29085, n29086, n29087,
         n29088, n29089, n29090, n29091, n29092, n29093, n29094, n29095,
         n29096, n29097, n29098, n29099, n29100, n29101, n29102, n29103,
         n29104, n29105, n29106, n29107, n29108, n29109, n29110, n29111,
         n29112, n29113, n29114, n29115, n29116, n29117, n29118, n29119,
         n29120, n29121, n29122, n29123, n29124, n29125, n29126, n29127,
         n29128, n29129, n29130, n29131, n29132, n29133, n29134, n29135,
         n29136, n29137, n29138, n29139, n29140, n29141, n29142, n29143,
         n29144, n29145, n29146, n29147, n29148, n29149, n29150, n29151,
         n29152, n29153, n29154, n29155, n29156, n29157, n29158, n29159,
         n29160, n29161, n29162, n29163, n29164, n29165, n29166, n29167,
         n29168, n29169, n29170, n29171, n29172, n29173, n29174, n29175,
         n29176, n29177, n29178, n29179, n29180, n29181, n29182, n29183,
         n29184, n29185, n29186, n29187, n29188, n29189, n29190, n29191,
         n29192, n29193, n29194, n29195, n29196, n29197, n29198, n29199,
         n29200, n29201, n29202, n29203, n29204, n29205, n29206, n29207,
         n29208, n29209, n29210, n29211, n29212, n29213, n29214, n29215,
         n29216, n29217, n29218, n29219, n29220, n29221, n29222, n29223,
         n29224, n29225, n29226, n29227, n29228, n29229, n29230, n29231,
         n29232, n29233, n29234, n29235, n29236, n29237, n29238, n29239,
         n29240, n29241, n29242, n29243, n29244, n29245, n29246, n29247,
         n29248, n29249, n29250, n29251, n29252, n29253, n29254, n29255,
         n29256, n29257, n29258, n29259, n29260, n29261, n29262, n29263,
         n29264, n29265, n29266, n29267, n29268, n29269, n29270, n29271,
         n29272, n29273, n29274, n29275, n29276, n29277, n29278, n29279,
         n29280, n29281, n29282, n29283, n29284, n29285, n29286, n29287,
         n29288, n29289, n29290, n29291, n29292, n29293, n29294, n29295,
         n29296, n29297, n29298, n29299, n29300, n29301, n29302, n29303,
         n29304, n29305, n29306, n29307, n29308, n29309, n29310, n29311,
         n29312, n29313, n29314, n29315, n29316, n29317, n29318, n29319,
         n29320, n29321, n29322, n29323, n29324, n29325, n29326, n29327,
         n29328, n29329, n29330, n29331, n29332, n29333, n29334, n29335,
         n29336, n29337, n29338, n29339, n29340, n29341, n29342, n29343,
         n29344, n29345, n29346, n29347, n29348, n29349, n29350, n29351,
         n29352, n29353, n29354, n29355, n29356, n29357, n29358, n29359,
         n29360, n29361, n29362, n29363, n29364, n29365, n29366, n29367,
         n29368, n29369, n29370, n29371, n29372, n29373, n29374, n29375,
         n29376, n29377, n29378, n29379, n29380, n29381, n29382, n29383,
         n29384, n29385, n29386, n29387, n29388, n29389, n29390, n29391,
         n29392, n29393, n29394, n29395, n29396, n29397, n29398, n29399,
         n29400, n29401, n29402, n29403, n29404, n29405, n29406, n29407,
         n29408, n29409, n29410, n29411, n29412, n29413, n29414, n29415,
         n29416, n29417, n29418, n29419, n29420, n29421, n29422, n29423,
         n29424, n29425, n29426, n29427, n29428, n29429, n29430, n29431,
         n29432, n29433, n29434, n29435, n29436, n29437, n29438, n29439,
         n29440, n29441, n29442, n29443, n29444, n29445, n29446, n29447,
         n29448, n29449, n29450, n29451, n29452, n29453, n29454, n29455,
         n29456, n29457, n29458, n29459, n29460, n29461, n29462, n29463,
         n29464, n29465, n29466, n29467, n29468, n29469, n29470, n29471,
         n29472, n29473, n29474, n29475, n29476, n29477, n29478, n29479,
         n29480, n29481, n29482, n29483, n29484, n29485, n29486, n29487,
         n29488, n29489, n29490, n29491, n29492, n29493, n29494, n29495,
         n29496, n29497, n29498, n29499, n29500, n29501, n29502, n29503,
         n29504, n29505, n29506, n29507, n29508, n29509, n29510, n29511,
         n29512, n29513, n29514, n29515, n29516, n29517, n29518, n29519,
         n29520, n29521, n29522, n29523, n29524, n29525, n29526, n29527,
         n29528, n29529, n29530, n29531, n29532, n29533, n29534, n29535,
         n29536, n29537, n29538, n29539, n29540, n29541, n29542, n29543,
         n29544, n29545, n29546, n29547, n29548, n29549, n29550, n29551,
         n29552, n29553, n29554, n29555, n29556, n29557, n29558, n29559,
         n29560, n29561, n29562, n29563, n29564, n29565, n29566, n29567,
         n29568, n29569, n29570, n29571, n29572, n29573, n29574, n29575,
         n29576, n29577, n29578, n29579, n29580, n29581, n29582, n29583,
         n29584, n29585, n29586, n29587, n29588, n29589, n29590, n29591,
         n29592, n29593, n29594, n29595, n29596, n29597, n29598, n29599,
         n29600, n29601, n29602, n29603, n29604, n29605, n29606, n29607,
         n29608, n29609, n29610, n29611, n29612, n29613, n29614, n29615,
         n29616, n29617, n29618, n29619, n29620, n29621, n29622, n29623,
         n29624, n29625, n29626, n29627, n29628, n29629, n29630, n29631,
         n29632, n29633, n29634, n29635, n29636, n29637, n29638, n29639,
         n29640, n29641, n29642, n29643, n29644, n29645, n29646, n29647,
         n29648, n29649, n29650, n29651, n29652, n29653, n29654, n29655,
         n29656, n29657, n29658, n29659, n29660, n29661, n29662, n29663,
         n29664, n29665, n29666, n29667, n29668, n29669, n29670, n29671,
         n29672, n29673, n29674, n29675, n29676, n29677, n29678, n29679,
         n29680, n29681, n29682, n29683, n29684, n29685, n29686, n29687,
         n29688, n29689, n29690, n29691, n29692, n29693, n29694, n29695,
         n29696, n29697, n29698, n29699, n29700, n29701, n29702, n29703,
         n29704, n29705, n29706, n29707, n29708, n29709, n29710, n29711,
         n29712, n29713, n29714, n29715, n29716, n29717, n29718, n29719,
         n29720, n29721, n29722, n29723, n29724, n29725, n29726, n29727,
         n29728, n29729, n29730, n29731, n29732, n29733, n29734, n29735,
         n29736, n29737, n29738, n29739, n29740, n29741, n29742, n29743,
         n29744, n29745, n29746, n29747, n29748, n29749, n29750, n29751,
         n29752, n29753, n29754, n29755, n29756, n29757, n29758, n29759,
         n29760, n29761, n29762, n29763, n29764, n29765, n29766, n29767,
         n29768, n29769, n29770, n29771, n29772, n29773, n29774, n29775,
         n29776, n29777, n29778, n29779, n29780, n29781, n29782, n29783,
         n29784, n29785, n29786, n29787, n29788, n29789, n29790, n29791,
         n29792, n29793, n29794, n29795, n29796, n29797, n29798, n29799,
         n29800, n29801, n29802, n29803, n29804, n29805, n29806, n29807,
         n29808, n29809, n29810, n29811, n29812, n29813, n29814, n29815,
         n29816, n29817, n29818, n29819, n29820, n29821, n29822, n29823,
         n29824, n29825, n29826, n29827, n29828, n29829, n29830, n29831,
         n29832, n29833, n29834, n29835, n29836, n29837, n29838, n29839,
         n29840, n29841, n29842, n29843, n29844, n29845, n29846, n29847,
         n29848, n29849, n29850, n29851, n29852, n29853, n29854, n29855,
         n29856, n29857, n29858, n29859, n29860, n29861, n29862, n29863,
         n29864, n29865, n29866, n29867, n29868, n29869, n29870, n29871,
         n29872, n29873, n29874, n29875, n29876, n29877, n29878, n29879,
         n29880, n29881, n29882, n29883, n29884, n29885, n29886, n29887,
         n29888, n29889, n29890, n29891, n29892, n29893, n29894, n29895,
         n29896, n29897, n29898, n29899, n29900, n29901, n29902, n29903,
         n29904, n29905, n29906, n29907, n29908, n29909, n29910, n29911,
         n29912, n29913, n29914, n29915, n29916, n29917, n29918, n29919,
         n29920, n29921, n29922, n29923, n29924, n29925, n29926, n29927,
         n29928, n29929, n29930, n29931, n29932, n29933, n29934, n29935,
         n29936, n29937, n29938, n29939, n29940, n29941, n29942, n29943,
         n29944, n29945, n29946, n29947, n29948, n29949, n29950, n29951,
         n29952, n29953, n29954, n29955, n29956, n29957, n29958, n29959,
         n29960, n29961, n29962, n29963, n29964, n29965, n29966, n29967,
         n29968, n29969, n29970, n29971, n29972, n29973, n29974, n29975,
         n29976, n29977, n29978, n29979, n29980, n29981, n29982, n29983,
         n29984, n29985, n29986, n29987, n29988, n29989, n29990, n29991,
         n29992, n29993, n29994, n29995, n29996, n29997, n29998, n29999,
         n30000, n30001, n30002, n30003, n30004, n30005, n30006, n30007,
         n30008, n30009, n30010, n30011, n30012, n30013, n30014, n30015,
         n30016, n30017, n30018, n30019, n30020, n30021, n30022, n30023,
         n30024, n30025, n30026, n30027, n30028, n30029, n30030, n30031,
         n30032, n30033, n30034, n30035, n30036, n30037, n30038, n30039,
         n30040, n30041, n30042, n30043, n30044, n30045, n30046, n30047,
         n30048, n30049, n30050, n30051, n30052, n30053, n30054, n30055,
         n30056, n30057, n30058, n30059, n30060, n30061, n30062, n30063,
         n30064, n30065, n30066, n30067, n30068, n30069, n30070, n30071,
         n30072, n30073, n30074, n30075, n30076, n30077, n30078, n30079,
         n30080, n30081, n30082, n30083, n30084, n30085, n30086, n30087,
         n30088, n30089, n30090, n30091, n30092, n30093, n30094, n30095,
         n30096, n30097, n30098, n30099, n30100, n30101, n30102, n30103,
         n30104, n30105, n30106, n30107, n30108, n30109, n30110, n30111,
         n30112, n30113, n30114, n30115, n30116, n30117, n30118, n30119,
         n30120, n30121, n30122, n30123, n30124, n30125, n30126, n30127,
         n30128, n30129, n30130, n30131, n30132, n30133, n30134, n30135,
         n30136, n30137, n30138, n30139, n30140, n30141, n30142, n30143,
         n30144, n30145, n30146, n30147, n30148, n30149, n30150, n30151,
         n30152, n30153, n30154, n30155, n30156, n30157, n30158, n30159,
         n30160, n30161, n30162, n30163, n30164, n30165, n30166, n30167,
         n30168, n30169, n30170, n30171, n30172, n30173, n30174, n30175,
         n30176, n30177, n30178, n30179, n30180, n30181, n30182, n30183,
         n30184, n30185, n30186, n30187, n30188, n30189, n30190, n30191,
         n30192, n30193, n30194, n30195, n30196, n30197, n30198, n30199,
         n30200, n30201, n30202, n30203, n30204, n30205, n30206, n30207,
         n30208, n30209, n30210, n30211, n30212, n30213, n30214, n30215,
         n30216, n30217, n30218, n30219, n30220, n30221, n30222, n30223,
         n30224, n30225, n30226, n30227, n30228, n30229, n30230, n30231,
         n30232, n30233, n30234, n30235, n30236, n30237, n30238, n30239,
         n30240, n30241, n30242, n30243, n30244, n30245, n30246, n30247,
         n30248, n30249, n30250, n30251, n30252, n30253, n30254, n30255,
         n30256, n30257, n30258, n30259, n30260, n30261, n30262, n30263,
         n30264, n30265, n30266, n30267, n30268, n30269, n30270, n30271,
         n30272, n30273, n30274, n30275, n30276, n30277, n30278, n30279,
         n30280, n30281, n30282, n30283, n30284, n30285, n30286, n30287,
         n30288, n30289, n30290, n30291, n30292, n30293, n30294, n30295,
         n30296, n30297, n30298, n30299, n30300, n30301, n30302, n30303,
         n30304, n30305, n30306, n30307, n30308, n30309, n30310, n30311,
         n30312, n30313, n30314, n30315, n30316, n30317, n30318, n30319,
         n30320, n30321, n30322, n30323, n30324, n30325, n30326, n30327,
         n30328, n30329, n30330, n30331, n30332, n30333, n30334, n30335,
         n30336, n30337, n30338, n30339, n30340, n30341, n30342, n30343,
         n30344, n30345, n30346, n30347, n30348, n30349, n30350, n30351,
         n30352, n30353, n30354, n30355, n30356, n30357, n30358, n30359,
         n30360, n30361, n30362, n30363, n30364, n30365, n30366, n30367,
         n30368, n30369, n30370, n30371, n30372, n30373, n30374, n30375,
         n30376, n30377, n30378, n30379, n30380, n30381, n30382, n30383,
         n30384, n30385, n30386, n30387, n30388, n30389, n30390, n30391,
         n30392, n30393, n30394, n30395, n30396, n30397, n30398, n30399,
         n30400, n30401, n30402, n30403, n30404, n30405, n30406, n30407,
         n30408, n30409, n30410, n30411, n30412, n30413, n30414, n30415,
         n30416, n30417, n30418, n30419, n30420, n30421, n30422, n30423,
         n30424, n30425, n30426, n30427, n30428, n30429, n30430, n30431,
         n30432, n30433, n30434, n30435, n30436, n30437, n30438, n30439,
         n30440, n30441, n30442, n30443, n30444, n30445, n30446, n30447,
         n30448, n30449, n30450, n30451, n30452, n30453, n30454, n30455,
         n30456, n30457, n30458, n30459, n30460, n30461, n30462, n30463,
         n30464, n30465, n30466, n30467, n30468, n30469, n30470, n30471,
         n30472, n30473, n30474, n30475, n30476, n30477, n30478, n30479,
         n30480, n30481, n30482, n30483, n30484, n30485, n30486, n30487,
         n30488, n30489, n30490, n30491, n30492, n30493, n30494, n30495,
         n30496, n30497, n30498, n30499, n30500, n30501, n30502, n30503,
         n30504, n30505, n30506, n30507, n30508, n30509, n30510, n30511,
         n30512, n30513, n30514, n30515, n30516, n30517, n30518, n30519,
         n30520, n30521, n30522, n30523, n30524, n30525, n30526, n30527,
         n30528, n30529, n30530, n30531, n30532, n30533, n30534, n30535,
         n30536, n30537, n30538, n30539, n30540, n30541, n30542, n30543,
         n30544, n30545, n30546, n30547, n30548, n30549, n30550, n30551,
         n30552, n30553, n30554, n30555, n30556, n30557, n30558, n30559,
         n30560, n30561, n30562, n30563, n30564, n30565, n30566, n30567,
         n30568, n30569, n30570, n30571, n30572, n30573, n30574, n30575,
         n30576, n30577, n30578, n30579, n30580, n30581, n30582, n30583,
         n30584, n30585, n30586, n30587, n30588, n30589, n30590, n30591,
         n30592, n30593, n30594, n30595, n30596, n30597, n30598, n30599,
         n30600, n30601, n30602, n30603, n30604, n30605, n30606, n30607,
         n30608, n30609, n30610, n30611, n30612, n30613, n30614, n30615,
         n30616, n30617, n30618, n30619, n30620, n30621, n30622, n30623,
         n30624, n30625, n30626, n30627, n30628, n30629, n30630, n30631,
         n30632, n30633, n30634, n30635, n30636, n30637, n30638, n30639,
         n30640, n30641, n30642, n30643, n30644, n30645, n30646, n30647,
         n30648, n30649, n30650, n30651, n30652, n30653, n30654, n30655,
         n30656, n30657, n30658, n30659, n30660, n30661, n30662, n30663,
         n30664, n30665, n30666, n30667, n30668, n30669, n30670, n30671,
         n30672, n30673, n30674, n30675, n30676, n30677, n30678, n30679,
         n30680, n30681, n30682, n30683, n30684, n30685, n30686, n30687,
         n30688, n30689, n30690, n30691, n30692, n30693, n30694, n30695,
         n30696, n30697, n30698, n30699, n30700, n30701, n30702, n30703,
         n30704, n30705, n30706, n30707, n30708, n30709, n30710, n30711,
         n30712, n30713, n30714, n30715, n30716, n30717, n30718, n30719,
         n30720, n30721, n30722, n30723, n30724, n30725, n30726, n30727,
         n30728, n30729, n30730, n30731, n30732, n30733, n30734, n30735,
         n30736, n30737, n30738, n30739, n30740, n30741, n30742, n30743,
         n30744, n30745, n30746, n30747, n30748, n30749, n30750, n30751,
         n30752, n30753, n30754, n30755, n30756, n30757, n30758, n30759,
         n30760, n30761, n30762, n30763, n30764, n30765, n30766, n30767,
         n30768, n30769, n30770, n30771, n30772, n30773, n30774, n30775,
         n30776, n30777, n30778, n30779, n30780, n30781, n30782, n30783,
         n30784, n30785, n30786, n30787, n30788, n30789, n30790, n30791,
         n30792, n30793, n30794, n30795, n30796, n30797, n30798, n30799,
         n30800, n30801, n30802, n30803, n30804, n30805, n30806, n30807,
         n30808, n30809, n30810, n30811, n30812, n30813, n30814, n30815,
         n30816, n30817, n30818, n30819, n30820, n30821, n30822, n30823,
         n30824, n30825, n30826, n30827, n30828, n30829, n30830, n30831,
         n30832, n30833, n30834, n30835, n30836, n30837, n30838, n30839,
         n30840, n30841, n30842, n30843, n30844, n30845, n30846, n30847,
         n30848, n30849, n30850, n30851, n30852, n30853, n30854, n30855,
         n30856, n30857, n30858, n30859, n30860, n30861, n30862, n30863,
         n30864, n30865, n30866, n30867, n30868, n30869, n30870, n30871,
         n30872, n30873, n30874, n30875, n30876, n30877, n30878, n30879,
         n30880, n30881, n30882, n30883, n30884, n30885, n30886, n30887,
         n30888, n30889, n30890, n30891, n30892, n30893, n30894, n30895,
         n30896, n30897, n30898, n30899, n30900, n30901, n30902, n30903,
         n30904, n30905, n30906, n30907, n30908, n30909, n30910, n30911,
         n30912, n30913, n30914, n30915, n30916, n30917, n30918, n30919,
         n30920, n30921, n30922, n30923, n30924, n30925, n30926, n30927,
         n30928, n30929, n30930, n30931, n30932, n30933, n30934, n30935,
         n30936, n30937, n30938, n30939, n30940, n30941, n30942, n30943,
         n30944, n30945, n30946, n30947, n30948, n30949, n30950, n30951,
         n30952, n30953, n30954, n30955, n30956, n30957, n30958, n30959,
         n30960, n30961, n30962, n30963, n30964, n30965, n30966, n30967,
         n30968, n30969, n30970, n30971, n30972, n30973, n30974, n30975,
         n30976, n30977, n30978, n30979, n30980, n30981, n30982, n30983,
         n30984, n30985, n30986, n30987, n30988, n30989, n30990, n30991,
         n30992, n30993, n30994, n30995, n30996, n30997, n30998, n30999,
         n31000, n31001, n31002, n31003, n31004, n31005, n31006, n31007,
         n31008, n31009, n31010, n31011, n31012, n31013, n31014, n31015,
         n31016, n31017, n31018, n31019, n31020, n31021, n31022, n31023,
         n31024, n31025, n31026, n31027, n31028, n31029, n31030, n31031,
         n31032, n31033, n31034, n31035, n31036, n31037, n31038, n31039,
         n31040, n31041, n31042, n31043, n31044, n31045, n31046, n31047,
         n31048, n31049, n31050, n31051, n31052, n31053, n31054, n31055,
         n31056, n31057, n31058, n31059, n31060, n31061, n31062, n31063,
         n31064, n31065, n31066, n31067, n31068, n31069, n31070, n31071,
         n31072, n31073, n31074, n31075, n31076, n31077, n31078, n31079,
         n31080, n31081, n31082, n31083, n31084, n31085, n31086, n31087,
         n31088, n31089, n31090, n31091, n31092, n31093, n31094, n31095,
         n31096, n31097, n31098, n31099, n31100, n31101, n31102, n31103,
         n31104, n31105, n31106, n31107, n31108, n31109, n31110, n31111,
         n31112, n31113, n31114, n31115, n31116, n31117, n31118, n31119,
         n31120, n31121, n31122, n31123, n31124, n31125, n31126, n31127,
         n31128, n31129, n31130, n31131, n31132, n31133, n31134, n31135,
         n31136, n31137, n31138, n31139, n31140, n31141, n31142, n31143,
         n31144, n31145, n31146, n31147, n31148, n31149, n31150, n31151,
         n31152, n31153, n31154, n31155, n31156, n31157, n31158, n31159,
         n31160, n31161, n31162, n31163, n31164, n31165, n31166, n31167,
         n31168, n31169, n31170, n31171, n31172, n31173, n31174, n31175,
         n31176, n31177, n31178, n31179, n31180, n31181, n31182, n31183,
         n31184, n31185, n31186, n31187, n31188, n31189, n31190, n31191,
         n31192, n31193, n31194, n31195, n31196, n31197, n31198, n31199,
         n31200, n31201, n31202, n31203, n31204, n31205, n31206, n31207,
         n31208, n31209, n31210, n31211, n31212, n31213, n31214, n31215,
         n31216, n31217, n31218, n31219, n31220, n31221, n31222, n31223,
         n31224, n31225, n31226, n31227, n31228, n31229, n31230, n31231,
         n31232, n31233, n31234, n31235, n31236, n31237, n31238, n31239,
         n31240, n31241, n31242, n31243, n31244, n31245, n31246, n31247,
         n31248, n31249, n31250, n31251, n31252, n31253, n31254, n31255,
         n31256, n31257, n31258, n31259, n31260, n31261, n31262, n31263,
         n31264, n31265, n31266, n31267, n31268, n31269, n31270, n31271,
         n31272, n31273, n31274, n31275, n31276, n31277, n31278, n31279,
         n31280, n31281, n31282, n31283, n31284, n31285, n31286, n31287,
         n31288, n31289, n31290, n31291, n31292, n31293, n31294, n31295,
         n31296, n31297, n31298, n31299, n31300, n31301, n31302, n31303,
         n31304, n31305, n31306, n31307, n31308, n31309, n31310, n31311,
         n31312, n31313, n31314, n31315, n31316, n31317, n31318, n31319,
         n31320, n31321, n31322, n31323, n31324, n31325, n31326, n31327,
         n31328, n31329, n31330, n31331, n31332, n31333, n31334, n31335,
         n31336, n31337, n31338, n31339, n31340, n31341, n31342, n31343,
         n31344, n31345, n31346, n31347, n31348, n31349, n31350, n31351,
         n31352, n31353, n31354, n31355, n31356, n31357, n31358, n31359,
         n31360, n31361, n31362, n31363, n31364, n31365, n31366, n31367,
         n31368, n31369, n31370, n31371, n31372, n31373, n31374, n31375,
         n31376, n31377, n31378, n31379, n31380, n31381, n31382, n31383,
         n31384, n31385, n31386, n31387, n31388, n31389, n31390, n31391,
         n31392, n31393, n31394, n31395, n31396, n31397, n31398, n31399,
         n31400, n31401, n31402, n31403, n31404, n31405, n31406, n31407,
         n31408, n31409, n31410, n31411, n31412, n31413, n31414, n31415,
         n31416, n31417, n31418, n31419, n31420, n31421, n31422, n31423,
         n31424, n31425, n31426, n31427, n31428, n31429, n31430, n31431,
         n31432, n31433, n31434, n31435, n31436, n31437, n31438, n31439,
         n31440, n31441, n31442, n31443, n31444, n31445, n31446, n31447,
         n31448, n31449, n31450, n31451, n31452, n31453, n31454, n31455,
         n31456, n31457, n31458, n31459, n31460, n31461, n31462, n31463,
         n31464, n31465, n31466, n31467, n31468, n31469, n31470, n31471,
         n31472, n31473, n31474, n31475, n31476, n31477, n31478, n31479,
         n31480, n31481, n31482, n31483, n31484, n31485, n31486, n31487,
         n31488, n31489, n31490, n31491, n31492, n31493, n31494, n31495,
         n31496, n31497, n31498, n31499, n31500, n31501, n31502, n31503,
         n31504, n31505, n31506, n31507, n31508, n31509, n31510, n31511,
         n31512, n31513, n31514, n31515, n31516, n31517, n31518, n31519,
         n31520, n31521, n31522, n31523, n31524, n31525, n31526, n31527,
         n31528, n31529, n31530, n31531, n31532, n31533, n31534, n31535,
         n31536, n31537, n31538, n31539, n31540, n31541, n31542, n31543,
         n31544, n31545, n31546, n31547, n31548, n31549, n31550, n31551,
         n31552, n31553, n31554, n31555, n31556, n31557, n31558, n31559,
         n31560, n31561, n31562, n31563, n31564, n31565, n31566, n31567,
         n31568, n31569, n31570, n31571, n31572, n31573, n31574, n31575,
         n31576, n31577, n31578, n31579, n31580, n31581, n31582, n31583,
         n31584, n31585, n31586, n31587, n31588, n31589, n31590, n31591,
         n31592, n31593, n31594, n31595, n31596, n31597, n31598, n31599,
         n31600, n31601, n31602, n31603, n31604, n31605, n31606, n31607,
         n31608, n31609, n31610, n31611, n31612, n31613, n31614, n31615,
         n31616, n31617, n31618, n31619, n31620, n31621, n31622, n31623,
         n31624, n31625, n31626, n31627, n31628, n31629, n31630, n31631,
         n31632, n31633, n31634, n31635, n31636, n31637, n31638, n31639,
         n31640, n31641, n31642, n31643, n31644, n31645, n31646, n31647,
         n31648, n31649, n31650, n31651, n31652, n31653, n31654, n31655,
         n31656, n31657, n31658, n31659, n31660, n31661, n31662, n31663,
         n31664, n31665, n31666, n31667, n31668, n31669, n31670, n31671,
         n31672, n31673, n31674, n31675, n31676, n31677, n31678, n31679,
         n31680, n31681, n31682, n31683, n31684, n31685, n31686, n31687,
         n31688, n31689, n31690, n31691, n31692, n31693, n31694, n31695,
         n31696, n31697, n31698, n31699, n31700, n31701, n31702, n31703,
         n31704, n31705, n31706, n31707, n31708, n31709, n31710, n31711,
         n31712, n31713, n31714, n31715, n31716, n31717, n31718, n31719,
         n31720, n31721, n31722, n31723, n31724, n31725, n31726, n31727,
         n31728, n31729, n31730, n31731, n31732, n31733, n31734, n31735,
         n31736, n31737, n31738, n31739, n31740, n31741, n31742, n31743,
         n31744, n31745, n31746, n31747, n31748, n31749, n31750, n31751,
         n31752, n31753, n31754, n31755, n31756, n31757, n31758, n31759,
         n31760, n31761, n31762, n31763, n31764, n31765, n31766, n31767,
         n31768, n31769, n31770, n31771, n31772, n31773, n31774, n31775,
         n31776, n31777, n31778, n31779, n31780, n31781, n31782, n31783,
         n31784, n31785, n31786, n31787, n31788, n31789, n31790, n31791,
         n31792, n31793, n31794, n31795, n31796, n31797, n31798, n31799,
         n31800, n31801, n31802, n31803, n31804, n31805, n31806, n31807,
         n31808, n31809, n31810, n31811, n31812, n31813, n31814, n31815,
         n31816, n31817, n31818, n31819, n31820, n31821, n31822, n31823,
         n31824, n31825, n31826, n31827, n31828, n31829, n31830, n31831,
         n31832, n31833, n31834, n31835, n31836, n31837, n31838, n31839,
         n31840, n31841, n31842, n31843, n31844, n31845, n31846, n31847,
         n31848, n31849, n31850, n31851, n31852, n31853, n31854, n31855,
         n31856, n31857, n31858, n31859, n31860, n31861, n31862, n31863,
         n31864, n31865, n31866, n31867, n31868, n31869, n31870, n31871,
         n31872, n31873, n31874, n31875, n31876, n31877, n31878, n31879,
         n31880, n31881, n31882, n31883, n31884, n31885, n31886, n31887,
         n31888, n31889, n31890, n31891, n31892, n31893, n31894, n31895,
         n31896, n31897, n31898, n31899, n31900, n31901, n31902, n31903,
         n31904, n31905, n31906, n31907, n31908, n31909, n31910, n31911,
         n31912, n31913, n31914, n31915, n31916, n31917, n31918, n31919,
         n31920, n31921, n31922, n31923, n31924, n31925, n31926, n31927,
         n31928, n31929, n31930, n31931, n31932, n31933, n31934, n31935,
         n31936, n31937, n31938, n31939, n31940, n31941, n31942, n31943,
         n31944, n31945, n31946, n31947, n31948, n31949, n31950, n31951,
         n31952, n31953, n31954, n31955, n31956, n31957, n31958, n31959,
         n31960, n31961, n31962, n31963, n31964, n31965, n31966, n31967,
         n31968, n31969, n31970, n31971, n31972, n31973, n31974, n31975,
         n31976, n31977, n31978, n31979, n31980, n31981, n31982, n31983,
         n31984, n31985, n31986, n31987, n31988, n31989, n31990, n31991,
         n31992, n31993, n31994, n31995, n31996, n31997, n31998, n31999,
         n32000, n32001, n32002, n32003, n32004, n32005, n32006, n32007,
         n32008, n32009, n32010, n32011, n32012, n32013, n32014, n32015,
         n32016, n32017, n32018, n32019, n32020, n32021, n32022, n32023,
         n32024, n32025, n32026, n32027, n32028, n32029, n32030, n32031,
         n32032, n32033, n32034, n32035, n32036, n32037, n32038, n32039,
         n32040, n32041, n32042, n32043, n32044, n32045, n32046, n32047,
         n32048, n32049, n32050, n32051, n32052, n32053, n32054, n32055,
         n32056, n32057, n32058, n32059, n32060, n32061, n32062, n32063,
         n32064, n32065, n32066, n32067, n32068, n32069, n32070, n32071,
         n32072, n32073, n32074, n32075, n32076, n32077, n32078, n32079,
         n32080, n32081, n32082, n32083, n32084, n32085, n32086, n32087,
         n32088, n32089, n32090, n32091, n32092, n32093, n32094, n32095,
         n32096, n32097, n32098, n32099, n32100, n32101, n32102, n32103,
         n32104, n32105, n32106, n32107, n32108, n32109, n32110, n32111,
         n32112, n32113, n32114, n32115, n32116, n32117, n32118, n32119,
         n32120, n32121, n32122, n32123, n32124, n32125, n32126, n32127,
         n32128, n32129, n32130, n32131, n32132, n32133, n32134, n32135,
         n32136, n32137, n32138, n32139, n32140, n32141, n32142, n32143,
         n32144, n32145, n32146, n32147, n32148, n32149, n32150, n32151,
         n32152, n32153, n32154, n32155, n32156, n32157, n32158, n32159,
         n32160, n32161, n32162, n32163, n32164, n32165, n32166, n32167,
         n32168, n32169, n32170, n32171, n32172, n32173, n32174, n32175,
         n32176, n32177, n32178, n32179, n32180, n32181, n32182, n32183,
         n32184, n32185, n32186, n32187, n32188, n32189, n32190, n32191,
         n32192, n32193, n32194, n32195, n32196, n32197, n32198, n32199,
         n32200, n32201, n32202, n32203, n32204, n32205, n32206, n32207,
         n32208, n32209, n32210, n32211, n32212, n32213, n32214, n32215,
         n32216, n32217, n32218, n32219, n32220, n32221, n32222, n32223,
         n32224, n32225, n32226, n32227, n32228, n32229, n32230, n32231,
         n32232, n32233, n32234, n32235, n32236, n32237, n32238, n32239,
         n32240, n32241, n32242, n32243, n32244, n32245, n32246, n32247,
         n32248, n32249, n32250, n32251, n32252, n32253, n32254, n32255,
         n32256, n32257, n32258, n32259, n32260, n32261, n32262, n32263,
         n32264, n32265, n32266, n32267, n32268, n32269, n32270, n32271,
         n32272, n32273, n32274, n32275, n32276, n32277, n32278, n32279,
         n32280, n32281, n32282, n32283, n32284, n32285, n32286, n32287,
         n32288, n32289, n32290, n32291, n32292, n32293, n32294, n32295,
         n32296, n32297, n32298, n32299, n32300, n32301, n32302, n32303,
         n32304, n32305, n32306, n32307, n32308, n32309, n32310, n32311,
         n32312, n32313, n32314, n32315, n32316, n32317, n32318, n32319,
         n32320, n32321, n32322, n32323, n32324, n32325, n32326, n32327,
         n32328, n32329, n32330, n32331, n32332, n32333, n32334, n32335,
         n32336, n32337, n32338, n32339, n32340, n32341, n32342, n32343,
         n32344, n32345, n32346, n32347, n32348, n32349, n32350, n32351,
         n32352, n32353, n32354, n32355, n32356, n32357, n32358, n32359,
         n32360, n32361, n32362, n32363, n32364, n32365, n32366, n32367,
         n32368, n32369, n32370, n32371, n32372, n32373, n32374, n32375,
         n32376, n32377, n32378, n32379, n32380, n32381, n32382, n32383,
         n32384, n32385, n32386, n32387, n32388, n32389, n32390, n32391,
         n32392, n32393, n32394, n32395, n32396, n32397, n32398, n32399,
         n32400, n32401, n32402, n32403, n32404, n32405, n32406, n32407,
         n32408, n32409, n32410, n32411, n32412, n32413, n32414, n32415,
         n32416, n32417, n32418, n32419, n32420, n32421, n32422, n32423,
         n32424, n32425, n32426, n32427, n32428, n32429, n32430, n32431,
         n32432, n32433, n32434, n32435, n32436, n32437, n32438, n32439,
         n32440, n32441, n32442, n32443, n32444, n32445, n32446, n32447,
         n32448, n32449, n32450, n32451, n32452, n32453, n32454, n32455,
         n32456, n32457, n32458, n32459, n32460, n32461, n32462, n32463,
         n32464, n32465, n32466, n32467, n32468, n32469, n32470, n32471,
         n32472, n32473, n32474, n32475, n32476, n32477, n32478, n32479,
         n32480, n32481, n32482, n32483, n32484, n32485, n32486, n32487,
         n32488, n32489, n32490, n32491, n32492, n32493, n32494, n32495,
         n32496, n32497, n32498, n32499, n32500, n32501, n32502, n32503,
         n32504, n32505, n32506, n32507, n32508, n32509, n32510, n32511,
         n32512, n32513, n32514, n32515, n32516, n32517, n32518, n32519,
         n32520, n32521, n32522, n32523, n32524, n32525, n32526, n32527,
         n32528, n32529, n32530, n32531, n32532, n32533, n32534, n32535,
         n32536, n32537, n32538, n32539, n32540, n32541, n32542, n32543,
         n32544, n32545, n32546, n32547, n32548, n32549, n32550, n32551,
         n32552, n32553, n32554, n32555, n32556, n32557, n32558, n32559,
         n32560, n32561, n32562, n32563, n32564, n32565, n32566, n32567,
         n32568, n32569, n32570, n32571, n32572, n32573, n32574, n32575,
         n32576, n32577, n32578, n32579, n32580, n32581, n32582, n32583,
         n32584, n32585, n32586, n32587, n32588, n32589, n32590, n32591,
         n32592, n32593, n32594, n32595, n32596, n32597, n32598, n32599,
         n32600, n32601, n32602, n32603, n32604, n32605, n32606, n32607,
         n32608, n32609, n32610, n32611, n32612, n32613, n32614, n32615,
         n32616, n32617, n32618, n32619, n32620, n32621, n32622, n32623,
         n32624, n32625, n32626, n32627, n32628, n32629, n32630, n32631,
         n32632, n32633, n32634, n32635, n32636, n32637, n32638, n32639,
         n32640, n32641, n32642, n32643, n32644, n32645, n32646, n32647,
         n32648, n32649, n32650, n32651, n32652, n32653, n32654, n32655,
         n32656, n32657, n32658, n32659, n32660, n32661, n32662, n32663,
         n32664, n32665, n32666, n32667, n32668, n32669, n32670, n32671,
         n32672, n32673, n32674, n32675, n32676, n32677, n32678, n32679,
         n32680, n32681, n32682, n32683, n32684, n32685, n32686, n32687,
         n32688, n32689, n32690, n32691, n32692, n32693, n32694, n32695,
         n32696, n32697, n32698, n32699, n32700, n32701, n32702, n32703,
         n32704, n32705, n32706, n32707, n32708, n32709, n32710, n32711,
         n32712, n32713, n32714, n32715, n32716, n32717, n32718, n32719,
         n32720, n32721, n32722, n32723, n32724, n32725, n32726, n32727,
         n32728, n32729, n32730, n32731, n32732, n32733, n32734, n32735,
         n32736, n32737, n32738, n32739, n32740, n32741, n32742, n32743,
         n32744, n32745, n32746, n32747, n32748, n32749, n32750, n32751,
         n32752, n32753, n32754, n32755, n32756, n32757, n32758, n32759,
         n32760, n32761, n32762, n32763, n32764, n32765, n32766, n32767,
         n32768, n32769, n32770, n32771, n32772, n32773, n32774, n32775,
         n32776, n32777, n32778, n32779, n32780, n32781, n32782, n32783,
         n32784, n32785, n32786, n32787, n32788, n32789, n32790, n32791,
         n32792, n32793, n32794, n32795, n32796, n32797, n32798, n32799,
         n32800, n32801, n32802, n32803, n32804, n32805, n32806, n32807,
         n32808, n32809, n32810, n32811, n32812, n32813, n32814, n32815,
         n32816, n32817, n32818, n32819, n32820, n32821, n32822, n32823,
         n32824, n32825, n32826, n32827, n32828, n32829, n32830, n32831,
         n32832, n32833, n32834, n32835, n32836, n32837, n32838, n32839,
         n32840, n32841, n32842, n32843, n32844, n32845, n32846, n32847,
         n32848, n32849, n32850, n32851, n32852, n32853, n32854, n32855,
         n32856, n32857, n32858, n32859, n32860, n32861, n32862, n32863,
         n32864, n32865, n32866, n32867, n32868, n32869, n32870, n32871,
         n32872, n32873, n32874, n32875, n32876, n32877, n32878, n32879,
         n32880, n32881, n32882, n32883, n32884, n32885, n32886, n32887,
         n32888, n32889, n32890, n32891, n32892, n32893, n32894, n32895,
         n32896, n32897, n32898, n32899, n32900, n32901, n32902, n32903,
         n32904, n32905, n32906, n32907, n32908, n32909, n32910, n32911,
         n32912, n32913, n32914, n32915, n32916, n32917, n32918, n32919,
         n32920, n32921, n32922, n32923, n32924, n32925, n32926, n32927,
         n32928, n32929, n32930, n32931, n32932, n32933, n32934, n32935,
         n32936, n32937, n32938, n32939, n32940, n32941, n32942, n32943,
         n32944, n32945, n32946, n32947, n32948, n32949, n32950, n32951,
         n32952, n32953, n32954, n32955, n32956, n32957, n32958, n32959,
         n32960, n32961, n32962, n32963, n32964, n32965, n32966, n32967,
         n32968, n32969, n32970, n32971, n32972, n32973, n32974, n32975,
         n32976, n32977, n32978, n32979, n32980, n32981, n32982, n32983,
         n32984, n32985, n32986, n32987, n32988, n32989, n32990, n32991,
         n32992, n32993, n32994, n32995, n32996, n32997, n32998, n32999,
         n33000, n33001, n33002, n33003, n33004, n33005, n33006, n33007,
         n33008, n33009, n33010, n33011, n33012, n33013, n33014, n33015,
         n33016, n33017, n33018, n33019, n33020, n33021, n33022, n33023,
         n33024, n33025, n33026, n33027, n33028, n33029, n33030, n33031,
         n33032, n33033, n33034, n33035, n33036, n33037, n33038, n33039,
         n33040, n33041, n33042, n33043, n33044, n33045, n33046, n33047,
         n33048, n33049, n33050, n33051, n33052, n33053, n33054, n33055,
         n33056, n33057, n33058, n33059, n33060, n33061, n33062, n33063,
         n33064, n33065, n33066, n33067, n33068, n33069, n33070, n33071,
         n33072, n33073, n33074, n33075, n33076, n33077, n33078, n33079,
         n33080, n33081, n33082, n33083, n33084, n33085, n33086, n33087,
         n33088, n33089, n33090, n33091, n33092, n33093, n33094, n33095,
         n33096, n33097, n33098, n33099, n33100, n33101, n33102, n33103,
         n33104, n33105, n33106, n33107, n33108, n33109, n33110, n33111,
         n33112, n33113, n33114, n33115, n33116, n33117, n33118, n33119,
         n33120, n33121, n33122, n33123, n33124, n33125, n33126, n33127,
         n33128, n33129, n33130, n33131, n33132, n33133, n33134, n33135,
         n33136, n33137, n33138, n33139, n33140, n33141, n33142, n33143,
         n33144, n33145, n33146, n33147, n33148, n33149, n33150, n33151,
         n33152, n33153, n33154, n33155, n33156, n33157, n33158, n33159,
         n33160, n33161, n33162, n33163, n33164, n33165, n33166, n33167,
         n33168, n33169, n33170, n33171, n33172, n33173, n33174, n33175,
         n33176, n33177, n33178, n33179, n33180, n33181, n33182, n33183,
         n33184, n33185, n33186, n33187, n33188, n33189, n33190, n33191,
         n33192, n33193, n33194, n33195, n33196, n33197, n33198, n33199,
         n33200, n33201, n33202, n33203, n33204, n33205, n33206, n33207,
         n33208, n33209, n33210, n33211, n33212, n33213, n33214, n33215,
         n33216, n33217, n33218, n33219, n33220, n33221, n33222, n33223,
         n33224, n33225, n33226, n33227, n33228, n33229, n33230, n33231,
         n33232, n33233, n33234, n33235, n33236, n33237, n33238, n33239,
         n33240, n33241, n33242, n33243, n33244, n33245, n33246, n33247,
         n33248, n33249, n33250, n33251, n33252, n33253, n33254, n33255,
         n33256, n33257, n33258, n33259, n33260, n33261, n33262, n33263,
         n33264, n33265, n33266, n33267, n33268, n33269, n33270, n33271,
         n33272, n33273, n33274, n33275, n33276, n33277, n33278, n33279,
         n33280, n33281, n33282, n33283, n33284, n33285, n33286, n33287,
         n33288, n33289, n33290, n33291, n33292, n33293, n33294, n33295,
         n33296, n33297, n33298, n33299, n33300, n33301, n33302, n33303,
         n33304, n33305, n33306, n33307, n33308, n33309, n33310, n33311,
         n33312, n33313, n33314, n33315, n33316, n33317, n33318, n33319,
         n33320, n33321, n33322, n33323, n33324, n33325, n33326, n33327,
         n33328, n33329, n33330, n33331, n33332, n33333, n33334, n33335,
         n33336, n33337, n33338, n33339, n33340, n33341, n33342, n33343,
         n33344, n33345, n33346, n33347, n33348, n33349, n33350, n33351,
         n33352, n33353, n33354, n33355, n33356, n33357, n33358, n33359,
         n33360, n33361, n33362, n33363, n33364, n33365, n33366, n33367,
         n33368, n33369, n33370, n33371, n33372, n33373, n33374, n33375,
         n33376, n33377, n33378, n33379, n33380, n33381, n33382, n33383,
         n33384, n33385, n33386, n33387, n33388, n33389, n33390, n33391,
         n33392, n33393, n33394, n33395, n33396, n33397, n33398, n33399,
         n33400, n33401, n33402, n33403, n33404, n33405, n33406, n33407,
         n33408, n33409, n33410, n33411, n33412, n33413, n33414, n33415,
         n33416, n33417, n33418, n33419, n33420, n33421, n33422, n33423,
         n33424, n33425, n33426, n33427, n33428, n33429, n33430, n33431,
         n33432, n33433, n33434, n33435, n33436, n33437, n33438, n33439,
         n33440, n33441, n33442, n33443, n33444, n33445, n33446, n33447,
         n33448, n33449, n33450, n33451, n33452, n33453, n33454, n33455,
         n33456, n33457, n33458, n33459, n33460, n33461, n33462, n33463,
         n33464, n33465, n33466, n33467, n33468, n33469, n33470, n33471,
         n33472, n33473, n33474, n33475, n33476, n33477, n33478, n33479,
         n33480, n33481, n33482, n33483, n33484, n33485, n33486, n33487,
         n33488, n33489, n33490, n33491, n33492, n33493, n33494, n33495,
         n33496, n33497, n33498, n33499, n33500, n33501, n33502, n33503,
         n33504, n33505, n33506, n33507, n33508, n33509, n33510, n33511,
         n33512, n33513, n33514, n33515, n33516, n33517, n33518, n33519,
         n33520, n33521, n33522, n33523, n33524, n33525, n33526, n33527,
         n33528, n33529, n33530, n33531, n33532, n33533, n33534, n33535,
         n33536, n33537, n33538, n33539, n33540, n33541, n33542, n33543,
         n33544, n33545, n33546, n33547, n33548, n33549, n33550, n33551,
         n33552, n33553, n33554, n33555, n33556, n33557, n33558, n33559,
         n33560, n33561, n33562, n33563, n33564, n33565, n33566, n33567,
         n33568, n33569, n33570, n33571, n33572, n33573, n33574, n33575,
         n33576, n33577, n33578, n33579, n33580, n33581, n33582, n33583,
         n33584, n33585, n33586, n33587, n33588, n33589, n33590, n33591,
         n33592, n33593, n33594, n33595, n33596, n33597, n33598, n33599,
         n33600, n33601, n33602, n33603, n33604, n33605, n33606, n33607,
         n33608, n33609, n33610, n33611, n33612, n33613, n33614, n33615,
         n33616, n33617, n33618, n33619, n33620, n33621, n33622, n33623,
         n33624, n33625, n33626, n33627, n33628, n33629, n33630, n33631,
         n33632, n33633, n33634, n33635, n33636, n33637, n33638, n33639,
         n33640, n33641, n33642, n33643, n33644, n33645, n33646, n33647,
         n33648, n33649, n33650, n33651, n33652, n33653, n33654, n33655,
         n33656, n33657, n33658, n33659, n33660, n33661, n33662, n33663,
         n33664, n33665, n33666, n33667, n33668, n33669, n33670, n33671,
         n33672, n33673, n33674, n33675, n33676, n33677, n33678, n33679,
         n33680, n33681, n33682, n33683, n33684, n33685, n33686, n33687,
         n33688, n33689, n33690, n33691, n33692, n33693, n33694, n33695,
         n33696, n33697, n33698, n33699, n33700, n33701, n33702, n33703,
         n33704, n33705, n33706, n33707, n33708, n33709, n33710, n33711,
         n33712, n33713, n33714, n33715, n33716, n33717, n33718, n33719,
         n33720, n33721, n33722, n33723, n33724, n33725, n33726, n33727,
         n33728, n33729, n33730, n33731, n33732, n33733, n33734, n33735,
         n33736, n33737, n33738, n33739, n33740, n33741, n33742, n33743,
         n33744, n33745, n33746, n33747, n33748, n33749, n33750, n33751,
         n33752, n33753, n33754, n33755, n33756, n33757, n33758, n33759,
         n33760, n33761, n33762, n33763, n33764, n33765, n33766, n33767,
         n33768, n33769, n33770, n33771, n33772, n33773, n33774, n33775,
         n33776, n33777, n33778, n33779, n33780, n33781, n33782, n33783,
         n33784, n33785, n33786, n33787, n33788, n33789, n33790, n33791,
         n33792, n33793, n33794, n33795, n33796, n33797, n33798, n33799,
         n33800, n33801, n33802, n33803, n33804, n33805, n33806, n33807,
         n33808, n33809, n33810, n33811, n33812, n33813, n33814, n33815,
         n33816, n33817, n33818, n33819, n33820, n33821, n33822, n33823,
         n33824, n33825, n33826, n33827, n33828, n33829, n33830, n33831,
         n33832, n33833, n33834, n33835, n33836, n33837, n33838, n33839,
         n33840, n33841, n33842, n33843, n33844, n33845, n33846, n33847,
         n33848, n33849, n33850, n33851, n33852, n33853, n33854, n33855,
         n33856, n33857, n33858, n33859, n33860, n33861, n33862, n33863,
         n33864, n33865, n33866, n33867, n33868, n33869, n33870, n33871,
         n33872, n33873, n33874, n33875, n33876, n33877, n33878, n33879,
         n33880, n33881, n33882, n33883, n33884, n33885, n33886, n33887,
         n33888, n33889, n33890, n33891, n33892, n33893, n33894, n33895,
         n33896, n33897, n33898, n33899, n33900, n33901, n33902, n33903,
         n33904, n33905, n33906, n33907, n33908, n33909, n33910, n33911,
         n33912, n33913, n33914, n33915, n33916, n33917, n33918, n33919,
         n33920, n33921, n33922, n33923, n33924, n33925, n33926, n33927,
         n33928, n33929, n33930, n33931, n33932, n33933, n33934, n33935,
         n33936, n33937, n33938, n33939, n33940, n33941, n33942, n33943,
         n33944, n33945, n33946, n33947, n33948, n33949, n33950, n33951,
         n33952, n33953, n33954, n33955, n33956, n33957, n33958, n33959,
         n33960, n33961, n33962, n33963, n33964, n33965, n33966, n33967,
         n33968, n33969, n33970, n33971, n33972, n33973, n33974, n33975,
         n33976, n33977, n33978, n33979, n33980, n33981, n33982, n33983,
         n33984, n33985, n33986, n33987, n33988, n33989, n33990, n33991,
         n33992, n33993, n33994, n33995, n33996, n33997, n33998, n33999,
         n34000, n34001, n34002, n34003, n34004, n34005, n34006, n34007,
         n34008, n34009, n34010, n34011, n34012, n34013, n34014, n34015,
         n34016, n34017, n34018, n34019, n34020, n34021, n34022, n34023,
         n34024, n34025, n34026, n34027, n34028, n34029, n34030, n34031,
         n34032, n34033, n34034, n34035, n34036, n34037, n34038, n34039,
         n34040, n34041, n34042, n34043, n34044, n34045, n34046, n34047,
         n34048, n34049, n34050, n34051, n34052, n34053, n34054, n34055,
         n34056, n34057, n34058, n34059, n34060, n34061, n34062, n34063,
         n34064, n34065, n34066, n34067, n34068, n34069, n34070, n34071,
         n34072, n34073, n34074, n34075, n34076, n34077, n34078, n34079,
         n34080, n34081, n34082, n34083, n34084, n34085, n34086, n34087,
         n34088, n34089, n34090, n34091, n34092, n34093, n34094, n34095,
         n34096, n34097, n34098, n34099, n34100, n34101, n34102, n34103,
         n34104, n34105, n34106, n34107, n34108, n34109, n34110, n34111,
         n34112, n34113, n34114, n34115, n34116, n34117, n34118, n34119,
         n34120, n34121, n34122, n34123, n34124, n34125, n34126, n34127,
         n34128, n34129, n34130, n34131, n34132, n34133, n34134, n34135,
         n34136, n34137, n34138, n34139, n34140, n34141, n34142, n34143,
         n34144, n34145, n34146, n34147, n34148, n34149, n34150, n34151,
         n34152, n34153, n34154, n34155, n34156, n34157, n34158, n34159,
         n34160, n34161, n34162, n34163, n34164, n34165, n34166, n34167,
         n34168, n34169, n34170, n34171, n34172, n34173, n34174, n34175,
         n34176, n34177, n34178, n34179, n34180, n34181, n34182, n34183,
         n34184, n34185, n34186, n34187, n34188, n34189, n34190, n34191,
         n34192, n34193, n34194, n34195, n34196, n34197, n34198, n34199,
         n34200, n34201, n34202, n34203, n34204, n34205, n34206, n34207,
         n34208, n34209, n34210, n34211, n34212, n34213, n34214, n34215,
         n34216, n34217, n34218, n34219, n34220, n34221, n34222, n34223,
         n34224, n34225, n34226, n34227, n34228, n34229, n34230, n34231,
         n34232, n34233, n34234, n34235, n34236, n34237, n34238, n34239,
         n34240, n34241, n34242, n34243, n34244, n34245, n34246, n34247,
         n34248, n34249, n34250, n34251, n34252, n34253, n34254, n34255,
         n34256, n34257, n34258, n34259, n34260, n34261, n34262, n34263,
         n34264, n34265, n34266, n34267, n34268, n34269, n34270, n34271,
         n34272, n34273, n34274, n34275, n34276, n34277, n34278, n34279,
         n34280, n34281, n34282, n34283, n34284, n34285, n34286, n34287,
         n34288, n34289, n34290, n34291, n34292, n34293, n34294, n34295,
         n34296, n34297, n34298, n34299, n34300, n34301, n34302, n34303,
         n34304, n34305, n34306, n34307, n34308, n34309, n34310, n34311,
         n34312, n34313, n34314, n34315, n34316, n34317, n34318, n34319,
         n34320, n34321, n34322, n34323, n34324, n34325, n34326, n34327,
         n34328, n34329, n34330, n34331, n34332, n34333, n34334, n34335,
         n34336, n34337, n34338, n34339, n34340, n34341, n34342, n34343,
         n34344, n34345, n34346, n34347, n34348, n34349, n34350, n34351,
         n34352, n34353, n34354, n34355, n34356, n34357, n34358, n34359,
         n34360, n34361, n34362, n34363, n34364, n34365, n34366, n34367,
         n34368, n34369, n34370, n34371, n34372, n34373, n34374, n34375,
         n34376, n34377, n34378, n34379, n34380, n34381, n34382, n34383,
         n34384, n34385, n34386, n34387, n34388, n34389, n34390, n34391,
         n34392, n34393, n34394, n34395, n34396, n34397, n34398, n34399,
         n34400, n34401, n34402, n34403, n34404, n34405, n34406, n34407,
         n34408, n34409, n34410, n34411, n34412, n34413, n34414, n34415,
         n34416, n34417, n34418, n34419, n34420, n34421, n34422, n34423,
         n34424, n34425, n34426, n34427, n34428, n34429, n34430, n34431,
         n34432, n34433, n34434, n34435, n34436, n34437, n34438, n34439,
         n34440, n34441, n34442, n34443, n34444, n34445, n34446, n34447,
         n34448, n34449, n34450, n34451, n34452, n34453, n34454, n34455,
         n34456, n34457, n34458, n34459, n34460, n34461, n34462, n34463,
         n34464, n34465, n34466, n34467, n34468, n34469, n34470, n34471,
         n34472, n34473, n34474, n34475, n34476, n34477, n34478, n34479,
         n34480, n34481, n34482, n34483, n34484, n34485, n34486, n34487,
         n34488, n34489, n34490, n34491, n34492, n34493, n34494, n34495,
         n34496, n34497, n34498, n34499, n34500, n34501, n34502, n34503,
         n34504, n34505, n34506, n34507, n34508, n34509, n34510, n34511,
         n34512, n34513, n34514, n34515, n34516, n34517, n34518, n34519,
         n34520, n34521, n34522, n34523, n34524, n34525, n34526, n34527,
         n34528, n34529, n34530, n34531, n34532, n34533, n34534, n34535,
         n34536, n34537, n34538, n34539, n34540, n34541, n34542, n34543,
         n34544, n34545, n34546, n34547, n34548, n34549, n34550, n34551,
         n34552, n34553, n34554, n34555, n34556, n34557, n34558, n34559,
         n34560, n34561, n34562, n34563, n34564, n34565, n34566, n34567,
         n34568, n34569, n34570, n34571, n34572, n34573, n34574, n34575,
         n34576, n34577, n34578, n34579, n34580, n34581, n34582, n34583,
         n34584, n34585, n34586, n34587, n34588, n34589, n34590, n34591,
         n34592, n34593, n34594, n34595, n34596, n34597, n34598, n34599,
         n34600, n34601, n34602, n34603, n34604, n34605, n34606, n34607,
         n34608, n34609, n34610, n34611, n34612, n34613, n34614, n34615,
         n34616, n34617, n34618, n34619, n34620, n34621, n34622, n34623,
         n34624, n34625, n34626, n34627, n34628, n34629, n34630, n34631,
         n34632, n34633, n34634, n34635, n34636, n34637, n34638, n34639,
         n34640, n34641, n34642, n34643, n34644, n34645, n34646, n34647,
         n34648, n34649, n34650, n34651, n34652, n34653, n34654, n34655,
         n34656, n34657, n34658, n34659, n34660, n34661, n34662, n34663,
         n34664, n34665, n34666, n34667, n34668, n34669, n34670, n34671,
         n34672, n34673, n34674, n34675, n34676, n34677, n34678, n34679,
         n34680, n34681, n34682, n34683, n34684, n34685, n34686, n34687,
         n34688, n34689, n34690, n34691, n34692, n34693, n34694, n34695,
         n34696, n34697, n34698, n34699, n34700, n34701, n34702, n34703,
         n34704, n34705, n34706, n34707, n34708, n34709, n34710, n34711,
         n34712, n34713, n34714, n34715, n34716, n34717, n34718, n34719,
         n34720, n34721, n34722, n34723, n34724, n34725, n34726, n34727,
         n34728, n34729, n34730, n34731, n34732, n34733, n34734, n34735,
         n34736, n34737, n34738, n34739, n34740, n34741, n34742, n34743,
         n34744, n34745, n34746, n34747, n34748, n34749, n34750, n34751,
         n34752, n34753, n34754, n34755, n34756, n34757, n34758, n34759,
         n34760, n34761, n34762, n34763, n34764, n34765, n34766, n34767,
         n34768, n34769, n34770, n34771, n34772, n34773, n34774, n34775,
         n34776, n34777, n34778, n34779, n34780, n34781, n34782, n34783,
         n34784, n34785, n34786, n34787, n34788, n34789, n34790, n34791,
         n34792, n34793, n34794, n34795, n34796, n34797, n34798, n34799,
         n34800, n34801, n34802, n34803, n34804, n34805, n34806, n34807,
         n34808, n34809, n34810, n34811, n34812, n34813, n34814, n34815,
         n34816, n34817, n34818, n34819, n34820, n34821, n34822, n34823,
         n34824, n34825, n34826, n34827, n34828, n34829, n34830, n34831,
         n34832, n34833, n34834, n34835, n34836, n34837, n34838, n34839,
         n34840, n34841, n34842, n34843, n34844, n34845, n34846, n34847,
         n34848, n34849, n34850, n34851, n34852, n34853, n34854, n34855,
         n34856, n34857, n34858, n34859, n34860, n34861, n34862, n34863,
         n34864, n34865, n34866, n34867, n34868, n34869, n34870, n34871,
         n34872, n34873, n34874, n34875, n34876, n34877, n34878, n34879,
         n34880, n34881, n34882, n34883, n34884, n34885, n34886, n34887,
         n34888, n34889, n34890, n34891, n34892, n34893, n34894, n34895,
         n34896, n34897, n34898, n34899, n34900, n34901, n34902, n34903,
         n34904, n34905, n34906, n34907, n34908, n34909, n34910, n34911,
         n34912, n34913, n34914, n34915, n34916, n34917, n34918, n34919,
         n34920, n34921, n34922, n34923, n34924, n34925, n34926, n34927,
         n34928, n34929, n34930, n34931, n34932, n34933, n34934, n34935,
         n34936, n34937, n34938, n34939, n34940, n34941, n34942, n34943,
         n34944, n34945, n34946, n34947, n34948, n34949, n34950, n34951,
         n34952, n34953, n34954, n34955, n34956, n34957, n34958, n34959,
         n34960, n34961, n34962, n34963, n34964, n34965, n34966, n34967,
         n34968, n34969, n34970, n34971, n34972, n34973, n34974, n34975,
         n34976, n34977, n34978, n34979, n34980, n34981, n34982, n34983,
         n34984, n34985, n34986, n34987, n34988, n34989, n34990, n34991,
         n34992, n34993, n34994, n34995, n34996, n34997, n34998, n34999,
         n35000, n35001, n35002, n35003, n35004, n35005, n35006, n35007,
         n35008, n35009, n35010, n35011, n35012, n35013, n35014, n35015,
         n35016, n35017, n35018, n35019, n35020, n35021, n35022, n35023,
         n35024, n35025, n35026, n35027, n35028, n35029, n35030, n35031,
         n35032, n35033, n35034, n35035, n35036, n35037, n35038, n35039,
         n35040, n35041, n35042, n35043, n35044, n35045, n35046, n35047,
         n35048, n35049, n35050, n35051, n35052, n35053, n35054, n35055,
         n35056, n35057, n35058, n35059, n35060, n35061, n35062, n35063,
         n35064, n35065, n35066, n35067, n35068, n35069, n35070, n35071,
         n35072, n35073, n35074, n35075, n35076, n35077, n35078, n35079,
         n35080, n35081, n35082, n35083, n35084, n35085, n35086, n35087,
         n35088, n35089, n35090, n35091, n35092, n35093, n35094, n35095,
         n35096, n35097, n35098, n35099, n35100, n35101, n35102, n35103,
         n35104, n35105, n35106, n35107, n35108, n35109, n35110, n35111,
         n35112, n35113, n35114, n35115, n35116, n35117, n35118, n35119,
         n35120, n35121, n35122, n35123, n35124, n35125, n35126, n35127,
         n35128, n35129, n35130, n35131, n35132, n35133, n35134, n35135,
         n35136, n35137, n35138, n35139, n35140, n35141, n35142, n35143,
         n35144, n35145, n35146, n35147, n35148, n35149, n35150, n35151,
         n35152, n35153, n35154, n35155, n35156, n35157, n35158, n35159,
         n35160, n35161, n35162, n35163, n35164, n35165, n35166, n35167,
         n35168, n35169, n35170, n35171, n35172, n35173, n35174, n35175,
         n35176, n35177, n35178, n35179, n35180, n35181, n35182, n35183,
         n35184, n35185, n35186, n35187, n35188, n35189, n35190, n35191,
         n35192, n35193, n35194, n35195, n35196, n35197, n35198, n35199,
         n35200, n35201, n35202, n35203, n35204, n35205, n35206, n35207,
         n35208, n35209, n35210, n35211, n35212, n35213, n35214, n35215,
         n35216, n35217, n35218, n35219, n35220, n35221, n35222, n35223,
         n35224, n35225, n35226, n35227, n35228, n35229, n35230, n35231,
         n35232, n35233, n35234, n35235, n35236, n35237, n35238, n35239,
         n35240, n35241, n35242, n35243, n35244, n35245, n35246, n35247,
         n35248, n35249, n35250, n35251, n35252, n35253, n35254, n35255,
         n35256, n35257, n35258, n35259, n35260, n35261, n35262, n35263,
         n35264, n35265, n35266, n35267, n35268, n35269, n35270, n35271,
         n35272, n35273, n35274, n35275, n35276, n35277, n35278, n35279,
         n35280, n35281, n35282, n35283, n35284, n35285, n35286, n35287,
         n35288, n35289, n35290, n35291, n35292, n35293, n35294, n35295,
         n35296, n35297, n35298, n35299, n35300, n35301, n35302, n35303,
         n35304, n35305, n35306, n35307, n35308, n35309, n35310, n35311,
         n35312, n35313, n35314, n35315, n35316, n35317, n35318, n35319,
         n35320, n35321, n35322, n35323, n35324, n35325, n35326, n35327,
         n35328, n35329, n35330, n35331, n35332, n35333, n35334, n35335,
         n35336, n35337, n35338, n35339, n35340, n35341, n35342, n35343,
         n35344, n35345, n35346, n35347, n35348, n35349, n35350, n35351,
         n35352, n35353, n35354, n35355, n35356, n35357, n35358, n35359,
         n35360, n35361, n35362, n35363, n35364, n35365, n35366, n35367,
         n35368, n35369, n35370, n35371, n35372, n35373, n35374, n35375,
         n35376, n35377, n35378, n35379, n35380, n35381, n35382, n35383,
         n35384, n35385, n35386, n35387, n35388, n35389, n35390, n35391,
         n35392, n35393, n35394, n35395, n35396, n35397, n35398, n35399,
         n35400, n35401, n35402, n35403, n35404, n35405, n35406, n35407,
         n35408, n35409, n35410, n35411, n35412, n35413, n35414, n35415,
         n35416, n35417, n35418, n35419, n35420, n35421, n35422, n35423,
         n35424, n35425, n35426, n35427, n35428, n35429, n35430, n35431,
         n35432, n35433, n35434, n35435, n35436, n35437, n35438, n35439,
         n35440, n35441, n35442, n35443, n35444, n35445, n35446, n35447,
         n35448, n35449, n35450, n35451, n35452, n35453, n35454, n35455,
         n35456, n35457, n35458, n35459, n35460, n35461, n35462, n35463,
         n35464, n35465, n35466, n35467, n35468, n35469, n35470, n35471,
         n35472, n35473, n35474, n35475, n35476, n35477, n35478, n35479,
         n35480, n35481, n35482, n35483, n35484, n35485, n35486, n35487,
         n35488, n35489, n35490, n35491, n35492, n35493, n35494, n35495,
         n35496, n35497, n35498, n35499, n35500, n35501, n35502, n35503,
         n35504, n35505, n35506, n35507, n35508, n35509, n35510, n35511,
         n35512, n35513, n35514, n35515, n35516, n35517, n35518, n35519,
         n35520, n35521, n35522, n35523, n35524, n35525, n35526, n35527,
         n35528, n35529, n35530, n35531, n35532, n35533, n35534, n35535,
         n35536, n35537, n35538, n35539, n35540, n35541, n35542, n35543,
         n35544, n35545, n35546, n35547, n35548, n35549, n35550, n35551,
         n35552, n35553, n35554, n35555, n35556, n35557, n35558, n35559,
         n35560, n35561, n35562, n35563, n35564, n35565, n35566, n35567,
         n35568, n35569, n35570, n35571, n35572, n35573, n35574, n35575,
         n35576, n35577, n35578, n35579, n35580, n35581, n35582, n35583,
         n35584, n35585, n35586, n35587, n35588, n35589, n35590, n35591,
         n35592, n35593, n35594, n35595, n35596, n35597, n35598, n35599,
         n35600, n35601, n35602, n35603, n35604, n35605, n35606, n35607,
         n35608, n35609, n35610, n35611, n35612, n35613, n35614, n35615,
         n35616, n35617, n35618, n35619, n35620, n35621, n35622, n35623,
         n35624, n35625, n35626, n35627, n35628, n35629, n35630, n35631,
         n35632, n35633, n35634, n35635, n35636, n35637, n35638, n35639,
         n35640, n35641, n35642, n35643, n35644, n35645, n35646, n35647,
         n35648, n35649, n35650, n35651, n35652, n35653, n35654, n35655,
         n35656, n35657, n35658, n35659, n35660, n35661, n35662, n35663,
         n35664, n35665, n35666, n35667, n35668, n35669, n35670, n35671,
         n35672, n35673, n35674, n35675, n35676, n35677, n35678, n35679,
         n35680, n35681, n35682, n35683, n35684, n35685, n35686, n35687,
         n35688, n35689, n35690, n35691, n35692, n35693, n35694, n35695,
         n35696, n35697, n35698, n35699, n35700, n35701, n35702, n35703,
         n35704, n35705, n35706, n35707, n35708, n35709, n35710, n35711,
         n35712, n35713, n35714, n35715, n35716, n35717, n35718, n35719,
         n35720, n35721, n35722, n35723, n35724, n35725, n35726, n35727,
         n35728, n35729, n35730, n35731, n35732, n35733, n35734, n35735,
         n35736, n35737, n35738, n35739, n35740, n35741, n35742, n35743,
         n35744, n35745, n35746, n35747, n35748, n35749, n35750, n35751,
         n35752, n35753, n35754, n35755, n35756, n35757, n35758, n35759,
         n35760, n35761, n35762, n35763, n35764, n35765, n35766, n35767,
         n35768, n35769, n35770, n35771, n35772, n35773, n35774, n35775,
         n35776, n35777, n35778, n35779, n35780, n35781, n35782, n35783,
         n35784, n35785, n35786, n35787, n35788, n35789, n35790, n35791,
         n35792, n35793, n35794, n35795, n35796, n35797, n35798, n35799,
         n35800, n35801, n35802, n35803, n35804, n35805, n35806, n35807,
         n35808, n35809, n35810, n35811, n35812, n35813, n35814, n35815,
         n35816, n35817, n35818, n35819, n35820, n35821, n35822, n35823,
         n35824, n35825, n35826, n35827, n35828, n35829, n35830, n35831,
         n35832, n35833, n35834, n35835, n35836, n35837, n35838, n35839,
         n35840, n35841, n35842, n35843, n35844, n35845, n35846, n35847,
         n35848, n35849, n35850, n35851, n35852, n35853, n35854, n35855,
         n35856, n35857, n35858, n35859, n35860, n35861, n35862, n35863,
         n35864, n35865, n35866, n35867, n35868, n35869, n35870, n35871,
         n35872, n35873, n35874, n35875, n35876, n35877, n35878, n35879,
         n35880, n35881, n35882, n35883, n35884, n35885, n35886, n35887,
         n35888, n35889, n35890, n35891, n35892, n35893, n35894, n35895,
         n35896, n35897, n35898, n35899, n35900, n35901, n35902, n35903,
         n35904, n35905, n35906, n35907, n35908, n35909, n35910, n35911,
         n35912, n35913, n35914, n35915, n35916, n35917, n35918, n35919,
         n35920, n35921, n35922, n35923, n35924, n35925, n35926, n35927,
         n35928, n35929, n35930, n35931, n35932, n35933, n35934, n35935,
         n35936, n35937, n35938, n35939, n35940, n35941, n35942, n35943,
         n35944, n35945, n35946, n35947, n35948, n35949, n35950, n35951,
         n35952, n35953, n35954, n35955, n35956, n35957, n35958, n35959,
         n35960, n35961, n35962, n35963, n35964, n35965, n35966, n35967,
         n35968, n35969, n35970, n35971, n35972, n35973, n35974, n35975,
         n35976, n35977, n35978, n35979, n35980, n35981, n35982, n35983,
         n35984, n35985, n35986, n35987, n35988, n35989, n35990, n35991,
         n35992, n35993, n35994, n35995, n35996, n35997, n35998, n35999,
         n36000, n36001, n36002, n36003, n36004, n36005, n36006, n36007,
         n36008, n36009, n36010, n36011, n36012, n36013, n36014, n36015,
         n36016, n36017, n36018, n36019, n36020, n36021, n36022, n36023,
         n36024, n36025, n36026, n36027, n36028, n36029, n36030, n36031,
         n36032, n36033, n36034, n36035, n36036, n36037, n36038, n36039,
         n36040, n36041, n36042, n36043, n36044, n36045, n36046, n36047,
         n36048, n36049, n36050, n36051, n36052, n36053, n36054, n36055,
         n36056, n36057, n36058, n36059, n36060, n36061, n36062, n36063,
         n36064, n36065, n36066, n36067, n36068, n36069, n36070, n36071,
         n36072, n36073, n36074, n36075, n36076, n36077, n36078, n36079,
         n36080, n36081, n36082, n36083, n36084, n36085, n36086, n36087,
         n36088, n36089, n36090, n36091, n36092, n36093, n36094, n36095,
         n36096, n36097, n36098, n36099, n36100, n36101, n36102, n36103,
         n36104, n36105, n36106, n36107, n36108, n36109, n36110, n36111,
         n36112, n36113, n36114, n36115, n36116, n36117, n36118, n36119,
         n36120, n36121, n36122, n36123, n36124, n36125, n36126, n36127,
         n36128, n36129, n36130, n36131, n36132, n36133, n36134, n36135,
         n36136, n36137, n36138, n36139, n36140, n36141, n36142, n36143,
         n36144, n36145, n36146, n36147, n36148, n36149, n36150, n36151,
         n36152, n36153, n36154, n36155, n36156, n36157, n36158, n36159,
         n36160, n36161, n36162, n36163, n36164, n36165, n36166, n36167,
         n36168, n36169, n36170, n36171, n36172, n36173, n36174, n36175,
         n36176, n36177, n36178, n36179, n36180, n36181, n36182, n36183,
         n36184, n36185, n36186, n36187, n36188, n36189, n36190, n36191,
         n36192, n36193, n36194, n36195, n36196, n36197, n36198, n36199,
         n36200, n36201, n36202, n36203, n36204, n36205, n36206, n36207,
         n36208, n36209, n36210, n36211, n36212, n36213, n36214, n36215,
         n36216, n36217, n36218, n36219, n36220, n36221, n36222, n36223,
         n36224, n36225, n36226, n36227, n36228, n36229, n36230, n36231,
         n36232, n36233, n36234, n36235, n36236, n36237, n36238, n36239,
         n36240, n36241, n36242, n36243, n36244, n36245, n36246, n36247,
         n36248, n36249, n36250, n36251, n36252, n36253, n36254, n36255,
         n36256, n36257, n36258, n36259, n36260, n36261, n36262, n36263,
         n36264, n36265, n36266, n36267, n36268, n36269, n36270, n36271,
         n36272, n36273, n36274, n36275, n36276, n36277, n36278, n36279,
         n36280, n36281, n36282, n36283, n36284, n36285, n36286, n36287,
         n36288, n36289, n36290, n36291, n36292, n36293, n36294, n36295,
         n36296, n36297, n36298, n36299, n36300, n36301, n36302, n36303,
         n36304, n36305, n36306, n36307, n36308, n36309, n36310, n36311,
         n36312, n36313, n36314, n36315, n36316, n36317, n36318, n36319,
         n36320, n36321, n36322, n36323, n36324, n36325, n36326, n36327,
         n36328, n36329, n36330, n36331, n36332, n36333, n36334, n36335,
         n36336, n36337, n36338, n36339, n36340, n36341, n36342, n36343,
         n36344, n36345, n36346, n36347, n36348, n36349, n36350, n36351,
         n36352, n36353, n36354, n36355, n36356, n36357, n36358, n36359,
         n36360, n36361, n36362, n36363, n36364, n36365, n36366, n36367,
         n36368, n36369, n36370, n36371, n36372, n36373, n36374, n36375,
         n36376, n36377, n36378, n36379, n36380, n36381, n36382, n36383,
         n36384, n36385, n36386, n36387, n36388, n36389, n36390, n36391,
         n36392, n36393, n36394, n36395, n36396, n36397, n36398, n36399,
         n36400, n36401, n36402, n36403, n36404, n36405, n36406, n36407,
         n36408, n36409, n36410, n36411, n36412, n36413, n36414, n36415,
         n36416, n36417, n36418, n36419, n36420, n36421, n36422, n36423,
         n36424, n36425, n36426, n36427, n36428, n36429, n36430, n36431,
         n36432, n36433, n36434, n36435, n36436, n36437, n36438, n36439,
         n36440, n36441, n36442, n36443, n36444, n36445, n36446, n36447,
         n36448, n36449, n36450, n36451, n36452, n36453, n36454, n36455,
         n36456, n36457, n36458, n36459, n36460, n36461, n36462, n36463,
         n36464, n36465, n36466, n36467, n36468, n36469, n36470, n36471,
         n36472, n36473, n36474, n36475, n36476, n36477, n36478, n36479,
         n36480, n36481, n36482, n36483, n36484, n36485, n36486, n36487,
         n36488, n36489, n36490, n36491, n36492, n36493, n36494, n36495,
         n36496, n36497, n36498, n36499, n36500, n36501, n36502, n36503,
         n36504, n36505, n36506, n36507, n36508, n36509, n36510, n36511,
         n36512, n36513, n36514, n36515, n36516, n36517, n36518, n36519,
         n36520, n36521, n36522, n36523, n36524, n36525, n36526, n36527,
         n36528, n36529, n36530, n36531, n36532, n36533, n36534, n36535,
         n36536, n36537, n36538, n36539, n36540, n36541, n36542, n36543,
         n36544, n36545, n36546, n36547, n36548, n36549, n36550, n36551,
         n36552, n36553, n36554, n36555, n36556, n36557, n36558, n36559,
         n36560, n36561, n36562, n36563, n36564, n36565, n36566, n36567,
         n36568, n36569, n36570, n36571, n36572, n36573, n36574, n36575,
         n36576, n36577, n36578, n36579, n36580, n36581, n36582, n36583,
         n36584, n36585, n36586, n36587, n36588, n36589, n36590, n36591,
         n36592, n36593, n36594, n36595, n36596, n36597, n36598, n36599,
         n36600, n36601, n36602, n36603, n36604, n36605, n36606, n36607,
         n36608, n36609, n36610, n36611, n36612, n36613, n36614, n36615,
         n36616, n36617, n36618, n36619, n36620, n36621, n36622, n36623,
         n36624, n36625, n36626, n36627, n36628, n36629, n36630, n36631,
         n36632, n36633, n36634, n36635, n36636, n36637, n36638, n36639,
         n36640, n36641, n36642, n36643, n36644, n36645, n36646, n36647,
         n36648, n36649, n36650, n36651, n36652, n36653, n36654, n36655,
         n36656, n36657, n36658, n36659, n36660, n36661, n36662, n36663,
         n36664, n36665, n36666, n36667, n36668, n36669, n36670, n36671,
         n36672, n36673, n36674, n36675, n36676, n36677, n36678, n36679,
         n36680, n36681, n36682, n36683, n36684, n36685, n36686, n36687,
         n36688, n36689, n36690, n36691, n36692, n36693, n36694, n36695,
         n36696, n36697, n36698, n36699, n36700, n36701, n36702, n36703,
         n36704, n36705, n36706, n36707, n36708, n36709, n36710, n36711,
         n36712, n36713, n36714, n36715, n36716, n36717, n36718, n36719,
         n36720, n36721, n36722, n36723, n36724, n36725, n36726, n36727,
         n36728, n36729, n36730, n36731, n36732, n36733, n36734, n36735,
         n36736, n36737, n36738, n36739, n36740, n36741, n36742, n36743,
         n36744, n36745, n36746, n36747, n36748, n36749, n36750, n36751,
         n36752, n36753, n36754, n36755, n36756, n36757, n36758, n36759,
         n36760, n36761, n36762, n36763, n36764, n36765, n36766, n36767,
         n36768, n36769, n36770, n36771, n36772, n36773, n36774, n36775,
         n36776, n36777, n36778, n36779, n36780, n36781, n36782, n36783,
         n36784, n36785, n36786, n36787, n36788, n36789, n36790, n36791,
         n36792, n36793, n36794, n36795, n36796, n36797, n36798, n36799,
         n36800, n36801, n36802, n36803, n36804, n36805, n36806, n36807,
         n36808, n36809, n36810, n36811, n36812, n36813, n36814, n36815,
         n36816, n36817, n36818, n36819, n36820, n36821, n36822, n36823,
         n36824, n36825, n36826, n36827, n36828, n36829, n36830, n36831,
         n36832, n36833, n36834, n36835, n36836, n36837, n36838, n36839,
         n36840, n36841, n36842, n36843, n36844, n36845, n36846, n36847,
         n36848, n36849, n36850, n36851, n36852, n36853, n36854, n36855,
         n36856, n36857, n36858, n36859, n36860, n36861, n36862, n36863,
         n36864, n36865, n36866, n36867, n36868, n36869, n36870, n36871,
         n36872, n36873, n36874, n36875, n36876, n36877, n36878, n36879,
         n36880, n36881, n36882, n36883, n36884, n36885, n36886, n36887,
         n36888, n36889, n36890, n36891, n36892, n36893, n36894, n36895,
         n36896, n36897, n36898, n36899, n36900, n36901, n36902, n36903,
         n36904, n36905, n36906, n36907, n36908, n36909, n36910, n36911,
         n36912, n36913, n36914, n36915, n36916, n36917, n36918, n36919,
         n36920, n36921, n36922, n36923, n36924, n36925, n36926, n36927,
         n36928, n36929, n36930, n36931, n36932, n36933, n36934, n36935,
         n36936, n36937, n36938, n36939, n36940, n36941, n36942, n36943,
         n36944, n36945, n36946, n36947, n36948, n36949, n36950, n36951,
         n36952, n36953, n36954, n36955, n36956, n36957, n36958, n36959,
         n36960, n36961, n36962, n36963, n36964, n36965, n36966, n36967,
         n36968, n36969, n36970, n36971, n36972, n36973, n36974, n36975,
         n36976, n36977, n36978, n36979, n36980, n36981, n36982, n36983,
         n36984, n36985, n36986, n36987, n36988, n36989, n36990, n36991,
         n36992, n36993, n36994, n36995, n36996, n36997, n36998, n36999,
         n37000, n37001, n37002, n37003, n37004, n37005, n37006, n37007,
         n37008, n37009, n37010, n37011, n37012, n37013, n37014, n37015,
         n37016, n37017, n37018, n37019, n37020, n37021, n37022, n37023,
         n37024, n37025, n37026, n37027, n37028, n37029, n37030, n37031,
         n37032, n37033, n37034, n37035, n37036, n37037, n37038, n37039,
         n37040, n37041, n37042, n37043, n37044, n37045, n37046, n37047,
         n37048, n37049, n37050, n37051, n37052, n37053, n37054, n37055,
         n37056, n37057, n37058, n37059, n37060, n37061, n37062, n37063,
         n37064, n37065, n37066, n37067, n37068, n37069, n37070, n37071,
         n37072, n37073, n37074, n37075, n37076, n37077, n37078, n37079,
         n37080, n37081, n37082, n37083, n37084, n37085, n37086, n37087,
         n37088, n37089, n37090, n37091, n37092, n37093, n37094, n37095,
         n37096, n37097, n37098, n37099, n37100, n37101, n37102, n37103,
         n37104, n37105, n37106, n37107, n37108, n37109, n37110, n37111,
         n37112, n37113, n37114, n37115, n37116, n37117, n37118, n37119,
         n37120, n37121, n37122, n37123, n37124, n37125, n37126, n37127,
         n37128, n37129, n37130, n37131, n37132, n37133, n37134, n37135,
         n37136, n37137, n37138, n37139, n37140, n37141, n37142, n37143,
         n37144, n37145, n37146, n37147, n37148, n37149, n37150, n37151,
         n37152, n37153, n37154, n37155, n37156, n37157, n37158, n37159,
         n37160, n37161, n37162, n37163, n37164, n37165, n37166, n37167,
         n37168, n37169, n37170, n37171, n37172, n37173, n37174, n37175,
         n37176, n37177, n37178, n37179, n37180, n37181, n37182, n37183,
         n37184, n37185, n37186, n37187, n37188, n37189, n37190, n37191,
         n37192, n37193, n37194, n37195, n37196, n37197, n37198, n37199,
         n37200, n37201, n37202, n37203, n37204, n37205, n37206, n37207,
         n37208, n37209, n37210, n37211, n37212, n37213, n37214, n37215,
         n37216, n37217, n37218, n37219, n37220, n37221, n37222, n37223,
         n37224, n37225, n37226, n37227, n37228, n37229, n37230, n37231,
         n37232, n37233, n37234, n37235, n37236, n37237, n37238, n37239,
         n37240, n37241, n37242, n37243, n37244, n37245, n37246, n37247,
         n37248, n37249, n37250, n37251, n37252, n37253, n37254, n37255,
         n37256, n37257, n37258, n37259, n37260, n37261, n37262, n37263,
         n37264, n37265, n37266, n37267, n37268, n37269, n37270, n37271,
         n37272, n37273, n37274, n37275, n37276, n37277, n37278, n37279,
         n37280, n37281, n37282, n37283, n37284, n37285, n37286, n37287,
         n37288, n37289, n37290, n37291, n37292, n37293, n37294, n37295,
         n37296, n37297, n37298, n37299, n37300, n37301, n37302, n37303,
         n37304, n37305, n37306, n37307, n37308, n37309, n37310, n37311,
         n37312, n37313, n37314, n37315, n37316, n37317, n37318, n37319,
         n37320, n37321, n37322, n37323, n37324, n37325, n37326, n37327,
         n37328, n37329, n37330, n37331, n37332, n37333, n37334, n37335,
         n37336, n37337, n37338, n37339, n37340, n37341, n37342, n37343,
         n37344, n37345, n37346, n37347, n37348, n37349, n37350, n37351,
         n37352, n37353, n37354, n37355, n37356, n37357, n37358, n37359,
         n37360, n37361, n37362, n37363, n37364, n37365, n37366, n37367,
         n37368, n37369, n37370, n37371, n37372, n37373, n37374, n37375,
         n37376, n37377, n37378, n37379, n37380, n37381, n37382, n37383,
         n37384, n37385, n37386, n37387, n37388, n37389, n37390, n37391,
         n37392, n37393, n37394, n37395, n37396, n37397, n37398, n37399,
         n37400, n37401, n37402, n37403, n37404, n37405, n37406, n37407,
         n37408, n37409, n37410, n37411, n37412, n37413, n37414, n37415,
         n37416, n37417, n37418, n37419, n37420, n37421, n37422, n37423,
         n37424, n37425, n37426, n37427, n37428, n37429, n37430, n37431,
         n37432, n37433, n37434, n37435, n37436, n37437, n37438, n37439,
         n37440, n37441, n37442, n37443, n37444, n37445, n37446, n37447,
         n37448, n37449, n37450, n37451, n37452, n37453, n37454, n37455,
         n37456, n37457, n37458, n37459, n37460, n37461, n37462, n37463,
         n37464, n37465, n37466, n37467, n37468, n37469, n37470, n37471,
         n37472, n37473, n37474, n37475, n37476, n37477, n37478, n37479,
         n37480, n37481, n37482, n37483, n37484, n37485, n37486, n37487,
         n37488, n37489, n37490, n37491, n37492, n37493, n37494, n37495,
         n37496, n37497, n37498, n37499, n37500, n37501, n37502, n37503,
         n37504, n37505, n37506, n37507, n37508, n37509, n37510, n37511,
         n37512, n37513, n37514, n37515, n37516, n37517, n37518, n37519,
         n37520, n37521, n37522, n37523, n37524, n37525, n37526, n37527,
         n37528, n37529, n37530, n37531, n37532, n37533, n37534, n37535,
         n37536, n37537, n37538, n37539, n37540, n37541, n37542, n37543,
         n37544, n37545, n37546, n37547, n37548, n37549, n37550, n37551,
         n37552, n37553, n37554, n37555, n37556, n37557, n37558, n37559,
         n37560, n37561, n37562, n37563, n37564, n37565, n37566, n37567,
         n37568, n37569, n37570, n37571, n37572, n37573, n37574, n37575,
         n37576, n37577, n37578, n37579, n37580, n37581, n37582, n37583,
         n37584, n37585, n37586, n37587, n37588, n37589, n37590, n37591,
         n37592, n37593, n37594, n37595, n37596, n37597, n37598, n37599,
         n37600, n37601, n37602, n37603, n37604, n37605, n37606, n37607,
         n37608, n37609, n37610, n37611, n37612, n37613, n37614, n37615,
         n37616, n37617, n37618, n37619, n37620, n37621, n37622, n37623,
         n37624, n37625, n37626, n37627, n37628, n37629, n37630, n37631,
         n37632, n37633, n37634, n37635, n37636, n37637, n37638, n37639,
         n37640, n37641, n37642, n37643, n37644, n37645, n37646, n37647,
         n37648, n37649, n37650, n37651, n37652, n37653, n37654, n37655,
         n37656, n37657, n37658, n37659, n37660, n37661, n37662, n37663,
         n37664, n37665, n37666, n37667, n37668, n37669, n37670, n37671,
         n37672, n37673, n37674, n37675, n37676, n37677, n37678, n37679,
         n37680, n37681, n37682, n37683, n37684, n37685, n37686, n37687,
         n37688, n37689, n37690, n37691, n37692, n37693, n37694, n37695,
         n37696, n37697, n37698, n37699, n37700, n37701, n37702, n37703,
         n37704, n37705, n37706, n37707, n37708, n37709, n37710, n37711,
         n37712, n37713, n37714, n37715, n37716, n37717, n37718, n37719,
         n37720, n37721, n37722, n37723, n37724, n37725, n37726, n37727,
         n37728, n37729, n37730, n37731, n37732, n37733, n37734, n37735,
         n37736, n37737, n37738, n37739, n37740, n37741, n37742, n37743,
         n37744, n37745, n37746, n37747, n37748, n37749, n37750, n37751,
         n37752, n37753, n37754, n37755, n37756, n37757, n37758, n37759,
         n37760, n37761, n37762, n37763, n37764, n37765, n37766, n37767,
         n37768, n37769, n37770, n37771, n37772, n37773, n37774, n37775,
         n37776, n37777, n37778, n37779, n37780, n37781, n37782, n37783,
         n37784, n37785, n37786, n37787, n37788, n37789, n37790, n37791,
         n37792, n37793, n37794, n37795, n37796, n37797, n37798, n37799,
         n37800, n37801, n37802, n37803, n37804, n37805, n37806, n37807,
         n37808, n37809, n37810, n37811, n37812, n37813, n37814, n37815,
         n37816, n37817, n37818, n37819, n37820, n37821, n37822, n37823,
         n37824, n37825, n37826, n37827, n37828, n37829, n37830, n37831,
         n37832, n37833, n37834, n37835, n37836, n37837, n37838, n37839,
         n37840, n37841, n37842, n37843, n37844, n37845, n37846, n37847,
         n37848, n37849, n37850, n37851, n37852, n37853, n37854, n37855,
         n37856, n37857, n37858, n37859, n37860, n37861, n37862, n37863,
         n37864, n37865, n37866, n37867, n37868, n37869, n37870, n37871,
         n37872, n37873, n37874, n37875, n37876, n37877, n37878, n37879,
         n37880, n37881, n37882, n37883, n37884, n37885, n37886, n37887,
         n37888, n37889, n37890, n37891, n37892, n37893, n37894, n37895,
         n37896, n37897, n37898, n37899, n37900, n37901, n37902, n37903,
         n37904, n37905, n37906, n37907, n37908, n37909, n37910, n37911,
         n37912, n37913, n37914, n37915, n37916, n37917, n37918, n37919,
         n37920, n37921, n37922, n37923, n37924, n37925, n37926, n37927,
         n37928, n37929, n37930, n37931, n37932, n37933, n37934, n37935,
         n37936, n37937, n37938, n37939, n37940, n37941, n37942, n37943,
         n37944, n37945, n37946, n37947, n37948, n37949, n37950, n37951,
         n37952, n37953, n37954, n37955, n37956, n37957, n37958, n37959,
         n37960, n37961, n37962, n37963, n37964, n37965, n37966, n37967,
         n37968, n37969, n37970, n37971, n37972, n37973, n37974, n37975,
         n37976, n37977, n37978, n37979, n37980, n37981, n37982, n37983,
         n37984, n37985, n37986, n37987, n37988, n37989, n37990, n37991,
         n37992, n37993, n37994, n37995, n37996, n37997, n37998, n37999,
         n38000, n38001, n38002, n38003, n38004, n38005, n38006, n38007,
         n38008, n38009, n38010, n38011, n38012, n38013, n38014, n38015,
         n38016, n38017, n38018, n38019, n38020, n38021, n38022, n38023,
         n38024, n38025, n38026, n38027, n38028, n38029, n38030, n38031,
         n38032, n38033, n38034, n38035, n38036, n38037, n38038, n38039,
         n38040, n38041, n38042, n38043, n38044, n38045, n38046, n38047,
         n38048, n38049, n38050, n38051, n38052, n38053, n38054, n38055,
         n38056, n38057, n38058, n38059, n38060, n38061, n38062, n38063,
         n38064, n38065, n38066, n38067, n38068, n38069, n38070, n38071,
         n38072, n38073, n38074, n38075, n38076, n38077, n38078, n38079,
         n38080, n38081, n38082, n38083, n38084, n38085, n38086, n38087,
         n38088, n38089, n38090, n38091, n38092, n38093, n38094, n38095,
         n38096, n38097, n38098, n38099, n38100, n38101, n38102, n38103,
         n38104, n38105, n38106, n38107, n38108, n38109, n38110, n38111,
         n38112, n38113, n38114, n38115, n38116, n38117, n38118, n38119,
         n38120, n38121, n38122, n38123, n38124, n38125, n38126, n38127,
         n38128, n38129, n38130, n38131, n38132, n38133, n38134, n38135,
         n38136, n38137, n38138, n38139, n38140, n38141, n38142, n38143,
         n38144, n38145, n38146, n38147, n38148, n38149, n38150, n38151,
         n38152, n38153, n38154, n38155, n38156, n38157, n38158, n38159,
         n38160, n38161, n38162, n38163, n38164, n38165, n38166, n38167,
         n38168, n38169, n38170, n38171, n38172, n38173, n38174, n38175,
         n38176, n38177, n38178, n38179, n38180, n38181, n38182, n38183,
         n38184, n38185, n38186, n38187, n38188, n38189, n38190, n38191,
         n38192, n38193, n38194, n38195, n38196, n38197, n38198, n38199,
         n38200, n38201, n38202, n38203, n38204, n38205, n38206, n38207,
         n38208, n38209, n38210, n38211, n38212, n38213, n38214, n38215,
         n38216, n38217, n38218, n38219, n38220, n38221, n38222, n38223,
         n38224, n38225, n38226, n38227, n38228, n38229, n38230, n38231,
         n38232, n38233, n38234, n38235, n38236, n38237, n38238, n38239,
         n38240, n38241, n38242, n38243, n38244, n38245, n38246, n38247,
         n38248, n38249, n38250, n38251, n38252, n38253, n38254, n38255,
         n38256, n38257, n38258, n38259, n38260, n38261, n38262, n38263,
         n38264, n38265, n38266, n38267, n38268, n38269, n38270, n38271,
         n38272, n38273, n38274, n38275, n38276, n38277, n38278, n38279,
         n38280, n38281, n38282, n38283, n38284, n38285, n38286, n38287,
         n38288, n38289, n38290, n38291, n38292, n38293, n38294, n38295,
         n38296, n38297, n38298, n38299, n38300, n38301, n38302, n38303,
         n38304, n38305, n38306, n38307, n38308, n38309, n38310, n38311,
         n38312, n38313, n38314, n38315, n38316, n38317, n38318, n38319,
         n38320, n38321, n38322, n38323, n38324, n38325, n38326, n38327,
         n38328, n38329, n38330, n38331, n38332, n38333, n38334, n38335,
         n38336, n38337, n38338, n38339, n38340, n38341, n38342, n38343,
         n38344, n38345, n38346, n38347, n38348, n38349, n38350, n38351,
         n38352, n38353, n38354, n38355, n38356, n38357, n38358, n38359,
         n38360, n38361, n38362, n38363, n38364, n38365, n38366, n38367,
         n38368, n38369, n38370, n38371, n38372, n38373, n38374, n38375,
         n38376, n38377, n38378, n38379, n38380, n38381, n38382, n38383,
         n38384, n38385, n38386, n38387, n38388, n38389, n38390, n38391,
         n38392, n38393, n38394, n38395, n38396, n38397, n38398, n38399,
         n38400, n38401, n38402, n38403, n38404, n38405, n38406, n38407,
         n38408, n38409, n38410, n38411, n38412, n38413, n38414, n38415,
         n38416, n38417, n38418, n38419, n38420, n38421, n38422, n38423,
         n38424, n38425, n38426, n38427, n38428, n38429, n38430, n38431,
         n38432, n38433, n38434, n38435, n38436, n38437, n38438, n38439,
         n38440, n38441, n38442, n38443, n38444, n38445, n38446, n38447,
         n38448, n38449, n38450, n38451, n38452, n38453, n38454, n38455,
         n38456, n38457, n38458, n38459, n38460, n38461, n38462, n38463,
         n38464, n38465, n38466, n38467, n38468, n38469, n38470, n38471,
         n38472, n38473, n38474, n38475, n38476, n38477, n38478, n38479,
         n38480, n38481, n38482, n38483, n38484, n38485, n38486, n38487,
         n38488, n38489, n38490, n38491, n38492, n38493, n38494, n38495,
         n38496, n38497, n38498, n38499, n38500, n38501, n38502, n38503,
         n38504, n38505, n38506, n38507, n38508, n38509, n38510, n38511,
         n38512, n38513, n38514, n38515, n38516, n38517, n38518, n38519,
         n38520, n38521, n38522, n38523, n38524, n38525, n38526, n38527,
         n38528, n38529, n38530, n38531, n38532, n38533, n38534, n38535,
         n38536, n38537, n38538, n38539, n38540, n38541, n38542, n38543,
         n38544, n38545, n38546, n38547, n38548, n38549, n38550, n38551,
         n38552, n38553, n38554, n38555, n38556, n38557, n38558, n38559,
         n38560, n38561, n38562, n38563, n38564, n38565, n38566, n38567,
         n38568, n38569, n38570, n38571, n38572, n38573, n38574, n38575,
         n38576, n38577, n38578, n38579, n38580, n38581, n38582, n38583,
         n38584, n38585, n38586, n38587, n38588, n38589, n38590, n38591,
         n38592, n38593, n38594, n38595, n38596, n38597, n38598, n38599,
         n38600, n38601, n38602, n38603, n38604, n38605, n38606, n38607,
         n38608, n38609, n38610, n38611, n38612, n38613, n38614, n38615,
         n38616, n38617, n38618, n38619, n38620, n38621, n38622, n38623,
         n38624, n38625, n38626, n38627, n38628, n38629, n38630, n38631,
         n38632, n38633, n38634, n38635, n38636, n38637, n38638, n38639,
         n38640, n38641, n38642, n38643, n38644, n38645, n38646, n38647,
         n38648, n38649, n38650, n38651, n38652, n38653, n38654, n38655,
         n38656, n38657, n38658, n38659, n38660, n38661, n38662, n38663,
         n38664, n38665, n38666, n38667, n38668, n38669, n38670, n38671,
         n38672, n38673, n38674, n38675, n38676, n38677, n38678, n38679,
         n38680, n38681, n38682, n38683, n38684, n38685, n38686, n38687,
         n38688, n38689, n38690, n38691, n38692, n38693, n38694, n38695,
         n38696, n38697, n38698, n38699, n38700, n38701, n38702, n38703,
         n38704, n38705, n38706, n38707, n38708, n38709, n38710, n38711,
         n38712, n38713, n38714, n38715, n38716, n38717, n38718, n38719,
         n38720, n38721, n38722, n38723, n38724, n38725, n38726, n38727,
         n38728, n38729, n38730, n38731, n38732, n38733, n38734, n38735,
         n38736, n38737, n38738, n38739, n38740, n38741, n38742, n38743,
         n38744, n38745, n38746, n38747, n38748, n38749, n38750, n38751,
         n38752, n38753, n38754, n38755, n38756, n38757, n38758, n38759,
         n38760, n38761, n38762, n38763, n38764, n38765, n38766, n38767,
         n38768, n38769, n38770, n38771, n38772, n38773, n38774, n38775,
         n38776, n38777, n38778, n38779, n38780, n38781, n38782, n38783,
         n38784, n38785, n38786, n38787, n38788, n38789, n38790, n38791,
         n38792, n38793, n38794, n38795, n38796, n38797, n38798, n38799,
         n38800, n38801, n38802, n38803, n38804, n38805, n38806, n38807,
         n38808, n38809, n38810, n38811, n38812, n38813, n38814, n38815,
         n38816, n38817, n38818, n38819, n38820, n38821, n38822, n38823,
         n38824, n38825, n38826, n38827, n38828, n38829, n38830, n38831,
         n38832, n38833, n38834, n38835, n38836, n38837, n38838, n38839,
         n38840, n38841, n38842, n38843, n38844, n38845, n38846, n38847,
         n38848, n38849, n38850, n38851, n38852, n38853, n38854, n38855,
         n38856, n38857, n38858, n38859, n38860, n38861, n38862, n38863,
         n38864, n38865, n38866, n38867, n38868, n38869, n38870, n38871,
         n38872, n38873, n38874, n38875, n38876, n38877, n38878, n38879,
         n38880, n38881, n38882, n38883, n38884, n38885, n38886, n38887,
         n38888, n38889, n38890, n38891, n38892, n38893, n38894, n38895,
         n38896, n38897, n38898, n38899, n38900, n38901, n38902, n38903,
         n38904, n38905, n38906, n38907, n38908, n38909, n38910, n38911,
         n38912, n38913, n38914, n38915, n38916, n38917, n38918, n38919,
         n38920, n38921, n38922, n38923, n38924, n38925, n38926, n38927,
         n38928, n38929, n38930, n38931, n38932, n38933, n38934, n38935,
         n38936, n38937, n38938, n38939, n38940, n38941, n38942, n38943,
         n38944, n38945, n38946, n38947, n38948, n38949, n38950, n38951,
         n38952, n38953, n38954, n38955, n38956, n38957, n38958, n38959,
         n38960, n38961, n38962, n38963, n38964, n38965, n38966, n38967,
         n38968, n38969, n38970, n38971, n38972, n38973, n38974, n38975,
         n38976, n38977, n38978, n38979, n38980, n38981, n38982, n38983,
         n38984, n38985, n38986, n38987, n38988, n38989, n38990, n38991,
         n38992, n38993, n38994, n38995, n38996, n38997, n38998, n38999,
         n39000, n39001, n39002, n39003, n39004, n39005, n39006, n39007,
         n39008, n39009, n39010, n39011, n39012, n39013, n39014, n39015,
         n39016, n39017, n39018, n39019, n39020, n39021, n39022, n39023,
         n39024, n39025, n39026, n39027, n39028, n39029, n39030, n39031,
         n39032, n39033, n39034, n39035, n39036, n39037, n39038, n39039,
         n39040, n39041, n39042, n39043, n39044, n39045, n39046, n39047,
         n39048, n39049, n39050, n39051, n39052, n39053, n39054, n39055,
         n39056, n39057, n39058, n39059, n39060, n39061, n39062, n39063,
         n39064, n39065, n39066, n39067, n39068, n39069, n39070, n39071,
         n39072, n39073, n39074, n39075, n39076, n39077, n39078, n39079,
         n39080, n39081, n39082, n39083, n39084, n39085, n39086, n39087,
         n39088, n39089, n39090, n39091, n39092, n39093, n39094, n39095,
         n39096, n39097, n39098, n39099, n39100, n39101, n39102, n39103,
         n39104, n39105, n39106, n39107, n39108, n39109, n39110, n39111,
         n39112, n39113, n39114, n39115, n39116, n39117, n39118, n39119,
         n39120, n39121, n39122, n39123, n39124, n39125, n39126, n39127,
         n39128, n39129, n39130, n39131, n39132, n39133, n39134, n39135,
         n39136, n39137, n39138, n39139, n39140, n39141, n39142, n39143,
         n39144, n39145, n39146, n39147, n39148, n39149, n39150, n39151,
         n39152, n39153, n39154, n39155, n39156, n39157, n39158, n39159,
         n39160, n39161, n39162, n39163, n39164, n39165, n39166, n39167,
         n39168, n39169, n39170, n39171, n39172, n39173, n39174, n39175,
         n39176, n39177, n39178, n39179, n39180, n39181, n39182, n39183,
         n39184, n39185, n39186, n39187, n39188, n39189, n39190, n39191,
         n39192, n39193, n39194, n39195, n39196, n39197, n39198, n39199,
         n39200, n39201, n39202, n39203, n39204, n39205, n39206, n39207,
         n39208, n39209, n39210, n39211, n39212, n39213, n39214, n39215,
         n39216, n39217, n39218, n39219, n39220, n39221, n39222, n39223,
         n39224, n39225, n39226, n39227, n39228, n39229, n39230, n39231,
         n39232, n39233, n39234, n39235, n39236, n39237, n39238, n39239,
         n39240, n39241, n39242, n39243, n39244, n39245, n39246, n39247,
         n39248, n39249, n39250, n39251, n39252, n39253, n39254, n39255,
         n39256, n39257, n39258, n39259, n39260, n39261, n39262, n39263,
         n39264, n39265, n39266, n39267, n39268, n39269, n39270, n39271,
         n39272, n39273, n39274, n39275, n39276, n39277, n39278, n39279,
         n39280, n39281, n39282, n39283, n39284, n39285, n39286, n39287,
         n39288, n39289, n39290, n39291, n39292, n39293, n39294, n39295,
         n39296, n39297, n39298, n39299, n39300, n39301, n39302, n39303,
         n39304, n39305, n39306, n39307, n39308, n39309, n39310, n39311,
         n39312, n39313, n39314, n39315, n39316, n39317, n39318, n39319,
         n39320, n39321, n39322, n39323, n39324, n39325, n39326, n39327,
         n39328, n39329, n39330, n39331, n39332, n39333, n39334, n39335,
         n39336, n39337, n39338, n39339, n39340, n39341, n39342, n39343,
         n39344, n39345, n39346, n39347, n39348, n39349, n39350, n39351,
         n39352, n39353, n39354, n39355, n39356, n39357, n39358, n39359,
         n39360, n39361, n39362, n39363, n39364, n39365, n39366, n39367,
         n39368, n39369, n39370, n39371, n39372, n39373, n39374, n39375,
         n39376, n39377, n39378, n39379, n39380, n39381, n39382, n39383,
         n39384, n39385, n39386, n39387, n39388, n39389, n39390, n39391,
         n39392, n39393, n39394, n39395, n39396, n39397, n39398, n39399,
         n39400, n39401, n39402, n39403, n39404, n39405, n39406, n39407,
         n39408, n39409, n39410, n39411, n39412, n39413, n39414, n39415,
         n39416, n39417, n39418, n39419, n39420, n39421, n39422, n39423,
         n39424, n39425, n39426, n39427, n39428, n39429, n39430, n39431,
         n39432, n39433, n39434, n39435, n39436, n39437, n39438, n39439,
         n39440, n39441, n39442, n39443, n39444, n39445, n39446, n39447,
         n39448, n39449, n39450, n39451, n39452, n39453, n39454, n39455,
         n39456, n39457, n39458, n39459, n39460, n39461, n39462, n39463,
         n39464, n39465, n39466, n39467, n39468, n39469, n39470, n39471,
         n39472, n39473, n39474, n39475, n39476, n39477, n39478, n39479,
         n39480, n39481, n39482, n39483, n39484, n39485, n39486, n39487,
         n39488, n39489, n39490, n39491, n39492, n39493, n39494, n39495,
         n39496, n39497, n39498, n39499, n39500, n39501, n39502, n39503,
         n39504, n39505, n39506, n39507, n39508, n39509, n39510, n39511,
         n39512, n39513, n39514, n39515, n39516, n39517, n39518, n39519,
         n39520, n39521, n39522, n39523, n39524, n39525, n39526, n39527,
         n39528, n39529, n39530, n39531, n39532, n39533, n39534, n39535,
         n39536, n39537, n39538, n39539, n39540, n39541, n39542, n39543,
         n39544, n39545, n39546, n39547, n39548, n39549, n39550, n39551,
         n39552, n39553, n39554, n39555, n39556, n39557, n39558, n39559,
         n39560, n39561, n39562, n39563, n39564, n39565, n39566, n39567,
         n39568, n39569, n39570, n39571, n39572, n39573, n39574, n39575,
         n39576, n39577, n39578, n39579, n39580, n39581, n39582, n39583,
         n39584, n39585, n39586, n39587, n39588, n39589, n39590, n39591,
         n39592, n39593, n39594, n39595, n39596, n39597, n39598, n39599,
         n39600, n39601, n39602, n39603, n39604, n39605, n39606, n39607,
         n39608, n39609, n39610, n39611, n39612, n39613, n39614, n39615,
         n39616, n39617, n39618, n39619, n39620, n39621, n39622, n39623,
         n39624, n39625, n39626, n39627, n39628, n39629, n39630, n39631,
         n39632, n39633, n39634, n39635, n39636, n39637, n39638, n39639,
         n39640, n39641, n39642, n39643, n39644, n39645, n39646, n39647,
         n39648, n39649, n39650, n39651, n39652, n39653, n39654, n39655,
         n39656, n39657, n39658, n39659, n39660, n39661, n39662, n39663,
         n39664, n39665, n39666, n39667, n39668, n39669, n39670, n39671,
         n39672, n39673, n39674, n39675, n39676, n39677, n39678, n39679,
         n39680, n39681, n39682, n39683, n39684, n39685, n39686, n39687,
         n39688, n39689, n39690, n39691, n39692, n39693, n39694, n39695,
         n39696, n39697, n39698, n39699, n39700, n39701, n39702, n39703,
         n39704, n39705, n39706, n39707, n39708, n39709, n39710, n39711,
         n39712, n39713, n39714, n39715, n39716, n39717, n39718, n39719,
         n39720, n39721, n39722, n39723, n39724, n39725, n39726, n39727,
         n39728, n39729, n39730, n39731, n39732, n39733, n39734, n39735,
         n39736, n39737, n39738, n39739, n39740, n39741, n39742, n39743,
         n39744, n39745, n39746, n39747, n39748, n39749, n39750, n39751,
         n39752, n39753, n39754, n39755, n39756, n39757, n39758, n39759,
         n39760, n39761, n39762, n39763, n39764, n39765, n39766, n39767,
         n39768, n39769, n39770, n39771, n39772, n39773, n39774, n39775,
         n39776, n39777, n39778, n39779, n39780, n39781, n39782, n39783,
         n39784, n39785, n39786, n39787, n39788, n39789, n39790, n39791,
         n39792, n39793, n39794, n39795, n39796, n39797, n39798, n39799,
         n39800, n39801, n39802, n39803, n39804, n39805, n39806, n39807,
         n39808, n39809, n39810, n39811, n39812, n39813, n39814, n39815,
         n39816, n39817, n39818, n39819, n39820, n39821, n39822, n39823,
         n39824, n39825, n39826, n39827, n39828, n39829, n39830, n39831,
         n39832, n39833, n39834, n39835, n39836, n39837, n39838, n39839,
         n39840, n39841, n39842, n39843, n39844, n39845, n39846, n39847,
         n39848, n39849, n39850, n39851, n39852, n39853, n39854, n39855,
         n39856, n39857, n39858, n39859, n39860, n39861, n39862, n39863,
         n39864, n39865, n39866, n39867, n39868, n39869, n39870, n39871,
         n39872, n39873, n39874, n39875, n39876, n39877, n39878, n39879,
         n39880, n39881, n39882, n39883, n39884, n39885, n39886, n39887,
         n39888, n39889, n39890, n39891, n39892, n39893, n39894, n39895,
         n39896, n39897, n39898, n39899, n39900, n39901, n39902, n39903,
         n39904, n39905, n39906, n39907, n39908, n39909, n39910, n39911,
         n39912, n39913, n39914, n39915, n39916, n39917, n39918, n39919,
         n39920, n39921, n39922, n39923, n39924, n39925, n39926, n39927,
         n39928, n39929, n39930, n39931, n39932, n39933, n39934, n39935,
         n39936, n39937, n39938, n39939, n39940, n39941, n39942, n39943,
         n39944, n39945, n39946, n39947, n39948, n39949, n39950, n39951,
         n39952, n39953, n39954, n39955, n39956, n39957, n39958, n39959,
         n39960, n39961, n39962, n39963, n39964, n39965, n39966, n39967,
         n39968, n39969, n39970, n39971, n39972, n39973, n39974, n39975,
         n39976, n39977, n39978, n39979, n39980, n39981, n39982, n39983,
         n39984, n39985, n39986, n39987, n39988, n39989, n39990, n39991,
         n39992, n39993, n39994, n39995, n39996, n39997, n39998, n39999,
         n40000, n40001, n40002, n40003, n40004, n40005, n40006, n40007,
         n40008, n40009, n40010, n40011, n40012, n40013, n40014, n40015,
         n40016, n40017, n40018, n40019, n40020, n40021, n40022, n40023,
         n40024, n40025, n40026, n40027, n40028, n40029, n40030, n40031,
         n40032, n40033, n40034, n40035, n40036, n40037, n40038, n40039,
         n40040, n40041, n40042, n40043, n40044, n40045, n40046, n40047,
         n40048, n40049, n40050, n40051, n40052, n40053, n40054, n40055,
         n40056, n40057, n40058, n40059, n40060, n40061, n40062, n40063,
         n40064, n40065, n40066, n40067, n40068, n40069, n40070, n40071,
         n40072, n40073, n40074, n40075, n40076, n40077, n40078, n40079,
         n40080, n40081, n40082, n40083, n40084, n40085, n40086, n40087,
         n40088, n40089, n40090, n40091, n40092, n40093, n40094, n40095,
         n40096, n40097, n40098, n40099, n40100, n40101, n40102, n40103,
         n40104, n40105, n40106, n40107, n40108, n40109, n40110, n40111,
         n40112, n40113, n40114, n40115, n40116, n40117, n40118, n40119,
         n40120, n40121, n40122, n40123, n40124, n40125, n40126, n40127,
         n40128, n40129, n40130, n40131, n40132, n40133, n40134, n40135,
         n40136, n40137, n40138, n40139, n40140, n40141, n40142, n40143,
         n40144, n40145, n40146, n40147, n40148, n40149, n40150, n40151,
         n40152, n40153, n40154, n40155, n40156, n40157, n40158, n40159,
         n40160, n40161, n40162, n40163, n40164, n40165, n40166, n40167,
         n40168, n40169, n40170, n40171, n40172, n40173, n40174, n40175,
         n40176, n40177, n40178, n40179, n40180, n40181, n40182, n40183,
         n40184, n40185, n40186, n40187, n40188, n40189, n40190, n40191,
         n40192, n40193, n40194, n40195, n40196, n40197, n40198, n40199,
         n40200, n40201, n40202, n40203, n40204, n40205, n40206, n40207,
         n40208, n40209, n40210, n40211, n40212, n40213, n40214, n40215,
         n40216, n40217, n40218, n40219, n40220, n40221, n40222, n40223,
         n40224, n40225, n40226, n40227, n40228, n40229, n40230, n40231,
         n40232, n40233, n40234, n40235, n40236, n40237, n40238, n40239,
         n40240, n40241, n40242, n40243, n40244, n40245, n40246, n40247,
         n40248, n40249, n40250, n40251, n40252, n40253, n40254, n40255,
         n40256, n40257, n40258, n40259, n40260, n40261, n40262, n40263,
         n40264, n40265, n40266, n40267, n40268, n40269, n40270, n40271,
         n40272, n40273, n40274, n40275, n40276, n40277, n40278, n40279,
         n40280, n40281, n40282, n40283, n40284, n40285, n40286, n40287,
         n40288, n40289, n40290, n40291, n40292, n40293, n40294, n40295,
         n40296, n40297, n40298, n40299, n40300, n40301, n40302, n40303,
         n40304, n40305, n40306, n40307, n40308, n40309, n40310, n40311,
         n40312, n40313, n40314, n40315, n40316, n40317, n40318, n40319,
         n40320, n40321, n40322, n40323, n40324, n40325, n40326, n40327,
         n40328, n40329, n40330, n40331, n40332, n40333, n40334, n40335,
         n40336, n40337, n40338, n40339, n40340, n40341, n40342, n40343,
         n40344, n40345, n40346, n40347, n40348, n40349, n40350, n40351,
         n40352, n40353, n40354, n40355, n40356, n40357, n40358, n40359,
         n40360, n40361, n40362, n40363, n40364, n40365, n40366, n40367,
         n40368, n40369, n40370, n40371, n40372, n40373, n40374, n40375,
         n40376, n40377, n40378, n40379, n40380, n40381, n40382, n40383,
         n40384, n40385, n40386, n40387, n40388, n40389, n40390, n40391,
         n40392, n40393, n40394, n40395, n40396, n40397, n40398, n40399,
         n40400, n40401, n40402, n40403, n40404, n40405, n40406, n40407,
         n40408, n40409, n40410, n40411, n40412, n40413, n40414, n40415,
         n40416, n40417, n40418, n40419, n40420, n40421, n40422, n40423,
         n40424, n40425, n40426, n40427, n40428, n40429, n40430, n40431,
         n40432, n40433, n40434, n40435, n40436, n40437, n40438, n40439,
         n40440, n40441, n40442, n40443, n40444, n40445, n40446, n40447,
         n40448, n40449, n40450, n40451, n40452, n40453, n40454, n40455,
         n40456, n40457, n40458, n40459, n40460, n40461, n40462, n40463,
         n40464, n40465, n40466, n40467, n40468, n40469, n40470, n40471,
         n40472, n40473, n40474, n40475, n40476, n40477, n40478, n40479,
         n40480, n40481, n40482, n40483, n40484, n40485, n40486, n40487,
         n40488, n40489, n40490, n40491, n40492, n40493, n40494, n40495,
         n40496, n40497, n40498, n40499, n40500, n40501, n40502, n40503,
         n40504, n40505, n40506, n40507, n40508, n40509, n40510, n40511,
         n40512, n40513, n40514, n40515, n40516, n40517, n40518, n40519,
         n40520, n40521, n40522, n40523, n40524, n40525, n40526, n40527,
         n40528, n40529, n40530, n40531, n40532, n40533, n40534, n40535,
         n40536, n40537, n40538, n40539, n40540, n40541, n40542, n40543,
         n40544, n40545, n40546, n40547, n40548, n40549, n40550, n40551,
         n40552, n40553, n40554, n40555, n40556, n40557, n40558, n40559,
         n40560, n40561, n40562, n40563, n40564, n40565, n40566, n40567,
         n40568, n40569, n40570, n40571, n40572, n40573, n40574, n40575,
         n40576, n40577, n40578, n40579, n40580, n40581, n40582, n40583,
         n40584, n40585, n40586, n40587, n40588, n40589, n40590, n40591,
         n40592, n40593, n40594, n40595, n40596, n40597, n40598, n40599,
         n40600, n40601, n40602, n40603, n40604, n40605, n40606, n40607,
         n40608, n40609, n40610, n40611, n40612, n40613, n40614, n40615,
         n40616, n40617, n40618, n40619, n40620, n40621, n40622, n40623,
         n40624, n40625, n40626, n40627, n40628, n40629, n40630, n40631,
         n40632, n40633, n40634, n40635, n40636, n40637, n40638, n40639,
         n40640, n40641, n40642, n40643, n40644, n40645, n40646, n40647,
         n40648, n40649, n40650, n40651, n40652, n40653, n40654, n40655,
         n40656, n40657, n40658, n40659, n40660, n40661, n40662, n40663,
         n40664, n40665, n40666, n40667, n40668, n40669, n40670, n40671,
         n40672, n40673, n40674, n40675, n40676, n40677, n40678, n40679,
         n40680, n40681, n40682, n40683, n40684, n40685, n40686, n40687,
         n40688, n40689, n40690, n40691, n40692, n40693, n40694, n40695,
         n40696, n40697, n40698, n40699, n40700, n40701, n40702, n40703,
         n40704, n40705, n40706, n40707, n40708, n40709, n40710, n40711,
         n40712, n40713, n40714, n40715, n40716, n40717, n40718, n40719,
         n40720, n40721, n40722, n40723, n40724, n40725, n40726, n40727,
         n40728, n40729, n40730, n40731, n40732, n40733, n40734, n40735,
         n40736, n40737, n40738, n40739, n40740, n40741, n40742, n40743,
         n40744, n40745, n40746, n40747, n40748, n40749, n40750, n40751,
         n40752, n40753, n40754, n40755, n40756, n40757, n40758, n40759,
         n40760, n40761, n40762, n40763, n40764, n40765, n40766, n40767,
         n40768, n40769, n40770, n40771, n40772, n40773, n40774, n40775,
         n40776, n40777, n40778, n40779, n40780, n40781, n40782, n40783,
         n40784, n40785, n40786, n40787, n40788, n40789, n40790, n40791,
         n40792, n40793, n40794, n40795, n40796, n40797, n40798, n40799,
         n40800, n40801, n40802, n40803, n40804, n40805, n40806, n40807,
         n40808, n40809, n40810, n40811, n40812, n40813, n40814, n40815,
         n40816, n40817, n40818, n40819, n40820, n40821, n40822, n40823,
         n40824, n40825, n40826, n40827, n40828, n40829, n40830, n40831,
         n40832, n40833, n40834, n40835, n40836, n40837, n40838, n40839,
         n40840, n40841, n40842, n40843, n40844, n40845, n40846, n40847,
         n40848, n40849, n40850, n40851, n40852, n40853, n40854, n40855,
         n40856, n40857, n40858, n40859, n40860, n40861, n40862, n40863,
         n40864, n40865, n40866, n40867, n40868, n40869, n40870, n40871,
         n40872, n40873, n40874, n40875, n40876, n40877, n40878, n40879,
         n40880, n40881, n40882, n40883, n40884, n40885, n40886, n40887,
         n40888, n40889, n40890, n40891, n40892, n40893, n40894, n40895,
         n40896, n40897, n40898, n40899, n40900, n40901, n40902, n40903,
         n40904, n40905, n40906, n40907, n40908, n40909, n40910, n40911,
         n40912, n40913, n40914, n40915, n40916, n40917, n40918, n40919,
         n40920, n40921, n40922, n40923, n40924, n40925, n40926, n40927,
         n40928, n40929, n40930, n40931, n40932, n40933, n40934, n40935,
         n40936, n40937, n40938, n40939, n40940, n40941, n40942, n40943,
         n40944, n40945, n40946, n40947, n40948, n40949, n40950, n40951,
         n40952, n40953, n40954, n40955, n40956, n40957, n40958, n40959,
         n40960, n40961, n40962, n40963, n40964, n40965, n40966, n40967,
         n40968, n40969, n40970, n40971, n40972, n40973, n40974, n40975,
         n40976, n40977, n40978, n40979, n40980, n40981, n40982, n40983,
         n40984, n40985, n40986, n40987, n40988, n40989, n40990, n40991,
         n40992, n40993, n40994, n40995, n40996, n40997, n40998, n40999,
         n41000, n41001, n41002, n41003, n41004, n41005, n41006, n41007,
         n41008, n41009, n41010, n41011, n41012, n41013, n41014, n41015,
         n41016, n41017, n41018, n41019, n41020, n41021, n41022, n41023,
         n41024, n41025, n41026, n41027, n41028, n41029, n41030, n41031,
         n41032, n41033, n41034, n41035, n41036, n41037, n41038, n41039,
         n41040, n41041, n41042, n41043, n41044, n41045, n41046, n41047,
         n41048, n41049, n41050, n41051, n41052, n41053, n41054, n41055,
         n41056, n41057, n41058, n41059, n41060, n41061, n41062, n41063,
         n41064, n41065, n41066, n41067, n41068, n41069, n41070, n41071,
         n41072, n41073, n41074, n41075, n41076, n41077, n41078, n41079,
         n41080, n41081, n41082, n41083, n41084, n41085, n41086, n41087,
         n41088, n41089, n41090, n41091, n41092, n41093, n41094, n41095,
         n41096, n41097, n41098, n41099, n41100, n41101, n41102, n41103,
         n41104, n41105, n41106, n41107, n41108, n41109, n41110, n41111,
         n41112, n41113, n41114, n41115, n41116, n41117, n41118, n41119,
         n41120, n41121, n41122, n41123, n41124, n41125, n41126, n41127,
         n41128, n41129, n41130, n41131, n41132, n41133, n41134, n41135,
         n41136, n41137, n41138, n41139, n41140, n41141, n41142, n41143,
         n41144, n41145, n41146, n41147, n41148, n41149, n41150, n41151,
         n41152, n41153, n41154, n41155, n41156, n41157, n41158, n41159,
         n41160, n41161, n41162, n41163, n41164, n41165, n41166, n41167,
         n41168, n41169, n41170, n41171, n41172, n41173, n41174, n41175,
         n41176, n41177, n41178, n41179, n41180, n41181, n41182, n41183,
         n41184, n41185, n41186, n41187, n41188, n41189, n41190, n41191,
         n41192, n41193, n41194, n41195, n41196, n41197, n41198, n41199,
         n41200, n41201, n41202, n41203, n41204, n41205, n41206, n41207,
         n41208, n41209, n41210, n41211, n41212, n41213, n41214, n41215,
         n41216, n41217, n41218, n41219, n41220, n41221, n41222, n41223,
         n41224, n41225, n41226, n41227, n41228, n41229, n41230, n41231,
         n41232, n41233, n41234, n41235, n41236, n41237, n41238, n41239,
         n41240, n41241, n41242, n41243, n41244, n41245, n41246, n41247,
         n41248, n41249, n41250, n41251, n41252, n41253, n41254, n41255,
         n41256, n41257, n41258, n41259, n41260, n41261, n41262, n41263,
         n41264, n41265, n41266, n41267, n41268, n41269, n41270, n41271,
         n41272, n41273, n41274, n41275, n41276, n41277, n41278, n41279,
         n41280, n41281, n41282, n41283, n41284, n41285, n41286, n41287,
         n41288, n41289, n41290, n41291, n41292, n41293, n41294, n41295,
         n41296, n41297, n41298, n41299, n41300, n41301, n41302, n41303,
         n41304, n41305, n41306, n41307, n41308, n41309, n41310, n41311,
         n41312, n41313, n41314, n41315, n41316, n41317, n41318, n41319,
         n41320, n41321, n41322, n41323, n41324, n41325, n41326, n41327,
         n41328, n41329, n41330, n41331, n41332, n41333, n41334, n41335,
         n41336, n41337, n41338, n41339, n41340, n41341, n41342, n41343,
         n41344, n41345, n41346, n41347, n41348, n41349, n41350, n41351,
         n41352, n41353, n41354, n41355, n41356, n41357, n41358, n41359,
         n41360, n41361, n41362, n41363, n41364, n41365, n41366, n41367,
         n41368, n41369, n41370, n41371, n41372, n41373, n41374, n41375,
         n41376, n41377, n41378, n41379, n41380, n41381, n41382, n41383,
         n41384, n41385, n41386, n41387, n41388, n41389, n41390, n41391,
         n41392, n41393, n41394, n41395, n41396, n41397, n41398, n41399,
         n41400, n41401, n41402, n41403, n41404, n41405, n41406, n41407,
         n41408, n41409, n41410, n41411, n41412, n41413, n41414, n41415,
         n41416, n41417, n41418, n41419, n41420, n41421, n41422, n41423,
         n41424, n41425, n41426, n41427, n41428, n41429, n41430, n41431,
         n41432, n41433, n41434, n41435, n41436, n41437, n41438, n41439,
         n41440, n41441, n41442, n41443, n41444, n41445, n41446, n41447,
         n41448, n41449, n41450, n41451, n41452, n41453, n41454, n41455,
         n41456, n41457, n41458, n41459, n41460, n41461, n41462, n41463,
         n41464, n41465, n41466, n41467, n41468, n41469, n41470, n41471,
         n41472, n41473, n41474, n41475, n41476, n41477, n41478, n41479,
         n41480, n41481, n41482, n41483, n41484, n41485, n41486, n41487,
         n41488, n41489, n41490, n41491, n41492, n41493, n41494, n41495,
         n41496, n41497, n41498, n41499, n41500, n41501, n41502, n41503,
         n41504, n41505, n41506, n41507, n41508, n41509, n41510, n41511,
         n41512, n41513, n41514, n41515, n41516, n41517, n41518, n41519,
         n41520, n41521, n41522, n41523, n41524, n41525, n41526, n41527,
         n41528, n41529, n41530, n41531, n41532, n41533, n41534, n41535,
         n41536, n41537, n41538, n41539, n41540, n41541, n41542, n41543,
         n41544, n41545, n41546, n41547, n41548, n41549, n41550, n41551,
         n41552, n41553, n41554, n41555, n41556, n41557, n41558, n41559,
         n41560, n41561, n41562, n41563, n41564, n41565, n41566, n41567,
         n41568, n41569, n41570, n41571, n41572, n41573, n41574, n41575,
         n41576, n41577, n41578, n41579, n41580, n41581, n41582, n41583,
         n41584, n41585, n41586, n41587, n41588, n41589, n41590, n41591,
         n41592, n41593, n41594, n41595, n41596, n41597, n41598, n41599,
         n41600, n41601, n41602, n41603, n41604, n41605, n41606, n41607,
         n41608, n41609, n41610, n41611, n41612, n41613, n41614, n41615,
         n41616, n41617, n41618, n41619, n41620, n41621, n41622, n41623,
         n41624, n41625, n41626, n41627, n41628, n41629, n41630, n41631,
         n41632, n41633, n41634, n41635, n41636, n41637, n41638, n41639,
         n41640, n41641, n41642, n41643, n41644, n41645, n41646, n41647,
         n41648, n41649, n41650, n41651, n41652, n41653, n41654, n41655,
         n41656, n41657, n41658, n41659, n41660, n41661, n41662, n41663,
         n41664, n41665, n41666, n41667, n41668, n41669, n41670, n41671,
         n41672, n41673, n41674, n41675, n41676, n41677, n41678, n41679,
         n41680, n41681, n41682, n41683, n41684, n41685, n41686, n41687,
         n41688, n41689, n41690, n41691, n41692, n41693, n41694, n41695,
         n41696, n41697, n41698, n41699, n41700, n41701, n41702, n41703,
         n41704, n41705, n41706, n41707, n41708, n41709, n41710, n41711,
         n41712, n41713, n41714, n41715, n41716, n41717, n41718, n41719,
         n41720, n41721, n41722, n41723, n41724, n41725, n41726, n41727,
         n41728, n41729, n41730, n41731, n41732, n41733, n41734, n41735,
         n41736, n41737, n41738, n41739, n41740, n41741, n41742, n41743,
         n41744, n41745, n41746, n41747, n41748, n41749, n41750, n41751,
         n41752, n41753, n41754, n41755, n41756, n41757, n41758, n41759,
         n41760, n41761, n41762, n41763, n41764, n41765, n41766, n41767,
         n41768, n41769, n41770, n41771, n41772, n41773, n41774, n41775,
         n41776, n41777, n41778, n41779, n41780, n41781, n41782, n41783,
         n41784, n41785, n41786, n41787, n41788, n41789, n41790, n41791,
         n41792, n41793, n41794, n41795, n41796, n41797, n41798, n41799,
         n41800, n41801, n41802, n41803, n41804, n41805, n41806, n41807,
         n41808, n41809, n41810, n41811, n41812, n41813, n41814, n41815,
         n41816, n41817, n41818, n41819, n41820, n41821, n41822, n41823,
         n41824, n41825, n41826, n41827, n41828, n41829, n41830, n41831,
         n41832, n41833, n41834, n41835, n41836, n41837, n41838, n41839,
         n41840, n41841, n41842, n41843, n41844, n41845, n41846, n41847,
         n41848, n41849, n41850, n41851, n41852, n41853, n41854, n41855,
         n41856, n41857, n41858, n41859, n41860, n41861, n41862, n41863,
         n41864, n41865, n41866, n41867, n41868, n41869, n41870, n41871,
         n41872, n41873, n41874, n41875, n41876, n41877, n41878, n41879,
         n41880, n41881, n41882, n41883, n41884, n41885, n41886, n41887,
         n41888, n41889, n41890, n41891, n41892, n41893, n41894, n41895,
         n41896, n41897, n41898, n41899, n41900, n41901, n41902, n41903,
         n41904, n41905, n41906, n41907, n41908, n41909, n41910, n41911,
         n41912, n41913, n41914, n41915, n41916, n41917, n41918, n41919,
         n41920, n41921, n41922, n41923, n41924, n41925, n41926, n41927,
         n41928, n41929, n41930, n41931, n41932, n41933, n41934, n41935,
         n41936, n41937, n41938, n41939, n41940, n41941, n41942, n41943,
         n41944, n41945, n41946, n41947, n41948, n41949, n41950, n41951,
         n41952, n41953, n41954, n41955, n41956, n41957, n41958, n41959,
         n41960, n41961, n41962, n41963, n41964, n41965, n41966, n41967,
         n41968, n41969, n41970, n41971, n41972, n41973, n41974, n41975,
         n41976, n41977, n41978, n41979, n41980, n41981, n41982, n41983,
         n41984, n41985, n41986, n41987, n41988, n41989;
  wire   [1023:0] start_in;
  wire   [1023:0] ein;
  wire   [1023:0] mod_mult_o;
  wire   [1023:0] creg;
  wire   [1023:0] ereg_next;

  DFF \start_reg_reg[0]  ( .D(start_in[1023]), .CLK(clk), .RST(rst), .I(1'b1), 
        .Q(start_in[0]) );
  DFF \start_reg_reg[1]  ( .D(start_in[0]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[1]) );
  DFF \start_reg_reg[2]  ( .D(start_in[1]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[2]) );
  DFF \start_reg_reg[3]  ( .D(start_in[2]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[3]) );
  DFF \start_reg_reg[4]  ( .D(start_in[3]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[4]) );
  DFF \start_reg_reg[5]  ( .D(start_in[4]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[5]) );
  DFF \start_reg_reg[6]  ( .D(start_in[5]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[6]) );
  DFF \start_reg_reg[7]  ( .D(start_in[6]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[7]) );
  DFF \start_reg_reg[8]  ( .D(start_in[7]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[8]) );
  DFF \start_reg_reg[9]  ( .D(start_in[8]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[9]) );
  DFF \start_reg_reg[10]  ( .D(start_in[9]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[10]) );
  DFF \start_reg_reg[11]  ( .D(start_in[10]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[11]) );
  DFF \start_reg_reg[12]  ( .D(start_in[11]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[12]) );
  DFF \start_reg_reg[13]  ( .D(start_in[12]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[13]) );
  DFF \start_reg_reg[14]  ( .D(start_in[13]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[14]) );
  DFF \start_reg_reg[15]  ( .D(start_in[14]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[15]) );
  DFF \start_reg_reg[16]  ( .D(start_in[15]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[16]) );
  DFF \start_reg_reg[17]  ( .D(start_in[16]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[17]) );
  DFF \start_reg_reg[18]  ( .D(start_in[17]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[18]) );
  DFF \start_reg_reg[19]  ( .D(start_in[18]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[19]) );
  DFF \start_reg_reg[20]  ( .D(start_in[19]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[20]) );
  DFF \start_reg_reg[21]  ( .D(start_in[20]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[21]) );
  DFF \start_reg_reg[22]  ( .D(start_in[21]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[22]) );
  DFF \start_reg_reg[23]  ( .D(start_in[22]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[23]) );
  DFF \start_reg_reg[24]  ( .D(start_in[23]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[24]) );
  DFF \start_reg_reg[25]  ( .D(start_in[24]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[25]) );
  DFF \start_reg_reg[26]  ( .D(start_in[25]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[26]) );
  DFF \start_reg_reg[27]  ( .D(start_in[26]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[27]) );
  DFF \start_reg_reg[28]  ( .D(start_in[27]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[28]) );
  DFF \start_reg_reg[29]  ( .D(start_in[28]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[29]) );
  DFF \start_reg_reg[30]  ( .D(start_in[29]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[30]) );
  DFF \start_reg_reg[31]  ( .D(start_in[30]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[31]) );
  DFF \start_reg_reg[32]  ( .D(start_in[31]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[32]) );
  DFF \start_reg_reg[33]  ( .D(start_in[32]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[33]) );
  DFF \start_reg_reg[34]  ( .D(start_in[33]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[34]) );
  DFF \start_reg_reg[35]  ( .D(start_in[34]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[35]) );
  DFF \start_reg_reg[36]  ( .D(start_in[35]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[36]) );
  DFF \start_reg_reg[37]  ( .D(start_in[36]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[37]) );
  DFF \start_reg_reg[38]  ( .D(start_in[37]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[38]) );
  DFF \start_reg_reg[39]  ( .D(start_in[38]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[39]) );
  DFF \start_reg_reg[40]  ( .D(start_in[39]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[40]) );
  DFF \start_reg_reg[41]  ( .D(start_in[40]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[41]) );
  DFF \start_reg_reg[42]  ( .D(start_in[41]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[42]) );
  DFF \start_reg_reg[43]  ( .D(start_in[42]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[43]) );
  DFF \start_reg_reg[44]  ( .D(start_in[43]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[44]) );
  DFF \start_reg_reg[45]  ( .D(start_in[44]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[45]) );
  DFF \start_reg_reg[46]  ( .D(start_in[45]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[46]) );
  DFF \start_reg_reg[47]  ( .D(start_in[46]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[47]) );
  DFF \start_reg_reg[48]  ( .D(start_in[47]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[48]) );
  DFF \start_reg_reg[49]  ( .D(start_in[48]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[49]) );
  DFF \start_reg_reg[50]  ( .D(start_in[49]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[50]) );
  DFF \start_reg_reg[51]  ( .D(start_in[50]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[51]) );
  DFF \start_reg_reg[52]  ( .D(start_in[51]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[52]) );
  DFF \start_reg_reg[53]  ( .D(start_in[52]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[53]) );
  DFF \start_reg_reg[54]  ( .D(start_in[53]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[54]) );
  DFF \start_reg_reg[55]  ( .D(start_in[54]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[55]) );
  DFF \start_reg_reg[56]  ( .D(start_in[55]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[56]) );
  DFF \start_reg_reg[57]  ( .D(start_in[56]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[57]) );
  DFF \start_reg_reg[58]  ( .D(start_in[57]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[58]) );
  DFF \start_reg_reg[59]  ( .D(start_in[58]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[59]) );
  DFF \start_reg_reg[60]  ( .D(start_in[59]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[60]) );
  DFF \start_reg_reg[61]  ( .D(start_in[60]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[61]) );
  DFF \start_reg_reg[62]  ( .D(start_in[61]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[62]) );
  DFF \start_reg_reg[63]  ( .D(start_in[62]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[63]) );
  DFF \start_reg_reg[64]  ( .D(start_in[63]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[64]) );
  DFF \start_reg_reg[65]  ( .D(start_in[64]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[65]) );
  DFF \start_reg_reg[66]  ( .D(start_in[65]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[66]) );
  DFF \start_reg_reg[67]  ( .D(start_in[66]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[67]) );
  DFF \start_reg_reg[68]  ( .D(start_in[67]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[68]) );
  DFF \start_reg_reg[69]  ( .D(start_in[68]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[69]) );
  DFF \start_reg_reg[70]  ( .D(start_in[69]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[70]) );
  DFF \start_reg_reg[71]  ( .D(start_in[70]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[71]) );
  DFF \start_reg_reg[72]  ( .D(start_in[71]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[72]) );
  DFF \start_reg_reg[73]  ( .D(start_in[72]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[73]) );
  DFF \start_reg_reg[74]  ( .D(start_in[73]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[74]) );
  DFF \start_reg_reg[75]  ( .D(start_in[74]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[75]) );
  DFF \start_reg_reg[76]  ( .D(start_in[75]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[76]) );
  DFF \start_reg_reg[77]  ( .D(start_in[76]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[77]) );
  DFF \start_reg_reg[78]  ( .D(start_in[77]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[78]) );
  DFF \start_reg_reg[79]  ( .D(start_in[78]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[79]) );
  DFF \start_reg_reg[80]  ( .D(start_in[79]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[80]) );
  DFF \start_reg_reg[81]  ( .D(start_in[80]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[81]) );
  DFF \start_reg_reg[82]  ( .D(start_in[81]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[82]) );
  DFF \start_reg_reg[83]  ( .D(start_in[82]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[83]) );
  DFF \start_reg_reg[84]  ( .D(start_in[83]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[84]) );
  DFF \start_reg_reg[85]  ( .D(start_in[84]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[85]) );
  DFF \start_reg_reg[86]  ( .D(start_in[85]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[86]) );
  DFF \start_reg_reg[87]  ( .D(start_in[86]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[87]) );
  DFF \start_reg_reg[88]  ( .D(start_in[87]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[88]) );
  DFF \start_reg_reg[89]  ( .D(start_in[88]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[89]) );
  DFF \start_reg_reg[90]  ( .D(start_in[89]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[90]) );
  DFF \start_reg_reg[91]  ( .D(start_in[90]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[91]) );
  DFF \start_reg_reg[92]  ( .D(start_in[91]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[92]) );
  DFF \start_reg_reg[93]  ( .D(start_in[92]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[93]) );
  DFF \start_reg_reg[94]  ( .D(start_in[93]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[94]) );
  DFF \start_reg_reg[95]  ( .D(start_in[94]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[95]) );
  DFF \start_reg_reg[96]  ( .D(start_in[95]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[96]) );
  DFF \start_reg_reg[97]  ( .D(start_in[96]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[97]) );
  DFF \start_reg_reg[98]  ( .D(start_in[97]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[98]) );
  DFF \start_reg_reg[99]  ( .D(start_in[98]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[99]) );
  DFF \start_reg_reg[100]  ( .D(start_in[99]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[100]) );
  DFF \start_reg_reg[101]  ( .D(start_in[100]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[101]) );
  DFF \start_reg_reg[102]  ( .D(start_in[101]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[102]) );
  DFF \start_reg_reg[103]  ( .D(start_in[102]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[103]) );
  DFF \start_reg_reg[104]  ( .D(start_in[103]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[104]) );
  DFF \start_reg_reg[105]  ( .D(start_in[104]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[105]) );
  DFF \start_reg_reg[106]  ( .D(start_in[105]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[106]) );
  DFF \start_reg_reg[107]  ( .D(start_in[106]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[107]) );
  DFF \start_reg_reg[108]  ( .D(start_in[107]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[108]) );
  DFF \start_reg_reg[109]  ( .D(start_in[108]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[109]) );
  DFF \start_reg_reg[110]  ( .D(start_in[109]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[110]) );
  DFF \start_reg_reg[111]  ( .D(start_in[110]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[111]) );
  DFF \start_reg_reg[112]  ( .D(start_in[111]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[112]) );
  DFF \start_reg_reg[113]  ( .D(start_in[112]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[113]) );
  DFF \start_reg_reg[114]  ( .D(start_in[113]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[114]) );
  DFF \start_reg_reg[115]  ( .D(start_in[114]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[115]) );
  DFF \start_reg_reg[116]  ( .D(start_in[115]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[116]) );
  DFF \start_reg_reg[117]  ( .D(start_in[116]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[117]) );
  DFF \start_reg_reg[118]  ( .D(start_in[117]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[118]) );
  DFF \start_reg_reg[119]  ( .D(start_in[118]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[119]) );
  DFF \start_reg_reg[120]  ( .D(start_in[119]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[120]) );
  DFF \start_reg_reg[121]  ( .D(start_in[120]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[121]) );
  DFF \start_reg_reg[122]  ( .D(start_in[121]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[122]) );
  DFF \start_reg_reg[123]  ( .D(start_in[122]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[123]) );
  DFF \start_reg_reg[124]  ( .D(start_in[123]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[124]) );
  DFF \start_reg_reg[125]  ( .D(start_in[124]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[125]) );
  DFF \start_reg_reg[126]  ( .D(start_in[125]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[126]) );
  DFF \start_reg_reg[127]  ( .D(start_in[126]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[127]) );
  DFF \start_reg_reg[128]  ( .D(start_in[127]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[128]) );
  DFF \start_reg_reg[129]  ( .D(start_in[128]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[129]) );
  DFF \start_reg_reg[130]  ( .D(start_in[129]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[130]) );
  DFF \start_reg_reg[131]  ( .D(start_in[130]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[131]) );
  DFF \start_reg_reg[132]  ( .D(start_in[131]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[132]) );
  DFF \start_reg_reg[133]  ( .D(start_in[132]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[133]) );
  DFF \start_reg_reg[134]  ( .D(start_in[133]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[134]) );
  DFF \start_reg_reg[135]  ( .D(start_in[134]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[135]) );
  DFF \start_reg_reg[136]  ( .D(start_in[135]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[136]) );
  DFF \start_reg_reg[137]  ( .D(start_in[136]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[137]) );
  DFF \start_reg_reg[138]  ( .D(start_in[137]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[138]) );
  DFF \start_reg_reg[139]  ( .D(start_in[138]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[139]) );
  DFF \start_reg_reg[140]  ( .D(start_in[139]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[140]) );
  DFF \start_reg_reg[141]  ( .D(start_in[140]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[141]) );
  DFF \start_reg_reg[142]  ( .D(start_in[141]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[142]) );
  DFF \start_reg_reg[143]  ( .D(start_in[142]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[143]) );
  DFF \start_reg_reg[144]  ( .D(start_in[143]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[144]) );
  DFF \start_reg_reg[145]  ( .D(start_in[144]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[145]) );
  DFF \start_reg_reg[146]  ( .D(start_in[145]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[146]) );
  DFF \start_reg_reg[147]  ( .D(start_in[146]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[147]) );
  DFF \start_reg_reg[148]  ( .D(start_in[147]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[148]) );
  DFF \start_reg_reg[149]  ( .D(start_in[148]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[149]) );
  DFF \start_reg_reg[150]  ( .D(start_in[149]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[150]) );
  DFF \start_reg_reg[151]  ( .D(start_in[150]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[151]) );
  DFF \start_reg_reg[152]  ( .D(start_in[151]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[152]) );
  DFF \start_reg_reg[153]  ( .D(start_in[152]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[153]) );
  DFF \start_reg_reg[154]  ( .D(start_in[153]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[154]) );
  DFF \start_reg_reg[155]  ( .D(start_in[154]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[155]) );
  DFF \start_reg_reg[156]  ( .D(start_in[155]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[156]) );
  DFF \start_reg_reg[157]  ( .D(start_in[156]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[157]) );
  DFF \start_reg_reg[158]  ( .D(start_in[157]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[158]) );
  DFF \start_reg_reg[159]  ( .D(start_in[158]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[159]) );
  DFF \start_reg_reg[160]  ( .D(start_in[159]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[160]) );
  DFF \start_reg_reg[161]  ( .D(start_in[160]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[161]) );
  DFF \start_reg_reg[162]  ( .D(start_in[161]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[162]) );
  DFF \start_reg_reg[163]  ( .D(start_in[162]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[163]) );
  DFF \start_reg_reg[164]  ( .D(start_in[163]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[164]) );
  DFF \start_reg_reg[165]  ( .D(start_in[164]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[165]) );
  DFF \start_reg_reg[166]  ( .D(start_in[165]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[166]) );
  DFF \start_reg_reg[167]  ( .D(start_in[166]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[167]) );
  DFF \start_reg_reg[168]  ( .D(start_in[167]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[168]) );
  DFF \start_reg_reg[169]  ( .D(start_in[168]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[169]) );
  DFF \start_reg_reg[170]  ( .D(start_in[169]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[170]) );
  DFF \start_reg_reg[171]  ( .D(start_in[170]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[171]) );
  DFF \start_reg_reg[172]  ( .D(start_in[171]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[172]) );
  DFF \start_reg_reg[173]  ( .D(start_in[172]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[173]) );
  DFF \start_reg_reg[174]  ( .D(start_in[173]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[174]) );
  DFF \start_reg_reg[175]  ( .D(start_in[174]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[175]) );
  DFF \start_reg_reg[176]  ( .D(start_in[175]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[176]) );
  DFF \start_reg_reg[177]  ( .D(start_in[176]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[177]) );
  DFF \start_reg_reg[178]  ( .D(start_in[177]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[178]) );
  DFF \start_reg_reg[179]  ( .D(start_in[178]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[179]) );
  DFF \start_reg_reg[180]  ( .D(start_in[179]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[180]) );
  DFF \start_reg_reg[181]  ( .D(start_in[180]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[181]) );
  DFF \start_reg_reg[182]  ( .D(start_in[181]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[182]) );
  DFF \start_reg_reg[183]  ( .D(start_in[182]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[183]) );
  DFF \start_reg_reg[184]  ( .D(start_in[183]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[184]) );
  DFF \start_reg_reg[185]  ( .D(start_in[184]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[185]) );
  DFF \start_reg_reg[186]  ( .D(start_in[185]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[186]) );
  DFF \start_reg_reg[187]  ( .D(start_in[186]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[187]) );
  DFF \start_reg_reg[188]  ( .D(start_in[187]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[188]) );
  DFF \start_reg_reg[189]  ( .D(start_in[188]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[189]) );
  DFF \start_reg_reg[190]  ( .D(start_in[189]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[190]) );
  DFF \start_reg_reg[191]  ( .D(start_in[190]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[191]) );
  DFF \start_reg_reg[192]  ( .D(start_in[191]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[192]) );
  DFF \start_reg_reg[193]  ( .D(start_in[192]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[193]) );
  DFF \start_reg_reg[194]  ( .D(start_in[193]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[194]) );
  DFF \start_reg_reg[195]  ( .D(start_in[194]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[195]) );
  DFF \start_reg_reg[196]  ( .D(start_in[195]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[196]) );
  DFF \start_reg_reg[197]  ( .D(start_in[196]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[197]) );
  DFF \start_reg_reg[198]  ( .D(start_in[197]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[198]) );
  DFF \start_reg_reg[199]  ( .D(start_in[198]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[199]) );
  DFF \start_reg_reg[200]  ( .D(start_in[199]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[200]) );
  DFF \start_reg_reg[201]  ( .D(start_in[200]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[201]) );
  DFF \start_reg_reg[202]  ( .D(start_in[201]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[202]) );
  DFF \start_reg_reg[203]  ( .D(start_in[202]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[203]) );
  DFF \start_reg_reg[204]  ( .D(start_in[203]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[204]) );
  DFF \start_reg_reg[205]  ( .D(start_in[204]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[205]) );
  DFF \start_reg_reg[206]  ( .D(start_in[205]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[206]) );
  DFF \start_reg_reg[207]  ( .D(start_in[206]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[207]) );
  DFF \start_reg_reg[208]  ( .D(start_in[207]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[208]) );
  DFF \start_reg_reg[209]  ( .D(start_in[208]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[209]) );
  DFF \start_reg_reg[210]  ( .D(start_in[209]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[210]) );
  DFF \start_reg_reg[211]  ( .D(start_in[210]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[211]) );
  DFF \start_reg_reg[212]  ( .D(start_in[211]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[212]) );
  DFF \start_reg_reg[213]  ( .D(start_in[212]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[213]) );
  DFF \start_reg_reg[214]  ( .D(start_in[213]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[214]) );
  DFF \start_reg_reg[215]  ( .D(start_in[214]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[215]) );
  DFF \start_reg_reg[216]  ( .D(start_in[215]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[216]) );
  DFF \start_reg_reg[217]  ( .D(start_in[216]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[217]) );
  DFF \start_reg_reg[218]  ( .D(start_in[217]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[218]) );
  DFF \start_reg_reg[219]  ( .D(start_in[218]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[219]) );
  DFF \start_reg_reg[220]  ( .D(start_in[219]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[220]) );
  DFF \start_reg_reg[221]  ( .D(start_in[220]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[221]) );
  DFF \start_reg_reg[222]  ( .D(start_in[221]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[222]) );
  DFF \start_reg_reg[223]  ( .D(start_in[222]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[223]) );
  DFF \start_reg_reg[224]  ( .D(start_in[223]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[224]) );
  DFF \start_reg_reg[225]  ( .D(start_in[224]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[225]) );
  DFF \start_reg_reg[226]  ( .D(start_in[225]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[226]) );
  DFF \start_reg_reg[227]  ( .D(start_in[226]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[227]) );
  DFF \start_reg_reg[228]  ( .D(start_in[227]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[228]) );
  DFF \start_reg_reg[229]  ( .D(start_in[228]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[229]) );
  DFF \start_reg_reg[230]  ( .D(start_in[229]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[230]) );
  DFF \start_reg_reg[231]  ( .D(start_in[230]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[231]) );
  DFF \start_reg_reg[232]  ( .D(start_in[231]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[232]) );
  DFF \start_reg_reg[233]  ( .D(start_in[232]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[233]) );
  DFF \start_reg_reg[234]  ( .D(start_in[233]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[234]) );
  DFF \start_reg_reg[235]  ( .D(start_in[234]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[235]) );
  DFF \start_reg_reg[236]  ( .D(start_in[235]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[236]) );
  DFF \start_reg_reg[237]  ( .D(start_in[236]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[237]) );
  DFF \start_reg_reg[238]  ( .D(start_in[237]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[238]) );
  DFF \start_reg_reg[239]  ( .D(start_in[238]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[239]) );
  DFF \start_reg_reg[240]  ( .D(start_in[239]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[240]) );
  DFF \start_reg_reg[241]  ( .D(start_in[240]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[241]) );
  DFF \start_reg_reg[242]  ( .D(start_in[241]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[242]) );
  DFF \start_reg_reg[243]  ( .D(start_in[242]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[243]) );
  DFF \start_reg_reg[244]  ( .D(start_in[243]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[244]) );
  DFF \start_reg_reg[245]  ( .D(start_in[244]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[245]) );
  DFF \start_reg_reg[246]  ( .D(start_in[245]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[246]) );
  DFF \start_reg_reg[247]  ( .D(start_in[246]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[247]) );
  DFF \start_reg_reg[248]  ( .D(start_in[247]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[248]) );
  DFF \start_reg_reg[249]  ( .D(start_in[248]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[249]) );
  DFF \start_reg_reg[250]  ( .D(start_in[249]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[250]) );
  DFF \start_reg_reg[251]  ( .D(start_in[250]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[251]) );
  DFF \start_reg_reg[252]  ( .D(start_in[251]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[252]) );
  DFF \start_reg_reg[253]  ( .D(start_in[252]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[253]) );
  DFF \start_reg_reg[254]  ( .D(start_in[253]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[254]) );
  DFF \start_reg_reg[255]  ( .D(start_in[254]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[255]) );
  DFF \start_reg_reg[256]  ( .D(start_in[255]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[256]) );
  DFF \start_reg_reg[257]  ( .D(start_in[256]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[257]) );
  DFF \start_reg_reg[258]  ( .D(start_in[257]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[258]) );
  DFF \start_reg_reg[259]  ( .D(start_in[258]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[259]) );
  DFF \start_reg_reg[260]  ( .D(start_in[259]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[260]) );
  DFF \start_reg_reg[261]  ( .D(start_in[260]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[261]) );
  DFF \start_reg_reg[262]  ( .D(start_in[261]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[262]) );
  DFF \start_reg_reg[263]  ( .D(start_in[262]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[263]) );
  DFF \start_reg_reg[264]  ( .D(start_in[263]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[264]) );
  DFF \start_reg_reg[265]  ( .D(start_in[264]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[265]) );
  DFF \start_reg_reg[266]  ( .D(start_in[265]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[266]) );
  DFF \start_reg_reg[267]  ( .D(start_in[266]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[267]) );
  DFF \start_reg_reg[268]  ( .D(start_in[267]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[268]) );
  DFF \start_reg_reg[269]  ( .D(start_in[268]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[269]) );
  DFF \start_reg_reg[270]  ( .D(start_in[269]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[270]) );
  DFF \start_reg_reg[271]  ( .D(start_in[270]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[271]) );
  DFF \start_reg_reg[272]  ( .D(start_in[271]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[272]) );
  DFF \start_reg_reg[273]  ( .D(start_in[272]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[273]) );
  DFF \start_reg_reg[274]  ( .D(start_in[273]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[274]) );
  DFF \start_reg_reg[275]  ( .D(start_in[274]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[275]) );
  DFF \start_reg_reg[276]  ( .D(start_in[275]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[276]) );
  DFF \start_reg_reg[277]  ( .D(start_in[276]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[277]) );
  DFF \start_reg_reg[278]  ( .D(start_in[277]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[278]) );
  DFF \start_reg_reg[279]  ( .D(start_in[278]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[279]) );
  DFF \start_reg_reg[280]  ( .D(start_in[279]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[280]) );
  DFF \start_reg_reg[281]  ( .D(start_in[280]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[281]) );
  DFF \start_reg_reg[282]  ( .D(start_in[281]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[282]) );
  DFF \start_reg_reg[283]  ( .D(start_in[282]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[283]) );
  DFF \start_reg_reg[284]  ( .D(start_in[283]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[284]) );
  DFF \start_reg_reg[285]  ( .D(start_in[284]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[285]) );
  DFF \start_reg_reg[286]  ( .D(start_in[285]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[286]) );
  DFF \start_reg_reg[287]  ( .D(start_in[286]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[287]) );
  DFF \start_reg_reg[288]  ( .D(start_in[287]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[288]) );
  DFF \start_reg_reg[289]  ( .D(start_in[288]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[289]) );
  DFF \start_reg_reg[290]  ( .D(start_in[289]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[290]) );
  DFF \start_reg_reg[291]  ( .D(start_in[290]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[291]) );
  DFF \start_reg_reg[292]  ( .D(start_in[291]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[292]) );
  DFF \start_reg_reg[293]  ( .D(start_in[292]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[293]) );
  DFF \start_reg_reg[294]  ( .D(start_in[293]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[294]) );
  DFF \start_reg_reg[295]  ( .D(start_in[294]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[295]) );
  DFF \start_reg_reg[296]  ( .D(start_in[295]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[296]) );
  DFF \start_reg_reg[297]  ( .D(start_in[296]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[297]) );
  DFF \start_reg_reg[298]  ( .D(start_in[297]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[298]) );
  DFF \start_reg_reg[299]  ( .D(start_in[298]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[299]) );
  DFF \start_reg_reg[300]  ( .D(start_in[299]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[300]) );
  DFF \start_reg_reg[301]  ( .D(start_in[300]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[301]) );
  DFF \start_reg_reg[302]  ( .D(start_in[301]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[302]) );
  DFF \start_reg_reg[303]  ( .D(start_in[302]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[303]) );
  DFF \start_reg_reg[304]  ( .D(start_in[303]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[304]) );
  DFF \start_reg_reg[305]  ( .D(start_in[304]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[305]) );
  DFF \start_reg_reg[306]  ( .D(start_in[305]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[306]) );
  DFF \start_reg_reg[307]  ( .D(start_in[306]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[307]) );
  DFF \start_reg_reg[308]  ( .D(start_in[307]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[308]) );
  DFF \start_reg_reg[309]  ( .D(start_in[308]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[309]) );
  DFF \start_reg_reg[310]  ( .D(start_in[309]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[310]) );
  DFF \start_reg_reg[311]  ( .D(start_in[310]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[311]) );
  DFF \start_reg_reg[312]  ( .D(start_in[311]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[312]) );
  DFF \start_reg_reg[313]  ( .D(start_in[312]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[313]) );
  DFF \start_reg_reg[314]  ( .D(start_in[313]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[314]) );
  DFF \start_reg_reg[315]  ( .D(start_in[314]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[315]) );
  DFF \start_reg_reg[316]  ( .D(start_in[315]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[316]) );
  DFF \start_reg_reg[317]  ( .D(start_in[316]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[317]) );
  DFF \start_reg_reg[318]  ( .D(start_in[317]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[318]) );
  DFF \start_reg_reg[319]  ( .D(start_in[318]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[319]) );
  DFF \start_reg_reg[320]  ( .D(start_in[319]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[320]) );
  DFF \start_reg_reg[321]  ( .D(start_in[320]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[321]) );
  DFF \start_reg_reg[322]  ( .D(start_in[321]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[322]) );
  DFF \start_reg_reg[323]  ( .D(start_in[322]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[323]) );
  DFF \start_reg_reg[324]  ( .D(start_in[323]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[324]) );
  DFF \start_reg_reg[325]  ( .D(start_in[324]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[325]) );
  DFF \start_reg_reg[326]  ( .D(start_in[325]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[326]) );
  DFF \start_reg_reg[327]  ( .D(start_in[326]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[327]) );
  DFF \start_reg_reg[328]  ( .D(start_in[327]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[328]) );
  DFF \start_reg_reg[329]  ( .D(start_in[328]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[329]) );
  DFF \start_reg_reg[330]  ( .D(start_in[329]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[330]) );
  DFF \start_reg_reg[331]  ( .D(start_in[330]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[331]) );
  DFF \start_reg_reg[332]  ( .D(start_in[331]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[332]) );
  DFF \start_reg_reg[333]  ( .D(start_in[332]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[333]) );
  DFF \start_reg_reg[334]  ( .D(start_in[333]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[334]) );
  DFF \start_reg_reg[335]  ( .D(start_in[334]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[335]) );
  DFF \start_reg_reg[336]  ( .D(start_in[335]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[336]) );
  DFF \start_reg_reg[337]  ( .D(start_in[336]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[337]) );
  DFF \start_reg_reg[338]  ( .D(start_in[337]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[338]) );
  DFF \start_reg_reg[339]  ( .D(start_in[338]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[339]) );
  DFF \start_reg_reg[340]  ( .D(start_in[339]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[340]) );
  DFF \start_reg_reg[341]  ( .D(start_in[340]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[341]) );
  DFF \start_reg_reg[342]  ( .D(start_in[341]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[342]) );
  DFF \start_reg_reg[343]  ( .D(start_in[342]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[343]) );
  DFF \start_reg_reg[344]  ( .D(start_in[343]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[344]) );
  DFF \start_reg_reg[345]  ( .D(start_in[344]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[345]) );
  DFF \start_reg_reg[346]  ( .D(start_in[345]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[346]) );
  DFF \start_reg_reg[347]  ( .D(start_in[346]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[347]) );
  DFF \start_reg_reg[348]  ( .D(start_in[347]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[348]) );
  DFF \start_reg_reg[349]  ( .D(start_in[348]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[349]) );
  DFF \start_reg_reg[350]  ( .D(start_in[349]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[350]) );
  DFF \start_reg_reg[351]  ( .D(start_in[350]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[351]) );
  DFF \start_reg_reg[352]  ( .D(start_in[351]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[352]) );
  DFF \start_reg_reg[353]  ( .D(start_in[352]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[353]) );
  DFF \start_reg_reg[354]  ( .D(start_in[353]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[354]) );
  DFF \start_reg_reg[355]  ( .D(start_in[354]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[355]) );
  DFF \start_reg_reg[356]  ( .D(start_in[355]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[356]) );
  DFF \start_reg_reg[357]  ( .D(start_in[356]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[357]) );
  DFF \start_reg_reg[358]  ( .D(start_in[357]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[358]) );
  DFF \start_reg_reg[359]  ( .D(start_in[358]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[359]) );
  DFF \start_reg_reg[360]  ( .D(start_in[359]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[360]) );
  DFF \start_reg_reg[361]  ( .D(start_in[360]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[361]) );
  DFF \start_reg_reg[362]  ( .D(start_in[361]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[362]) );
  DFF \start_reg_reg[363]  ( .D(start_in[362]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[363]) );
  DFF \start_reg_reg[364]  ( .D(start_in[363]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[364]) );
  DFF \start_reg_reg[365]  ( .D(start_in[364]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[365]) );
  DFF \start_reg_reg[366]  ( .D(start_in[365]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[366]) );
  DFF \start_reg_reg[367]  ( .D(start_in[366]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[367]) );
  DFF \start_reg_reg[368]  ( .D(start_in[367]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[368]) );
  DFF \start_reg_reg[369]  ( .D(start_in[368]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[369]) );
  DFF \start_reg_reg[370]  ( .D(start_in[369]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[370]) );
  DFF \start_reg_reg[371]  ( .D(start_in[370]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[371]) );
  DFF \start_reg_reg[372]  ( .D(start_in[371]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[372]) );
  DFF \start_reg_reg[373]  ( .D(start_in[372]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[373]) );
  DFF \start_reg_reg[374]  ( .D(start_in[373]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[374]) );
  DFF \start_reg_reg[375]  ( .D(start_in[374]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[375]) );
  DFF \start_reg_reg[376]  ( .D(start_in[375]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[376]) );
  DFF \start_reg_reg[377]  ( .D(start_in[376]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[377]) );
  DFF \start_reg_reg[378]  ( .D(start_in[377]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[378]) );
  DFF \start_reg_reg[379]  ( .D(start_in[378]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[379]) );
  DFF \start_reg_reg[380]  ( .D(start_in[379]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[380]) );
  DFF \start_reg_reg[381]  ( .D(start_in[380]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[381]) );
  DFF \start_reg_reg[382]  ( .D(start_in[381]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[382]) );
  DFF \start_reg_reg[383]  ( .D(start_in[382]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[383]) );
  DFF \start_reg_reg[384]  ( .D(start_in[383]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[384]) );
  DFF \start_reg_reg[385]  ( .D(start_in[384]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[385]) );
  DFF \start_reg_reg[386]  ( .D(start_in[385]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[386]) );
  DFF \start_reg_reg[387]  ( .D(start_in[386]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[387]) );
  DFF \start_reg_reg[388]  ( .D(start_in[387]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[388]) );
  DFF \start_reg_reg[389]  ( .D(start_in[388]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[389]) );
  DFF \start_reg_reg[390]  ( .D(start_in[389]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[390]) );
  DFF \start_reg_reg[391]  ( .D(start_in[390]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[391]) );
  DFF \start_reg_reg[392]  ( .D(start_in[391]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[392]) );
  DFF \start_reg_reg[393]  ( .D(start_in[392]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[393]) );
  DFF \start_reg_reg[394]  ( .D(start_in[393]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[394]) );
  DFF \start_reg_reg[395]  ( .D(start_in[394]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[395]) );
  DFF \start_reg_reg[396]  ( .D(start_in[395]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[396]) );
  DFF \start_reg_reg[397]  ( .D(start_in[396]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[397]) );
  DFF \start_reg_reg[398]  ( .D(start_in[397]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[398]) );
  DFF \start_reg_reg[399]  ( .D(start_in[398]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[399]) );
  DFF \start_reg_reg[400]  ( .D(start_in[399]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[400]) );
  DFF \start_reg_reg[401]  ( .D(start_in[400]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[401]) );
  DFF \start_reg_reg[402]  ( .D(start_in[401]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[402]) );
  DFF \start_reg_reg[403]  ( .D(start_in[402]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[403]) );
  DFF \start_reg_reg[404]  ( .D(start_in[403]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[404]) );
  DFF \start_reg_reg[405]  ( .D(start_in[404]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[405]) );
  DFF \start_reg_reg[406]  ( .D(start_in[405]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[406]) );
  DFF \start_reg_reg[407]  ( .D(start_in[406]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[407]) );
  DFF \start_reg_reg[408]  ( .D(start_in[407]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[408]) );
  DFF \start_reg_reg[409]  ( .D(start_in[408]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[409]) );
  DFF \start_reg_reg[410]  ( .D(start_in[409]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[410]) );
  DFF \start_reg_reg[411]  ( .D(start_in[410]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[411]) );
  DFF \start_reg_reg[412]  ( .D(start_in[411]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[412]) );
  DFF \start_reg_reg[413]  ( .D(start_in[412]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[413]) );
  DFF \start_reg_reg[414]  ( .D(start_in[413]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[414]) );
  DFF \start_reg_reg[415]  ( .D(start_in[414]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[415]) );
  DFF \start_reg_reg[416]  ( .D(start_in[415]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[416]) );
  DFF \start_reg_reg[417]  ( .D(start_in[416]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[417]) );
  DFF \start_reg_reg[418]  ( .D(start_in[417]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[418]) );
  DFF \start_reg_reg[419]  ( .D(start_in[418]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[419]) );
  DFF \start_reg_reg[420]  ( .D(start_in[419]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[420]) );
  DFF \start_reg_reg[421]  ( .D(start_in[420]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[421]) );
  DFF \start_reg_reg[422]  ( .D(start_in[421]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[422]) );
  DFF \start_reg_reg[423]  ( .D(start_in[422]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[423]) );
  DFF \start_reg_reg[424]  ( .D(start_in[423]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[424]) );
  DFF \start_reg_reg[425]  ( .D(start_in[424]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[425]) );
  DFF \start_reg_reg[426]  ( .D(start_in[425]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[426]) );
  DFF \start_reg_reg[427]  ( .D(start_in[426]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[427]) );
  DFF \start_reg_reg[428]  ( .D(start_in[427]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[428]) );
  DFF \start_reg_reg[429]  ( .D(start_in[428]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[429]) );
  DFF \start_reg_reg[430]  ( .D(start_in[429]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[430]) );
  DFF \start_reg_reg[431]  ( .D(start_in[430]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[431]) );
  DFF \start_reg_reg[432]  ( .D(start_in[431]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[432]) );
  DFF \start_reg_reg[433]  ( .D(start_in[432]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[433]) );
  DFF \start_reg_reg[434]  ( .D(start_in[433]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[434]) );
  DFF \start_reg_reg[435]  ( .D(start_in[434]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[435]) );
  DFF \start_reg_reg[436]  ( .D(start_in[435]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[436]) );
  DFF \start_reg_reg[437]  ( .D(start_in[436]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[437]) );
  DFF \start_reg_reg[438]  ( .D(start_in[437]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[438]) );
  DFF \start_reg_reg[439]  ( .D(start_in[438]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[439]) );
  DFF \start_reg_reg[440]  ( .D(start_in[439]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[440]) );
  DFF \start_reg_reg[441]  ( .D(start_in[440]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[441]) );
  DFF \start_reg_reg[442]  ( .D(start_in[441]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[442]) );
  DFF \start_reg_reg[443]  ( .D(start_in[442]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[443]) );
  DFF \start_reg_reg[444]  ( .D(start_in[443]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[444]) );
  DFF \start_reg_reg[445]  ( .D(start_in[444]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[445]) );
  DFF \start_reg_reg[446]  ( .D(start_in[445]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[446]) );
  DFF \start_reg_reg[447]  ( .D(start_in[446]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[447]) );
  DFF \start_reg_reg[448]  ( .D(start_in[447]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[448]) );
  DFF \start_reg_reg[449]  ( .D(start_in[448]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[449]) );
  DFF \start_reg_reg[450]  ( .D(start_in[449]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[450]) );
  DFF \start_reg_reg[451]  ( .D(start_in[450]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[451]) );
  DFF \start_reg_reg[452]  ( .D(start_in[451]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[452]) );
  DFF \start_reg_reg[453]  ( .D(start_in[452]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[453]) );
  DFF \start_reg_reg[454]  ( .D(start_in[453]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[454]) );
  DFF \start_reg_reg[455]  ( .D(start_in[454]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[455]) );
  DFF \start_reg_reg[456]  ( .D(start_in[455]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[456]) );
  DFF \start_reg_reg[457]  ( .D(start_in[456]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[457]) );
  DFF \start_reg_reg[458]  ( .D(start_in[457]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[458]) );
  DFF \start_reg_reg[459]  ( .D(start_in[458]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[459]) );
  DFF \start_reg_reg[460]  ( .D(start_in[459]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[460]) );
  DFF \start_reg_reg[461]  ( .D(start_in[460]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[461]) );
  DFF \start_reg_reg[462]  ( .D(start_in[461]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[462]) );
  DFF \start_reg_reg[463]  ( .D(start_in[462]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[463]) );
  DFF \start_reg_reg[464]  ( .D(start_in[463]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[464]) );
  DFF \start_reg_reg[465]  ( .D(start_in[464]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[465]) );
  DFF \start_reg_reg[466]  ( .D(start_in[465]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[466]) );
  DFF \start_reg_reg[467]  ( .D(start_in[466]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[467]) );
  DFF \start_reg_reg[468]  ( .D(start_in[467]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[468]) );
  DFF \start_reg_reg[469]  ( .D(start_in[468]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[469]) );
  DFF \start_reg_reg[470]  ( .D(start_in[469]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[470]) );
  DFF \start_reg_reg[471]  ( .D(start_in[470]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[471]) );
  DFF \start_reg_reg[472]  ( .D(start_in[471]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[472]) );
  DFF \start_reg_reg[473]  ( .D(start_in[472]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[473]) );
  DFF \start_reg_reg[474]  ( .D(start_in[473]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[474]) );
  DFF \start_reg_reg[475]  ( .D(start_in[474]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[475]) );
  DFF \start_reg_reg[476]  ( .D(start_in[475]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[476]) );
  DFF \start_reg_reg[477]  ( .D(start_in[476]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[477]) );
  DFF \start_reg_reg[478]  ( .D(start_in[477]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[478]) );
  DFF \start_reg_reg[479]  ( .D(start_in[478]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[479]) );
  DFF \start_reg_reg[480]  ( .D(start_in[479]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[480]) );
  DFF \start_reg_reg[481]  ( .D(start_in[480]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[481]) );
  DFF \start_reg_reg[482]  ( .D(start_in[481]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[482]) );
  DFF \start_reg_reg[483]  ( .D(start_in[482]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[483]) );
  DFF \start_reg_reg[484]  ( .D(start_in[483]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[484]) );
  DFF \start_reg_reg[485]  ( .D(start_in[484]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[485]) );
  DFF \start_reg_reg[486]  ( .D(start_in[485]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[486]) );
  DFF \start_reg_reg[487]  ( .D(start_in[486]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[487]) );
  DFF \start_reg_reg[488]  ( .D(start_in[487]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[488]) );
  DFF \start_reg_reg[489]  ( .D(start_in[488]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[489]) );
  DFF \start_reg_reg[490]  ( .D(start_in[489]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[490]) );
  DFF \start_reg_reg[491]  ( .D(start_in[490]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[491]) );
  DFF \start_reg_reg[492]  ( .D(start_in[491]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[492]) );
  DFF \start_reg_reg[493]  ( .D(start_in[492]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[493]) );
  DFF \start_reg_reg[494]  ( .D(start_in[493]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[494]) );
  DFF \start_reg_reg[495]  ( .D(start_in[494]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[495]) );
  DFF \start_reg_reg[496]  ( .D(start_in[495]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[496]) );
  DFF \start_reg_reg[497]  ( .D(start_in[496]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[497]) );
  DFF \start_reg_reg[498]  ( .D(start_in[497]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[498]) );
  DFF \start_reg_reg[499]  ( .D(start_in[498]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[499]) );
  DFF \start_reg_reg[500]  ( .D(start_in[499]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[500]) );
  DFF \start_reg_reg[501]  ( .D(start_in[500]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[501]) );
  DFF \start_reg_reg[502]  ( .D(start_in[501]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[502]) );
  DFF \start_reg_reg[503]  ( .D(start_in[502]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[503]) );
  DFF \start_reg_reg[504]  ( .D(start_in[503]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[504]) );
  DFF \start_reg_reg[505]  ( .D(start_in[504]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[505]) );
  DFF \start_reg_reg[506]  ( .D(start_in[505]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[506]) );
  DFF \start_reg_reg[507]  ( .D(start_in[506]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[507]) );
  DFF \start_reg_reg[508]  ( .D(start_in[507]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[508]) );
  DFF \start_reg_reg[509]  ( .D(start_in[508]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[509]) );
  DFF \start_reg_reg[510]  ( .D(start_in[509]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[510]) );
  DFF \start_reg_reg[511]  ( .D(start_in[510]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[511]) );
  DFF \start_reg_reg[512]  ( .D(start_in[511]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[512]) );
  DFF \start_reg_reg[513]  ( .D(start_in[512]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[513]) );
  DFF \start_reg_reg[514]  ( .D(start_in[513]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[514]) );
  DFF \start_reg_reg[515]  ( .D(start_in[514]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[515]) );
  DFF \start_reg_reg[516]  ( .D(start_in[515]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[516]) );
  DFF \start_reg_reg[517]  ( .D(start_in[516]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[517]) );
  DFF \start_reg_reg[518]  ( .D(start_in[517]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[518]) );
  DFF \start_reg_reg[519]  ( .D(start_in[518]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[519]) );
  DFF \start_reg_reg[520]  ( .D(start_in[519]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[520]) );
  DFF \start_reg_reg[521]  ( .D(start_in[520]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[521]) );
  DFF \start_reg_reg[522]  ( .D(start_in[521]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[522]) );
  DFF \start_reg_reg[523]  ( .D(start_in[522]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[523]) );
  DFF \start_reg_reg[524]  ( .D(start_in[523]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[524]) );
  DFF \start_reg_reg[525]  ( .D(start_in[524]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[525]) );
  DFF \start_reg_reg[526]  ( .D(start_in[525]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[526]) );
  DFF \start_reg_reg[527]  ( .D(start_in[526]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[527]) );
  DFF \start_reg_reg[528]  ( .D(start_in[527]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[528]) );
  DFF \start_reg_reg[529]  ( .D(start_in[528]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[529]) );
  DFF \start_reg_reg[530]  ( .D(start_in[529]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[530]) );
  DFF \start_reg_reg[531]  ( .D(start_in[530]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[531]) );
  DFF \start_reg_reg[532]  ( .D(start_in[531]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[532]) );
  DFF \start_reg_reg[533]  ( .D(start_in[532]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[533]) );
  DFF \start_reg_reg[534]  ( .D(start_in[533]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[534]) );
  DFF \start_reg_reg[535]  ( .D(start_in[534]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[535]) );
  DFF \start_reg_reg[536]  ( .D(start_in[535]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[536]) );
  DFF \start_reg_reg[537]  ( .D(start_in[536]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[537]) );
  DFF \start_reg_reg[538]  ( .D(start_in[537]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[538]) );
  DFF \start_reg_reg[539]  ( .D(start_in[538]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[539]) );
  DFF \start_reg_reg[540]  ( .D(start_in[539]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[540]) );
  DFF \start_reg_reg[541]  ( .D(start_in[540]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[541]) );
  DFF \start_reg_reg[542]  ( .D(start_in[541]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[542]) );
  DFF \start_reg_reg[543]  ( .D(start_in[542]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[543]) );
  DFF \start_reg_reg[544]  ( .D(start_in[543]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[544]) );
  DFF \start_reg_reg[545]  ( .D(start_in[544]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[545]) );
  DFF \start_reg_reg[546]  ( .D(start_in[545]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[546]) );
  DFF \start_reg_reg[547]  ( .D(start_in[546]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[547]) );
  DFF \start_reg_reg[548]  ( .D(start_in[547]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[548]) );
  DFF \start_reg_reg[549]  ( .D(start_in[548]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[549]) );
  DFF \start_reg_reg[550]  ( .D(start_in[549]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[550]) );
  DFF \start_reg_reg[551]  ( .D(start_in[550]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[551]) );
  DFF \start_reg_reg[552]  ( .D(start_in[551]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[552]) );
  DFF \start_reg_reg[553]  ( .D(start_in[552]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[553]) );
  DFF \start_reg_reg[554]  ( .D(start_in[553]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[554]) );
  DFF \start_reg_reg[555]  ( .D(start_in[554]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[555]) );
  DFF \start_reg_reg[556]  ( .D(start_in[555]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[556]) );
  DFF \start_reg_reg[557]  ( .D(start_in[556]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[557]) );
  DFF \start_reg_reg[558]  ( .D(start_in[557]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[558]) );
  DFF \start_reg_reg[559]  ( .D(start_in[558]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[559]) );
  DFF \start_reg_reg[560]  ( .D(start_in[559]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[560]) );
  DFF \start_reg_reg[561]  ( .D(start_in[560]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[561]) );
  DFF \start_reg_reg[562]  ( .D(start_in[561]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[562]) );
  DFF \start_reg_reg[563]  ( .D(start_in[562]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[563]) );
  DFF \start_reg_reg[564]  ( .D(start_in[563]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[564]) );
  DFF \start_reg_reg[565]  ( .D(start_in[564]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[565]) );
  DFF \start_reg_reg[566]  ( .D(start_in[565]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[566]) );
  DFF \start_reg_reg[567]  ( .D(start_in[566]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[567]) );
  DFF \start_reg_reg[568]  ( .D(start_in[567]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[568]) );
  DFF \start_reg_reg[569]  ( .D(start_in[568]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[569]) );
  DFF \start_reg_reg[570]  ( .D(start_in[569]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[570]) );
  DFF \start_reg_reg[571]  ( .D(start_in[570]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[571]) );
  DFF \start_reg_reg[572]  ( .D(start_in[571]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[572]) );
  DFF \start_reg_reg[573]  ( .D(start_in[572]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[573]) );
  DFF \start_reg_reg[574]  ( .D(start_in[573]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[574]) );
  DFF \start_reg_reg[575]  ( .D(start_in[574]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[575]) );
  DFF \start_reg_reg[576]  ( .D(start_in[575]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[576]) );
  DFF \start_reg_reg[577]  ( .D(start_in[576]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[577]) );
  DFF \start_reg_reg[578]  ( .D(start_in[577]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[578]) );
  DFF \start_reg_reg[579]  ( .D(start_in[578]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[579]) );
  DFF \start_reg_reg[580]  ( .D(start_in[579]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[580]) );
  DFF \start_reg_reg[581]  ( .D(start_in[580]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[581]) );
  DFF \start_reg_reg[582]  ( .D(start_in[581]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[582]) );
  DFF \start_reg_reg[583]  ( .D(start_in[582]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[583]) );
  DFF \start_reg_reg[584]  ( .D(start_in[583]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[584]) );
  DFF \start_reg_reg[585]  ( .D(start_in[584]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[585]) );
  DFF \start_reg_reg[586]  ( .D(start_in[585]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[586]) );
  DFF \start_reg_reg[587]  ( .D(start_in[586]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[587]) );
  DFF \start_reg_reg[588]  ( .D(start_in[587]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[588]) );
  DFF \start_reg_reg[589]  ( .D(start_in[588]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[589]) );
  DFF \start_reg_reg[590]  ( .D(start_in[589]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[590]) );
  DFF \start_reg_reg[591]  ( .D(start_in[590]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[591]) );
  DFF \start_reg_reg[592]  ( .D(start_in[591]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[592]) );
  DFF \start_reg_reg[593]  ( .D(start_in[592]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[593]) );
  DFF \start_reg_reg[594]  ( .D(start_in[593]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[594]) );
  DFF \start_reg_reg[595]  ( .D(start_in[594]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[595]) );
  DFF \start_reg_reg[596]  ( .D(start_in[595]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[596]) );
  DFF \start_reg_reg[597]  ( .D(start_in[596]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[597]) );
  DFF \start_reg_reg[598]  ( .D(start_in[597]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[598]) );
  DFF \start_reg_reg[599]  ( .D(start_in[598]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[599]) );
  DFF \start_reg_reg[600]  ( .D(start_in[599]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[600]) );
  DFF \start_reg_reg[601]  ( .D(start_in[600]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[601]) );
  DFF \start_reg_reg[602]  ( .D(start_in[601]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[602]) );
  DFF \start_reg_reg[603]  ( .D(start_in[602]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[603]) );
  DFF \start_reg_reg[604]  ( .D(start_in[603]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[604]) );
  DFF \start_reg_reg[605]  ( .D(start_in[604]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[605]) );
  DFF \start_reg_reg[606]  ( .D(start_in[605]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[606]) );
  DFF \start_reg_reg[607]  ( .D(start_in[606]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[607]) );
  DFF \start_reg_reg[608]  ( .D(start_in[607]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[608]) );
  DFF \start_reg_reg[609]  ( .D(start_in[608]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[609]) );
  DFF \start_reg_reg[610]  ( .D(start_in[609]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[610]) );
  DFF \start_reg_reg[611]  ( .D(start_in[610]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[611]) );
  DFF \start_reg_reg[612]  ( .D(start_in[611]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[612]) );
  DFF \start_reg_reg[613]  ( .D(start_in[612]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[613]) );
  DFF \start_reg_reg[614]  ( .D(start_in[613]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[614]) );
  DFF \start_reg_reg[615]  ( .D(start_in[614]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[615]) );
  DFF \start_reg_reg[616]  ( .D(start_in[615]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[616]) );
  DFF \start_reg_reg[617]  ( .D(start_in[616]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[617]) );
  DFF \start_reg_reg[618]  ( .D(start_in[617]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[618]) );
  DFF \start_reg_reg[619]  ( .D(start_in[618]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[619]) );
  DFF \start_reg_reg[620]  ( .D(start_in[619]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[620]) );
  DFF \start_reg_reg[621]  ( .D(start_in[620]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[621]) );
  DFF \start_reg_reg[622]  ( .D(start_in[621]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[622]) );
  DFF \start_reg_reg[623]  ( .D(start_in[622]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[623]) );
  DFF \start_reg_reg[624]  ( .D(start_in[623]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[624]) );
  DFF \start_reg_reg[625]  ( .D(start_in[624]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[625]) );
  DFF \start_reg_reg[626]  ( .D(start_in[625]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[626]) );
  DFF \start_reg_reg[627]  ( .D(start_in[626]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[627]) );
  DFF \start_reg_reg[628]  ( .D(start_in[627]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[628]) );
  DFF \start_reg_reg[629]  ( .D(start_in[628]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[629]) );
  DFF \start_reg_reg[630]  ( .D(start_in[629]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[630]) );
  DFF \start_reg_reg[631]  ( .D(start_in[630]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[631]) );
  DFF \start_reg_reg[632]  ( .D(start_in[631]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[632]) );
  DFF \start_reg_reg[633]  ( .D(start_in[632]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[633]) );
  DFF \start_reg_reg[634]  ( .D(start_in[633]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[634]) );
  DFF \start_reg_reg[635]  ( .D(start_in[634]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[635]) );
  DFF \start_reg_reg[636]  ( .D(start_in[635]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[636]) );
  DFF \start_reg_reg[637]  ( .D(start_in[636]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[637]) );
  DFF \start_reg_reg[638]  ( .D(start_in[637]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[638]) );
  DFF \start_reg_reg[639]  ( .D(start_in[638]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[639]) );
  DFF \start_reg_reg[640]  ( .D(start_in[639]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[640]) );
  DFF \start_reg_reg[641]  ( .D(start_in[640]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[641]) );
  DFF \start_reg_reg[642]  ( .D(start_in[641]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[642]) );
  DFF \start_reg_reg[643]  ( .D(start_in[642]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[643]) );
  DFF \start_reg_reg[644]  ( .D(start_in[643]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[644]) );
  DFF \start_reg_reg[645]  ( .D(start_in[644]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[645]) );
  DFF \start_reg_reg[646]  ( .D(start_in[645]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[646]) );
  DFF \start_reg_reg[647]  ( .D(start_in[646]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[647]) );
  DFF \start_reg_reg[648]  ( .D(start_in[647]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[648]) );
  DFF \start_reg_reg[649]  ( .D(start_in[648]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[649]) );
  DFF \start_reg_reg[650]  ( .D(start_in[649]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[650]) );
  DFF \start_reg_reg[651]  ( .D(start_in[650]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[651]) );
  DFF \start_reg_reg[652]  ( .D(start_in[651]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[652]) );
  DFF \start_reg_reg[653]  ( .D(start_in[652]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[653]) );
  DFF \start_reg_reg[654]  ( .D(start_in[653]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[654]) );
  DFF \start_reg_reg[655]  ( .D(start_in[654]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[655]) );
  DFF \start_reg_reg[656]  ( .D(start_in[655]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[656]) );
  DFF \start_reg_reg[657]  ( .D(start_in[656]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[657]) );
  DFF \start_reg_reg[658]  ( .D(start_in[657]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[658]) );
  DFF \start_reg_reg[659]  ( .D(start_in[658]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[659]) );
  DFF \start_reg_reg[660]  ( .D(start_in[659]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[660]) );
  DFF \start_reg_reg[661]  ( .D(start_in[660]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[661]) );
  DFF \start_reg_reg[662]  ( .D(start_in[661]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[662]) );
  DFF \start_reg_reg[663]  ( .D(start_in[662]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[663]) );
  DFF \start_reg_reg[664]  ( .D(start_in[663]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[664]) );
  DFF \start_reg_reg[665]  ( .D(start_in[664]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[665]) );
  DFF \start_reg_reg[666]  ( .D(start_in[665]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[666]) );
  DFF \start_reg_reg[667]  ( .D(start_in[666]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[667]) );
  DFF \start_reg_reg[668]  ( .D(start_in[667]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[668]) );
  DFF \start_reg_reg[669]  ( .D(start_in[668]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[669]) );
  DFF \start_reg_reg[670]  ( .D(start_in[669]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[670]) );
  DFF \start_reg_reg[671]  ( .D(start_in[670]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[671]) );
  DFF \start_reg_reg[672]  ( .D(start_in[671]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[672]) );
  DFF \start_reg_reg[673]  ( .D(start_in[672]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[673]) );
  DFF \start_reg_reg[674]  ( .D(start_in[673]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[674]) );
  DFF \start_reg_reg[675]  ( .D(start_in[674]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[675]) );
  DFF \start_reg_reg[676]  ( .D(start_in[675]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[676]) );
  DFF \start_reg_reg[677]  ( .D(start_in[676]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[677]) );
  DFF \start_reg_reg[678]  ( .D(start_in[677]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[678]) );
  DFF \start_reg_reg[679]  ( .D(start_in[678]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[679]) );
  DFF \start_reg_reg[680]  ( .D(start_in[679]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[680]) );
  DFF \start_reg_reg[681]  ( .D(start_in[680]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[681]) );
  DFF \start_reg_reg[682]  ( .D(start_in[681]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[682]) );
  DFF \start_reg_reg[683]  ( .D(start_in[682]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[683]) );
  DFF \start_reg_reg[684]  ( .D(start_in[683]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[684]) );
  DFF \start_reg_reg[685]  ( .D(start_in[684]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[685]) );
  DFF \start_reg_reg[686]  ( .D(start_in[685]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[686]) );
  DFF \start_reg_reg[687]  ( .D(start_in[686]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[687]) );
  DFF \start_reg_reg[688]  ( .D(start_in[687]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[688]) );
  DFF \start_reg_reg[689]  ( .D(start_in[688]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[689]) );
  DFF \start_reg_reg[690]  ( .D(start_in[689]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[690]) );
  DFF \start_reg_reg[691]  ( .D(start_in[690]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[691]) );
  DFF \start_reg_reg[692]  ( .D(start_in[691]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[692]) );
  DFF \start_reg_reg[693]  ( .D(start_in[692]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[693]) );
  DFF \start_reg_reg[694]  ( .D(start_in[693]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[694]) );
  DFF \start_reg_reg[695]  ( .D(start_in[694]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[695]) );
  DFF \start_reg_reg[696]  ( .D(start_in[695]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[696]) );
  DFF \start_reg_reg[697]  ( .D(start_in[696]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[697]) );
  DFF \start_reg_reg[698]  ( .D(start_in[697]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[698]) );
  DFF \start_reg_reg[699]  ( .D(start_in[698]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[699]) );
  DFF \start_reg_reg[700]  ( .D(start_in[699]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[700]) );
  DFF \start_reg_reg[701]  ( .D(start_in[700]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[701]) );
  DFF \start_reg_reg[702]  ( .D(start_in[701]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[702]) );
  DFF \start_reg_reg[703]  ( .D(start_in[702]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[703]) );
  DFF \start_reg_reg[704]  ( .D(start_in[703]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[704]) );
  DFF \start_reg_reg[705]  ( .D(start_in[704]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[705]) );
  DFF \start_reg_reg[706]  ( .D(start_in[705]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[706]) );
  DFF \start_reg_reg[707]  ( .D(start_in[706]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[707]) );
  DFF \start_reg_reg[708]  ( .D(start_in[707]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[708]) );
  DFF \start_reg_reg[709]  ( .D(start_in[708]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[709]) );
  DFF \start_reg_reg[710]  ( .D(start_in[709]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[710]) );
  DFF \start_reg_reg[711]  ( .D(start_in[710]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[711]) );
  DFF \start_reg_reg[712]  ( .D(start_in[711]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[712]) );
  DFF \start_reg_reg[713]  ( .D(start_in[712]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[713]) );
  DFF \start_reg_reg[714]  ( .D(start_in[713]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[714]) );
  DFF \start_reg_reg[715]  ( .D(start_in[714]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[715]) );
  DFF \start_reg_reg[716]  ( .D(start_in[715]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[716]) );
  DFF \start_reg_reg[717]  ( .D(start_in[716]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[717]) );
  DFF \start_reg_reg[718]  ( .D(start_in[717]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[718]) );
  DFF \start_reg_reg[719]  ( .D(start_in[718]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[719]) );
  DFF \start_reg_reg[720]  ( .D(start_in[719]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[720]) );
  DFF \start_reg_reg[721]  ( .D(start_in[720]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[721]) );
  DFF \start_reg_reg[722]  ( .D(start_in[721]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[722]) );
  DFF \start_reg_reg[723]  ( .D(start_in[722]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[723]) );
  DFF \start_reg_reg[724]  ( .D(start_in[723]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[724]) );
  DFF \start_reg_reg[725]  ( .D(start_in[724]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[725]) );
  DFF \start_reg_reg[726]  ( .D(start_in[725]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[726]) );
  DFF \start_reg_reg[727]  ( .D(start_in[726]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[727]) );
  DFF \start_reg_reg[728]  ( .D(start_in[727]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[728]) );
  DFF \start_reg_reg[729]  ( .D(start_in[728]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[729]) );
  DFF \start_reg_reg[730]  ( .D(start_in[729]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[730]) );
  DFF \start_reg_reg[731]  ( .D(start_in[730]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[731]) );
  DFF \start_reg_reg[732]  ( .D(start_in[731]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[732]) );
  DFF \start_reg_reg[733]  ( .D(start_in[732]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[733]) );
  DFF \start_reg_reg[734]  ( .D(start_in[733]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[734]) );
  DFF \start_reg_reg[735]  ( .D(start_in[734]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[735]) );
  DFF \start_reg_reg[736]  ( .D(start_in[735]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[736]) );
  DFF \start_reg_reg[737]  ( .D(start_in[736]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[737]) );
  DFF \start_reg_reg[738]  ( .D(start_in[737]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[738]) );
  DFF \start_reg_reg[739]  ( .D(start_in[738]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[739]) );
  DFF \start_reg_reg[740]  ( .D(start_in[739]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[740]) );
  DFF \start_reg_reg[741]  ( .D(start_in[740]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[741]) );
  DFF \start_reg_reg[742]  ( .D(start_in[741]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[742]) );
  DFF \start_reg_reg[743]  ( .D(start_in[742]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[743]) );
  DFF \start_reg_reg[744]  ( .D(start_in[743]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[744]) );
  DFF \start_reg_reg[745]  ( .D(start_in[744]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[745]) );
  DFF \start_reg_reg[746]  ( .D(start_in[745]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[746]) );
  DFF \start_reg_reg[747]  ( .D(start_in[746]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[747]) );
  DFF \start_reg_reg[748]  ( .D(start_in[747]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[748]) );
  DFF \start_reg_reg[749]  ( .D(start_in[748]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[749]) );
  DFF \start_reg_reg[750]  ( .D(start_in[749]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[750]) );
  DFF \start_reg_reg[751]  ( .D(start_in[750]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[751]) );
  DFF \start_reg_reg[752]  ( .D(start_in[751]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[752]) );
  DFF \start_reg_reg[753]  ( .D(start_in[752]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[753]) );
  DFF \start_reg_reg[754]  ( .D(start_in[753]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[754]) );
  DFF \start_reg_reg[755]  ( .D(start_in[754]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[755]) );
  DFF \start_reg_reg[756]  ( .D(start_in[755]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[756]) );
  DFF \start_reg_reg[757]  ( .D(start_in[756]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[757]) );
  DFF \start_reg_reg[758]  ( .D(start_in[757]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[758]) );
  DFF \start_reg_reg[759]  ( .D(start_in[758]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[759]) );
  DFF \start_reg_reg[760]  ( .D(start_in[759]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[760]) );
  DFF \start_reg_reg[761]  ( .D(start_in[760]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[761]) );
  DFF \start_reg_reg[762]  ( .D(start_in[761]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[762]) );
  DFF \start_reg_reg[763]  ( .D(start_in[762]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[763]) );
  DFF \start_reg_reg[764]  ( .D(start_in[763]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[764]) );
  DFF \start_reg_reg[765]  ( .D(start_in[764]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[765]) );
  DFF \start_reg_reg[766]  ( .D(start_in[765]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[766]) );
  DFF \start_reg_reg[767]  ( .D(start_in[766]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[767]) );
  DFF \start_reg_reg[768]  ( .D(start_in[767]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[768]) );
  DFF \start_reg_reg[769]  ( .D(start_in[768]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[769]) );
  DFF \start_reg_reg[770]  ( .D(start_in[769]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[770]) );
  DFF \start_reg_reg[771]  ( .D(start_in[770]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[771]) );
  DFF \start_reg_reg[772]  ( .D(start_in[771]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[772]) );
  DFF \start_reg_reg[773]  ( .D(start_in[772]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[773]) );
  DFF \start_reg_reg[774]  ( .D(start_in[773]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[774]) );
  DFF \start_reg_reg[775]  ( .D(start_in[774]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[775]) );
  DFF \start_reg_reg[776]  ( .D(start_in[775]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[776]) );
  DFF \start_reg_reg[777]  ( .D(start_in[776]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[777]) );
  DFF \start_reg_reg[778]  ( .D(start_in[777]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[778]) );
  DFF \start_reg_reg[779]  ( .D(start_in[778]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[779]) );
  DFF \start_reg_reg[780]  ( .D(start_in[779]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[780]) );
  DFF \start_reg_reg[781]  ( .D(start_in[780]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[781]) );
  DFF \start_reg_reg[782]  ( .D(start_in[781]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[782]) );
  DFF \start_reg_reg[783]  ( .D(start_in[782]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[783]) );
  DFF \start_reg_reg[784]  ( .D(start_in[783]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[784]) );
  DFF \start_reg_reg[785]  ( .D(start_in[784]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[785]) );
  DFF \start_reg_reg[786]  ( .D(start_in[785]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[786]) );
  DFF \start_reg_reg[787]  ( .D(start_in[786]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[787]) );
  DFF \start_reg_reg[788]  ( .D(start_in[787]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[788]) );
  DFF \start_reg_reg[789]  ( .D(start_in[788]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[789]) );
  DFF \start_reg_reg[790]  ( .D(start_in[789]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[790]) );
  DFF \start_reg_reg[791]  ( .D(start_in[790]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[791]) );
  DFF \start_reg_reg[792]  ( .D(start_in[791]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[792]) );
  DFF \start_reg_reg[793]  ( .D(start_in[792]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[793]) );
  DFF \start_reg_reg[794]  ( .D(start_in[793]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[794]) );
  DFF \start_reg_reg[795]  ( .D(start_in[794]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[795]) );
  DFF \start_reg_reg[796]  ( .D(start_in[795]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[796]) );
  DFF \start_reg_reg[797]  ( .D(start_in[796]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[797]) );
  DFF \start_reg_reg[798]  ( .D(start_in[797]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[798]) );
  DFF \start_reg_reg[799]  ( .D(start_in[798]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[799]) );
  DFF \start_reg_reg[800]  ( .D(start_in[799]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[800]) );
  DFF \start_reg_reg[801]  ( .D(start_in[800]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[801]) );
  DFF \start_reg_reg[802]  ( .D(start_in[801]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[802]) );
  DFF \start_reg_reg[803]  ( .D(start_in[802]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[803]) );
  DFF \start_reg_reg[804]  ( .D(start_in[803]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[804]) );
  DFF \start_reg_reg[805]  ( .D(start_in[804]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[805]) );
  DFF \start_reg_reg[806]  ( .D(start_in[805]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[806]) );
  DFF \start_reg_reg[807]  ( .D(start_in[806]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[807]) );
  DFF \start_reg_reg[808]  ( .D(start_in[807]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[808]) );
  DFF \start_reg_reg[809]  ( .D(start_in[808]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[809]) );
  DFF \start_reg_reg[810]  ( .D(start_in[809]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[810]) );
  DFF \start_reg_reg[811]  ( .D(start_in[810]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[811]) );
  DFF \start_reg_reg[812]  ( .D(start_in[811]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[812]) );
  DFF \start_reg_reg[813]  ( .D(start_in[812]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[813]) );
  DFF \start_reg_reg[814]  ( .D(start_in[813]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[814]) );
  DFF \start_reg_reg[815]  ( .D(start_in[814]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[815]) );
  DFF \start_reg_reg[816]  ( .D(start_in[815]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[816]) );
  DFF \start_reg_reg[817]  ( .D(start_in[816]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[817]) );
  DFF \start_reg_reg[818]  ( .D(start_in[817]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[818]) );
  DFF \start_reg_reg[819]  ( .D(start_in[818]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[819]) );
  DFF \start_reg_reg[820]  ( .D(start_in[819]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[820]) );
  DFF \start_reg_reg[821]  ( .D(start_in[820]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[821]) );
  DFF \start_reg_reg[822]  ( .D(start_in[821]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[822]) );
  DFF \start_reg_reg[823]  ( .D(start_in[822]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[823]) );
  DFF \start_reg_reg[824]  ( .D(start_in[823]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[824]) );
  DFF \start_reg_reg[825]  ( .D(start_in[824]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[825]) );
  DFF \start_reg_reg[826]  ( .D(start_in[825]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[826]) );
  DFF \start_reg_reg[827]  ( .D(start_in[826]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[827]) );
  DFF \start_reg_reg[828]  ( .D(start_in[827]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[828]) );
  DFF \start_reg_reg[829]  ( .D(start_in[828]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[829]) );
  DFF \start_reg_reg[830]  ( .D(start_in[829]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[830]) );
  DFF \start_reg_reg[831]  ( .D(start_in[830]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[831]) );
  DFF \start_reg_reg[832]  ( .D(start_in[831]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[832]) );
  DFF \start_reg_reg[833]  ( .D(start_in[832]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[833]) );
  DFF \start_reg_reg[834]  ( .D(start_in[833]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[834]) );
  DFF \start_reg_reg[835]  ( .D(start_in[834]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[835]) );
  DFF \start_reg_reg[836]  ( .D(start_in[835]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[836]) );
  DFF \start_reg_reg[837]  ( .D(start_in[836]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[837]) );
  DFF \start_reg_reg[838]  ( .D(start_in[837]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[838]) );
  DFF \start_reg_reg[839]  ( .D(start_in[838]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[839]) );
  DFF \start_reg_reg[840]  ( .D(start_in[839]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[840]) );
  DFF \start_reg_reg[841]  ( .D(start_in[840]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[841]) );
  DFF \start_reg_reg[842]  ( .D(start_in[841]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[842]) );
  DFF \start_reg_reg[843]  ( .D(start_in[842]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[843]) );
  DFF \start_reg_reg[844]  ( .D(start_in[843]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[844]) );
  DFF \start_reg_reg[845]  ( .D(start_in[844]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[845]) );
  DFF \start_reg_reg[846]  ( .D(start_in[845]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[846]) );
  DFF \start_reg_reg[847]  ( .D(start_in[846]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[847]) );
  DFF \start_reg_reg[848]  ( .D(start_in[847]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[848]) );
  DFF \start_reg_reg[849]  ( .D(start_in[848]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[849]) );
  DFF \start_reg_reg[850]  ( .D(start_in[849]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[850]) );
  DFF \start_reg_reg[851]  ( .D(start_in[850]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[851]) );
  DFF \start_reg_reg[852]  ( .D(start_in[851]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[852]) );
  DFF \start_reg_reg[853]  ( .D(start_in[852]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[853]) );
  DFF \start_reg_reg[854]  ( .D(start_in[853]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[854]) );
  DFF \start_reg_reg[855]  ( .D(start_in[854]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[855]) );
  DFF \start_reg_reg[856]  ( .D(start_in[855]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[856]) );
  DFF \start_reg_reg[857]  ( .D(start_in[856]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[857]) );
  DFF \start_reg_reg[858]  ( .D(start_in[857]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[858]) );
  DFF \start_reg_reg[859]  ( .D(start_in[858]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[859]) );
  DFF \start_reg_reg[860]  ( .D(start_in[859]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[860]) );
  DFF \start_reg_reg[861]  ( .D(start_in[860]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[861]) );
  DFF \start_reg_reg[862]  ( .D(start_in[861]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[862]) );
  DFF \start_reg_reg[863]  ( .D(start_in[862]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[863]) );
  DFF \start_reg_reg[864]  ( .D(start_in[863]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[864]) );
  DFF \start_reg_reg[865]  ( .D(start_in[864]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[865]) );
  DFF \start_reg_reg[866]  ( .D(start_in[865]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[866]) );
  DFF \start_reg_reg[867]  ( .D(start_in[866]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[867]) );
  DFF \start_reg_reg[868]  ( .D(start_in[867]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[868]) );
  DFF \start_reg_reg[869]  ( .D(start_in[868]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[869]) );
  DFF \start_reg_reg[870]  ( .D(start_in[869]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[870]) );
  DFF \start_reg_reg[871]  ( .D(start_in[870]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[871]) );
  DFF \start_reg_reg[872]  ( .D(start_in[871]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[872]) );
  DFF \start_reg_reg[873]  ( .D(start_in[872]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[873]) );
  DFF \start_reg_reg[874]  ( .D(start_in[873]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[874]) );
  DFF \start_reg_reg[875]  ( .D(start_in[874]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[875]) );
  DFF \start_reg_reg[876]  ( .D(start_in[875]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[876]) );
  DFF \start_reg_reg[877]  ( .D(start_in[876]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[877]) );
  DFF \start_reg_reg[878]  ( .D(start_in[877]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[878]) );
  DFF \start_reg_reg[879]  ( .D(start_in[878]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[879]) );
  DFF \start_reg_reg[880]  ( .D(start_in[879]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[880]) );
  DFF \start_reg_reg[881]  ( .D(start_in[880]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[881]) );
  DFF \start_reg_reg[882]  ( .D(start_in[881]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[882]) );
  DFF \start_reg_reg[883]  ( .D(start_in[882]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[883]) );
  DFF \start_reg_reg[884]  ( .D(start_in[883]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[884]) );
  DFF \start_reg_reg[885]  ( .D(start_in[884]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[885]) );
  DFF \start_reg_reg[886]  ( .D(start_in[885]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[886]) );
  DFF \start_reg_reg[887]  ( .D(start_in[886]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[887]) );
  DFF \start_reg_reg[888]  ( .D(start_in[887]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[888]) );
  DFF \start_reg_reg[889]  ( .D(start_in[888]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[889]) );
  DFF \start_reg_reg[890]  ( .D(start_in[889]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[890]) );
  DFF \start_reg_reg[891]  ( .D(start_in[890]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[891]) );
  DFF \start_reg_reg[892]  ( .D(start_in[891]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[892]) );
  DFF \start_reg_reg[893]  ( .D(start_in[892]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[893]) );
  DFF \start_reg_reg[894]  ( .D(start_in[893]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[894]) );
  DFF \start_reg_reg[895]  ( .D(start_in[894]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[895]) );
  DFF \start_reg_reg[896]  ( .D(start_in[895]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[896]) );
  DFF \start_reg_reg[897]  ( .D(start_in[896]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[897]) );
  DFF \start_reg_reg[898]  ( .D(start_in[897]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[898]) );
  DFF \start_reg_reg[899]  ( .D(start_in[898]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[899]) );
  DFF \start_reg_reg[900]  ( .D(start_in[899]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[900]) );
  DFF \start_reg_reg[901]  ( .D(start_in[900]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[901]) );
  DFF \start_reg_reg[902]  ( .D(start_in[901]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[902]) );
  DFF \start_reg_reg[903]  ( .D(start_in[902]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[903]) );
  DFF \start_reg_reg[904]  ( .D(start_in[903]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[904]) );
  DFF \start_reg_reg[905]  ( .D(start_in[904]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[905]) );
  DFF \start_reg_reg[906]  ( .D(start_in[905]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[906]) );
  DFF \start_reg_reg[907]  ( .D(start_in[906]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[907]) );
  DFF \start_reg_reg[908]  ( .D(start_in[907]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[908]) );
  DFF \start_reg_reg[909]  ( .D(start_in[908]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[909]) );
  DFF \start_reg_reg[910]  ( .D(start_in[909]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[910]) );
  DFF \start_reg_reg[911]  ( .D(start_in[910]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[911]) );
  DFF \start_reg_reg[912]  ( .D(start_in[911]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[912]) );
  DFF \start_reg_reg[913]  ( .D(start_in[912]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[913]) );
  DFF \start_reg_reg[914]  ( .D(start_in[913]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[914]) );
  DFF \start_reg_reg[915]  ( .D(start_in[914]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[915]) );
  DFF \start_reg_reg[916]  ( .D(start_in[915]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[916]) );
  DFF \start_reg_reg[917]  ( .D(start_in[916]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[917]) );
  DFF \start_reg_reg[918]  ( .D(start_in[917]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[918]) );
  DFF \start_reg_reg[919]  ( .D(start_in[918]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[919]) );
  DFF \start_reg_reg[920]  ( .D(start_in[919]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[920]) );
  DFF \start_reg_reg[921]  ( .D(start_in[920]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[921]) );
  DFF \start_reg_reg[922]  ( .D(start_in[921]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[922]) );
  DFF \start_reg_reg[923]  ( .D(start_in[922]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[923]) );
  DFF \start_reg_reg[924]  ( .D(start_in[923]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[924]) );
  DFF \start_reg_reg[925]  ( .D(start_in[924]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[925]) );
  DFF \start_reg_reg[926]  ( .D(start_in[925]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[926]) );
  DFF \start_reg_reg[927]  ( .D(start_in[926]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[927]) );
  DFF \start_reg_reg[928]  ( .D(start_in[927]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[928]) );
  DFF \start_reg_reg[929]  ( .D(start_in[928]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[929]) );
  DFF \start_reg_reg[930]  ( .D(start_in[929]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[930]) );
  DFF \start_reg_reg[931]  ( .D(start_in[930]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[931]) );
  DFF \start_reg_reg[932]  ( .D(start_in[931]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[932]) );
  DFF \start_reg_reg[933]  ( .D(start_in[932]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[933]) );
  DFF \start_reg_reg[934]  ( .D(start_in[933]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[934]) );
  DFF \start_reg_reg[935]  ( .D(start_in[934]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[935]) );
  DFF \start_reg_reg[936]  ( .D(start_in[935]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[936]) );
  DFF \start_reg_reg[937]  ( .D(start_in[936]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[937]) );
  DFF \start_reg_reg[938]  ( .D(start_in[937]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[938]) );
  DFF \start_reg_reg[939]  ( .D(start_in[938]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[939]) );
  DFF \start_reg_reg[940]  ( .D(start_in[939]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[940]) );
  DFF \start_reg_reg[941]  ( .D(start_in[940]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[941]) );
  DFF \start_reg_reg[942]  ( .D(start_in[941]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[942]) );
  DFF \start_reg_reg[943]  ( .D(start_in[942]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[943]) );
  DFF \start_reg_reg[944]  ( .D(start_in[943]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[944]) );
  DFF \start_reg_reg[945]  ( .D(start_in[944]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[945]) );
  DFF \start_reg_reg[946]  ( .D(start_in[945]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[946]) );
  DFF \start_reg_reg[947]  ( .D(start_in[946]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[947]) );
  DFF \start_reg_reg[948]  ( .D(start_in[947]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[948]) );
  DFF \start_reg_reg[949]  ( .D(start_in[948]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[949]) );
  DFF \start_reg_reg[950]  ( .D(start_in[949]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[950]) );
  DFF \start_reg_reg[951]  ( .D(start_in[950]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[951]) );
  DFF \start_reg_reg[952]  ( .D(start_in[951]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[952]) );
  DFF \start_reg_reg[953]  ( .D(start_in[952]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[953]) );
  DFF \start_reg_reg[954]  ( .D(start_in[953]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[954]) );
  DFF \start_reg_reg[955]  ( .D(start_in[954]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[955]) );
  DFF \start_reg_reg[956]  ( .D(start_in[955]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[956]) );
  DFF \start_reg_reg[957]  ( .D(start_in[956]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[957]) );
  DFF \start_reg_reg[958]  ( .D(start_in[957]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[958]) );
  DFF \start_reg_reg[959]  ( .D(start_in[958]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[959]) );
  DFF \start_reg_reg[960]  ( .D(start_in[959]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[960]) );
  DFF \start_reg_reg[961]  ( .D(start_in[960]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[961]) );
  DFF \start_reg_reg[962]  ( .D(start_in[961]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[962]) );
  DFF \start_reg_reg[963]  ( .D(start_in[962]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[963]) );
  DFF \start_reg_reg[964]  ( .D(start_in[963]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[964]) );
  DFF \start_reg_reg[965]  ( .D(start_in[964]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[965]) );
  DFF \start_reg_reg[966]  ( .D(start_in[965]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[966]) );
  DFF \start_reg_reg[967]  ( .D(start_in[966]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[967]) );
  DFF \start_reg_reg[968]  ( .D(start_in[967]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[968]) );
  DFF \start_reg_reg[969]  ( .D(start_in[968]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[969]) );
  DFF \start_reg_reg[970]  ( .D(start_in[969]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[970]) );
  DFF \start_reg_reg[971]  ( .D(start_in[970]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[971]) );
  DFF \start_reg_reg[972]  ( .D(start_in[971]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[972]) );
  DFF \start_reg_reg[973]  ( .D(start_in[972]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[973]) );
  DFF \start_reg_reg[974]  ( .D(start_in[973]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[974]) );
  DFF \start_reg_reg[975]  ( .D(start_in[974]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[975]) );
  DFF \start_reg_reg[976]  ( .D(start_in[975]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[976]) );
  DFF \start_reg_reg[977]  ( .D(start_in[976]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[977]) );
  DFF \start_reg_reg[978]  ( .D(start_in[977]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[978]) );
  DFF \start_reg_reg[979]  ( .D(start_in[978]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[979]) );
  DFF \start_reg_reg[980]  ( .D(start_in[979]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[980]) );
  DFF \start_reg_reg[981]  ( .D(start_in[980]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[981]) );
  DFF \start_reg_reg[982]  ( .D(start_in[981]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[982]) );
  DFF \start_reg_reg[983]  ( .D(start_in[982]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[983]) );
  DFF \start_reg_reg[984]  ( .D(start_in[983]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[984]) );
  DFF \start_reg_reg[985]  ( .D(start_in[984]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[985]) );
  DFF \start_reg_reg[986]  ( .D(start_in[985]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[986]) );
  DFF \start_reg_reg[987]  ( .D(start_in[986]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[987]) );
  DFF \start_reg_reg[988]  ( .D(start_in[987]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[988]) );
  DFF \start_reg_reg[989]  ( .D(start_in[988]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[989]) );
  DFF \start_reg_reg[990]  ( .D(start_in[989]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[990]) );
  DFF \start_reg_reg[991]  ( .D(start_in[990]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[991]) );
  DFF \start_reg_reg[992]  ( .D(start_in[991]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[992]) );
  DFF \start_reg_reg[993]  ( .D(start_in[992]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[993]) );
  DFF \start_reg_reg[994]  ( .D(start_in[993]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[994]) );
  DFF \start_reg_reg[995]  ( .D(start_in[994]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[995]) );
  DFF \start_reg_reg[996]  ( .D(start_in[995]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[996]) );
  DFF \start_reg_reg[997]  ( .D(start_in[996]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[997]) );
  DFF \start_reg_reg[998]  ( .D(start_in[997]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[998]) );
  DFF \start_reg_reg[999]  ( .D(start_in[998]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[999]) );
  DFF \start_reg_reg[1000]  ( .D(start_in[999]), .CLK(clk), .RST(rst), .I(1'b0), .Q(start_in[1000]) );
  DFF \start_reg_reg[1001]  ( .D(start_in[1000]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1001]) );
  DFF \start_reg_reg[1002]  ( .D(start_in[1001]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1002]) );
  DFF \start_reg_reg[1003]  ( .D(start_in[1002]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1003]) );
  DFF \start_reg_reg[1004]  ( .D(start_in[1003]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1004]) );
  DFF \start_reg_reg[1005]  ( .D(start_in[1004]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1005]) );
  DFF \start_reg_reg[1006]  ( .D(start_in[1005]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1006]) );
  DFF \start_reg_reg[1007]  ( .D(start_in[1006]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1007]) );
  DFF \start_reg_reg[1008]  ( .D(start_in[1007]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1008]) );
  DFF \start_reg_reg[1009]  ( .D(start_in[1008]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1009]) );
  DFF \start_reg_reg[1010]  ( .D(start_in[1009]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1010]) );
  DFF \start_reg_reg[1011]  ( .D(start_in[1010]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1011]) );
  DFF \start_reg_reg[1012]  ( .D(start_in[1011]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1012]) );
  DFF \start_reg_reg[1013]  ( .D(start_in[1012]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1013]) );
  DFF \start_reg_reg[1014]  ( .D(start_in[1013]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1014]) );
  DFF \start_reg_reg[1015]  ( .D(start_in[1014]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1015]) );
  DFF \start_reg_reg[1016]  ( .D(start_in[1015]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1016]) );
  DFF \start_reg_reg[1017]  ( .D(start_in[1016]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1017]) );
  DFF \start_reg_reg[1018]  ( .D(start_in[1017]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1018]) );
  DFF \start_reg_reg[1019]  ( .D(start_in[1018]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1019]) );
  DFF \start_reg_reg[1020]  ( .D(start_in[1019]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1020]) );
  DFF \start_reg_reg[1021]  ( .D(start_in[1020]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1021]) );
  DFF \start_reg_reg[1022]  ( .D(start_in[1021]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1022]) );
  DFF \start_reg_reg[1023]  ( .D(start_in[1022]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1023]) );
  DFF mul_pow_reg ( .D(n8), .CLK(clk), .RST(rst), .I(1'b0), .Q(mul_pow) );
  DFF \ereg_reg[0]  ( .D(ereg_next[0]), .CLK(clk), .RST(rst), .I(e_init[0]), 
        .Q(ein[0]) );
  DFF \ereg_reg[1]  ( .D(ereg_next[1]), .CLK(clk), .RST(rst), .I(e_init[1]), 
        .Q(ein[1]) );
  DFF \ereg_reg[2]  ( .D(ereg_next[2]), .CLK(clk), .RST(rst), .I(e_init[2]), 
        .Q(ein[2]) );
  DFF \ereg_reg[3]  ( .D(ereg_next[3]), .CLK(clk), .RST(rst), .I(e_init[3]), 
        .Q(ein[3]) );
  DFF \ereg_reg[4]  ( .D(ereg_next[4]), .CLK(clk), .RST(rst), .I(e_init[4]), 
        .Q(ein[4]) );
  DFF \ereg_reg[5]  ( .D(ereg_next[5]), .CLK(clk), .RST(rst), .I(e_init[5]), 
        .Q(ein[5]) );
  DFF \ereg_reg[6]  ( .D(ereg_next[6]), .CLK(clk), .RST(rst), .I(e_init[6]), 
        .Q(ein[6]) );
  DFF \ereg_reg[7]  ( .D(ereg_next[7]), .CLK(clk), .RST(rst), .I(e_init[7]), 
        .Q(ein[7]) );
  DFF \ereg_reg[8]  ( .D(ereg_next[8]), .CLK(clk), .RST(rst), .I(e_init[8]), 
        .Q(ein[8]) );
  DFF \ereg_reg[9]  ( .D(ereg_next[9]), .CLK(clk), .RST(rst), .I(e_init[9]), 
        .Q(ein[9]) );
  DFF \ereg_reg[10]  ( .D(ereg_next[10]), .CLK(clk), .RST(rst), .I(e_init[10]), 
        .Q(ein[10]) );
  DFF \ereg_reg[11]  ( .D(ereg_next[11]), .CLK(clk), .RST(rst), .I(e_init[11]), 
        .Q(ein[11]) );
  DFF \ereg_reg[12]  ( .D(ereg_next[12]), .CLK(clk), .RST(rst), .I(e_init[12]), 
        .Q(ein[12]) );
  DFF \ereg_reg[13]  ( .D(ereg_next[13]), .CLK(clk), .RST(rst), .I(e_init[13]), 
        .Q(ein[13]) );
  DFF \ereg_reg[14]  ( .D(ereg_next[14]), .CLK(clk), .RST(rst), .I(e_init[14]), 
        .Q(ein[14]) );
  DFF \ereg_reg[15]  ( .D(ereg_next[15]), .CLK(clk), .RST(rst), .I(e_init[15]), 
        .Q(ein[15]) );
  DFF \ereg_reg[16]  ( .D(ereg_next[16]), .CLK(clk), .RST(rst), .I(e_init[16]), 
        .Q(ein[16]) );
  DFF \ereg_reg[17]  ( .D(ereg_next[17]), .CLK(clk), .RST(rst), .I(e_init[17]), 
        .Q(ein[17]) );
  DFF \ereg_reg[18]  ( .D(ereg_next[18]), .CLK(clk), .RST(rst), .I(e_init[18]), 
        .Q(ein[18]) );
  DFF \ereg_reg[19]  ( .D(ereg_next[19]), .CLK(clk), .RST(rst), .I(e_init[19]), 
        .Q(ein[19]) );
  DFF \ereg_reg[20]  ( .D(ereg_next[20]), .CLK(clk), .RST(rst), .I(e_init[20]), 
        .Q(ein[20]) );
  DFF \ereg_reg[21]  ( .D(ereg_next[21]), .CLK(clk), .RST(rst), .I(e_init[21]), 
        .Q(ein[21]) );
  DFF \ereg_reg[22]  ( .D(ereg_next[22]), .CLK(clk), .RST(rst), .I(e_init[22]), 
        .Q(ein[22]) );
  DFF \ereg_reg[23]  ( .D(ereg_next[23]), .CLK(clk), .RST(rst), .I(e_init[23]), 
        .Q(ein[23]) );
  DFF \ereg_reg[24]  ( .D(ereg_next[24]), .CLK(clk), .RST(rst), .I(e_init[24]), 
        .Q(ein[24]) );
  DFF \ereg_reg[25]  ( .D(ereg_next[25]), .CLK(clk), .RST(rst), .I(e_init[25]), 
        .Q(ein[25]) );
  DFF \ereg_reg[26]  ( .D(ereg_next[26]), .CLK(clk), .RST(rst), .I(e_init[26]), 
        .Q(ein[26]) );
  DFF \ereg_reg[27]  ( .D(ereg_next[27]), .CLK(clk), .RST(rst), .I(e_init[27]), 
        .Q(ein[27]) );
  DFF \ereg_reg[28]  ( .D(ereg_next[28]), .CLK(clk), .RST(rst), .I(e_init[28]), 
        .Q(ein[28]) );
  DFF \ereg_reg[29]  ( .D(ereg_next[29]), .CLK(clk), .RST(rst), .I(e_init[29]), 
        .Q(ein[29]) );
  DFF \ereg_reg[30]  ( .D(ereg_next[30]), .CLK(clk), .RST(rst), .I(e_init[30]), 
        .Q(ein[30]) );
  DFF \ereg_reg[31]  ( .D(ereg_next[31]), .CLK(clk), .RST(rst), .I(e_init[31]), 
        .Q(ein[31]) );
  DFF \ereg_reg[32]  ( .D(ereg_next[32]), .CLK(clk), .RST(rst), .I(e_init[32]), 
        .Q(ein[32]) );
  DFF \ereg_reg[33]  ( .D(ereg_next[33]), .CLK(clk), .RST(rst), .I(e_init[33]), 
        .Q(ein[33]) );
  DFF \ereg_reg[34]  ( .D(ereg_next[34]), .CLK(clk), .RST(rst), .I(e_init[34]), 
        .Q(ein[34]) );
  DFF \ereg_reg[35]  ( .D(ereg_next[35]), .CLK(clk), .RST(rst), .I(e_init[35]), 
        .Q(ein[35]) );
  DFF \ereg_reg[36]  ( .D(ereg_next[36]), .CLK(clk), .RST(rst), .I(e_init[36]), 
        .Q(ein[36]) );
  DFF \ereg_reg[37]  ( .D(ereg_next[37]), .CLK(clk), .RST(rst), .I(e_init[37]), 
        .Q(ein[37]) );
  DFF \ereg_reg[38]  ( .D(ereg_next[38]), .CLK(clk), .RST(rst), .I(e_init[38]), 
        .Q(ein[38]) );
  DFF \ereg_reg[39]  ( .D(ereg_next[39]), .CLK(clk), .RST(rst), .I(e_init[39]), 
        .Q(ein[39]) );
  DFF \ereg_reg[40]  ( .D(ereg_next[40]), .CLK(clk), .RST(rst), .I(e_init[40]), 
        .Q(ein[40]) );
  DFF \ereg_reg[41]  ( .D(ereg_next[41]), .CLK(clk), .RST(rst), .I(e_init[41]), 
        .Q(ein[41]) );
  DFF \ereg_reg[42]  ( .D(ereg_next[42]), .CLK(clk), .RST(rst), .I(e_init[42]), 
        .Q(ein[42]) );
  DFF \ereg_reg[43]  ( .D(ereg_next[43]), .CLK(clk), .RST(rst), .I(e_init[43]), 
        .Q(ein[43]) );
  DFF \ereg_reg[44]  ( .D(ereg_next[44]), .CLK(clk), .RST(rst), .I(e_init[44]), 
        .Q(ein[44]) );
  DFF \ereg_reg[45]  ( .D(ereg_next[45]), .CLK(clk), .RST(rst), .I(e_init[45]), 
        .Q(ein[45]) );
  DFF \ereg_reg[46]  ( .D(ereg_next[46]), .CLK(clk), .RST(rst), .I(e_init[46]), 
        .Q(ein[46]) );
  DFF \ereg_reg[47]  ( .D(ereg_next[47]), .CLK(clk), .RST(rst), .I(e_init[47]), 
        .Q(ein[47]) );
  DFF \ereg_reg[48]  ( .D(ereg_next[48]), .CLK(clk), .RST(rst), .I(e_init[48]), 
        .Q(ein[48]) );
  DFF \ereg_reg[49]  ( .D(ereg_next[49]), .CLK(clk), .RST(rst), .I(e_init[49]), 
        .Q(ein[49]) );
  DFF \ereg_reg[50]  ( .D(ereg_next[50]), .CLK(clk), .RST(rst), .I(e_init[50]), 
        .Q(ein[50]) );
  DFF \ereg_reg[51]  ( .D(ereg_next[51]), .CLK(clk), .RST(rst), .I(e_init[51]), 
        .Q(ein[51]) );
  DFF \ereg_reg[52]  ( .D(ereg_next[52]), .CLK(clk), .RST(rst), .I(e_init[52]), 
        .Q(ein[52]) );
  DFF \ereg_reg[53]  ( .D(ereg_next[53]), .CLK(clk), .RST(rst), .I(e_init[53]), 
        .Q(ein[53]) );
  DFF \ereg_reg[54]  ( .D(ereg_next[54]), .CLK(clk), .RST(rst), .I(e_init[54]), 
        .Q(ein[54]) );
  DFF \ereg_reg[55]  ( .D(ereg_next[55]), .CLK(clk), .RST(rst), .I(e_init[55]), 
        .Q(ein[55]) );
  DFF \ereg_reg[56]  ( .D(ereg_next[56]), .CLK(clk), .RST(rst), .I(e_init[56]), 
        .Q(ein[56]) );
  DFF \ereg_reg[57]  ( .D(ereg_next[57]), .CLK(clk), .RST(rst), .I(e_init[57]), 
        .Q(ein[57]) );
  DFF \ereg_reg[58]  ( .D(ereg_next[58]), .CLK(clk), .RST(rst), .I(e_init[58]), 
        .Q(ein[58]) );
  DFF \ereg_reg[59]  ( .D(ereg_next[59]), .CLK(clk), .RST(rst), .I(e_init[59]), 
        .Q(ein[59]) );
  DFF \ereg_reg[60]  ( .D(ereg_next[60]), .CLK(clk), .RST(rst), .I(e_init[60]), 
        .Q(ein[60]) );
  DFF \ereg_reg[61]  ( .D(ereg_next[61]), .CLK(clk), .RST(rst), .I(e_init[61]), 
        .Q(ein[61]) );
  DFF \ereg_reg[62]  ( .D(ereg_next[62]), .CLK(clk), .RST(rst), .I(e_init[62]), 
        .Q(ein[62]) );
  DFF \ereg_reg[63]  ( .D(ereg_next[63]), .CLK(clk), .RST(rst), .I(e_init[63]), 
        .Q(ein[63]) );
  DFF \ereg_reg[64]  ( .D(ereg_next[64]), .CLK(clk), .RST(rst), .I(e_init[64]), 
        .Q(ein[64]) );
  DFF \ereg_reg[65]  ( .D(ereg_next[65]), .CLK(clk), .RST(rst), .I(e_init[65]), 
        .Q(ein[65]) );
  DFF \ereg_reg[66]  ( .D(ereg_next[66]), .CLK(clk), .RST(rst), .I(e_init[66]), 
        .Q(ein[66]) );
  DFF \ereg_reg[67]  ( .D(ereg_next[67]), .CLK(clk), .RST(rst), .I(e_init[67]), 
        .Q(ein[67]) );
  DFF \ereg_reg[68]  ( .D(ereg_next[68]), .CLK(clk), .RST(rst), .I(e_init[68]), 
        .Q(ein[68]) );
  DFF \ereg_reg[69]  ( .D(ereg_next[69]), .CLK(clk), .RST(rst), .I(e_init[69]), 
        .Q(ein[69]) );
  DFF \ereg_reg[70]  ( .D(ereg_next[70]), .CLK(clk), .RST(rst), .I(e_init[70]), 
        .Q(ein[70]) );
  DFF \ereg_reg[71]  ( .D(ereg_next[71]), .CLK(clk), .RST(rst), .I(e_init[71]), 
        .Q(ein[71]) );
  DFF \ereg_reg[72]  ( .D(ereg_next[72]), .CLK(clk), .RST(rst), .I(e_init[72]), 
        .Q(ein[72]) );
  DFF \ereg_reg[73]  ( .D(ereg_next[73]), .CLK(clk), .RST(rst), .I(e_init[73]), 
        .Q(ein[73]) );
  DFF \ereg_reg[74]  ( .D(ereg_next[74]), .CLK(clk), .RST(rst), .I(e_init[74]), 
        .Q(ein[74]) );
  DFF \ereg_reg[75]  ( .D(ereg_next[75]), .CLK(clk), .RST(rst), .I(e_init[75]), 
        .Q(ein[75]) );
  DFF \ereg_reg[76]  ( .D(ereg_next[76]), .CLK(clk), .RST(rst), .I(e_init[76]), 
        .Q(ein[76]) );
  DFF \ereg_reg[77]  ( .D(ereg_next[77]), .CLK(clk), .RST(rst), .I(e_init[77]), 
        .Q(ein[77]) );
  DFF \ereg_reg[78]  ( .D(ereg_next[78]), .CLK(clk), .RST(rst), .I(e_init[78]), 
        .Q(ein[78]) );
  DFF \ereg_reg[79]  ( .D(ereg_next[79]), .CLK(clk), .RST(rst), .I(e_init[79]), 
        .Q(ein[79]) );
  DFF \ereg_reg[80]  ( .D(ereg_next[80]), .CLK(clk), .RST(rst), .I(e_init[80]), 
        .Q(ein[80]) );
  DFF \ereg_reg[81]  ( .D(ereg_next[81]), .CLK(clk), .RST(rst), .I(e_init[81]), 
        .Q(ein[81]) );
  DFF \ereg_reg[82]  ( .D(ereg_next[82]), .CLK(clk), .RST(rst), .I(e_init[82]), 
        .Q(ein[82]) );
  DFF \ereg_reg[83]  ( .D(ereg_next[83]), .CLK(clk), .RST(rst), .I(e_init[83]), 
        .Q(ein[83]) );
  DFF \ereg_reg[84]  ( .D(ereg_next[84]), .CLK(clk), .RST(rst), .I(e_init[84]), 
        .Q(ein[84]) );
  DFF \ereg_reg[85]  ( .D(ereg_next[85]), .CLK(clk), .RST(rst), .I(e_init[85]), 
        .Q(ein[85]) );
  DFF \ereg_reg[86]  ( .D(ereg_next[86]), .CLK(clk), .RST(rst), .I(e_init[86]), 
        .Q(ein[86]) );
  DFF \ereg_reg[87]  ( .D(ereg_next[87]), .CLK(clk), .RST(rst), .I(e_init[87]), 
        .Q(ein[87]) );
  DFF \ereg_reg[88]  ( .D(ereg_next[88]), .CLK(clk), .RST(rst), .I(e_init[88]), 
        .Q(ein[88]) );
  DFF \ereg_reg[89]  ( .D(ereg_next[89]), .CLK(clk), .RST(rst), .I(e_init[89]), 
        .Q(ein[89]) );
  DFF \ereg_reg[90]  ( .D(ereg_next[90]), .CLK(clk), .RST(rst), .I(e_init[90]), 
        .Q(ein[90]) );
  DFF \ereg_reg[91]  ( .D(ereg_next[91]), .CLK(clk), .RST(rst), .I(e_init[91]), 
        .Q(ein[91]) );
  DFF \ereg_reg[92]  ( .D(ereg_next[92]), .CLK(clk), .RST(rst), .I(e_init[92]), 
        .Q(ein[92]) );
  DFF \ereg_reg[93]  ( .D(ereg_next[93]), .CLK(clk), .RST(rst), .I(e_init[93]), 
        .Q(ein[93]) );
  DFF \ereg_reg[94]  ( .D(ereg_next[94]), .CLK(clk), .RST(rst), .I(e_init[94]), 
        .Q(ein[94]) );
  DFF \ereg_reg[95]  ( .D(ereg_next[95]), .CLK(clk), .RST(rst), .I(e_init[95]), 
        .Q(ein[95]) );
  DFF \ereg_reg[96]  ( .D(ereg_next[96]), .CLK(clk), .RST(rst), .I(e_init[96]), 
        .Q(ein[96]) );
  DFF \ereg_reg[97]  ( .D(ereg_next[97]), .CLK(clk), .RST(rst), .I(e_init[97]), 
        .Q(ein[97]) );
  DFF \ereg_reg[98]  ( .D(ereg_next[98]), .CLK(clk), .RST(rst), .I(e_init[98]), 
        .Q(ein[98]) );
  DFF \ereg_reg[99]  ( .D(ereg_next[99]), .CLK(clk), .RST(rst), .I(e_init[99]), 
        .Q(ein[99]) );
  DFF \ereg_reg[100]  ( .D(ereg_next[100]), .CLK(clk), .RST(rst), .I(
        e_init[100]), .Q(ein[100]) );
  DFF \ereg_reg[101]  ( .D(ereg_next[101]), .CLK(clk), .RST(rst), .I(
        e_init[101]), .Q(ein[101]) );
  DFF \ereg_reg[102]  ( .D(ereg_next[102]), .CLK(clk), .RST(rst), .I(
        e_init[102]), .Q(ein[102]) );
  DFF \ereg_reg[103]  ( .D(ereg_next[103]), .CLK(clk), .RST(rst), .I(
        e_init[103]), .Q(ein[103]) );
  DFF \ereg_reg[104]  ( .D(ereg_next[104]), .CLK(clk), .RST(rst), .I(
        e_init[104]), .Q(ein[104]) );
  DFF \ereg_reg[105]  ( .D(ereg_next[105]), .CLK(clk), .RST(rst), .I(
        e_init[105]), .Q(ein[105]) );
  DFF \ereg_reg[106]  ( .D(ereg_next[106]), .CLK(clk), .RST(rst), .I(
        e_init[106]), .Q(ein[106]) );
  DFF \ereg_reg[107]  ( .D(ereg_next[107]), .CLK(clk), .RST(rst), .I(
        e_init[107]), .Q(ein[107]) );
  DFF \ereg_reg[108]  ( .D(ereg_next[108]), .CLK(clk), .RST(rst), .I(
        e_init[108]), .Q(ein[108]) );
  DFF \ereg_reg[109]  ( .D(ereg_next[109]), .CLK(clk), .RST(rst), .I(
        e_init[109]), .Q(ein[109]) );
  DFF \ereg_reg[110]  ( .D(ereg_next[110]), .CLK(clk), .RST(rst), .I(
        e_init[110]), .Q(ein[110]) );
  DFF \ereg_reg[111]  ( .D(ereg_next[111]), .CLK(clk), .RST(rst), .I(
        e_init[111]), .Q(ein[111]) );
  DFF \ereg_reg[112]  ( .D(ereg_next[112]), .CLK(clk), .RST(rst), .I(
        e_init[112]), .Q(ein[112]) );
  DFF \ereg_reg[113]  ( .D(ereg_next[113]), .CLK(clk), .RST(rst), .I(
        e_init[113]), .Q(ein[113]) );
  DFF \ereg_reg[114]  ( .D(ereg_next[114]), .CLK(clk), .RST(rst), .I(
        e_init[114]), .Q(ein[114]) );
  DFF \ereg_reg[115]  ( .D(ereg_next[115]), .CLK(clk), .RST(rst), .I(
        e_init[115]), .Q(ein[115]) );
  DFF \ereg_reg[116]  ( .D(ereg_next[116]), .CLK(clk), .RST(rst), .I(
        e_init[116]), .Q(ein[116]) );
  DFF \ereg_reg[117]  ( .D(ereg_next[117]), .CLK(clk), .RST(rst), .I(
        e_init[117]), .Q(ein[117]) );
  DFF \ereg_reg[118]  ( .D(ereg_next[118]), .CLK(clk), .RST(rst), .I(
        e_init[118]), .Q(ein[118]) );
  DFF \ereg_reg[119]  ( .D(ereg_next[119]), .CLK(clk), .RST(rst), .I(
        e_init[119]), .Q(ein[119]) );
  DFF \ereg_reg[120]  ( .D(ereg_next[120]), .CLK(clk), .RST(rst), .I(
        e_init[120]), .Q(ein[120]) );
  DFF \ereg_reg[121]  ( .D(ereg_next[121]), .CLK(clk), .RST(rst), .I(
        e_init[121]), .Q(ein[121]) );
  DFF \ereg_reg[122]  ( .D(ereg_next[122]), .CLK(clk), .RST(rst), .I(
        e_init[122]), .Q(ein[122]) );
  DFF \ereg_reg[123]  ( .D(ereg_next[123]), .CLK(clk), .RST(rst), .I(
        e_init[123]), .Q(ein[123]) );
  DFF \ereg_reg[124]  ( .D(ereg_next[124]), .CLK(clk), .RST(rst), .I(
        e_init[124]), .Q(ein[124]) );
  DFF \ereg_reg[125]  ( .D(ereg_next[125]), .CLK(clk), .RST(rst), .I(
        e_init[125]), .Q(ein[125]) );
  DFF \ereg_reg[126]  ( .D(ereg_next[126]), .CLK(clk), .RST(rst), .I(
        e_init[126]), .Q(ein[126]) );
  DFF \ereg_reg[127]  ( .D(ereg_next[127]), .CLK(clk), .RST(rst), .I(
        e_init[127]), .Q(ein[127]) );
  DFF \ereg_reg[128]  ( .D(ereg_next[128]), .CLK(clk), .RST(rst), .I(
        e_init[128]), .Q(ein[128]) );
  DFF \ereg_reg[129]  ( .D(ereg_next[129]), .CLK(clk), .RST(rst), .I(
        e_init[129]), .Q(ein[129]) );
  DFF \ereg_reg[130]  ( .D(ereg_next[130]), .CLK(clk), .RST(rst), .I(
        e_init[130]), .Q(ein[130]) );
  DFF \ereg_reg[131]  ( .D(ereg_next[131]), .CLK(clk), .RST(rst), .I(
        e_init[131]), .Q(ein[131]) );
  DFF \ereg_reg[132]  ( .D(ereg_next[132]), .CLK(clk), .RST(rst), .I(
        e_init[132]), .Q(ein[132]) );
  DFF \ereg_reg[133]  ( .D(ereg_next[133]), .CLK(clk), .RST(rst), .I(
        e_init[133]), .Q(ein[133]) );
  DFF \ereg_reg[134]  ( .D(ereg_next[134]), .CLK(clk), .RST(rst), .I(
        e_init[134]), .Q(ein[134]) );
  DFF \ereg_reg[135]  ( .D(ereg_next[135]), .CLK(clk), .RST(rst), .I(
        e_init[135]), .Q(ein[135]) );
  DFF \ereg_reg[136]  ( .D(ereg_next[136]), .CLK(clk), .RST(rst), .I(
        e_init[136]), .Q(ein[136]) );
  DFF \ereg_reg[137]  ( .D(ereg_next[137]), .CLK(clk), .RST(rst), .I(
        e_init[137]), .Q(ein[137]) );
  DFF \ereg_reg[138]  ( .D(ereg_next[138]), .CLK(clk), .RST(rst), .I(
        e_init[138]), .Q(ein[138]) );
  DFF \ereg_reg[139]  ( .D(ereg_next[139]), .CLK(clk), .RST(rst), .I(
        e_init[139]), .Q(ein[139]) );
  DFF \ereg_reg[140]  ( .D(ereg_next[140]), .CLK(clk), .RST(rst), .I(
        e_init[140]), .Q(ein[140]) );
  DFF \ereg_reg[141]  ( .D(ereg_next[141]), .CLK(clk), .RST(rst), .I(
        e_init[141]), .Q(ein[141]) );
  DFF \ereg_reg[142]  ( .D(ereg_next[142]), .CLK(clk), .RST(rst), .I(
        e_init[142]), .Q(ein[142]) );
  DFF \ereg_reg[143]  ( .D(ereg_next[143]), .CLK(clk), .RST(rst), .I(
        e_init[143]), .Q(ein[143]) );
  DFF \ereg_reg[144]  ( .D(ereg_next[144]), .CLK(clk), .RST(rst), .I(
        e_init[144]), .Q(ein[144]) );
  DFF \ereg_reg[145]  ( .D(ereg_next[145]), .CLK(clk), .RST(rst), .I(
        e_init[145]), .Q(ein[145]) );
  DFF \ereg_reg[146]  ( .D(ereg_next[146]), .CLK(clk), .RST(rst), .I(
        e_init[146]), .Q(ein[146]) );
  DFF \ereg_reg[147]  ( .D(ereg_next[147]), .CLK(clk), .RST(rst), .I(
        e_init[147]), .Q(ein[147]) );
  DFF \ereg_reg[148]  ( .D(ereg_next[148]), .CLK(clk), .RST(rst), .I(
        e_init[148]), .Q(ein[148]) );
  DFF \ereg_reg[149]  ( .D(ereg_next[149]), .CLK(clk), .RST(rst), .I(
        e_init[149]), .Q(ein[149]) );
  DFF \ereg_reg[150]  ( .D(ereg_next[150]), .CLK(clk), .RST(rst), .I(
        e_init[150]), .Q(ein[150]) );
  DFF \ereg_reg[151]  ( .D(ereg_next[151]), .CLK(clk), .RST(rst), .I(
        e_init[151]), .Q(ein[151]) );
  DFF \ereg_reg[152]  ( .D(ereg_next[152]), .CLK(clk), .RST(rst), .I(
        e_init[152]), .Q(ein[152]) );
  DFF \ereg_reg[153]  ( .D(ereg_next[153]), .CLK(clk), .RST(rst), .I(
        e_init[153]), .Q(ein[153]) );
  DFF \ereg_reg[154]  ( .D(ereg_next[154]), .CLK(clk), .RST(rst), .I(
        e_init[154]), .Q(ein[154]) );
  DFF \ereg_reg[155]  ( .D(ereg_next[155]), .CLK(clk), .RST(rst), .I(
        e_init[155]), .Q(ein[155]) );
  DFF \ereg_reg[156]  ( .D(ereg_next[156]), .CLK(clk), .RST(rst), .I(
        e_init[156]), .Q(ein[156]) );
  DFF \ereg_reg[157]  ( .D(ereg_next[157]), .CLK(clk), .RST(rst), .I(
        e_init[157]), .Q(ein[157]) );
  DFF \ereg_reg[158]  ( .D(ereg_next[158]), .CLK(clk), .RST(rst), .I(
        e_init[158]), .Q(ein[158]) );
  DFF \ereg_reg[159]  ( .D(ereg_next[159]), .CLK(clk), .RST(rst), .I(
        e_init[159]), .Q(ein[159]) );
  DFF \ereg_reg[160]  ( .D(ereg_next[160]), .CLK(clk), .RST(rst), .I(
        e_init[160]), .Q(ein[160]) );
  DFF \ereg_reg[161]  ( .D(ereg_next[161]), .CLK(clk), .RST(rst), .I(
        e_init[161]), .Q(ein[161]) );
  DFF \ereg_reg[162]  ( .D(ereg_next[162]), .CLK(clk), .RST(rst), .I(
        e_init[162]), .Q(ein[162]) );
  DFF \ereg_reg[163]  ( .D(ereg_next[163]), .CLK(clk), .RST(rst), .I(
        e_init[163]), .Q(ein[163]) );
  DFF \ereg_reg[164]  ( .D(ereg_next[164]), .CLK(clk), .RST(rst), .I(
        e_init[164]), .Q(ein[164]) );
  DFF \ereg_reg[165]  ( .D(ereg_next[165]), .CLK(clk), .RST(rst), .I(
        e_init[165]), .Q(ein[165]) );
  DFF \ereg_reg[166]  ( .D(ereg_next[166]), .CLK(clk), .RST(rst), .I(
        e_init[166]), .Q(ein[166]) );
  DFF \ereg_reg[167]  ( .D(ereg_next[167]), .CLK(clk), .RST(rst), .I(
        e_init[167]), .Q(ein[167]) );
  DFF \ereg_reg[168]  ( .D(ereg_next[168]), .CLK(clk), .RST(rst), .I(
        e_init[168]), .Q(ein[168]) );
  DFF \ereg_reg[169]  ( .D(ereg_next[169]), .CLK(clk), .RST(rst), .I(
        e_init[169]), .Q(ein[169]) );
  DFF \ereg_reg[170]  ( .D(ereg_next[170]), .CLK(clk), .RST(rst), .I(
        e_init[170]), .Q(ein[170]) );
  DFF \ereg_reg[171]  ( .D(ereg_next[171]), .CLK(clk), .RST(rst), .I(
        e_init[171]), .Q(ein[171]) );
  DFF \ereg_reg[172]  ( .D(ereg_next[172]), .CLK(clk), .RST(rst), .I(
        e_init[172]), .Q(ein[172]) );
  DFF \ereg_reg[173]  ( .D(ereg_next[173]), .CLK(clk), .RST(rst), .I(
        e_init[173]), .Q(ein[173]) );
  DFF \ereg_reg[174]  ( .D(ereg_next[174]), .CLK(clk), .RST(rst), .I(
        e_init[174]), .Q(ein[174]) );
  DFF \ereg_reg[175]  ( .D(ereg_next[175]), .CLK(clk), .RST(rst), .I(
        e_init[175]), .Q(ein[175]) );
  DFF \ereg_reg[176]  ( .D(ereg_next[176]), .CLK(clk), .RST(rst), .I(
        e_init[176]), .Q(ein[176]) );
  DFF \ereg_reg[177]  ( .D(ereg_next[177]), .CLK(clk), .RST(rst), .I(
        e_init[177]), .Q(ein[177]) );
  DFF \ereg_reg[178]  ( .D(ereg_next[178]), .CLK(clk), .RST(rst), .I(
        e_init[178]), .Q(ein[178]) );
  DFF \ereg_reg[179]  ( .D(ereg_next[179]), .CLK(clk), .RST(rst), .I(
        e_init[179]), .Q(ein[179]) );
  DFF \ereg_reg[180]  ( .D(ereg_next[180]), .CLK(clk), .RST(rst), .I(
        e_init[180]), .Q(ein[180]) );
  DFF \ereg_reg[181]  ( .D(ereg_next[181]), .CLK(clk), .RST(rst), .I(
        e_init[181]), .Q(ein[181]) );
  DFF \ereg_reg[182]  ( .D(ereg_next[182]), .CLK(clk), .RST(rst), .I(
        e_init[182]), .Q(ein[182]) );
  DFF \ereg_reg[183]  ( .D(ereg_next[183]), .CLK(clk), .RST(rst), .I(
        e_init[183]), .Q(ein[183]) );
  DFF \ereg_reg[184]  ( .D(ereg_next[184]), .CLK(clk), .RST(rst), .I(
        e_init[184]), .Q(ein[184]) );
  DFF \ereg_reg[185]  ( .D(ereg_next[185]), .CLK(clk), .RST(rst), .I(
        e_init[185]), .Q(ein[185]) );
  DFF \ereg_reg[186]  ( .D(ereg_next[186]), .CLK(clk), .RST(rst), .I(
        e_init[186]), .Q(ein[186]) );
  DFF \ereg_reg[187]  ( .D(ereg_next[187]), .CLK(clk), .RST(rst), .I(
        e_init[187]), .Q(ein[187]) );
  DFF \ereg_reg[188]  ( .D(ereg_next[188]), .CLK(clk), .RST(rst), .I(
        e_init[188]), .Q(ein[188]) );
  DFF \ereg_reg[189]  ( .D(ereg_next[189]), .CLK(clk), .RST(rst), .I(
        e_init[189]), .Q(ein[189]) );
  DFF \ereg_reg[190]  ( .D(ereg_next[190]), .CLK(clk), .RST(rst), .I(
        e_init[190]), .Q(ein[190]) );
  DFF \ereg_reg[191]  ( .D(ereg_next[191]), .CLK(clk), .RST(rst), .I(
        e_init[191]), .Q(ein[191]) );
  DFF \ereg_reg[192]  ( .D(ereg_next[192]), .CLK(clk), .RST(rst), .I(
        e_init[192]), .Q(ein[192]) );
  DFF \ereg_reg[193]  ( .D(ereg_next[193]), .CLK(clk), .RST(rst), .I(
        e_init[193]), .Q(ein[193]) );
  DFF \ereg_reg[194]  ( .D(ereg_next[194]), .CLK(clk), .RST(rst), .I(
        e_init[194]), .Q(ein[194]) );
  DFF \ereg_reg[195]  ( .D(ereg_next[195]), .CLK(clk), .RST(rst), .I(
        e_init[195]), .Q(ein[195]) );
  DFF \ereg_reg[196]  ( .D(ereg_next[196]), .CLK(clk), .RST(rst), .I(
        e_init[196]), .Q(ein[196]) );
  DFF \ereg_reg[197]  ( .D(ereg_next[197]), .CLK(clk), .RST(rst), .I(
        e_init[197]), .Q(ein[197]) );
  DFF \ereg_reg[198]  ( .D(ereg_next[198]), .CLK(clk), .RST(rst), .I(
        e_init[198]), .Q(ein[198]) );
  DFF \ereg_reg[199]  ( .D(ereg_next[199]), .CLK(clk), .RST(rst), .I(
        e_init[199]), .Q(ein[199]) );
  DFF \ereg_reg[200]  ( .D(ereg_next[200]), .CLK(clk), .RST(rst), .I(
        e_init[200]), .Q(ein[200]) );
  DFF \ereg_reg[201]  ( .D(ereg_next[201]), .CLK(clk), .RST(rst), .I(
        e_init[201]), .Q(ein[201]) );
  DFF \ereg_reg[202]  ( .D(ereg_next[202]), .CLK(clk), .RST(rst), .I(
        e_init[202]), .Q(ein[202]) );
  DFF \ereg_reg[203]  ( .D(ereg_next[203]), .CLK(clk), .RST(rst), .I(
        e_init[203]), .Q(ein[203]) );
  DFF \ereg_reg[204]  ( .D(ereg_next[204]), .CLK(clk), .RST(rst), .I(
        e_init[204]), .Q(ein[204]) );
  DFF \ereg_reg[205]  ( .D(ereg_next[205]), .CLK(clk), .RST(rst), .I(
        e_init[205]), .Q(ein[205]) );
  DFF \ereg_reg[206]  ( .D(ereg_next[206]), .CLK(clk), .RST(rst), .I(
        e_init[206]), .Q(ein[206]) );
  DFF \ereg_reg[207]  ( .D(ereg_next[207]), .CLK(clk), .RST(rst), .I(
        e_init[207]), .Q(ein[207]) );
  DFF \ereg_reg[208]  ( .D(ereg_next[208]), .CLK(clk), .RST(rst), .I(
        e_init[208]), .Q(ein[208]) );
  DFF \ereg_reg[209]  ( .D(ereg_next[209]), .CLK(clk), .RST(rst), .I(
        e_init[209]), .Q(ein[209]) );
  DFF \ereg_reg[210]  ( .D(ereg_next[210]), .CLK(clk), .RST(rst), .I(
        e_init[210]), .Q(ein[210]) );
  DFF \ereg_reg[211]  ( .D(ereg_next[211]), .CLK(clk), .RST(rst), .I(
        e_init[211]), .Q(ein[211]) );
  DFF \ereg_reg[212]  ( .D(ereg_next[212]), .CLK(clk), .RST(rst), .I(
        e_init[212]), .Q(ein[212]) );
  DFF \ereg_reg[213]  ( .D(ereg_next[213]), .CLK(clk), .RST(rst), .I(
        e_init[213]), .Q(ein[213]) );
  DFF \ereg_reg[214]  ( .D(ereg_next[214]), .CLK(clk), .RST(rst), .I(
        e_init[214]), .Q(ein[214]) );
  DFF \ereg_reg[215]  ( .D(ereg_next[215]), .CLK(clk), .RST(rst), .I(
        e_init[215]), .Q(ein[215]) );
  DFF \ereg_reg[216]  ( .D(ereg_next[216]), .CLK(clk), .RST(rst), .I(
        e_init[216]), .Q(ein[216]) );
  DFF \ereg_reg[217]  ( .D(ereg_next[217]), .CLK(clk), .RST(rst), .I(
        e_init[217]), .Q(ein[217]) );
  DFF \ereg_reg[218]  ( .D(ereg_next[218]), .CLK(clk), .RST(rst), .I(
        e_init[218]), .Q(ein[218]) );
  DFF \ereg_reg[219]  ( .D(ereg_next[219]), .CLK(clk), .RST(rst), .I(
        e_init[219]), .Q(ein[219]) );
  DFF \ereg_reg[220]  ( .D(ereg_next[220]), .CLK(clk), .RST(rst), .I(
        e_init[220]), .Q(ein[220]) );
  DFF \ereg_reg[221]  ( .D(ereg_next[221]), .CLK(clk), .RST(rst), .I(
        e_init[221]), .Q(ein[221]) );
  DFF \ereg_reg[222]  ( .D(ereg_next[222]), .CLK(clk), .RST(rst), .I(
        e_init[222]), .Q(ein[222]) );
  DFF \ereg_reg[223]  ( .D(ereg_next[223]), .CLK(clk), .RST(rst), .I(
        e_init[223]), .Q(ein[223]) );
  DFF \ereg_reg[224]  ( .D(ereg_next[224]), .CLK(clk), .RST(rst), .I(
        e_init[224]), .Q(ein[224]) );
  DFF \ereg_reg[225]  ( .D(ereg_next[225]), .CLK(clk), .RST(rst), .I(
        e_init[225]), .Q(ein[225]) );
  DFF \ereg_reg[226]  ( .D(ereg_next[226]), .CLK(clk), .RST(rst), .I(
        e_init[226]), .Q(ein[226]) );
  DFF \ereg_reg[227]  ( .D(ereg_next[227]), .CLK(clk), .RST(rst), .I(
        e_init[227]), .Q(ein[227]) );
  DFF \ereg_reg[228]  ( .D(ereg_next[228]), .CLK(clk), .RST(rst), .I(
        e_init[228]), .Q(ein[228]) );
  DFF \ereg_reg[229]  ( .D(ereg_next[229]), .CLK(clk), .RST(rst), .I(
        e_init[229]), .Q(ein[229]) );
  DFF \ereg_reg[230]  ( .D(ereg_next[230]), .CLK(clk), .RST(rst), .I(
        e_init[230]), .Q(ein[230]) );
  DFF \ereg_reg[231]  ( .D(ereg_next[231]), .CLK(clk), .RST(rst), .I(
        e_init[231]), .Q(ein[231]) );
  DFF \ereg_reg[232]  ( .D(ereg_next[232]), .CLK(clk), .RST(rst), .I(
        e_init[232]), .Q(ein[232]) );
  DFF \ereg_reg[233]  ( .D(ereg_next[233]), .CLK(clk), .RST(rst), .I(
        e_init[233]), .Q(ein[233]) );
  DFF \ereg_reg[234]  ( .D(ereg_next[234]), .CLK(clk), .RST(rst), .I(
        e_init[234]), .Q(ein[234]) );
  DFF \ereg_reg[235]  ( .D(ereg_next[235]), .CLK(clk), .RST(rst), .I(
        e_init[235]), .Q(ein[235]) );
  DFF \ereg_reg[236]  ( .D(ereg_next[236]), .CLK(clk), .RST(rst), .I(
        e_init[236]), .Q(ein[236]) );
  DFF \ereg_reg[237]  ( .D(ereg_next[237]), .CLK(clk), .RST(rst), .I(
        e_init[237]), .Q(ein[237]) );
  DFF \ereg_reg[238]  ( .D(ereg_next[238]), .CLK(clk), .RST(rst), .I(
        e_init[238]), .Q(ein[238]) );
  DFF \ereg_reg[239]  ( .D(ereg_next[239]), .CLK(clk), .RST(rst), .I(
        e_init[239]), .Q(ein[239]) );
  DFF \ereg_reg[240]  ( .D(ereg_next[240]), .CLK(clk), .RST(rst), .I(
        e_init[240]), .Q(ein[240]) );
  DFF \ereg_reg[241]  ( .D(ereg_next[241]), .CLK(clk), .RST(rst), .I(
        e_init[241]), .Q(ein[241]) );
  DFF \ereg_reg[242]  ( .D(ereg_next[242]), .CLK(clk), .RST(rst), .I(
        e_init[242]), .Q(ein[242]) );
  DFF \ereg_reg[243]  ( .D(ereg_next[243]), .CLK(clk), .RST(rst), .I(
        e_init[243]), .Q(ein[243]) );
  DFF \ereg_reg[244]  ( .D(ereg_next[244]), .CLK(clk), .RST(rst), .I(
        e_init[244]), .Q(ein[244]) );
  DFF \ereg_reg[245]  ( .D(ereg_next[245]), .CLK(clk), .RST(rst), .I(
        e_init[245]), .Q(ein[245]) );
  DFF \ereg_reg[246]  ( .D(ereg_next[246]), .CLK(clk), .RST(rst), .I(
        e_init[246]), .Q(ein[246]) );
  DFF \ereg_reg[247]  ( .D(ereg_next[247]), .CLK(clk), .RST(rst), .I(
        e_init[247]), .Q(ein[247]) );
  DFF \ereg_reg[248]  ( .D(ereg_next[248]), .CLK(clk), .RST(rst), .I(
        e_init[248]), .Q(ein[248]) );
  DFF \ereg_reg[249]  ( .D(ereg_next[249]), .CLK(clk), .RST(rst), .I(
        e_init[249]), .Q(ein[249]) );
  DFF \ereg_reg[250]  ( .D(ereg_next[250]), .CLK(clk), .RST(rst), .I(
        e_init[250]), .Q(ein[250]) );
  DFF \ereg_reg[251]  ( .D(ereg_next[251]), .CLK(clk), .RST(rst), .I(
        e_init[251]), .Q(ein[251]) );
  DFF \ereg_reg[252]  ( .D(ereg_next[252]), .CLK(clk), .RST(rst), .I(
        e_init[252]), .Q(ein[252]) );
  DFF \ereg_reg[253]  ( .D(ereg_next[253]), .CLK(clk), .RST(rst), .I(
        e_init[253]), .Q(ein[253]) );
  DFF \ereg_reg[254]  ( .D(ereg_next[254]), .CLK(clk), .RST(rst), .I(
        e_init[254]), .Q(ein[254]) );
  DFF \ereg_reg[255]  ( .D(ereg_next[255]), .CLK(clk), .RST(rst), .I(
        e_init[255]), .Q(ein[255]) );
  DFF \ereg_reg[256]  ( .D(ereg_next[256]), .CLK(clk), .RST(rst), .I(
        e_init[256]), .Q(ein[256]) );
  DFF \ereg_reg[257]  ( .D(ereg_next[257]), .CLK(clk), .RST(rst), .I(
        e_init[257]), .Q(ein[257]) );
  DFF \ereg_reg[258]  ( .D(ereg_next[258]), .CLK(clk), .RST(rst), .I(
        e_init[258]), .Q(ein[258]) );
  DFF \ereg_reg[259]  ( .D(ereg_next[259]), .CLK(clk), .RST(rst), .I(
        e_init[259]), .Q(ein[259]) );
  DFF \ereg_reg[260]  ( .D(ereg_next[260]), .CLK(clk), .RST(rst), .I(
        e_init[260]), .Q(ein[260]) );
  DFF \ereg_reg[261]  ( .D(ereg_next[261]), .CLK(clk), .RST(rst), .I(
        e_init[261]), .Q(ein[261]) );
  DFF \ereg_reg[262]  ( .D(ereg_next[262]), .CLK(clk), .RST(rst), .I(
        e_init[262]), .Q(ein[262]) );
  DFF \ereg_reg[263]  ( .D(ereg_next[263]), .CLK(clk), .RST(rst), .I(
        e_init[263]), .Q(ein[263]) );
  DFF \ereg_reg[264]  ( .D(ereg_next[264]), .CLK(clk), .RST(rst), .I(
        e_init[264]), .Q(ein[264]) );
  DFF \ereg_reg[265]  ( .D(ereg_next[265]), .CLK(clk), .RST(rst), .I(
        e_init[265]), .Q(ein[265]) );
  DFF \ereg_reg[266]  ( .D(ereg_next[266]), .CLK(clk), .RST(rst), .I(
        e_init[266]), .Q(ein[266]) );
  DFF \ereg_reg[267]  ( .D(ereg_next[267]), .CLK(clk), .RST(rst), .I(
        e_init[267]), .Q(ein[267]) );
  DFF \ereg_reg[268]  ( .D(ereg_next[268]), .CLK(clk), .RST(rst), .I(
        e_init[268]), .Q(ein[268]) );
  DFF \ereg_reg[269]  ( .D(ereg_next[269]), .CLK(clk), .RST(rst), .I(
        e_init[269]), .Q(ein[269]) );
  DFF \ereg_reg[270]  ( .D(ereg_next[270]), .CLK(clk), .RST(rst), .I(
        e_init[270]), .Q(ein[270]) );
  DFF \ereg_reg[271]  ( .D(ereg_next[271]), .CLK(clk), .RST(rst), .I(
        e_init[271]), .Q(ein[271]) );
  DFF \ereg_reg[272]  ( .D(ereg_next[272]), .CLK(clk), .RST(rst), .I(
        e_init[272]), .Q(ein[272]) );
  DFF \ereg_reg[273]  ( .D(ereg_next[273]), .CLK(clk), .RST(rst), .I(
        e_init[273]), .Q(ein[273]) );
  DFF \ereg_reg[274]  ( .D(ereg_next[274]), .CLK(clk), .RST(rst), .I(
        e_init[274]), .Q(ein[274]) );
  DFF \ereg_reg[275]  ( .D(ereg_next[275]), .CLK(clk), .RST(rst), .I(
        e_init[275]), .Q(ein[275]) );
  DFF \ereg_reg[276]  ( .D(ereg_next[276]), .CLK(clk), .RST(rst), .I(
        e_init[276]), .Q(ein[276]) );
  DFF \ereg_reg[277]  ( .D(ereg_next[277]), .CLK(clk), .RST(rst), .I(
        e_init[277]), .Q(ein[277]) );
  DFF \ereg_reg[278]  ( .D(ereg_next[278]), .CLK(clk), .RST(rst), .I(
        e_init[278]), .Q(ein[278]) );
  DFF \ereg_reg[279]  ( .D(ereg_next[279]), .CLK(clk), .RST(rst), .I(
        e_init[279]), .Q(ein[279]) );
  DFF \ereg_reg[280]  ( .D(ereg_next[280]), .CLK(clk), .RST(rst), .I(
        e_init[280]), .Q(ein[280]) );
  DFF \ereg_reg[281]  ( .D(ereg_next[281]), .CLK(clk), .RST(rst), .I(
        e_init[281]), .Q(ein[281]) );
  DFF \ereg_reg[282]  ( .D(ereg_next[282]), .CLK(clk), .RST(rst), .I(
        e_init[282]), .Q(ein[282]) );
  DFF \ereg_reg[283]  ( .D(ereg_next[283]), .CLK(clk), .RST(rst), .I(
        e_init[283]), .Q(ein[283]) );
  DFF \ereg_reg[284]  ( .D(ereg_next[284]), .CLK(clk), .RST(rst), .I(
        e_init[284]), .Q(ein[284]) );
  DFF \ereg_reg[285]  ( .D(ereg_next[285]), .CLK(clk), .RST(rst), .I(
        e_init[285]), .Q(ein[285]) );
  DFF \ereg_reg[286]  ( .D(ereg_next[286]), .CLK(clk), .RST(rst), .I(
        e_init[286]), .Q(ein[286]) );
  DFF \ereg_reg[287]  ( .D(ereg_next[287]), .CLK(clk), .RST(rst), .I(
        e_init[287]), .Q(ein[287]) );
  DFF \ereg_reg[288]  ( .D(ereg_next[288]), .CLK(clk), .RST(rst), .I(
        e_init[288]), .Q(ein[288]) );
  DFF \ereg_reg[289]  ( .D(ereg_next[289]), .CLK(clk), .RST(rst), .I(
        e_init[289]), .Q(ein[289]) );
  DFF \ereg_reg[290]  ( .D(ereg_next[290]), .CLK(clk), .RST(rst), .I(
        e_init[290]), .Q(ein[290]) );
  DFF \ereg_reg[291]  ( .D(ereg_next[291]), .CLK(clk), .RST(rst), .I(
        e_init[291]), .Q(ein[291]) );
  DFF \ereg_reg[292]  ( .D(ereg_next[292]), .CLK(clk), .RST(rst), .I(
        e_init[292]), .Q(ein[292]) );
  DFF \ereg_reg[293]  ( .D(ereg_next[293]), .CLK(clk), .RST(rst), .I(
        e_init[293]), .Q(ein[293]) );
  DFF \ereg_reg[294]  ( .D(ereg_next[294]), .CLK(clk), .RST(rst), .I(
        e_init[294]), .Q(ein[294]) );
  DFF \ereg_reg[295]  ( .D(ereg_next[295]), .CLK(clk), .RST(rst), .I(
        e_init[295]), .Q(ein[295]) );
  DFF \ereg_reg[296]  ( .D(ereg_next[296]), .CLK(clk), .RST(rst), .I(
        e_init[296]), .Q(ein[296]) );
  DFF \ereg_reg[297]  ( .D(ereg_next[297]), .CLK(clk), .RST(rst), .I(
        e_init[297]), .Q(ein[297]) );
  DFF \ereg_reg[298]  ( .D(ereg_next[298]), .CLK(clk), .RST(rst), .I(
        e_init[298]), .Q(ein[298]) );
  DFF \ereg_reg[299]  ( .D(ereg_next[299]), .CLK(clk), .RST(rst), .I(
        e_init[299]), .Q(ein[299]) );
  DFF \ereg_reg[300]  ( .D(ereg_next[300]), .CLK(clk), .RST(rst), .I(
        e_init[300]), .Q(ein[300]) );
  DFF \ereg_reg[301]  ( .D(ereg_next[301]), .CLK(clk), .RST(rst), .I(
        e_init[301]), .Q(ein[301]) );
  DFF \ereg_reg[302]  ( .D(ereg_next[302]), .CLK(clk), .RST(rst), .I(
        e_init[302]), .Q(ein[302]) );
  DFF \ereg_reg[303]  ( .D(ereg_next[303]), .CLK(clk), .RST(rst), .I(
        e_init[303]), .Q(ein[303]) );
  DFF \ereg_reg[304]  ( .D(ereg_next[304]), .CLK(clk), .RST(rst), .I(
        e_init[304]), .Q(ein[304]) );
  DFF \ereg_reg[305]  ( .D(ereg_next[305]), .CLK(clk), .RST(rst), .I(
        e_init[305]), .Q(ein[305]) );
  DFF \ereg_reg[306]  ( .D(ereg_next[306]), .CLK(clk), .RST(rst), .I(
        e_init[306]), .Q(ein[306]) );
  DFF \ereg_reg[307]  ( .D(ereg_next[307]), .CLK(clk), .RST(rst), .I(
        e_init[307]), .Q(ein[307]) );
  DFF \ereg_reg[308]  ( .D(ereg_next[308]), .CLK(clk), .RST(rst), .I(
        e_init[308]), .Q(ein[308]) );
  DFF \ereg_reg[309]  ( .D(ereg_next[309]), .CLK(clk), .RST(rst), .I(
        e_init[309]), .Q(ein[309]) );
  DFF \ereg_reg[310]  ( .D(ereg_next[310]), .CLK(clk), .RST(rst), .I(
        e_init[310]), .Q(ein[310]) );
  DFF \ereg_reg[311]  ( .D(ereg_next[311]), .CLK(clk), .RST(rst), .I(
        e_init[311]), .Q(ein[311]) );
  DFF \ereg_reg[312]  ( .D(ereg_next[312]), .CLK(clk), .RST(rst), .I(
        e_init[312]), .Q(ein[312]) );
  DFF \ereg_reg[313]  ( .D(ereg_next[313]), .CLK(clk), .RST(rst), .I(
        e_init[313]), .Q(ein[313]) );
  DFF \ereg_reg[314]  ( .D(ereg_next[314]), .CLK(clk), .RST(rst), .I(
        e_init[314]), .Q(ein[314]) );
  DFF \ereg_reg[315]  ( .D(ereg_next[315]), .CLK(clk), .RST(rst), .I(
        e_init[315]), .Q(ein[315]) );
  DFF \ereg_reg[316]  ( .D(ereg_next[316]), .CLK(clk), .RST(rst), .I(
        e_init[316]), .Q(ein[316]) );
  DFF \ereg_reg[317]  ( .D(ereg_next[317]), .CLK(clk), .RST(rst), .I(
        e_init[317]), .Q(ein[317]) );
  DFF \ereg_reg[318]  ( .D(ereg_next[318]), .CLK(clk), .RST(rst), .I(
        e_init[318]), .Q(ein[318]) );
  DFF \ereg_reg[319]  ( .D(ereg_next[319]), .CLK(clk), .RST(rst), .I(
        e_init[319]), .Q(ein[319]) );
  DFF \ereg_reg[320]  ( .D(ereg_next[320]), .CLK(clk), .RST(rst), .I(
        e_init[320]), .Q(ein[320]) );
  DFF \ereg_reg[321]  ( .D(ereg_next[321]), .CLK(clk), .RST(rst), .I(
        e_init[321]), .Q(ein[321]) );
  DFF \ereg_reg[322]  ( .D(ereg_next[322]), .CLK(clk), .RST(rst), .I(
        e_init[322]), .Q(ein[322]) );
  DFF \ereg_reg[323]  ( .D(ereg_next[323]), .CLK(clk), .RST(rst), .I(
        e_init[323]), .Q(ein[323]) );
  DFF \ereg_reg[324]  ( .D(ereg_next[324]), .CLK(clk), .RST(rst), .I(
        e_init[324]), .Q(ein[324]) );
  DFF \ereg_reg[325]  ( .D(ereg_next[325]), .CLK(clk), .RST(rst), .I(
        e_init[325]), .Q(ein[325]) );
  DFF \ereg_reg[326]  ( .D(ereg_next[326]), .CLK(clk), .RST(rst), .I(
        e_init[326]), .Q(ein[326]) );
  DFF \ereg_reg[327]  ( .D(ereg_next[327]), .CLK(clk), .RST(rst), .I(
        e_init[327]), .Q(ein[327]) );
  DFF \ereg_reg[328]  ( .D(ereg_next[328]), .CLK(clk), .RST(rst), .I(
        e_init[328]), .Q(ein[328]) );
  DFF \ereg_reg[329]  ( .D(ereg_next[329]), .CLK(clk), .RST(rst), .I(
        e_init[329]), .Q(ein[329]) );
  DFF \ereg_reg[330]  ( .D(ereg_next[330]), .CLK(clk), .RST(rst), .I(
        e_init[330]), .Q(ein[330]) );
  DFF \ereg_reg[331]  ( .D(ereg_next[331]), .CLK(clk), .RST(rst), .I(
        e_init[331]), .Q(ein[331]) );
  DFF \ereg_reg[332]  ( .D(ereg_next[332]), .CLK(clk), .RST(rst), .I(
        e_init[332]), .Q(ein[332]) );
  DFF \ereg_reg[333]  ( .D(ereg_next[333]), .CLK(clk), .RST(rst), .I(
        e_init[333]), .Q(ein[333]) );
  DFF \ereg_reg[334]  ( .D(ereg_next[334]), .CLK(clk), .RST(rst), .I(
        e_init[334]), .Q(ein[334]) );
  DFF \ereg_reg[335]  ( .D(ereg_next[335]), .CLK(clk), .RST(rst), .I(
        e_init[335]), .Q(ein[335]) );
  DFF \ereg_reg[336]  ( .D(ereg_next[336]), .CLK(clk), .RST(rst), .I(
        e_init[336]), .Q(ein[336]) );
  DFF \ereg_reg[337]  ( .D(ereg_next[337]), .CLK(clk), .RST(rst), .I(
        e_init[337]), .Q(ein[337]) );
  DFF \ereg_reg[338]  ( .D(ereg_next[338]), .CLK(clk), .RST(rst), .I(
        e_init[338]), .Q(ein[338]) );
  DFF \ereg_reg[339]  ( .D(ereg_next[339]), .CLK(clk), .RST(rst), .I(
        e_init[339]), .Q(ein[339]) );
  DFF \ereg_reg[340]  ( .D(ereg_next[340]), .CLK(clk), .RST(rst), .I(
        e_init[340]), .Q(ein[340]) );
  DFF \ereg_reg[341]  ( .D(ereg_next[341]), .CLK(clk), .RST(rst), .I(
        e_init[341]), .Q(ein[341]) );
  DFF \ereg_reg[342]  ( .D(ereg_next[342]), .CLK(clk), .RST(rst), .I(
        e_init[342]), .Q(ein[342]) );
  DFF \ereg_reg[343]  ( .D(ereg_next[343]), .CLK(clk), .RST(rst), .I(
        e_init[343]), .Q(ein[343]) );
  DFF \ereg_reg[344]  ( .D(ereg_next[344]), .CLK(clk), .RST(rst), .I(
        e_init[344]), .Q(ein[344]) );
  DFF \ereg_reg[345]  ( .D(ereg_next[345]), .CLK(clk), .RST(rst), .I(
        e_init[345]), .Q(ein[345]) );
  DFF \ereg_reg[346]  ( .D(ereg_next[346]), .CLK(clk), .RST(rst), .I(
        e_init[346]), .Q(ein[346]) );
  DFF \ereg_reg[347]  ( .D(ereg_next[347]), .CLK(clk), .RST(rst), .I(
        e_init[347]), .Q(ein[347]) );
  DFF \ereg_reg[348]  ( .D(ereg_next[348]), .CLK(clk), .RST(rst), .I(
        e_init[348]), .Q(ein[348]) );
  DFF \ereg_reg[349]  ( .D(ereg_next[349]), .CLK(clk), .RST(rst), .I(
        e_init[349]), .Q(ein[349]) );
  DFF \ereg_reg[350]  ( .D(ereg_next[350]), .CLK(clk), .RST(rst), .I(
        e_init[350]), .Q(ein[350]) );
  DFF \ereg_reg[351]  ( .D(ereg_next[351]), .CLK(clk), .RST(rst), .I(
        e_init[351]), .Q(ein[351]) );
  DFF \ereg_reg[352]  ( .D(ereg_next[352]), .CLK(clk), .RST(rst), .I(
        e_init[352]), .Q(ein[352]) );
  DFF \ereg_reg[353]  ( .D(ereg_next[353]), .CLK(clk), .RST(rst), .I(
        e_init[353]), .Q(ein[353]) );
  DFF \ereg_reg[354]  ( .D(ereg_next[354]), .CLK(clk), .RST(rst), .I(
        e_init[354]), .Q(ein[354]) );
  DFF \ereg_reg[355]  ( .D(ereg_next[355]), .CLK(clk), .RST(rst), .I(
        e_init[355]), .Q(ein[355]) );
  DFF \ereg_reg[356]  ( .D(ereg_next[356]), .CLK(clk), .RST(rst), .I(
        e_init[356]), .Q(ein[356]) );
  DFF \ereg_reg[357]  ( .D(ereg_next[357]), .CLK(clk), .RST(rst), .I(
        e_init[357]), .Q(ein[357]) );
  DFF \ereg_reg[358]  ( .D(ereg_next[358]), .CLK(clk), .RST(rst), .I(
        e_init[358]), .Q(ein[358]) );
  DFF \ereg_reg[359]  ( .D(ereg_next[359]), .CLK(clk), .RST(rst), .I(
        e_init[359]), .Q(ein[359]) );
  DFF \ereg_reg[360]  ( .D(ereg_next[360]), .CLK(clk), .RST(rst), .I(
        e_init[360]), .Q(ein[360]) );
  DFF \ereg_reg[361]  ( .D(ereg_next[361]), .CLK(clk), .RST(rst), .I(
        e_init[361]), .Q(ein[361]) );
  DFF \ereg_reg[362]  ( .D(ereg_next[362]), .CLK(clk), .RST(rst), .I(
        e_init[362]), .Q(ein[362]) );
  DFF \ereg_reg[363]  ( .D(ereg_next[363]), .CLK(clk), .RST(rst), .I(
        e_init[363]), .Q(ein[363]) );
  DFF \ereg_reg[364]  ( .D(ereg_next[364]), .CLK(clk), .RST(rst), .I(
        e_init[364]), .Q(ein[364]) );
  DFF \ereg_reg[365]  ( .D(ereg_next[365]), .CLK(clk), .RST(rst), .I(
        e_init[365]), .Q(ein[365]) );
  DFF \ereg_reg[366]  ( .D(ereg_next[366]), .CLK(clk), .RST(rst), .I(
        e_init[366]), .Q(ein[366]) );
  DFF \ereg_reg[367]  ( .D(ereg_next[367]), .CLK(clk), .RST(rst), .I(
        e_init[367]), .Q(ein[367]) );
  DFF \ereg_reg[368]  ( .D(ereg_next[368]), .CLK(clk), .RST(rst), .I(
        e_init[368]), .Q(ein[368]) );
  DFF \ereg_reg[369]  ( .D(ereg_next[369]), .CLK(clk), .RST(rst), .I(
        e_init[369]), .Q(ein[369]) );
  DFF \ereg_reg[370]  ( .D(ereg_next[370]), .CLK(clk), .RST(rst), .I(
        e_init[370]), .Q(ein[370]) );
  DFF \ereg_reg[371]  ( .D(ereg_next[371]), .CLK(clk), .RST(rst), .I(
        e_init[371]), .Q(ein[371]) );
  DFF \ereg_reg[372]  ( .D(ereg_next[372]), .CLK(clk), .RST(rst), .I(
        e_init[372]), .Q(ein[372]) );
  DFF \ereg_reg[373]  ( .D(ereg_next[373]), .CLK(clk), .RST(rst), .I(
        e_init[373]), .Q(ein[373]) );
  DFF \ereg_reg[374]  ( .D(ereg_next[374]), .CLK(clk), .RST(rst), .I(
        e_init[374]), .Q(ein[374]) );
  DFF \ereg_reg[375]  ( .D(ereg_next[375]), .CLK(clk), .RST(rst), .I(
        e_init[375]), .Q(ein[375]) );
  DFF \ereg_reg[376]  ( .D(ereg_next[376]), .CLK(clk), .RST(rst), .I(
        e_init[376]), .Q(ein[376]) );
  DFF \ereg_reg[377]  ( .D(ereg_next[377]), .CLK(clk), .RST(rst), .I(
        e_init[377]), .Q(ein[377]) );
  DFF \ereg_reg[378]  ( .D(ereg_next[378]), .CLK(clk), .RST(rst), .I(
        e_init[378]), .Q(ein[378]) );
  DFF \ereg_reg[379]  ( .D(ereg_next[379]), .CLK(clk), .RST(rst), .I(
        e_init[379]), .Q(ein[379]) );
  DFF \ereg_reg[380]  ( .D(ereg_next[380]), .CLK(clk), .RST(rst), .I(
        e_init[380]), .Q(ein[380]) );
  DFF \ereg_reg[381]  ( .D(ereg_next[381]), .CLK(clk), .RST(rst), .I(
        e_init[381]), .Q(ein[381]) );
  DFF \ereg_reg[382]  ( .D(ereg_next[382]), .CLK(clk), .RST(rst), .I(
        e_init[382]), .Q(ein[382]) );
  DFF \ereg_reg[383]  ( .D(ereg_next[383]), .CLK(clk), .RST(rst), .I(
        e_init[383]), .Q(ein[383]) );
  DFF \ereg_reg[384]  ( .D(ereg_next[384]), .CLK(clk), .RST(rst), .I(
        e_init[384]), .Q(ein[384]) );
  DFF \ereg_reg[385]  ( .D(ereg_next[385]), .CLK(clk), .RST(rst), .I(
        e_init[385]), .Q(ein[385]) );
  DFF \ereg_reg[386]  ( .D(ereg_next[386]), .CLK(clk), .RST(rst), .I(
        e_init[386]), .Q(ein[386]) );
  DFF \ereg_reg[387]  ( .D(ereg_next[387]), .CLK(clk), .RST(rst), .I(
        e_init[387]), .Q(ein[387]) );
  DFF \ereg_reg[388]  ( .D(ereg_next[388]), .CLK(clk), .RST(rst), .I(
        e_init[388]), .Q(ein[388]) );
  DFF \ereg_reg[389]  ( .D(ereg_next[389]), .CLK(clk), .RST(rst), .I(
        e_init[389]), .Q(ein[389]) );
  DFF \ereg_reg[390]  ( .D(ereg_next[390]), .CLK(clk), .RST(rst), .I(
        e_init[390]), .Q(ein[390]) );
  DFF \ereg_reg[391]  ( .D(ereg_next[391]), .CLK(clk), .RST(rst), .I(
        e_init[391]), .Q(ein[391]) );
  DFF \ereg_reg[392]  ( .D(ereg_next[392]), .CLK(clk), .RST(rst), .I(
        e_init[392]), .Q(ein[392]) );
  DFF \ereg_reg[393]  ( .D(ereg_next[393]), .CLK(clk), .RST(rst), .I(
        e_init[393]), .Q(ein[393]) );
  DFF \ereg_reg[394]  ( .D(ereg_next[394]), .CLK(clk), .RST(rst), .I(
        e_init[394]), .Q(ein[394]) );
  DFF \ereg_reg[395]  ( .D(ereg_next[395]), .CLK(clk), .RST(rst), .I(
        e_init[395]), .Q(ein[395]) );
  DFF \ereg_reg[396]  ( .D(ereg_next[396]), .CLK(clk), .RST(rst), .I(
        e_init[396]), .Q(ein[396]) );
  DFF \ereg_reg[397]  ( .D(ereg_next[397]), .CLK(clk), .RST(rst), .I(
        e_init[397]), .Q(ein[397]) );
  DFF \ereg_reg[398]  ( .D(ereg_next[398]), .CLK(clk), .RST(rst), .I(
        e_init[398]), .Q(ein[398]) );
  DFF \ereg_reg[399]  ( .D(ereg_next[399]), .CLK(clk), .RST(rst), .I(
        e_init[399]), .Q(ein[399]) );
  DFF \ereg_reg[400]  ( .D(ereg_next[400]), .CLK(clk), .RST(rst), .I(
        e_init[400]), .Q(ein[400]) );
  DFF \ereg_reg[401]  ( .D(ereg_next[401]), .CLK(clk), .RST(rst), .I(
        e_init[401]), .Q(ein[401]) );
  DFF \ereg_reg[402]  ( .D(ereg_next[402]), .CLK(clk), .RST(rst), .I(
        e_init[402]), .Q(ein[402]) );
  DFF \ereg_reg[403]  ( .D(ereg_next[403]), .CLK(clk), .RST(rst), .I(
        e_init[403]), .Q(ein[403]) );
  DFF \ereg_reg[404]  ( .D(ereg_next[404]), .CLK(clk), .RST(rst), .I(
        e_init[404]), .Q(ein[404]) );
  DFF \ereg_reg[405]  ( .D(ereg_next[405]), .CLK(clk), .RST(rst), .I(
        e_init[405]), .Q(ein[405]) );
  DFF \ereg_reg[406]  ( .D(ereg_next[406]), .CLK(clk), .RST(rst), .I(
        e_init[406]), .Q(ein[406]) );
  DFF \ereg_reg[407]  ( .D(ereg_next[407]), .CLK(clk), .RST(rst), .I(
        e_init[407]), .Q(ein[407]) );
  DFF \ereg_reg[408]  ( .D(ereg_next[408]), .CLK(clk), .RST(rst), .I(
        e_init[408]), .Q(ein[408]) );
  DFF \ereg_reg[409]  ( .D(ereg_next[409]), .CLK(clk), .RST(rst), .I(
        e_init[409]), .Q(ein[409]) );
  DFF \ereg_reg[410]  ( .D(ereg_next[410]), .CLK(clk), .RST(rst), .I(
        e_init[410]), .Q(ein[410]) );
  DFF \ereg_reg[411]  ( .D(ereg_next[411]), .CLK(clk), .RST(rst), .I(
        e_init[411]), .Q(ein[411]) );
  DFF \ereg_reg[412]  ( .D(ereg_next[412]), .CLK(clk), .RST(rst), .I(
        e_init[412]), .Q(ein[412]) );
  DFF \ereg_reg[413]  ( .D(ereg_next[413]), .CLK(clk), .RST(rst), .I(
        e_init[413]), .Q(ein[413]) );
  DFF \ereg_reg[414]  ( .D(ereg_next[414]), .CLK(clk), .RST(rst), .I(
        e_init[414]), .Q(ein[414]) );
  DFF \ereg_reg[415]  ( .D(ereg_next[415]), .CLK(clk), .RST(rst), .I(
        e_init[415]), .Q(ein[415]) );
  DFF \ereg_reg[416]  ( .D(ereg_next[416]), .CLK(clk), .RST(rst), .I(
        e_init[416]), .Q(ein[416]) );
  DFF \ereg_reg[417]  ( .D(ereg_next[417]), .CLK(clk), .RST(rst), .I(
        e_init[417]), .Q(ein[417]) );
  DFF \ereg_reg[418]  ( .D(ereg_next[418]), .CLK(clk), .RST(rst), .I(
        e_init[418]), .Q(ein[418]) );
  DFF \ereg_reg[419]  ( .D(ereg_next[419]), .CLK(clk), .RST(rst), .I(
        e_init[419]), .Q(ein[419]) );
  DFF \ereg_reg[420]  ( .D(ereg_next[420]), .CLK(clk), .RST(rst), .I(
        e_init[420]), .Q(ein[420]) );
  DFF \ereg_reg[421]  ( .D(ereg_next[421]), .CLK(clk), .RST(rst), .I(
        e_init[421]), .Q(ein[421]) );
  DFF \ereg_reg[422]  ( .D(ereg_next[422]), .CLK(clk), .RST(rst), .I(
        e_init[422]), .Q(ein[422]) );
  DFF \ereg_reg[423]  ( .D(ereg_next[423]), .CLK(clk), .RST(rst), .I(
        e_init[423]), .Q(ein[423]) );
  DFF \ereg_reg[424]  ( .D(ereg_next[424]), .CLK(clk), .RST(rst), .I(
        e_init[424]), .Q(ein[424]) );
  DFF \ereg_reg[425]  ( .D(ereg_next[425]), .CLK(clk), .RST(rst), .I(
        e_init[425]), .Q(ein[425]) );
  DFF \ereg_reg[426]  ( .D(ereg_next[426]), .CLK(clk), .RST(rst), .I(
        e_init[426]), .Q(ein[426]) );
  DFF \ereg_reg[427]  ( .D(ereg_next[427]), .CLK(clk), .RST(rst), .I(
        e_init[427]), .Q(ein[427]) );
  DFF \ereg_reg[428]  ( .D(ereg_next[428]), .CLK(clk), .RST(rst), .I(
        e_init[428]), .Q(ein[428]) );
  DFF \ereg_reg[429]  ( .D(ereg_next[429]), .CLK(clk), .RST(rst), .I(
        e_init[429]), .Q(ein[429]) );
  DFF \ereg_reg[430]  ( .D(ereg_next[430]), .CLK(clk), .RST(rst), .I(
        e_init[430]), .Q(ein[430]) );
  DFF \ereg_reg[431]  ( .D(ereg_next[431]), .CLK(clk), .RST(rst), .I(
        e_init[431]), .Q(ein[431]) );
  DFF \ereg_reg[432]  ( .D(ereg_next[432]), .CLK(clk), .RST(rst), .I(
        e_init[432]), .Q(ein[432]) );
  DFF \ereg_reg[433]  ( .D(ereg_next[433]), .CLK(clk), .RST(rst), .I(
        e_init[433]), .Q(ein[433]) );
  DFF \ereg_reg[434]  ( .D(ereg_next[434]), .CLK(clk), .RST(rst), .I(
        e_init[434]), .Q(ein[434]) );
  DFF \ereg_reg[435]  ( .D(ereg_next[435]), .CLK(clk), .RST(rst), .I(
        e_init[435]), .Q(ein[435]) );
  DFF \ereg_reg[436]  ( .D(ereg_next[436]), .CLK(clk), .RST(rst), .I(
        e_init[436]), .Q(ein[436]) );
  DFF \ereg_reg[437]  ( .D(ereg_next[437]), .CLK(clk), .RST(rst), .I(
        e_init[437]), .Q(ein[437]) );
  DFF \ereg_reg[438]  ( .D(ereg_next[438]), .CLK(clk), .RST(rst), .I(
        e_init[438]), .Q(ein[438]) );
  DFF \ereg_reg[439]  ( .D(ereg_next[439]), .CLK(clk), .RST(rst), .I(
        e_init[439]), .Q(ein[439]) );
  DFF \ereg_reg[440]  ( .D(ereg_next[440]), .CLK(clk), .RST(rst), .I(
        e_init[440]), .Q(ein[440]) );
  DFF \ereg_reg[441]  ( .D(ereg_next[441]), .CLK(clk), .RST(rst), .I(
        e_init[441]), .Q(ein[441]) );
  DFF \ereg_reg[442]  ( .D(ereg_next[442]), .CLK(clk), .RST(rst), .I(
        e_init[442]), .Q(ein[442]) );
  DFF \ereg_reg[443]  ( .D(ereg_next[443]), .CLK(clk), .RST(rst), .I(
        e_init[443]), .Q(ein[443]) );
  DFF \ereg_reg[444]  ( .D(ereg_next[444]), .CLK(clk), .RST(rst), .I(
        e_init[444]), .Q(ein[444]) );
  DFF \ereg_reg[445]  ( .D(ereg_next[445]), .CLK(clk), .RST(rst), .I(
        e_init[445]), .Q(ein[445]) );
  DFF \ereg_reg[446]  ( .D(ereg_next[446]), .CLK(clk), .RST(rst), .I(
        e_init[446]), .Q(ein[446]) );
  DFF \ereg_reg[447]  ( .D(ereg_next[447]), .CLK(clk), .RST(rst), .I(
        e_init[447]), .Q(ein[447]) );
  DFF \ereg_reg[448]  ( .D(ereg_next[448]), .CLK(clk), .RST(rst), .I(
        e_init[448]), .Q(ein[448]) );
  DFF \ereg_reg[449]  ( .D(ereg_next[449]), .CLK(clk), .RST(rst), .I(
        e_init[449]), .Q(ein[449]) );
  DFF \ereg_reg[450]  ( .D(ereg_next[450]), .CLK(clk), .RST(rst), .I(
        e_init[450]), .Q(ein[450]) );
  DFF \ereg_reg[451]  ( .D(ereg_next[451]), .CLK(clk), .RST(rst), .I(
        e_init[451]), .Q(ein[451]) );
  DFF \ereg_reg[452]  ( .D(ereg_next[452]), .CLK(clk), .RST(rst), .I(
        e_init[452]), .Q(ein[452]) );
  DFF \ereg_reg[453]  ( .D(ereg_next[453]), .CLK(clk), .RST(rst), .I(
        e_init[453]), .Q(ein[453]) );
  DFF \ereg_reg[454]  ( .D(ereg_next[454]), .CLK(clk), .RST(rst), .I(
        e_init[454]), .Q(ein[454]) );
  DFF \ereg_reg[455]  ( .D(ereg_next[455]), .CLK(clk), .RST(rst), .I(
        e_init[455]), .Q(ein[455]) );
  DFF \ereg_reg[456]  ( .D(ereg_next[456]), .CLK(clk), .RST(rst), .I(
        e_init[456]), .Q(ein[456]) );
  DFF \ereg_reg[457]  ( .D(ereg_next[457]), .CLK(clk), .RST(rst), .I(
        e_init[457]), .Q(ein[457]) );
  DFF \ereg_reg[458]  ( .D(ereg_next[458]), .CLK(clk), .RST(rst), .I(
        e_init[458]), .Q(ein[458]) );
  DFF \ereg_reg[459]  ( .D(ereg_next[459]), .CLK(clk), .RST(rst), .I(
        e_init[459]), .Q(ein[459]) );
  DFF \ereg_reg[460]  ( .D(ereg_next[460]), .CLK(clk), .RST(rst), .I(
        e_init[460]), .Q(ein[460]) );
  DFF \ereg_reg[461]  ( .D(ereg_next[461]), .CLK(clk), .RST(rst), .I(
        e_init[461]), .Q(ein[461]) );
  DFF \ereg_reg[462]  ( .D(ereg_next[462]), .CLK(clk), .RST(rst), .I(
        e_init[462]), .Q(ein[462]) );
  DFF \ereg_reg[463]  ( .D(ereg_next[463]), .CLK(clk), .RST(rst), .I(
        e_init[463]), .Q(ein[463]) );
  DFF \ereg_reg[464]  ( .D(ereg_next[464]), .CLK(clk), .RST(rst), .I(
        e_init[464]), .Q(ein[464]) );
  DFF \ereg_reg[465]  ( .D(ereg_next[465]), .CLK(clk), .RST(rst), .I(
        e_init[465]), .Q(ein[465]) );
  DFF \ereg_reg[466]  ( .D(ereg_next[466]), .CLK(clk), .RST(rst), .I(
        e_init[466]), .Q(ein[466]) );
  DFF \ereg_reg[467]  ( .D(ereg_next[467]), .CLK(clk), .RST(rst), .I(
        e_init[467]), .Q(ein[467]) );
  DFF \ereg_reg[468]  ( .D(ereg_next[468]), .CLK(clk), .RST(rst), .I(
        e_init[468]), .Q(ein[468]) );
  DFF \ereg_reg[469]  ( .D(ereg_next[469]), .CLK(clk), .RST(rst), .I(
        e_init[469]), .Q(ein[469]) );
  DFF \ereg_reg[470]  ( .D(ereg_next[470]), .CLK(clk), .RST(rst), .I(
        e_init[470]), .Q(ein[470]) );
  DFF \ereg_reg[471]  ( .D(ereg_next[471]), .CLK(clk), .RST(rst), .I(
        e_init[471]), .Q(ein[471]) );
  DFF \ereg_reg[472]  ( .D(ereg_next[472]), .CLK(clk), .RST(rst), .I(
        e_init[472]), .Q(ein[472]) );
  DFF \ereg_reg[473]  ( .D(ereg_next[473]), .CLK(clk), .RST(rst), .I(
        e_init[473]), .Q(ein[473]) );
  DFF \ereg_reg[474]  ( .D(ereg_next[474]), .CLK(clk), .RST(rst), .I(
        e_init[474]), .Q(ein[474]) );
  DFF \ereg_reg[475]  ( .D(ereg_next[475]), .CLK(clk), .RST(rst), .I(
        e_init[475]), .Q(ein[475]) );
  DFF \ereg_reg[476]  ( .D(ereg_next[476]), .CLK(clk), .RST(rst), .I(
        e_init[476]), .Q(ein[476]) );
  DFF \ereg_reg[477]  ( .D(ereg_next[477]), .CLK(clk), .RST(rst), .I(
        e_init[477]), .Q(ein[477]) );
  DFF \ereg_reg[478]  ( .D(ereg_next[478]), .CLK(clk), .RST(rst), .I(
        e_init[478]), .Q(ein[478]) );
  DFF \ereg_reg[479]  ( .D(ereg_next[479]), .CLK(clk), .RST(rst), .I(
        e_init[479]), .Q(ein[479]) );
  DFF \ereg_reg[480]  ( .D(ereg_next[480]), .CLK(clk), .RST(rst), .I(
        e_init[480]), .Q(ein[480]) );
  DFF \ereg_reg[481]  ( .D(ereg_next[481]), .CLK(clk), .RST(rst), .I(
        e_init[481]), .Q(ein[481]) );
  DFF \ereg_reg[482]  ( .D(ereg_next[482]), .CLK(clk), .RST(rst), .I(
        e_init[482]), .Q(ein[482]) );
  DFF \ereg_reg[483]  ( .D(ereg_next[483]), .CLK(clk), .RST(rst), .I(
        e_init[483]), .Q(ein[483]) );
  DFF \ereg_reg[484]  ( .D(ereg_next[484]), .CLK(clk), .RST(rst), .I(
        e_init[484]), .Q(ein[484]) );
  DFF \ereg_reg[485]  ( .D(ereg_next[485]), .CLK(clk), .RST(rst), .I(
        e_init[485]), .Q(ein[485]) );
  DFF \ereg_reg[486]  ( .D(ereg_next[486]), .CLK(clk), .RST(rst), .I(
        e_init[486]), .Q(ein[486]) );
  DFF \ereg_reg[487]  ( .D(ereg_next[487]), .CLK(clk), .RST(rst), .I(
        e_init[487]), .Q(ein[487]) );
  DFF \ereg_reg[488]  ( .D(ereg_next[488]), .CLK(clk), .RST(rst), .I(
        e_init[488]), .Q(ein[488]) );
  DFF \ereg_reg[489]  ( .D(ereg_next[489]), .CLK(clk), .RST(rst), .I(
        e_init[489]), .Q(ein[489]) );
  DFF \ereg_reg[490]  ( .D(ereg_next[490]), .CLK(clk), .RST(rst), .I(
        e_init[490]), .Q(ein[490]) );
  DFF \ereg_reg[491]  ( .D(ereg_next[491]), .CLK(clk), .RST(rst), .I(
        e_init[491]), .Q(ein[491]) );
  DFF \ereg_reg[492]  ( .D(ereg_next[492]), .CLK(clk), .RST(rst), .I(
        e_init[492]), .Q(ein[492]) );
  DFF \ereg_reg[493]  ( .D(ereg_next[493]), .CLK(clk), .RST(rst), .I(
        e_init[493]), .Q(ein[493]) );
  DFF \ereg_reg[494]  ( .D(ereg_next[494]), .CLK(clk), .RST(rst), .I(
        e_init[494]), .Q(ein[494]) );
  DFF \ereg_reg[495]  ( .D(ereg_next[495]), .CLK(clk), .RST(rst), .I(
        e_init[495]), .Q(ein[495]) );
  DFF \ereg_reg[496]  ( .D(ereg_next[496]), .CLK(clk), .RST(rst), .I(
        e_init[496]), .Q(ein[496]) );
  DFF \ereg_reg[497]  ( .D(ereg_next[497]), .CLK(clk), .RST(rst), .I(
        e_init[497]), .Q(ein[497]) );
  DFF \ereg_reg[498]  ( .D(ereg_next[498]), .CLK(clk), .RST(rst), .I(
        e_init[498]), .Q(ein[498]) );
  DFF \ereg_reg[499]  ( .D(ereg_next[499]), .CLK(clk), .RST(rst), .I(
        e_init[499]), .Q(ein[499]) );
  DFF \ereg_reg[500]  ( .D(ereg_next[500]), .CLK(clk), .RST(rst), .I(
        e_init[500]), .Q(ein[500]) );
  DFF \ereg_reg[501]  ( .D(ereg_next[501]), .CLK(clk), .RST(rst), .I(
        e_init[501]), .Q(ein[501]) );
  DFF \ereg_reg[502]  ( .D(ereg_next[502]), .CLK(clk), .RST(rst), .I(
        e_init[502]), .Q(ein[502]) );
  DFF \ereg_reg[503]  ( .D(ereg_next[503]), .CLK(clk), .RST(rst), .I(
        e_init[503]), .Q(ein[503]) );
  DFF \ereg_reg[504]  ( .D(ereg_next[504]), .CLK(clk), .RST(rst), .I(
        e_init[504]), .Q(ein[504]) );
  DFF \ereg_reg[505]  ( .D(ereg_next[505]), .CLK(clk), .RST(rst), .I(
        e_init[505]), .Q(ein[505]) );
  DFF \ereg_reg[506]  ( .D(ereg_next[506]), .CLK(clk), .RST(rst), .I(
        e_init[506]), .Q(ein[506]) );
  DFF \ereg_reg[507]  ( .D(ereg_next[507]), .CLK(clk), .RST(rst), .I(
        e_init[507]), .Q(ein[507]) );
  DFF \ereg_reg[508]  ( .D(ereg_next[508]), .CLK(clk), .RST(rst), .I(
        e_init[508]), .Q(ein[508]) );
  DFF \ereg_reg[509]  ( .D(ereg_next[509]), .CLK(clk), .RST(rst), .I(
        e_init[509]), .Q(ein[509]) );
  DFF \ereg_reg[510]  ( .D(ereg_next[510]), .CLK(clk), .RST(rst), .I(
        e_init[510]), .Q(ein[510]) );
  DFF \ereg_reg[511]  ( .D(ereg_next[511]), .CLK(clk), .RST(rst), .I(
        e_init[511]), .Q(ein[511]) );
  DFF \ereg_reg[512]  ( .D(ereg_next[512]), .CLK(clk), .RST(rst), .I(
        e_init[512]), .Q(ein[512]) );
  DFF \ereg_reg[513]  ( .D(ereg_next[513]), .CLK(clk), .RST(rst), .I(
        e_init[513]), .Q(ein[513]) );
  DFF \ereg_reg[514]  ( .D(ereg_next[514]), .CLK(clk), .RST(rst), .I(
        e_init[514]), .Q(ein[514]) );
  DFF \ereg_reg[515]  ( .D(ereg_next[515]), .CLK(clk), .RST(rst), .I(
        e_init[515]), .Q(ein[515]) );
  DFF \ereg_reg[516]  ( .D(ereg_next[516]), .CLK(clk), .RST(rst), .I(
        e_init[516]), .Q(ein[516]) );
  DFF \ereg_reg[517]  ( .D(ereg_next[517]), .CLK(clk), .RST(rst), .I(
        e_init[517]), .Q(ein[517]) );
  DFF \ereg_reg[518]  ( .D(ereg_next[518]), .CLK(clk), .RST(rst), .I(
        e_init[518]), .Q(ein[518]) );
  DFF \ereg_reg[519]  ( .D(ereg_next[519]), .CLK(clk), .RST(rst), .I(
        e_init[519]), .Q(ein[519]) );
  DFF \ereg_reg[520]  ( .D(ereg_next[520]), .CLK(clk), .RST(rst), .I(
        e_init[520]), .Q(ein[520]) );
  DFF \ereg_reg[521]  ( .D(ereg_next[521]), .CLK(clk), .RST(rst), .I(
        e_init[521]), .Q(ein[521]) );
  DFF \ereg_reg[522]  ( .D(ereg_next[522]), .CLK(clk), .RST(rst), .I(
        e_init[522]), .Q(ein[522]) );
  DFF \ereg_reg[523]  ( .D(ereg_next[523]), .CLK(clk), .RST(rst), .I(
        e_init[523]), .Q(ein[523]) );
  DFF \ereg_reg[524]  ( .D(ereg_next[524]), .CLK(clk), .RST(rst), .I(
        e_init[524]), .Q(ein[524]) );
  DFF \ereg_reg[525]  ( .D(ereg_next[525]), .CLK(clk), .RST(rst), .I(
        e_init[525]), .Q(ein[525]) );
  DFF \ereg_reg[526]  ( .D(ereg_next[526]), .CLK(clk), .RST(rst), .I(
        e_init[526]), .Q(ein[526]) );
  DFF \ereg_reg[527]  ( .D(ereg_next[527]), .CLK(clk), .RST(rst), .I(
        e_init[527]), .Q(ein[527]) );
  DFF \ereg_reg[528]  ( .D(ereg_next[528]), .CLK(clk), .RST(rst), .I(
        e_init[528]), .Q(ein[528]) );
  DFF \ereg_reg[529]  ( .D(ereg_next[529]), .CLK(clk), .RST(rst), .I(
        e_init[529]), .Q(ein[529]) );
  DFF \ereg_reg[530]  ( .D(ereg_next[530]), .CLK(clk), .RST(rst), .I(
        e_init[530]), .Q(ein[530]) );
  DFF \ereg_reg[531]  ( .D(ereg_next[531]), .CLK(clk), .RST(rst), .I(
        e_init[531]), .Q(ein[531]) );
  DFF \ereg_reg[532]  ( .D(ereg_next[532]), .CLK(clk), .RST(rst), .I(
        e_init[532]), .Q(ein[532]) );
  DFF \ereg_reg[533]  ( .D(ereg_next[533]), .CLK(clk), .RST(rst), .I(
        e_init[533]), .Q(ein[533]) );
  DFF \ereg_reg[534]  ( .D(ereg_next[534]), .CLK(clk), .RST(rst), .I(
        e_init[534]), .Q(ein[534]) );
  DFF \ereg_reg[535]  ( .D(ereg_next[535]), .CLK(clk), .RST(rst), .I(
        e_init[535]), .Q(ein[535]) );
  DFF \ereg_reg[536]  ( .D(ereg_next[536]), .CLK(clk), .RST(rst), .I(
        e_init[536]), .Q(ein[536]) );
  DFF \ereg_reg[537]  ( .D(ereg_next[537]), .CLK(clk), .RST(rst), .I(
        e_init[537]), .Q(ein[537]) );
  DFF \ereg_reg[538]  ( .D(ereg_next[538]), .CLK(clk), .RST(rst), .I(
        e_init[538]), .Q(ein[538]) );
  DFF \ereg_reg[539]  ( .D(ereg_next[539]), .CLK(clk), .RST(rst), .I(
        e_init[539]), .Q(ein[539]) );
  DFF \ereg_reg[540]  ( .D(ereg_next[540]), .CLK(clk), .RST(rst), .I(
        e_init[540]), .Q(ein[540]) );
  DFF \ereg_reg[541]  ( .D(ereg_next[541]), .CLK(clk), .RST(rst), .I(
        e_init[541]), .Q(ein[541]) );
  DFF \ereg_reg[542]  ( .D(ereg_next[542]), .CLK(clk), .RST(rst), .I(
        e_init[542]), .Q(ein[542]) );
  DFF \ereg_reg[543]  ( .D(ereg_next[543]), .CLK(clk), .RST(rst), .I(
        e_init[543]), .Q(ein[543]) );
  DFF \ereg_reg[544]  ( .D(ereg_next[544]), .CLK(clk), .RST(rst), .I(
        e_init[544]), .Q(ein[544]) );
  DFF \ereg_reg[545]  ( .D(ereg_next[545]), .CLK(clk), .RST(rst), .I(
        e_init[545]), .Q(ein[545]) );
  DFF \ereg_reg[546]  ( .D(ereg_next[546]), .CLK(clk), .RST(rst), .I(
        e_init[546]), .Q(ein[546]) );
  DFF \ereg_reg[547]  ( .D(ereg_next[547]), .CLK(clk), .RST(rst), .I(
        e_init[547]), .Q(ein[547]) );
  DFF \ereg_reg[548]  ( .D(ereg_next[548]), .CLK(clk), .RST(rst), .I(
        e_init[548]), .Q(ein[548]) );
  DFF \ereg_reg[549]  ( .D(ereg_next[549]), .CLK(clk), .RST(rst), .I(
        e_init[549]), .Q(ein[549]) );
  DFF \ereg_reg[550]  ( .D(ereg_next[550]), .CLK(clk), .RST(rst), .I(
        e_init[550]), .Q(ein[550]) );
  DFF \ereg_reg[551]  ( .D(ereg_next[551]), .CLK(clk), .RST(rst), .I(
        e_init[551]), .Q(ein[551]) );
  DFF \ereg_reg[552]  ( .D(ereg_next[552]), .CLK(clk), .RST(rst), .I(
        e_init[552]), .Q(ein[552]) );
  DFF \ereg_reg[553]  ( .D(ereg_next[553]), .CLK(clk), .RST(rst), .I(
        e_init[553]), .Q(ein[553]) );
  DFF \ereg_reg[554]  ( .D(ereg_next[554]), .CLK(clk), .RST(rst), .I(
        e_init[554]), .Q(ein[554]) );
  DFF \ereg_reg[555]  ( .D(ereg_next[555]), .CLK(clk), .RST(rst), .I(
        e_init[555]), .Q(ein[555]) );
  DFF \ereg_reg[556]  ( .D(ereg_next[556]), .CLK(clk), .RST(rst), .I(
        e_init[556]), .Q(ein[556]) );
  DFF \ereg_reg[557]  ( .D(ereg_next[557]), .CLK(clk), .RST(rst), .I(
        e_init[557]), .Q(ein[557]) );
  DFF \ereg_reg[558]  ( .D(ereg_next[558]), .CLK(clk), .RST(rst), .I(
        e_init[558]), .Q(ein[558]) );
  DFF \ereg_reg[559]  ( .D(ereg_next[559]), .CLK(clk), .RST(rst), .I(
        e_init[559]), .Q(ein[559]) );
  DFF \ereg_reg[560]  ( .D(ereg_next[560]), .CLK(clk), .RST(rst), .I(
        e_init[560]), .Q(ein[560]) );
  DFF \ereg_reg[561]  ( .D(ereg_next[561]), .CLK(clk), .RST(rst), .I(
        e_init[561]), .Q(ein[561]) );
  DFF \ereg_reg[562]  ( .D(ereg_next[562]), .CLK(clk), .RST(rst), .I(
        e_init[562]), .Q(ein[562]) );
  DFF \ereg_reg[563]  ( .D(ereg_next[563]), .CLK(clk), .RST(rst), .I(
        e_init[563]), .Q(ein[563]) );
  DFF \ereg_reg[564]  ( .D(ereg_next[564]), .CLK(clk), .RST(rst), .I(
        e_init[564]), .Q(ein[564]) );
  DFF \ereg_reg[565]  ( .D(ereg_next[565]), .CLK(clk), .RST(rst), .I(
        e_init[565]), .Q(ein[565]) );
  DFF \ereg_reg[566]  ( .D(ereg_next[566]), .CLK(clk), .RST(rst), .I(
        e_init[566]), .Q(ein[566]) );
  DFF \ereg_reg[567]  ( .D(ereg_next[567]), .CLK(clk), .RST(rst), .I(
        e_init[567]), .Q(ein[567]) );
  DFF \ereg_reg[568]  ( .D(ereg_next[568]), .CLK(clk), .RST(rst), .I(
        e_init[568]), .Q(ein[568]) );
  DFF \ereg_reg[569]  ( .D(ereg_next[569]), .CLK(clk), .RST(rst), .I(
        e_init[569]), .Q(ein[569]) );
  DFF \ereg_reg[570]  ( .D(ereg_next[570]), .CLK(clk), .RST(rst), .I(
        e_init[570]), .Q(ein[570]) );
  DFF \ereg_reg[571]  ( .D(ereg_next[571]), .CLK(clk), .RST(rst), .I(
        e_init[571]), .Q(ein[571]) );
  DFF \ereg_reg[572]  ( .D(ereg_next[572]), .CLK(clk), .RST(rst), .I(
        e_init[572]), .Q(ein[572]) );
  DFF \ereg_reg[573]  ( .D(ereg_next[573]), .CLK(clk), .RST(rst), .I(
        e_init[573]), .Q(ein[573]) );
  DFF \ereg_reg[574]  ( .D(ereg_next[574]), .CLK(clk), .RST(rst), .I(
        e_init[574]), .Q(ein[574]) );
  DFF \ereg_reg[575]  ( .D(ereg_next[575]), .CLK(clk), .RST(rst), .I(
        e_init[575]), .Q(ein[575]) );
  DFF \ereg_reg[576]  ( .D(ereg_next[576]), .CLK(clk), .RST(rst), .I(
        e_init[576]), .Q(ein[576]) );
  DFF \ereg_reg[577]  ( .D(ereg_next[577]), .CLK(clk), .RST(rst), .I(
        e_init[577]), .Q(ein[577]) );
  DFF \ereg_reg[578]  ( .D(ereg_next[578]), .CLK(clk), .RST(rst), .I(
        e_init[578]), .Q(ein[578]) );
  DFF \ereg_reg[579]  ( .D(ereg_next[579]), .CLK(clk), .RST(rst), .I(
        e_init[579]), .Q(ein[579]) );
  DFF \ereg_reg[580]  ( .D(ereg_next[580]), .CLK(clk), .RST(rst), .I(
        e_init[580]), .Q(ein[580]) );
  DFF \ereg_reg[581]  ( .D(ereg_next[581]), .CLK(clk), .RST(rst), .I(
        e_init[581]), .Q(ein[581]) );
  DFF \ereg_reg[582]  ( .D(ereg_next[582]), .CLK(clk), .RST(rst), .I(
        e_init[582]), .Q(ein[582]) );
  DFF \ereg_reg[583]  ( .D(ereg_next[583]), .CLK(clk), .RST(rst), .I(
        e_init[583]), .Q(ein[583]) );
  DFF \ereg_reg[584]  ( .D(ereg_next[584]), .CLK(clk), .RST(rst), .I(
        e_init[584]), .Q(ein[584]) );
  DFF \ereg_reg[585]  ( .D(ereg_next[585]), .CLK(clk), .RST(rst), .I(
        e_init[585]), .Q(ein[585]) );
  DFF \ereg_reg[586]  ( .D(ereg_next[586]), .CLK(clk), .RST(rst), .I(
        e_init[586]), .Q(ein[586]) );
  DFF \ereg_reg[587]  ( .D(ereg_next[587]), .CLK(clk), .RST(rst), .I(
        e_init[587]), .Q(ein[587]) );
  DFF \ereg_reg[588]  ( .D(ereg_next[588]), .CLK(clk), .RST(rst), .I(
        e_init[588]), .Q(ein[588]) );
  DFF \ereg_reg[589]  ( .D(ereg_next[589]), .CLK(clk), .RST(rst), .I(
        e_init[589]), .Q(ein[589]) );
  DFF \ereg_reg[590]  ( .D(ereg_next[590]), .CLK(clk), .RST(rst), .I(
        e_init[590]), .Q(ein[590]) );
  DFF \ereg_reg[591]  ( .D(ereg_next[591]), .CLK(clk), .RST(rst), .I(
        e_init[591]), .Q(ein[591]) );
  DFF \ereg_reg[592]  ( .D(ereg_next[592]), .CLK(clk), .RST(rst), .I(
        e_init[592]), .Q(ein[592]) );
  DFF \ereg_reg[593]  ( .D(ereg_next[593]), .CLK(clk), .RST(rst), .I(
        e_init[593]), .Q(ein[593]) );
  DFF \ereg_reg[594]  ( .D(ereg_next[594]), .CLK(clk), .RST(rst), .I(
        e_init[594]), .Q(ein[594]) );
  DFF \ereg_reg[595]  ( .D(ereg_next[595]), .CLK(clk), .RST(rst), .I(
        e_init[595]), .Q(ein[595]) );
  DFF \ereg_reg[596]  ( .D(ereg_next[596]), .CLK(clk), .RST(rst), .I(
        e_init[596]), .Q(ein[596]) );
  DFF \ereg_reg[597]  ( .D(ereg_next[597]), .CLK(clk), .RST(rst), .I(
        e_init[597]), .Q(ein[597]) );
  DFF \ereg_reg[598]  ( .D(ereg_next[598]), .CLK(clk), .RST(rst), .I(
        e_init[598]), .Q(ein[598]) );
  DFF \ereg_reg[599]  ( .D(ereg_next[599]), .CLK(clk), .RST(rst), .I(
        e_init[599]), .Q(ein[599]) );
  DFF \ereg_reg[600]  ( .D(ereg_next[600]), .CLK(clk), .RST(rst), .I(
        e_init[600]), .Q(ein[600]) );
  DFF \ereg_reg[601]  ( .D(ereg_next[601]), .CLK(clk), .RST(rst), .I(
        e_init[601]), .Q(ein[601]) );
  DFF \ereg_reg[602]  ( .D(ereg_next[602]), .CLK(clk), .RST(rst), .I(
        e_init[602]), .Q(ein[602]) );
  DFF \ereg_reg[603]  ( .D(ereg_next[603]), .CLK(clk), .RST(rst), .I(
        e_init[603]), .Q(ein[603]) );
  DFF \ereg_reg[604]  ( .D(ereg_next[604]), .CLK(clk), .RST(rst), .I(
        e_init[604]), .Q(ein[604]) );
  DFF \ereg_reg[605]  ( .D(ereg_next[605]), .CLK(clk), .RST(rst), .I(
        e_init[605]), .Q(ein[605]) );
  DFF \ereg_reg[606]  ( .D(ereg_next[606]), .CLK(clk), .RST(rst), .I(
        e_init[606]), .Q(ein[606]) );
  DFF \ereg_reg[607]  ( .D(ereg_next[607]), .CLK(clk), .RST(rst), .I(
        e_init[607]), .Q(ein[607]) );
  DFF \ereg_reg[608]  ( .D(ereg_next[608]), .CLK(clk), .RST(rst), .I(
        e_init[608]), .Q(ein[608]) );
  DFF \ereg_reg[609]  ( .D(ereg_next[609]), .CLK(clk), .RST(rst), .I(
        e_init[609]), .Q(ein[609]) );
  DFF \ereg_reg[610]  ( .D(ereg_next[610]), .CLK(clk), .RST(rst), .I(
        e_init[610]), .Q(ein[610]) );
  DFF \ereg_reg[611]  ( .D(ereg_next[611]), .CLK(clk), .RST(rst), .I(
        e_init[611]), .Q(ein[611]) );
  DFF \ereg_reg[612]  ( .D(ereg_next[612]), .CLK(clk), .RST(rst), .I(
        e_init[612]), .Q(ein[612]) );
  DFF \ereg_reg[613]  ( .D(ereg_next[613]), .CLK(clk), .RST(rst), .I(
        e_init[613]), .Q(ein[613]) );
  DFF \ereg_reg[614]  ( .D(ereg_next[614]), .CLK(clk), .RST(rst), .I(
        e_init[614]), .Q(ein[614]) );
  DFF \ereg_reg[615]  ( .D(ereg_next[615]), .CLK(clk), .RST(rst), .I(
        e_init[615]), .Q(ein[615]) );
  DFF \ereg_reg[616]  ( .D(ereg_next[616]), .CLK(clk), .RST(rst), .I(
        e_init[616]), .Q(ein[616]) );
  DFF \ereg_reg[617]  ( .D(ereg_next[617]), .CLK(clk), .RST(rst), .I(
        e_init[617]), .Q(ein[617]) );
  DFF \ereg_reg[618]  ( .D(ereg_next[618]), .CLK(clk), .RST(rst), .I(
        e_init[618]), .Q(ein[618]) );
  DFF \ereg_reg[619]  ( .D(ereg_next[619]), .CLK(clk), .RST(rst), .I(
        e_init[619]), .Q(ein[619]) );
  DFF \ereg_reg[620]  ( .D(ereg_next[620]), .CLK(clk), .RST(rst), .I(
        e_init[620]), .Q(ein[620]) );
  DFF \ereg_reg[621]  ( .D(ereg_next[621]), .CLK(clk), .RST(rst), .I(
        e_init[621]), .Q(ein[621]) );
  DFF \ereg_reg[622]  ( .D(ereg_next[622]), .CLK(clk), .RST(rst), .I(
        e_init[622]), .Q(ein[622]) );
  DFF \ereg_reg[623]  ( .D(ereg_next[623]), .CLK(clk), .RST(rst), .I(
        e_init[623]), .Q(ein[623]) );
  DFF \ereg_reg[624]  ( .D(ereg_next[624]), .CLK(clk), .RST(rst), .I(
        e_init[624]), .Q(ein[624]) );
  DFF \ereg_reg[625]  ( .D(ereg_next[625]), .CLK(clk), .RST(rst), .I(
        e_init[625]), .Q(ein[625]) );
  DFF \ereg_reg[626]  ( .D(ereg_next[626]), .CLK(clk), .RST(rst), .I(
        e_init[626]), .Q(ein[626]) );
  DFF \ereg_reg[627]  ( .D(ereg_next[627]), .CLK(clk), .RST(rst), .I(
        e_init[627]), .Q(ein[627]) );
  DFF \ereg_reg[628]  ( .D(ereg_next[628]), .CLK(clk), .RST(rst), .I(
        e_init[628]), .Q(ein[628]) );
  DFF \ereg_reg[629]  ( .D(ereg_next[629]), .CLK(clk), .RST(rst), .I(
        e_init[629]), .Q(ein[629]) );
  DFF \ereg_reg[630]  ( .D(ereg_next[630]), .CLK(clk), .RST(rst), .I(
        e_init[630]), .Q(ein[630]) );
  DFF \ereg_reg[631]  ( .D(ereg_next[631]), .CLK(clk), .RST(rst), .I(
        e_init[631]), .Q(ein[631]) );
  DFF \ereg_reg[632]  ( .D(ereg_next[632]), .CLK(clk), .RST(rst), .I(
        e_init[632]), .Q(ein[632]) );
  DFF \ereg_reg[633]  ( .D(ereg_next[633]), .CLK(clk), .RST(rst), .I(
        e_init[633]), .Q(ein[633]) );
  DFF \ereg_reg[634]  ( .D(ereg_next[634]), .CLK(clk), .RST(rst), .I(
        e_init[634]), .Q(ein[634]) );
  DFF \ereg_reg[635]  ( .D(ereg_next[635]), .CLK(clk), .RST(rst), .I(
        e_init[635]), .Q(ein[635]) );
  DFF \ereg_reg[636]  ( .D(ereg_next[636]), .CLK(clk), .RST(rst), .I(
        e_init[636]), .Q(ein[636]) );
  DFF \ereg_reg[637]  ( .D(ereg_next[637]), .CLK(clk), .RST(rst), .I(
        e_init[637]), .Q(ein[637]) );
  DFF \ereg_reg[638]  ( .D(ereg_next[638]), .CLK(clk), .RST(rst), .I(
        e_init[638]), .Q(ein[638]) );
  DFF \ereg_reg[639]  ( .D(ereg_next[639]), .CLK(clk), .RST(rst), .I(
        e_init[639]), .Q(ein[639]) );
  DFF \ereg_reg[640]  ( .D(ereg_next[640]), .CLK(clk), .RST(rst), .I(
        e_init[640]), .Q(ein[640]) );
  DFF \ereg_reg[641]  ( .D(ereg_next[641]), .CLK(clk), .RST(rst), .I(
        e_init[641]), .Q(ein[641]) );
  DFF \ereg_reg[642]  ( .D(ereg_next[642]), .CLK(clk), .RST(rst), .I(
        e_init[642]), .Q(ein[642]) );
  DFF \ereg_reg[643]  ( .D(ereg_next[643]), .CLK(clk), .RST(rst), .I(
        e_init[643]), .Q(ein[643]) );
  DFF \ereg_reg[644]  ( .D(ereg_next[644]), .CLK(clk), .RST(rst), .I(
        e_init[644]), .Q(ein[644]) );
  DFF \ereg_reg[645]  ( .D(ereg_next[645]), .CLK(clk), .RST(rst), .I(
        e_init[645]), .Q(ein[645]) );
  DFF \ereg_reg[646]  ( .D(ereg_next[646]), .CLK(clk), .RST(rst), .I(
        e_init[646]), .Q(ein[646]) );
  DFF \ereg_reg[647]  ( .D(ereg_next[647]), .CLK(clk), .RST(rst), .I(
        e_init[647]), .Q(ein[647]) );
  DFF \ereg_reg[648]  ( .D(ereg_next[648]), .CLK(clk), .RST(rst), .I(
        e_init[648]), .Q(ein[648]) );
  DFF \ereg_reg[649]  ( .D(ereg_next[649]), .CLK(clk), .RST(rst), .I(
        e_init[649]), .Q(ein[649]) );
  DFF \ereg_reg[650]  ( .D(ereg_next[650]), .CLK(clk), .RST(rst), .I(
        e_init[650]), .Q(ein[650]) );
  DFF \ereg_reg[651]  ( .D(ereg_next[651]), .CLK(clk), .RST(rst), .I(
        e_init[651]), .Q(ein[651]) );
  DFF \ereg_reg[652]  ( .D(ereg_next[652]), .CLK(clk), .RST(rst), .I(
        e_init[652]), .Q(ein[652]) );
  DFF \ereg_reg[653]  ( .D(ereg_next[653]), .CLK(clk), .RST(rst), .I(
        e_init[653]), .Q(ein[653]) );
  DFF \ereg_reg[654]  ( .D(ereg_next[654]), .CLK(clk), .RST(rst), .I(
        e_init[654]), .Q(ein[654]) );
  DFF \ereg_reg[655]  ( .D(ereg_next[655]), .CLK(clk), .RST(rst), .I(
        e_init[655]), .Q(ein[655]) );
  DFF \ereg_reg[656]  ( .D(ereg_next[656]), .CLK(clk), .RST(rst), .I(
        e_init[656]), .Q(ein[656]) );
  DFF \ereg_reg[657]  ( .D(ereg_next[657]), .CLK(clk), .RST(rst), .I(
        e_init[657]), .Q(ein[657]) );
  DFF \ereg_reg[658]  ( .D(ereg_next[658]), .CLK(clk), .RST(rst), .I(
        e_init[658]), .Q(ein[658]) );
  DFF \ereg_reg[659]  ( .D(ereg_next[659]), .CLK(clk), .RST(rst), .I(
        e_init[659]), .Q(ein[659]) );
  DFF \ereg_reg[660]  ( .D(ereg_next[660]), .CLK(clk), .RST(rst), .I(
        e_init[660]), .Q(ein[660]) );
  DFF \ereg_reg[661]  ( .D(ereg_next[661]), .CLK(clk), .RST(rst), .I(
        e_init[661]), .Q(ein[661]) );
  DFF \ereg_reg[662]  ( .D(ereg_next[662]), .CLK(clk), .RST(rst), .I(
        e_init[662]), .Q(ein[662]) );
  DFF \ereg_reg[663]  ( .D(ereg_next[663]), .CLK(clk), .RST(rst), .I(
        e_init[663]), .Q(ein[663]) );
  DFF \ereg_reg[664]  ( .D(ereg_next[664]), .CLK(clk), .RST(rst), .I(
        e_init[664]), .Q(ein[664]) );
  DFF \ereg_reg[665]  ( .D(ereg_next[665]), .CLK(clk), .RST(rst), .I(
        e_init[665]), .Q(ein[665]) );
  DFF \ereg_reg[666]  ( .D(ereg_next[666]), .CLK(clk), .RST(rst), .I(
        e_init[666]), .Q(ein[666]) );
  DFF \ereg_reg[667]  ( .D(ereg_next[667]), .CLK(clk), .RST(rst), .I(
        e_init[667]), .Q(ein[667]) );
  DFF \ereg_reg[668]  ( .D(ereg_next[668]), .CLK(clk), .RST(rst), .I(
        e_init[668]), .Q(ein[668]) );
  DFF \ereg_reg[669]  ( .D(ereg_next[669]), .CLK(clk), .RST(rst), .I(
        e_init[669]), .Q(ein[669]) );
  DFF \ereg_reg[670]  ( .D(ereg_next[670]), .CLK(clk), .RST(rst), .I(
        e_init[670]), .Q(ein[670]) );
  DFF \ereg_reg[671]  ( .D(ereg_next[671]), .CLK(clk), .RST(rst), .I(
        e_init[671]), .Q(ein[671]) );
  DFF \ereg_reg[672]  ( .D(ereg_next[672]), .CLK(clk), .RST(rst), .I(
        e_init[672]), .Q(ein[672]) );
  DFF \ereg_reg[673]  ( .D(ereg_next[673]), .CLK(clk), .RST(rst), .I(
        e_init[673]), .Q(ein[673]) );
  DFF \ereg_reg[674]  ( .D(ereg_next[674]), .CLK(clk), .RST(rst), .I(
        e_init[674]), .Q(ein[674]) );
  DFF \ereg_reg[675]  ( .D(ereg_next[675]), .CLK(clk), .RST(rst), .I(
        e_init[675]), .Q(ein[675]) );
  DFF \ereg_reg[676]  ( .D(ereg_next[676]), .CLK(clk), .RST(rst), .I(
        e_init[676]), .Q(ein[676]) );
  DFF \ereg_reg[677]  ( .D(ereg_next[677]), .CLK(clk), .RST(rst), .I(
        e_init[677]), .Q(ein[677]) );
  DFF \ereg_reg[678]  ( .D(ereg_next[678]), .CLK(clk), .RST(rst), .I(
        e_init[678]), .Q(ein[678]) );
  DFF \ereg_reg[679]  ( .D(ereg_next[679]), .CLK(clk), .RST(rst), .I(
        e_init[679]), .Q(ein[679]) );
  DFF \ereg_reg[680]  ( .D(ereg_next[680]), .CLK(clk), .RST(rst), .I(
        e_init[680]), .Q(ein[680]) );
  DFF \ereg_reg[681]  ( .D(ereg_next[681]), .CLK(clk), .RST(rst), .I(
        e_init[681]), .Q(ein[681]) );
  DFF \ereg_reg[682]  ( .D(ereg_next[682]), .CLK(clk), .RST(rst), .I(
        e_init[682]), .Q(ein[682]) );
  DFF \ereg_reg[683]  ( .D(ereg_next[683]), .CLK(clk), .RST(rst), .I(
        e_init[683]), .Q(ein[683]) );
  DFF \ereg_reg[684]  ( .D(ereg_next[684]), .CLK(clk), .RST(rst), .I(
        e_init[684]), .Q(ein[684]) );
  DFF \ereg_reg[685]  ( .D(ereg_next[685]), .CLK(clk), .RST(rst), .I(
        e_init[685]), .Q(ein[685]) );
  DFF \ereg_reg[686]  ( .D(ereg_next[686]), .CLK(clk), .RST(rst), .I(
        e_init[686]), .Q(ein[686]) );
  DFF \ereg_reg[687]  ( .D(ereg_next[687]), .CLK(clk), .RST(rst), .I(
        e_init[687]), .Q(ein[687]) );
  DFF \ereg_reg[688]  ( .D(ereg_next[688]), .CLK(clk), .RST(rst), .I(
        e_init[688]), .Q(ein[688]) );
  DFF \ereg_reg[689]  ( .D(ereg_next[689]), .CLK(clk), .RST(rst), .I(
        e_init[689]), .Q(ein[689]) );
  DFF \ereg_reg[690]  ( .D(ereg_next[690]), .CLK(clk), .RST(rst), .I(
        e_init[690]), .Q(ein[690]) );
  DFF \ereg_reg[691]  ( .D(ereg_next[691]), .CLK(clk), .RST(rst), .I(
        e_init[691]), .Q(ein[691]) );
  DFF \ereg_reg[692]  ( .D(ereg_next[692]), .CLK(clk), .RST(rst), .I(
        e_init[692]), .Q(ein[692]) );
  DFF \ereg_reg[693]  ( .D(ereg_next[693]), .CLK(clk), .RST(rst), .I(
        e_init[693]), .Q(ein[693]) );
  DFF \ereg_reg[694]  ( .D(ereg_next[694]), .CLK(clk), .RST(rst), .I(
        e_init[694]), .Q(ein[694]) );
  DFF \ereg_reg[695]  ( .D(ereg_next[695]), .CLK(clk), .RST(rst), .I(
        e_init[695]), .Q(ein[695]) );
  DFF \ereg_reg[696]  ( .D(ereg_next[696]), .CLK(clk), .RST(rst), .I(
        e_init[696]), .Q(ein[696]) );
  DFF \ereg_reg[697]  ( .D(ereg_next[697]), .CLK(clk), .RST(rst), .I(
        e_init[697]), .Q(ein[697]) );
  DFF \ereg_reg[698]  ( .D(ereg_next[698]), .CLK(clk), .RST(rst), .I(
        e_init[698]), .Q(ein[698]) );
  DFF \ereg_reg[699]  ( .D(ereg_next[699]), .CLK(clk), .RST(rst), .I(
        e_init[699]), .Q(ein[699]) );
  DFF \ereg_reg[700]  ( .D(ereg_next[700]), .CLK(clk), .RST(rst), .I(
        e_init[700]), .Q(ein[700]) );
  DFF \ereg_reg[701]  ( .D(ereg_next[701]), .CLK(clk), .RST(rst), .I(
        e_init[701]), .Q(ein[701]) );
  DFF \ereg_reg[702]  ( .D(ereg_next[702]), .CLK(clk), .RST(rst), .I(
        e_init[702]), .Q(ein[702]) );
  DFF \ereg_reg[703]  ( .D(ereg_next[703]), .CLK(clk), .RST(rst), .I(
        e_init[703]), .Q(ein[703]) );
  DFF \ereg_reg[704]  ( .D(ereg_next[704]), .CLK(clk), .RST(rst), .I(
        e_init[704]), .Q(ein[704]) );
  DFF \ereg_reg[705]  ( .D(ereg_next[705]), .CLK(clk), .RST(rst), .I(
        e_init[705]), .Q(ein[705]) );
  DFF \ereg_reg[706]  ( .D(ereg_next[706]), .CLK(clk), .RST(rst), .I(
        e_init[706]), .Q(ein[706]) );
  DFF \ereg_reg[707]  ( .D(ereg_next[707]), .CLK(clk), .RST(rst), .I(
        e_init[707]), .Q(ein[707]) );
  DFF \ereg_reg[708]  ( .D(ereg_next[708]), .CLK(clk), .RST(rst), .I(
        e_init[708]), .Q(ein[708]) );
  DFF \ereg_reg[709]  ( .D(ereg_next[709]), .CLK(clk), .RST(rst), .I(
        e_init[709]), .Q(ein[709]) );
  DFF \ereg_reg[710]  ( .D(ereg_next[710]), .CLK(clk), .RST(rst), .I(
        e_init[710]), .Q(ein[710]) );
  DFF \ereg_reg[711]  ( .D(ereg_next[711]), .CLK(clk), .RST(rst), .I(
        e_init[711]), .Q(ein[711]) );
  DFF \ereg_reg[712]  ( .D(ereg_next[712]), .CLK(clk), .RST(rst), .I(
        e_init[712]), .Q(ein[712]) );
  DFF \ereg_reg[713]  ( .D(ereg_next[713]), .CLK(clk), .RST(rst), .I(
        e_init[713]), .Q(ein[713]) );
  DFF \ereg_reg[714]  ( .D(ereg_next[714]), .CLK(clk), .RST(rst), .I(
        e_init[714]), .Q(ein[714]) );
  DFF \ereg_reg[715]  ( .D(ereg_next[715]), .CLK(clk), .RST(rst), .I(
        e_init[715]), .Q(ein[715]) );
  DFF \ereg_reg[716]  ( .D(ereg_next[716]), .CLK(clk), .RST(rst), .I(
        e_init[716]), .Q(ein[716]) );
  DFF \ereg_reg[717]  ( .D(ereg_next[717]), .CLK(clk), .RST(rst), .I(
        e_init[717]), .Q(ein[717]) );
  DFF \ereg_reg[718]  ( .D(ereg_next[718]), .CLK(clk), .RST(rst), .I(
        e_init[718]), .Q(ein[718]) );
  DFF \ereg_reg[719]  ( .D(ereg_next[719]), .CLK(clk), .RST(rst), .I(
        e_init[719]), .Q(ein[719]) );
  DFF \ereg_reg[720]  ( .D(ereg_next[720]), .CLK(clk), .RST(rst), .I(
        e_init[720]), .Q(ein[720]) );
  DFF \ereg_reg[721]  ( .D(ereg_next[721]), .CLK(clk), .RST(rst), .I(
        e_init[721]), .Q(ein[721]) );
  DFF \ereg_reg[722]  ( .D(ereg_next[722]), .CLK(clk), .RST(rst), .I(
        e_init[722]), .Q(ein[722]) );
  DFF \ereg_reg[723]  ( .D(ereg_next[723]), .CLK(clk), .RST(rst), .I(
        e_init[723]), .Q(ein[723]) );
  DFF \ereg_reg[724]  ( .D(ereg_next[724]), .CLK(clk), .RST(rst), .I(
        e_init[724]), .Q(ein[724]) );
  DFF \ereg_reg[725]  ( .D(ereg_next[725]), .CLK(clk), .RST(rst), .I(
        e_init[725]), .Q(ein[725]) );
  DFF \ereg_reg[726]  ( .D(ereg_next[726]), .CLK(clk), .RST(rst), .I(
        e_init[726]), .Q(ein[726]) );
  DFF \ereg_reg[727]  ( .D(ereg_next[727]), .CLK(clk), .RST(rst), .I(
        e_init[727]), .Q(ein[727]) );
  DFF \ereg_reg[728]  ( .D(ereg_next[728]), .CLK(clk), .RST(rst), .I(
        e_init[728]), .Q(ein[728]) );
  DFF \ereg_reg[729]  ( .D(ereg_next[729]), .CLK(clk), .RST(rst), .I(
        e_init[729]), .Q(ein[729]) );
  DFF \ereg_reg[730]  ( .D(ereg_next[730]), .CLK(clk), .RST(rst), .I(
        e_init[730]), .Q(ein[730]) );
  DFF \ereg_reg[731]  ( .D(ereg_next[731]), .CLK(clk), .RST(rst), .I(
        e_init[731]), .Q(ein[731]) );
  DFF \ereg_reg[732]  ( .D(ereg_next[732]), .CLK(clk), .RST(rst), .I(
        e_init[732]), .Q(ein[732]) );
  DFF \ereg_reg[733]  ( .D(ereg_next[733]), .CLK(clk), .RST(rst), .I(
        e_init[733]), .Q(ein[733]) );
  DFF \ereg_reg[734]  ( .D(ereg_next[734]), .CLK(clk), .RST(rst), .I(
        e_init[734]), .Q(ein[734]) );
  DFF \ereg_reg[735]  ( .D(ereg_next[735]), .CLK(clk), .RST(rst), .I(
        e_init[735]), .Q(ein[735]) );
  DFF \ereg_reg[736]  ( .D(ereg_next[736]), .CLK(clk), .RST(rst), .I(
        e_init[736]), .Q(ein[736]) );
  DFF \ereg_reg[737]  ( .D(ereg_next[737]), .CLK(clk), .RST(rst), .I(
        e_init[737]), .Q(ein[737]) );
  DFF \ereg_reg[738]  ( .D(ereg_next[738]), .CLK(clk), .RST(rst), .I(
        e_init[738]), .Q(ein[738]) );
  DFF \ereg_reg[739]  ( .D(ereg_next[739]), .CLK(clk), .RST(rst), .I(
        e_init[739]), .Q(ein[739]) );
  DFF \ereg_reg[740]  ( .D(ereg_next[740]), .CLK(clk), .RST(rst), .I(
        e_init[740]), .Q(ein[740]) );
  DFF \ereg_reg[741]  ( .D(ereg_next[741]), .CLK(clk), .RST(rst), .I(
        e_init[741]), .Q(ein[741]) );
  DFF \ereg_reg[742]  ( .D(ereg_next[742]), .CLK(clk), .RST(rst), .I(
        e_init[742]), .Q(ein[742]) );
  DFF \ereg_reg[743]  ( .D(ereg_next[743]), .CLK(clk), .RST(rst), .I(
        e_init[743]), .Q(ein[743]) );
  DFF \ereg_reg[744]  ( .D(ereg_next[744]), .CLK(clk), .RST(rst), .I(
        e_init[744]), .Q(ein[744]) );
  DFF \ereg_reg[745]  ( .D(ereg_next[745]), .CLK(clk), .RST(rst), .I(
        e_init[745]), .Q(ein[745]) );
  DFF \ereg_reg[746]  ( .D(ereg_next[746]), .CLK(clk), .RST(rst), .I(
        e_init[746]), .Q(ein[746]) );
  DFF \ereg_reg[747]  ( .D(ereg_next[747]), .CLK(clk), .RST(rst), .I(
        e_init[747]), .Q(ein[747]) );
  DFF \ereg_reg[748]  ( .D(ereg_next[748]), .CLK(clk), .RST(rst), .I(
        e_init[748]), .Q(ein[748]) );
  DFF \ereg_reg[749]  ( .D(ereg_next[749]), .CLK(clk), .RST(rst), .I(
        e_init[749]), .Q(ein[749]) );
  DFF \ereg_reg[750]  ( .D(ereg_next[750]), .CLK(clk), .RST(rst), .I(
        e_init[750]), .Q(ein[750]) );
  DFF \ereg_reg[751]  ( .D(ereg_next[751]), .CLK(clk), .RST(rst), .I(
        e_init[751]), .Q(ein[751]) );
  DFF \ereg_reg[752]  ( .D(ereg_next[752]), .CLK(clk), .RST(rst), .I(
        e_init[752]), .Q(ein[752]) );
  DFF \ereg_reg[753]  ( .D(ereg_next[753]), .CLK(clk), .RST(rst), .I(
        e_init[753]), .Q(ein[753]) );
  DFF \ereg_reg[754]  ( .D(ereg_next[754]), .CLK(clk), .RST(rst), .I(
        e_init[754]), .Q(ein[754]) );
  DFF \ereg_reg[755]  ( .D(ereg_next[755]), .CLK(clk), .RST(rst), .I(
        e_init[755]), .Q(ein[755]) );
  DFF \ereg_reg[756]  ( .D(ereg_next[756]), .CLK(clk), .RST(rst), .I(
        e_init[756]), .Q(ein[756]) );
  DFF \ereg_reg[757]  ( .D(ereg_next[757]), .CLK(clk), .RST(rst), .I(
        e_init[757]), .Q(ein[757]) );
  DFF \ereg_reg[758]  ( .D(ereg_next[758]), .CLK(clk), .RST(rst), .I(
        e_init[758]), .Q(ein[758]) );
  DFF \ereg_reg[759]  ( .D(ereg_next[759]), .CLK(clk), .RST(rst), .I(
        e_init[759]), .Q(ein[759]) );
  DFF \ereg_reg[760]  ( .D(ereg_next[760]), .CLK(clk), .RST(rst), .I(
        e_init[760]), .Q(ein[760]) );
  DFF \ereg_reg[761]  ( .D(ereg_next[761]), .CLK(clk), .RST(rst), .I(
        e_init[761]), .Q(ein[761]) );
  DFF \ereg_reg[762]  ( .D(ereg_next[762]), .CLK(clk), .RST(rst), .I(
        e_init[762]), .Q(ein[762]) );
  DFF \ereg_reg[763]  ( .D(ereg_next[763]), .CLK(clk), .RST(rst), .I(
        e_init[763]), .Q(ein[763]) );
  DFF \ereg_reg[764]  ( .D(ereg_next[764]), .CLK(clk), .RST(rst), .I(
        e_init[764]), .Q(ein[764]) );
  DFF \ereg_reg[765]  ( .D(ereg_next[765]), .CLK(clk), .RST(rst), .I(
        e_init[765]), .Q(ein[765]) );
  DFF \ereg_reg[766]  ( .D(ereg_next[766]), .CLK(clk), .RST(rst), .I(
        e_init[766]), .Q(ein[766]) );
  DFF \ereg_reg[767]  ( .D(ereg_next[767]), .CLK(clk), .RST(rst), .I(
        e_init[767]), .Q(ein[767]) );
  DFF \ereg_reg[768]  ( .D(ereg_next[768]), .CLK(clk), .RST(rst), .I(
        e_init[768]), .Q(ein[768]) );
  DFF \ereg_reg[769]  ( .D(ereg_next[769]), .CLK(clk), .RST(rst), .I(
        e_init[769]), .Q(ein[769]) );
  DFF \ereg_reg[770]  ( .D(ereg_next[770]), .CLK(clk), .RST(rst), .I(
        e_init[770]), .Q(ein[770]) );
  DFF \ereg_reg[771]  ( .D(ereg_next[771]), .CLK(clk), .RST(rst), .I(
        e_init[771]), .Q(ein[771]) );
  DFF \ereg_reg[772]  ( .D(ereg_next[772]), .CLK(clk), .RST(rst), .I(
        e_init[772]), .Q(ein[772]) );
  DFF \ereg_reg[773]  ( .D(ereg_next[773]), .CLK(clk), .RST(rst), .I(
        e_init[773]), .Q(ein[773]) );
  DFF \ereg_reg[774]  ( .D(ereg_next[774]), .CLK(clk), .RST(rst), .I(
        e_init[774]), .Q(ein[774]) );
  DFF \ereg_reg[775]  ( .D(ereg_next[775]), .CLK(clk), .RST(rst), .I(
        e_init[775]), .Q(ein[775]) );
  DFF \ereg_reg[776]  ( .D(ereg_next[776]), .CLK(clk), .RST(rst), .I(
        e_init[776]), .Q(ein[776]) );
  DFF \ereg_reg[777]  ( .D(ereg_next[777]), .CLK(clk), .RST(rst), .I(
        e_init[777]), .Q(ein[777]) );
  DFF \ereg_reg[778]  ( .D(ereg_next[778]), .CLK(clk), .RST(rst), .I(
        e_init[778]), .Q(ein[778]) );
  DFF \ereg_reg[779]  ( .D(ereg_next[779]), .CLK(clk), .RST(rst), .I(
        e_init[779]), .Q(ein[779]) );
  DFF \ereg_reg[780]  ( .D(ereg_next[780]), .CLK(clk), .RST(rst), .I(
        e_init[780]), .Q(ein[780]) );
  DFF \ereg_reg[781]  ( .D(ereg_next[781]), .CLK(clk), .RST(rst), .I(
        e_init[781]), .Q(ein[781]) );
  DFF \ereg_reg[782]  ( .D(ereg_next[782]), .CLK(clk), .RST(rst), .I(
        e_init[782]), .Q(ein[782]) );
  DFF \ereg_reg[783]  ( .D(ereg_next[783]), .CLK(clk), .RST(rst), .I(
        e_init[783]), .Q(ein[783]) );
  DFF \ereg_reg[784]  ( .D(ereg_next[784]), .CLK(clk), .RST(rst), .I(
        e_init[784]), .Q(ein[784]) );
  DFF \ereg_reg[785]  ( .D(ereg_next[785]), .CLK(clk), .RST(rst), .I(
        e_init[785]), .Q(ein[785]) );
  DFF \ereg_reg[786]  ( .D(ereg_next[786]), .CLK(clk), .RST(rst), .I(
        e_init[786]), .Q(ein[786]) );
  DFF \ereg_reg[787]  ( .D(ereg_next[787]), .CLK(clk), .RST(rst), .I(
        e_init[787]), .Q(ein[787]) );
  DFF \ereg_reg[788]  ( .D(ereg_next[788]), .CLK(clk), .RST(rst), .I(
        e_init[788]), .Q(ein[788]) );
  DFF \ereg_reg[789]  ( .D(ereg_next[789]), .CLK(clk), .RST(rst), .I(
        e_init[789]), .Q(ein[789]) );
  DFF \ereg_reg[790]  ( .D(ereg_next[790]), .CLK(clk), .RST(rst), .I(
        e_init[790]), .Q(ein[790]) );
  DFF \ereg_reg[791]  ( .D(ereg_next[791]), .CLK(clk), .RST(rst), .I(
        e_init[791]), .Q(ein[791]) );
  DFF \ereg_reg[792]  ( .D(ereg_next[792]), .CLK(clk), .RST(rst), .I(
        e_init[792]), .Q(ein[792]) );
  DFF \ereg_reg[793]  ( .D(ereg_next[793]), .CLK(clk), .RST(rst), .I(
        e_init[793]), .Q(ein[793]) );
  DFF \ereg_reg[794]  ( .D(ereg_next[794]), .CLK(clk), .RST(rst), .I(
        e_init[794]), .Q(ein[794]) );
  DFF \ereg_reg[795]  ( .D(ereg_next[795]), .CLK(clk), .RST(rst), .I(
        e_init[795]), .Q(ein[795]) );
  DFF \ereg_reg[796]  ( .D(ereg_next[796]), .CLK(clk), .RST(rst), .I(
        e_init[796]), .Q(ein[796]) );
  DFF \ereg_reg[797]  ( .D(ereg_next[797]), .CLK(clk), .RST(rst), .I(
        e_init[797]), .Q(ein[797]) );
  DFF \ereg_reg[798]  ( .D(ereg_next[798]), .CLK(clk), .RST(rst), .I(
        e_init[798]), .Q(ein[798]) );
  DFF \ereg_reg[799]  ( .D(ereg_next[799]), .CLK(clk), .RST(rst), .I(
        e_init[799]), .Q(ein[799]) );
  DFF \ereg_reg[800]  ( .D(ereg_next[800]), .CLK(clk), .RST(rst), .I(
        e_init[800]), .Q(ein[800]) );
  DFF \ereg_reg[801]  ( .D(ereg_next[801]), .CLK(clk), .RST(rst), .I(
        e_init[801]), .Q(ein[801]) );
  DFF \ereg_reg[802]  ( .D(ereg_next[802]), .CLK(clk), .RST(rst), .I(
        e_init[802]), .Q(ein[802]) );
  DFF \ereg_reg[803]  ( .D(ereg_next[803]), .CLK(clk), .RST(rst), .I(
        e_init[803]), .Q(ein[803]) );
  DFF \ereg_reg[804]  ( .D(ereg_next[804]), .CLK(clk), .RST(rst), .I(
        e_init[804]), .Q(ein[804]) );
  DFF \ereg_reg[805]  ( .D(ereg_next[805]), .CLK(clk), .RST(rst), .I(
        e_init[805]), .Q(ein[805]) );
  DFF \ereg_reg[806]  ( .D(ereg_next[806]), .CLK(clk), .RST(rst), .I(
        e_init[806]), .Q(ein[806]) );
  DFF \ereg_reg[807]  ( .D(ereg_next[807]), .CLK(clk), .RST(rst), .I(
        e_init[807]), .Q(ein[807]) );
  DFF \ereg_reg[808]  ( .D(ereg_next[808]), .CLK(clk), .RST(rst), .I(
        e_init[808]), .Q(ein[808]) );
  DFF \ereg_reg[809]  ( .D(ereg_next[809]), .CLK(clk), .RST(rst), .I(
        e_init[809]), .Q(ein[809]) );
  DFF \ereg_reg[810]  ( .D(ereg_next[810]), .CLK(clk), .RST(rst), .I(
        e_init[810]), .Q(ein[810]) );
  DFF \ereg_reg[811]  ( .D(ereg_next[811]), .CLK(clk), .RST(rst), .I(
        e_init[811]), .Q(ein[811]) );
  DFF \ereg_reg[812]  ( .D(ereg_next[812]), .CLK(clk), .RST(rst), .I(
        e_init[812]), .Q(ein[812]) );
  DFF \ereg_reg[813]  ( .D(ereg_next[813]), .CLK(clk), .RST(rst), .I(
        e_init[813]), .Q(ein[813]) );
  DFF \ereg_reg[814]  ( .D(ereg_next[814]), .CLK(clk), .RST(rst), .I(
        e_init[814]), .Q(ein[814]) );
  DFF \ereg_reg[815]  ( .D(ereg_next[815]), .CLK(clk), .RST(rst), .I(
        e_init[815]), .Q(ein[815]) );
  DFF \ereg_reg[816]  ( .D(ereg_next[816]), .CLK(clk), .RST(rst), .I(
        e_init[816]), .Q(ein[816]) );
  DFF \ereg_reg[817]  ( .D(ereg_next[817]), .CLK(clk), .RST(rst), .I(
        e_init[817]), .Q(ein[817]) );
  DFF \ereg_reg[818]  ( .D(ereg_next[818]), .CLK(clk), .RST(rst), .I(
        e_init[818]), .Q(ein[818]) );
  DFF \ereg_reg[819]  ( .D(ereg_next[819]), .CLK(clk), .RST(rst), .I(
        e_init[819]), .Q(ein[819]) );
  DFF \ereg_reg[820]  ( .D(ereg_next[820]), .CLK(clk), .RST(rst), .I(
        e_init[820]), .Q(ein[820]) );
  DFF \ereg_reg[821]  ( .D(ereg_next[821]), .CLK(clk), .RST(rst), .I(
        e_init[821]), .Q(ein[821]) );
  DFF \ereg_reg[822]  ( .D(ereg_next[822]), .CLK(clk), .RST(rst), .I(
        e_init[822]), .Q(ein[822]) );
  DFF \ereg_reg[823]  ( .D(ereg_next[823]), .CLK(clk), .RST(rst), .I(
        e_init[823]), .Q(ein[823]) );
  DFF \ereg_reg[824]  ( .D(ereg_next[824]), .CLK(clk), .RST(rst), .I(
        e_init[824]), .Q(ein[824]) );
  DFF \ereg_reg[825]  ( .D(ereg_next[825]), .CLK(clk), .RST(rst), .I(
        e_init[825]), .Q(ein[825]) );
  DFF \ereg_reg[826]  ( .D(ereg_next[826]), .CLK(clk), .RST(rst), .I(
        e_init[826]), .Q(ein[826]) );
  DFF \ereg_reg[827]  ( .D(ereg_next[827]), .CLK(clk), .RST(rst), .I(
        e_init[827]), .Q(ein[827]) );
  DFF \ereg_reg[828]  ( .D(ereg_next[828]), .CLK(clk), .RST(rst), .I(
        e_init[828]), .Q(ein[828]) );
  DFF \ereg_reg[829]  ( .D(ereg_next[829]), .CLK(clk), .RST(rst), .I(
        e_init[829]), .Q(ein[829]) );
  DFF \ereg_reg[830]  ( .D(ereg_next[830]), .CLK(clk), .RST(rst), .I(
        e_init[830]), .Q(ein[830]) );
  DFF \ereg_reg[831]  ( .D(ereg_next[831]), .CLK(clk), .RST(rst), .I(
        e_init[831]), .Q(ein[831]) );
  DFF \ereg_reg[832]  ( .D(ereg_next[832]), .CLK(clk), .RST(rst), .I(
        e_init[832]), .Q(ein[832]) );
  DFF \ereg_reg[833]  ( .D(ereg_next[833]), .CLK(clk), .RST(rst), .I(
        e_init[833]), .Q(ein[833]) );
  DFF \ereg_reg[834]  ( .D(ereg_next[834]), .CLK(clk), .RST(rst), .I(
        e_init[834]), .Q(ein[834]) );
  DFF \ereg_reg[835]  ( .D(ereg_next[835]), .CLK(clk), .RST(rst), .I(
        e_init[835]), .Q(ein[835]) );
  DFF \ereg_reg[836]  ( .D(ereg_next[836]), .CLK(clk), .RST(rst), .I(
        e_init[836]), .Q(ein[836]) );
  DFF \ereg_reg[837]  ( .D(ereg_next[837]), .CLK(clk), .RST(rst), .I(
        e_init[837]), .Q(ein[837]) );
  DFF \ereg_reg[838]  ( .D(ereg_next[838]), .CLK(clk), .RST(rst), .I(
        e_init[838]), .Q(ein[838]) );
  DFF \ereg_reg[839]  ( .D(ereg_next[839]), .CLK(clk), .RST(rst), .I(
        e_init[839]), .Q(ein[839]) );
  DFF \ereg_reg[840]  ( .D(ereg_next[840]), .CLK(clk), .RST(rst), .I(
        e_init[840]), .Q(ein[840]) );
  DFF \ereg_reg[841]  ( .D(ereg_next[841]), .CLK(clk), .RST(rst), .I(
        e_init[841]), .Q(ein[841]) );
  DFF \ereg_reg[842]  ( .D(ereg_next[842]), .CLK(clk), .RST(rst), .I(
        e_init[842]), .Q(ein[842]) );
  DFF \ereg_reg[843]  ( .D(ereg_next[843]), .CLK(clk), .RST(rst), .I(
        e_init[843]), .Q(ein[843]) );
  DFF \ereg_reg[844]  ( .D(ereg_next[844]), .CLK(clk), .RST(rst), .I(
        e_init[844]), .Q(ein[844]) );
  DFF \ereg_reg[845]  ( .D(ereg_next[845]), .CLK(clk), .RST(rst), .I(
        e_init[845]), .Q(ein[845]) );
  DFF \ereg_reg[846]  ( .D(ereg_next[846]), .CLK(clk), .RST(rst), .I(
        e_init[846]), .Q(ein[846]) );
  DFF \ereg_reg[847]  ( .D(ereg_next[847]), .CLK(clk), .RST(rst), .I(
        e_init[847]), .Q(ein[847]) );
  DFF \ereg_reg[848]  ( .D(ereg_next[848]), .CLK(clk), .RST(rst), .I(
        e_init[848]), .Q(ein[848]) );
  DFF \ereg_reg[849]  ( .D(ereg_next[849]), .CLK(clk), .RST(rst), .I(
        e_init[849]), .Q(ein[849]) );
  DFF \ereg_reg[850]  ( .D(ereg_next[850]), .CLK(clk), .RST(rst), .I(
        e_init[850]), .Q(ein[850]) );
  DFF \ereg_reg[851]  ( .D(ereg_next[851]), .CLK(clk), .RST(rst), .I(
        e_init[851]), .Q(ein[851]) );
  DFF \ereg_reg[852]  ( .D(ereg_next[852]), .CLK(clk), .RST(rst), .I(
        e_init[852]), .Q(ein[852]) );
  DFF \ereg_reg[853]  ( .D(ereg_next[853]), .CLK(clk), .RST(rst), .I(
        e_init[853]), .Q(ein[853]) );
  DFF \ereg_reg[854]  ( .D(ereg_next[854]), .CLK(clk), .RST(rst), .I(
        e_init[854]), .Q(ein[854]) );
  DFF \ereg_reg[855]  ( .D(ereg_next[855]), .CLK(clk), .RST(rst), .I(
        e_init[855]), .Q(ein[855]) );
  DFF \ereg_reg[856]  ( .D(ereg_next[856]), .CLK(clk), .RST(rst), .I(
        e_init[856]), .Q(ein[856]) );
  DFF \ereg_reg[857]  ( .D(ereg_next[857]), .CLK(clk), .RST(rst), .I(
        e_init[857]), .Q(ein[857]) );
  DFF \ereg_reg[858]  ( .D(ereg_next[858]), .CLK(clk), .RST(rst), .I(
        e_init[858]), .Q(ein[858]) );
  DFF \ereg_reg[859]  ( .D(ereg_next[859]), .CLK(clk), .RST(rst), .I(
        e_init[859]), .Q(ein[859]) );
  DFF \ereg_reg[860]  ( .D(ereg_next[860]), .CLK(clk), .RST(rst), .I(
        e_init[860]), .Q(ein[860]) );
  DFF \ereg_reg[861]  ( .D(ereg_next[861]), .CLK(clk), .RST(rst), .I(
        e_init[861]), .Q(ein[861]) );
  DFF \ereg_reg[862]  ( .D(ereg_next[862]), .CLK(clk), .RST(rst), .I(
        e_init[862]), .Q(ein[862]) );
  DFF \ereg_reg[863]  ( .D(ereg_next[863]), .CLK(clk), .RST(rst), .I(
        e_init[863]), .Q(ein[863]) );
  DFF \ereg_reg[864]  ( .D(ereg_next[864]), .CLK(clk), .RST(rst), .I(
        e_init[864]), .Q(ein[864]) );
  DFF \ereg_reg[865]  ( .D(ereg_next[865]), .CLK(clk), .RST(rst), .I(
        e_init[865]), .Q(ein[865]) );
  DFF \ereg_reg[866]  ( .D(ereg_next[866]), .CLK(clk), .RST(rst), .I(
        e_init[866]), .Q(ein[866]) );
  DFF \ereg_reg[867]  ( .D(ereg_next[867]), .CLK(clk), .RST(rst), .I(
        e_init[867]), .Q(ein[867]) );
  DFF \ereg_reg[868]  ( .D(ereg_next[868]), .CLK(clk), .RST(rst), .I(
        e_init[868]), .Q(ein[868]) );
  DFF \ereg_reg[869]  ( .D(ereg_next[869]), .CLK(clk), .RST(rst), .I(
        e_init[869]), .Q(ein[869]) );
  DFF \ereg_reg[870]  ( .D(ereg_next[870]), .CLK(clk), .RST(rst), .I(
        e_init[870]), .Q(ein[870]) );
  DFF \ereg_reg[871]  ( .D(ereg_next[871]), .CLK(clk), .RST(rst), .I(
        e_init[871]), .Q(ein[871]) );
  DFF \ereg_reg[872]  ( .D(ereg_next[872]), .CLK(clk), .RST(rst), .I(
        e_init[872]), .Q(ein[872]) );
  DFF \ereg_reg[873]  ( .D(ereg_next[873]), .CLK(clk), .RST(rst), .I(
        e_init[873]), .Q(ein[873]) );
  DFF \ereg_reg[874]  ( .D(ereg_next[874]), .CLK(clk), .RST(rst), .I(
        e_init[874]), .Q(ein[874]) );
  DFF \ereg_reg[875]  ( .D(ereg_next[875]), .CLK(clk), .RST(rst), .I(
        e_init[875]), .Q(ein[875]) );
  DFF \ereg_reg[876]  ( .D(ereg_next[876]), .CLK(clk), .RST(rst), .I(
        e_init[876]), .Q(ein[876]) );
  DFF \ereg_reg[877]  ( .D(ereg_next[877]), .CLK(clk), .RST(rst), .I(
        e_init[877]), .Q(ein[877]) );
  DFF \ereg_reg[878]  ( .D(ereg_next[878]), .CLK(clk), .RST(rst), .I(
        e_init[878]), .Q(ein[878]) );
  DFF \ereg_reg[879]  ( .D(ereg_next[879]), .CLK(clk), .RST(rst), .I(
        e_init[879]), .Q(ein[879]) );
  DFF \ereg_reg[880]  ( .D(ereg_next[880]), .CLK(clk), .RST(rst), .I(
        e_init[880]), .Q(ein[880]) );
  DFF \ereg_reg[881]  ( .D(ereg_next[881]), .CLK(clk), .RST(rst), .I(
        e_init[881]), .Q(ein[881]) );
  DFF \ereg_reg[882]  ( .D(ereg_next[882]), .CLK(clk), .RST(rst), .I(
        e_init[882]), .Q(ein[882]) );
  DFF \ereg_reg[883]  ( .D(ereg_next[883]), .CLK(clk), .RST(rst), .I(
        e_init[883]), .Q(ein[883]) );
  DFF \ereg_reg[884]  ( .D(ereg_next[884]), .CLK(clk), .RST(rst), .I(
        e_init[884]), .Q(ein[884]) );
  DFF \ereg_reg[885]  ( .D(ereg_next[885]), .CLK(clk), .RST(rst), .I(
        e_init[885]), .Q(ein[885]) );
  DFF \ereg_reg[886]  ( .D(ereg_next[886]), .CLK(clk), .RST(rst), .I(
        e_init[886]), .Q(ein[886]) );
  DFF \ereg_reg[887]  ( .D(ereg_next[887]), .CLK(clk), .RST(rst), .I(
        e_init[887]), .Q(ein[887]) );
  DFF \ereg_reg[888]  ( .D(ereg_next[888]), .CLK(clk), .RST(rst), .I(
        e_init[888]), .Q(ein[888]) );
  DFF \ereg_reg[889]  ( .D(ereg_next[889]), .CLK(clk), .RST(rst), .I(
        e_init[889]), .Q(ein[889]) );
  DFF \ereg_reg[890]  ( .D(ereg_next[890]), .CLK(clk), .RST(rst), .I(
        e_init[890]), .Q(ein[890]) );
  DFF \ereg_reg[891]  ( .D(ereg_next[891]), .CLK(clk), .RST(rst), .I(
        e_init[891]), .Q(ein[891]) );
  DFF \ereg_reg[892]  ( .D(ereg_next[892]), .CLK(clk), .RST(rst), .I(
        e_init[892]), .Q(ein[892]) );
  DFF \ereg_reg[893]  ( .D(ereg_next[893]), .CLK(clk), .RST(rst), .I(
        e_init[893]), .Q(ein[893]) );
  DFF \ereg_reg[894]  ( .D(ereg_next[894]), .CLK(clk), .RST(rst), .I(
        e_init[894]), .Q(ein[894]) );
  DFF \ereg_reg[895]  ( .D(ereg_next[895]), .CLK(clk), .RST(rst), .I(
        e_init[895]), .Q(ein[895]) );
  DFF \ereg_reg[896]  ( .D(ereg_next[896]), .CLK(clk), .RST(rst), .I(
        e_init[896]), .Q(ein[896]) );
  DFF \ereg_reg[897]  ( .D(ereg_next[897]), .CLK(clk), .RST(rst), .I(
        e_init[897]), .Q(ein[897]) );
  DFF \ereg_reg[898]  ( .D(ereg_next[898]), .CLK(clk), .RST(rst), .I(
        e_init[898]), .Q(ein[898]) );
  DFF \ereg_reg[899]  ( .D(ereg_next[899]), .CLK(clk), .RST(rst), .I(
        e_init[899]), .Q(ein[899]) );
  DFF \ereg_reg[900]  ( .D(ereg_next[900]), .CLK(clk), .RST(rst), .I(
        e_init[900]), .Q(ein[900]) );
  DFF \ereg_reg[901]  ( .D(ereg_next[901]), .CLK(clk), .RST(rst), .I(
        e_init[901]), .Q(ein[901]) );
  DFF \ereg_reg[902]  ( .D(ereg_next[902]), .CLK(clk), .RST(rst), .I(
        e_init[902]), .Q(ein[902]) );
  DFF \ereg_reg[903]  ( .D(ereg_next[903]), .CLK(clk), .RST(rst), .I(
        e_init[903]), .Q(ein[903]) );
  DFF \ereg_reg[904]  ( .D(ereg_next[904]), .CLK(clk), .RST(rst), .I(
        e_init[904]), .Q(ein[904]) );
  DFF \ereg_reg[905]  ( .D(ereg_next[905]), .CLK(clk), .RST(rst), .I(
        e_init[905]), .Q(ein[905]) );
  DFF \ereg_reg[906]  ( .D(ereg_next[906]), .CLK(clk), .RST(rst), .I(
        e_init[906]), .Q(ein[906]) );
  DFF \ereg_reg[907]  ( .D(ereg_next[907]), .CLK(clk), .RST(rst), .I(
        e_init[907]), .Q(ein[907]) );
  DFF \ereg_reg[908]  ( .D(ereg_next[908]), .CLK(clk), .RST(rst), .I(
        e_init[908]), .Q(ein[908]) );
  DFF \ereg_reg[909]  ( .D(ereg_next[909]), .CLK(clk), .RST(rst), .I(
        e_init[909]), .Q(ein[909]) );
  DFF \ereg_reg[910]  ( .D(ereg_next[910]), .CLK(clk), .RST(rst), .I(
        e_init[910]), .Q(ein[910]) );
  DFF \ereg_reg[911]  ( .D(ereg_next[911]), .CLK(clk), .RST(rst), .I(
        e_init[911]), .Q(ein[911]) );
  DFF \ereg_reg[912]  ( .D(ereg_next[912]), .CLK(clk), .RST(rst), .I(
        e_init[912]), .Q(ein[912]) );
  DFF \ereg_reg[913]  ( .D(ereg_next[913]), .CLK(clk), .RST(rst), .I(
        e_init[913]), .Q(ein[913]) );
  DFF \ereg_reg[914]  ( .D(ereg_next[914]), .CLK(clk), .RST(rst), .I(
        e_init[914]), .Q(ein[914]) );
  DFF \ereg_reg[915]  ( .D(ereg_next[915]), .CLK(clk), .RST(rst), .I(
        e_init[915]), .Q(ein[915]) );
  DFF \ereg_reg[916]  ( .D(ereg_next[916]), .CLK(clk), .RST(rst), .I(
        e_init[916]), .Q(ein[916]) );
  DFF \ereg_reg[917]  ( .D(ereg_next[917]), .CLK(clk), .RST(rst), .I(
        e_init[917]), .Q(ein[917]) );
  DFF \ereg_reg[918]  ( .D(ereg_next[918]), .CLK(clk), .RST(rst), .I(
        e_init[918]), .Q(ein[918]) );
  DFF \ereg_reg[919]  ( .D(ereg_next[919]), .CLK(clk), .RST(rst), .I(
        e_init[919]), .Q(ein[919]) );
  DFF \ereg_reg[920]  ( .D(ereg_next[920]), .CLK(clk), .RST(rst), .I(
        e_init[920]), .Q(ein[920]) );
  DFF \ereg_reg[921]  ( .D(ereg_next[921]), .CLK(clk), .RST(rst), .I(
        e_init[921]), .Q(ein[921]) );
  DFF \ereg_reg[922]  ( .D(ereg_next[922]), .CLK(clk), .RST(rst), .I(
        e_init[922]), .Q(ein[922]) );
  DFF \ereg_reg[923]  ( .D(ereg_next[923]), .CLK(clk), .RST(rst), .I(
        e_init[923]), .Q(ein[923]) );
  DFF \ereg_reg[924]  ( .D(ereg_next[924]), .CLK(clk), .RST(rst), .I(
        e_init[924]), .Q(ein[924]) );
  DFF \ereg_reg[925]  ( .D(ereg_next[925]), .CLK(clk), .RST(rst), .I(
        e_init[925]), .Q(ein[925]) );
  DFF \ereg_reg[926]  ( .D(ereg_next[926]), .CLK(clk), .RST(rst), .I(
        e_init[926]), .Q(ein[926]) );
  DFF \ereg_reg[927]  ( .D(ereg_next[927]), .CLK(clk), .RST(rst), .I(
        e_init[927]), .Q(ein[927]) );
  DFF \ereg_reg[928]  ( .D(ereg_next[928]), .CLK(clk), .RST(rst), .I(
        e_init[928]), .Q(ein[928]) );
  DFF \ereg_reg[929]  ( .D(ereg_next[929]), .CLK(clk), .RST(rst), .I(
        e_init[929]), .Q(ein[929]) );
  DFF \ereg_reg[930]  ( .D(ereg_next[930]), .CLK(clk), .RST(rst), .I(
        e_init[930]), .Q(ein[930]) );
  DFF \ereg_reg[931]  ( .D(ereg_next[931]), .CLK(clk), .RST(rst), .I(
        e_init[931]), .Q(ein[931]) );
  DFF \ereg_reg[932]  ( .D(ereg_next[932]), .CLK(clk), .RST(rst), .I(
        e_init[932]), .Q(ein[932]) );
  DFF \ereg_reg[933]  ( .D(ereg_next[933]), .CLK(clk), .RST(rst), .I(
        e_init[933]), .Q(ein[933]) );
  DFF \ereg_reg[934]  ( .D(ereg_next[934]), .CLK(clk), .RST(rst), .I(
        e_init[934]), .Q(ein[934]) );
  DFF \ereg_reg[935]  ( .D(ereg_next[935]), .CLK(clk), .RST(rst), .I(
        e_init[935]), .Q(ein[935]) );
  DFF \ereg_reg[936]  ( .D(ereg_next[936]), .CLK(clk), .RST(rst), .I(
        e_init[936]), .Q(ein[936]) );
  DFF \ereg_reg[937]  ( .D(ereg_next[937]), .CLK(clk), .RST(rst), .I(
        e_init[937]), .Q(ein[937]) );
  DFF \ereg_reg[938]  ( .D(ereg_next[938]), .CLK(clk), .RST(rst), .I(
        e_init[938]), .Q(ein[938]) );
  DFF \ereg_reg[939]  ( .D(ereg_next[939]), .CLK(clk), .RST(rst), .I(
        e_init[939]), .Q(ein[939]) );
  DFF \ereg_reg[940]  ( .D(ereg_next[940]), .CLK(clk), .RST(rst), .I(
        e_init[940]), .Q(ein[940]) );
  DFF \ereg_reg[941]  ( .D(ereg_next[941]), .CLK(clk), .RST(rst), .I(
        e_init[941]), .Q(ein[941]) );
  DFF \ereg_reg[942]  ( .D(ereg_next[942]), .CLK(clk), .RST(rst), .I(
        e_init[942]), .Q(ein[942]) );
  DFF \ereg_reg[943]  ( .D(ereg_next[943]), .CLK(clk), .RST(rst), .I(
        e_init[943]), .Q(ein[943]) );
  DFF \ereg_reg[944]  ( .D(ereg_next[944]), .CLK(clk), .RST(rst), .I(
        e_init[944]), .Q(ein[944]) );
  DFF \ereg_reg[945]  ( .D(ereg_next[945]), .CLK(clk), .RST(rst), .I(
        e_init[945]), .Q(ein[945]) );
  DFF \ereg_reg[946]  ( .D(ereg_next[946]), .CLK(clk), .RST(rst), .I(
        e_init[946]), .Q(ein[946]) );
  DFF \ereg_reg[947]  ( .D(ereg_next[947]), .CLK(clk), .RST(rst), .I(
        e_init[947]), .Q(ein[947]) );
  DFF \ereg_reg[948]  ( .D(ereg_next[948]), .CLK(clk), .RST(rst), .I(
        e_init[948]), .Q(ein[948]) );
  DFF \ereg_reg[949]  ( .D(ereg_next[949]), .CLK(clk), .RST(rst), .I(
        e_init[949]), .Q(ein[949]) );
  DFF \ereg_reg[950]  ( .D(ereg_next[950]), .CLK(clk), .RST(rst), .I(
        e_init[950]), .Q(ein[950]) );
  DFF \ereg_reg[951]  ( .D(ereg_next[951]), .CLK(clk), .RST(rst), .I(
        e_init[951]), .Q(ein[951]) );
  DFF \ereg_reg[952]  ( .D(ereg_next[952]), .CLK(clk), .RST(rst), .I(
        e_init[952]), .Q(ein[952]) );
  DFF \ereg_reg[953]  ( .D(ereg_next[953]), .CLK(clk), .RST(rst), .I(
        e_init[953]), .Q(ein[953]) );
  DFF \ereg_reg[954]  ( .D(ereg_next[954]), .CLK(clk), .RST(rst), .I(
        e_init[954]), .Q(ein[954]) );
  DFF \ereg_reg[955]  ( .D(ereg_next[955]), .CLK(clk), .RST(rst), .I(
        e_init[955]), .Q(ein[955]) );
  DFF \ereg_reg[956]  ( .D(ereg_next[956]), .CLK(clk), .RST(rst), .I(
        e_init[956]), .Q(ein[956]) );
  DFF \ereg_reg[957]  ( .D(ereg_next[957]), .CLK(clk), .RST(rst), .I(
        e_init[957]), .Q(ein[957]) );
  DFF \ereg_reg[958]  ( .D(ereg_next[958]), .CLK(clk), .RST(rst), .I(
        e_init[958]), .Q(ein[958]) );
  DFF \ereg_reg[959]  ( .D(ereg_next[959]), .CLK(clk), .RST(rst), .I(
        e_init[959]), .Q(ein[959]) );
  DFF \ereg_reg[960]  ( .D(ereg_next[960]), .CLK(clk), .RST(rst), .I(
        e_init[960]), .Q(ein[960]) );
  DFF \ereg_reg[961]  ( .D(ereg_next[961]), .CLK(clk), .RST(rst), .I(
        e_init[961]), .Q(ein[961]) );
  DFF \ereg_reg[962]  ( .D(ereg_next[962]), .CLK(clk), .RST(rst), .I(
        e_init[962]), .Q(ein[962]) );
  DFF \ereg_reg[963]  ( .D(ereg_next[963]), .CLK(clk), .RST(rst), .I(
        e_init[963]), .Q(ein[963]) );
  DFF \ereg_reg[964]  ( .D(ereg_next[964]), .CLK(clk), .RST(rst), .I(
        e_init[964]), .Q(ein[964]) );
  DFF \ereg_reg[965]  ( .D(ereg_next[965]), .CLK(clk), .RST(rst), .I(
        e_init[965]), .Q(ein[965]) );
  DFF \ereg_reg[966]  ( .D(ereg_next[966]), .CLK(clk), .RST(rst), .I(
        e_init[966]), .Q(ein[966]) );
  DFF \ereg_reg[967]  ( .D(ereg_next[967]), .CLK(clk), .RST(rst), .I(
        e_init[967]), .Q(ein[967]) );
  DFF \ereg_reg[968]  ( .D(ereg_next[968]), .CLK(clk), .RST(rst), .I(
        e_init[968]), .Q(ein[968]) );
  DFF \ereg_reg[969]  ( .D(ereg_next[969]), .CLK(clk), .RST(rst), .I(
        e_init[969]), .Q(ein[969]) );
  DFF \ereg_reg[970]  ( .D(ereg_next[970]), .CLK(clk), .RST(rst), .I(
        e_init[970]), .Q(ein[970]) );
  DFF \ereg_reg[971]  ( .D(ereg_next[971]), .CLK(clk), .RST(rst), .I(
        e_init[971]), .Q(ein[971]) );
  DFF \ereg_reg[972]  ( .D(ereg_next[972]), .CLK(clk), .RST(rst), .I(
        e_init[972]), .Q(ein[972]) );
  DFF \ereg_reg[973]  ( .D(ereg_next[973]), .CLK(clk), .RST(rst), .I(
        e_init[973]), .Q(ein[973]) );
  DFF \ereg_reg[974]  ( .D(ereg_next[974]), .CLK(clk), .RST(rst), .I(
        e_init[974]), .Q(ein[974]) );
  DFF \ereg_reg[975]  ( .D(ereg_next[975]), .CLK(clk), .RST(rst), .I(
        e_init[975]), .Q(ein[975]) );
  DFF \ereg_reg[976]  ( .D(ereg_next[976]), .CLK(clk), .RST(rst), .I(
        e_init[976]), .Q(ein[976]) );
  DFF \ereg_reg[977]  ( .D(ereg_next[977]), .CLK(clk), .RST(rst), .I(
        e_init[977]), .Q(ein[977]) );
  DFF \ereg_reg[978]  ( .D(ereg_next[978]), .CLK(clk), .RST(rst), .I(
        e_init[978]), .Q(ein[978]) );
  DFF \ereg_reg[979]  ( .D(ereg_next[979]), .CLK(clk), .RST(rst), .I(
        e_init[979]), .Q(ein[979]) );
  DFF \ereg_reg[980]  ( .D(ereg_next[980]), .CLK(clk), .RST(rst), .I(
        e_init[980]), .Q(ein[980]) );
  DFF \ereg_reg[981]  ( .D(ereg_next[981]), .CLK(clk), .RST(rst), .I(
        e_init[981]), .Q(ein[981]) );
  DFF \ereg_reg[982]  ( .D(ereg_next[982]), .CLK(clk), .RST(rst), .I(
        e_init[982]), .Q(ein[982]) );
  DFF \ereg_reg[983]  ( .D(ereg_next[983]), .CLK(clk), .RST(rst), .I(
        e_init[983]), .Q(ein[983]) );
  DFF \ereg_reg[984]  ( .D(ereg_next[984]), .CLK(clk), .RST(rst), .I(
        e_init[984]), .Q(ein[984]) );
  DFF \ereg_reg[985]  ( .D(ereg_next[985]), .CLK(clk), .RST(rst), .I(
        e_init[985]), .Q(ein[985]) );
  DFF \ereg_reg[986]  ( .D(ereg_next[986]), .CLK(clk), .RST(rst), .I(
        e_init[986]), .Q(ein[986]) );
  DFF \ereg_reg[987]  ( .D(ereg_next[987]), .CLK(clk), .RST(rst), .I(
        e_init[987]), .Q(ein[987]) );
  DFF \ereg_reg[988]  ( .D(ereg_next[988]), .CLK(clk), .RST(rst), .I(
        e_init[988]), .Q(ein[988]) );
  DFF \ereg_reg[989]  ( .D(ereg_next[989]), .CLK(clk), .RST(rst), .I(
        e_init[989]), .Q(ein[989]) );
  DFF \ereg_reg[990]  ( .D(ereg_next[990]), .CLK(clk), .RST(rst), .I(
        e_init[990]), .Q(ein[990]) );
  DFF \ereg_reg[991]  ( .D(ereg_next[991]), .CLK(clk), .RST(rst), .I(
        e_init[991]), .Q(ein[991]) );
  DFF \ereg_reg[992]  ( .D(ereg_next[992]), .CLK(clk), .RST(rst), .I(
        e_init[992]), .Q(ein[992]) );
  DFF \ereg_reg[993]  ( .D(ereg_next[993]), .CLK(clk), .RST(rst), .I(
        e_init[993]), .Q(ein[993]) );
  DFF \ereg_reg[994]  ( .D(ereg_next[994]), .CLK(clk), .RST(rst), .I(
        e_init[994]), .Q(ein[994]) );
  DFF \ereg_reg[995]  ( .D(ereg_next[995]), .CLK(clk), .RST(rst), .I(
        e_init[995]), .Q(ein[995]) );
  DFF \ereg_reg[996]  ( .D(ereg_next[996]), .CLK(clk), .RST(rst), .I(
        e_init[996]), .Q(ein[996]) );
  DFF \ereg_reg[997]  ( .D(ereg_next[997]), .CLK(clk), .RST(rst), .I(
        e_init[997]), .Q(ein[997]) );
  DFF \ereg_reg[998]  ( .D(ereg_next[998]), .CLK(clk), .RST(rst), .I(
        e_init[998]), .Q(ein[998]) );
  DFF \ereg_reg[999]  ( .D(ereg_next[999]), .CLK(clk), .RST(rst), .I(
        e_init[999]), .Q(ein[999]) );
  DFF \ereg_reg[1000]  ( .D(ereg_next[1000]), .CLK(clk), .RST(rst), .I(
        e_init[1000]), .Q(ein[1000]) );
  DFF \ereg_reg[1001]  ( .D(ereg_next[1001]), .CLK(clk), .RST(rst), .I(
        e_init[1001]), .Q(ein[1001]) );
  DFF \ereg_reg[1002]  ( .D(ereg_next[1002]), .CLK(clk), .RST(rst), .I(
        e_init[1002]), .Q(ein[1002]) );
  DFF \ereg_reg[1003]  ( .D(ereg_next[1003]), .CLK(clk), .RST(rst), .I(
        e_init[1003]), .Q(ein[1003]) );
  DFF \ereg_reg[1004]  ( .D(ereg_next[1004]), .CLK(clk), .RST(rst), .I(
        e_init[1004]), .Q(ein[1004]) );
  DFF \ereg_reg[1005]  ( .D(ereg_next[1005]), .CLK(clk), .RST(rst), .I(
        e_init[1005]), .Q(ein[1005]) );
  DFF \ereg_reg[1006]  ( .D(ereg_next[1006]), .CLK(clk), .RST(rst), .I(
        e_init[1006]), .Q(ein[1006]) );
  DFF \ereg_reg[1007]  ( .D(ereg_next[1007]), .CLK(clk), .RST(rst), .I(
        e_init[1007]), .Q(ein[1007]) );
  DFF \ereg_reg[1008]  ( .D(ereg_next[1008]), .CLK(clk), .RST(rst), .I(
        e_init[1008]), .Q(ein[1008]) );
  DFF \ereg_reg[1009]  ( .D(ereg_next[1009]), .CLK(clk), .RST(rst), .I(
        e_init[1009]), .Q(ein[1009]) );
  DFF \ereg_reg[1010]  ( .D(ereg_next[1010]), .CLK(clk), .RST(rst), .I(
        e_init[1010]), .Q(ein[1010]) );
  DFF \ereg_reg[1011]  ( .D(ereg_next[1011]), .CLK(clk), .RST(rst), .I(
        e_init[1011]), .Q(ein[1011]) );
  DFF \ereg_reg[1012]  ( .D(ereg_next[1012]), .CLK(clk), .RST(rst), .I(
        e_init[1012]), .Q(ein[1012]) );
  DFF \ereg_reg[1013]  ( .D(ereg_next[1013]), .CLK(clk), .RST(rst), .I(
        e_init[1013]), .Q(ein[1013]) );
  DFF \ereg_reg[1014]  ( .D(ereg_next[1014]), .CLK(clk), .RST(rst), .I(
        e_init[1014]), .Q(ein[1014]) );
  DFF \ereg_reg[1015]  ( .D(ereg_next[1015]), .CLK(clk), .RST(rst), .I(
        e_init[1015]), .Q(ein[1015]) );
  DFF \ereg_reg[1016]  ( .D(ereg_next[1016]), .CLK(clk), .RST(rst), .I(
        e_init[1016]), .Q(ein[1016]) );
  DFF \ereg_reg[1017]  ( .D(ereg_next[1017]), .CLK(clk), .RST(rst), .I(
        e_init[1017]), .Q(ein[1017]) );
  DFF \ereg_reg[1018]  ( .D(ereg_next[1018]), .CLK(clk), .RST(rst), .I(
        e_init[1018]), .Q(ein[1018]) );
  DFF \ereg_reg[1019]  ( .D(ereg_next[1019]), .CLK(clk), .RST(rst), .I(
        e_init[1019]), .Q(ein[1019]) );
  DFF \ereg_reg[1020]  ( .D(ereg_next[1020]), .CLK(clk), .RST(rst), .I(
        e_init[1020]), .Q(ein[1020]) );
  DFF \ereg_reg[1021]  ( .D(ereg_next[1021]), .CLK(clk), .RST(rst), .I(
        e_init[1021]), .Q(ein[1021]) );
  DFF \ereg_reg[1022]  ( .D(ereg_next[1022]), .CLK(clk), .RST(rst), .I(
        e_init[1022]), .Q(ein[1022]) );
  DFF \ereg_reg[1023]  ( .D(ereg_next[1023]), .CLK(clk), .RST(rst), .I(
        e_init[1023]), .Q(ein[1023]) );
  DFF first_one_reg ( .D(n6), .CLK(clk), .RST(rst), .I(1'b0), .Q(first_one) );
  DFF \creg_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .I(g_init[0]), .Q(
        creg[0]) );
  DFF \creg_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .I(g_init[1]), .Q(
        creg[1]) );
  DFF \creg_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .I(g_init[2]), .Q(
        creg[2]) );
  DFF \creg_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .I(g_init[3]), .Q(
        creg[3]) );
  DFF \creg_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .I(g_init[4]), .Q(
        creg[4]) );
  DFF \creg_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .I(g_init[5]), .Q(
        creg[5]) );
  DFF \creg_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .I(g_init[6]), .Q(
        creg[6]) );
  DFF \creg_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .I(g_init[7]), .Q(
        creg[7]) );
  DFF \creg_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .I(g_init[8]), .Q(
        creg[8]) );
  DFF \creg_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .I(g_init[9]), .Q(
        creg[9]) );
  DFF \creg_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .I(g_init[10]), .Q(
        creg[10]) );
  DFF \creg_reg[11]  ( .D(o[11]), .CLK(clk), .RST(rst), .I(g_init[11]), .Q(
        creg[11]) );
  DFF \creg_reg[12]  ( .D(o[12]), .CLK(clk), .RST(rst), .I(g_init[12]), .Q(
        creg[12]) );
  DFF \creg_reg[13]  ( .D(o[13]), .CLK(clk), .RST(rst), .I(g_init[13]), .Q(
        creg[13]) );
  DFF \creg_reg[14]  ( .D(o[14]), .CLK(clk), .RST(rst), .I(g_init[14]), .Q(
        creg[14]) );
  DFF \creg_reg[15]  ( .D(o[15]), .CLK(clk), .RST(rst), .I(g_init[15]), .Q(
        creg[15]) );
  DFF \creg_reg[16]  ( .D(o[16]), .CLK(clk), .RST(rst), .I(g_init[16]), .Q(
        creg[16]) );
  DFF \creg_reg[17]  ( .D(o[17]), .CLK(clk), .RST(rst), .I(g_init[17]), .Q(
        creg[17]) );
  DFF \creg_reg[18]  ( .D(o[18]), .CLK(clk), .RST(rst), .I(g_init[18]), .Q(
        creg[18]) );
  DFF \creg_reg[19]  ( .D(o[19]), .CLK(clk), .RST(rst), .I(g_init[19]), .Q(
        creg[19]) );
  DFF \creg_reg[20]  ( .D(o[20]), .CLK(clk), .RST(rst), .I(g_init[20]), .Q(
        creg[20]) );
  DFF \creg_reg[21]  ( .D(o[21]), .CLK(clk), .RST(rst), .I(g_init[21]), .Q(
        creg[21]) );
  DFF \creg_reg[22]  ( .D(o[22]), .CLK(clk), .RST(rst), .I(g_init[22]), .Q(
        creg[22]) );
  DFF \creg_reg[23]  ( .D(o[23]), .CLK(clk), .RST(rst), .I(g_init[23]), .Q(
        creg[23]) );
  DFF \creg_reg[24]  ( .D(o[24]), .CLK(clk), .RST(rst), .I(g_init[24]), .Q(
        creg[24]) );
  DFF \creg_reg[25]  ( .D(o[25]), .CLK(clk), .RST(rst), .I(g_init[25]), .Q(
        creg[25]) );
  DFF \creg_reg[26]  ( .D(o[26]), .CLK(clk), .RST(rst), .I(g_init[26]), .Q(
        creg[26]) );
  DFF \creg_reg[27]  ( .D(o[27]), .CLK(clk), .RST(rst), .I(g_init[27]), .Q(
        creg[27]) );
  DFF \creg_reg[28]  ( .D(o[28]), .CLK(clk), .RST(rst), .I(g_init[28]), .Q(
        creg[28]) );
  DFF \creg_reg[29]  ( .D(o[29]), .CLK(clk), .RST(rst), .I(g_init[29]), .Q(
        creg[29]) );
  DFF \creg_reg[30]  ( .D(o[30]), .CLK(clk), .RST(rst), .I(g_init[30]), .Q(
        creg[30]) );
  DFF \creg_reg[31]  ( .D(o[31]), .CLK(clk), .RST(rst), .I(g_init[31]), .Q(
        creg[31]) );
  DFF \creg_reg[32]  ( .D(o[32]), .CLK(clk), .RST(rst), .I(g_init[32]), .Q(
        creg[32]) );
  DFF \creg_reg[33]  ( .D(o[33]), .CLK(clk), .RST(rst), .I(g_init[33]), .Q(
        creg[33]) );
  DFF \creg_reg[34]  ( .D(o[34]), .CLK(clk), .RST(rst), .I(g_init[34]), .Q(
        creg[34]) );
  DFF \creg_reg[35]  ( .D(o[35]), .CLK(clk), .RST(rst), .I(g_init[35]), .Q(
        creg[35]) );
  DFF \creg_reg[36]  ( .D(o[36]), .CLK(clk), .RST(rst), .I(g_init[36]), .Q(
        creg[36]) );
  DFF \creg_reg[37]  ( .D(o[37]), .CLK(clk), .RST(rst), .I(g_init[37]), .Q(
        creg[37]) );
  DFF \creg_reg[38]  ( .D(o[38]), .CLK(clk), .RST(rst), .I(g_init[38]), .Q(
        creg[38]) );
  DFF \creg_reg[39]  ( .D(o[39]), .CLK(clk), .RST(rst), .I(g_init[39]), .Q(
        creg[39]) );
  DFF \creg_reg[40]  ( .D(o[40]), .CLK(clk), .RST(rst), .I(g_init[40]), .Q(
        creg[40]) );
  DFF \creg_reg[41]  ( .D(o[41]), .CLK(clk), .RST(rst), .I(g_init[41]), .Q(
        creg[41]) );
  DFF \creg_reg[42]  ( .D(o[42]), .CLK(clk), .RST(rst), .I(g_init[42]), .Q(
        creg[42]) );
  DFF \creg_reg[43]  ( .D(o[43]), .CLK(clk), .RST(rst), .I(g_init[43]), .Q(
        creg[43]) );
  DFF \creg_reg[44]  ( .D(o[44]), .CLK(clk), .RST(rst), .I(g_init[44]), .Q(
        creg[44]) );
  DFF \creg_reg[45]  ( .D(o[45]), .CLK(clk), .RST(rst), .I(g_init[45]), .Q(
        creg[45]) );
  DFF \creg_reg[46]  ( .D(o[46]), .CLK(clk), .RST(rst), .I(g_init[46]), .Q(
        creg[46]) );
  DFF \creg_reg[47]  ( .D(o[47]), .CLK(clk), .RST(rst), .I(g_init[47]), .Q(
        creg[47]) );
  DFF \creg_reg[48]  ( .D(o[48]), .CLK(clk), .RST(rst), .I(g_init[48]), .Q(
        creg[48]) );
  DFF \creg_reg[49]  ( .D(o[49]), .CLK(clk), .RST(rst), .I(g_init[49]), .Q(
        creg[49]) );
  DFF \creg_reg[50]  ( .D(o[50]), .CLK(clk), .RST(rst), .I(g_init[50]), .Q(
        creg[50]) );
  DFF \creg_reg[51]  ( .D(o[51]), .CLK(clk), .RST(rst), .I(g_init[51]), .Q(
        creg[51]) );
  DFF \creg_reg[52]  ( .D(o[52]), .CLK(clk), .RST(rst), .I(g_init[52]), .Q(
        creg[52]) );
  DFF \creg_reg[53]  ( .D(o[53]), .CLK(clk), .RST(rst), .I(g_init[53]), .Q(
        creg[53]) );
  DFF \creg_reg[54]  ( .D(o[54]), .CLK(clk), .RST(rst), .I(g_init[54]), .Q(
        creg[54]) );
  DFF \creg_reg[55]  ( .D(o[55]), .CLK(clk), .RST(rst), .I(g_init[55]), .Q(
        creg[55]) );
  DFF \creg_reg[56]  ( .D(o[56]), .CLK(clk), .RST(rst), .I(g_init[56]), .Q(
        creg[56]) );
  DFF \creg_reg[57]  ( .D(o[57]), .CLK(clk), .RST(rst), .I(g_init[57]), .Q(
        creg[57]) );
  DFF \creg_reg[58]  ( .D(o[58]), .CLK(clk), .RST(rst), .I(g_init[58]), .Q(
        creg[58]) );
  DFF \creg_reg[59]  ( .D(o[59]), .CLK(clk), .RST(rst), .I(g_init[59]), .Q(
        creg[59]) );
  DFF \creg_reg[60]  ( .D(o[60]), .CLK(clk), .RST(rst), .I(g_init[60]), .Q(
        creg[60]) );
  DFF \creg_reg[61]  ( .D(o[61]), .CLK(clk), .RST(rst), .I(g_init[61]), .Q(
        creg[61]) );
  DFF \creg_reg[62]  ( .D(o[62]), .CLK(clk), .RST(rst), .I(g_init[62]), .Q(
        creg[62]) );
  DFF \creg_reg[63]  ( .D(o[63]), .CLK(clk), .RST(rst), .I(g_init[63]), .Q(
        creg[63]) );
  DFF \creg_reg[64]  ( .D(o[64]), .CLK(clk), .RST(rst), .I(g_init[64]), .Q(
        creg[64]) );
  DFF \creg_reg[65]  ( .D(o[65]), .CLK(clk), .RST(rst), .I(g_init[65]), .Q(
        creg[65]) );
  DFF \creg_reg[66]  ( .D(o[66]), .CLK(clk), .RST(rst), .I(g_init[66]), .Q(
        creg[66]) );
  DFF \creg_reg[67]  ( .D(o[67]), .CLK(clk), .RST(rst), .I(g_init[67]), .Q(
        creg[67]) );
  DFF \creg_reg[68]  ( .D(o[68]), .CLK(clk), .RST(rst), .I(g_init[68]), .Q(
        creg[68]) );
  DFF \creg_reg[69]  ( .D(o[69]), .CLK(clk), .RST(rst), .I(g_init[69]), .Q(
        creg[69]) );
  DFF \creg_reg[70]  ( .D(o[70]), .CLK(clk), .RST(rst), .I(g_init[70]), .Q(
        creg[70]) );
  DFF \creg_reg[71]  ( .D(o[71]), .CLK(clk), .RST(rst), .I(g_init[71]), .Q(
        creg[71]) );
  DFF \creg_reg[72]  ( .D(o[72]), .CLK(clk), .RST(rst), .I(g_init[72]), .Q(
        creg[72]) );
  DFF \creg_reg[73]  ( .D(o[73]), .CLK(clk), .RST(rst), .I(g_init[73]), .Q(
        creg[73]) );
  DFF \creg_reg[74]  ( .D(o[74]), .CLK(clk), .RST(rst), .I(g_init[74]), .Q(
        creg[74]) );
  DFF \creg_reg[75]  ( .D(o[75]), .CLK(clk), .RST(rst), .I(g_init[75]), .Q(
        creg[75]) );
  DFF \creg_reg[76]  ( .D(o[76]), .CLK(clk), .RST(rst), .I(g_init[76]), .Q(
        creg[76]) );
  DFF \creg_reg[77]  ( .D(o[77]), .CLK(clk), .RST(rst), .I(g_init[77]), .Q(
        creg[77]) );
  DFF \creg_reg[78]  ( .D(o[78]), .CLK(clk), .RST(rst), .I(g_init[78]), .Q(
        creg[78]) );
  DFF \creg_reg[79]  ( .D(o[79]), .CLK(clk), .RST(rst), .I(g_init[79]), .Q(
        creg[79]) );
  DFF \creg_reg[80]  ( .D(o[80]), .CLK(clk), .RST(rst), .I(g_init[80]), .Q(
        creg[80]) );
  DFF \creg_reg[81]  ( .D(o[81]), .CLK(clk), .RST(rst), .I(g_init[81]), .Q(
        creg[81]) );
  DFF \creg_reg[82]  ( .D(o[82]), .CLK(clk), .RST(rst), .I(g_init[82]), .Q(
        creg[82]) );
  DFF \creg_reg[83]  ( .D(o[83]), .CLK(clk), .RST(rst), .I(g_init[83]), .Q(
        creg[83]) );
  DFF \creg_reg[84]  ( .D(o[84]), .CLK(clk), .RST(rst), .I(g_init[84]), .Q(
        creg[84]) );
  DFF \creg_reg[85]  ( .D(o[85]), .CLK(clk), .RST(rst), .I(g_init[85]), .Q(
        creg[85]) );
  DFF \creg_reg[86]  ( .D(o[86]), .CLK(clk), .RST(rst), .I(g_init[86]), .Q(
        creg[86]) );
  DFF \creg_reg[87]  ( .D(o[87]), .CLK(clk), .RST(rst), .I(g_init[87]), .Q(
        creg[87]) );
  DFF \creg_reg[88]  ( .D(o[88]), .CLK(clk), .RST(rst), .I(g_init[88]), .Q(
        creg[88]) );
  DFF \creg_reg[89]  ( .D(o[89]), .CLK(clk), .RST(rst), .I(g_init[89]), .Q(
        creg[89]) );
  DFF \creg_reg[90]  ( .D(o[90]), .CLK(clk), .RST(rst), .I(g_init[90]), .Q(
        creg[90]) );
  DFF \creg_reg[91]  ( .D(o[91]), .CLK(clk), .RST(rst), .I(g_init[91]), .Q(
        creg[91]) );
  DFF \creg_reg[92]  ( .D(o[92]), .CLK(clk), .RST(rst), .I(g_init[92]), .Q(
        creg[92]) );
  DFF \creg_reg[93]  ( .D(o[93]), .CLK(clk), .RST(rst), .I(g_init[93]), .Q(
        creg[93]) );
  DFF \creg_reg[94]  ( .D(o[94]), .CLK(clk), .RST(rst), .I(g_init[94]), .Q(
        creg[94]) );
  DFF \creg_reg[95]  ( .D(o[95]), .CLK(clk), .RST(rst), .I(g_init[95]), .Q(
        creg[95]) );
  DFF \creg_reg[96]  ( .D(o[96]), .CLK(clk), .RST(rst), .I(g_init[96]), .Q(
        creg[96]) );
  DFF \creg_reg[97]  ( .D(o[97]), .CLK(clk), .RST(rst), .I(g_init[97]), .Q(
        creg[97]) );
  DFF \creg_reg[98]  ( .D(o[98]), .CLK(clk), .RST(rst), .I(g_init[98]), .Q(
        creg[98]) );
  DFF \creg_reg[99]  ( .D(o[99]), .CLK(clk), .RST(rst), .I(g_init[99]), .Q(
        creg[99]) );
  DFF \creg_reg[100]  ( .D(o[100]), .CLK(clk), .RST(rst), .I(g_init[100]), .Q(
        creg[100]) );
  DFF \creg_reg[101]  ( .D(o[101]), .CLK(clk), .RST(rst), .I(g_init[101]), .Q(
        creg[101]) );
  DFF \creg_reg[102]  ( .D(o[102]), .CLK(clk), .RST(rst), .I(g_init[102]), .Q(
        creg[102]) );
  DFF \creg_reg[103]  ( .D(o[103]), .CLK(clk), .RST(rst), .I(g_init[103]), .Q(
        creg[103]) );
  DFF \creg_reg[104]  ( .D(o[104]), .CLK(clk), .RST(rst), .I(g_init[104]), .Q(
        creg[104]) );
  DFF \creg_reg[105]  ( .D(o[105]), .CLK(clk), .RST(rst), .I(g_init[105]), .Q(
        creg[105]) );
  DFF \creg_reg[106]  ( .D(o[106]), .CLK(clk), .RST(rst), .I(g_init[106]), .Q(
        creg[106]) );
  DFF \creg_reg[107]  ( .D(o[107]), .CLK(clk), .RST(rst), .I(g_init[107]), .Q(
        creg[107]) );
  DFF \creg_reg[108]  ( .D(o[108]), .CLK(clk), .RST(rst), .I(g_init[108]), .Q(
        creg[108]) );
  DFF \creg_reg[109]  ( .D(o[109]), .CLK(clk), .RST(rst), .I(g_init[109]), .Q(
        creg[109]) );
  DFF \creg_reg[110]  ( .D(o[110]), .CLK(clk), .RST(rst), .I(g_init[110]), .Q(
        creg[110]) );
  DFF \creg_reg[111]  ( .D(o[111]), .CLK(clk), .RST(rst), .I(g_init[111]), .Q(
        creg[111]) );
  DFF \creg_reg[112]  ( .D(o[112]), .CLK(clk), .RST(rst), .I(g_init[112]), .Q(
        creg[112]) );
  DFF \creg_reg[113]  ( .D(o[113]), .CLK(clk), .RST(rst), .I(g_init[113]), .Q(
        creg[113]) );
  DFF \creg_reg[114]  ( .D(o[114]), .CLK(clk), .RST(rst), .I(g_init[114]), .Q(
        creg[114]) );
  DFF \creg_reg[115]  ( .D(o[115]), .CLK(clk), .RST(rst), .I(g_init[115]), .Q(
        creg[115]) );
  DFF \creg_reg[116]  ( .D(o[116]), .CLK(clk), .RST(rst), .I(g_init[116]), .Q(
        creg[116]) );
  DFF \creg_reg[117]  ( .D(o[117]), .CLK(clk), .RST(rst), .I(g_init[117]), .Q(
        creg[117]) );
  DFF \creg_reg[118]  ( .D(o[118]), .CLK(clk), .RST(rst), .I(g_init[118]), .Q(
        creg[118]) );
  DFF \creg_reg[119]  ( .D(o[119]), .CLK(clk), .RST(rst), .I(g_init[119]), .Q(
        creg[119]) );
  DFF \creg_reg[120]  ( .D(o[120]), .CLK(clk), .RST(rst), .I(g_init[120]), .Q(
        creg[120]) );
  DFF \creg_reg[121]  ( .D(o[121]), .CLK(clk), .RST(rst), .I(g_init[121]), .Q(
        creg[121]) );
  DFF \creg_reg[122]  ( .D(o[122]), .CLK(clk), .RST(rst), .I(g_init[122]), .Q(
        creg[122]) );
  DFF \creg_reg[123]  ( .D(o[123]), .CLK(clk), .RST(rst), .I(g_init[123]), .Q(
        creg[123]) );
  DFF \creg_reg[124]  ( .D(o[124]), .CLK(clk), .RST(rst), .I(g_init[124]), .Q(
        creg[124]) );
  DFF \creg_reg[125]  ( .D(o[125]), .CLK(clk), .RST(rst), .I(g_init[125]), .Q(
        creg[125]) );
  DFF \creg_reg[126]  ( .D(o[126]), .CLK(clk), .RST(rst), .I(g_init[126]), .Q(
        creg[126]) );
  DFF \creg_reg[127]  ( .D(o[127]), .CLK(clk), .RST(rst), .I(g_init[127]), .Q(
        creg[127]) );
  DFF \creg_reg[128]  ( .D(o[128]), .CLK(clk), .RST(rst), .I(g_init[128]), .Q(
        creg[128]) );
  DFF \creg_reg[129]  ( .D(o[129]), .CLK(clk), .RST(rst), .I(g_init[129]), .Q(
        creg[129]) );
  DFF \creg_reg[130]  ( .D(o[130]), .CLK(clk), .RST(rst), .I(g_init[130]), .Q(
        creg[130]) );
  DFF \creg_reg[131]  ( .D(o[131]), .CLK(clk), .RST(rst), .I(g_init[131]), .Q(
        creg[131]) );
  DFF \creg_reg[132]  ( .D(o[132]), .CLK(clk), .RST(rst), .I(g_init[132]), .Q(
        creg[132]) );
  DFF \creg_reg[133]  ( .D(o[133]), .CLK(clk), .RST(rst), .I(g_init[133]), .Q(
        creg[133]) );
  DFF \creg_reg[134]  ( .D(o[134]), .CLK(clk), .RST(rst), .I(g_init[134]), .Q(
        creg[134]) );
  DFF \creg_reg[135]  ( .D(o[135]), .CLK(clk), .RST(rst), .I(g_init[135]), .Q(
        creg[135]) );
  DFF \creg_reg[136]  ( .D(o[136]), .CLK(clk), .RST(rst), .I(g_init[136]), .Q(
        creg[136]) );
  DFF \creg_reg[137]  ( .D(o[137]), .CLK(clk), .RST(rst), .I(g_init[137]), .Q(
        creg[137]) );
  DFF \creg_reg[138]  ( .D(o[138]), .CLK(clk), .RST(rst), .I(g_init[138]), .Q(
        creg[138]) );
  DFF \creg_reg[139]  ( .D(o[139]), .CLK(clk), .RST(rst), .I(g_init[139]), .Q(
        creg[139]) );
  DFF \creg_reg[140]  ( .D(o[140]), .CLK(clk), .RST(rst), .I(g_init[140]), .Q(
        creg[140]) );
  DFF \creg_reg[141]  ( .D(o[141]), .CLK(clk), .RST(rst), .I(g_init[141]), .Q(
        creg[141]) );
  DFF \creg_reg[142]  ( .D(o[142]), .CLK(clk), .RST(rst), .I(g_init[142]), .Q(
        creg[142]) );
  DFF \creg_reg[143]  ( .D(o[143]), .CLK(clk), .RST(rst), .I(g_init[143]), .Q(
        creg[143]) );
  DFF \creg_reg[144]  ( .D(o[144]), .CLK(clk), .RST(rst), .I(g_init[144]), .Q(
        creg[144]) );
  DFF \creg_reg[145]  ( .D(o[145]), .CLK(clk), .RST(rst), .I(g_init[145]), .Q(
        creg[145]) );
  DFF \creg_reg[146]  ( .D(o[146]), .CLK(clk), .RST(rst), .I(g_init[146]), .Q(
        creg[146]) );
  DFF \creg_reg[147]  ( .D(o[147]), .CLK(clk), .RST(rst), .I(g_init[147]), .Q(
        creg[147]) );
  DFF \creg_reg[148]  ( .D(o[148]), .CLK(clk), .RST(rst), .I(g_init[148]), .Q(
        creg[148]) );
  DFF \creg_reg[149]  ( .D(o[149]), .CLK(clk), .RST(rst), .I(g_init[149]), .Q(
        creg[149]) );
  DFF \creg_reg[150]  ( .D(o[150]), .CLK(clk), .RST(rst), .I(g_init[150]), .Q(
        creg[150]) );
  DFF \creg_reg[151]  ( .D(o[151]), .CLK(clk), .RST(rst), .I(g_init[151]), .Q(
        creg[151]) );
  DFF \creg_reg[152]  ( .D(o[152]), .CLK(clk), .RST(rst), .I(g_init[152]), .Q(
        creg[152]) );
  DFF \creg_reg[153]  ( .D(o[153]), .CLK(clk), .RST(rst), .I(g_init[153]), .Q(
        creg[153]) );
  DFF \creg_reg[154]  ( .D(o[154]), .CLK(clk), .RST(rst), .I(g_init[154]), .Q(
        creg[154]) );
  DFF \creg_reg[155]  ( .D(o[155]), .CLK(clk), .RST(rst), .I(g_init[155]), .Q(
        creg[155]) );
  DFF \creg_reg[156]  ( .D(o[156]), .CLK(clk), .RST(rst), .I(g_init[156]), .Q(
        creg[156]) );
  DFF \creg_reg[157]  ( .D(o[157]), .CLK(clk), .RST(rst), .I(g_init[157]), .Q(
        creg[157]) );
  DFF \creg_reg[158]  ( .D(o[158]), .CLK(clk), .RST(rst), .I(g_init[158]), .Q(
        creg[158]) );
  DFF \creg_reg[159]  ( .D(o[159]), .CLK(clk), .RST(rst), .I(g_init[159]), .Q(
        creg[159]) );
  DFF \creg_reg[160]  ( .D(o[160]), .CLK(clk), .RST(rst), .I(g_init[160]), .Q(
        creg[160]) );
  DFF \creg_reg[161]  ( .D(o[161]), .CLK(clk), .RST(rst), .I(g_init[161]), .Q(
        creg[161]) );
  DFF \creg_reg[162]  ( .D(o[162]), .CLK(clk), .RST(rst), .I(g_init[162]), .Q(
        creg[162]) );
  DFF \creg_reg[163]  ( .D(o[163]), .CLK(clk), .RST(rst), .I(g_init[163]), .Q(
        creg[163]) );
  DFF \creg_reg[164]  ( .D(o[164]), .CLK(clk), .RST(rst), .I(g_init[164]), .Q(
        creg[164]) );
  DFF \creg_reg[165]  ( .D(o[165]), .CLK(clk), .RST(rst), .I(g_init[165]), .Q(
        creg[165]) );
  DFF \creg_reg[166]  ( .D(o[166]), .CLK(clk), .RST(rst), .I(g_init[166]), .Q(
        creg[166]) );
  DFF \creg_reg[167]  ( .D(o[167]), .CLK(clk), .RST(rst), .I(g_init[167]), .Q(
        creg[167]) );
  DFF \creg_reg[168]  ( .D(o[168]), .CLK(clk), .RST(rst), .I(g_init[168]), .Q(
        creg[168]) );
  DFF \creg_reg[169]  ( .D(o[169]), .CLK(clk), .RST(rst), .I(g_init[169]), .Q(
        creg[169]) );
  DFF \creg_reg[170]  ( .D(o[170]), .CLK(clk), .RST(rst), .I(g_init[170]), .Q(
        creg[170]) );
  DFF \creg_reg[171]  ( .D(o[171]), .CLK(clk), .RST(rst), .I(g_init[171]), .Q(
        creg[171]) );
  DFF \creg_reg[172]  ( .D(o[172]), .CLK(clk), .RST(rst), .I(g_init[172]), .Q(
        creg[172]) );
  DFF \creg_reg[173]  ( .D(o[173]), .CLK(clk), .RST(rst), .I(g_init[173]), .Q(
        creg[173]) );
  DFF \creg_reg[174]  ( .D(o[174]), .CLK(clk), .RST(rst), .I(g_init[174]), .Q(
        creg[174]) );
  DFF \creg_reg[175]  ( .D(o[175]), .CLK(clk), .RST(rst), .I(g_init[175]), .Q(
        creg[175]) );
  DFF \creg_reg[176]  ( .D(o[176]), .CLK(clk), .RST(rst), .I(g_init[176]), .Q(
        creg[176]) );
  DFF \creg_reg[177]  ( .D(o[177]), .CLK(clk), .RST(rst), .I(g_init[177]), .Q(
        creg[177]) );
  DFF \creg_reg[178]  ( .D(o[178]), .CLK(clk), .RST(rst), .I(g_init[178]), .Q(
        creg[178]) );
  DFF \creg_reg[179]  ( .D(o[179]), .CLK(clk), .RST(rst), .I(g_init[179]), .Q(
        creg[179]) );
  DFF \creg_reg[180]  ( .D(o[180]), .CLK(clk), .RST(rst), .I(g_init[180]), .Q(
        creg[180]) );
  DFF \creg_reg[181]  ( .D(o[181]), .CLK(clk), .RST(rst), .I(g_init[181]), .Q(
        creg[181]) );
  DFF \creg_reg[182]  ( .D(o[182]), .CLK(clk), .RST(rst), .I(g_init[182]), .Q(
        creg[182]) );
  DFF \creg_reg[183]  ( .D(o[183]), .CLK(clk), .RST(rst), .I(g_init[183]), .Q(
        creg[183]) );
  DFF \creg_reg[184]  ( .D(o[184]), .CLK(clk), .RST(rst), .I(g_init[184]), .Q(
        creg[184]) );
  DFF \creg_reg[185]  ( .D(o[185]), .CLK(clk), .RST(rst), .I(g_init[185]), .Q(
        creg[185]) );
  DFF \creg_reg[186]  ( .D(o[186]), .CLK(clk), .RST(rst), .I(g_init[186]), .Q(
        creg[186]) );
  DFF \creg_reg[187]  ( .D(o[187]), .CLK(clk), .RST(rst), .I(g_init[187]), .Q(
        creg[187]) );
  DFF \creg_reg[188]  ( .D(o[188]), .CLK(clk), .RST(rst), .I(g_init[188]), .Q(
        creg[188]) );
  DFF \creg_reg[189]  ( .D(o[189]), .CLK(clk), .RST(rst), .I(g_init[189]), .Q(
        creg[189]) );
  DFF \creg_reg[190]  ( .D(o[190]), .CLK(clk), .RST(rst), .I(g_init[190]), .Q(
        creg[190]) );
  DFF \creg_reg[191]  ( .D(o[191]), .CLK(clk), .RST(rst), .I(g_init[191]), .Q(
        creg[191]) );
  DFF \creg_reg[192]  ( .D(o[192]), .CLK(clk), .RST(rst), .I(g_init[192]), .Q(
        creg[192]) );
  DFF \creg_reg[193]  ( .D(o[193]), .CLK(clk), .RST(rst), .I(g_init[193]), .Q(
        creg[193]) );
  DFF \creg_reg[194]  ( .D(o[194]), .CLK(clk), .RST(rst), .I(g_init[194]), .Q(
        creg[194]) );
  DFF \creg_reg[195]  ( .D(o[195]), .CLK(clk), .RST(rst), .I(g_init[195]), .Q(
        creg[195]) );
  DFF \creg_reg[196]  ( .D(o[196]), .CLK(clk), .RST(rst), .I(g_init[196]), .Q(
        creg[196]) );
  DFF \creg_reg[197]  ( .D(o[197]), .CLK(clk), .RST(rst), .I(g_init[197]), .Q(
        creg[197]) );
  DFF \creg_reg[198]  ( .D(o[198]), .CLK(clk), .RST(rst), .I(g_init[198]), .Q(
        creg[198]) );
  DFF \creg_reg[199]  ( .D(o[199]), .CLK(clk), .RST(rst), .I(g_init[199]), .Q(
        creg[199]) );
  DFF \creg_reg[200]  ( .D(o[200]), .CLK(clk), .RST(rst), .I(g_init[200]), .Q(
        creg[200]) );
  DFF \creg_reg[201]  ( .D(o[201]), .CLK(clk), .RST(rst), .I(g_init[201]), .Q(
        creg[201]) );
  DFF \creg_reg[202]  ( .D(o[202]), .CLK(clk), .RST(rst), .I(g_init[202]), .Q(
        creg[202]) );
  DFF \creg_reg[203]  ( .D(o[203]), .CLK(clk), .RST(rst), .I(g_init[203]), .Q(
        creg[203]) );
  DFF \creg_reg[204]  ( .D(o[204]), .CLK(clk), .RST(rst), .I(g_init[204]), .Q(
        creg[204]) );
  DFF \creg_reg[205]  ( .D(o[205]), .CLK(clk), .RST(rst), .I(g_init[205]), .Q(
        creg[205]) );
  DFF \creg_reg[206]  ( .D(o[206]), .CLK(clk), .RST(rst), .I(g_init[206]), .Q(
        creg[206]) );
  DFF \creg_reg[207]  ( .D(o[207]), .CLK(clk), .RST(rst), .I(g_init[207]), .Q(
        creg[207]) );
  DFF \creg_reg[208]  ( .D(o[208]), .CLK(clk), .RST(rst), .I(g_init[208]), .Q(
        creg[208]) );
  DFF \creg_reg[209]  ( .D(o[209]), .CLK(clk), .RST(rst), .I(g_init[209]), .Q(
        creg[209]) );
  DFF \creg_reg[210]  ( .D(o[210]), .CLK(clk), .RST(rst), .I(g_init[210]), .Q(
        creg[210]) );
  DFF \creg_reg[211]  ( .D(o[211]), .CLK(clk), .RST(rst), .I(g_init[211]), .Q(
        creg[211]) );
  DFF \creg_reg[212]  ( .D(o[212]), .CLK(clk), .RST(rst), .I(g_init[212]), .Q(
        creg[212]) );
  DFF \creg_reg[213]  ( .D(o[213]), .CLK(clk), .RST(rst), .I(g_init[213]), .Q(
        creg[213]) );
  DFF \creg_reg[214]  ( .D(o[214]), .CLK(clk), .RST(rst), .I(g_init[214]), .Q(
        creg[214]) );
  DFF \creg_reg[215]  ( .D(o[215]), .CLK(clk), .RST(rst), .I(g_init[215]), .Q(
        creg[215]) );
  DFF \creg_reg[216]  ( .D(o[216]), .CLK(clk), .RST(rst), .I(g_init[216]), .Q(
        creg[216]) );
  DFF \creg_reg[217]  ( .D(o[217]), .CLK(clk), .RST(rst), .I(g_init[217]), .Q(
        creg[217]) );
  DFF \creg_reg[218]  ( .D(o[218]), .CLK(clk), .RST(rst), .I(g_init[218]), .Q(
        creg[218]) );
  DFF \creg_reg[219]  ( .D(o[219]), .CLK(clk), .RST(rst), .I(g_init[219]), .Q(
        creg[219]) );
  DFF \creg_reg[220]  ( .D(o[220]), .CLK(clk), .RST(rst), .I(g_init[220]), .Q(
        creg[220]) );
  DFF \creg_reg[221]  ( .D(o[221]), .CLK(clk), .RST(rst), .I(g_init[221]), .Q(
        creg[221]) );
  DFF \creg_reg[222]  ( .D(o[222]), .CLK(clk), .RST(rst), .I(g_init[222]), .Q(
        creg[222]) );
  DFF \creg_reg[223]  ( .D(o[223]), .CLK(clk), .RST(rst), .I(g_init[223]), .Q(
        creg[223]) );
  DFF \creg_reg[224]  ( .D(o[224]), .CLK(clk), .RST(rst), .I(g_init[224]), .Q(
        creg[224]) );
  DFF \creg_reg[225]  ( .D(o[225]), .CLK(clk), .RST(rst), .I(g_init[225]), .Q(
        creg[225]) );
  DFF \creg_reg[226]  ( .D(o[226]), .CLK(clk), .RST(rst), .I(g_init[226]), .Q(
        creg[226]) );
  DFF \creg_reg[227]  ( .D(o[227]), .CLK(clk), .RST(rst), .I(g_init[227]), .Q(
        creg[227]) );
  DFF \creg_reg[228]  ( .D(o[228]), .CLK(clk), .RST(rst), .I(g_init[228]), .Q(
        creg[228]) );
  DFF \creg_reg[229]  ( .D(o[229]), .CLK(clk), .RST(rst), .I(g_init[229]), .Q(
        creg[229]) );
  DFF \creg_reg[230]  ( .D(o[230]), .CLK(clk), .RST(rst), .I(g_init[230]), .Q(
        creg[230]) );
  DFF \creg_reg[231]  ( .D(o[231]), .CLK(clk), .RST(rst), .I(g_init[231]), .Q(
        creg[231]) );
  DFF \creg_reg[232]  ( .D(o[232]), .CLK(clk), .RST(rst), .I(g_init[232]), .Q(
        creg[232]) );
  DFF \creg_reg[233]  ( .D(o[233]), .CLK(clk), .RST(rst), .I(g_init[233]), .Q(
        creg[233]) );
  DFF \creg_reg[234]  ( .D(o[234]), .CLK(clk), .RST(rst), .I(g_init[234]), .Q(
        creg[234]) );
  DFF \creg_reg[235]  ( .D(o[235]), .CLK(clk), .RST(rst), .I(g_init[235]), .Q(
        creg[235]) );
  DFF \creg_reg[236]  ( .D(o[236]), .CLK(clk), .RST(rst), .I(g_init[236]), .Q(
        creg[236]) );
  DFF \creg_reg[237]  ( .D(o[237]), .CLK(clk), .RST(rst), .I(g_init[237]), .Q(
        creg[237]) );
  DFF \creg_reg[238]  ( .D(o[238]), .CLK(clk), .RST(rst), .I(g_init[238]), .Q(
        creg[238]) );
  DFF \creg_reg[239]  ( .D(o[239]), .CLK(clk), .RST(rst), .I(g_init[239]), .Q(
        creg[239]) );
  DFF \creg_reg[240]  ( .D(o[240]), .CLK(clk), .RST(rst), .I(g_init[240]), .Q(
        creg[240]) );
  DFF \creg_reg[241]  ( .D(o[241]), .CLK(clk), .RST(rst), .I(g_init[241]), .Q(
        creg[241]) );
  DFF \creg_reg[242]  ( .D(o[242]), .CLK(clk), .RST(rst), .I(g_init[242]), .Q(
        creg[242]) );
  DFF \creg_reg[243]  ( .D(o[243]), .CLK(clk), .RST(rst), .I(g_init[243]), .Q(
        creg[243]) );
  DFF \creg_reg[244]  ( .D(o[244]), .CLK(clk), .RST(rst), .I(g_init[244]), .Q(
        creg[244]) );
  DFF \creg_reg[245]  ( .D(o[245]), .CLK(clk), .RST(rst), .I(g_init[245]), .Q(
        creg[245]) );
  DFF \creg_reg[246]  ( .D(o[246]), .CLK(clk), .RST(rst), .I(g_init[246]), .Q(
        creg[246]) );
  DFF \creg_reg[247]  ( .D(o[247]), .CLK(clk), .RST(rst), .I(g_init[247]), .Q(
        creg[247]) );
  DFF \creg_reg[248]  ( .D(o[248]), .CLK(clk), .RST(rst), .I(g_init[248]), .Q(
        creg[248]) );
  DFF \creg_reg[249]  ( .D(o[249]), .CLK(clk), .RST(rst), .I(g_init[249]), .Q(
        creg[249]) );
  DFF \creg_reg[250]  ( .D(o[250]), .CLK(clk), .RST(rst), .I(g_init[250]), .Q(
        creg[250]) );
  DFF \creg_reg[251]  ( .D(o[251]), .CLK(clk), .RST(rst), .I(g_init[251]), .Q(
        creg[251]) );
  DFF \creg_reg[252]  ( .D(o[252]), .CLK(clk), .RST(rst), .I(g_init[252]), .Q(
        creg[252]) );
  DFF \creg_reg[253]  ( .D(o[253]), .CLK(clk), .RST(rst), .I(g_init[253]), .Q(
        creg[253]) );
  DFF \creg_reg[254]  ( .D(o[254]), .CLK(clk), .RST(rst), .I(g_init[254]), .Q(
        creg[254]) );
  DFF \creg_reg[255]  ( .D(o[255]), .CLK(clk), .RST(rst), .I(g_init[255]), .Q(
        creg[255]) );
  DFF \creg_reg[256]  ( .D(o[256]), .CLK(clk), .RST(rst), .I(g_init[256]), .Q(
        creg[256]) );
  DFF \creg_reg[257]  ( .D(o[257]), .CLK(clk), .RST(rst), .I(g_init[257]), .Q(
        creg[257]) );
  DFF \creg_reg[258]  ( .D(o[258]), .CLK(clk), .RST(rst), .I(g_init[258]), .Q(
        creg[258]) );
  DFF \creg_reg[259]  ( .D(o[259]), .CLK(clk), .RST(rst), .I(g_init[259]), .Q(
        creg[259]) );
  DFF \creg_reg[260]  ( .D(o[260]), .CLK(clk), .RST(rst), .I(g_init[260]), .Q(
        creg[260]) );
  DFF \creg_reg[261]  ( .D(o[261]), .CLK(clk), .RST(rst), .I(g_init[261]), .Q(
        creg[261]) );
  DFF \creg_reg[262]  ( .D(o[262]), .CLK(clk), .RST(rst), .I(g_init[262]), .Q(
        creg[262]) );
  DFF \creg_reg[263]  ( .D(o[263]), .CLK(clk), .RST(rst), .I(g_init[263]), .Q(
        creg[263]) );
  DFF \creg_reg[264]  ( .D(o[264]), .CLK(clk), .RST(rst), .I(g_init[264]), .Q(
        creg[264]) );
  DFF \creg_reg[265]  ( .D(o[265]), .CLK(clk), .RST(rst), .I(g_init[265]), .Q(
        creg[265]) );
  DFF \creg_reg[266]  ( .D(o[266]), .CLK(clk), .RST(rst), .I(g_init[266]), .Q(
        creg[266]) );
  DFF \creg_reg[267]  ( .D(o[267]), .CLK(clk), .RST(rst), .I(g_init[267]), .Q(
        creg[267]) );
  DFF \creg_reg[268]  ( .D(o[268]), .CLK(clk), .RST(rst), .I(g_init[268]), .Q(
        creg[268]) );
  DFF \creg_reg[269]  ( .D(o[269]), .CLK(clk), .RST(rst), .I(g_init[269]), .Q(
        creg[269]) );
  DFF \creg_reg[270]  ( .D(o[270]), .CLK(clk), .RST(rst), .I(g_init[270]), .Q(
        creg[270]) );
  DFF \creg_reg[271]  ( .D(o[271]), .CLK(clk), .RST(rst), .I(g_init[271]), .Q(
        creg[271]) );
  DFF \creg_reg[272]  ( .D(o[272]), .CLK(clk), .RST(rst), .I(g_init[272]), .Q(
        creg[272]) );
  DFF \creg_reg[273]  ( .D(o[273]), .CLK(clk), .RST(rst), .I(g_init[273]), .Q(
        creg[273]) );
  DFF \creg_reg[274]  ( .D(o[274]), .CLK(clk), .RST(rst), .I(g_init[274]), .Q(
        creg[274]) );
  DFF \creg_reg[275]  ( .D(o[275]), .CLK(clk), .RST(rst), .I(g_init[275]), .Q(
        creg[275]) );
  DFF \creg_reg[276]  ( .D(o[276]), .CLK(clk), .RST(rst), .I(g_init[276]), .Q(
        creg[276]) );
  DFF \creg_reg[277]  ( .D(o[277]), .CLK(clk), .RST(rst), .I(g_init[277]), .Q(
        creg[277]) );
  DFF \creg_reg[278]  ( .D(o[278]), .CLK(clk), .RST(rst), .I(g_init[278]), .Q(
        creg[278]) );
  DFF \creg_reg[279]  ( .D(o[279]), .CLK(clk), .RST(rst), .I(g_init[279]), .Q(
        creg[279]) );
  DFF \creg_reg[280]  ( .D(o[280]), .CLK(clk), .RST(rst), .I(g_init[280]), .Q(
        creg[280]) );
  DFF \creg_reg[281]  ( .D(o[281]), .CLK(clk), .RST(rst), .I(g_init[281]), .Q(
        creg[281]) );
  DFF \creg_reg[282]  ( .D(o[282]), .CLK(clk), .RST(rst), .I(g_init[282]), .Q(
        creg[282]) );
  DFF \creg_reg[283]  ( .D(o[283]), .CLK(clk), .RST(rst), .I(g_init[283]), .Q(
        creg[283]) );
  DFF \creg_reg[284]  ( .D(o[284]), .CLK(clk), .RST(rst), .I(g_init[284]), .Q(
        creg[284]) );
  DFF \creg_reg[285]  ( .D(o[285]), .CLK(clk), .RST(rst), .I(g_init[285]), .Q(
        creg[285]) );
  DFF \creg_reg[286]  ( .D(o[286]), .CLK(clk), .RST(rst), .I(g_init[286]), .Q(
        creg[286]) );
  DFF \creg_reg[287]  ( .D(o[287]), .CLK(clk), .RST(rst), .I(g_init[287]), .Q(
        creg[287]) );
  DFF \creg_reg[288]  ( .D(o[288]), .CLK(clk), .RST(rst), .I(g_init[288]), .Q(
        creg[288]) );
  DFF \creg_reg[289]  ( .D(o[289]), .CLK(clk), .RST(rst), .I(g_init[289]), .Q(
        creg[289]) );
  DFF \creg_reg[290]  ( .D(o[290]), .CLK(clk), .RST(rst), .I(g_init[290]), .Q(
        creg[290]) );
  DFF \creg_reg[291]  ( .D(o[291]), .CLK(clk), .RST(rst), .I(g_init[291]), .Q(
        creg[291]) );
  DFF \creg_reg[292]  ( .D(o[292]), .CLK(clk), .RST(rst), .I(g_init[292]), .Q(
        creg[292]) );
  DFF \creg_reg[293]  ( .D(o[293]), .CLK(clk), .RST(rst), .I(g_init[293]), .Q(
        creg[293]) );
  DFF \creg_reg[294]  ( .D(o[294]), .CLK(clk), .RST(rst), .I(g_init[294]), .Q(
        creg[294]) );
  DFF \creg_reg[295]  ( .D(o[295]), .CLK(clk), .RST(rst), .I(g_init[295]), .Q(
        creg[295]) );
  DFF \creg_reg[296]  ( .D(o[296]), .CLK(clk), .RST(rst), .I(g_init[296]), .Q(
        creg[296]) );
  DFF \creg_reg[297]  ( .D(o[297]), .CLK(clk), .RST(rst), .I(g_init[297]), .Q(
        creg[297]) );
  DFF \creg_reg[298]  ( .D(o[298]), .CLK(clk), .RST(rst), .I(g_init[298]), .Q(
        creg[298]) );
  DFF \creg_reg[299]  ( .D(o[299]), .CLK(clk), .RST(rst), .I(g_init[299]), .Q(
        creg[299]) );
  DFF \creg_reg[300]  ( .D(o[300]), .CLK(clk), .RST(rst), .I(g_init[300]), .Q(
        creg[300]) );
  DFF \creg_reg[301]  ( .D(o[301]), .CLK(clk), .RST(rst), .I(g_init[301]), .Q(
        creg[301]) );
  DFF \creg_reg[302]  ( .D(o[302]), .CLK(clk), .RST(rst), .I(g_init[302]), .Q(
        creg[302]) );
  DFF \creg_reg[303]  ( .D(o[303]), .CLK(clk), .RST(rst), .I(g_init[303]), .Q(
        creg[303]) );
  DFF \creg_reg[304]  ( .D(o[304]), .CLK(clk), .RST(rst), .I(g_init[304]), .Q(
        creg[304]) );
  DFF \creg_reg[305]  ( .D(o[305]), .CLK(clk), .RST(rst), .I(g_init[305]), .Q(
        creg[305]) );
  DFF \creg_reg[306]  ( .D(o[306]), .CLK(clk), .RST(rst), .I(g_init[306]), .Q(
        creg[306]) );
  DFF \creg_reg[307]  ( .D(o[307]), .CLK(clk), .RST(rst), .I(g_init[307]), .Q(
        creg[307]) );
  DFF \creg_reg[308]  ( .D(o[308]), .CLK(clk), .RST(rst), .I(g_init[308]), .Q(
        creg[308]) );
  DFF \creg_reg[309]  ( .D(o[309]), .CLK(clk), .RST(rst), .I(g_init[309]), .Q(
        creg[309]) );
  DFF \creg_reg[310]  ( .D(o[310]), .CLK(clk), .RST(rst), .I(g_init[310]), .Q(
        creg[310]) );
  DFF \creg_reg[311]  ( .D(o[311]), .CLK(clk), .RST(rst), .I(g_init[311]), .Q(
        creg[311]) );
  DFF \creg_reg[312]  ( .D(o[312]), .CLK(clk), .RST(rst), .I(g_init[312]), .Q(
        creg[312]) );
  DFF \creg_reg[313]  ( .D(o[313]), .CLK(clk), .RST(rst), .I(g_init[313]), .Q(
        creg[313]) );
  DFF \creg_reg[314]  ( .D(o[314]), .CLK(clk), .RST(rst), .I(g_init[314]), .Q(
        creg[314]) );
  DFF \creg_reg[315]  ( .D(o[315]), .CLK(clk), .RST(rst), .I(g_init[315]), .Q(
        creg[315]) );
  DFF \creg_reg[316]  ( .D(o[316]), .CLK(clk), .RST(rst), .I(g_init[316]), .Q(
        creg[316]) );
  DFF \creg_reg[317]  ( .D(o[317]), .CLK(clk), .RST(rst), .I(g_init[317]), .Q(
        creg[317]) );
  DFF \creg_reg[318]  ( .D(o[318]), .CLK(clk), .RST(rst), .I(g_init[318]), .Q(
        creg[318]) );
  DFF \creg_reg[319]  ( .D(o[319]), .CLK(clk), .RST(rst), .I(g_init[319]), .Q(
        creg[319]) );
  DFF \creg_reg[320]  ( .D(o[320]), .CLK(clk), .RST(rst), .I(g_init[320]), .Q(
        creg[320]) );
  DFF \creg_reg[321]  ( .D(o[321]), .CLK(clk), .RST(rst), .I(g_init[321]), .Q(
        creg[321]) );
  DFF \creg_reg[322]  ( .D(o[322]), .CLK(clk), .RST(rst), .I(g_init[322]), .Q(
        creg[322]) );
  DFF \creg_reg[323]  ( .D(o[323]), .CLK(clk), .RST(rst), .I(g_init[323]), .Q(
        creg[323]) );
  DFF \creg_reg[324]  ( .D(o[324]), .CLK(clk), .RST(rst), .I(g_init[324]), .Q(
        creg[324]) );
  DFF \creg_reg[325]  ( .D(o[325]), .CLK(clk), .RST(rst), .I(g_init[325]), .Q(
        creg[325]) );
  DFF \creg_reg[326]  ( .D(o[326]), .CLK(clk), .RST(rst), .I(g_init[326]), .Q(
        creg[326]) );
  DFF \creg_reg[327]  ( .D(o[327]), .CLK(clk), .RST(rst), .I(g_init[327]), .Q(
        creg[327]) );
  DFF \creg_reg[328]  ( .D(o[328]), .CLK(clk), .RST(rst), .I(g_init[328]), .Q(
        creg[328]) );
  DFF \creg_reg[329]  ( .D(o[329]), .CLK(clk), .RST(rst), .I(g_init[329]), .Q(
        creg[329]) );
  DFF \creg_reg[330]  ( .D(o[330]), .CLK(clk), .RST(rst), .I(g_init[330]), .Q(
        creg[330]) );
  DFF \creg_reg[331]  ( .D(o[331]), .CLK(clk), .RST(rst), .I(g_init[331]), .Q(
        creg[331]) );
  DFF \creg_reg[332]  ( .D(o[332]), .CLK(clk), .RST(rst), .I(g_init[332]), .Q(
        creg[332]) );
  DFF \creg_reg[333]  ( .D(o[333]), .CLK(clk), .RST(rst), .I(g_init[333]), .Q(
        creg[333]) );
  DFF \creg_reg[334]  ( .D(o[334]), .CLK(clk), .RST(rst), .I(g_init[334]), .Q(
        creg[334]) );
  DFF \creg_reg[335]  ( .D(o[335]), .CLK(clk), .RST(rst), .I(g_init[335]), .Q(
        creg[335]) );
  DFF \creg_reg[336]  ( .D(o[336]), .CLK(clk), .RST(rst), .I(g_init[336]), .Q(
        creg[336]) );
  DFF \creg_reg[337]  ( .D(o[337]), .CLK(clk), .RST(rst), .I(g_init[337]), .Q(
        creg[337]) );
  DFF \creg_reg[338]  ( .D(o[338]), .CLK(clk), .RST(rst), .I(g_init[338]), .Q(
        creg[338]) );
  DFF \creg_reg[339]  ( .D(o[339]), .CLK(clk), .RST(rst), .I(g_init[339]), .Q(
        creg[339]) );
  DFF \creg_reg[340]  ( .D(o[340]), .CLK(clk), .RST(rst), .I(g_init[340]), .Q(
        creg[340]) );
  DFF \creg_reg[341]  ( .D(o[341]), .CLK(clk), .RST(rst), .I(g_init[341]), .Q(
        creg[341]) );
  DFF \creg_reg[342]  ( .D(o[342]), .CLK(clk), .RST(rst), .I(g_init[342]), .Q(
        creg[342]) );
  DFF \creg_reg[343]  ( .D(o[343]), .CLK(clk), .RST(rst), .I(g_init[343]), .Q(
        creg[343]) );
  DFF \creg_reg[344]  ( .D(o[344]), .CLK(clk), .RST(rst), .I(g_init[344]), .Q(
        creg[344]) );
  DFF \creg_reg[345]  ( .D(o[345]), .CLK(clk), .RST(rst), .I(g_init[345]), .Q(
        creg[345]) );
  DFF \creg_reg[346]  ( .D(o[346]), .CLK(clk), .RST(rst), .I(g_init[346]), .Q(
        creg[346]) );
  DFF \creg_reg[347]  ( .D(o[347]), .CLK(clk), .RST(rst), .I(g_init[347]), .Q(
        creg[347]) );
  DFF \creg_reg[348]  ( .D(o[348]), .CLK(clk), .RST(rst), .I(g_init[348]), .Q(
        creg[348]) );
  DFF \creg_reg[349]  ( .D(o[349]), .CLK(clk), .RST(rst), .I(g_init[349]), .Q(
        creg[349]) );
  DFF \creg_reg[350]  ( .D(o[350]), .CLK(clk), .RST(rst), .I(g_init[350]), .Q(
        creg[350]) );
  DFF \creg_reg[351]  ( .D(o[351]), .CLK(clk), .RST(rst), .I(g_init[351]), .Q(
        creg[351]) );
  DFF \creg_reg[352]  ( .D(o[352]), .CLK(clk), .RST(rst), .I(g_init[352]), .Q(
        creg[352]) );
  DFF \creg_reg[353]  ( .D(o[353]), .CLK(clk), .RST(rst), .I(g_init[353]), .Q(
        creg[353]) );
  DFF \creg_reg[354]  ( .D(o[354]), .CLK(clk), .RST(rst), .I(g_init[354]), .Q(
        creg[354]) );
  DFF \creg_reg[355]  ( .D(o[355]), .CLK(clk), .RST(rst), .I(g_init[355]), .Q(
        creg[355]) );
  DFF \creg_reg[356]  ( .D(o[356]), .CLK(clk), .RST(rst), .I(g_init[356]), .Q(
        creg[356]) );
  DFF \creg_reg[357]  ( .D(o[357]), .CLK(clk), .RST(rst), .I(g_init[357]), .Q(
        creg[357]) );
  DFF \creg_reg[358]  ( .D(o[358]), .CLK(clk), .RST(rst), .I(g_init[358]), .Q(
        creg[358]) );
  DFF \creg_reg[359]  ( .D(o[359]), .CLK(clk), .RST(rst), .I(g_init[359]), .Q(
        creg[359]) );
  DFF \creg_reg[360]  ( .D(o[360]), .CLK(clk), .RST(rst), .I(g_init[360]), .Q(
        creg[360]) );
  DFF \creg_reg[361]  ( .D(o[361]), .CLK(clk), .RST(rst), .I(g_init[361]), .Q(
        creg[361]) );
  DFF \creg_reg[362]  ( .D(o[362]), .CLK(clk), .RST(rst), .I(g_init[362]), .Q(
        creg[362]) );
  DFF \creg_reg[363]  ( .D(o[363]), .CLK(clk), .RST(rst), .I(g_init[363]), .Q(
        creg[363]) );
  DFF \creg_reg[364]  ( .D(o[364]), .CLK(clk), .RST(rst), .I(g_init[364]), .Q(
        creg[364]) );
  DFF \creg_reg[365]  ( .D(o[365]), .CLK(clk), .RST(rst), .I(g_init[365]), .Q(
        creg[365]) );
  DFF \creg_reg[366]  ( .D(o[366]), .CLK(clk), .RST(rst), .I(g_init[366]), .Q(
        creg[366]) );
  DFF \creg_reg[367]  ( .D(o[367]), .CLK(clk), .RST(rst), .I(g_init[367]), .Q(
        creg[367]) );
  DFF \creg_reg[368]  ( .D(o[368]), .CLK(clk), .RST(rst), .I(g_init[368]), .Q(
        creg[368]) );
  DFF \creg_reg[369]  ( .D(o[369]), .CLK(clk), .RST(rst), .I(g_init[369]), .Q(
        creg[369]) );
  DFF \creg_reg[370]  ( .D(o[370]), .CLK(clk), .RST(rst), .I(g_init[370]), .Q(
        creg[370]) );
  DFF \creg_reg[371]  ( .D(o[371]), .CLK(clk), .RST(rst), .I(g_init[371]), .Q(
        creg[371]) );
  DFF \creg_reg[372]  ( .D(o[372]), .CLK(clk), .RST(rst), .I(g_init[372]), .Q(
        creg[372]) );
  DFF \creg_reg[373]  ( .D(o[373]), .CLK(clk), .RST(rst), .I(g_init[373]), .Q(
        creg[373]) );
  DFF \creg_reg[374]  ( .D(o[374]), .CLK(clk), .RST(rst), .I(g_init[374]), .Q(
        creg[374]) );
  DFF \creg_reg[375]  ( .D(o[375]), .CLK(clk), .RST(rst), .I(g_init[375]), .Q(
        creg[375]) );
  DFF \creg_reg[376]  ( .D(o[376]), .CLK(clk), .RST(rst), .I(g_init[376]), .Q(
        creg[376]) );
  DFF \creg_reg[377]  ( .D(o[377]), .CLK(clk), .RST(rst), .I(g_init[377]), .Q(
        creg[377]) );
  DFF \creg_reg[378]  ( .D(o[378]), .CLK(clk), .RST(rst), .I(g_init[378]), .Q(
        creg[378]) );
  DFF \creg_reg[379]  ( .D(o[379]), .CLK(clk), .RST(rst), .I(g_init[379]), .Q(
        creg[379]) );
  DFF \creg_reg[380]  ( .D(o[380]), .CLK(clk), .RST(rst), .I(g_init[380]), .Q(
        creg[380]) );
  DFF \creg_reg[381]  ( .D(o[381]), .CLK(clk), .RST(rst), .I(g_init[381]), .Q(
        creg[381]) );
  DFF \creg_reg[382]  ( .D(o[382]), .CLK(clk), .RST(rst), .I(g_init[382]), .Q(
        creg[382]) );
  DFF \creg_reg[383]  ( .D(o[383]), .CLK(clk), .RST(rst), .I(g_init[383]), .Q(
        creg[383]) );
  DFF \creg_reg[384]  ( .D(o[384]), .CLK(clk), .RST(rst), .I(g_init[384]), .Q(
        creg[384]) );
  DFF \creg_reg[385]  ( .D(o[385]), .CLK(clk), .RST(rst), .I(g_init[385]), .Q(
        creg[385]) );
  DFF \creg_reg[386]  ( .D(o[386]), .CLK(clk), .RST(rst), .I(g_init[386]), .Q(
        creg[386]) );
  DFF \creg_reg[387]  ( .D(o[387]), .CLK(clk), .RST(rst), .I(g_init[387]), .Q(
        creg[387]) );
  DFF \creg_reg[388]  ( .D(o[388]), .CLK(clk), .RST(rst), .I(g_init[388]), .Q(
        creg[388]) );
  DFF \creg_reg[389]  ( .D(o[389]), .CLK(clk), .RST(rst), .I(g_init[389]), .Q(
        creg[389]) );
  DFF \creg_reg[390]  ( .D(o[390]), .CLK(clk), .RST(rst), .I(g_init[390]), .Q(
        creg[390]) );
  DFF \creg_reg[391]  ( .D(o[391]), .CLK(clk), .RST(rst), .I(g_init[391]), .Q(
        creg[391]) );
  DFF \creg_reg[392]  ( .D(o[392]), .CLK(clk), .RST(rst), .I(g_init[392]), .Q(
        creg[392]) );
  DFF \creg_reg[393]  ( .D(o[393]), .CLK(clk), .RST(rst), .I(g_init[393]), .Q(
        creg[393]) );
  DFF \creg_reg[394]  ( .D(o[394]), .CLK(clk), .RST(rst), .I(g_init[394]), .Q(
        creg[394]) );
  DFF \creg_reg[395]  ( .D(o[395]), .CLK(clk), .RST(rst), .I(g_init[395]), .Q(
        creg[395]) );
  DFF \creg_reg[396]  ( .D(o[396]), .CLK(clk), .RST(rst), .I(g_init[396]), .Q(
        creg[396]) );
  DFF \creg_reg[397]  ( .D(o[397]), .CLK(clk), .RST(rst), .I(g_init[397]), .Q(
        creg[397]) );
  DFF \creg_reg[398]  ( .D(o[398]), .CLK(clk), .RST(rst), .I(g_init[398]), .Q(
        creg[398]) );
  DFF \creg_reg[399]  ( .D(o[399]), .CLK(clk), .RST(rst), .I(g_init[399]), .Q(
        creg[399]) );
  DFF \creg_reg[400]  ( .D(o[400]), .CLK(clk), .RST(rst), .I(g_init[400]), .Q(
        creg[400]) );
  DFF \creg_reg[401]  ( .D(o[401]), .CLK(clk), .RST(rst), .I(g_init[401]), .Q(
        creg[401]) );
  DFF \creg_reg[402]  ( .D(o[402]), .CLK(clk), .RST(rst), .I(g_init[402]), .Q(
        creg[402]) );
  DFF \creg_reg[403]  ( .D(o[403]), .CLK(clk), .RST(rst), .I(g_init[403]), .Q(
        creg[403]) );
  DFF \creg_reg[404]  ( .D(o[404]), .CLK(clk), .RST(rst), .I(g_init[404]), .Q(
        creg[404]) );
  DFF \creg_reg[405]  ( .D(o[405]), .CLK(clk), .RST(rst), .I(g_init[405]), .Q(
        creg[405]) );
  DFF \creg_reg[406]  ( .D(o[406]), .CLK(clk), .RST(rst), .I(g_init[406]), .Q(
        creg[406]) );
  DFF \creg_reg[407]  ( .D(o[407]), .CLK(clk), .RST(rst), .I(g_init[407]), .Q(
        creg[407]) );
  DFF \creg_reg[408]  ( .D(o[408]), .CLK(clk), .RST(rst), .I(g_init[408]), .Q(
        creg[408]) );
  DFF \creg_reg[409]  ( .D(o[409]), .CLK(clk), .RST(rst), .I(g_init[409]), .Q(
        creg[409]) );
  DFF \creg_reg[410]  ( .D(o[410]), .CLK(clk), .RST(rst), .I(g_init[410]), .Q(
        creg[410]) );
  DFF \creg_reg[411]  ( .D(o[411]), .CLK(clk), .RST(rst), .I(g_init[411]), .Q(
        creg[411]) );
  DFF \creg_reg[412]  ( .D(o[412]), .CLK(clk), .RST(rst), .I(g_init[412]), .Q(
        creg[412]) );
  DFF \creg_reg[413]  ( .D(o[413]), .CLK(clk), .RST(rst), .I(g_init[413]), .Q(
        creg[413]) );
  DFF \creg_reg[414]  ( .D(o[414]), .CLK(clk), .RST(rst), .I(g_init[414]), .Q(
        creg[414]) );
  DFF \creg_reg[415]  ( .D(o[415]), .CLK(clk), .RST(rst), .I(g_init[415]), .Q(
        creg[415]) );
  DFF \creg_reg[416]  ( .D(o[416]), .CLK(clk), .RST(rst), .I(g_init[416]), .Q(
        creg[416]) );
  DFF \creg_reg[417]  ( .D(o[417]), .CLK(clk), .RST(rst), .I(g_init[417]), .Q(
        creg[417]) );
  DFF \creg_reg[418]  ( .D(o[418]), .CLK(clk), .RST(rst), .I(g_init[418]), .Q(
        creg[418]) );
  DFF \creg_reg[419]  ( .D(o[419]), .CLK(clk), .RST(rst), .I(g_init[419]), .Q(
        creg[419]) );
  DFF \creg_reg[420]  ( .D(o[420]), .CLK(clk), .RST(rst), .I(g_init[420]), .Q(
        creg[420]) );
  DFF \creg_reg[421]  ( .D(o[421]), .CLK(clk), .RST(rst), .I(g_init[421]), .Q(
        creg[421]) );
  DFF \creg_reg[422]  ( .D(o[422]), .CLK(clk), .RST(rst), .I(g_init[422]), .Q(
        creg[422]) );
  DFF \creg_reg[423]  ( .D(o[423]), .CLK(clk), .RST(rst), .I(g_init[423]), .Q(
        creg[423]) );
  DFF \creg_reg[424]  ( .D(o[424]), .CLK(clk), .RST(rst), .I(g_init[424]), .Q(
        creg[424]) );
  DFF \creg_reg[425]  ( .D(o[425]), .CLK(clk), .RST(rst), .I(g_init[425]), .Q(
        creg[425]) );
  DFF \creg_reg[426]  ( .D(o[426]), .CLK(clk), .RST(rst), .I(g_init[426]), .Q(
        creg[426]) );
  DFF \creg_reg[427]  ( .D(o[427]), .CLK(clk), .RST(rst), .I(g_init[427]), .Q(
        creg[427]) );
  DFF \creg_reg[428]  ( .D(o[428]), .CLK(clk), .RST(rst), .I(g_init[428]), .Q(
        creg[428]) );
  DFF \creg_reg[429]  ( .D(o[429]), .CLK(clk), .RST(rst), .I(g_init[429]), .Q(
        creg[429]) );
  DFF \creg_reg[430]  ( .D(o[430]), .CLK(clk), .RST(rst), .I(g_init[430]), .Q(
        creg[430]) );
  DFF \creg_reg[431]  ( .D(o[431]), .CLK(clk), .RST(rst), .I(g_init[431]), .Q(
        creg[431]) );
  DFF \creg_reg[432]  ( .D(o[432]), .CLK(clk), .RST(rst), .I(g_init[432]), .Q(
        creg[432]) );
  DFF \creg_reg[433]  ( .D(o[433]), .CLK(clk), .RST(rst), .I(g_init[433]), .Q(
        creg[433]) );
  DFF \creg_reg[434]  ( .D(o[434]), .CLK(clk), .RST(rst), .I(g_init[434]), .Q(
        creg[434]) );
  DFF \creg_reg[435]  ( .D(o[435]), .CLK(clk), .RST(rst), .I(g_init[435]), .Q(
        creg[435]) );
  DFF \creg_reg[436]  ( .D(o[436]), .CLK(clk), .RST(rst), .I(g_init[436]), .Q(
        creg[436]) );
  DFF \creg_reg[437]  ( .D(o[437]), .CLK(clk), .RST(rst), .I(g_init[437]), .Q(
        creg[437]) );
  DFF \creg_reg[438]  ( .D(o[438]), .CLK(clk), .RST(rst), .I(g_init[438]), .Q(
        creg[438]) );
  DFF \creg_reg[439]  ( .D(o[439]), .CLK(clk), .RST(rst), .I(g_init[439]), .Q(
        creg[439]) );
  DFF \creg_reg[440]  ( .D(o[440]), .CLK(clk), .RST(rst), .I(g_init[440]), .Q(
        creg[440]) );
  DFF \creg_reg[441]  ( .D(o[441]), .CLK(clk), .RST(rst), .I(g_init[441]), .Q(
        creg[441]) );
  DFF \creg_reg[442]  ( .D(o[442]), .CLK(clk), .RST(rst), .I(g_init[442]), .Q(
        creg[442]) );
  DFF \creg_reg[443]  ( .D(o[443]), .CLK(clk), .RST(rst), .I(g_init[443]), .Q(
        creg[443]) );
  DFF \creg_reg[444]  ( .D(o[444]), .CLK(clk), .RST(rst), .I(g_init[444]), .Q(
        creg[444]) );
  DFF \creg_reg[445]  ( .D(o[445]), .CLK(clk), .RST(rst), .I(g_init[445]), .Q(
        creg[445]) );
  DFF \creg_reg[446]  ( .D(o[446]), .CLK(clk), .RST(rst), .I(g_init[446]), .Q(
        creg[446]) );
  DFF \creg_reg[447]  ( .D(o[447]), .CLK(clk), .RST(rst), .I(g_init[447]), .Q(
        creg[447]) );
  DFF \creg_reg[448]  ( .D(o[448]), .CLK(clk), .RST(rst), .I(g_init[448]), .Q(
        creg[448]) );
  DFF \creg_reg[449]  ( .D(o[449]), .CLK(clk), .RST(rst), .I(g_init[449]), .Q(
        creg[449]) );
  DFF \creg_reg[450]  ( .D(o[450]), .CLK(clk), .RST(rst), .I(g_init[450]), .Q(
        creg[450]) );
  DFF \creg_reg[451]  ( .D(o[451]), .CLK(clk), .RST(rst), .I(g_init[451]), .Q(
        creg[451]) );
  DFF \creg_reg[452]  ( .D(o[452]), .CLK(clk), .RST(rst), .I(g_init[452]), .Q(
        creg[452]) );
  DFF \creg_reg[453]  ( .D(o[453]), .CLK(clk), .RST(rst), .I(g_init[453]), .Q(
        creg[453]) );
  DFF \creg_reg[454]  ( .D(o[454]), .CLK(clk), .RST(rst), .I(g_init[454]), .Q(
        creg[454]) );
  DFF \creg_reg[455]  ( .D(o[455]), .CLK(clk), .RST(rst), .I(g_init[455]), .Q(
        creg[455]) );
  DFF \creg_reg[456]  ( .D(o[456]), .CLK(clk), .RST(rst), .I(g_init[456]), .Q(
        creg[456]) );
  DFF \creg_reg[457]  ( .D(o[457]), .CLK(clk), .RST(rst), .I(g_init[457]), .Q(
        creg[457]) );
  DFF \creg_reg[458]  ( .D(o[458]), .CLK(clk), .RST(rst), .I(g_init[458]), .Q(
        creg[458]) );
  DFF \creg_reg[459]  ( .D(o[459]), .CLK(clk), .RST(rst), .I(g_init[459]), .Q(
        creg[459]) );
  DFF \creg_reg[460]  ( .D(o[460]), .CLK(clk), .RST(rst), .I(g_init[460]), .Q(
        creg[460]) );
  DFF \creg_reg[461]  ( .D(o[461]), .CLK(clk), .RST(rst), .I(g_init[461]), .Q(
        creg[461]) );
  DFF \creg_reg[462]  ( .D(o[462]), .CLK(clk), .RST(rst), .I(g_init[462]), .Q(
        creg[462]) );
  DFF \creg_reg[463]  ( .D(o[463]), .CLK(clk), .RST(rst), .I(g_init[463]), .Q(
        creg[463]) );
  DFF \creg_reg[464]  ( .D(o[464]), .CLK(clk), .RST(rst), .I(g_init[464]), .Q(
        creg[464]) );
  DFF \creg_reg[465]  ( .D(o[465]), .CLK(clk), .RST(rst), .I(g_init[465]), .Q(
        creg[465]) );
  DFF \creg_reg[466]  ( .D(o[466]), .CLK(clk), .RST(rst), .I(g_init[466]), .Q(
        creg[466]) );
  DFF \creg_reg[467]  ( .D(o[467]), .CLK(clk), .RST(rst), .I(g_init[467]), .Q(
        creg[467]) );
  DFF \creg_reg[468]  ( .D(o[468]), .CLK(clk), .RST(rst), .I(g_init[468]), .Q(
        creg[468]) );
  DFF \creg_reg[469]  ( .D(o[469]), .CLK(clk), .RST(rst), .I(g_init[469]), .Q(
        creg[469]) );
  DFF \creg_reg[470]  ( .D(o[470]), .CLK(clk), .RST(rst), .I(g_init[470]), .Q(
        creg[470]) );
  DFF \creg_reg[471]  ( .D(o[471]), .CLK(clk), .RST(rst), .I(g_init[471]), .Q(
        creg[471]) );
  DFF \creg_reg[472]  ( .D(o[472]), .CLK(clk), .RST(rst), .I(g_init[472]), .Q(
        creg[472]) );
  DFF \creg_reg[473]  ( .D(o[473]), .CLK(clk), .RST(rst), .I(g_init[473]), .Q(
        creg[473]) );
  DFF \creg_reg[474]  ( .D(o[474]), .CLK(clk), .RST(rst), .I(g_init[474]), .Q(
        creg[474]) );
  DFF \creg_reg[475]  ( .D(o[475]), .CLK(clk), .RST(rst), .I(g_init[475]), .Q(
        creg[475]) );
  DFF \creg_reg[476]  ( .D(o[476]), .CLK(clk), .RST(rst), .I(g_init[476]), .Q(
        creg[476]) );
  DFF \creg_reg[477]  ( .D(o[477]), .CLK(clk), .RST(rst), .I(g_init[477]), .Q(
        creg[477]) );
  DFF \creg_reg[478]  ( .D(o[478]), .CLK(clk), .RST(rst), .I(g_init[478]), .Q(
        creg[478]) );
  DFF \creg_reg[479]  ( .D(o[479]), .CLK(clk), .RST(rst), .I(g_init[479]), .Q(
        creg[479]) );
  DFF \creg_reg[480]  ( .D(o[480]), .CLK(clk), .RST(rst), .I(g_init[480]), .Q(
        creg[480]) );
  DFF \creg_reg[481]  ( .D(o[481]), .CLK(clk), .RST(rst), .I(g_init[481]), .Q(
        creg[481]) );
  DFF \creg_reg[482]  ( .D(o[482]), .CLK(clk), .RST(rst), .I(g_init[482]), .Q(
        creg[482]) );
  DFF \creg_reg[483]  ( .D(o[483]), .CLK(clk), .RST(rst), .I(g_init[483]), .Q(
        creg[483]) );
  DFF \creg_reg[484]  ( .D(o[484]), .CLK(clk), .RST(rst), .I(g_init[484]), .Q(
        creg[484]) );
  DFF \creg_reg[485]  ( .D(o[485]), .CLK(clk), .RST(rst), .I(g_init[485]), .Q(
        creg[485]) );
  DFF \creg_reg[486]  ( .D(o[486]), .CLK(clk), .RST(rst), .I(g_init[486]), .Q(
        creg[486]) );
  DFF \creg_reg[487]  ( .D(o[487]), .CLK(clk), .RST(rst), .I(g_init[487]), .Q(
        creg[487]) );
  DFF \creg_reg[488]  ( .D(o[488]), .CLK(clk), .RST(rst), .I(g_init[488]), .Q(
        creg[488]) );
  DFF \creg_reg[489]  ( .D(o[489]), .CLK(clk), .RST(rst), .I(g_init[489]), .Q(
        creg[489]) );
  DFF \creg_reg[490]  ( .D(o[490]), .CLK(clk), .RST(rst), .I(g_init[490]), .Q(
        creg[490]) );
  DFF \creg_reg[491]  ( .D(o[491]), .CLK(clk), .RST(rst), .I(g_init[491]), .Q(
        creg[491]) );
  DFF \creg_reg[492]  ( .D(o[492]), .CLK(clk), .RST(rst), .I(g_init[492]), .Q(
        creg[492]) );
  DFF \creg_reg[493]  ( .D(o[493]), .CLK(clk), .RST(rst), .I(g_init[493]), .Q(
        creg[493]) );
  DFF \creg_reg[494]  ( .D(o[494]), .CLK(clk), .RST(rst), .I(g_init[494]), .Q(
        creg[494]) );
  DFF \creg_reg[495]  ( .D(o[495]), .CLK(clk), .RST(rst), .I(g_init[495]), .Q(
        creg[495]) );
  DFF \creg_reg[496]  ( .D(o[496]), .CLK(clk), .RST(rst), .I(g_init[496]), .Q(
        creg[496]) );
  DFF \creg_reg[497]  ( .D(o[497]), .CLK(clk), .RST(rst), .I(g_init[497]), .Q(
        creg[497]) );
  DFF \creg_reg[498]  ( .D(o[498]), .CLK(clk), .RST(rst), .I(g_init[498]), .Q(
        creg[498]) );
  DFF \creg_reg[499]  ( .D(o[499]), .CLK(clk), .RST(rst), .I(g_init[499]), .Q(
        creg[499]) );
  DFF \creg_reg[500]  ( .D(o[500]), .CLK(clk), .RST(rst), .I(g_init[500]), .Q(
        creg[500]) );
  DFF \creg_reg[501]  ( .D(o[501]), .CLK(clk), .RST(rst), .I(g_init[501]), .Q(
        creg[501]) );
  DFF \creg_reg[502]  ( .D(o[502]), .CLK(clk), .RST(rst), .I(g_init[502]), .Q(
        creg[502]) );
  DFF \creg_reg[503]  ( .D(o[503]), .CLK(clk), .RST(rst), .I(g_init[503]), .Q(
        creg[503]) );
  DFF \creg_reg[504]  ( .D(o[504]), .CLK(clk), .RST(rst), .I(g_init[504]), .Q(
        creg[504]) );
  DFF \creg_reg[505]  ( .D(o[505]), .CLK(clk), .RST(rst), .I(g_init[505]), .Q(
        creg[505]) );
  DFF \creg_reg[506]  ( .D(o[506]), .CLK(clk), .RST(rst), .I(g_init[506]), .Q(
        creg[506]) );
  DFF \creg_reg[507]  ( .D(o[507]), .CLK(clk), .RST(rst), .I(g_init[507]), .Q(
        creg[507]) );
  DFF \creg_reg[508]  ( .D(o[508]), .CLK(clk), .RST(rst), .I(g_init[508]), .Q(
        creg[508]) );
  DFF \creg_reg[509]  ( .D(o[509]), .CLK(clk), .RST(rst), .I(g_init[509]), .Q(
        creg[509]) );
  DFF \creg_reg[510]  ( .D(o[510]), .CLK(clk), .RST(rst), .I(g_init[510]), .Q(
        creg[510]) );
  DFF \creg_reg[511]  ( .D(o[511]), .CLK(clk), .RST(rst), .I(g_init[511]), .Q(
        creg[511]) );
  DFF \creg_reg[512]  ( .D(o[512]), .CLK(clk), .RST(rst), .I(g_init[512]), .Q(
        creg[512]) );
  DFF \creg_reg[513]  ( .D(o[513]), .CLK(clk), .RST(rst), .I(g_init[513]), .Q(
        creg[513]) );
  DFF \creg_reg[514]  ( .D(o[514]), .CLK(clk), .RST(rst), .I(g_init[514]), .Q(
        creg[514]) );
  DFF \creg_reg[515]  ( .D(o[515]), .CLK(clk), .RST(rst), .I(g_init[515]), .Q(
        creg[515]) );
  DFF \creg_reg[516]  ( .D(o[516]), .CLK(clk), .RST(rst), .I(g_init[516]), .Q(
        creg[516]) );
  DFF \creg_reg[517]  ( .D(o[517]), .CLK(clk), .RST(rst), .I(g_init[517]), .Q(
        creg[517]) );
  DFF \creg_reg[518]  ( .D(o[518]), .CLK(clk), .RST(rst), .I(g_init[518]), .Q(
        creg[518]) );
  DFF \creg_reg[519]  ( .D(o[519]), .CLK(clk), .RST(rst), .I(g_init[519]), .Q(
        creg[519]) );
  DFF \creg_reg[520]  ( .D(o[520]), .CLK(clk), .RST(rst), .I(g_init[520]), .Q(
        creg[520]) );
  DFF \creg_reg[521]  ( .D(o[521]), .CLK(clk), .RST(rst), .I(g_init[521]), .Q(
        creg[521]) );
  DFF \creg_reg[522]  ( .D(o[522]), .CLK(clk), .RST(rst), .I(g_init[522]), .Q(
        creg[522]) );
  DFF \creg_reg[523]  ( .D(o[523]), .CLK(clk), .RST(rst), .I(g_init[523]), .Q(
        creg[523]) );
  DFF \creg_reg[524]  ( .D(o[524]), .CLK(clk), .RST(rst), .I(g_init[524]), .Q(
        creg[524]) );
  DFF \creg_reg[525]  ( .D(o[525]), .CLK(clk), .RST(rst), .I(g_init[525]), .Q(
        creg[525]) );
  DFF \creg_reg[526]  ( .D(o[526]), .CLK(clk), .RST(rst), .I(g_init[526]), .Q(
        creg[526]) );
  DFF \creg_reg[527]  ( .D(o[527]), .CLK(clk), .RST(rst), .I(g_init[527]), .Q(
        creg[527]) );
  DFF \creg_reg[528]  ( .D(o[528]), .CLK(clk), .RST(rst), .I(g_init[528]), .Q(
        creg[528]) );
  DFF \creg_reg[529]  ( .D(o[529]), .CLK(clk), .RST(rst), .I(g_init[529]), .Q(
        creg[529]) );
  DFF \creg_reg[530]  ( .D(o[530]), .CLK(clk), .RST(rst), .I(g_init[530]), .Q(
        creg[530]) );
  DFF \creg_reg[531]  ( .D(o[531]), .CLK(clk), .RST(rst), .I(g_init[531]), .Q(
        creg[531]) );
  DFF \creg_reg[532]  ( .D(o[532]), .CLK(clk), .RST(rst), .I(g_init[532]), .Q(
        creg[532]) );
  DFF \creg_reg[533]  ( .D(o[533]), .CLK(clk), .RST(rst), .I(g_init[533]), .Q(
        creg[533]) );
  DFF \creg_reg[534]  ( .D(o[534]), .CLK(clk), .RST(rst), .I(g_init[534]), .Q(
        creg[534]) );
  DFF \creg_reg[535]  ( .D(o[535]), .CLK(clk), .RST(rst), .I(g_init[535]), .Q(
        creg[535]) );
  DFF \creg_reg[536]  ( .D(o[536]), .CLK(clk), .RST(rst), .I(g_init[536]), .Q(
        creg[536]) );
  DFF \creg_reg[537]  ( .D(o[537]), .CLK(clk), .RST(rst), .I(g_init[537]), .Q(
        creg[537]) );
  DFF \creg_reg[538]  ( .D(o[538]), .CLK(clk), .RST(rst), .I(g_init[538]), .Q(
        creg[538]) );
  DFF \creg_reg[539]  ( .D(o[539]), .CLK(clk), .RST(rst), .I(g_init[539]), .Q(
        creg[539]) );
  DFF \creg_reg[540]  ( .D(o[540]), .CLK(clk), .RST(rst), .I(g_init[540]), .Q(
        creg[540]) );
  DFF \creg_reg[541]  ( .D(o[541]), .CLK(clk), .RST(rst), .I(g_init[541]), .Q(
        creg[541]) );
  DFF \creg_reg[542]  ( .D(o[542]), .CLK(clk), .RST(rst), .I(g_init[542]), .Q(
        creg[542]) );
  DFF \creg_reg[543]  ( .D(o[543]), .CLK(clk), .RST(rst), .I(g_init[543]), .Q(
        creg[543]) );
  DFF \creg_reg[544]  ( .D(o[544]), .CLK(clk), .RST(rst), .I(g_init[544]), .Q(
        creg[544]) );
  DFF \creg_reg[545]  ( .D(o[545]), .CLK(clk), .RST(rst), .I(g_init[545]), .Q(
        creg[545]) );
  DFF \creg_reg[546]  ( .D(o[546]), .CLK(clk), .RST(rst), .I(g_init[546]), .Q(
        creg[546]) );
  DFF \creg_reg[547]  ( .D(o[547]), .CLK(clk), .RST(rst), .I(g_init[547]), .Q(
        creg[547]) );
  DFF \creg_reg[548]  ( .D(o[548]), .CLK(clk), .RST(rst), .I(g_init[548]), .Q(
        creg[548]) );
  DFF \creg_reg[549]  ( .D(o[549]), .CLK(clk), .RST(rst), .I(g_init[549]), .Q(
        creg[549]) );
  DFF \creg_reg[550]  ( .D(o[550]), .CLK(clk), .RST(rst), .I(g_init[550]), .Q(
        creg[550]) );
  DFF \creg_reg[551]  ( .D(o[551]), .CLK(clk), .RST(rst), .I(g_init[551]), .Q(
        creg[551]) );
  DFF \creg_reg[552]  ( .D(o[552]), .CLK(clk), .RST(rst), .I(g_init[552]), .Q(
        creg[552]) );
  DFF \creg_reg[553]  ( .D(o[553]), .CLK(clk), .RST(rst), .I(g_init[553]), .Q(
        creg[553]) );
  DFF \creg_reg[554]  ( .D(o[554]), .CLK(clk), .RST(rst), .I(g_init[554]), .Q(
        creg[554]) );
  DFF \creg_reg[555]  ( .D(o[555]), .CLK(clk), .RST(rst), .I(g_init[555]), .Q(
        creg[555]) );
  DFF \creg_reg[556]  ( .D(o[556]), .CLK(clk), .RST(rst), .I(g_init[556]), .Q(
        creg[556]) );
  DFF \creg_reg[557]  ( .D(o[557]), .CLK(clk), .RST(rst), .I(g_init[557]), .Q(
        creg[557]) );
  DFF \creg_reg[558]  ( .D(o[558]), .CLK(clk), .RST(rst), .I(g_init[558]), .Q(
        creg[558]) );
  DFF \creg_reg[559]  ( .D(o[559]), .CLK(clk), .RST(rst), .I(g_init[559]), .Q(
        creg[559]) );
  DFF \creg_reg[560]  ( .D(o[560]), .CLK(clk), .RST(rst), .I(g_init[560]), .Q(
        creg[560]) );
  DFF \creg_reg[561]  ( .D(o[561]), .CLK(clk), .RST(rst), .I(g_init[561]), .Q(
        creg[561]) );
  DFF \creg_reg[562]  ( .D(o[562]), .CLK(clk), .RST(rst), .I(g_init[562]), .Q(
        creg[562]) );
  DFF \creg_reg[563]  ( .D(o[563]), .CLK(clk), .RST(rst), .I(g_init[563]), .Q(
        creg[563]) );
  DFF \creg_reg[564]  ( .D(o[564]), .CLK(clk), .RST(rst), .I(g_init[564]), .Q(
        creg[564]) );
  DFF \creg_reg[565]  ( .D(o[565]), .CLK(clk), .RST(rst), .I(g_init[565]), .Q(
        creg[565]) );
  DFF \creg_reg[566]  ( .D(o[566]), .CLK(clk), .RST(rst), .I(g_init[566]), .Q(
        creg[566]) );
  DFF \creg_reg[567]  ( .D(o[567]), .CLK(clk), .RST(rst), .I(g_init[567]), .Q(
        creg[567]) );
  DFF \creg_reg[568]  ( .D(o[568]), .CLK(clk), .RST(rst), .I(g_init[568]), .Q(
        creg[568]) );
  DFF \creg_reg[569]  ( .D(o[569]), .CLK(clk), .RST(rst), .I(g_init[569]), .Q(
        creg[569]) );
  DFF \creg_reg[570]  ( .D(o[570]), .CLK(clk), .RST(rst), .I(g_init[570]), .Q(
        creg[570]) );
  DFF \creg_reg[571]  ( .D(o[571]), .CLK(clk), .RST(rst), .I(g_init[571]), .Q(
        creg[571]) );
  DFF \creg_reg[572]  ( .D(o[572]), .CLK(clk), .RST(rst), .I(g_init[572]), .Q(
        creg[572]) );
  DFF \creg_reg[573]  ( .D(o[573]), .CLK(clk), .RST(rst), .I(g_init[573]), .Q(
        creg[573]) );
  DFF \creg_reg[574]  ( .D(o[574]), .CLK(clk), .RST(rst), .I(g_init[574]), .Q(
        creg[574]) );
  DFF \creg_reg[575]  ( .D(o[575]), .CLK(clk), .RST(rst), .I(g_init[575]), .Q(
        creg[575]) );
  DFF \creg_reg[576]  ( .D(o[576]), .CLK(clk), .RST(rst), .I(g_init[576]), .Q(
        creg[576]) );
  DFF \creg_reg[577]  ( .D(o[577]), .CLK(clk), .RST(rst), .I(g_init[577]), .Q(
        creg[577]) );
  DFF \creg_reg[578]  ( .D(o[578]), .CLK(clk), .RST(rst), .I(g_init[578]), .Q(
        creg[578]) );
  DFF \creg_reg[579]  ( .D(o[579]), .CLK(clk), .RST(rst), .I(g_init[579]), .Q(
        creg[579]) );
  DFF \creg_reg[580]  ( .D(o[580]), .CLK(clk), .RST(rst), .I(g_init[580]), .Q(
        creg[580]) );
  DFF \creg_reg[581]  ( .D(o[581]), .CLK(clk), .RST(rst), .I(g_init[581]), .Q(
        creg[581]) );
  DFF \creg_reg[582]  ( .D(o[582]), .CLK(clk), .RST(rst), .I(g_init[582]), .Q(
        creg[582]) );
  DFF \creg_reg[583]  ( .D(o[583]), .CLK(clk), .RST(rst), .I(g_init[583]), .Q(
        creg[583]) );
  DFF \creg_reg[584]  ( .D(o[584]), .CLK(clk), .RST(rst), .I(g_init[584]), .Q(
        creg[584]) );
  DFF \creg_reg[585]  ( .D(o[585]), .CLK(clk), .RST(rst), .I(g_init[585]), .Q(
        creg[585]) );
  DFF \creg_reg[586]  ( .D(o[586]), .CLK(clk), .RST(rst), .I(g_init[586]), .Q(
        creg[586]) );
  DFF \creg_reg[587]  ( .D(o[587]), .CLK(clk), .RST(rst), .I(g_init[587]), .Q(
        creg[587]) );
  DFF \creg_reg[588]  ( .D(o[588]), .CLK(clk), .RST(rst), .I(g_init[588]), .Q(
        creg[588]) );
  DFF \creg_reg[589]  ( .D(o[589]), .CLK(clk), .RST(rst), .I(g_init[589]), .Q(
        creg[589]) );
  DFF \creg_reg[590]  ( .D(o[590]), .CLK(clk), .RST(rst), .I(g_init[590]), .Q(
        creg[590]) );
  DFF \creg_reg[591]  ( .D(o[591]), .CLK(clk), .RST(rst), .I(g_init[591]), .Q(
        creg[591]) );
  DFF \creg_reg[592]  ( .D(o[592]), .CLK(clk), .RST(rst), .I(g_init[592]), .Q(
        creg[592]) );
  DFF \creg_reg[593]  ( .D(o[593]), .CLK(clk), .RST(rst), .I(g_init[593]), .Q(
        creg[593]) );
  DFF \creg_reg[594]  ( .D(o[594]), .CLK(clk), .RST(rst), .I(g_init[594]), .Q(
        creg[594]) );
  DFF \creg_reg[595]  ( .D(o[595]), .CLK(clk), .RST(rst), .I(g_init[595]), .Q(
        creg[595]) );
  DFF \creg_reg[596]  ( .D(o[596]), .CLK(clk), .RST(rst), .I(g_init[596]), .Q(
        creg[596]) );
  DFF \creg_reg[597]  ( .D(o[597]), .CLK(clk), .RST(rst), .I(g_init[597]), .Q(
        creg[597]) );
  DFF \creg_reg[598]  ( .D(o[598]), .CLK(clk), .RST(rst), .I(g_init[598]), .Q(
        creg[598]) );
  DFF \creg_reg[599]  ( .D(o[599]), .CLK(clk), .RST(rst), .I(g_init[599]), .Q(
        creg[599]) );
  DFF \creg_reg[600]  ( .D(o[600]), .CLK(clk), .RST(rst), .I(g_init[600]), .Q(
        creg[600]) );
  DFF \creg_reg[601]  ( .D(o[601]), .CLK(clk), .RST(rst), .I(g_init[601]), .Q(
        creg[601]) );
  DFF \creg_reg[602]  ( .D(o[602]), .CLK(clk), .RST(rst), .I(g_init[602]), .Q(
        creg[602]) );
  DFF \creg_reg[603]  ( .D(o[603]), .CLK(clk), .RST(rst), .I(g_init[603]), .Q(
        creg[603]) );
  DFF \creg_reg[604]  ( .D(o[604]), .CLK(clk), .RST(rst), .I(g_init[604]), .Q(
        creg[604]) );
  DFF \creg_reg[605]  ( .D(o[605]), .CLK(clk), .RST(rst), .I(g_init[605]), .Q(
        creg[605]) );
  DFF \creg_reg[606]  ( .D(o[606]), .CLK(clk), .RST(rst), .I(g_init[606]), .Q(
        creg[606]) );
  DFF \creg_reg[607]  ( .D(o[607]), .CLK(clk), .RST(rst), .I(g_init[607]), .Q(
        creg[607]) );
  DFF \creg_reg[608]  ( .D(o[608]), .CLK(clk), .RST(rst), .I(g_init[608]), .Q(
        creg[608]) );
  DFF \creg_reg[609]  ( .D(o[609]), .CLK(clk), .RST(rst), .I(g_init[609]), .Q(
        creg[609]) );
  DFF \creg_reg[610]  ( .D(o[610]), .CLK(clk), .RST(rst), .I(g_init[610]), .Q(
        creg[610]) );
  DFF \creg_reg[611]  ( .D(o[611]), .CLK(clk), .RST(rst), .I(g_init[611]), .Q(
        creg[611]) );
  DFF \creg_reg[612]  ( .D(o[612]), .CLK(clk), .RST(rst), .I(g_init[612]), .Q(
        creg[612]) );
  DFF \creg_reg[613]  ( .D(o[613]), .CLK(clk), .RST(rst), .I(g_init[613]), .Q(
        creg[613]) );
  DFF \creg_reg[614]  ( .D(o[614]), .CLK(clk), .RST(rst), .I(g_init[614]), .Q(
        creg[614]) );
  DFF \creg_reg[615]  ( .D(o[615]), .CLK(clk), .RST(rst), .I(g_init[615]), .Q(
        creg[615]) );
  DFF \creg_reg[616]  ( .D(o[616]), .CLK(clk), .RST(rst), .I(g_init[616]), .Q(
        creg[616]) );
  DFF \creg_reg[617]  ( .D(o[617]), .CLK(clk), .RST(rst), .I(g_init[617]), .Q(
        creg[617]) );
  DFF \creg_reg[618]  ( .D(o[618]), .CLK(clk), .RST(rst), .I(g_init[618]), .Q(
        creg[618]) );
  DFF \creg_reg[619]  ( .D(o[619]), .CLK(clk), .RST(rst), .I(g_init[619]), .Q(
        creg[619]) );
  DFF \creg_reg[620]  ( .D(o[620]), .CLK(clk), .RST(rst), .I(g_init[620]), .Q(
        creg[620]) );
  DFF \creg_reg[621]  ( .D(o[621]), .CLK(clk), .RST(rst), .I(g_init[621]), .Q(
        creg[621]) );
  DFF \creg_reg[622]  ( .D(o[622]), .CLK(clk), .RST(rst), .I(g_init[622]), .Q(
        creg[622]) );
  DFF \creg_reg[623]  ( .D(o[623]), .CLK(clk), .RST(rst), .I(g_init[623]), .Q(
        creg[623]) );
  DFF \creg_reg[624]  ( .D(o[624]), .CLK(clk), .RST(rst), .I(g_init[624]), .Q(
        creg[624]) );
  DFF \creg_reg[625]  ( .D(o[625]), .CLK(clk), .RST(rst), .I(g_init[625]), .Q(
        creg[625]) );
  DFF \creg_reg[626]  ( .D(o[626]), .CLK(clk), .RST(rst), .I(g_init[626]), .Q(
        creg[626]) );
  DFF \creg_reg[627]  ( .D(o[627]), .CLK(clk), .RST(rst), .I(g_init[627]), .Q(
        creg[627]) );
  DFF \creg_reg[628]  ( .D(o[628]), .CLK(clk), .RST(rst), .I(g_init[628]), .Q(
        creg[628]) );
  DFF \creg_reg[629]  ( .D(o[629]), .CLK(clk), .RST(rst), .I(g_init[629]), .Q(
        creg[629]) );
  DFF \creg_reg[630]  ( .D(o[630]), .CLK(clk), .RST(rst), .I(g_init[630]), .Q(
        creg[630]) );
  DFF \creg_reg[631]  ( .D(o[631]), .CLK(clk), .RST(rst), .I(g_init[631]), .Q(
        creg[631]) );
  DFF \creg_reg[632]  ( .D(o[632]), .CLK(clk), .RST(rst), .I(g_init[632]), .Q(
        creg[632]) );
  DFF \creg_reg[633]  ( .D(o[633]), .CLK(clk), .RST(rst), .I(g_init[633]), .Q(
        creg[633]) );
  DFF \creg_reg[634]  ( .D(o[634]), .CLK(clk), .RST(rst), .I(g_init[634]), .Q(
        creg[634]) );
  DFF \creg_reg[635]  ( .D(o[635]), .CLK(clk), .RST(rst), .I(g_init[635]), .Q(
        creg[635]) );
  DFF \creg_reg[636]  ( .D(o[636]), .CLK(clk), .RST(rst), .I(g_init[636]), .Q(
        creg[636]) );
  DFF \creg_reg[637]  ( .D(o[637]), .CLK(clk), .RST(rst), .I(g_init[637]), .Q(
        creg[637]) );
  DFF \creg_reg[638]  ( .D(o[638]), .CLK(clk), .RST(rst), .I(g_init[638]), .Q(
        creg[638]) );
  DFF \creg_reg[639]  ( .D(o[639]), .CLK(clk), .RST(rst), .I(g_init[639]), .Q(
        creg[639]) );
  DFF \creg_reg[640]  ( .D(o[640]), .CLK(clk), .RST(rst), .I(g_init[640]), .Q(
        creg[640]) );
  DFF \creg_reg[641]  ( .D(o[641]), .CLK(clk), .RST(rst), .I(g_init[641]), .Q(
        creg[641]) );
  DFF \creg_reg[642]  ( .D(o[642]), .CLK(clk), .RST(rst), .I(g_init[642]), .Q(
        creg[642]) );
  DFF \creg_reg[643]  ( .D(o[643]), .CLK(clk), .RST(rst), .I(g_init[643]), .Q(
        creg[643]) );
  DFF \creg_reg[644]  ( .D(o[644]), .CLK(clk), .RST(rst), .I(g_init[644]), .Q(
        creg[644]) );
  DFF \creg_reg[645]  ( .D(o[645]), .CLK(clk), .RST(rst), .I(g_init[645]), .Q(
        creg[645]) );
  DFF \creg_reg[646]  ( .D(o[646]), .CLK(clk), .RST(rst), .I(g_init[646]), .Q(
        creg[646]) );
  DFF \creg_reg[647]  ( .D(o[647]), .CLK(clk), .RST(rst), .I(g_init[647]), .Q(
        creg[647]) );
  DFF \creg_reg[648]  ( .D(o[648]), .CLK(clk), .RST(rst), .I(g_init[648]), .Q(
        creg[648]) );
  DFF \creg_reg[649]  ( .D(o[649]), .CLK(clk), .RST(rst), .I(g_init[649]), .Q(
        creg[649]) );
  DFF \creg_reg[650]  ( .D(o[650]), .CLK(clk), .RST(rst), .I(g_init[650]), .Q(
        creg[650]) );
  DFF \creg_reg[651]  ( .D(o[651]), .CLK(clk), .RST(rst), .I(g_init[651]), .Q(
        creg[651]) );
  DFF \creg_reg[652]  ( .D(o[652]), .CLK(clk), .RST(rst), .I(g_init[652]), .Q(
        creg[652]) );
  DFF \creg_reg[653]  ( .D(o[653]), .CLK(clk), .RST(rst), .I(g_init[653]), .Q(
        creg[653]) );
  DFF \creg_reg[654]  ( .D(o[654]), .CLK(clk), .RST(rst), .I(g_init[654]), .Q(
        creg[654]) );
  DFF \creg_reg[655]  ( .D(o[655]), .CLK(clk), .RST(rst), .I(g_init[655]), .Q(
        creg[655]) );
  DFF \creg_reg[656]  ( .D(o[656]), .CLK(clk), .RST(rst), .I(g_init[656]), .Q(
        creg[656]) );
  DFF \creg_reg[657]  ( .D(o[657]), .CLK(clk), .RST(rst), .I(g_init[657]), .Q(
        creg[657]) );
  DFF \creg_reg[658]  ( .D(o[658]), .CLK(clk), .RST(rst), .I(g_init[658]), .Q(
        creg[658]) );
  DFF \creg_reg[659]  ( .D(o[659]), .CLK(clk), .RST(rst), .I(g_init[659]), .Q(
        creg[659]) );
  DFF \creg_reg[660]  ( .D(o[660]), .CLK(clk), .RST(rst), .I(g_init[660]), .Q(
        creg[660]) );
  DFF \creg_reg[661]  ( .D(o[661]), .CLK(clk), .RST(rst), .I(g_init[661]), .Q(
        creg[661]) );
  DFF \creg_reg[662]  ( .D(o[662]), .CLK(clk), .RST(rst), .I(g_init[662]), .Q(
        creg[662]) );
  DFF \creg_reg[663]  ( .D(o[663]), .CLK(clk), .RST(rst), .I(g_init[663]), .Q(
        creg[663]) );
  DFF \creg_reg[664]  ( .D(o[664]), .CLK(clk), .RST(rst), .I(g_init[664]), .Q(
        creg[664]) );
  DFF \creg_reg[665]  ( .D(o[665]), .CLK(clk), .RST(rst), .I(g_init[665]), .Q(
        creg[665]) );
  DFF \creg_reg[666]  ( .D(o[666]), .CLK(clk), .RST(rst), .I(g_init[666]), .Q(
        creg[666]) );
  DFF \creg_reg[667]  ( .D(o[667]), .CLK(clk), .RST(rst), .I(g_init[667]), .Q(
        creg[667]) );
  DFF \creg_reg[668]  ( .D(o[668]), .CLK(clk), .RST(rst), .I(g_init[668]), .Q(
        creg[668]) );
  DFF \creg_reg[669]  ( .D(o[669]), .CLK(clk), .RST(rst), .I(g_init[669]), .Q(
        creg[669]) );
  DFF \creg_reg[670]  ( .D(o[670]), .CLK(clk), .RST(rst), .I(g_init[670]), .Q(
        creg[670]) );
  DFF \creg_reg[671]  ( .D(o[671]), .CLK(clk), .RST(rst), .I(g_init[671]), .Q(
        creg[671]) );
  DFF \creg_reg[672]  ( .D(o[672]), .CLK(clk), .RST(rst), .I(g_init[672]), .Q(
        creg[672]) );
  DFF \creg_reg[673]  ( .D(o[673]), .CLK(clk), .RST(rst), .I(g_init[673]), .Q(
        creg[673]) );
  DFF \creg_reg[674]  ( .D(o[674]), .CLK(clk), .RST(rst), .I(g_init[674]), .Q(
        creg[674]) );
  DFF \creg_reg[675]  ( .D(o[675]), .CLK(clk), .RST(rst), .I(g_init[675]), .Q(
        creg[675]) );
  DFF \creg_reg[676]  ( .D(o[676]), .CLK(clk), .RST(rst), .I(g_init[676]), .Q(
        creg[676]) );
  DFF \creg_reg[677]  ( .D(o[677]), .CLK(clk), .RST(rst), .I(g_init[677]), .Q(
        creg[677]) );
  DFF \creg_reg[678]  ( .D(o[678]), .CLK(clk), .RST(rst), .I(g_init[678]), .Q(
        creg[678]) );
  DFF \creg_reg[679]  ( .D(o[679]), .CLK(clk), .RST(rst), .I(g_init[679]), .Q(
        creg[679]) );
  DFF \creg_reg[680]  ( .D(o[680]), .CLK(clk), .RST(rst), .I(g_init[680]), .Q(
        creg[680]) );
  DFF \creg_reg[681]  ( .D(o[681]), .CLK(clk), .RST(rst), .I(g_init[681]), .Q(
        creg[681]) );
  DFF \creg_reg[682]  ( .D(o[682]), .CLK(clk), .RST(rst), .I(g_init[682]), .Q(
        creg[682]) );
  DFF \creg_reg[683]  ( .D(o[683]), .CLK(clk), .RST(rst), .I(g_init[683]), .Q(
        creg[683]) );
  DFF \creg_reg[684]  ( .D(o[684]), .CLK(clk), .RST(rst), .I(g_init[684]), .Q(
        creg[684]) );
  DFF \creg_reg[685]  ( .D(o[685]), .CLK(clk), .RST(rst), .I(g_init[685]), .Q(
        creg[685]) );
  DFF \creg_reg[686]  ( .D(o[686]), .CLK(clk), .RST(rst), .I(g_init[686]), .Q(
        creg[686]) );
  DFF \creg_reg[687]  ( .D(o[687]), .CLK(clk), .RST(rst), .I(g_init[687]), .Q(
        creg[687]) );
  DFF \creg_reg[688]  ( .D(o[688]), .CLK(clk), .RST(rst), .I(g_init[688]), .Q(
        creg[688]) );
  DFF \creg_reg[689]  ( .D(o[689]), .CLK(clk), .RST(rst), .I(g_init[689]), .Q(
        creg[689]) );
  DFF \creg_reg[690]  ( .D(o[690]), .CLK(clk), .RST(rst), .I(g_init[690]), .Q(
        creg[690]) );
  DFF \creg_reg[691]  ( .D(o[691]), .CLK(clk), .RST(rst), .I(g_init[691]), .Q(
        creg[691]) );
  DFF \creg_reg[692]  ( .D(o[692]), .CLK(clk), .RST(rst), .I(g_init[692]), .Q(
        creg[692]) );
  DFF \creg_reg[693]  ( .D(o[693]), .CLK(clk), .RST(rst), .I(g_init[693]), .Q(
        creg[693]) );
  DFF \creg_reg[694]  ( .D(o[694]), .CLK(clk), .RST(rst), .I(g_init[694]), .Q(
        creg[694]) );
  DFF \creg_reg[695]  ( .D(o[695]), .CLK(clk), .RST(rst), .I(g_init[695]), .Q(
        creg[695]) );
  DFF \creg_reg[696]  ( .D(o[696]), .CLK(clk), .RST(rst), .I(g_init[696]), .Q(
        creg[696]) );
  DFF \creg_reg[697]  ( .D(o[697]), .CLK(clk), .RST(rst), .I(g_init[697]), .Q(
        creg[697]) );
  DFF \creg_reg[698]  ( .D(o[698]), .CLK(clk), .RST(rst), .I(g_init[698]), .Q(
        creg[698]) );
  DFF \creg_reg[699]  ( .D(o[699]), .CLK(clk), .RST(rst), .I(g_init[699]), .Q(
        creg[699]) );
  DFF \creg_reg[700]  ( .D(o[700]), .CLK(clk), .RST(rst), .I(g_init[700]), .Q(
        creg[700]) );
  DFF \creg_reg[701]  ( .D(o[701]), .CLK(clk), .RST(rst), .I(g_init[701]), .Q(
        creg[701]) );
  DFF \creg_reg[702]  ( .D(o[702]), .CLK(clk), .RST(rst), .I(g_init[702]), .Q(
        creg[702]) );
  DFF \creg_reg[703]  ( .D(o[703]), .CLK(clk), .RST(rst), .I(g_init[703]), .Q(
        creg[703]) );
  DFF \creg_reg[704]  ( .D(o[704]), .CLK(clk), .RST(rst), .I(g_init[704]), .Q(
        creg[704]) );
  DFF \creg_reg[705]  ( .D(o[705]), .CLK(clk), .RST(rst), .I(g_init[705]), .Q(
        creg[705]) );
  DFF \creg_reg[706]  ( .D(o[706]), .CLK(clk), .RST(rst), .I(g_init[706]), .Q(
        creg[706]) );
  DFF \creg_reg[707]  ( .D(o[707]), .CLK(clk), .RST(rst), .I(g_init[707]), .Q(
        creg[707]) );
  DFF \creg_reg[708]  ( .D(o[708]), .CLK(clk), .RST(rst), .I(g_init[708]), .Q(
        creg[708]) );
  DFF \creg_reg[709]  ( .D(o[709]), .CLK(clk), .RST(rst), .I(g_init[709]), .Q(
        creg[709]) );
  DFF \creg_reg[710]  ( .D(o[710]), .CLK(clk), .RST(rst), .I(g_init[710]), .Q(
        creg[710]) );
  DFF \creg_reg[711]  ( .D(o[711]), .CLK(clk), .RST(rst), .I(g_init[711]), .Q(
        creg[711]) );
  DFF \creg_reg[712]  ( .D(o[712]), .CLK(clk), .RST(rst), .I(g_init[712]), .Q(
        creg[712]) );
  DFF \creg_reg[713]  ( .D(o[713]), .CLK(clk), .RST(rst), .I(g_init[713]), .Q(
        creg[713]) );
  DFF \creg_reg[714]  ( .D(o[714]), .CLK(clk), .RST(rst), .I(g_init[714]), .Q(
        creg[714]) );
  DFF \creg_reg[715]  ( .D(o[715]), .CLK(clk), .RST(rst), .I(g_init[715]), .Q(
        creg[715]) );
  DFF \creg_reg[716]  ( .D(o[716]), .CLK(clk), .RST(rst), .I(g_init[716]), .Q(
        creg[716]) );
  DFF \creg_reg[717]  ( .D(o[717]), .CLK(clk), .RST(rst), .I(g_init[717]), .Q(
        creg[717]) );
  DFF \creg_reg[718]  ( .D(o[718]), .CLK(clk), .RST(rst), .I(g_init[718]), .Q(
        creg[718]) );
  DFF \creg_reg[719]  ( .D(o[719]), .CLK(clk), .RST(rst), .I(g_init[719]), .Q(
        creg[719]) );
  DFF \creg_reg[720]  ( .D(o[720]), .CLK(clk), .RST(rst), .I(g_init[720]), .Q(
        creg[720]) );
  DFF \creg_reg[721]  ( .D(o[721]), .CLK(clk), .RST(rst), .I(g_init[721]), .Q(
        creg[721]) );
  DFF \creg_reg[722]  ( .D(o[722]), .CLK(clk), .RST(rst), .I(g_init[722]), .Q(
        creg[722]) );
  DFF \creg_reg[723]  ( .D(o[723]), .CLK(clk), .RST(rst), .I(g_init[723]), .Q(
        creg[723]) );
  DFF \creg_reg[724]  ( .D(o[724]), .CLK(clk), .RST(rst), .I(g_init[724]), .Q(
        creg[724]) );
  DFF \creg_reg[725]  ( .D(o[725]), .CLK(clk), .RST(rst), .I(g_init[725]), .Q(
        creg[725]) );
  DFF \creg_reg[726]  ( .D(o[726]), .CLK(clk), .RST(rst), .I(g_init[726]), .Q(
        creg[726]) );
  DFF \creg_reg[727]  ( .D(o[727]), .CLK(clk), .RST(rst), .I(g_init[727]), .Q(
        creg[727]) );
  DFF \creg_reg[728]  ( .D(o[728]), .CLK(clk), .RST(rst), .I(g_init[728]), .Q(
        creg[728]) );
  DFF \creg_reg[729]  ( .D(o[729]), .CLK(clk), .RST(rst), .I(g_init[729]), .Q(
        creg[729]) );
  DFF \creg_reg[730]  ( .D(o[730]), .CLK(clk), .RST(rst), .I(g_init[730]), .Q(
        creg[730]) );
  DFF \creg_reg[731]  ( .D(o[731]), .CLK(clk), .RST(rst), .I(g_init[731]), .Q(
        creg[731]) );
  DFF \creg_reg[732]  ( .D(o[732]), .CLK(clk), .RST(rst), .I(g_init[732]), .Q(
        creg[732]) );
  DFF \creg_reg[733]  ( .D(o[733]), .CLK(clk), .RST(rst), .I(g_init[733]), .Q(
        creg[733]) );
  DFF \creg_reg[734]  ( .D(o[734]), .CLK(clk), .RST(rst), .I(g_init[734]), .Q(
        creg[734]) );
  DFF \creg_reg[735]  ( .D(o[735]), .CLK(clk), .RST(rst), .I(g_init[735]), .Q(
        creg[735]) );
  DFF \creg_reg[736]  ( .D(o[736]), .CLK(clk), .RST(rst), .I(g_init[736]), .Q(
        creg[736]) );
  DFF \creg_reg[737]  ( .D(o[737]), .CLK(clk), .RST(rst), .I(g_init[737]), .Q(
        creg[737]) );
  DFF \creg_reg[738]  ( .D(o[738]), .CLK(clk), .RST(rst), .I(g_init[738]), .Q(
        creg[738]) );
  DFF \creg_reg[739]  ( .D(o[739]), .CLK(clk), .RST(rst), .I(g_init[739]), .Q(
        creg[739]) );
  DFF \creg_reg[740]  ( .D(o[740]), .CLK(clk), .RST(rst), .I(g_init[740]), .Q(
        creg[740]) );
  DFF \creg_reg[741]  ( .D(o[741]), .CLK(clk), .RST(rst), .I(g_init[741]), .Q(
        creg[741]) );
  DFF \creg_reg[742]  ( .D(o[742]), .CLK(clk), .RST(rst), .I(g_init[742]), .Q(
        creg[742]) );
  DFF \creg_reg[743]  ( .D(o[743]), .CLK(clk), .RST(rst), .I(g_init[743]), .Q(
        creg[743]) );
  DFF \creg_reg[744]  ( .D(o[744]), .CLK(clk), .RST(rst), .I(g_init[744]), .Q(
        creg[744]) );
  DFF \creg_reg[745]  ( .D(o[745]), .CLK(clk), .RST(rst), .I(g_init[745]), .Q(
        creg[745]) );
  DFF \creg_reg[746]  ( .D(o[746]), .CLK(clk), .RST(rst), .I(g_init[746]), .Q(
        creg[746]) );
  DFF \creg_reg[747]  ( .D(o[747]), .CLK(clk), .RST(rst), .I(g_init[747]), .Q(
        creg[747]) );
  DFF \creg_reg[748]  ( .D(o[748]), .CLK(clk), .RST(rst), .I(g_init[748]), .Q(
        creg[748]) );
  DFF \creg_reg[749]  ( .D(o[749]), .CLK(clk), .RST(rst), .I(g_init[749]), .Q(
        creg[749]) );
  DFF \creg_reg[750]  ( .D(o[750]), .CLK(clk), .RST(rst), .I(g_init[750]), .Q(
        creg[750]) );
  DFF \creg_reg[751]  ( .D(o[751]), .CLK(clk), .RST(rst), .I(g_init[751]), .Q(
        creg[751]) );
  DFF \creg_reg[752]  ( .D(o[752]), .CLK(clk), .RST(rst), .I(g_init[752]), .Q(
        creg[752]) );
  DFF \creg_reg[753]  ( .D(o[753]), .CLK(clk), .RST(rst), .I(g_init[753]), .Q(
        creg[753]) );
  DFF \creg_reg[754]  ( .D(o[754]), .CLK(clk), .RST(rst), .I(g_init[754]), .Q(
        creg[754]) );
  DFF \creg_reg[755]  ( .D(o[755]), .CLK(clk), .RST(rst), .I(g_init[755]), .Q(
        creg[755]) );
  DFF \creg_reg[756]  ( .D(o[756]), .CLK(clk), .RST(rst), .I(g_init[756]), .Q(
        creg[756]) );
  DFF \creg_reg[757]  ( .D(o[757]), .CLK(clk), .RST(rst), .I(g_init[757]), .Q(
        creg[757]) );
  DFF \creg_reg[758]  ( .D(o[758]), .CLK(clk), .RST(rst), .I(g_init[758]), .Q(
        creg[758]) );
  DFF \creg_reg[759]  ( .D(o[759]), .CLK(clk), .RST(rst), .I(g_init[759]), .Q(
        creg[759]) );
  DFF \creg_reg[760]  ( .D(o[760]), .CLK(clk), .RST(rst), .I(g_init[760]), .Q(
        creg[760]) );
  DFF \creg_reg[761]  ( .D(o[761]), .CLK(clk), .RST(rst), .I(g_init[761]), .Q(
        creg[761]) );
  DFF \creg_reg[762]  ( .D(o[762]), .CLK(clk), .RST(rst), .I(g_init[762]), .Q(
        creg[762]) );
  DFF \creg_reg[763]  ( .D(o[763]), .CLK(clk), .RST(rst), .I(g_init[763]), .Q(
        creg[763]) );
  DFF \creg_reg[764]  ( .D(o[764]), .CLK(clk), .RST(rst), .I(g_init[764]), .Q(
        creg[764]) );
  DFF \creg_reg[765]  ( .D(o[765]), .CLK(clk), .RST(rst), .I(g_init[765]), .Q(
        creg[765]) );
  DFF \creg_reg[766]  ( .D(o[766]), .CLK(clk), .RST(rst), .I(g_init[766]), .Q(
        creg[766]) );
  DFF \creg_reg[767]  ( .D(o[767]), .CLK(clk), .RST(rst), .I(g_init[767]), .Q(
        creg[767]) );
  DFF \creg_reg[768]  ( .D(o[768]), .CLK(clk), .RST(rst), .I(g_init[768]), .Q(
        creg[768]) );
  DFF \creg_reg[769]  ( .D(o[769]), .CLK(clk), .RST(rst), .I(g_init[769]), .Q(
        creg[769]) );
  DFF \creg_reg[770]  ( .D(o[770]), .CLK(clk), .RST(rst), .I(g_init[770]), .Q(
        creg[770]) );
  DFF \creg_reg[771]  ( .D(o[771]), .CLK(clk), .RST(rst), .I(g_init[771]), .Q(
        creg[771]) );
  DFF \creg_reg[772]  ( .D(o[772]), .CLK(clk), .RST(rst), .I(g_init[772]), .Q(
        creg[772]) );
  DFF \creg_reg[773]  ( .D(o[773]), .CLK(clk), .RST(rst), .I(g_init[773]), .Q(
        creg[773]) );
  DFF \creg_reg[774]  ( .D(o[774]), .CLK(clk), .RST(rst), .I(g_init[774]), .Q(
        creg[774]) );
  DFF \creg_reg[775]  ( .D(o[775]), .CLK(clk), .RST(rst), .I(g_init[775]), .Q(
        creg[775]) );
  DFF \creg_reg[776]  ( .D(o[776]), .CLK(clk), .RST(rst), .I(g_init[776]), .Q(
        creg[776]) );
  DFF \creg_reg[777]  ( .D(o[777]), .CLK(clk), .RST(rst), .I(g_init[777]), .Q(
        creg[777]) );
  DFF \creg_reg[778]  ( .D(o[778]), .CLK(clk), .RST(rst), .I(g_init[778]), .Q(
        creg[778]) );
  DFF \creg_reg[779]  ( .D(o[779]), .CLK(clk), .RST(rst), .I(g_init[779]), .Q(
        creg[779]) );
  DFF \creg_reg[780]  ( .D(o[780]), .CLK(clk), .RST(rst), .I(g_init[780]), .Q(
        creg[780]) );
  DFF \creg_reg[781]  ( .D(o[781]), .CLK(clk), .RST(rst), .I(g_init[781]), .Q(
        creg[781]) );
  DFF \creg_reg[782]  ( .D(o[782]), .CLK(clk), .RST(rst), .I(g_init[782]), .Q(
        creg[782]) );
  DFF \creg_reg[783]  ( .D(o[783]), .CLK(clk), .RST(rst), .I(g_init[783]), .Q(
        creg[783]) );
  DFF \creg_reg[784]  ( .D(o[784]), .CLK(clk), .RST(rst), .I(g_init[784]), .Q(
        creg[784]) );
  DFF \creg_reg[785]  ( .D(o[785]), .CLK(clk), .RST(rst), .I(g_init[785]), .Q(
        creg[785]) );
  DFF \creg_reg[786]  ( .D(o[786]), .CLK(clk), .RST(rst), .I(g_init[786]), .Q(
        creg[786]) );
  DFF \creg_reg[787]  ( .D(o[787]), .CLK(clk), .RST(rst), .I(g_init[787]), .Q(
        creg[787]) );
  DFF \creg_reg[788]  ( .D(o[788]), .CLK(clk), .RST(rst), .I(g_init[788]), .Q(
        creg[788]) );
  DFF \creg_reg[789]  ( .D(o[789]), .CLK(clk), .RST(rst), .I(g_init[789]), .Q(
        creg[789]) );
  DFF \creg_reg[790]  ( .D(o[790]), .CLK(clk), .RST(rst), .I(g_init[790]), .Q(
        creg[790]) );
  DFF \creg_reg[791]  ( .D(o[791]), .CLK(clk), .RST(rst), .I(g_init[791]), .Q(
        creg[791]) );
  DFF \creg_reg[792]  ( .D(o[792]), .CLK(clk), .RST(rst), .I(g_init[792]), .Q(
        creg[792]) );
  DFF \creg_reg[793]  ( .D(o[793]), .CLK(clk), .RST(rst), .I(g_init[793]), .Q(
        creg[793]) );
  DFF \creg_reg[794]  ( .D(o[794]), .CLK(clk), .RST(rst), .I(g_init[794]), .Q(
        creg[794]) );
  DFF \creg_reg[795]  ( .D(o[795]), .CLK(clk), .RST(rst), .I(g_init[795]), .Q(
        creg[795]) );
  DFF \creg_reg[796]  ( .D(o[796]), .CLK(clk), .RST(rst), .I(g_init[796]), .Q(
        creg[796]) );
  DFF \creg_reg[797]  ( .D(o[797]), .CLK(clk), .RST(rst), .I(g_init[797]), .Q(
        creg[797]) );
  DFF \creg_reg[798]  ( .D(o[798]), .CLK(clk), .RST(rst), .I(g_init[798]), .Q(
        creg[798]) );
  DFF \creg_reg[799]  ( .D(o[799]), .CLK(clk), .RST(rst), .I(g_init[799]), .Q(
        creg[799]) );
  DFF \creg_reg[800]  ( .D(o[800]), .CLK(clk), .RST(rst), .I(g_init[800]), .Q(
        creg[800]) );
  DFF \creg_reg[801]  ( .D(o[801]), .CLK(clk), .RST(rst), .I(g_init[801]), .Q(
        creg[801]) );
  DFF \creg_reg[802]  ( .D(o[802]), .CLK(clk), .RST(rst), .I(g_init[802]), .Q(
        creg[802]) );
  DFF \creg_reg[803]  ( .D(o[803]), .CLK(clk), .RST(rst), .I(g_init[803]), .Q(
        creg[803]) );
  DFF \creg_reg[804]  ( .D(o[804]), .CLK(clk), .RST(rst), .I(g_init[804]), .Q(
        creg[804]) );
  DFF \creg_reg[805]  ( .D(o[805]), .CLK(clk), .RST(rst), .I(g_init[805]), .Q(
        creg[805]) );
  DFF \creg_reg[806]  ( .D(o[806]), .CLK(clk), .RST(rst), .I(g_init[806]), .Q(
        creg[806]) );
  DFF \creg_reg[807]  ( .D(o[807]), .CLK(clk), .RST(rst), .I(g_init[807]), .Q(
        creg[807]) );
  DFF \creg_reg[808]  ( .D(o[808]), .CLK(clk), .RST(rst), .I(g_init[808]), .Q(
        creg[808]) );
  DFF \creg_reg[809]  ( .D(o[809]), .CLK(clk), .RST(rst), .I(g_init[809]), .Q(
        creg[809]) );
  DFF \creg_reg[810]  ( .D(o[810]), .CLK(clk), .RST(rst), .I(g_init[810]), .Q(
        creg[810]) );
  DFF \creg_reg[811]  ( .D(o[811]), .CLK(clk), .RST(rst), .I(g_init[811]), .Q(
        creg[811]) );
  DFF \creg_reg[812]  ( .D(o[812]), .CLK(clk), .RST(rst), .I(g_init[812]), .Q(
        creg[812]) );
  DFF \creg_reg[813]  ( .D(o[813]), .CLK(clk), .RST(rst), .I(g_init[813]), .Q(
        creg[813]) );
  DFF \creg_reg[814]  ( .D(o[814]), .CLK(clk), .RST(rst), .I(g_init[814]), .Q(
        creg[814]) );
  DFF \creg_reg[815]  ( .D(o[815]), .CLK(clk), .RST(rst), .I(g_init[815]), .Q(
        creg[815]) );
  DFF \creg_reg[816]  ( .D(o[816]), .CLK(clk), .RST(rst), .I(g_init[816]), .Q(
        creg[816]) );
  DFF \creg_reg[817]  ( .D(o[817]), .CLK(clk), .RST(rst), .I(g_init[817]), .Q(
        creg[817]) );
  DFF \creg_reg[818]  ( .D(o[818]), .CLK(clk), .RST(rst), .I(g_init[818]), .Q(
        creg[818]) );
  DFF \creg_reg[819]  ( .D(o[819]), .CLK(clk), .RST(rst), .I(g_init[819]), .Q(
        creg[819]) );
  DFF \creg_reg[820]  ( .D(o[820]), .CLK(clk), .RST(rst), .I(g_init[820]), .Q(
        creg[820]) );
  DFF \creg_reg[821]  ( .D(o[821]), .CLK(clk), .RST(rst), .I(g_init[821]), .Q(
        creg[821]) );
  DFF \creg_reg[822]  ( .D(o[822]), .CLK(clk), .RST(rst), .I(g_init[822]), .Q(
        creg[822]) );
  DFF \creg_reg[823]  ( .D(o[823]), .CLK(clk), .RST(rst), .I(g_init[823]), .Q(
        creg[823]) );
  DFF \creg_reg[824]  ( .D(o[824]), .CLK(clk), .RST(rst), .I(g_init[824]), .Q(
        creg[824]) );
  DFF \creg_reg[825]  ( .D(o[825]), .CLK(clk), .RST(rst), .I(g_init[825]), .Q(
        creg[825]) );
  DFF \creg_reg[826]  ( .D(o[826]), .CLK(clk), .RST(rst), .I(g_init[826]), .Q(
        creg[826]) );
  DFF \creg_reg[827]  ( .D(o[827]), .CLK(clk), .RST(rst), .I(g_init[827]), .Q(
        creg[827]) );
  DFF \creg_reg[828]  ( .D(o[828]), .CLK(clk), .RST(rst), .I(g_init[828]), .Q(
        creg[828]) );
  DFF \creg_reg[829]  ( .D(o[829]), .CLK(clk), .RST(rst), .I(g_init[829]), .Q(
        creg[829]) );
  DFF \creg_reg[830]  ( .D(o[830]), .CLK(clk), .RST(rst), .I(g_init[830]), .Q(
        creg[830]) );
  DFF \creg_reg[831]  ( .D(o[831]), .CLK(clk), .RST(rst), .I(g_init[831]), .Q(
        creg[831]) );
  DFF \creg_reg[832]  ( .D(o[832]), .CLK(clk), .RST(rst), .I(g_init[832]), .Q(
        creg[832]) );
  DFF \creg_reg[833]  ( .D(o[833]), .CLK(clk), .RST(rst), .I(g_init[833]), .Q(
        creg[833]) );
  DFF \creg_reg[834]  ( .D(o[834]), .CLK(clk), .RST(rst), .I(g_init[834]), .Q(
        creg[834]) );
  DFF \creg_reg[835]  ( .D(o[835]), .CLK(clk), .RST(rst), .I(g_init[835]), .Q(
        creg[835]) );
  DFF \creg_reg[836]  ( .D(o[836]), .CLK(clk), .RST(rst), .I(g_init[836]), .Q(
        creg[836]) );
  DFF \creg_reg[837]  ( .D(o[837]), .CLK(clk), .RST(rst), .I(g_init[837]), .Q(
        creg[837]) );
  DFF \creg_reg[838]  ( .D(o[838]), .CLK(clk), .RST(rst), .I(g_init[838]), .Q(
        creg[838]) );
  DFF \creg_reg[839]  ( .D(o[839]), .CLK(clk), .RST(rst), .I(g_init[839]), .Q(
        creg[839]) );
  DFF \creg_reg[840]  ( .D(o[840]), .CLK(clk), .RST(rst), .I(g_init[840]), .Q(
        creg[840]) );
  DFF \creg_reg[841]  ( .D(o[841]), .CLK(clk), .RST(rst), .I(g_init[841]), .Q(
        creg[841]) );
  DFF \creg_reg[842]  ( .D(o[842]), .CLK(clk), .RST(rst), .I(g_init[842]), .Q(
        creg[842]) );
  DFF \creg_reg[843]  ( .D(o[843]), .CLK(clk), .RST(rst), .I(g_init[843]), .Q(
        creg[843]) );
  DFF \creg_reg[844]  ( .D(o[844]), .CLK(clk), .RST(rst), .I(g_init[844]), .Q(
        creg[844]) );
  DFF \creg_reg[845]  ( .D(o[845]), .CLK(clk), .RST(rst), .I(g_init[845]), .Q(
        creg[845]) );
  DFF \creg_reg[846]  ( .D(o[846]), .CLK(clk), .RST(rst), .I(g_init[846]), .Q(
        creg[846]) );
  DFF \creg_reg[847]  ( .D(o[847]), .CLK(clk), .RST(rst), .I(g_init[847]), .Q(
        creg[847]) );
  DFF \creg_reg[848]  ( .D(o[848]), .CLK(clk), .RST(rst), .I(g_init[848]), .Q(
        creg[848]) );
  DFF \creg_reg[849]  ( .D(o[849]), .CLK(clk), .RST(rst), .I(g_init[849]), .Q(
        creg[849]) );
  DFF \creg_reg[850]  ( .D(o[850]), .CLK(clk), .RST(rst), .I(g_init[850]), .Q(
        creg[850]) );
  DFF \creg_reg[851]  ( .D(o[851]), .CLK(clk), .RST(rst), .I(g_init[851]), .Q(
        creg[851]) );
  DFF \creg_reg[852]  ( .D(o[852]), .CLK(clk), .RST(rst), .I(g_init[852]), .Q(
        creg[852]) );
  DFF \creg_reg[853]  ( .D(o[853]), .CLK(clk), .RST(rst), .I(g_init[853]), .Q(
        creg[853]) );
  DFF \creg_reg[854]  ( .D(o[854]), .CLK(clk), .RST(rst), .I(g_init[854]), .Q(
        creg[854]) );
  DFF \creg_reg[855]  ( .D(o[855]), .CLK(clk), .RST(rst), .I(g_init[855]), .Q(
        creg[855]) );
  DFF \creg_reg[856]  ( .D(o[856]), .CLK(clk), .RST(rst), .I(g_init[856]), .Q(
        creg[856]) );
  DFF \creg_reg[857]  ( .D(o[857]), .CLK(clk), .RST(rst), .I(g_init[857]), .Q(
        creg[857]) );
  DFF \creg_reg[858]  ( .D(o[858]), .CLK(clk), .RST(rst), .I(g_init[858]), .Q(
        creg[858]) );
  DFF \creg_reg[859]  ( .D(o[859]), .CLK(clk), .RST(rst), .I(g_init[859]), .Q(
        creg[859]) );
  DFF \creg_reg[860]  ( .D(o[860]), .CLK(clk), .RST(rst), .I(g_init[860]), .Q(
        creg[860]) );
  DFF \creg_reg[861]  ( .D(o[861]), .CLK(clk), .RST(rst), .I(g_init[861]), .Q(
        creg[861]) );
  DFF \creg_reg[862]  ( .D(o[862]), .CLK(clk), .RST(rst), .I(g_init[862]), .Q(
        creg[862]) );
  DFF \creg_reg[863]  ( .D(o[863]), .CLK(clk), .RST(rst), .I(g_init[863]), .Q(
        creg[863]) );
  DFF \creg_reg[864]  ( .D(o[864]), .CLK(clk), .RST(rst), .I(g_init[864]), .Q(
        creg[864]) );
  DFF \creg_reg[865]  ( .D(o[865]), .CLK(clk), .RST(rst), .I(g_init[865]), .Q(
        creg[865]) );
  DFF \creg_reg[866]  ( .D(o[866]), .CLK(clk), .RST(rst), .I(g_init[866]), .Q(
        creg[866]) );
  DFF \creg_reg[867]  ( .D(o[867]), .CLK(clk), .RST(rst), .I(g_init[867]), .Q(
        creg[867]) );
  DFF \creg_reg[868]  ( .D(o[868]), .CLK(clk), .RST(rst), .I(g_init[868]), .Q(
        creg[868]) );
  DFF \creg_reg[869]  ( .D(o[869]), .CLK(clk), .RST(rst), .I(g_init[869]), .Q(
        creg[869]) );
  DFF \creg_reg[870]  ( .D(o[870]), .CLK(clk), .RST(rst), .I(g_init[870]), .Q(
        creg[870]) );
  DFF \creg_reg[871]  ( .D(o[871]), .CLK(clk), .RST(rst), .I(g_init[871]), .Q(
        creg[871]) );
  DFF \creg_reg[872]  ( .D(o[872]), .CLK(clk), .RST(rst), .I(g_init[872]), .Q(
        creg[872]) );
  DFF \creg_reg[873]  ( .D(o[873]), .CLK(clk), .RST(rst), .I(g_init[873]), .Q(
        creg[873]) );
  DFF \creg_reg[874]  ( .D(o[874]), .CLK(clk), .RST(rst), .I(g_init[874]), .Q(
        creg[874]) );
  DFF \creg_reg[875]  ( .D(o[875]), .CLK(clk), .RST(rst), .I(g_init[875]), .Q(
        creg[875]) );
  DFF \creg_reg[876]  ( .D(o[876]), .CLK(clk), .RST(rst), .I(g_init[876]), .Q(
        creg[876]) );
  DFF \creg_reg[877]  ( .D(o[877]), .CLK(clk), .RST(rst), .I(g_init[877]), .Q(
        creg[877]) );
  DFF \creg_reg[878]  ( .D(o[878]), .CLK(clk), .RST(rst), .I(g_init[878]), .Q(
        creg[878]) );
  DFF \creg_reg[879]  ( .D(o[879]), .CLK(clk), .RST(rst), .I(g_init[879]), .Q(
        creg[879]) );
  DFF \creg_reg[880]  ( .D(o[880]), .CLK(clk), .RST(rst), .I(g_init[880]), .Q(
        creg[880]) );
  DFF \creg_reg[881]  ( .D(o[881]), .CLK(clk), .RST(rst), .I(g_init[881]), .Q(
        creg[881]) );
  DFF \creg_reg[882]  ( .D(o[882]), .CLK(clk), .RST(rst), .I(g_init[882]), .Q(
        creg[882]) );
  DFF \creg_reg[883]  ( .D(o[883]), .CLK(clk), .RST(rst), .I(g_init[883]), .Q(
        creg[883]) );
  DFF \creg_reg[884]  ( .D(o[884]), .CLK(clk), .RST(rst), .I(g_init[884]), .Q(
        creg[884]) );
  DFF \creg_reg[885]  ( .D(o[885]), .CLK(clk), .RST(rst), .I(g_init[885]), .Q(
        creg[885]) );
  DFF \creg_reg[886]  ( .D(o[886]), .CLK(clk), .RST(rst), .I(g_init[886]), .Q(
        creg[886]) );
  DFF \creg_reg[887]  ( .D(o[887]), .CLK(clk), .RST(rst), .I(g_init[887]), .Q(
        creg[887]) );
  DFF \creg_reg[888]  ( .D(o[888]), .CLK(clk), .RST(rst), .I(g_init[888]), .Q(
        creg[888]) );
  DFF \creg_reg[889]  ( .D(o[889]), .CLK(clk), .RST(rst), .I(g_init[889]), .Q(
        creg[889]) );
  DFF \creg_reg[890]  ( .D(o[890]), .CLK(clk), .RST(rst), .I(g_init[890]), .Q(
        creg[890]) );
  DFF \creg_reg[891]  ( .D(o[891]), .CLK(clk), .RST(rst), .I(g_init[891]), .Q(
        creg[891]) );
  DFF \creg_reg[892]  ( .D(o[892]), .CLK(clk), .RST(rst), .I(g_init[892]), .Q(
        creg[892]) );
  DFF \creg_reg[893]  ( .D(o[893]), .CLK(clk), .RST(rst), .I(g_init[893]), .Q(
        creg[893]) );
  DFF \creg_reg[894]  ( .D(o[894]), .CLK(clk), .RST(rst), .I(g_init[894]), .Q(
        creg[894]) );
  DFF \creg_reg[895]  ( .D(o[895]), .CLK(clk), .RST(rst), .I(g_init[895]), .Q(
        creg[895]) );
  DFF \creg_reg[896]  ( .D(o[896]), .CLK(clk), .RST(rst), .I(g_init[896]), .Q(
        creg[896]) );
  DFF \creg_reg[897]  ( .D(o[897]), .CLK(clk), .RST(rst), .I(g_init[897]), .Q(
        creg[897]) );
  DFF \creg_reg[898]  ( .D(o[898]), .CLK(clk), .RST(rst), .I(g_init[898]), .Q(
        creg[898]) );
  DFF \creg_reg[899]  ( .D(o[899]), .CLK(clk), .RST(rst), .I(g_init[899]), .Q(
        creg[899]) );
  DFF \creg_reg[900]  ( .D(o[900]), .CLK(clk), .RST(rst), .I(g_init[900]), .Q(
        creg[900]) );
  DFF \creg_reg[901]  ( .D(o[901]), .CLK(clk), .RST(rst), .I(g_init[901]), .Q(
        creg[901]) );
  DFF \creg_reg[902]  ( .D(o[902]), .CLK(clk), .RST(rst), .I(g_init[902]), .Q(
        creg[902]) );
  DFF \creg_reg[903]  ( .D(o[903]), .CLK(clk), .RST(rst), .I(g_init[903]), .Q(
        creg[903]) );
  DFF \creg_reg[904]  ( .D(o[904]), .CLK(clk), .RST(rst), .I(g_init[904]), .Q(
        creg[904]) );
  DFF \creg_reg[905]  ( .D(o[905]), .CLK(clk), .RST(rst), .I(g_init[905]), .Q(
        creg[905]) );
  DFF \creg_reg[906]  ( .D(o[906]), .CLK(clk), .RST(rst), .I(g_init[906]), .Q(
        creg[906]) );
  DFF \creg_reg[907]  ( .D(o[907]), .CLK(clk), .RST(rst), .I(g_init[907]), .Q(
        creg[907]) );
  DFF \creg_reg[908]  ( .D(o[908]), .CLK(clk), .RST(rst), .I(g_init[908]), .Q(
        creg[908]) );
  DFF \creg_reg[909]  ( .D(o[909]), .CLK(clk), .RST(rst), .I(g_init[909]), .Q(
        creg[909]) );
  DFF \creg_reg[910]  ( .D(o[910]), .CLK(clk), .RST(rst), .I(g_init[910]), .Q(
        creg[910]) );
  DFF \creg_reg[911]  ( .D(o[911]), .CLK(clk), .RST(rst), .I(g_init[911]), .Q(
        creg[911]) );
  DFF \creg_reg[912]  ( .D(o[912]), .CLK(clk), .RST(rst), .I(g_init[912]), .Q(
        creg[912]) );
  DFF \creg_reg[913]  ( .D(o[913]), .CLK(clk), .RST(rst), .I(g_init[913]), .Q(
        creg[913]) );
  DFF \creg_reg[914]  ( .D(o[914]), .CLK(clk), .RST(rst), .I(g_init[914]), .Q(
        creg[914]) );
  DFF \creg_reg[915]  ( .D(o[915]), .CLK(clk), .RST(rst), .I(g_init[915]), .Q(
        creg[915]) );
  DFF \creg_reg[916]  ( .D(o[916]), .CLK(clk), .RST(rst), .I(g_init[916]), .Q(
        creg[916]) );
  DFF \creg_reg[917]  ( .D(o[917]), .CLK(clk), .RST(rst), .I(g_init[917]), .Q(
        creg[917]) );
  DFF \creg_reg[918]  ( .D(o[918]), .CLK(clk), .RST(rst), .I(g_init[918]), .Q(
        creg[918]) );
  DFF \creg_reg[919]  ( .D(o[919]), .CLK(clk), .RST(rst), .I(g_init[919]), .Q(
        creg[919]) );
  DFF \creg_reg[920]  ( .D(o[920]), .CLK(clk), .RST(rst), .I(g_init[920]), .Q(
        creg[920]) );
  DFF \creg_reg[921]  ( .D(o[921]), .CLK(clk), .RST(rst), .I(g_init[921]), .Q(
        creg[921]) );
  DFF \creg_reg[922]  ( .D(o[922]), .CLK(clk), .RST(rst), .I(g_init[922]), .Q(
        creg[922]) );
  DFF \creg_reg[923]  ( .D(o[923]), .CLK(clk), .RST(rst), .I(g_init[923]), .Q(
        creg[923]) );
  DFF \creg_reg[924]  ( .D(o[924]), .CLK(clk), .RST(rst), .I(g_init[924]), .Q(
        creg[924]) );
  DFF \creg_reg[925]  ( .D(o[925]), .CLK(clk), .RST(rst), .I(g_init[925]), .Q(
        creg[925]) );
  DFF \creg_reg[926]  ( .D(o[926]), .CLK(clk), .RST(rst), .I(g_init[926]), .Q(
        creg[926]) );
  DFF \creg_reg[927]  ( .D(o[927]), .CLK(clk), .RST(rst), .I(g_init[927]), .Q(
        creg[927]) );
  DFF \creg_reg[928]  ( .D(o[928]), .CLK(clk), .RST(rst), .I(g_init[928]), .Q(
        creg[928]) );
  DFF \creg_reg[929]  ( .D(o[929]), .CLK(clk), .RST(rst), .I(g_init[929]), .Q(
        creg[929]) );
  DFF \creg_reg[930]  ( .D(o[930]), .CLK(clk), .RST(rst), .I(g_init[930]), .Q(
        creg[930]) );
  DFF \creg_reg[931]  ( .D(o[931]), .CLK(clk), .RST(rst), .I(g_init[931]), .Q(
        creg[931]) );
  DFF \creg_reg[932]  ( .D(o[932]), .CLK(clk), .RST(rst), .I(g_init[932]), .Q(
        creg[932]) );
  DFF \creg_reg[933]  ( .D(o[933]), .CLK(clk), .RST(rst), .I(g_init[933]), .Q(
        creg[933]) );
  DFF \creg_reg[934]  ( .D(o[934]), .CLK(clk), .RST(rst), .I(g_init[934]), .Q(
        creg[934]) );
  DFF \creg_reg[935]  ( .D(o[935]), .CLK(clk), .RST(rst), .I(g_init[935]), .Q(
        creg[935]) );
  DFF \creg_reg[936]  ( .D(o[936]), .CLK(clk), .RST(rst), .I(g_init[936]), .Q(
        creg[936]) );
  DFF \creg_reg[937]  ( .D(o[937]), .CLK(clk), .RST(rst), .I(g_init[937]), .Q(
        creg[937]) );
  DFF \creg_reg[938]  ( .D(o[938]), .CLK(clk), .RST(rst), .I(g_init[938]), .Q(
        creg[938]) );
  DFF \creg_reg[939]  ( .D(o[939]), .CLK(clk), .RST(rst), .I(g_init[939]), .Q(
        creg[939]) );
  DFF \creg_reg[940]  ( .D(o[940]), .CLK(clk), .RST(rst), .I(g_init[940]), .Q(
        creg[940]) );
  DFF \creg_reg[941]  ( .D(o[941]), .CLK(clk), .RST(rst), .I(g_init[941]), .Q(
        creg[941]) );
  DFF \creg_reg[942]  ( .D(o[942]), .CLK(clk), .RST(rst), .I(g_init[942]), .Q(
        creg[942]) );
  DFF \creg_reg[943]  ( .D(o[943]), .CLK(clk), .RST(rst), .I(g_init[943]), .Q(
        creg[943]) );
  DFF \creg_reg[944]  ( .D(o[944]), .CLK(clk), .RST(rst), .I(g_init[944]), .Q(
        creg[944]) );
  DFF \creg_reg[945]  ( .D(o[945]), .CLK(clk), .RST(rst), .I(g_init[945]), .Q(
        creg[945]) );
  DFF \creg_reg[946]  ( .D(o[946]), .CLK(clk), .RST(rst), .I(g_init[946]), .Q(
        creg[946]) );
  DFF \creg_reg[947]  ( .D(o[947]), .CLK(clk), .RST(rst), .I(g_init[947]), .Q(
        creg[947]) );
  DFF \creg_reg[948]  ( .D(o[948]), .CLK(clk), .RST(rst), .I(g_init[948]), .Q(
        creg[948]) );
  DFF \creg_reg[949]  ( .D(o[949]), .CLK(clk), .RST(rst), .I(g_init[949]), .Q(
        creg[949]) );
  DFF \creg_reg[950]  ( .D(o[950]), .CLK(clk), .RST(rst), .I(g_init[950]), .Q(
        creg[950]) );
  DFF \creg_reg[951]  ( .D(o[951]), .CLK(clk), .RST(rst), .I(g_init[951]), .Q(
        creg[951]) );
  DFF \creg_reg[952]  ( .D(o[952]), .CLK(clk), .RST(rst), .I(g_init[952]), .Q(
        creg[952]) );
  DFF \creg_reg[953]  ( .D(o[953]), .CLK(clk), .RST(rst), .I(g_init[953]), .Q(
        creg[953]) );
  DFF \creg_reg[954]  ( .D(o[954]), .CLK(clk), .RST(rst), .I(g_init[954]), .Q(
        creg[954]) );
  DFF \creg_reg[955]  ( .D(o[955]), .CLK(clk), .RST(rst), .I(g_init[955]), .Q(
        creg[955]) );
  DFF \creg_reg[956]  ( .D(o[956]), .CLK(clk), .RST(rst), .I(g_init[956]), .Q(
        creg[956]) );
  DFF \creg_reg[957]  ( .D(o[957]), .CLK(clk), .RST(rst), .I(g_init[957]), .Q(
        creg[957]) );
  DFF \creg_reg[958]  ( .D(o[958]), .CLK(clk), .RST(rst), .I(g_init[958]), .Q(
        creg[958]) );
  DFF \creg_reg[959]  ( .D(o[959]), .CLK(clk), .RST(rst), .I(g_init[959]), .Q(
        creg[959]) );
  DFF \creg_reg[960]  ( .D(o[960]), .CLK(clk), .RST(rst), .I(g_init[960]), .Q(
        creg[960]) );
  DFF \creg_reg[961]  ( .D(o[961]), .CLK(clk), .RST(rst), .I(g_init[961]), .Q(
        creg[961]) );
  DFF \creg_reg[962]  ( .D(o[962]), .CLK(clk), .RST(rst), .I(g_init[962]), .Q(
        creg[962]) );
  DFF \creg_reg[963]  ( .D(o[963]), .CLK(clk), .RST(rst), .I(g_init[963]), .Q(
        creg[963]) );
  DFF \creg_reg[964]  ( .D(o[964]), .CLK(clk), .RST(rst), .I(g_init[964]), .Q(
        creg[964]) );
  DFF \creg_reg[965]  ( .D(o[965]), .CLK(clk), .RST(rst), .I(g_init[965]), .Q(
        creg[965]) );
  DFF \creg_reg[966]  ( .D(o[966]), .CLK(clk), .RST(rst), .I(g_init[966]), .Q(
        creg[966]) );
  DFF \creg_reg[967]  ( .D(o[967]), .CLK(clk), .RST(rst), .I(g_init[967]), .Q(
        creg[967]) );
  DFF \creg_reg[968]  ( .D(o[968]), .CLK(clk), .RST(rst), .I(g_init[968]), .Q(
        creg[968]) );
  DFF \creg_reg[969]  ( .D(o[969]), .CLK(clk), .RST(rst), .I(g_init[969]), .Q(
        creg[969]) );
  DFF \creg_reg[970]  ( .D(o[970]), .CLK(clk), .RST(rst), .I(g_init[970]), .Q(
        creg[970]) );
  DFF \creg_reg[971]  ( .D(o[971]), .CLK(clk), .RST(rst), .I(g_init[971]), .Q(
        creg[971]) );
  DFF \creg_reg[972]  ( .D(o[972]), .CLK(clk), .RST(rst), .I(g_init[972]), .Q(
        creg[972]) );
  DFF \creg_reg[973]  ( .D(o[973]), .CLK(clk), .RST(rst), .I(g_init[973]), .Q(
        creg[973]) );
  DFF \creg_reg[974]  ( .D(o[974]), .CLK(clk), .RST(rst), .I(g_init[974]), .Q(
        creg[974]) );
  DFF \creg_reg[975]  ( .D(o[975]), .CLK(clk), .RST(rst), .I(g_init[975]), .Q(
        creg[975]) );
  DFF \creg_reg[976]  ( .D(o[976]), .CLK(clk), .RST(rst), .I(g_init[976]), .Q(
        creg[976]) );
  DFF \creg_reg[977]  ( .D(o[977]), .CLK(clk), .RST(rst), .I(g_init[977]), .Q(
        creg[977]) );
  DFF \creg_reg[978]  ( .D(o[978]), .CLK(clk), .RST(rst), .I(g_init[978]), .Q(
        creg[978]) );
  DFF \creg_reg[979]  ( .D(o[979]), .CLK(clk), .RST(rst), .I(g_init[979]), .Q(
        creg[979]) );
  DFF \creg_reg[980]  ( .D(o[980]), .CLK(clk), .RST(rst), .I(g_init[980]), .Q(
        creg[980]) );
  DFF \creg_reg[981]  ( .D(o[981]), .CLK(clk), .RST(rst), .I(g_init[981]), .Q(
        creg[981]) );
  DFF \creg_reg[982]  ( .D(o[982]), .CLK(clk), .RST(rst), .I(g_init[982]), .Q(
        creg[982]) );
  DFF \creg_reg[983]  ( .D(o[983]), .CLK(clk), .RST(rst), .I(g_init[983]), .Q(
        creg[983]) );
  DFF \creg_reg[984]  ( .D(o[984]), .CLK(clk), .RST(rst), .I(g_init[984]), .Q(
        creg[984]) );
  DFF \creg_reg[985]  ( .D(o[985]), .CLK(clk), .RST(rst), .I(g_init[985]), .Q(
        creg[985]) );
  DFF \creg_reg[986]  ( .D(o[986]), .CLK(clk), .RST(rst), .I(g_init[986]), .Q(
        creg[986]) );
  DFF \creg_reg[987]  ( .D(o[987]), .CLK(clk), .RST(rst), .I(g_init[987]), .Q(
        creg[987]) );
  DFF \creg_reg[988]  ( .D(o[988]), .CLK(clk), .RST(rst), .I(g_init[988]), .Q(
        creg[988]) );
  DFF \creg_reg[989]  ( .D(o[989]), .CLK(clk), .RST(rst), .I(g_init[989]), .Q(
        creg[989]) );
  DFF \creg_reg[990]  ( .D(o[990]), .CLK(clk), .RST(rst), .I(g_init[990]), .Q(
        creg[990]) );
  DFF \creg_reg[991]  ( .D(o[991]), .CLK(clk), .RST(rst), .I(g_init[991]), .Q(
        creg[991]) );
  DFF \creg_reg[992]  ( .D(o[992]), .CLK(clk), .RST(rst), .I(g_init[992]), .Q(
        creg[992]) );
  DFF \creg_reg[993]  ( .D(o[993]), .CLK(clk), .RST(rst), .I(g_init[993]), .Q(
        creg[993]) );
  DFF \creg_reg[994]  ( .D(o[994]), .CLK(clk), .RST(rst), .I(g_init[994]), .Q(
        creg[994]) );
  DFF \creg_reg[995]  ( .D(o[995]), .CLK(clk), .RST(rst), .I(g_init[995]), .Q(
        creg[995]) );
  DFF \creg_reg[996]  ( .D(o[996]), .CLK(clk), .RST(rst), .I(g_init[996]), .Q(
        creg[996]) );
  DFF \creg_reg[997]  ( .D(o[997]), .CLK(clk), .RST(rst), .I(g_init[997]), .Q(
        creg[997]) );
  DFF \creg_reg[998]  ( .D(o[998]), .CLK(clk), .RST(rst), .I(g_init[998]), .Q(
        creg[998]) );
  DFF \creg_reg[999]  ( .D(o[999]), .CLK(clk), .RST(rst), .I(g_init[999]), .Q(
        creg[999]) );
  DFF \creg_reg[1000]  ( .D(o[1000]), .CLK(clk), .RST(rst), .I(g_init[1000]), 
        .Q(creg[1000]) );
  DFF \creg_reg[1001]  ( .D(o[1001]), .CLK(clk), .RST(rst), .I(g_init[1001]), 
        .Q(creg[1001]) );
  DFF \creg_reg[1002]  ( .D(o[1002]), .CLK(clk), .RST(rst), .I(g_init[1002]), 
        .Q(creg[1002]) );
  DFF \creg_reg[1003]  ( .D(o[1003]), .CLK(clk), .RST(rst), .I(g_init[1003]), 
        .Q(creg[1003]) );
  DFF \creg_reg[1004]  ( .D(o[1004]), .CLK(clk), .RST(rst), .I(g_init[1004]), 
        .Q(creg[1004]) );
  DFF \creg_reg[1005]  ( .D(o[1005]), .CLK(clk), .RST(rst), .I(g_init[1005]), 
        .Q(creg[1005]) );
  DFF \creg_reg[1006]  ( .D(o[1006]), .CLK(clk), .RST(rst), .I(g_init[1006]), 
        .Q(creg[1006]) );
  DFF \creg_reg[1007]  ( .D(o[1007]), .CLK(clk), .RST(rst), .I(g_init[1007]), 
        .Q(creg[1007]) );
  DFF \creg_reg[1008]  ( .D(o[1008]), .CLK(clk), .RST(rst), .I(g_init[1008]), 
        .Q(creg[1008]) );
  DFF \creg_reg[1009]  ( .D(o[1009]), .CLK(clk), .RST(rst), .I(g_init[1009]), 
        .Q(creg[1009]) );
  DFF \creg_reg[1010]  ( .D(o[1010]), .CLK(clk), .RST(rst), .I(g_init[1010]), 
        .Q(creg[1010]) );
  DFF \creg_reg[1011]  ( .D(o[1011]), .CLK(clk), .RST(rst), .I(g_init[1011]), 
        .Q(creg[1011]) );
  DFF \creg_reg[1012]  ( .D(o[1012]), .CLK(clk), .RST(rst), .I(g_init[1012]), 
        .Q(creg[1012]) );
  DFF \creg_reg[1013]  ( .D(o[1013]), .CLK(clk), .RST(rst), .I(g_init[1013]), 
        .Q(creg[1013]) );
  DFF \creg_reg[1014]  ( .D(o[1014]), .CLK(clk), .RST(rst), .I(g_init[1014]), 
        .Q(creg[1014]) );
  DFF \creg_reg[1015]  ( .D(o[1015]), .CLK(clk), .RST(rst), .I(g_init[1015]), 
        .Q(creg[1015]) );
  DFF \creg_reg[1016]  ( .D(o[1016]), .CLK(clk), .RST(rst), .I(g_init[1016]), 
        .Q(creg[1016]) );
  DFF \creg_reg[1017]  ( .D(o[1017]), .CLK(clk), .RST(rst), .I(g_init[1017]), 
        .Q(creg[1017]) );
  DFF \creg_reg[1018]  ( .D(o[1018]), .CLK(clk), .RST(rst), .I(g_init[1018]), 
        .Q(creg[1018]) );
  DFF \creg_reg[1019]  ( .D(o[1019]), .CLK(clk), .RST(rst), .I(g_init[1019]), 
        .Q(creg[1019]) );
  DFF \creg_reg[1020]  ( .D(o[1020]), .CLK(clk), .RST(rst), .I(g_init[1020]), 
        .Q(creg[1020]) );
  DFF \creg_reg[1021]  ( .D(o[1021]), .CLK(clk), .RST(rst), .I(g_init[1021]), 
        .Q(creg[1021]) );
  DFF \creg_reg[1022]  ( .D(o[1022]), .CLK(clk), .RST(rst), .I(g_init[1022]), 
        .Q(creg[1022]) );
  DFF \creg_reg[1023]  ( .D(o[1023]), .CLK(clk), .RST(rst), .I(g_init[1023]), 
        .Q(creg[1023]) );
  DFF \modmult_1/zreg_reg[1024]  ( .D(\modmult_1/zout[0][1024] ), .CLK(clk), 
        .RST(start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][1024] ) );
  DFF \modmult_1/zreg_reg[1023]  ( .D(mod_mult_o[1023]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][1023] ) );
  DFF \modmult_1/zreg_reg[1022]  ( .D(mod_mult_o[1022]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][1022] ) );
  DFF \modmult_1/zreg_reg[1021]  ( .D(mod_mult_o[1021]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][1021] ) );
  DFF \modmult_1/zreg_reg[1020]  ( .D(mod_mult_o[1020]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][1020] ) );
  DFF \modmult_1/zreg_reg[1019]  ( .D(mod_mult_o[1019]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][1019] ) );
  DFF \modmult_1/zreg_reg[1018]  ( .D(mod_mult_o[1018]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][1018] ) );
  DFF \modmult_1/zreg_reg[1017]  ( .D(mod_mult_o[1017]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][1017] ) );
  DFF \modmult_1/zreg_reg[1016]  ( .D(mod_mult_o[1016]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][1016] ) );
  DFF \modmult_1/zreg_reg[1015]  ( .D(mod_mult_o[1015]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][1015] ) );
  DFF \modmult_1/zreg_reg[1014]  ( .D(mod_mult_o[1014]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][1014] ) );
  DFF \modmult_1/zreg_reg[1013]  ( .D(mod_mult_o[1013]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][1013] ) );
  DFF \modmult_1/zreg_reg[1012]  ( .D(mod_mult_o[1012]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][1012] ) );
  DFF \modmult_1/zreg_reg[1011]  ( .D(mod_mult_o[1011]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][1011] ) );
  DFF \modmult_1/zreg_reg[1010]  ( .D(mod_mult_o[1010]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][1010] ) );
  DFF \modmult_1/zreg_reg[1009]  ( .D(mod_mult_o[1009]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][1009] ) );
  DFF \modmult_1/zreg_reg[1008]  ( .D(mod_mult_o[1008]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][1008] ) );
  DFF \modmult_1/zreg_reg[1007]  ( .D(mod_mult_o[1007]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][1007] ) );
  DFF \modmult_1/zreg_reg[1006]  ( .D(mod_mult_o[1006]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][1006] ) );
  DFF \modmult_1/zreg_reg[1005]  ( .D(mod_mult_o[1005]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][1005] ) );
  DFF \modmult_1/zreg_reg[1004]  ( .D(mod_mult_o[1004]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][1004] ) );
  DFF \modmult_1/zreg_reg[1003]  ( .D(mod_mult_o[1003]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][1003] ) );
  DFF \modmult_1/zreg_reg[1002]  ( .D(mod_mult_o[1002]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][1002] ) );
  DFF \modmult_1/zreg_reg[1001]  ( .D(mod_mult_o[1001]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][1001] ) );
  DFF \modmult_1/zreg_reg[1000]  ( .D(mod_mult_o[1000]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][1000] ) );
  DFF \modmult_1/zreg_reg[999]  ( .D(mod_mult_o[999]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][999] ) );
  DFF \modmult_1/zreg_reg[998]  ( .D(mod_mult_o[998]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][998] ) );
  DFF \modmult_1/zreg_reg[997]  ( .D(mod_mult_o[997]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][997] ) );
  DFF \modmult_1/zreg_reg[996]  ( .D(mod_mult_o[996]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][996] ) );
  DFF \modmult_1/zreg_reg[995]  ( .D(mod_mult_o[995]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][995] ) );
  DFF \modmult_1/zreg_reg[994]  ( .D(mod_mult_o[994]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][994] ) );
  DFF \modmult_1/zreg_reg[993]  ( .D(mod_mult_o[993]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][993] ) );
  DFF \modmult_1/zreg_reg[992]  ( .D(mod_mult_o[992]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][992] ) );
  DFF \modmult_1/zreg_reg[991]  ( .D(mod_mult_o[991]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][991] ) );
  DFF \modmult_1/zreg_reg[990]  ( .D(mod_mult_o[990]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][990] ) );
  DFF \modmult_1/zreg_reg[989]  ( .D(mod_mult_o[989]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][989] ) );
  DFF \modmult_1/zreg_reg[988]  ( .D(mod_mult_o[988]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][988] ) );
  DFF \modmult_1/zreg_reg[987]  ( .D(mod_mult_o[987]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][987] ) );
  DFF \modmult_1/zreg_reg[986]  ( .D(mod_mult_o[986]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][986] ) );
  DFF \modmult_1/zreg_reg[985]  ( .D(mod_mult_o[985]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][985] ) );
  DFF \modmult_1/zreg_reg[984]  ( .D(mod_mult_o[984]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][984] ) );
  DFF \modmult_1/zreg_reg[983]  ( .D(mod_mult_o[983]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][983] ) );
  DFF \modmult_1/zreg_reg[982]  ( .D(mod_mult_o[982]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][982] ) );
  DFF \modmult_1/zreg_reg[981]  ( .D(mod_mult_o[981]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][981] ) );
  DFF \modmult_1/zreg_reg[980]  ( .D(mod_mult_o[980]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][980] ) );
  DFF \modmult_1/zreg_reg[979]  ( .D(mod_mult_o[979]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][979] ) );
  DFF \modmult_1/zreg_reg[978]  ( .D(mod_mult_o[978]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][978] ) );
  DFF \modmult_1/zreg_reg[977]  ( .D(mod_mult_o[977]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][977] ) );
  DFF \modmult_1/zreg_reg[976]  ( .D(mod_mult_o[976]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][976] ) );
  DFF \modmult_1/zreg_reg[975]  ( .D(mod_mult_o[975]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][975] ) );
  DFF \modmult_1/zreg_reg[974]  ( .D(mod_mult_o[974]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][974] ) );
  DFF \modmult_1/zreg_reg[973]  ( .D(mod_mult_o[973]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][973] ) );
  DFF \modmult_1/zreg_reg[972]  ( .D(mod_mult_o[972]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][972] ) );
  DFF \modmult_1/zreg_reg[971]  ( .D(mod_mult_o[971]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][971] ) );
  DFF \modmult_1/zreg_reg[970]  ( .D(mod_mult_o[970]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][970] ) );
  DFF \modmult_1/zreg_reg[969]  ( .D(mod_mult_o[969]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][969] ) );
  DFF \modmult_1/zreg_reg[968]  ( .D(mod_mult_o[968]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][968] ) );
  DFF \modmult_1/zreg_reg[967]  ( .D(mod_mult_o[967]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][967] ) );
  DFF \modmult_1/zreg_reg[966]  ( .D(mod_mult_o[966]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][966] ) );
  DFF \modmult_1/zreg_reg[965]  ( .D(mod_mult_o[965]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][965] ) );
  DFF \modmult_1/zreg_reg[964]  ( .D(mod_mult_o[964]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][964] ) );
  DFF \modmult_1/zreg_reg[963]  ( .D(mod_mult_o[963]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][963] ) );
  DFF \modmult_1/zreg_reg[962]  ( .D(mod_mult_o[962]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][962] ) );
  DFF \modmult_1/zreg_reg[961]  ( .D(mod_mult_o[961]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][961] ) );
  DFF \modmult_1/zreg_reg[960]  ( .D(mod_mult_o[960]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][960] ) );
  DFF \modmult_1/zreg_reg[959]  ( .D(mod_mult_o[959]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][959] ) );
  DFF \modmult_1/zreg_reg[958]  ( .D(mod_mult_o[958]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][958] ) );
  DFF \modmult_1/zreg_reg[957]  ( .D(mod_mult_o[957]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][957] ) );
  DFF \modmult_1/zreg_reg[956]  ( .D(mod_mult_o[956]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][956] ) );
  DFF \modmult_1/zreg_reg[955]  ( .D(mod_mult_o[955]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][955] ) );
  DFF \modmult_1/zreg_reg[954]  ( .D(mod_mult_o[954]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][954] ) );
  DFF \modmult_1/zreg_reg[953]  ( .D(mod_mult_o[953]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][953] ) );
  DFF \modmult_1/zreg_reg[952]  ( .D(mod_mult_o[952]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][952] ) );
  DFF \modmult_1/zreg_reg[951]  ( .D(mod_mult_o[951]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][951] ) );
  DFF \modmult_1/zreg_reg[950]  ( .D(mod_mult_o[950]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][950] ) );
  DFF \modmult_1/zreg_reg[949]  ( .D(mod_mult_o[949]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][949] ) );
  DFF \modmult_1/zreg_reg[948]  ( .D(mod_mult_o[948]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][948] ) );
  DFF \modmult_1/zreg_reg[947]  ( .D(mod_mult_o[947]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][947] ) );
  DFF \modmult_1/zreg_reg[946]  ( .D(mod_mult_o[946]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][946] ) );
  DFF \modmult_1/zreg_reg[945]  ( .D(mod_mult_o[945]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][945] ) );
  DFF \modmult_1/zreg_reg[944]  ( .D(mod_mult_o[944]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][944] ) );
  DFF \modmult_1/zreg_reg[943]  ( .D(mod_mult_o[943]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][943] ) );
  DFF \modmult_1/zreg_reg[942]  ( .D(mod_mult_o[942]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][942] ) );
  DFF \modmult_1/zreg_reg[941]  ( .D(mod_mult_o[941]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][941] ) );
  DFF \modmult_1/zreg_reg[940]  ( .D(mod_mult_o[940]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][940] ) );
  DFF \modmult_1/zreg_reg[939]  ( .D(mod_mult_o[939]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][939] ) );
  DFF \modmult_1/zreg_reg[938]  ( .D(mod_mult_o[938]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][938] ) );
  DFF \modmult_1/zreg_reg[937]  ( .D(mod_mult_o[937]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][937] ) );
  DFF \modmult_1/zreg_reg[936]  ( .D(mod_mult_o[936]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][936] ) );
  DFF \modmult_1/zreg_reg[935]  ( .D(mod_mult_o[935]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][935] ) );
  DFF \modmult_1/zreg_reg[934]  ( .D(mod_mult_o[934]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][934] ) );
  DFF \modmult_1/zreg_reg[933]  ( .D(mod_mult_o[933]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][933] ) );
  DFF \modmult_1/zreg_reg[932]  ( .D(mod_mult_o[932]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][932] ) );
  DFF \modmult_1/zreg_reg[931]  ( .D(mod_mult_o[931]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][931] ) );
  DFF \modmult_1/zreg_reg[930]  ( .D(mod_mult_o[930]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][930] ) );
  DFF \modmult_1/zreg_reg[929]  ( .D(mod_mult_o[929]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][929] ) );
  DFF \modmult_1/zreg_reg[928]  ( .D(mod_mult_o[928]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][928] ) );
  DFF \modmult_1/zreg_reg[927]  ( .D(mod_mult_o[927]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][927] ) );
  DFF \modmult_1/zreg_reg[926]  ( .D(mod_mult_o[926]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][926] ) );
  DFF \modmult_1/zreg_reg[925]  ( .D(mod_mult_o[925]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][925] ) );
  DFF \modmult_1/zreg_reg[924]  ( .D(mod_mult_o[924]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][924] ) );
  DFF \modmult_1/zreg_reg[923]  ( .D(mod_mult_o[923]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][923] ) );
  DFF \modmult_1/zreg_reg[922]  ( .D(mod_mult_o[922]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][922] ) );
  DFF \modmult_1/zreg_reg[921]  ( .D(mod_mult_o[921]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][921] ) );
  DFF \modmult_1/zreg_reg[920]  ( .D(mod_mult_o[920]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][920] ) );
  DFF \modmult_1/zreg_reg[919]  ( .D(mod_mult_o[919]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][919] ) );
  DFF \modmult_1/zreg_reg[918]  ( .D(mod_mult_o[918]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][918] ) );
  DFF \modmult_1/zreg_reg[917]  ( .D(mod_mult_o[917]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][917] ) );
  DFF \modmult_1/zreg_reg[916]  ( .D(mod_mult_o[916]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][916] ) );
  DFF \modmult_1/zreg_reg[915]  ( .D(mod_mult_o[915]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][915] ) );
  DFF \modmult_1/zreg_reg[914]  ( .D(mod_mult_o[914]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][914] ) );
  DFF \modmult_1/zreg_reg[913]  ( .D(mod_mult_o[913]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][913] ) );
  DFF \modmult_1/zreg_reg[912]  ( .D(mod_mult_o[912]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][912] ) );
  DFF \modmult_1/zreg_reg[911]  ( .D(mod_mult_o[911]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][911] ) );
  DFF \modmult_1/zreg_reg[910]  ( .D(mod_mult_o[910]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][910] ) );
  DFF \modmult_1/zreg_reg[909]  ( .D(mod_mult_o[909]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][909] ) );
  DFF \modmult_1/zreg_reg[908]  ( .D(mod_mult_o[908]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][908] ) );
  DFF \modmult_1/zreg_reg[907]  ( .D(mod_mult_o[907]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][907] ) );
  DFF \modmult_1/zreg_reg[906]  ( .D(mod_mult_o[906]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][906] ) );
  DFF \modmult_1/zreg_reg[905]  ( .D(mod_mult_o[905]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][905] ) );
  DFF \modmult_1/zreg_reg[904]  ( .D(mod_mult_o[904]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][904] ) );
  DFF \modmult_1/zreg_reg[903]  ( .D(mod_mult_o[903]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][903] ) );
  DFF \modmult_1/zreg_reg[902]  ( .D(mod_mult_o[902]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][902] ) );
  DFF \modmult_1/zreg_reg[901]  ( .D(mod_mult_o[901]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][901] ) );
  DFF \modmult_1/zreg_reg[900]  ( .D(mod_mult_o[900]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][900] ) );
  DFF \modmult_1/zreg_reg[899]  ( .D(mod_mult_o[899]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][899] ) );
  DFF \modmult_1/zreg_reg[898]  ( .D(mod_mult_o[898]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][898] ) );
  DFF \modmult_1/zreg_reg[897]  ( .D(mod_mult_o[897]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][897] ) );
  DFF \modmult_1/zreg_reg[896]  ( .D(mod_mult_o[896]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][896] ) );
  DFF \modmult_1/zreg_reg[895]  ( .D(mod_mult_o[895]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][895] ) );
  DFF \modmult_1/zreg_reg[894]  ( .D(mod_mult_o[894]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][894] ) );
  DFF \modmult_1/zreg_reg[893]  ( .D(mod_mult_o[893]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][893] ) );
  DFF \modmult_1/zreg_reg[892]  ( .D(mod_mult_o[892]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][892] ) );
  DFF \modmult_1/zreg_reg[891]  ( .D(mod_mult_o[891]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][891] ) );
  DFF \modmult_1/zreg_reg[890]  ( .D(mod_mult_o[890]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][890] ) );
  DFF \modmult_1/zreg_reg[889]  ( .D(mod_mult_o[889]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][889] ) );
  DFF \modmult_1/zreg_reg[888]  ( .D(mod_mult_o[888]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][888] ) );
  DFF \modmult_1/zreg_reg[887]  ( .D(mod_mult_o[887]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][887] ) );
  DFF \modmult_1/zreg_reg[886]  ( .D(mod_mult_o[886]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][886] ) );
  DFF \modmult_1/zreg_reg[885]  ( .D(mod_mult_o[885]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][885] ) );
  DFF \modmult_1/zreg_reg[884]  ( .D(mod_mult_o[884]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][884] ) );
  DFF \modmult_1/zreg_reg[883]  ( .D(mod_mult_o[883]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][883] ) );
  DFF \modmult_1/zreg_reg[882]  ( .D(mod_mult_o[882]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][882] ) );
  DFF \modmult_1/zreg_reg[881]  ( .D(mod_mult_o[881]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][881] ) );
  DFF \modmult_1/zreg_reg[880]  ( .D(mod_mult_o[880]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][880] ) );
  DFF \modmult_1/zreg_reg[879]  ( .D(mod_mult_o[879]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][879] ) );
  DFF \modmult_1/zreg_reg[878]  ( .D(mod_mult_o[878]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][878] ) );
  DFF \modmult_1/zreg_reg[877]  ( .D(mod_mult_o[877]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][877] ) );
  DFF \modmult_1/zreg_reg[876]  ( .D(mod_mult_o[876]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][876] ) );
  DFF \modmult_1/zreg_reg[875]  ( .D(mod_mult_o[875]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][875] ) );
  DFF \modmult_1/zreg_reg[874]  ( .D(mod_mult_o[874]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][874] ) );
  DFF \modmult_1/zreg_reg[873]  ( .D(mod_mult_o[873]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][873] ) );
  DFF \modmult_1/zreg_reg[872]  ( .D(mod_mult_o[872]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][872] ) );
  DFF \modmult_1/zreg_reg[871]  ( .D(mod_mult_o[871]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][871] ) );
  DFF \modmult_1/zreg_reg[870]  ( .D(mod_mult_o[870]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][870] ) );
  DFF \modmult_1/zreg_reg[869]  ( .D(mod_mult_o[869]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][869] ) );
  DFF \modmult_1/zreg_reg[868]  ( .D(mod_mult_o[868]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][868] ) );
  DFF \modmult_1/zreg_reg[867]  ( .D(mod_mult_o[867]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][867] ) );
  DFF \modmult_1/zreg_reg[866]  ( .D(mod_mult_o[866]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][866] ) );
  DFF \modmult_1/zreg_reg[865]  ( .D(mod_mult_o[865]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][865] ) );
  DFF \modmult_1/zreg_reg[864]  ( .D(mod_mult_o[864]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][864] ) );
  DFF \modmult_1/zreg_reg[863]  ( .D(mod_mult_o[863]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][863] ) );
  DFF \modmult_1/zreg_reg[862]  ( .D(mod_mult_o[862]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][862] ) );
  DFF \modmult_1/zreg_reg[861]  ( .D(mod_mult_o[861]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][861] ) );
  DFF \modmult_1/zreg_reg[860]  ( .D(mod_mult_o[860]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][860] ) );
  DFF \modmult_1/zreg_reg[859]  ( .D(mod_mult_o[859]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][859] ) );
  DFF \modmult_1/zreg_reg[858]  ( .D(mod_mult_o[858]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][858] ) );
  DFF \modmult_1/zreg_reg[857]  ( .D(mod_mult_o[857]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][857] ) );
  DFF \modmult_1/zreg_reg[856]  ( .D(mod_mult_o[856]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][856] ) );
  DFF \modmult_1/zreg_reg[855]  ( .D(mod_mult_o[855]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][855] ) );
  DFF \modmult_1/zreg_reg[854]  ( .D(mod_mult_o[854]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][854] ) );
  DFF \modmult_1/zreg_reg[853]  ( .D(mod_mult_o[853]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][853] ) );
  DFF \modmult_1/zreg_reg[852]  ( .D(mod_mult_o[852]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][852] ) );
  DFF \modmult_1/zreg_reg[851]  ( .D(mod_mult_o[851]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][851] ) );
  DFF \modmult_1/zreg_reg[850]  ( .D(mod_mult_o[850]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][850] ) );
  DFF \modmult_1/zreg_reg[849]  ( .D(mod_mult_o[849]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][849] ) );
  DFF \modmult_1/zreg_reg[848]  ( .D(mod_mult_o[848]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][848] ) );
  DFF \modmult_1/zreg_reg[847]  ( .D(mod_mult_o[847]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][847] ) );
  DFF \modmult_1/zreg_reg[846]  ( .D(mod_mult_o[846]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][846] ) );
  DFF \modmult_1/zreg_reg[845]  ( .D(mod_mult_o[845]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][845] ) );
  DFF \modmult_1/zreg_reg[844]  ( .D(mod_mult_o[844]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][844] ) );
  DFF \modmult_1/zreg_reg[843]  ( .D(mod_mult_o[843]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][843] ) );
  DFF \modmult_1/zreg_reg[842]  ( .D(mod_mult_o[842]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][842] ) );
  DFF \modmult_1/zreg_reg[841]  ( .D(mod_mult_o[841]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][841] ) );
  DFF \modmult_1/zreg_reg[840]  ( .D(mod_mult_o[840]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][840] ) );
  DFF \modmult_1/zreg_reg[839]  ( .D(mod_mult_o[839]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][839] ) );
  DFF \modmult_1/zreg_reg[838]  ( .D(mod_mult_o[838]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][838] ) );
  DFF \modmult_1/zreg_reg[837]  ( .D(mod_mult_o[837]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][837] ) );
  DFF \modmult_1/zreg_reg[836]  ( .D(mod_mult_o[836]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][836] ) );
  DFF \modmult_1/zreg_reg[835]  ( .D(mod_mult_o[835]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][835] ) );
  DFF \modmult_1/zreg_reg[834]  ( .D(mod_mult_o[834]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][834] ) );
  DFF \modmult_1/zreg_reg[833]  ( .D(mod_mult_o[833]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][833] ) );
  DFF \modmult_1/zreg_reg[832]  ( .D(mod_mult_o[832]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][832] ) );
  DFF \modmult_1/zreg_reg[831]  ( .D(mod_mult_o[831]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][831] ) );
  DFF \modmult_1/zreg_reg[830]  ( .D(mod_mult_o[830]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][830] ) );
  DFF \modmult_1/zreg_reg[829]  ( .D(mod_mult_o[829]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][829] ) );
  DFF \modmult_1/zreg_reg[828]  ( .D(mod_mult_o[828]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][828] ) );
  DFF \modmult_1/zreg_reg[827]  ( .D(mod_mult_o[827]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][827] ) );
  DFF \modmult_1/zreg_reg[826]  ( .D(mod_mult_o[826]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][826] ) );
  DFF \modmult_1/zreg_reg[825]  ( .D(mod_mult_o[825]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][825] ) );
  DFF \modmult_1/zreg_reg[824]  ( .D(mod_mult_o[824]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][824] ) );
  DFF \modmult_1/zreg_reg[823]  ( .D(mod_mult_o[823]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][823] ) );
  DFF \modmult_1/zreg_reg[822]  ( .D(mod_mult_o[822]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][822] ) );
  DFF \modmult_1/zreg_reg[821]  ( .D(mod_mult_o[821]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][821] ) );
  DFF \modmult_1/zreg_reg[820]  ( .D(mod_mult_o[820]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][820] ) );
  DFF \modmult_1/zreg_reg[819]  ( .D(mod_mult_o[819]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][819] ) );
  DFF \modmult_1/zreg_reg[818]  ( .D(mod_mult_o[818]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][818] ) );
  DFF \modmult_1/zreg_reg[817]  ( .D(mod_mult_o[817]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][817] ) );
  DFF \modmult_1/zreg_reg[816]  ( .D(mod_mult_o[816]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][816] ) );
  DFF \modmult_1/zreg_reg[815]  ( .D(mod_mult_o[815]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][815] ) );
  DFF \modmult_1/zreg_reg[814]  ( .D(mod_mult_o[814]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][814] ) );
  DFF \modmult_1/zreg_reg[813]  ( .D(mod_mult_o[813]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][813] ) );
  DFF \modmult_1/zreg_reg[812]  ( .D(mod_mult_o[812]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][812] ) );
  DFF \modmult_1/zreg_reg[811]  ( .D(mod_mult_o[811]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][811] ) );
  DFF \modmult_1/zreg_reg[810]  ( .D(mod_mult_o[810]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][810] ) );
  DFF \modmult_1/zreg_reg[809]  ( .D(mod_mult_o[809]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][809] ) );
  DFF \modmult_1/zreg_reg[808]  ( .D(mod_mult_o[808]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][808] ) );
  DFF \modmult_1/zreg_reg[807]  ( .D(mod_mult_o[807]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][807] ) );
  DFF \modmult_1/zreg_reg[806]  ( .D(mod_mult_o[806]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][806] ) );
  DFF \modmult_1/zreg_reg[805]  ( .D(mod_mult_o[805]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][805] ) );
  DFF \modmult_1/zreg_reg[804]  ( .D(mod_mult_o[804]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][804] ) );
  DFF \modmult_1/zreg_reg[803]  ( .D(mod_mult_o[803]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][803] ) );
  DFF \modmult_1/zreg_reg[802]  ( .D(mod_mult_o[802]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][802] ) );
  DFF \modmult_1/zreg_reg[801]  ( .D(mod_mult_o[801]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][801] ) );
  DFF \modmult_1/zreg_reg[800]  ( .D(mod_mult_o[800]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][800] ) );
  DFF \modmult_1/zreg_reg[799]  ( .D(mod_mult_o[799]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][799] ) );
  DFF \modmult_1/zreg_reg[798]  ( .D(mod_mult_o[798]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][798] ) );
  DFF \modmult_1/zreg_reg[797]  ( .D(mod_mult_o[797]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][797] ) );
  DFF \modmult_1/zreg_reg[796]  ( .D(mod_mult_o[796]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][796] ) );
  DFF \modmult_1/zreg_reg[795]  ( .D(mod_mult_o[795]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][795] ) );
  DFF \modmult_1/zreg_reg[794]  ( .D(mod_mult_o[794]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][794] ) );
  DFF \modmult_1/zreg_reg[793]  ( .D(mod_mult_o[793]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][793] ) );
  DFF \modmult_1/zreg_reg[792]  ( .D(mod_mult_o[792]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][792] ) );
  DFF \modmult_1/zreg_reg[791]  ( .D(mod_mult_o[791]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][791] ) );
  DFF \modmult_1/zreg_reg[790]  ( .D(mod_mult_o[790]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][790] ) );
  DFF \modmult_1/zreg_reg[789]  ( .D(mod_mult_o[789]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][789] ) );
  DFF \modmult_1/zreg_reg[788]  ( .D(mod_mult_o[788]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][788] ) );
  DFF \modmult_1/zreg_reg[787]  ( .D(mod_mult_o[787]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][787] ) );
  DFF \modmult_1/zreg_reg[786]  ( .D(mod_mult_o[786]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][786] ) );
  DFF \modmult_1/zreg_reg[785]  ( .D(mod_mult_o[785]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][785] ) );
  DFF \modmult_1/zreg_reg[784]  ( .D(mod_mult_o[784]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][784] ) );
  DFF \modmult_1/zreg_reg[783]  ( .D(mod_mult_o[783]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][783] ) );
  DFF \modmult_1/zreg_reg[782]  ( .D(mod_mult_o[782]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][782] ) );
  DFF \modmult_1/zreg_reg[781]  ( .D(mod_mult_o[781]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][781] ) );
  DFF \modmult_1/zreg_reg[780]  ( .D(mod_mult_o[780]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][780] ) );
  DFF \modmult_1/zreg_reg[779]  ( .D(mod_mult_o[779]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][779] ) );
  DFF \modmult_1/zreg_reg[778]  ( .D(mod_mult_o[778]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][778] ) );
  DFF \modmult_1/zreg_reg[777]  ( .D(mod_mult_o[777]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][777] ) );
  DFF \modmult_1/zreg_reg[776]  ( .D(mod_mult_o[776]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][776] ) );
  DFF \modmult_1/zreg_reg[775]  ( .D(mod_mult_o[775]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][775] ) );
  DFF \modmult_1/zreg_reg[774]  ( .D(mod_mult_o[774]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][774] ) );
  DFF \modmult_1/zreg_reg[773]  ( .D(mod_mult_o[773]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][773] ) );
  DFF \modmult_1/zreg_reg[772]  ( .D(mod_mult_o[772]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][772] ) );
  DFF \modmult_1/zreg_reg[771]  ( .D(mod_mult_o[771]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][771] ) );
  DFF \modmult_1/zreg_reg[770]  ( .D(mod_mult_o[770]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][770] ) );
  DFF \modmult_1/zreg_reg[769]  ( .D(mod_mult_o[769]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][769] ) );
  DFF \modmult_1/zreg_reg[768]  ( .D(mod_mult_o[768]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][768] ) );
  DFF \modmult_1/zreg_reg[767]  ( .D(mod_mult_o[767]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][767] ) );
  DFF \modmult_1/zreg_reg[766]  ( .D(mod_mult_o[766]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][766] ) );
  DFF \modmult_1/zreg_reg[765]  ( .D(mod_mult_o[765]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][765] ) );
  DFF \modmult_1/zreg_reg[764]  ( .D(mod_mult_o[764]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][764] ) );
  DFF \modmult_1/zreg_reg[763]  ( .D(mod_mult_o[763]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][763] ) );
  DFF \modmult_1/zreg_reg[762]  ( .D(mod_mult_o[762]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][762] ) );
  DFF \modmult_1/zreg_reg[761]  ( .D(mod_mult_o[761]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][761] ) );
  DFF \modmult_1/zreg_reg[760]  ( .D(mod_mult_o[760]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][760] ) );
  DFF \modmult_1/zreg_reg[759]  ( .D(mod_mult_o[759]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][759] ) );
  DFF \modmult_1/zreg_reg[758]  ( .D(mod_mult_o[758]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][758] ) );
  DFF \modmult_1/zreg_reg[757]  ( .D(mod_mult_o[757]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][757] ) );
  DFF \modmult_1/zreg_reg[756]  ( .D(mod_mult_o[756]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][756] ) );
  DFF \modmult_1/zreg_reg[755]  ( .D(mod_mult_o[755]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][755] ) );
  DFF \modmult_1/zreg_reg[754]  ( .D(mod_mult_o[754]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][754] ) );
  DFF \modmult_1/zreg_reg[753]  ( .D(mod_mult_o[753]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][753] ) );
  DFF \modmult_1/zreg_reg[752]  ( .D(mod_mult_o[752]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][752] ) );
  DFF \modmult_1/zreg_reg[751]  ( .D(mod_mult_o[751]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][751] ) );
  DFF \modmult_1/zreg_reg[750]  ( .D(mod_mult_o[750]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][750] ) );
  DFF \modmult_1/zreg_reg[749]  ( .D(mod_mult_o[749]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][749] ) );
  DFF \modmult_1/zreg_reg[748]  ( .D(mod_mult_o[748]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][748] ) );
  DFF \modmult_1/zreg_reg[747]  ( .D(mod_mult_o[747]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][747] ) );
  DFF \modmult_1/zreg_reg[746]  ( .D(mod_mult_o[746]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][746] ) );
  DFF \modmult_1/zreg_reg[745]  ( .D(mod_mult_o[745]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][745] ) );
  DFF \modmult_1/zreg_reg[744]  ( .D(mod_mult_o[744]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][744] ) );
  DFF \modmult_1/zreg_reg[743]  ( .D(mod_mult_o[743]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][743] ) );
  DFF \modmult_1/zreg_reg[742]  ( .D(mod_mult_o[742]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][742] ) );
  DFF \modmult_1/zreg_reg[741]  ( .D(mod_mult_o[741]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][741] ) );
  DFF \modmult_1/zreg_reg[740]  ( .D(mod_mult_o[740]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][740] ) );
  DFF \modmult_1/zreg_reg[739]  ( .D(mod_mult_o[739]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][739] ) );
  DFF \modmult_1/zreg_reg[738]  ( .D(mod_mult_o[738]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][738] ) );
  DFF \modmult_1/zreg_reg[737]  ( .D(mod_mult_o[737]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][737] ) );
  DFF \modmult_1/zreg_reg[736]  ( .D(mod_mult_o[736]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][736] ) );
  DFF \modmult_1/zreg_reg[735]  ( .D(mod_mult_o[735]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][735] ) );
  DFF \modmult_1/zreg_reg[734]  ( .D(mod_mult_o[734]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][734] ) );
  DFF \modmult_1/zreg_reg[733]  ( .D(mod_mult_o[733]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][733] ) );
  DFF \modmult_1/zreg_reg[732]  ( .D(mod_mult_o[732]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][732] ) );
  DFF \modmult_1/zreg_reg[731]  ( .D(mod_mult_o[731]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][731] ) );
  DFF \modmult_1/zreg_reg[730]  ( .D(mod_mult_o[730]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][730] ) );
  DFF \modmult_1/zreg_reg[729]  ( .D(mod_mult_o[729]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][729] ) );
  DFF \modmult_1/zreg_reg[728]  ( .D(mod_mult_o[728]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][728] ) );
  DFF \modmult_1/zreg_reg[727]  ( .D(mod_mult_o[727]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][727] ) );
  DFF \modmult_1/zreg_reg[726]  ( .D(mod_mult_o[726]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][726] ) );
  DFF \modmult_1/zreg_reg[725]  ( .D(mod_mult_o[725]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][725] ) );
  DFF \modmult_1/zreg_reg[724]  ( .D(mod_mult_o[724]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][724] ) );
  DFF \modmult_1/zreg_reg[723]  ( .D(mod_mult_o[723]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][723] ) );
  DFF \modmult_1/zreg_reg[722]  ( .D(mod_mult_o[722]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][722] ) );
  DFF \modmult_1/zreg_reg[721]  ( .D(mod_mult_o[721]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][721] ) );
  DFF \modmult_1/zreg_reg[720]  ( .D(mod_mult_o[720]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][720] ) );
  DFF \modmult_1/zreg_reg[719]  ( .D(mod_mult_o[719]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][719] ) );
  DFF \modmult_1/zreg_reg[718]  ( .D(mod_mult_o[718]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][718] ) );
  DFF \modmult_1/zreg_reg[717]  ( .D(mod_mult_o[717]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][717] ) );
  DFF \modmult_1/zreg_reg[716]  ( .D(mod_mult_o[716]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][716] ) );
  DFF \modmult_1/zreg_reg[715]  ( .D(mod_mult_o[715]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][715] ) );
  DFF \modmult_1/zreg_reg[714]  ( .D(mod_mult_o[714]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][714] ) );
  DFF \modmult_1/zreg_reg[713]  ( .D(mod_mult_o[713]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][713] ) );
  DFF \modmult_1/zreg_reg[712]  ( .D(mod_mult_o[712]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][712] ) );
  DFF \modmult_1/zreg_reg[711]  ( .D(mod_mult_o[711]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][711] ) );
  DFF \modmult_1/zreg_reg[710]  ( .D(mod_mult_o[710]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][710] ) );
  DFF \modmult_1/zreg_reg[709]  ( .D(mod_mult_o[709]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][709] ) );
  DFF \modmult_1/zreg_reg[708]  ( .D(mod_mult_o[708]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][708] ) );
  DFF \modmult_1/zreg_reg[707]  ( .D(mod_mult_o[707]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][707] ) );
  DFF \modmult_1/zreg_reg[706]  ( .D(mod_mult_o[706]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][706] ) );
  DFF \modmult_1/zreg_reg[705]  ( .D(mod_mult_o[705]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][705] ) );
  DFF \modmult_1/zreg_reg[704]  ( .D(mod_mult_o[704]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][704] ) );
  DFF \modmult_1/zreg_reg[703]  ( .D(mod_mult_o[703]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][703] ) );
  DFF \modmult_1/zreg_reg[702]  ( .D(mod_mult_o[702]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][702] ) );
  DFF \modmult_1/zreg_reg[701]  ( .D(mod_mult_o[701]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][701] ) );
  DFF \modmult_1/zreg_reg[700]  ( .D(mod_mult_o[700]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][700] ) );
  DFF \modmult_1/zreg_reg[699]  ( .D(mod_mult_o[699]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][699] ) );
  DFF \modmult_1/zreg_reg[698]  ( .D(mod_mult_o[698]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][698] ) );
  DFF \modmult_1/zreg_reg[697]  ( .D(mod_mult_o[697]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][697] ) );
  DFF \modmult_1/zreg_reg[696]  ( .D(mod_mult_o[696]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][696] ) );
  DFF \modmult_1/zreg_reg[695]  ( .D(mod_mult_o[695]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][695] ) );
  DFF \modmult_1/zreg_reg[694]  ( .D(mod_mult_o[694]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][694] ) );
  DFF \modmult_1/zreg_reg[693]  ( .D(mod_mult_o[693]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][693] ) );
  DFF \modmult_1/zreg_reg[692]  ( .D(mod_mult_o[692]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][692] ) );
  DFF \modmult_1/zreg_reg[691]  ( .D(mod_mult_o[691]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][691] ) );
  DFF \modmult_1/zreg_reg[690]  ( .D(mod_mult_o[690]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][690] ) );
  DFF \modmult_1/zreg_reg[689]  ( .D(mod_mult_o[689]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][689] ) );
  DFF \modmult_1/zreg_reg[688]  ( .D(mod_mult_o[688]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][688] ) );
  DFF \modmult_1/zreg_reg[687]  ( .D(mod_mult_o[687]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][687] ) );
  DFF \modmult_1/zreg_reg[686]  ( .D(mod_mult_o[686]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][686] ) );
  DFF \modmult_1/zreg_reg[685]  ( .D(mod_mult_o[685]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][685] ) );
  DFF \modmult_1/zreg_reg[684]  ( .D(mod_mult_o[684]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][684] ) );
  DFF \modmult_1/zreg_reg[683]  ( .D(mod_mult_o[683]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][683] ) );
  DFF \modmult_1/zreg_reg[682]  ( .D(mod_mult_o[682]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][682] ) );
  DFF \modmult_1/zreg_reg[681]  ( .D(mod_mult_o[681]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][681] ) );
  DFF \modmult_1/zreg_reg[680]  ( .D(mod_mult_o[680]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][680] ) );
  DFF \modmult_1/zreg_reg[679]  ( .D(mod_mult_o[679]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][679] ) );
  DFF \modmult_1/zreg_reg[678]  ( .D(mod_mult_o[678]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][678] ) );
  DFF \modmult_1/zreg_reg[677]  ( .D(mod_mult_o[677]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][677] ) );
  DFF \modmult_1/zreg_reg[676]  ( .D(mod_mult_o[676]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][676] ) );
  DFF \modmult_1/zreg_reg[675]  ( .D(mod_mult_o[675]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][675] ) );
  DFF \modmult_1/zreg_reg[674]  ( .D(mod_mult_o[674]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][674] ) );
  DFF \modmult_1/zreg_reg[673]  ( .D(mod_mult_o[673]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][673] ) );
  DFF \modmult_1/zreg_reg[672]  ( .D(mod_mult_o[672]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][672] ) );
  DFF \modmult_1/zreg_reg[671]  ( .D(mod_mult_o[671]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][671] ) );
  DFF \modmult_1/zreg_reg[670]  ( .D(mod_mult_o[670]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][670] ) );
  DFF \modmult_1/zreg_reg[669]  ( .D(mod_mult_o[669]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][669] ) );
  DFF \modmult_1/zreg_reg[668]  ( .D(mod_mult_o[668]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][668] ) );
  DFF \modmult_1/zreg_reg[667]  ( .D(mod_mult_o[667]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][667] ) );
  DFF \modmult_1/zreg_reg[666]  ( .D(mod_mult_o[666]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][666] ) );
  DFF \modmult_1/zreg_reg[665]  ( .D(mod_mult_o[665]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][665] ) );
  DFF \modmult_1/zreg_reg[664]  ( .D(mod_mult_o[664]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][664] ) );
  DFF \modmult_1/zreg_reg[663]  ( .D(mod_mult_o[663]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][663] ) );
  DFF \modmult_1/zreg_reg[662]  ( .D(mod_mult_o[662]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][662] ) );
  DFF \modmult_1/zreg_reg[661]  ( .D(mod_mult_o[661]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][661] ) );
  DFF \modmult_1/zreg_reg[660]  ( .D(mod_mult_o[660]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][660] ) );
  DFF \modmult_1/zreg_reg[659]  ( .D(mod_mult_o[659]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][659] ) );
  DFF \modmult_1/zreg_reg[658]  ( .D(mod_mult_o[658]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][658] ) );
  DFF \modmult_1/zreg_reg[657]  ( .D(mod_mult_o[657]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][657] ) );
  DFF \modmult_1/zreg_reg[656]  ( .D(mod_mult_o[656]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][656] ) );
  DFF \modmult_1/zreg_reg[655]  ( .D(mod_mult_o[655]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][655] ) );
  DFF \modmult_1/zreg_reg[654]  ( .D(mod_mult_o[654]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][654] ) );
  DFF \modmult_1/zreg_reg[653]  ( .D(mod_mult_o[653]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][653] ) );
  DFF \modmult_1/zreg_reg[652]  ( .D(mod_mult_o[652]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][652] ) );
  DFF \modmult_1/zreg_reg[651]  ( .D(mod_mult_o[651]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][651] ) );
  DFF \modmult_1/zreg_reg[650]  ( .D(mod_mult_o[650]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][650] ) );
  DFF \modmult_1/zreg_reg[649]  ( .D(mod_mult_o[649]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][649] ) );
  DFF \modmult_1/zreg_reg[648]  ( .D(mod_mult_o[648]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][648] ) );
  DFF \modmult_1/zreg_reg[647]  ( .D(mod_mult_o[647]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][647] ) );
  DFF \modmult_1/zreg_reg[646]  ( .D(mod_mult_o[646]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][646] ) );
  DFF \modmult_1/zreg_reg[645]  ( .D(mod_mult_o[645]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][645] ) );
  DFF \modmult_1/zreg_reg[644]  ( .D(mod_mult_o[644]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][644] ) );
  DFF \modmult_1/zreg_reg[643]  ( .D(mod_mult_o[643]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][643] ) );
  DFF \modmult_1/zreg_reg[642]  ( .D(mod_mult_o[642]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][642] ) );
  DFF \modmult_1/zreg_reg[641]  ( .D(mod_mult_o[641]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][641] ) );
  DFF \modmult_1/zreg_reg[640]  ( .D(mod_mult_o[640]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][640] ) );
  DFF \modmult_1/zreg_reg[639]  ( .D(mod_mult_o[639]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][639] ) );
  DFF \modmult_1/zreg_reg[638]  ( .D(mod_mult_o[638]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][638] ) );
  DFF \modmult_1/zreg_reg[637]  ( .D(mod_mult_o[637]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][637] ) );
  DFF \modmult_1/zreg_reg[636]  ( .D(mod_mult_o[636]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][636] ) );
  DFF \modmult_1/zreg_reg[635]  ( .D(mod_mult_o[635]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][635] ) );
  DFF \modmult_1/zreg_reg[634]  ( .D(mod_mult_o[634]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][634] ) );
  DFF \modmult_1/zreg_reg[633]  ( .D(mod_mult_o[633]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][633] ) );
  DFF \modmult_1/zreg_reg[632]  ( .D(mod_mult_o[632]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][632] ) );
  DFF \modmult_1/zreg_reg[631]  ( .D(mod_mult_o[631]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][631] ) );
  DFF \modmult_1/zreg_reg[630]  ( .D(mod_mult_o[630]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][630] ) );
  DFF \modmult_1/zreg_reg[629]  ( .D(mod_mult_o[629]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][629] ) );
  DFF \modmult_1/zreg_reg[628]  ( .D(mod_mult_o[628]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][628] ) );
  DFF \modmult_1/zreg_reg[627]  ( .D(mod_mult_o[627]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][627] ) );
  DFF \modmult_1/zreg_reg[626]  ( .D(mod_mult_o[626]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][626] ) );
  DFF \modmult_1/zreg_reg[625]  ( .D(mod_mult_o[625]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][625] ) );
  DFF \modmult_1/zreg_reg[624]  ( .D(mod_mult_o[624]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][624] ) );
  DFF \modmult_1/zreg_reg[623]  ( .D(mod_mult_o[623]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][623] ) );
  DFF \modmult_1/zreg_reg[622]  ( .D(mod_mult_o[622]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][622] ) );
  DFF \modmult_1/zreg_reg[621]  ( .D(mod_mult_o[621]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][621] ) );
  DFF \modmult_1/zreg_reg[620]  ( .D(mod_mult_o[620]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][620] ) );
  DFF \modmult_1/zreg_reg[619]  ( .D(mod_mult_o[619]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][619] ) );
  DFF \modmult_1/zreg_reg[618]  ( .D(mod_mult_o[618]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][618] ) );
  DFF \modmult_1/zreg_reg[617]  ( .D(mod_mult_o[617]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][617] ) );
  DFF \modmult_1/zreg_reg[616]  ( .D(mod_mult_o[616]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][616] ) );
  DFF \modmult_1/zreg_reg[615]  ( .D(mod_mult_o[615]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][615] ) );
  DFF \modmult_1/zreg_reg[614]  ( .D(mod_mult_o[614]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][614] ) );
  DFF \modmult_1/zreg_reg[613]  ( .D(mod_mult_o[613]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][613] ) );
  DFF \modmult_1/zreg_reg[612]  ( .D(mod_mult_o[612]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][612] ) );
  DFF \modmult_1/zreg_reg[611]  ( .D(mod_mult_o[611]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][611] ) );
  DFF \modmult_1/zreg_reg[610]  ( .D(mod_mult_o[610]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][610] ) );
  DFF \modmult_1/zreg_reg[609]  ( .D(mod_mult_o[609]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][609] ) );
  DFF \modmult_1/zreg_reg[608]  ( .D(mod_mult_o[608]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][608] ) );
  DFF \modmult_1/zreg_reg[607]  ( .D(mod_mult_o[607]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][607] ) );
  DFF \modmult_1/zreg_reg[606]  ( .D(mod_mult_o[606]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][606] ) );
  DFF \modmult_1/zreg_reg[605]  ( .D(mod_mult_o[605]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][605] ) );
  DFF \modmult_1/zreg_reg[604]  ( .D(mod_mult_o[604]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][604] ) );
  DFF \modmult_1/zreg_reg[603]  ( .D(mod_mult_o[603]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][603] ) );
  DFF \modmult_1/zreg_reg[602]  ( .D(mod_mult_o[602]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][602] ) );
  DFF \modmult_1/zreg_reg[601]  ( .D(mod_mult_o[601]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][601] ) );
  DFF \modmult_1/zreg_reg[600]  ( .D(mod_mult_o[600]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][600] ) );
  DFF \modmult_1/zreg_reg[599]  ( .D(mod_mult_o[599]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][599] ) );
  DFF \modmult_1/zreg_reg[598]  ( .D(mod_mult_o[598]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][598] ) );
  DFF \modmult_1/zreg_reg[597]  ( .D(mod_mult_o[597]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][597] ) );
  DFF \modmult_1/zreg_reg[596]  ( .D(mod_mult_o[596]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][596] ) );
  DFF \modmult_1/zreg_reg[595]  ( .D(mod_mult_o[595]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][595] ) );
  DFF \modmult_1/zreg_reg[594]  ( .D(mod_mult_o[594]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][594] ) );
  DFF \modmult_1/zreg_reg[593]  ( .D(mod_mult_o[593]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][593] ) );
  DFF \modmult_1/zreg_reg[592]  ( .D(mod_mult_o[592]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][592] ) );
  DFF \modmult_1/zreg_reg[591]  ( .D(mod_mult_o[591]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][591] ) );
  DFF \modmult_1/zreg_reg[590]  ( .D(mod_mult_o[590]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][590] ) );
  DFF \modmult_1/zreg_reg[589]  ( .D(mod_mult_o[589]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][589] ) );
  DFF \modmult_1/zreg_reg[588]  ( .D(mod_mult_o[588]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][588] ) );
  DFF \modmult_1/zreg_reg[587]  ( .D(mod_mult_o[587]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][587] ) );
  DFF \modmult_1/zreg_reg[586]  ( .D(mod_mult_o[586]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][586] ) );
  DFF \modmult_1/zreg_reg[585]  ( .D(mod_mult_o[585]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][585] ) );
  DFF \modmult_1/zreg_reg[584]  ( .D(mod_mult_o[584]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][584] ) );
  DFF \modmult_1/zreg_reg[583]  ( .D(mod_mult_o[583]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][583] ) );
  DFF \modmult_1/zreg_reg[582]  ( .D(mod_mult_o[582]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][582] ) );
  DFF \modmult_1/zreg_reg[581]  ( .D(mod_mult_o[581]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][581] ) );
  DFF \modmult_1/zreg_reg[580]  ( .D(mod_mult_o[580]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][580] ) );
  DFF \modmult_1/zreg_reg[579]  ( .D(mod_mult_o[579]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][579] ) );
  DFF \modmult_1/zreg_reg[578]  ( .D(mod_mult_o[578]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][578] ) );
  DFF \modmult_1/zreg_reg[577]  ( .D(mod_mult_o[577]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][577] ) );
  DFF \modmult_1/zreg_reg[576]  ( .D(mod_mult_o[576]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][576] ) );
  DFF \modmult_1/zreg_reg[575]  ( .D(mod_mult_o[575]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][575] ) );
  DFF \modmult_1/zreg_reg[574]  ( .D(mod_mult_o[574]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][574] ) );
  DFF \modmult_1/zreg_reg[573]  ( .D(mod_mult_o[573]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][573] ) );
  DFF \modmult_1/zreg_reg[572]  ( .D(mod_mult_o[572]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][572] ) );
  DFF \modmult_1/zreg_reg[571]  ( .D(mod_mult_o[571]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][571] ) );
  DFF \modmult_1/zreg_reg[570]  ( .D(mod_mult_o[570]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][570] ) );
  DFF \modmult_1/zreg_reg[569]  ( .D(mod_mult_o[569]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][569] ) );
  DFF \modmult_1/zreg_reg[568]  ( .D(mod_mult_o[568]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][568] ) );
  DFF \modmult_1/zreg_reg[567]  ( .D(mod_mult_o[567]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][567] ) );
  DFF \modmult_1/zreg_reg[566]  ( .D(mod_mult_o[566]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][566] ) );
  DFF \modmult_1/zreg_reg[565]  ( .D(mod_mult_o[565]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][565] ) );
  DFF \modmult_1/zreg_reg[564]  ( .D(mod_mult_o[564]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][564] ) );
  DFF \modmult_1/zreg_reg[563]  ( .D(mod_mult_o[563]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][563] ) );
  DFF \modmult_1/zreg_reg[562]  ( .D(mod_mult_o[562]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][562] ) );
  DFF \modmult_1/zreg_reg[561]  ( .D(mod_mult_o[561]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][561] ) );
  DFF \modmult_1/zreg_reg[560]  ( .D(mod_mult_o[560]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][560] ) );
  DFF \modmult_1/zreg_reg[559]  ( .D(mod_mult_o[559]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][559] ) );
  DFF \modmult_1/zreg_reg[558]  ( .D(mod_mult_o[558]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][558] ) );
  DFF \modmult_1/zreg_reg[557]  ( .D(mod_mult_o[557]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][557] ) );
  DFF \modmult_1/zreg_reg[556]  ( .D(mod_mult_o[556]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][556] ) );
  DFF \modmult_1/zreg_reg[555]  ( .D(mod_mult_o[555]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][555] ) );
  DFF \modmult_1/zreg_reg[554]  ( .D(mod_mult_o[554]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][554] ) );
  DFF \modmult_1/zreg_reg[553]  ( .D(mod_mult_o[553]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][553] ) );
  DFF \modmult_1/zreg_reg[552]  ( .D(mod_mult_o[552]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][552] ) );
  DFF \modmult_1/zreg_reg[551]  ( .D(mod_mult_o[551]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][551] ) );
  DFF \modmult_1/zreg_reg[550]  ( .D(mod_mult_o[550]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][550] ) );
  DFF \modmult_1/zreg_reg[549]  ( .D(mod_mult_o[549]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][549] ) );
  DFF \modmult_1/zreg_reg[548]  ( .D(mod_mult_o[548]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][548] ) );
  DFF \modmult_1/zreg_reg[547]  ( .D(mod_mult_o[547]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][547] ) );
  DFF \modmult_1/zreg_reg[546]  ( .D(mod_mult_o[546]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][546] ) );
  DFF \modmult_1/zreg_reg[545]  ( .D(mod_mult_o[545]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][545] ) );
  DFF \modmult_1/zreg_reg[544]  ( .D(mod_mult_o[544]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][544] ) );
  DFF \modmult_1/zreg_reg[543]  ( .D(mod_mult_o[543]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][543] ) );
  DFF \modmult_1/zreg_reg[542]  ( .D(mod_mult_o[542]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][542] ) );
  DFF \modmult_1/zreg_reg[541]  ( .D(mod_mult_o[541]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][541] ) );
  DFF \modmult_1/zreg_reg[540]  ( .D(mod_mult_o[540]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][540] ) );
  DFF \modmult_1/zreg_reg[539]  ( .D(mod_mult_o[539]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][539] ) );
  DFF \modmult_1/zreg_reg[538]  ( .D(mod_mult_o[538]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][538] ) );
  DFF \modmult_1/zreg_reg[537]  ( .D(mod_mult_o[537]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][537] ) );
  DFF \modmult_1/zreg_reg[536]  ( .D(mod_mult_o[536]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][536] ) );
  DFF \modmult_1/zreg_reg[535]  ( .D(mod_mult_o[535]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][535] ) );
  DFF \modmult_1/zreg_reg[534]  ( .D(mod_mult_o[534]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][534] ) );
  DFF \modmult_1/zreg_reg[533]  ( .D(mod_mult_o[533]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][533] ) );
  DFF \modmult_1/zreg_reg[532]  ( .D(mod_mult_o[532]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][532] ) );
  DFF \modmult_1/zreg_reg[531]  ( .D(mod_mult_o[531]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][531] ) );
  DFF \modmult_1/zreg_reg[530]  ( .D(mod_mult_o[530]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][530] ) );
  DFF \modmult_1/zreg_reg[529]  ( .D(mod_mult_o[529]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][529] ) );
  DFF \modmult_1/zreg_reg[528]  ( .D(mod_mult_o[528]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][528] ) );
  DFF \modmult_1/zreg_reg[527]  ( .D(mod_mult_o[527]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][527] ) );
  DFF \modmult_1/zreg_reg[526]  ( .D(mod_mult_o[526]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][526] ) );
  DFF \modmult_1/zreg_reg[525]  ( .D(mod_mult_o[525]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][525] ) );
  DFF \modmult_1/zreg_reg[524]  ( .D(mod_mult_o[524]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][524] ) );
  DFF \modmult_1/zreg_reg[523]  ( .D(mod_mult_o[523]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][523] ) );
  DFF \modmult_1/zreg_reg[522]  ( .D(mod_mult_o[522]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][522] ) );
  DFF \modmult_1/zreg_reg[521]  ( .D(mod_mult_o[521]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][521] ) );
  DFF \modmult_1/zreg_reg[520]  ( .D(mod_mult_o[520]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][520] ) );
  DFF \modmult_1/zreg_reg[519]  ( .D(mod_mult_o[519]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][519] ) );
  DFF \modmult_1/zreg_reg[518]  ( .D(mod_mult_o[518]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][518] ) );
  DFF \modmult_1/zreg_reg[517]  ( .D(mod_mult_o[517]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][517] ) );
  DFF \modmult_1/zreg_reg[516]  ( .D(mod_mult_o[516]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][516] ) );
  DFF \modmult_1/zreg_reg[515]  ( .D(mod_mult_o[515]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][515] ) );
  DFF \modmult_1/zreg_reg[514]  ( .D(mod_mult_o[514]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][514] ) );
  DFF \modmult_1/zreg_reg[513]  ( .D(mod_mult_o[513]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][513] ) );
  DFF \modmult_1/zreg_reg[512]  ( .D(mod_mult_o[512]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][512] ) );
  DFF \modmult_1/zreg_reg[511]  ( .D(mod_mult_o[511]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][511] ) );
  DFF \modmult_1/zreg_reg[510]  ( .D(mod_mult_o[510]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][510] ) );
  DFF \modmult_1/zreg_reg[509]  ( .D(mod_mult_o[509]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][509] ) );
  DFF \modmult_1/zreg_reg[508]  ( .D(mod_mult_o[508]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][508] ) );
  DFF \modmult_1/zreg_reg[507]  ( .D(mod_mult_o[507]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][507] ) );
  DFF \modmult_1/zreg_reg[506]  ( .D(mod_mult_o[506]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][506] ) );
  DFF \modmult_1/zreg_reg[505]  ( .D(mod_mult_o[505]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][505] ) );
  DFF \modmult_1/zreg_reg[504]  ( .D(mod_mult_o[504]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][504] ) );
  DFF \modmult_1/zreg_reg[503]  ( .D(mod_mult_o[503]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][503] ) );
  DFF \modmult_1/zreg_reg[502]  ( .D(mod_mult_o[502]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][502] ) );
  DFF \modmult_1/zreg_reg[501]  ( .D(mod_mult_o[501]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][501] ) );
  DFF \modmult_1/zreg_reg[500]  ( .D(mod_mult_o[500]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][500] ) );
  DFF \modmult_1/zreg_reg[499]  ( .D(mod_mult_o[499]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][499] ) );
  DFF \modmult_1/zreg_reg[498]  ( .D(mod_mult_o[498]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][498] ) );
  DFF \modmult_1/zreg_reg[497]  ( .D(mod_mult_o[497]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][497] ) );
  DFF \modmult_1/zreg_reg[496]  ( .D(mod_mult_o[496]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][496] ) );
  DFF \modmult_1/zreg_reg[495]  ( .D(mod_mult_o[495]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][495] ) );
  DFF \modmult_1/zreg_reg[494]  ( .D(mod_mult_o[494]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][494] ) );
  DFF \modmult_1/zreg_reg[493]  ( .D(mod_mult_o[493]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][493] ) );
  DFF \modmult_1/zreg_reg[492]  ( .D(mod_mult_o[492]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][492] ) );
  DFF \modmult_1/zreg_reg[491]  ( .D(mod_mult_o[491]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][491] ) );
  DFF \modmult_1/zreg_reg[490]  ( .D(mod_mult_o[490]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][490] ) );
  DFF \modmult_1/zreg_reg[489]  ( .D(mod_mult_o[489]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][489] ) );
  DFF \modmult_1/zreg_reg[488]  ( .D(mod_mult_o[488]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][488] ) );
  DFF \modmult_1/zreg_reg[487]  ( .D(mod_mult_o[487]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][487] ) );
  DFF \modmult_1/zreg_reg[486]  ( .D(mod_mult_o[486]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][486] ) );
  DFF \modmult_1/zreg_reg[485]  ( .D(mod_mult_o[485]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][485] ) );
  DFF \modmult_1/zreg_reg[484]  ( .D(mod_mult_o[484]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][484] ) );
  DFF \modmult_1/zreg_reg[483]  ( .D(mod_mult_o[483]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][483] ) );
  DFF \modmult_1/zreg_reg[482]  ( .D(mod_mult_o[482]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][482] ) );
  DFF \modmult_1/zreg_reg[481]  ( .D(mod_mult_o[481]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][481] ) );
  DFF \modmult_1/zreg_reg[480]  ( .D(mod_mult_o[480]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][480] ) );
  DFF \modmult_1/zreg_reg[479]  ( .D(mod_mult_o[479]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][479] ) );
  DFF \modmult_1/zreg_reg[478]  ( .D(mod_mult_o[478]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][478] ) );
  DFF \modmult_1/zreg_reg[477]  ( .D(mod_mult_o[477]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][477] ) );
  DFF \modmult_1/zreg_reg[476]  ( .D(mod_mult_o[476]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][476] ) );
  DFF \modmult_1/zreg_reg[475]  ( .D(mod_mult_o[475]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][475] ) );
  DFF \modmult_1/zreg_reg[474]  ( .D(mod_mult_o[474]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][474] ) );
  DFF \modmult_1/zreg_reg[473]  ( .D(mod_mult_o[473]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][473] ) );
  DFF \modmult_1/zreg_reg[472]  ( .D(mod_mult_o[472]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][472] ) );
  DFF \modmult_1/zreg_reg[471]  ( .D(mod_mult_o[471]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][471] ) );
  DFF \modmult_1/zreg_reg[470]  ( .D(mod_mult_o[470]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][470] ) );
  DFF \modmult_1/zreg_reg[469]  ( .D(mod_mult_o[469]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][469] ) );
  DFF \modmult_1/zreg_reg[468]  ( .D(mod_mult_o[468]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][468] ) );
  DFF \modmult_1/zreg_reg[467]  ( .D(mod_mult_o[467]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][467] ) );
  DFF \modmult_1/zreg_reg[466]  ( .D(mod_mult_o[466]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][466] ) );
  DFF \modmult_1/zreg_reg[465]  ( .D(mod_mult_o[465]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][465] ) );
  DFF \modmult_1/zreg_reg[464]  ( .D(mod_mult_o[464]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][464] ) );
  DFF \modmult_1/zreg_reg[463]  ( .D(mod_mult_o[463]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][463] ) );
  DFF \modmult_1/zreg_reg[462]  ( .D(mod_mult_o[462]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][462] ) );
  DFF \modmult_1/zreg_reg[461]  ( .D(mod_mult_o[461]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][461] ) );
  DFF \modmult_1/zreg_reg[460]  ( .D(mod_mult_o[460]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][460] ) );
  DFF \modmult_1/zreg_reg[459]  ( .D(mod_mult_o[459]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][459] ) );
  DFF \modmult_1/zreg_reg[458]  ( .D(mod_mult_o[458]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][458] ) );
  DFF \modmult_1/zreg_reg[457]  ( .D(mod_mult_o[457]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][457] ) );
  DFF \modmult_1/zreg_reg[456]  ( .D(mod_mult_o[456]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][456] ) );
  DFF \modmult_1/zreg_reg[455]  ( .D(mod_mult_o[455]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][455] ) );
  DFF \modmult_1/zreg_reg[454]  ( .D(mod_mult_o[454]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][454] ) );
  DFF \modmult_1/zreg_reg[453]  ( .D(mod_mult_o[453]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][453] ) );
  DFF \modmult_1/zreg_reg[452]  ( .D(mod_mult_o[452]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][452] ) );
  DFF \modmult_1/zreg_reg[451]  ( .D(mod_mult_o[451]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][451] ) );
  DFF \modmult_1/zreg_reg[450]  ( .D(mod_mult_o[450]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][450] ) );
  DFF \modmult_1/zreg_reg[449]  ( .D(mod_mult_o[449]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][449] ) );
  DFF \modmult_1/zreg_reg[448]  ( .D(mod_mult_o[448]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][448] ) );
  DFF \modmult_1/zreg_reg[447]  ( .D(mod_mult_o[447]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][447] ) );
  DFF \modmult_1/zreg_reg[446]  ( .D(mod_mult_o[446]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][446] ) );
  DFF \modmult_1/zreg_reg[445]  ( .D(mod_mult_o[445]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][445] ) );
  DFF \modmult_1/zreg_reg[444]  ( .D(mod_mult_o[444]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][444] ) );
  DFF \modmult_1/zreg_reg[443]  ( .D(mod_mult_o[443]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][443] ) );
  DFF \modmult_1/zreg_reg[442]  ( .D(mod_mult_o[442]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][442] ) );
  DFF \modmult_1/zreg_reg[441]  ( .D(mod_mult_o[441]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][441] ) );
  DFF \modmult_1/zreg_reg[440]  ( .D(mod_mult_o[440]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][440] ) );
  DFF \modmult_1/zreg_reg[439]  ( .D(mod_mult_o[439]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][439] ) );
  DFF \modmult_1/zreg_reg[438]  ( .D(mod_mult_o[438]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][438] ) );
  DFF \modmult_1/zreg_reg[437]  ( .D(mod_mult_o[437]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][437] ) );
  DFF \modmult_1/zreg_reg[436]  ( .D(mod_mult_o[436]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][436] ) );
  DFF \modmult_1/zreg_reg[435]  ( .D(mod_mult_o[435]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][435] ) );
  DFF \modmult_1/zreg_reg[434]  ( .D(mod_mult_o[434]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][434] ) );
  DFF \modmult_1/zreg_reg[433]  ( .D(mod_mult_o[433]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][433] ) );
  DFF \modmult_1/zreg_reg[432]  ( .D(mod_mult_o[432]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][432] ) );
  DFF \modmult_1/zreg_reg[431]  ( .D(mod_mult_o[431]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][431] ) );
  DFF \modmult_1/zreg_reg[430]  ( .D(mod_mult_o[430]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][430] ) );
  DFF \modmult_1/zreg_reg[429]  ( .D(mod_mult_o[429]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][429] ) );
  DFF \modmult_1/zreg_reg[428]  ( .D(mod_mult_o[428]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][428] ) );
  DFF \modmult_1/zreg_reg[427]  ( .D(mod_mult_o[427]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][427] ) );
  DFF \modmult_1/zreg_reg[426]  ( .D(mod_mult_o[426]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][426] ) );
  DFF \modmult_1/zreg_reg[425]  ( .D(mod_mult_o[425]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][425] ) );
  DFF \modmult_1/zreg_reg[424]  ( .D(mod_mult_o[424]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][424] ) );
  DFF \modmult_1/zreg_reg[423]  ( .D(mod_mult_o[423]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][423] ) );
  DFF \modmult_1/zreg_reg[422]  ( .D(mod_mult_o[422]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][422] ) );
  DFF \modmult_1/zreg_reg[421]  ( .D(mod_mult_o[421]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][421] ) );
  DFF \modmult_1/zreg_reg[420]  ( .D(mod_mult_o[420]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][420] ) );
  DFF \modmult_1/zreg_reg[419]  ( .D(mod_mult_o[419]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][419] ) );
  DFF \modmult_1/zreg_reg[418]  ( .D(mod_mult_o[418]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][418] ) );
  DFF \modmult_1/zreg_reg[417]  ( .D(mod_mult_o[417]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][417] ) );
  DFF \modmult_1/zreg_reg[416]  ( .D(mod_mult_o[416]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][416] ) );
  DFF \modmult_1/zreg_reg[415]  ( .D(mod_mult_o[415]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][415] ) );
  DFF \modmult_1/zreg_reg[414]  ( .D(mod_mult_o[414]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][414] ) );
  DFF \modmult_1/zreg_reg[413]  ( .D(mod_mult_o[413]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][413] ) );
  DFF \modmult_1/zreg_reg[412]  ( .D(mod_mult_o[412]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][412] ) );
  DFF \modmult_1/zreg_reg[411]  ( .D(mod_mult_o[411]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][411] ) );
  DFF \modmult_1/zreg_reg[410]  ( .D(mod_mult_o[410]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][410] ) );
  DFF \modmult_1/zreg_reg[409]  ( .D(mod_mult_o[409]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][409] ) );
  DFF \modmult_1/zreg_reg[408]  ( .D(mod_mult_o[408]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][408] ) );
  DFF \modmult_1/zreg_reg[407]  ( .D(mod_mult_o[407]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][407] ) );
  DFF \modmult_1/zreg_reg[406]  ( .D(mod_mult_o[406]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][406] ) );
  DFF \modmult_1/zreg_reg[405]  ( .D(mod_mult_o[405]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][405] ) );
  DFF \modmult_1/zreg_reg[404]  ( .D(mod_mult_o[404]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][404] ) );
  DFF \modmult_1/zreg_reg[403]  ( .D(mod_mult_o[403]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][403] ) );
  DFF \modmult_1/zreg_reg[402]  ( .D(mod_mult_o[402]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][402] ) );
  DFF \modmult_1/zreg_reg[401]  ( .D(mod_mult_o[401]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][401] ) );
  DFF \modmult_1/zreg_reg[400]  ( .D(mod_mult_o[400]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][400] ) );
  DFF \modmult_1/zreg_reg[399]  ( .D(mod_mult_o[399]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][399] ) );
  DFF \modmult_1/zreg_reg[398]  ( .D(mod_mult_o[398]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][398] ) );
  DFF \modmult_1/zreg_reg[397]  ( .D(mod_mult_o[397]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][397] ) );
  DFF \modmult_1/zreg_reg[396]  ( .D(mod_mult_o[396]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][396] ) );
  DFF \modmult_1/zreg_reg[395]  ( .D(mod_mult_o[395]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][395] ) );
  DFF \modmult_1/zreg_reg[394]  ( .D(mod_mult_o[394]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][394] ) );
  DFF \modmult_1/zreg_reg[393]  ( .D(mod_mult_o[393]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][393] ) );
  DFF \modmult_1/zreg_reg[392]  ( .D(mod_mult_o[392]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][392] ) );
  DFF \modmult_1/zreg_reg[391]  ( .D(mod_mult_o[391]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][391] ) );
  DFF \modmult_1/zreg_reg[390]  ( .D(mod_mult_o[390]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][390] ) );
  DFF \modmult_1/zreg_reg[389]  ( .D(mod_mult_o[389]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][389] ) );
  DFF \modmult_1/zreg_reg[388]  ( .D(mod_mult_o[388]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][388] ) );
  DFF \modmult_1/zreg_reg[387]  ( .D(mod_mult_o[387]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][387] ) );
  DFF \modmult_1/zreg_reg[386]  ( .D(mod_mult_o[386]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][386] ) );
  DFF \modmult_1/zreg_reg[385]  ( .D(mod_mult_o[385]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][385] ) );
  DFF \modmult_1/zreg_reg[384]  ( .D(mod_mult_o[384]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][384] ) );
  DFF \modmult_1/zreg_reg[383]  ( .D(mod_mult_o[383]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][383] ) );
  DFF \modmult_1/zreg_reg[382]  ( .D(mod_mult_o[382]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][382] ) );
  DFF \modmult_1/zreg_reg[381]  ( .D(mod_mult_o[381]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][381] ) );
  DFF \modmult_1/zreg_reg[380]  ( .D(mod_mult_o[380]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][380] ) );
  DFF \modmult_1/zreg_reg[379]  ( .D(mod_mult_o[379]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][379] ) );
  DFF \modmult_1/zreg_reg[378]  ( .D(mod_mult_o[378]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][378] ) );
  DFF \modmult_1/zreg_reg[377]  ( .D(mod_mult_o[377]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][377] ) );
  DFF \modmult_1/zreg_reg[376]  ( .D(mod_mult_o[376]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][376] ) );
  DFF \modmult_1/zreg_reg[375]  ( .D(mod_mult_o[375]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][375] ) );
  DFF \modmult_1/zreg_reg[374]  ( .D(mod_mult_o[374]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][374] ) );
  DFF \modmult_1/zreg_reg[373]  ( .D(mod_mult_o[373]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][373] ) );
  DFF \modmult_1/zreg_reg[372]  ( .D(mod_mult_o[372]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][372] ) );
  DFF \modmult_1/zreg_reg[371]  ( .D(mod_mult_o[371]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][371] ) );
  DFF \modmult_1/zreg_reg[370]  ( .D(mod_mult_o[370]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][370] ) );
  DFF \modmult_1/zreg_reg[369]  ( .D(mod_mult_o[369]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][369] ) );
  DFF \modmult_1/zreg_reg[368]  ( .D(mod_mult_o[368]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][368] ) );
  DFF \modmult_1/zreg_reg[367]  ( .D(mod_mult_o[367]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][367] ) );
  DFF \modmult_1/zreg_reg[366]  ( .D(mod_mult_o[366]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][366] ) );
  DFF \modmult_1/zreg_reg[365]  ( .D(mod_mult_o[365]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][365] ) );
  DFF \modmult_1/zreg_reg[364]  ( .D(mod_mult_o[364]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][364] ) );
  DFF \modmult_1/zreg_reg[363]  ( .D(mod_mult_o[363]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][363] ) );
  DFF \modmult_1/zreg_reg[362]  ( .D(mod_mult_o[362]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][362] ) );
  DFF \modmult_1/zreg_reg[361]  ( .D(mod_mult_o[361]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][361] ) );
  DFF \modmult_1/zreg_reg[360]  ( .D(mod_mult_o[360]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][360] ) );
  DFF \modmult_1/zreg_reg[359]  ( .D(mod_mult_o[359]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][359] ) );
  DFF \modmult_1/zreg_reg[358]  ( .D(mod_mult_o[358]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][358] ) );
  DFF \modmult_1/zreg_reg[357]  ( .D(mod_mult_o[357]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][357] ) );
  DFF \modmult_1/zreg_reg[356]  ( .D(mod_mult_o[356]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][356] ) );
  DFF \modmult_1/zreg_reg[355]  ( .D(mod_mult_o[355]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][355] ) );
  DFF \modmult_1/zreg_reg[354]  ( .D(mod_mult_o[354]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][354] ) );
  DFF \modmult_1/zreg_reg[353]  ( .D(mod_mult_o[353]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][353] ) );
  DFF \modmult_1/zreg_reg[352]  ( .D(mod_mult_o[352]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][352] ) );
  DFF \modmult_1/zreg_reg[351]  ( .D(mod_mult_o[351]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][351] ) );
  DFF \modmult_1/zreg_reg[350]  ( .D(mod_mult_o[350]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][350] ) );
  DFF \modmult_1/zreg_reg[349]  ( .D(mod_mult_o[349]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][349] ) );
  DFF \modmult_1/zreg_reg[348]  ( .D(mod_mult_o[348]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][348] ) );
  DFF \modmult_1/zreg_reg[347]  ( .D(mod_mult_o[347]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][347] ) );
  DFF \modmult_1/zreg_reg[346]  ( .D(mod_mult_o[346]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][346] ) );
  DFF \modmult_1/zreg_reg[345]  ( .D(mod_mult_o[345]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][345] ) );
  DFF \modmult_1/zreg_reg[344]  ( .D(mod_mult_o[344]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][344] ) );
  DFF \modmult_1/zreg_reg[343]  ( .D(mod_mult_o[343]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][343] ) );
  DFF \modmult_1/zreg_reg[342]  ( .D(mod_mult_o[342]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][342] ) );
  DFF \modmult_1/zreg_reg[341]  ( .D(mod_mult_o[341]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][341] ) );
  DFF \modmult_1/zreg_reg[340]  ( .D(mod_mult_o[340]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][340] ) );
  DFF \modmult_1/zreg_reg[339]  ( .D(mod_mult_o[339]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][339] ) );
  DFF \modmult_1/zreg_reg[338]  ( .D(mod_mult_o[338]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][338] ) );
  DFF \modmult_1/zreg_reg[337]  ( .D(mod_mult_o[337]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][337] ) );
  DFF \modmult_1/zreg_reg[336]  ( .D(mod_mult_o[336]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][336] ) );
  DFF \modmult_1/zreg_reg[335]  ( .D(mod_mult_o[335]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][335] ) );
  DFF \modmult_1/zreg_reg[334]  ( .D(mod_mult_o[334]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][334] ) );
  DFF \modmult_1/zreg_reg[333]  ( .D(mod_mult_o[333]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][333] ) );
  DFF \modmult_1/zreg_reg[332]  ( .D(mod_mult_o[332]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][332] ) );
  DFF \modmult_1/zreg_reg[331]  ( .D(mod_mult_o[331]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][331] ) );
  DFF \modmult_1/zreg_reg[330]  ( .D(mod_mult_o[330]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][330] ) );
  DFF \modmult_1/zreg_reg[329]  ( .D(mod_mult_o[329]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][329] ) );
  DFF \modmult_1/zreg_reg[328]  ( .D(mod_mult_o[328]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][328] ) );
  DFF \modmult_1/zreg_reg[327]  ( .D(mod_mult_o[327]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][327] ) );
  DFF \modmult_1/zreg_reg[326]  ( .D(mod_mult_o[326]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][326] ) );
  DFF \modmult_1/zreg_reg[325]  ( .D(mod_mult_o[325]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][325] ) );
  DFF \modmult_1/zreg_reg[324]  ( .D(mod_mult_o[324]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][324] ) );
  DFF \modmult_1/zreg_reg[323]  ( .D(mod_mult_o[323]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][323] ) );
  DFF \modmult_1/zreg_reg[322]  ( .D(mod_mult_o[322]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][322] ) );
  DFF \modmult_1/zreg_reg[321]  ( .D(mod_mult_o[321]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][321] ) );
  DFF \modmult_1/zreg_reg[320]  ( .D(mod_mult_o[320]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][320] ) );
  DFF \modmult_1/zreg_reg[319]  ( .D(mod_mult_o[319]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][319] ) );
  DFF \modmult_1/zreg_reg[318]  ( .D(mod_mult_o[318]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][318] ) );
  DFF \modmult_1/zreg_reg[317]  ( .D(mod_mult_o[317]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][317] ) );
  DFF \modmult_1/zreg_reg[316]  ( .D(mod_mult_o[316]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][316] ) );
  DFF \modmult_1/zreg_reg[315]  ( .D(mod_mult_o[315]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][315] ) );
  DFF \modmult_1/zreg_reg[314]  ( .D(mod_mult_o[314]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][314] ) );
  DFF \modmult_1/zreg_reg[313]  ( .D(mod_mult_o[313]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][313] ) );
  DFF \modmult_1/zreg_reg[312]  ( .D(mod_mult_o[312]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][312] ) );
  DFF \modmult_1/zreg_reg[311]  ( .D(mod_mult_o[311]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][311] ) );
  DFF \modmult_1/zreg_reg[310]  ( .D(mod_mult_o[310]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][310] ) );
  DFF \modmult_1/zreg_reg[309]  ( .D(mod_mult_o[309]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][309] ) );
  DFF \modmult_1/zreg_reg[308]  ( .D(mod_mult_o[308]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][308] ) );
  DFF \modmult_1/zreg_reg[307]  ( .D(mod_mult_o[307]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][307] ) );
  DFF \modmult_1/zreg_reg[306]  ( .D(mod_mult_o[306]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][306] ) );
  DFF \modmult_1/zreg_reg[305]  ( .D(mod_mult_o[305]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][305] ) );
  DFF \modmult_1/zreg_reg[304]  ( .D(mod_mult_o[304]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][304] ) );
  DFF \modmult_1/zreg_reg[303]  ( .D(mod_mult_o[303]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][303] ) );
  DFF \modmult_1/zreg_reg[302]  ( .D(mod_mult_o[302]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][302] ) );
  DFF \modmult_1/zreg_reg[301]  ( .D(mod_mult_o[301]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][301] ) );
  DFF \modmult_1/zreg_reg[300]  ( .D(mod_mult_o[300]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][300] ) );
  DFF \modmult_1/zreg_reg[299]  ( .D(mod_mult_o[299]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][299] ) );
  DFF \modmult_1/zreg_reg[298]  ( .D(mod_mult_o[298]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][298] ) );
  DFF \modmult_1/zreg_reg[297]  ( .D(mod_mult_o[297]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][297] ) );
  DFF \modmult_1/zreg_reg[296]  ( .D(mod_mult_o[296]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][296] ) );
  DFF \modmult_1/zreg_reg[295]  ( .D(mod_mult_o[295]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][295] ) );
  DFF \modmult_1/zreg_reg[294]  ( .D(mod_mult_o[294]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][294] ) );
  DFF \modmult_1/zreg_reg[293]  ( .D(mod_mult_o[293]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][293] ) );
  DFF \modmult_1/zreg_reg[292]  ( .D(mod_mult_o[292]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][292] ) );
  DFF \modmult_1/zreg_reg[291]  ( .D(mod_mult_o[291]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][291] ) );
  DFF \modmult_1/zreg_reg[290]  ( .D(mod_mult_o[290]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][290] ) );
  DFF \modmult_1/zreg_reg[289]  ( .D(mod_mult_o[289]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][289] ) );
  DFF \modmult_1/zreg_reg[288]  ( .D(mod_mult_o[288]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][288] ) );
  DFF \modmult_1/zreg_reg[287]  ( .D(mod_mult_o[287]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][287] ) );
  DFF \modmult_1/zreg_reg[286]  ( .D(mod_mult_o[286]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][286] ) );
  DFF \modmult_1/zreg_reg[285]  ( .D(mod_mult_o[285]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][285] ) );
  DFF \modmult_1/zreg_reg[284]  ( .D(mod_mult_o[284]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][284] ) );
  DFF \modmult_1/zreg_reg[283]  ( .D(mod_mult_o[283]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][283] ) );
  DFF \modmult_1/zreg_reg[282]  ( .D(mod_mult_o[282]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][282] ) );
  DFF \modmult_1/zreg_reg[281]  ( .D(mod_mult_o[281]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][281] ) );
  DFF \modmult_1/zreg_reg[280]  ( .D(mod_mult_o[280]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][280] ) );
  DFF \modmult_1/zreg_reg[279]  ( .D(mod_mult_o[279]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][279] ) );
  DFF \modmult_1/zreg_reg[278]  ( .D(mod_mult_o[278]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][278] ) );
  DFF \modmult_1/zreg_reg[277]  ( .D(mod_mult_o[277]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][277] ) );
  DFF \modmult_1/zreg_reg[276]  ( .D(mod_mult_o[276]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][276] ) );
  DFF \modmult_1/zreg_reg[275]  ( .D(mod_mult_o[275]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][275] ) );
  DFF \modmult_1/zreg_reg[274]  ( .D(mod_mult_o[274]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][274] ) );
  DFF \modmult_1/zreg_reg[273]  ( .D(mod_mult_o[273]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][273] ) );
  DFF \modmult_1/zreg_reg[272]  ( .D(mod_mult_o[272]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][272] ) );
  DFF \modmult_1/zreg_reg[271]  ( .D(mod_mult_o[271]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][271] ) );
  DFF \modmult_1/zreg_reg[270]  ( .D(mod_mult_o[270]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][270] ) );
  DFF \modmult_1/zreg_reg[269]  ( .D(mod_mult_o[269]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][269] ) );
  DFF \modmult_1/zreg_reg[268]  ( .D(mod_mult_o[268]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][268] ) );
  DFF \modmult_1/zreg_reg[267]  ( .D(mod_mult_o[267]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][267] ) );
  DFF \modmult_1/zreg_reg[266]  ( .D(mod_mult_o[266]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][266] ) );
  DFF \modmult_1/zreg_reg[265]  ( .D(mod_mult_o[265]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][265] ) );
  DFF \modmult_1/zreg_reg[264]  ( .D(mod_mult_o[264]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][264] ) );
  DFF \modmult_1/zreg_reg[263]  ( .D(mod_mult_o[263]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][263] ) );
  DFF \modmult_1/zreg_reg[262]  ( .D(mod_mult_o[262]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][262] ) );
  DFF \modmult_1/zreg_reg[261]  ( .D(mod_mult_o[261]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][261] ) );
  DFF \modmult_1/zreg_reg[260]  ( .D(mod_mult_o[260]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][260] ) );
  DFF \modmult_1/zreg_reg[259]  ( .D(mod_mult_o[259]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][259] ) );
  DFF \modmult_1/zreg_reg[258]  ( .D(mod_mult_o[258]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][258] ) );
  DFF \modmult_1/zreg_reg[257]  ( .D(mod_mult_o[257]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][257] ) );
  DFF \modmult_1/zreg_reg[256]  ( .D(mod_mult_o[256]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][256] ) );
  DFF \modmult_1/zreg_reg[255]  ( .D(mod_mult_o[255]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][255] ) );
  DFF \modmult_1/zreg_reg[254]  ( .D(mod_mult_o[254]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][254] ) );
  DFF \modmult_1/zreg_reg[253]  ( .D(mod_mult_o[253]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][253] ) );
  DFF \modmult_1/zreg_reg[252]  ( .D(mod_mult_o[252]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][252] ) );
  DFF \modmult_1/zreg_reg[251]  ( .D(mod_mult_o[251]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][251] ) );
  DFF \modmult_1/zreg_reg[250]  ( .D(mod_mult_o[250]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][250] ) );
  DFF \modmult_1/zreg_reg[249]  ( .D(mod_mult_o[249]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][249] ) );
  DFF \modmult_1/zreg_reg[248]  ( .D(mod_mult_o[248]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][248] ) );
  DFF \modmult_1/zreg_reg[247]  ( .D(mod_mult_o[247]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][247] ) );
  DFF \modmult_1/zreg_reg[246]  ( .D(mod_mult_o[246]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][246] ) );
  DFF \modmult_1/zreg_reg[245]  ( .D(mod_mult_o[245]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][245] ) );
  DFF \modmult_1/zreg_reg[244]  ( .D(mod_mult_o[244]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][244] ) );
  DFF \modmult_1/zreg_reg[243]  ( .D(mod_mult_o[243]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][243] ) );
  DFF \modmult_1/zreg_reg[242]  ( .D(mod_mult_o[242]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][242] ) );
  DFF \modmult_1/zreg_reg[241]  ( .D(mod_mult_o[241]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][241] ) );
  DFF \modmult_1/zreg_reg[240]  ( .D(mod_mult_o[240]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][240] ) );
  DFF \modmult_1/zreg_reg[239]  ( .D(mod_mult_o[239]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][239] ) );
  DFF \modmult_1/zreg_reg[238]  ( .D(mod_mult_o[238]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][238] ) );
  DFF \modmult_1/zreg_reg[237]  ( .D(mod_mult_o[237]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][237] ) );
  DFF \modmult_1/zreg_reg[236]  ( .D(mod_mult_o[236]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][236] ) );
  DFF \modmult_1/zreg_reg[235]  ( .D(mod_mult_o[235]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][235] ) );
  DFF \modmult_1/zreg_reg[234]  ( .D(mod_mult_o[234]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][234] ) );
  DFF \modmult_1/zreg_reg[233]  ( .D(mod_mult_o[233]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][233] ) );
  DFF \modmult_1/zreg_reg[232]  ( .D(mod_mult_o[232]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][232] ) );
  DFF \modmult_1/zreg_reg[231]  ( .D(mod_mult_o[231]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][231] ) );
  DFF \modmult_1/zreg_reg[230]  ( .D(mod_mult_o[230]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][230] ) );
  DFF \modmult_1/zreg_reg[229]  ( .D(mod_mult_o[229]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][229] ) );
  DFF \modmult_1/zreg_reg[228]  ( .D(mod_mult_o[228]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][228] ) );
  DFF \modmult_1/zreg_reg[227]  ( .D(mod_mult_o[227]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][227] ) );
  DFF \modmult_1/zreg_reg[226]  ( .D(mod_mult_o[226]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][226] ) );
  DFF \modmult_1/zreg_reg[225]  ( .D(mod_mult_o[225]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][225] ) );
  DFF \modmult_1/zreg_reg[224]  ( .D(mod_mult_o[224]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][224] ) );
  DFF \modmult_1/zreg_reg[223]  ( .D(mod_mult_o[223]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][223] ) );
  DFF \modmult_1/zreg_reg[222]  ( .D(mod_mult_o[222]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][222] ) );
  DFF \modmult_1/zreg_reg[221]  ( .D(mod_mult_o[221]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][221] ) );
  DFF \modmult_1/zreg_reg[220]  ( .D(mod_mult_o[220]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][220] ) );
  DFF \modmult_1/zreg_reg[219]  ( .D(mod_mult_o[219]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][219] ) );
  DFF \modmult_1/zreg_reg[218]  ( .D(mod_mult_o[218]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][218] ) );
  DFF \modmult_1/zreg_reg[217]  ( .D(mod_mult_o[217]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][217] ) );
  DFF \modmult_1/zreg_reg[216]  ( .D(mod_mult_o[216]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][216] ) );
  DFF \modmult_1/zreg_reg[215]  ( .D(mod_mult_o[215]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][215] ) );
  DFF \modmult_1/zreg_reg[214]  ( .D(mod_mult_o[214]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][214] ) );
  DFF \modmult_1/zreg_reg[213]  ( .D(mod_mult_o[213]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][213] ) );
  DFF \modmult_1/zreg_reg[212]  ( .D(mod_mult_o[212]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][212] ) );
  DFF \modmult_1/zreg_reg[211]  ( .D(mod_mult_o[211]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][211] ) );
  DFF \modmult_1/zreg_reg[210]  ( .D(mod_mult_o[210]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][210] ) );
  DFF \modmult_1/zreg_reg[209]  ( .D(mod_mult_o[209]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][209] ) );
  DFF \modmult_1/zreg_reg[208]  ( .D(mod_mult_o[208]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][208] ) );
  DFF \modmult_1/zreg_reg[207]  ( .D(mod_mult_o[207]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][207] ) );
  DFF \modmult_1/zreg_reg[206]  ( .D(mod_mult_o[206]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][206] ) );
  DFF \modmult_1/zreg_reg[205]  ( .D(mod_mult_o[205]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][205] ) );
  DFF \modmult_1/zreg_reg[204]  ( .D(mod_mult_o[204]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][204] ) );
  DFF \modmult_1/zreg_reg[203]  ( .D(mod_mult_o[203]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][203] ) );
  DFF \modmult_1/zreg_reg[202]  ( .D(mod_mult_o[202]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][202] ) );
  DFF \modmult_1/zreg_reg[201]  ( .D(mod_mult_o[201]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][201] ) );
  DFF \modmult_1/zreg_reg[200]  ( .D(mod_mult_o[200]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][200] ) );
  DFF \modmult_1/zreg_reg[199]  ( .D(mod_mult_o[199]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][199] ) );
  DFF \modmult_1/zreg_reg[198]  ( .D(mod_mult_o[198]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][198] ) );
  DFF \modmult_1/zreg_reg[197]  ( .D(mod_mult_o[197]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][197] ) );
  DFF \modmult_1/zreg_reg[196]  ( .D(mod_mult_o[196]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][196] ) );
  DFF \modmult_1/zreg_reg[195]  ( .D(mod_mult_o[195]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][195] ) );
  DFF \modmult_1/zreg_reg[194]  ( .D(mod_mult_o[194]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][194] ) );
  DFF \modmult_1/zreg_reg[193]  ( .D(mod_mult_o[193]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][193] ) );
  DFF \modmult_1/zreg_reg[192]  ( .D(mod_mult_o[192]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][192] ) );
  DFF \modmult_1/zreg_reg[191]  ( .D(mod_mult_o[191]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][191] ) );
  DFF \modmult_1/zreg_reg[190]  ( .D(mod_mult_o[190]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][190] ) );
  DFF \modmult_1/zreg_reg[189]  ( .D(mod_mult_o[189]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][189] ) );
  DFF \modmult_1/zreg_reg[188]  ( .D(mod_mult_o[188]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][188] ) );
  DFF \modmult_1/zreg_reg[187]  ( .D(mod_mult_o[187]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][187] ) );
  DFF \modmult_1/zreg_reg[186]  ( .D(mod_mult_o[186]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][186] ) );
  DFF \modmult_1/zreg_reg[185]  ( .D(mod_mult_o[185]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][185] ) );
  DFF \modmult_1/zreg_reg[184]  ( .D(mod_mult_o[184]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][184] ) );
  DFF \modmult_1/zreg_reg[183]  ( .D(mod_mult_o[183]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][183] ) );
  DFF \modmult_1/zreg_reg[182]  ( .D(mod_mult_o[182]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][182] ) );
  DFF \modmult_1/zreg_reg[181]  ( .D(mod_mult_o[181]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][181] ) );
  DFF \modmult_1/zreg_reg[180]  ( .D(mod_mult_o[180]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][180] ) );
  DFF \modmult_1/zreg_reg[179]  ( .D(mod_mult_o[179]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][179] ) );
  DFF \modmult_1/zreg_reg[178]  ( .D(mod_mult_o[178]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][178] ) );
  DFF \modmult_1/zreg_reg[177]  ( .D(mod_mult_o[177]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][177] ) );
  DFF \modmult_1/zreg_reg[176]  ( .D(mod_mult_o[176]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][176] ) );
  DFF \modmult_1/zreg_reg[175]  ( .D(mod_mult_o[175]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][175] ) );
  DFF \modmult_1/zreg_reg[174]  ( .D(mod_mult_o[174]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][174] ) );
  DFF \modmult_1/zreg_reg[173]  ( .D(mod_mult_o[173]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][173] ) );
  DFF \modmult_1/zreg_reg[172]  ( .D(mod_mult_o[172]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][172] ) );
  DFF \modmult_1/zreg_reg[171]  ( .D(mod_mult_o[171]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][171] ) );
  DFF \modmult_1/zreg_reg[170]  ( .D(mod_mult_o[170]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][170] ) );
  DFF \modmult_1/zreg_reg[169]  ( .D(mod_mult_o[169]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][169] ) );
  DFF \modmult_1/zreg_reg[168]  ( .D(mod_mult_o[168]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][168] ) );
  DFF \modmult_1/zreg_reg[167]  ( .D(mod_mult_o[167]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][167] ) );
  DFF \modmult_1/zreg_reg[166]  ( .D(mod_mult_o[166]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][166] ) );
  DFF \modmult_1/zreg_reg[165]  ( .D(mod_mult_o[165]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][165] ) );
  DFF \modmult_1/zreg_reg[164]  ( .D(mod_mult_o[164]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][164] ) );
  DFF \modmult_1/zreg_reg[163]  ( .D(mod_mult_o[163]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][163] ) );
  DFF \modmult_1/zreg_reg[162]  ( .D(mod_mult_o[162]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][162] ) );
  DFF \modmult_1/zreg_reg[161]  ( .D(mod_mult_o[161]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][161] ) );
  DFF \modmult_1/zreg_reg[160]  ( .D(mod_mult_o[160]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][160] ) );
  DFF \modmult_1/zreg_reg[159]  ( .D(mod_mult_o[159]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][159] ) );
  DFF \modmult_1/zreg_reg[158]  ( .D(mod_mult_o[158]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][158] ) );
  DFF \modmult_1/zreg_reg[157]  ( .D(mod_mult_o[157]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][157] ) );
  DFF \modmult_1/zreg_reg[156]  ( .D(mod_mult_o[156]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][156] ) );
  DFF \modmult_1/zreg_reg[155]  ( .D(mod_mult_o[155]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][155] ) );
  DFF \modmult_1/zreg_reg[154]  ( .D(mod_mult_o[154]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][154] ) );
  DFF \modmult_1/zreg_reg[153]  ( .D(mod_mult_o[153]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][153] ) );
  DFF \modmult_1/zreg_reg[152]  ( .D(mod_mult_o[152]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][152] ) );
  DFF \modmult_1/zreg_reg[151]  ( .D(mod_mult_o[151]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][151] ) );
  DFF \modmult_1/zreg_reg[150]  ( .D(mod_mult_o[150]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][150] ) );
  DFF \modmult_1/zreg_reg[149]  ( .D(mod_mult_o[149]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][149] ) );
  DFF \modmult_1/zreg_reg[148]  ( .D(mod_mult_o[148]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][148] ) );
  DFF \modmult_1/zreg_reg[147]  ( .D(mod_mult_o[147]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][147] ) );
  DFF \modmult_1/zreg_reg[146]  ( .D(mod_mult_o[146]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][146] ) );
  DFF \modmult_1/zreg_reg[145]  ( .D(mod_mult_o[145]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][145] ) );
  DFF \modmult_1/zreg_reg[144]  ( .D(mod_mult_o[144]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][144] ) );
  DFF \modmult_1/zreg_reg[143]  ( .D(mod_mult_o[143]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][143] ) );
  DFF \modmult_1/zreg_reg[142]  ( .D(mod_mult_o[142]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][142] ) );
  DFF \modmult_1/zreg_reg[141]  ( .D(mod_mult_o[141]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][141] ) );
  DFF \modmult_1/zreg_reg[140]  ( .D(mod_mult_o[140]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][140] ) );
  DFF \modmult_1/zreg_reg[139]  ( .D(mod_mult_o[139]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][139] ) );
  DFF \modmult_1/zreg_reg[138]  ( .D(mod_mult_o[138]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][138] ) );
  DFF \modmult_1/zreg_reg[137]  ( .D(mod_mult_o[137]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][137] ) );
  DFF \modmult_1/zreg_reg[136]  ( .D(mod_mult_o[136]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][136] ) );
  DFF \modmult_1/zreg_reg[135]  ( .D(mod_mult_o[135]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][135] ) );
  DFF \modmult_1/zreg_reg[134]  ( .D(mod_mult_o[134]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][134] ) );
  DFF \modmult_1/zreg_reg[133]  ( .D(mod_mult_o[133]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][133] ) );
  DFF \modmult_1/zreg_reg[132]  ( .D(mod_mult_o[132]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][132] ) );
  DFF \modmult_1/zreg_reg[131]  ( .D(mod_mult_o[131]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][131] ) );
  DFF \modmult_1/zreg_reg[130]  ( .D(mod_mult_o[130]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][130] ) );
  DFF \modmult_1/zreg_reg[129]  ( .D(mod_mult_o[129]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][129] ) );
  DFF \modmult_1/zreg_reg[128]  ( .D(mod_mult_o[128]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][128] ) );
  DFF \modmult_1/zreg_reg[127]  ( .D(mod_mult_o[127]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][127] ) );
  DFF \modmult_1/zreg_reg[126]  ( .D(mod_mult_o[126]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][126] ) );
  DFF \modmult_1/zreg_reg[125]  ( .D(mod_mult_o[125]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][125] ) );
  DFF \modmult_1/zreg_reg[124]  ( .D(mod_mult_o[124]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][124] ) );
  DFF \modmult_1/zreg_reg[123]  ( .D(mod_mult_o[123]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][123] ) );
  DFF \modmult_1/zreg_reg[122]  ( .D(mod_mult_o[122]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][122] ) );
  DFF \modmult_1/zreg_reg[121]  ( .D(mod_mult_o[121]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][121] ) );
  DFF \modmult_1/zreg_reg[120]  ( .D(mod_mult_o[120]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][120] ) );
  DFF \modmult_1/zreg_reg[119]  ( .D(mod_mult_o[119]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][119] ) );
  DFF \modmult_1/zreg_reg[118]  ( .D(mod_mult_o[118]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][118] ) );
  DFF \modmult_1/zreg_reg[117]  ( .D(mod_mult_o[117]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][117] ) );
  DFF \modmult_1/zreg_reg[116]  ( .D(mod_mult_o[116]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][116] ) );
  DFF \modmult_1/zreg_reg[115]  ( .D(mod_mult_o[115]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][115] ) );
  DFF \modmult_1/zreg_reg[114]  ( .D(mod_mult_o[114]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][114] ) );
  DFF \modmult_1/zreg_reg[113]  ( .D(mod_mult_o[113]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][113] ) );
  DFF \modmult_1/zreg_reg[112]  ( .D(mod_mult_o[112]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][112] ) );
  DFF \modmult_1/zreg_reg[111]  ( .D(mod_mult_o[111]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][111] ) );
  DFF \modmult_1/zreg_reg[110]  ( .D(mod_mult_o[110]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][110] ) );
  DFF \modmult_1/zreg_reg[109]  ( .D(mod_mult_o[109]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][109] ) );
  DFF \modmult_1/zreg_reg[108]  ( .D(mod_mult_o[108]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][108] ) );
  DFF \modmult_1/zreg_reg[107]  ( .D(mod_mult_o[107]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][107] ) );
  DFF \modmult_1/zreg_reg[106]  ( .D(mod_mult_o[106]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][106] ) );
  DFF \modmult_1/zreg_reg[105]  ( .D(mod_mult_o[105]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][105] ) );
  DFF \modmult_1/zreg_reg[104]  ( .D(mod_mult_o[104]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][104] ) );
  DFF \modmult_1/zreg_reg[103]  ( .D(mod_mult_o[103]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][103] ) );
  DFF \modmult_1/zreg_reg[102]  ( .D(mod_mult_o[102]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][102] ) );
  DFF \modmult_1/zreg_reg[101]  ( .D(mod_mult_o[101]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][101] ) );
  DFF \modmult_1/zreg_reg[100]  ( .D(mod_mult_o[100]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][100] ) );
  DFF \modmult_1/zreg_reg[99]  ( .D(mod_mult_o[99]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][99] ) );
  DFF \modmult_1/zreg_reg[98]  ( .D(mod_mult_o[98]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][98] ) );
  DFF \modmult_1/zreg_reg[97]  ( .D(mod_mult_o[97]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][97] ) );
  DFF \modmult_1/zreg_reg[96]  ( .D(mod_mult_o[96]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][96] ) );
  DFF \modmult_1/zreg_reg[95]  ( .D(mod_mult_o[95]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][95] ) );
  DFF \modmult_1/zreg_reg[94]  ( .D(mod_mult_o[94]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][94] ) );
  DFF \modmult_1/zreg_reg[93]  ( .D(mod_mult_o[93]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][93] ) );
  DFF \modmult_1/zreg_reg[92]  ( .D(mod_mult_o[92]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][92] ) );
  DFF \modmult_1/zreg_reg[91]  ( .D(mod_mult_o[91]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][91] ) );
  DFF \modmult_1/zreg_reg[90]  ( .D(mod_mult_o[90]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][90] ) );
  DFF \modmult_1/zreg_reg[89]  ( .D(mod_mult_o[89]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][89] ) );
  DFF \modmult_1/zreg_reg[88]  ( .D(mod_mult_o[88]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][88] ) );
  DFF \modmult_1/zreg_reg[87]  ( .D(mod_mult_o[87]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][87] ) );
  DFF \modmult_1/zreg_reg[86]  ( .D(mod_mult_o[86]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][86] ) );
  DFF \modmult_1/zreg_reg[85]  ( .D(mod_mult_o[85]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][85] ) );
  DFF \modmult_1/zreg_reg[84]  ( .D(mod_mult_o[84]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][84] ) );
  DFF \modmult_1/zreg_reg[83]  ( .D(mod_mult_o[83]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][83] ) );
  DFF \modmult_1/zreg_reg[82]  ( .D(mod_mult_o[82]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][82] ) );
  DFF \modmult_1/zreg_reg[81]  ( .D(mod_mult_o[81]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][81] ) );
  DFF \modmult_1/zreg_reg[80]  ( .D(mod_mult_o[80]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][80] ) );
  DFF \modmult_1/zreg_reg[79]  ( .D(mod_mult_o[79]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][79] ) );
  DFF \modmult_1/zreg_reg[78]  ( .D(mod_mult_o[78]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][78] ) );
  DFF \modmult_1/zreg_reg[77]  ( .D(mod_mult_o[77]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][77] ) );
  DFF \modmult_1/zreg_reg[76]  ( .D(mod_mult_o[76]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][76] ) );
  DFF \modmult_1/zreg_reg[75]  ( .D(mod_mult_o[75]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][75] ) );
  DFF \modmult_1/zreg_reg[74]  ( .D(mod_mult_o[74]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][74] ) );
  DFF \modmult_1/zreg_reg[73]  ( .D(mod_mult_o[73]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][73] ) );
  DFF \modmult_1/zreg_reg[72]  ( .D(mod_mult_o[72]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][72] ) );
  DFF \modmult_1/zreg_reg[71]  ( .D(mod_mult_o[71]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][71] ) );
  DFF \modmult_1/zreg_reg[70]  ( .D(mod_mult_o[70]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][70] ) );
  DFF \modmult_1/zreg_reg[69]  ( .D(mod_mult_o[69]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][69] ) );
  DFF \modmult_1/zreg_reg[68]  ( .D(mod_mult_o[68]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][68] ) );
  DFF \modmult_1/zreg_reg[67]  ( .D(mod_mult_o[67]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][67] ) );
  DFF \modmult_1/zreg_reg[66]  ( .D(mod_mult_o[66]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][66] ) );
  DFF \modmult_1/zreg_reg[65]  ( .D(mod_mult_o[65]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][65] ) );
  DFF \modmult_1/zreg_reg[64]  ( .D(mod_mult_o[64]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][64] ) );
  DFF \modmult_1/zreg_reg[63]  ( .D(mod_mult_o[63]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][63] ) );
  DFF \modmult_1/zreg_reg[62]  ( .D(mod_mult_o[62]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][62] ) );
  DFF \modmult_1/zreg_reg[61]  ( .D(mod_mult_o[61]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][61] ) );
  DFF \modmult_1/zreg_reg[60]  ( .D(mod_mult_o[60]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][60] ) );
  DFF \modmult_1/zreg_reg[59]  ( .D(mod_mult_o[59]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][59] ) );
  DFF \modmult_1/zreg_reg[58]  ( .D(mod_mult_o[58]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][58] ) );
  DFF \modmult_1/zreg_reg[57]  ( .D(mod_mult_o[57]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][57] ) );
  DFF \modmult_1/zreg_reg[56]  ( .D(mod_mult_o[56]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][56] ) );
  DFF \modmult_1/zreg_reg[55]  ( .D(mod_mult_o[55]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][55] ) );
  DFF \modmult_1/zreg_reg[54]  ( .D(mod_mult_o[54]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][54] ) );
  DFF \modmult_1/zreg_reg[53]  ( .D(mod_mult_o[53]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][53] ) );
  DFF \modmult_1/zreg_reg[52]  ( .D(mod_mult_o[52]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][52] ) );
  DFF \modmult_1/zreg_reg[51]  ( .D(mod_mult_o[51]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][51] ) );
  DFF \modmult_1/zreg_reg[50]  ( .D(mod_mult_o[50]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][50] ) );
  DFF \modmult_1/zreg_reg[49]  ( .D(mod_mult_o[49]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][49] ) );
  DFF \modmult_1/zreg_reg[48]  ( .D(mod_mult_o[48]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][48] ) );
  DFF \modmult_1/zreg_reg[47]  ( .D(mod_mult_o[47]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][47] ) );
  DFF \modmult_1/zreg_reg[46]  ( .D(mod_mult_o[46]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][46] ) );
  DFF \modmult_1/zreg_reg[45]  ( .D(mod_mult_o[45]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][45] ) );
  DFF \modmult_1/zreg_reg[44]  ( .D(mod_mult_o[44]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][44] ) );
  DFF \modmult_1/zreg_reg[43]  ( .D(mod_mult_o[43]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][43] ) );
  DFF \modmult_1/zreg_reg[42]  ( .D(mod_mult_o[42]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][42] ) );
  DFF \modmult_1/zreg_reg[41]  ( .D(mod_mult_o[41]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][41] ) );
  DFF \modmult_1/zreg_reg[40]  ( .D(mod_mult_o[40]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][40] ) );
  DFF \modmult_1/zreg_reg[39]  ( .D(mod_mult_o[39]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][39] ) );
  DFF \modmult_1/zreg_reg[38]  ( .D(mod_mult_o[38]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][38] ) );
  DFF \modmult_1/zreg_reg[37]  ( .D(mod_mult_o[37]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][37] ) );
  DFF \modmult_1/zreg_reg[36]  ( .D(mod_mult_o[36]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][36] ) );
  DFF \modmult_1/zreg_reg[35]  ( .D(mod_mult_o[35]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][35] ) );
  DFF \modmult_1/zreg_reg[34]  ( .D(mod_mult_o[34]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][34] ) );
  DFF \modmult_1/zreg_reg[33]  ( .D(mod_mult_o[33]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][33] ) );
  DFF \modmult_1/zreg_reg[32]  ( .D(mod_mult_o[32]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][32] ) );
  DFF \modmult_1/zreg_reg[31]  ( .D(mod_mult_o[31]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][31] ) );
  DFF \modmult_1/zreg_reg[30]  ( .D(mod_mult_o[30]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][30] ) );
  DFF \modmult_1/zreg_reg[29]  ( .D(mod_mult_o[29]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][29] ) );
  DFF \modmult_1/zreg_reg[28]  ( .D(mod_mult_o[28]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][28] ) );
  DFF \modmult_1/zreg_reg[27]  ( .D(mod_mult_o[27]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][27] ) );
  DFF \modmult_1/zreg_reg[26]  ( .D(mod_mult_o[26]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][26] ) );
  DFF \modmult_1/zreg_reg[25]  ( .D(mod_mult_o[25]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][25] ) );
  DFF \modmult_1/zreg_reg[24]  ( .D(mod_mult_o[24]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][24] ) );
  DFF \modmult_1/zreg_reg[23]  ( .D(mod_mult_o[23]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][23] ) );
  DFF \modmult_1/zreg_reg[22]  ( .D(mod_mult_o[22]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][22] ) );
  DFF \modmult_1/zreg_reg[21]  ( .D(mod_mult_o[21]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][21] ) );
  DFF \modmult_1/zreg_reg[20]  ( .D(mod_mult_o[20]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][20] ) );
  DFF \modmult_1/zreg_reg[19]  ( .D(mod_mult_o[19]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][19] ) );
  DFF \modmult_1/zreg_reg[18]  ( .D(mod_mult_o[18]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][18] ) );
  DFF \modmult_1/zreg_reg[17]  ( .D(mod_mult_o[17]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][17] ) );
  DFF \modmult_1/zreg_reg[16]  ( .D(mod_mult_o[16]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][16] ) );
  DFF \modmult_1/zreg_reg[15]  ( .D(mod_mult_o[15]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][15] ) );
  DFF \modmult_1/zreg_reg[14]  ( .D(mod_mult_o[14]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][14] ) );
  DFF \modmult_1/zreg_reg[13]  ( .D(mod_mult_o[13]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][13] ) );
  DFF \modmult_1/zreg_reg[12]  ( .D(mod_mult_o[12]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][12] ) );
  DFF \modmult_1/zreg_reg[11]  ( .D(mod_mult_o[11]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][11] ) );
  DFF \modmult_1/zreg_reg[10]  ( .D(mod_mult_o[10]), .CLK(clk), .RST(
        start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][10] ) );
  DFF \modmult_1/zreg_reg[9]  ( .D(mod_mult_o[9]), .CLK(clk), .RST(start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][9] ) );
  DFF \modmult_1/zreg_reg[8]  ( .D(mod_mult_o[8]), .CLK(clk), .RST(start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][8] ) );
  DFF \modmult_1/zreg_reg[7]  ( .D(mod_mult_o[7]), .CLK(clk), .RST(start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][7] ) );
  DFF \modmult_1/zreg_reg[6]  ( .D(mod_mult_o[6]), .CLK(clk), .RST(start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][6] ) );
  DFF \modmult_1/zreg_reg[5]  ( .D(mod_mult_o[5]), .CLK(clk), .RST(start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][5] ) );
  DFF \modmult_1/zreg_reg[4]  ( .D(mod_mult_o[4]), .CLK(clk), .RST(start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][4] ) );
  DFF \modmult_1/zreg_reg[3]  ( .D(mod_mult_o[3]), .CLK(clk), .RST(start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][3] ) );
  DFF \modmult_1/zreg_reg[2]  ( .D(mod_mult_o[2]), .CLK(clk), .RST(start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][2] ) );
  DFF \modmult_1/zreg_reg[1]  ( .D(mod_mult_o[1]), .CLK(clk), .RST(start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][1] ) );
  DFF \modmult_1/zreg_reg[0]  ( .D(mod_mult_o[0]), .CLK(clk), .RST(start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][0] ) );
  DFF \modmult_1/xreg_reg[1023]  ( .D(\modmult_1/xin[1022] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[1023]), .Q(\modmult_1/xin[1023] ) );
  DFF \modmult_1/xreg_reg[1022]  ( .D(\modmult_1/xin[1021] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[1022]), .Q(\modmult_1/xin[1022] ) );
  DFF \modmult_1/xreg_reg[1021]  ( .D(\modmult_1/xin[1020] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[1021]), .Q(\modmult_1/xin[1021] ) );
  DFF \modmult_1/xreg_reg[1020]  ( .D(\modmult_1/xin[1019] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[1020]), .Q(\modmult_1/xin[1020] ) );
  DFF \modmult_1/xreg_reg[1019]  ( .D(\modmult_1/xin[1018] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[1019]), .Q(\modmult_1/xin[1019] ) );
  DFF \modmult_1/xreg_reg[1018]  ( .D(\modmult_1/xin[1017] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[1018]), .Q(\modmult_1/xin[1018] ) );
  DFF \modmult_1/xreg_reg[1017]  ( .D(\modmult_1/xin[1016] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[1017]), .Q(\modmult_1/xin[1017] ) );
  DFF \modmult_1/xreg_reg[1016]  ( .D(\modmult_1/xin[1015] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[1016]), .Q(\modmult_1/xin[1016] ) );
  DFF \modmult_1/xreg_reg[1015]  ( .D(\modmult_1/xin[1014] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[1015]), .Q(\modmult_1/xin[1015] ) );
  DFF \modmult_1/xreg_reg[1014]  ( .D(\modmult_1/xin[1013] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[1014]), .Q(\modmult_1/xin[1014] ) );
  DFF \modmult_1/xreg_reg[1013]  ( .D(\modmult_1/xin[1012] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[1013]), .Q(\modmult_1/xin[1013] ) );
  DFF \modmult_1/xreg_reg[1012]  ( .D(\modmult_1/xin[1011] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[1012]), .Q(\modmult_1/xin[1012] ) );
  DFF \modmult_1/xreg_reg[1011]  ( .D(\modmult_1/xin[1010] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[1011]), .Q(\modmult_1/xin[1011] ) );
  DFF \modmult_1/xreg_reg[1010]  ( .D(\modmult_1/xin[1009] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[1010]), .Q(\modmult_1/xin[1010] ) );
  DFF \modmult_1/xreg_reg[1009]  ( .D(\modmult_1/xin[1008] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[1009]), .Q(\modmult_1/xin[1009] ) );
  DFF \modmult_1/xreg_reg[1008]  ( .D(\modmult_1/xin[1007] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[1008]), .Q(\modmult_1/xin[1008] ) );
  DFF \modmult_1/xreg_reg[1007]  ( .D(\modmult_1/xin[1006] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[1007]), .Q(\modmult_1/xin[1007] ) );
  DFF \modmult_1/xreg_reg[1006]  ( .D(\modmult_1/xin[1005] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[1006]), .Q(\modmult_1/xin[1006] ) );
  DFF \modmult_1/xreg_reg[1005]  ( .D(\modmult_1/xin[1004] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[1005]), .Q(\modmult_1/xin[1005] ) );
  DFF \modmult_1/xreg_reg[1004]  ( .D(\modmult_1/xin[1003] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[1004]), .Q(\modmult_1/xin[1004] ) );
  DFF \modmult_1/xreg_reg[1003]  ( .D(\modmult_1/xin[1002] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[1003]), .Q(\modmult_1/xin[1003] ) );
  DFF \modmult_1/xreg_reg[1002]  ( .D(\modmult_1/xin[1001] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[1002]), .Q(\modmult_1/xin[1002] ) );
  DFF \modmult_1/xreg_reg[1001]  ( .D(\modmult_1/xin[1000] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[1001]), .Q(\modmult_1/xin[1001] ) );
  DFF \modmult_1/xreg_reg[1000]  ( .D(\modmult_1/xin[999] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[1000]), .Q(\modmult_1/xin[1000] ) );
  DFF \modmult_1/xreg_reg[999]  ( .D(\modmult_1/xin[998] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[999]), .Q(\modmult_1/xin[999] ) );
  DFF \modmult_1/xreg_reg[998]  ( .D(\modmult_1/xin[997] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[998]), .Q(\modmult_1/xin[998] ) );
  DFF \modmult_1/xreg_reg[997]  ( .D(\modmult_1/xin[996] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[997]), .Q(\modmult_1/xin[997] ) );
  DFF \modmult_1/xreg_reg[996]  ( .D(\modmult_1/xin[995] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[996]), .Q(\modmult_1/xin[996] ) );
  DFF \modmult_1/xreg_reg[995]  ( .D(\modmult_1/xin[994] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[995]), .Q(\modmult_1/xin[995] ) );
  DFF \modmult_1/xreg_reg[994]  ( .D(\modmult_1/xin[993] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[994]), .Q(\modmult_1/xin[994] ) );
  DFF \modmult_1/xreg_reg[993]  ( .D(\modmult_1/xin[992] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[993]), .Q(\modmult_1/xin[993] ) );
  DFF \modmult_1/xreg_reg[992]  ( .D(\modmult_1/xin[991] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[992]), .Q(\modmult_1/xin[992] ) );
  DFF \modmult_1/xreg_reg[991]  ( .D(\modmult_1/xin[990] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[991]), .Q(\modmult_1/xin[991] ) );
  DFF \modmult_1/xreg_reg[990]  ( .D(\modmult_1/xin[989] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[990]), .Q(\modmult_1/xin[990] ) );
  DFF \modmult_1/xreg_reg[989]  ( .D(\modmult_1/xin[988] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[989]), .Q(\modmult_1/xin[989] ) );
  DFF \modmult_1/xreg_reg[988]  ( .D(\modmult_1/xin[987] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[988]), .Q(\modmult_1/xin[988] ) );
  DFF \modmult_1/xreg_reg[987]  ( .D(\modmult_1/xin[986] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[987]), .Q(\modmult_1/xin[987] ) );
  DFF \modmult_1/xreg_reg[986]  ( .D(\modmult_1/xin[985] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[986]), .Q(\modmult_1/xin[986] ) );
  DFF \modmult_1/xreg_reg[985]  ( .D(\modmult_1/xin[984] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[985]), .Q(\modmult_1/xin[985] ) );
  DFF \modmult_1/xreg_reg[984]  ( .D(\modmult_1/xin[983] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[984]), .Q(\modmult_1/xin[984] ) );
  DFF \modmult_1/xreg_reg[983]  ( .D(\modmult_1/xin[982] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[983]), .Q(\modmult_1/xin[983] ) );
  DFF \modmult_1/xreg_reg[982]  ( .D(\modmult_1/xin[981] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[982]), .Q(\modmult_1/xin[982] ) );
  DFF \modmult_1/xreg_reg[981]  ( .D(\modmult_1/xin[980] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[981]), .Q(\modmult_1/xin[981] ) );
  DFF \modmult_1/xreg_reg[980]  ( .D(\modmult_1/xin[979] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[980]), .Q(\modmult_1/xin[980] ) );
  DFF \modmult_1/xreg_reg[979]  ( .D(\modmult_1/xin[978] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[979]), .Q(\modmult_1/xin[979] ) );
  DFF \modmult_1/xreg_reg[978]  ( .D(\modmult_1/xin[977] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[978]), .Q(\modmult_1/xin[978] ) );
  DFF \modmult_1/xreg_reg[977]  ( .D(\modmult_1/xin[976] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[977]), .Q(\modmult_1/xin[977] ) );
  DFF \modmult_1/xreg_reg[976]  ( .D(\modmult_1/xin[975] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[976]), .Q(\modmult_1/xin[976] ) );
  DFF \modmult_1/xreg_reg[975]  ( .D(\modmult_1/xin[974] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[975]), .Q(\modmult_1/xin[975] ) );
  DFF \modmult_1/xreg_reg[974]  ( .D(\modmult_1/xin[973] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[974]), .Q(\modmult_1/xin[974] ) );
  DFF \modmult_1/xreg_reg[973]  ( .D(\modmult_1/xin[972] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[973]), .Q(\modmult_1/xin[973] ) );
  DFF \modmult_1/xreg_reg[972]  ( .D(\modmult_1/xin[971] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[972]), .Q(\modmult_1/xin[972] ) );
  DFF \modmult_1/xreg_reg[971]  ( .D(\modmult_1/xin[970] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[971]), .Q(\modmult_1/xin[971] ) );
  DFF \modmult_1/xreg_reg[970]  ( .D(\modmult_1/xin[969] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[970]), .Q(\modmult_1/xin[970] ) );
  DFF \modmult_1/xreg_reg[969]  ( .D(\modmult_1/xin[968] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[969]), .Q(\modmult_1/xin[969] ) );
  DFF \modmult_1/xreg_reg[968]  ( .D(\modmult_1/xin[967] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[968]), .Q(\modmult_1/xin[968] ) );
  DFF \modmult_1/xreg_reg[967]  ( .D(\modmult_1/xin[966] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[967]), .Q(\modmult_1/xin[967] ) );
  DFF \modmult_1/xreg_reg[966]  ( .D(\modmult_1/xin[965] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[966]), .Q(\modmult_1/xin[966] ) );
  DFF \modmult_1/xreg_reg[965]  ( .D(\modmult_1/xin[964] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[965]), .Q(\modmult_1/xin[965] ) );
  DFF \modmult_1/xreg_reg[964]  ( .D(\modmult_1/xin[963] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[964]), .Q(\modmult_1/xin[964] ) );
  DFF \modmult_1/xreg_reg[963]  ( .D(\modmult_1/xin[962] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[963]), .Q(\modmult_1/xin[963] ) );
  DFF \modmult_1/xreg_reg[962]  ( .D(\modmult_1/xin[961] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[962]), .Q(\modmult_1/xin[962] ) );
  DFF \modmult_1/xreg_reg[961]  ( .D(\modmult_1/xin[960] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[961]), .Q(\modmult_1/xin[961] ) );
  DFF \modmult_1/xreg_reg[960]  ( .D(\modmult_1/xin[959] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[960]), .Q(\modmult_1/xin[960] ) );
  DFF \modmult_1/xreg_reg[959]  ( .D(\modmult_1/xin[958] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[959]), .Q(\modmult_1/xin[959] ) );
  DFF \modmult_1/xreg_reg[958]  ( .D(\modmult_1/xin[957] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[958]), .Q(\modmult_1/xin[958] ) );
  DFF \modmult_1/xreg_reg[957]  ( .D(\modmult_1/xin[956] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[957]), .Q(\modmult_1/xin[957] ) );
  DFF \modmult_1/xreg_reg[956]  ( .D(\modmult_1/xin[955] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[956]), .Q(\modmult_1/xin[956] ) );
  DFF \modmult_1/xreg_reg[955]  ( .D(\modmult_1/xin[954] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[955]), .Q(\modmult_1/xin[955] ) );
  DFF \modmult_1/xreg_reg[954]  ( .D(\modmult_1/xin[953] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[954]), .Q(\modmult_1/xin[954] ) );
  DFF \modmult_1/xreg_reg[953]  ( .D(\modmult_1/xin[952] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[953]), .Q(\modmult_1/xin[953] ) );
  DFF \modmult_1/xreg_reg[952]  ( .D(\modmult_1/xin[951] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[952]), .Q(\modmult_1/xin[952] ) );
  DFF \modmult_1/xreg_reg[951]  ( .D(\modmult_1/xin[950] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[951]), .Q(\modmult_1/xin[951] ) );
  DFF \modmult_1/xreg_reg[950]  ( .D(\modmult_1/xin[949] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[950]), .Q(\modmult_1/xin[950] ) );
  DFF \modmult_1/xreg_reg[949]  ( .D(\modmult_1/xin[948] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[949]), .Q(\modmult_1/xin[949] ) );
  DFF \modmult_1/xreg_reg[948]  ( .D(\modmult_1/xin[947] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[948]), .Q(\modmult_1/xin[948] ) );
  DFF \modmult_1/xreg_reg[947]  ( .D(\modmult_1/xin[946] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[947]), .Q(\modmult_1/xin[947] ) );
  DFF \modmult_1/xreg_reg[946]  ( .D(\modmult_1/xin[945] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[946]), .Q(\modmult_1/xin[946] ) );
  DFF \modmult_1/xreg_reg[945]  ( .D(\modmult_1/xin[944] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[945]), .Q(\modmult_1/xin[945] ) );
  DFF \modmult_1/xreg_reg[944]  ( .D(\modmult_1/xin[943] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[944]), .Q(\modmult_1/xin[944] ) );
  DFF \modmult_1/xreg_reg[943]  ( .D(\modmult_1/xin[942] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[943]), .Q(\modmult_1/xin[943] ) );
  DFF \modmult_1/xreg_reg[942]  ( .D(\modmult_1/xin[941] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[942]), .Q(\modmult_1/xin[942] ) );
  DFF \modmult_1/xreg_reg[941]  ( .D(\modmult_1/xin[940] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[941]), .Q(\modmult_1/xin[941] ) );
  DFF \modmult_1/xreg_reg[940]  ( .D(\modmult_1/xin[939] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[940]), .Q(\modmult_1/xin[940] ) );
  DFF \modmult_1/xreg_reg[939]  ( .D(\modmult_1/xin[938] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[939]), .Q(\modmult_1/xin[939] ) );
  DFF \modmult_1/xreg_reg[938]  ( .D(\modmult_1/xin[937] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[938]), .Q(\modmult_1/xin[938] ) );
  DFF \modmult_1/xreg_reg[937]  ( .D(\modmult_1/xin[936] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[937]), .Q(\modmult_1/xin[937] ) );
  DFF \modmult_1/xreg_reg[936]  ( .D(\modmult_1/xin[935] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[936]), .Q(\modmult_1/xin[936] ) );
  DFF \modmult_1/xreg_reg[935]  ( .D(\modmult_1/xin[934] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[935]), .Q(\modmult_1/xin[935] ) );
  DFF \modmult_1/xreg_reg[934]  ( .D(\modmult_1/xin[933] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[934]), .Q(\modmult_1/xin[934] ) );
  DFF \modmult_1/xreg_reg[933]  ( .D(\modmult_1/xin[932] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[933]), .Q(\modmult_1/xin[933] ) );
  DFF \modmult_1/xreg_reg[932]  ( .D(\modmult_1/xin[931] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[932]), .Q(\modmult_1/xin[932] ) );
  DFF \modmult_1/xreg_reg[931]  ( .D(\modmult_1/xin[930] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[931]), .Q(\modmult_1/xin[931] ) );
  DFF \modmult_1/xreg_reg[930]  ( .D(\modmult_1/xin[929] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[930]), .Q(\modmult_1/xin[930] ) );
  DFF \modmult_1/xreg_reg[929]  ( .D(\modmult_1/xin[928] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[929]), .Q(\modmult_1/xin[929] ) );
  DFF \modmult_1/xreg_reg[928]  ( .D(\modmult_1/xin[927] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[928]), .Q(\modmult_1/xin[928] ) );
  DFF \modmult_1/xreg_reg[927]  ( .D(\modmult_1/xin[926] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[927]), .Q(\modmult_1/xin[927] ) );
  DFF \modmult_1/xreg_reg[926]  ( .D(\modmult_1/xin[925] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[926]), .Q(\modmult_1/xin[926] ) );
  DFF \modmult_1/xreg_reg[925]  ( .D(\modmult_1/xin[924] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[925]), .Q(\modmult_1/xin[925] ) );
  DFF \modmult_1/xreg_reg[924]  ( .D(\modmult_1/xin[923] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[924]), .Q(\modmult_1/xin[924] ) );
  DFF \modmult_1/xreg_reg[923]  ( .D(\modmult_1/xin[922] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[923]), .Q(\modmult_1/xin[923] ) );
  DFF \modmult_1/xreg_reg[922]  ( .D(\modmult_1/xin[921] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[922]), .Q(\modmult_1/xin[922] ) );
  DFF \modmult_1/xreg_reg[921]  ( .D(\modmult_1/xin[920] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[921]), .Q(\modmult_1/xin[921] ) );
  DFF \modmult_1/xreg_reg[920]  ( .D(\modmult_1/xin[919] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[920]), .Q(\modmult_1/xin[920] ) );
  DFF \modmult_1/xreg_reg[919]  ( .D(\modmult_1/xin[918] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[919]), .Q(\modmult_1/xin[919] ) );
  DFF \modmult_1/xreg_reg[918]  ( .D(\modmult_1/xin[917] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[918]), .Q(\modmult_1/xin[918] ) );
  DFF \modmult_1/xreg_reg[917]  ( .D(\modmult_1/xin[916] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[917]), .Q(\modmult_1/xin[917] ) );
  DFF \modmult_1/xreg_reg[916]  ( .D(\modmult_1/xin[915] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[916]), .Q(\modmult_1/xin[916] ) );
  DFF \modmult_1/xreg_reg[915]  ( .D(\modmult_1/xin[914] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[915]), .Q(\modmult_1/xin[915] ) );
  DFF \modmult_1/xreg_reg[914]  ( .D(\modmult_1/xin[913] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[914]), .Q(\modmult_1/xin[914] ) );
  DFF \modmult_1/xreg_reg[913]  ( .D(\modmult_1/xin[912] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[913]), .Q(\modmult_1/xin[913] ) );
  DFF \modmult_1/xreg_reg[912]  ( .D(\modmult_1/xin[911] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[912]), .Q(\modmult_1/xin[912] ) );
  DFF \modmult_1/xreg_reg[911]  ( .D(\modmult_1/xin[910] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[911]), .Q(\modmult_1/xin[911] ) );
  DFF \modmult_1/xreg_reg[910]  ( .D(\modmult_1/xin[909] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[910]), .Q(\modmult_1/xin[910] ) );
  DFF \modmult_1/xreg_reg[909]  ( .D(\modmult_1/xin[908] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[909]), .Q(\modmult_1/xin[909] ) );
  DFF \modmult_1/xreg_reg[908]  ( .D(\modmult_1/xin[907] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[908]), .Q(\modmult_1/xin[908] ) );
  DFF \modmult_1/xreg_reg[907]  ( .D(\modmult_1/xin[906] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[907]), .Q(\modmult_1/xin[907] ) );
  DFF \modmult_1/xreg_reg[906]  ( .D(\modmult_1/xin[905] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[906]), .Q(\modmult_1/xin[906] ) );
  DFF \modmult_1/xreg_reg[905]  ( .D(\modmult_1/xin[904] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[905]), .Q(\modmult_1/xin[905] ) );
  DFF \modmult_1/xreg_reg[904]  ( .D(\modmult_1/xin[903] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[904]), .Q(\modmult_1/xin[904] ) );
  DFF \modmult_1/xreg_reg[903]  ( .D(\modmult_1/xin[902] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[903]), .Q(\modmult_1/xin[903] ) );
  DFF \modmult_1/xreg_reg[902]  ( .D(\modmult_1/xin[901] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[902]), .Q(\modmult_1/xin[902] ) );
  DFF \modmult_1/xreg_reg[901]  ( .D(\modmult_1/xin[900] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[901]), .Q(\modmult_1/xin[901] ) );
  DFF \modmult_1/xreg_reg[900]  ( .D(\modmult_1/xin[899] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[900]), .Q(\modmult_1/xin[900] ) );
  DFF \modmult_1/xreg_reg[899]  ( .D(\modmult_1/xin[898] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[899]), .Q(\modmult_1/xin[899] ) );
  DFF \modmult_1/xreg_reg[898]  ( .D(\modmult_1/xin[897] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[898]), .Q(\modmult_1/xin[898] ) );
  DFF \modmult_1/xreg_reg[897]  ( .D(\modmult_1/xin[896] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[897]), .Q(\modmult_1/xin[897] ) );
  DFF \modmult_1/xreg_reg[896]  ( .D(\modmult_1/xin[895] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[896]), .Q(\modmult_1/xin[896] ) );
  DFF \modmult_1/xreg_reg[895]  ( .D(\modmult_1/xin[894] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[895]), .Q(\modmult_1/xin[895] ) );
  DFF \modmult_1/xreg_reg[894]  ( .D(\modmult_1/xin[893] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[894]), .Q(\modmult_1/xin[894] ) );
  DFF \modmult_1/xreg_reg[893]  ( .D(\modmult_1/xin[892] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[893]), .Q(\modmult_1/xin[893] ) );
  DFF \modmult_1/xreg_reg[892]  ( .D(\modmult_1/xin[891] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[892]), .Q(\modmult_1/xin[892] ) );
  DFF \modmult_1/xreg_reg[891]  ( .D(\modmult_1/xin[890] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[891]), .Q(\modmult_1/xin[891] ) );
  DFF \modmult_1/xreg_reg[890]  ( .D(\modmult_1/xin[889] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[890]), .Q(\modmult_1/xin[890] ) );
  DFF \modmult_1/xreg_reg[889]  ( .D(\modmult_1/xin[888] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[889]), .Q(\modmult_1/xin[889] ) );
  DFF \modmult_1/xreg_reg[888]  ( .D(\modmult_1/xin[887] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[888]), .Q(\modmult_1/xin[888] ) );
  DFF \modmult_1/xreg_reg[887]  ( .D(\modmult_1/xin[886] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[887]), .Q(\modmult_1/xin[887] ) );
  DFF \modmult_1/xreg_reg[886]  ( .D(\modmult_1/xin[885] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[886]), .Q(\modmult_1/xin[886] ) );
  DFF \modmult_1/xreg_reg[885]  ( .D(\modmult_1/xin[884] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[885]), .Q(\modmult_1/xin[885] ) );
  DFF \modmult_1/xreg_reg[884]  ( .D(\modmult_1/xin[883] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[884]), .Q(\modmult_1/xin[884] ) );
  DFF \modmult_1/xreg_reg[883]  ( .D(\modmult_1/xin[882] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[883]), .Q(\modmult_1/xin[883] ) );
  DFF \modmult_1/xreg_reg[882]  ( .D(\modmult_1/xin[881] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[882]), .Q(\modmult_1/xin[882] ) );
  DFF \modmult_1/xreg_reg[881]  ( .D(\modmult_1/xin[880] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[881]), .Q(\modmult_1/xin[881] ) );
  DFF \modmult_1/xreg_reg[880]  ( .D(\modmult_1/xin[879] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[880]), .Q(\modmult_1/xin[880] ) );
  DFF \modmult_1/xreg_reg[879]  ( .D(\modmult_1/xin[878] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[879]), .Q(\modmult_1/xin[879] ) );
  DFF \modmult_1/xreg_reg[878]  ( .D(\modmult_1/xin[877] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[878]), .Q(\modmult_1/xin[878] ) );
  DFF \modmult_1/xreg_reg[877]  ( .D(\modmult_1/xin[876] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[877]), .Q(\modmult_1/xin[877] ) );
  DFF \modmult_1/xreg_reg[876]  ( .D(\modmult_1/xin[875] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[876]), .Q(\modmult_1/xin[876] ) );
  DFF \modmult_1/xreg_reg[875]  ( .D(\modmult_1/xin[874] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[875]), .Q(\modmult_1/xin[875] ) );
  DFF \modmult_1/xreg_reg[874]  ( .D(\modmult_1/xin[873] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[874]), .Q(\modmult_1/xin[874] ) );
  DFF \modmult_1/xreg_reg[873]  ( .D(\modmult_1/xin[872] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[873]), .Q(\modmult_1/xin[873] ) );
  DFF \modmult_1/xreg_reg[872]  ( .D(\modmult_1/xin[871] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[872]), .Q(\modmult_1/xin[872] ) );
  DFF \modmult_1/xreg_reg[871]  ( .D(\modmult_1/xin[870] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[871]), .Q(\modmult_1/xin[871] ) );
  DFF \modmult_1/xreg_reg[870]  ( .D(\modmult_1/xin[869] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[870]), .Q(\modmult_1/xin[870] ) );
  DFF \modmult_1/xreg_reg[869]  ( .D(\modmult_1/xin[868] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[869]), .Q(\modmult_1/xin[869] ) );
  DFF \modmult_1/xreg_reg[868]  ( .D(\modmult_1/xin[867] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[868]), .Q(\modmult_1/xin[868] ) );
  DFF \modmult_1/xreg_reg[867]  ( .D(\modmult_1/xin[866] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[867]), .Q(\modmult_1/xin[867] ) );
  DFF \modmult_1/xreg_reg[866]  ( .D(\modmult_1/xin[865] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[866]), .Q(\modmult_1/xin[866] ) );
  DFF \modmult_1/xreg_reg[865]  ( .D(\modmult_1/xin[864] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[865]), .Q(\modmult_1/xin[865] ) );
  DFF \modmult_1/xreg_reg[864]  ( .D(\modmult_1/xin[863] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[864]), .Q(\modmult_1/xin[864] ) );
  DFF \modmult_1/xreg_reg[863]  ( .D(\modmult_1/xin[862] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[863]), .Q(\modmult_1/xin[863] ) );
  DFF \modmult_1/xreg_reg[862]  ( .D(\modmult_1/xin[861] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[862]), .Q(\modmult_1/xin[862] ) );
  DFF \modmult_1/xreg_reg[861]  ( .D(\modmult_1/xin[860] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[861]), .Q(\modmult_1/xin[861] ) );
  DFF \modmult_1/xreg_reg[860]  ( .D(\modmult_1/xin[859] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[860]), .Q(\modmult_1/xin[860] ) );
  DFF \modmult_1/xreg_reg[859]  ( .D(\modmult_1/xin[858] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[859]), .Q(\modmult_1/xin[859] ) );
  DFF \modmult_1/xreg_reg[858]  ( .D(\modmult_1/xin[857] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[858]), .Q(\modmult_1/xin[858] ) );
  DFF \modmult_1/xreg_reg[857]  ( .D(\modmult_1/xin[856] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[857]), .Q(\modmult_1/xin[857] ) );
  DFF \modmult_1/xreg_reg[856]  ( .D(\modmult_1/xin[855] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[856]), .Q(\modmult_1/xin[856] ) );
  DFF \modmult_1/xreg_reg[855]  ( .D(\modmult_1/xin[854] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[855]), .Q(\modmult_1/xin[855] ) );
  DFF \modmult_1/xreg_reg[854]  ( .D(\modmult_1/xin[853] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[854]), .Q(\modmult_1/xin[854] ) );
  DFF \modmult_1/xreg_reg[853]  ( .D(\modmult_1/xin[852] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[853]), .Q(\modmult_1/xin[853] ) );
  DFF \modmult_1/xreg_reg[852]  ( .D(\modmult_1/xin[851] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[852]), .Q(\modmult_1/xin[852] ) );
  DFF \modmult_1/xreg_reg[851]  ( .D(\modmult_1/xin[850] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[851]), .Q(\modmult_1/xin[851] ) );
  DFF \modmult_1/xreg_reg[850]  ( .D(\modmult_1/xin[849] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[850]), .Q(\modmult_1/xin[850] ) );
  DFF \modmult_1/xreg_reg[849]  ( .D(\modmult_1/xin[848] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[849]), .Q(\modmult_1/xin[849] ) );
  DFF \modmult_1/xreg_reg[848]  ( .D(\modmult_1/xin[847] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[848]), .Q(\modmult_1/xin[848] ) );
  DFF \modmult_1/xreg_reg[847]  ( .D(\modmult_1/xin[846] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[847]), .Q(\modmult_1/xin[847] ) );
  DFF \modmult_1/xreg_reg[846]  ( .D(\modmult_1/xin[845] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[846]), .Q(\modmult_1/xin[846] ) );
  DFF \modmult_1/xreg_reg[845]  ( .D(\modmult_1/xin[844] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[845]), .Q(\modmult_1/xin[845] ) );
  DFF \modmult_1/xreg_reg[844]  ( .D(\modmult_1/xin[843] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[844]), .Q(\modmult_1/xin[844] ) );
  DFF \modmult_1/xreg_reg[843]  ( .D(\modmult_1/xin[842] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[843]), .Q(\modmult_1/xin[843] ) );
  DFF \modmult_1/xreg_reg[842]  ( .D(\modmult_1/xin[841] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[842]), .Q(\modmult_1/xin[842] ) );
  DFF \modmult_1/xreg_reg[841]  ( .D(\modmult_1/xin[840] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[841]), .Q(\modmult_1/xin[841] ) );
  DFF \modmult_1/xreg_reg[840]  ( .D(\modmult_1/xin[839] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[840]), .Q(\modmult_1/xin[840] ) );
  DFF \modmult_1/xreg_reg[839]  ( .D(\modmult_1/xin[838] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[839]), .Q(\modmult_1/xin[839] ) );
  DFF \modmult_1/xreg_reg[838]  ( .D(\modmult_1/xin[837] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[838]), .Q(\modmult_1/xin[838] ) );
  DFF \modmult_1/xreg_reg[837]  ( .D(\modmult_1/xin[836] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[837]), .Q(\modmult_1/xin[837] ) );
  DFF \modmult_1/xreg_reg[836]  ( .D(\modmult_1/xin[835] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[836]), .Q(\modmult_1/xin[836] ) );
  DFF \modmult_1/xreg_reg[835]  ( .D(\modmult_1/xin[834] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[835]), .Q(\modmult_1/xin[835] ) );
  DFF \modmult_1/xreg_reg[834]  ( .D(\modmult_1/xin[833] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[834]), .Q(\modmult_1/xin[834] ) );
  DFF \modmult_1/xreg_reg[833]  ( .D(\modmult_1/xin[832] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[833]), .Q(\modmult_1/xin[833] ) );
  DFF \modmult_1/xreg_reg[832]  ( .D(\modmult_1/xin[831] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[832]), .Q(\modmult_1/xin[832] ) );
  DFF \modmult_1/xreg_reg[831]  ( .D(\modmult_1/xin[830] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[831]), .Q(\modmult_1/xin[831] ) );
  DFF \modmult_1/xreg_reg[830]  ( .D(\modmult_1/xin[829] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[830]), .Q(\modmult_1/xin[830] ) );
  DFF \modmult_1/xreg_reg[829]  ( .D(\modmult_1/xin[828] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[829]), .Q(\modmult_1/xin[829] ) );
  DFF \modmult_1/xreg_reg[828]  ( .D(\modmult_1/xin[827] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[828]), .Q(\modmult_1/xin[828] ) );
  DFF \modmult_1/xreg_reg[827]  ( .D(\modmult_1/xin[826] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[827]), .Q(\modmult_1/xin[827] ) );
  DFF \modmult_1/xreg_reg[826]  ( .D(\modmult_1/xin[825] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[826]), .Q(\modmult_1/xin[826] ) );
  DFF \modmult_1/xreg_reg[825]  ( .D(\modmult_1/xin[824] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[825]), .Q(\modmult_1/xin[825] ) );
  DFF \modmult_1/xreg_reg[824]  ( .D(\modmult_1/xin[823] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[824]), .Q(\modmult_1/xin[824] ) );
  DFF \modmult_1/xreg_reg[823]  ( .D(\modmult_1/xin[822] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[823]), .Q(\modmult_1/xin[823] ) );
  DFF \modmult_1/xreg_reg[822]  ( .D(\modmult_1/xin[821] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[822]), .Q(\modmult_1/xin[822] ) );
  DFF \modmult_1/xreg_reg[821]  ( .D(\modmult_1/xin[820] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[821]), .Q(\modmult_1/xin[821] ) );
  DFF \modmult_1/xreg_reg[820]  ( .D(\modmult_1/xin[819] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[820]), .Q(\modmult_1/xin[820] ) );
  DFF \modmult_1/xreg_reg[819]  ( .D(\modmult_1/xin[818] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[819]), .Q(\modmult_1/xin[819] ) );
  DFF \modmult_1/xreg_reg[818]  ( .D(\modmult_1/xin[817] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[818]), .Q(\modmult_1/xin[818] ) );
  DFF \modmult_1/xreg_reg[817]  ( .D(\modmult_1/xin[816] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[817]), .Q(\modmult_1/xin[817] ) );
  DFF \modmult_1/xreg_reg[816]  ( .D(\modmult_1/xin[815] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[816]), .Q(\modmult_1/xin[816] ) );
  DFF \modmult_1/xreg_reg[815]  ( .D(\modmult_1/xin[814] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[815]), .Q(\modmult_1/xin[815] ) );
  DFF \modmult_1/xreg_reg[814]  ( .D(\modmult_1/xin[813] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[814]), .Q(\modmult_1/xin[814] ) );
  DFF \modmult_1/xreg_reg[813]  ( .D(\modmult_1/xin[812] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[813]), .Q(\modmult_1/xin[813] ) );
  DFF \modmult_1/xreg_reg[812]  ( .D(\modmult_1/xin[811] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[812]), .Q(\modmult_1/xin[812] ) );
  DFF \modmult_1/xreg_reg[811]  ( .D(\modmult_1/xin[810] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[811]), .Q(\modmult_1/xin[811] ) );
  DFF \modmult_1/xreg_reg[810]  ( .D(\modmult_1/xin[809] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[810]), .Q(\modmult_1/xin[810] ) );
  DFF \modmult_1/xreg_reg[809]  ( .D(\modmult_1/xin[808] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[809]), .Q(\modmult_1/xin[809] ) );
  DFF \modmult_1/xreg_reg[808]  ( .D(\modmult_1/xin[807] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[808]), .Q(\modmult_1/xin[808] ) );
  DFF \modmult_1/xreg_reg[807]  ( .D(\modmult_1/xin[806] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[807]), .Q(\modmult_1/xin[807] ) );
  DFF \modmult_1/xreg_reg[806]  ( .D(\modmult_1/xin[805] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[806]), .Q(\modmult_1/xin[806] ) );
  DFF \modmult_1/xreg_reg[805]  ( .D(\modmult_1/xin[804] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[805]), .Q(\modmult_1/xin[805] ) );
  DFF \modmult_1/xreg_reg[804]  ( .D(\modmult_1/xin[803] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[804]), .Q(\modmult_1/xin[804] ) );
  DFF \modmult_1/xreg_reg[803]  ( .D(\modmult_1/xin[802] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[803]), .Q(\modmult_1/xin[803] ) );
  DFF \modmult_1/xreg_reg[802]  ( .D(\modmult_1/xin[801] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[802]), .Q(\modmult_1/xin[802] ) );
  DFF \modmult_1/xreg_reg[801]  ( .D(\modmult_1/xin[800] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[801]), .Q(\modmult_1/xin[801] ) );
  DFF \modmult_1/xreg_reg[800]  ( .D(\modmult_1/xin[799] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[800]), .Q(\modmult_1/xin[800] ) );
  DFF \modmult_1/xreg_reg[799]  ( .D(\modmult_1/xin[798] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[799]), .Q(\modmult_1/xin[799] ) );
  DFF \modmult_1/xreg_reg[798]  ( .D(\modmult_1/xin[797] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[798]), .Q(\modmult_1/xin[798] ) );
  DFF \modmult_1/xreg_reg[797]  ( .D(\modmult_1/xin[796] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[797]), .Q(\modmult_1/xin[797] ) );
  DFF \modmult_1/xreg_reg[796]  ( .D(\modmult_1/xin[795] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[796]), .Q(\modmult_1/xin[796] ) );
  DFF \modmult_1/xreg_reg[795]  ( .D(\modmult_1/xin[794] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[795]), .Q(\modmult_1/xin[795] ) );
  DFF \modmult_1/xreg_reg[794]  ( .D(\modmult_1/xin[793] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[794]), .Q(\modmult_1/xin[794] ) );
  DFF \modmult_1/xreg_reg[793]  ( .D(\modmult_1/xin[792] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[793]), .Q(\modmult_1/xin[793] ) );
  DFF \modmult_1/xreg_reg[792]  ( .D(\modmult_1/xin[791] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[792]), .Q(\modmult_1/xin[792] ) );
  DFF \modmult_1/xreg_reg[791]  ( .D(\modmult_1/xin[790] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[791]), .Q(\modmult_1/xin[791] ) );
  DFF \modmult_1/xreg_reg[790]  ( .D(\modmult_1/xin[789] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[790]), .Q(\modmult_1/xin[790] ) );
  DFF \modmult_1/xreg_reg[789]  ( .D(\modmult_1/xin[788] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[789]), .Q(\modmult_1/xin[789] ) );
  DFF \modmult_1/xreg_reg[788]  ( .D(\modmult_1/xin[787] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[788]), .Q(\modmult_1/xin[788] ) );
  DFF \modmult_1/xreg_reg[787]  ( .D(\modmult_1/xin[786] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[787]), .Q(\modmult_1/xin[787] ) );
  DFF \modmult_1/xreg_reg[786]  ( .D(\modmult_1/xin[785] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[786]), .Q(\modmult_1/xin[786] ) );
  DFF \modmult_1/xreg_reg[785]  ( .D(\modmult_1/xin[784] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[785]), .Q(\modmult_1/xin[785] ) );
  DFF \modmult_1/xreg_reg[784]  ( .D(\modmult_1/xin[783] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[784]), .Q(\modmult_1/xin[784] ) );
  DFF \modmult_1/xreg_reg[783]  ( .D(\modmult_1/xin[782] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[783]), .Q(\modmult_1/xin[783] ) );
  DFF \modmult_1/xreg_reg[782]  ( .D(\modmult_1/xin[781] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[782]), .Q(\modmult_1/xin[782] ) );
  DFF \modmult_1/xreg_reg[781]  ( .D(\modmult_1/xin[780] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[781]), .Q(\modmult_1/xin[781] ) );
  DFF \modmult_1/xreg_reg[780]  ( .D(\modmult_1/xin[779] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[780]), .Q(\modmult_1/xin[780] ) );
  DFF \modmult_1/xreg_reg[779]  ( .D(\modmult_1/xin[778] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[779]), .Q(\modmult_1/xin[779] ) );
  DFF \modmult_1/xreg_reg[778]  ( .D(\modmult_1/xin[777] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[778]), .Q(\modmult_1/xin[778] ) );
  DFF \modmult_1/xreg_reg[777]  ( .D(\modmult_1/xin[776] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[777]), .Q(\modmult_1/xin[777] ) );
  DFF \modmult_1/xreg_reg[776]  ( .D(\modmult_1/xin[775] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[776]), .Q(\modmult_1/xin[776] ) );
  DFF \modmult_1/xreg_reg[775]  ( .D(\modmult_1/xin[774] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[775]), .Q(\modmult_1/xin[775] ) );
  DFF \modmult_1/xreg_reg[774]  ( .D(\modmult_1/xin[773] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[774]), .Q(\modmult_1/xin[774] ) );
  DFF \modmult_1/xreg_reg[773]  ( .D(\modmult_1/xin[772] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[773]), .Q(\modmult_1/xin[773] ) );
  DFF \modmult_1/xreg_reg[772]  ( .D(\modmult_1/xin[771] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[772]), .Q(\modmult_1/xin[772] ) );
  DFF \modmult_1/xreg_reg[771]  ( .D(\modmult_1/xin[770] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[771]), .Q(\modmult_1/xin[771] ) );
  DFF \modmult_1/xreg_reg[770]  ( .D(\modmult_1/xin[769] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[770]), .Q(\modmult_1/xin[770] ) );
  DFF \modmult_1/xreg_reg[769]  ( .D(\modmult_1/xin[768] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[769]), .Q(\modmult_1/xin[769] ) );
  DFF \modmult_1/xreg_reg[768]  ( .D(\modmult_1/xin[767] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[768]), .Q(\modmult_1/xin[768] ) );
  DFF \modmult_1/xreg_reg[767]  ( .D(\modmult_1/xin[766] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[767]), .Q(\modmult_1/xin[767] ) );
  DFF \modmult_1/xreg_reg[766]  ( .D(\modmult_1/xin[765] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[766]), .Q(\modmult_1/xin[766] ) );
  DFF \modmult_1/xreg_reg[765]  ( .D(\modmult_1/xin[764] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[765]), .Q(\modmult_1/xin[765] ) );
  DFF \modmult_1/xreg_reg[764]  ( .D(\modmult_1/xin[763] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[764]), .Q(\modmult_1/xin[764] ) );
  DFF \modmult_1/xreg_reg[763]  ( .D(\modmult_1/xin[762] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[763]), .Q(\modmult_1/xin[763] ) );
  DFF \modmult_1/xreg_reg[762]  ( .D(\modmult_1/xin[761] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[762]), .Q(\modmult_1/xin[762] ) );
  DFF \modmult_1/xreg_reg[761]  ( .D(\modmult_1/xin[760] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[761]), .Q(\modmult_1/xin[761] ) );
  DFF \modmult_1/xreg_reg[760]  ( .D(\modmult_1/xin[759] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[760]), .Q(\modmult_1/xin[760] ) );
  DFF \modmult_1/xreg_reg[759]  ( .D(\modmult_1/xin[758] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[759]), .Q(\modmult_1/xin[759] ) );
  DFF \modmult_1/xreg_reg[758]  ( .D(\modmult_1/xin[757] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[758]), .Q(\modmult_1/xin[758] ) );
  DFF \modmult_1/xreg_reg[757]  ( .D(\modmult_1/xin[756] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[757]), .Q(\modmult_1/xin[757] ) );
  DFF \modmult_1/xreg_reg[756]  ( .D(\modmult_1/xin[755] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[756]), .Q(\modmult_1/xin[756] ) );
  DFF \modmult_1/xreg_reg[755]  ( .D(\modmult_1/xin[754] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[755]), .Q(\modmult_1/xin[755] ) );
  DFF \modmult_1/xreg_reg[754]  ( .D(\modmult_1/xin[753] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[754]), .Q(\modmult_1/xin[754] ) );
  DFF \modmult_1/xreg_reg[753]  ( .D(\modmult_1/xin[752] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[753]), .Q(\modmult_1/xin[753] ) );
  DFF \modmult_1/xreg_reg[752]  ( .D(\modmult_1/xin[751] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[752]), .Q(\modmult_1/xin[752] ) );
  DFF \modmult_1/xreg_reg[751]  ( .D(\modmult_1/xin[750] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[751]), .Q(\modmult_1/xin[751] ) );
  DFF \modmult_1/xreg_reg[750]  ( .D(\modmult_1/xin[749] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[750]), .Q(\modmult_1/xin[750] ) );
  DFF \modmult_1/xreg_reg[749]  ( .D(\modmult_1/xin[748] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[749]), .Q(\modmult_1/xin[749] ) );
  DFF \modmult_1/xreg_reg[748]  ( .D(\modmult_1/xin[747] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[748]), .Q(\modmult_1/xin[748] ) );
  DFF \modmult_1/xreg_reg[747]  ( .D(\modmult_1/xin[746] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[747]), .Q(\modmult_1/xin[747] ) );
  DFF \modmult_1/xreg_reg[746]  ( .D(\modmult_1/xin[745] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[746]), .Q(\modmult_1/xin[746] ) );
  DFF \modmult_1/xreg_reg[745]  ( .D(\modmult_1/xin[744] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[745]), .Q(\modmult_1/xin[745] ) );
  DFF \modmult_1/xreg_reg[744]  ( .D(\modmult_1/xin[743] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[744]), .Q(\modmult_1/xin[744] ) );
  DFF \modmult_1/xreg_reg[743]  ( .D(\modmult_1/xin[742] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[743]), .Q(\modmult_1/xin[743] ) );
  DFF \modmult_1/xreg_reg[742]  ( .D(\modmult_1/xin[741] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[742]), .Q(\modmult_1/xin[742] ) );
  DFF \modmult_1/xreg_reg[741]  ( .D(\modmult_1/xin[740] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[741]), .Q(\modmult_1/xin[741] ) );
  DFF \modmult_1/xreg_reg[740]  ( .D(\modmult_1/xin[739] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[740]), .Q(\modmult_1/xin[740] ) );
  DFF \modmult_1/xreg_reg[739]  ( .D(\modmult_1/xin[738] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[739]), .Q(\modmult_1/xin[739] ) );
  DFF \modmult_1/xreg_reg[738]  ( .D(\modmult_1/xin[737] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[738]), .Q(\modmult_1/xin[738] ) );
  DFF \modmult_1/xreg_reg[737]  ( .D(\modmult_1/xin[736] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[737]), .Q(\modmult_1/xin[737] ) );
  DFF \modmult_1/xreg_reg[736]  ( .D(\modmult_1/xin[735] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[736]), .Q(\modmult_1/xin[736] ) );
  DFF \modmult_1/xreg_reg[735]  ( .D(\modmult_1/xin[734] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[735]), .Q(\modmult_1/xin[735] ) );
  DFF \modmult_1/xreg_reg[734]  ( .D(\modmult_1/xin[733] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[734]), .Q(\modmult_1/xin[734] ) );
  DFF \modmult_1/xreg_reg[733]  ( .D(\modmult_1/xin[732] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[733]), .Q(\modmult_1/xin[733] ) );
  DFF \modmult_1/xreg_reg[732]  ( .D(\modmult_1/xin[731] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[732]), .Q(\modmult_1/xin[732] ) );
  DFF \modmult_1/xreg_reg[731]  ( .D(\modmult_1/xin[730] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[731]), .Q(\modmult_1/xin[731] ) );
  DFF \modmult_1/xreg_reg[730]  ( .D(\modmult_1/xin[729] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[730]), .Q(\modmult_1/xin[730] ) );
  DFF \modmult_1/xreg_reg[729]  ( .D(\modmult_1/xin[728] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[729]), .Q(\modmult_1/xin[729] ) );
  DFF \modmult_1/xreg_reg[728]  ( .D(\modmult_1/xin[727] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[728]), .Q(\modmult_1/xin[728] ) );
  DFF \modmult_1/xreg_reg[727]  ( .D(\modmult_1/xin[726] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[727]), .Q(\modmult_1/xin[727] ) );
  DFF \modmult_1/xreg_reg[726]  ( .D(\modmult_1/xin[725] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[726]), .Q(\modmult_1/xin[726] ) );
  DFF \modmult_1/xreg_reg[725]  ( .D(\modmult_1/xin[724] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[725]), .Q(\modmult_1/xin[725] ) );
  DFF \modmult_1/xreg_reg[724]  ( .D(\modmult_1/xin[723] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[724]), .Q(\modmult_1/xin[724] ) );
  DFF \modmult_1/xreg_reg[723]  ( .D(\modmult_1/xin[722] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[723]), .Q(\modmult_1/xin[723] ) );
  DFF \modmult_1/xreg_reg[722]  ( .D(\modmult_1/xin[721] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[722]), .Q(\modmult_1/xin[722] ) );
  DFF \modmult_1/xreg_reg[721]  ( .D(\modmult_1/xin[720] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[721]), .Q(\modmult_1/xin[721] ) );
  DFF \modmult_1/xreg_reg[720]  ( .D(\modmult_1/xin[719] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[720]), .Q(\modmult_1/xin[720] ) );
  DFF \modmult_1/xreg_reg[719]  ( .D(\modmult_1/xin[718] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[719]), .Q(\modmult_1/xin[719] ) );
  DFF \modmult_1/xreg_reg[718]  ( .D(\modmult_1/xin[717] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[718]), .Q(\modmult_1/xin[718] ) );
  DFF \modmult_1/xreg_reg[717]  ( .D(\modmult_1/xin[716] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[717]), .Q(\modmult_1/xin[717] ) );
  DFF \modmult_1/xreg_reg[716]  ( .D(\modmult_1/xin[715] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[716]), .Q(\modmult_1/xin[716] ) );
  DFF \modmult_1/xreg_reg[715]  ( .D(\modmult_1/xin[714] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[715]), .Q(\modmult_1/xin[715] ) );
  DFF \modmult_1/xreg_reg[714]  ( .D(\modmult_1/xin[713] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[714]), .Q(\modmult_1/xin[714] ) );
  DFF \modmult_1/xreg_reg[713]  ( .D(\modmult_1/xin[712] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[713]), .Q(\modmult_1/xin[713] ) );
  DFF \modmult_1/xreg_reg[712]  ( .D(\modmult_1/xin[711] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[712]), .Q(\modmult_1/xin[712] ) );
  DFF \modmult_1/xreg_reg[711]  ( .D(\modmult_1/xin[710] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[711]), .Q(\modmult_1/xin[711] ) );
  DFF \modmult_1/xreg_reg[710]  ( .D(\modmult_1/xin[709] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[710]), .Q(\modmult_1/xin[710] ) );
  DFF \modmult_1/xreg_reg[709]  ( .D(\modmult_1/xin[708] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[709]), .Q(\modmult_1/xin[709] ) );
  DFF \modmult_1/xreg_reg[708]  ( .D(\modmult_1/xin[707] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[708]), .Q(\modmult_1/xin[708] ) );
  DFF \modmult_1/xreg_reg[707]  ( .D(\modmult_1/xin[706] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[707]), .Q(\modmult_1/xin[707] ) );
  DFF \modmult_1/xreg_reg[706]  ( .D(\modmult_1/xin[705] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[706]), .Q(\modmult_1/xin[706] ) );
  DFF \modmult_1/xreg_reg[705]  ( .D(\modmult_1/xin[704] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[705]), .Q(\modmult_1/xin[705] ) );
  DFF \modmult_1/xreg_reg[704]  ( .D(\modmult_1/xin[703] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[704]), .Q(\modmult_1/xin[704] ) );
  DFF \modmult_1/xreg_reg[703]  ( .D(\modmult_1/xin[702] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[703]), .Q(\modmult_1/xin[703] ) );
  DFF \modmult_1/xreg_reg[702]  ( .D(\modmult_1/xin[701] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[702]), .Q(\modmult_1/xin[702] ) );
  DFF \modmult_1/xreg_reg[701]  ( .D(\modmult_1/xin[700] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[701]), .Q(\modmult_1/xin[701] ) );
  DFF \modmult_1/xreg_reg[700]  ( .D(\modmult_1/xin[699] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[700]), .Q(\modmult_1/xin[700] ) );
  DFF \modmult_1/xreg_reg[699]  ( .D(\modmult_1/xin[698] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[699]), .Q(\modmult_1/xin[699] ) );
  DFF \modmult_1/xreg_reg[698]  ( .D(\modmult_1/xin[697] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[698]), .Q(\modmult_1/xin[698] ) );
  DFF \modmult_1/xreg_reg[697]  ( .D(\modmult_1/xin[696] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[697]), .Q(\modmult_1/xin[697] ) );
  DFF \modmult_1/xreg_reg[696]  ( .D(\modmult_1/xin[695] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[696]), .Q(\modmult_1/xin[696] ) );
  DFF \modmult_1/xreg_reg[695]  ( .D(\modmult_1/xin[694] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[695]), .Q(\modmult_1/xin[695] ) );
  DFF \modmult_1/xreg_reg[694]  ( .D(\modmult_1/xin[693] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[694]), .Q(\modmult_1/xin[694] ) );
  DFF \modmult_1/xreg_reg[693]  ( .D(\modmult_1/xin[692] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[693]), .Q(\modmult_1/xin[693] ) );
  DFF \modmult_1/xreg_reg[692]  ( .D(\modmult_1/xin[691] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[692]), .Q(\modmult_1/xin[692] ) );
  DFF \modmult_1/xreg_reg[691]  ( .D(\modmult_1/xin[690] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[691]), .Q(\modmult_1/xin[691] ) );
  DFF \modmult_1/xreg_reg[690]  ( .D(\modmult_1/xin[689] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[690]), .Q(\modmult_1/xin[690] ) );
  DFF \modmult_1/xreg_reg[689]  ( .D(\modmult_1/xin[688] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[689]), .Q(\modmult_1/xin[689] ) );
  DFF \modmult_1/xreg_reg[688]  ( .D(\modmult_1/xin[687] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[688]), .Q(\modmult_1/xin[688] ) );
  DFF \modmult_1/xreg_reg[687]  ( .D(\modmult_1/xin[686] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[687]), .Q(\modmult_1/xin[687] ) );
  DFF \modmult_1/xreg_reg[686]  ( .D(\modmult_1/xin[685] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[686]), .Q(\modmult_1/xin[686] ) );
  DFF \modmult_1/xreg_reg[685]  ( .D(\modmult_1/xin[684] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[685]), .Q(\modmult_1/xin[685] ) );
  DFF \modmult_1/xreg_reg[684]  ( .D(\modmult_1/xin[683] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[684]), .Q(\modmult_1/xin[684] ) );
  DFF \modmult_1/xreg_reg[683]  ( .D(\modmult_1/xin[682] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[683]), .Q(\modmult_1/xin[683] ) );
  DFF \modmult_1/xreg_reg[682]  ( .D(\modmult_1/xin[681] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[682]), .Q(\modmult_1/xin[682] ) );
  DFF \modmult_1/xreg_reg[681]  ( .D(\modmult_1/xin[680] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[681]), .Q(\modmult_1/xin[681] ) );
  DFF \modmult_1/xreg_reg[680]  ( .D(\modmult_1/xin[679] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[680]), .Q(\modmult_1/xin[680] ) );
  DFF \modmult_1/xreg_reg[679]  ( .D(\modmult_1/xin[678] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[679]), .Q(\modmult_1/xin[679] ) );
  DFF \modmult_1/xreg_reg[678]  ( .D(\modmult_1/xin[677] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[678]), .Q(\modmult_1/xin[678] ) );
  DFF \modmult_1/xreg_reg[677]  ( .D(\modmult_1/xin[676] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[677]), .Q(\modmult_1/xin[677] ) );
  DFF \modmult_1/xreg_reg[676]  ( .D(\modmult_1/xin[675] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[676]), .Q(\modmult_1/xin[676] ) );
  DFF \modmult_1/xreg_reg[675]  ( .D(\modmult_1/xin[674] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[675]), .Q(\modmult_1/xin[675] ) );
  DFF \modmult_1/xreg_reg[674]  ( .D(\modmult_1/xin[673] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[674]), .Q(\modmult_1/xin[674] ) );
  DFF \modmult_1/xreg_reg[673]  ( .D(\modmult_1/xin[672] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[673]), .Q(\modmult_1/xin[673] ) );
  DFF \modmult_1/xreg_reg[672]  ( .D(\modmult_1/xin[671] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[672]), .Q(\modmult_1/xin[672] ) );
  DFF \modmult_1/xreg_reg[671]  ( .D(\modmult_1/xin[670] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[671]), .Q(\modmult_1/xin[671] ) );
  DFF \modmult_1/xreg_reg[670]  ( .D(\modmult_1/xin[669] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[670]), .Q(\modmult_1/xin[670] ) );
  DFF \modmult_1/xreg_reg[669]  ( .D(\modmult_1/xin[668] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[669]), .Q(\modmult_1/xin[669] ) );
  DFF \modmult_1/xreg_reg[668]  ( .D(\modmult_1/xin[667] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[668]), .Q(\modmult_1/xin[668] ) );
  DFF \modmult_1/xreg_reg[667]  ( .D(\modmult_1/xin[666] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[667]), .Q(\modmult_1/xin[667] ) );
  DFF \modmult_1/xreg_reg[666]  ( .D(\modmult_1/xin[665] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[666]), .Q(\modmult_1/xin[666] ) );
  DFF \modmult_1/xreg_reg[665]  ( .D(\modmult_1/xin[664] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[665]), .Q(\modmult_1/xin[665] ) );
  DFF \modmult_1/xreg_reg[664]  ( .D(\modmult_1/xin[663] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[664]), .Q(\modmult_1/xin[664] ) );
  DFF \modmult_1/xreg_reg[663]  ( .D(\modmult_1/xin[662] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[663]), .Q(\modmult_1/xin[663] ) );
  DFF \modmult_1/xreg_reg[662]  ( .D(\modmult_1/xin[661] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[662]), .Q(\modmult_1/xin[662] ) );
  DFF \modmult_1/xreg_reg[661]  ( .D(\modmult_1/xin[660] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[661]), .Q(\modmult_1/xin[661] ) );
  DFF \modmult_1/xreg_reg[660]  ( .D(\modmult_1/xin[659] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[660]), .Q(\modmult_1/xin[660] ) );
  DFF \modmult_1/xreg_reg[659]  ( .D(\modmult_1/xin[658] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[659]), .Q(\modmult_1/xin[659] ) );
  DFF \modmult_1/xreg_reg[658]  ( .D(\modmult_1/xin[657] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[658]), .Q(\modmult_1/xin[658] ) );
  DFF \modmult_1/xreg_reg[657]  ( .D(\modmult_1/xin[656] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[657]), .Q(\modmult_1/xin[657] ) );
  DFF \modmult_1/xreg_reg[656]  ( .D(\modmult_1/xin[655] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[656]), .Q(\modmult_1/xin[656] ) );
  DFF \modmult_1/xreg_reg[655]  ( .D(\modmult_1/xin[654] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[655]), .Q(\modmult_1/xin[655] ) );
  DFF \modmult_1/xreg_reg[654]  ( .D(\modmult_1/xin[653] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[654]), .Q(\modmult_1/xin[654] ) );
  DFF \modmult_1/xreg_reg[653]  ( .D(\modmult_1/xin[652] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[653]), .Q(\modmult_1/xin[653] ) );
  DFF \modmult_1/xreg_reg[652]  ( .D(\modmult_1/xin[651] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[652]), .Q(\modmult_1/xin[652] ) );
  DFF \modmult_1/xreg_reg[651]  ( .D(\modmult_1/xin[650] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[651]), .Q(\modmult_1/xin[651] ) );
  DFF \modmult_1/xreg_reg[650]  ( .D(\modmult_1/xin[649] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[650]), .Q(\modmult_1/xin[650] ) );
  DFF \modmult_1/xreg_reg[649]  ( .D(\modmult_1/xin[648] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[649]), .Q(\modmult_1/xin[649] ) );
  DFF \modmult_1/xreg_reg[648]  ( .D(\modmult_1/xin[647] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[648]), .Q(\modmult_1/xin[648] ) );
  DFF \modmult_1/xreg_reg[647]  ( .D(\modmult_1/xin[646] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[647]), .Q(\modmult_1/xin[647] ) );
  DFF \modmult_1/xreg_reg[646]  ( .D(\modmult_1/xin[645] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[646]), .Q(\modmult_1/xin[646] ) );
  DFF \modmult_1/xreg_reg[645]  ( .D(\modmult_1/xin[644] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[645]), .Q(\modmult_1/xin[645] ) );
  DFF \modmult_1/xreg_reg[644]  ( .D(\modmult_1/xin[643] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[644]), .Q(\modmult_1/xin[644] ) );
  DFF \modmult_1/xreg_reg[643]  ( .D(\modmult_1/xin[642] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[643]), .Q(\modmult_1/xin[643] ) );
  DFF \modmult_1/xreg_reg[642]  ( .D(\modmult_1/xin[641] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[642]), .Q(\modmult_1/xin[642] ) );
  DFF \modmult_1/xreg_reg[641]  ( .D(\modmult_1/xin[640] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[641]), .Q(\modmult_1/xin[641] ) );
  DFF \modmult_1/xreg_reg[640]  ( .D(\modmult_1/xin[639] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[640]), .Q(\modmult_1/xin[640] ) );
  DFF \modmult_1/xreg_reg[639]  ( .D(\modmult_1/xin[638] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[639]), .Q(\modmult_1/xin[639] ) );
  DFF \modmult_1/xreg_reg[638]  ( .D(\modmult_1/xin[637] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[638]), .Q(\modmult_1/xin[638] ) );
  DFF \modmult_1/xreg_reg[637]  ( .D(\modmult_1/xin[636] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[637]), .Q(\modmult_1/xin[637] ) );
  DFF \modmult_1/xreg_reg[636]  ( .D(\modmult_1/xin[635] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[636]), .Q(\modmult_1/xin[636] ) );
  DFF \modmult_1/xreg_reg[635]  ( .D(\modmult_1/xin[634] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[635]), .Q(\modmult_1/xin[635] ) );
  DFF \modmult_1/xreg_reg[634]  ( .D(\modmult_1/xin[633] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[634]), .Q(\modmult_1/xin[634] ) );
  DFF \modmult_1/xreg_reg[633]  ( .D(\modmult_1/xin[632] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[633]), .Q(\modmult_1/xin[633] ) );
  DFF \modmult_1/xreg_reg[632]  ( .D(\modmult_1/xin[631] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[632]), .Q(\modmult_1/xin[632] ) );
  DFF \modmult_1/xreg_reg[631]  ( .D(\modmult_1/xin[630] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[631]), .Q(\modmult_1/xin[631] ) );
  DFF \modmult_1/xreg_reg[630]  ( .D(\modmult_1/xin[629] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[630]), .Q(\modmult_1/xin[630] ) );
  DFF \modmult_1/xreg_reg[629]  ( .D(\modmult_1/xin[628] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[629]), .Q(\modmult_1/xin[629] ) );
  DFF \modmult_1/xreg_reg[628]  ( .D(\modmult_1/xin[627] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[628]), .Q(\modmult_1/xin[628] ) );
  DFF \modmult_1/xreg_reg[627]  ( .D(\modmult_1/xin[626] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[627]), .Q(\modmult_1/xin[627] ) );
  DFF \modmult_1/xreg_reg[626]  ( .D(\modmult_1/xin[625] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[626]), .Q(\modmult_1/xin[626] ) );
  DFF \modmult_1/xreg_reg[625]  ( .D(\modmult_1/xin[624] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[625]), .Q(\modmult_1/xin[625] ) );
  DFF \modmult_1/xreg_reg[624]  ( .D(\modmult_1/xin[623] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[624]), .Q(\modmult_1/xin[624] ) );
  DFF \modmult_1/xreg_reg[623]  ( .D(\modmult_1/xin[622] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[623]), .Q(\modmult_1/xin[623] ) );
  DFF \modmult_1/xreg_reg[622]  ( .D(\modmult_1/xin[621] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[622]), .Q(\modmult_1/xin[622] ) );
  DFF \modmult_1/xreg_reg[621]  ( .D(\modmult_1/xin[620] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[621]), .Q(\modmult_1/xin[621] ) );
  DFF \modmult_1/xreg_reg[620]  ( .D(\modmult_1/xin[619] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[620]), .Q(\modmult_1/xin[620] ) );
  DFF \modmult_1/xreg_reg[619]  ( .D(\modmult_1/xin[618] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[619]), .Q(\modmult_1/xin[619] ) );
  DFF \modmult_1/xreg_reg[618]  ( .D(\modmult_1/xin[617] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[618]), .Q(\modmult_1/xin[618] ) );
  DFF \modmult_1/xreg_reg[617]  ( .D(\modmult_1/xin[616] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[617]), .Q(\modmult_1/xin[617] ) );
  DFF \modmult_1/xreg_reg[616]  ( .D(\modmult_1/xin[615] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[616]), .Q(\modmult_1/xin[616] ) );
  DFF \modmult_1/xreg_reg[615]  ( .D(\modmult_1/xin[614] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[615]), .Q(\modmult_1/xin[615] ) );
  DFF \modmult_1/xreg_reg[614]  ( .D(\modmult_1/xin[613] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[614]), .Q(\modmult_1/xin[614] ) );
  DFF \modmult_1/xreg_reg[613]  ( .D(\modmult_1/xin[612] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[613]), .Q(\modmult_1/xin[613] ) );
  DFF \modmult_1/xreg_reg[612]  ( .D(\modmult_1/xin[611] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[612]), .Q(\modmult_1/xin[612] ) );
  DFF \modmult_1/xreg_reg[611]  ( .D(\modmult_1/xin[610] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[611]), .Q(\modmult_1/xin[611] ) );
  DFF \modmult_1/xreg_reg[610]  ( .D(\modmult_1/xin[609] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[610]), .Q(\modmult_1/xin[610] ) );
  DFF \modmult_1/xreg_reg[609]  ( .D(\modmult_1/xin[608] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[609]), .Q(\modmult_1/xin[609] ) );
  DFF \modmult_1/xreg_reg[608]  ( .D(\modmult_1/xin[607] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[608]), .Q(\modmult_1/xin[608] ) );
  DFF \modmult_1/xreg_reg[607]  ( .D(\modmult_1/xin[606] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[607]), .Q(\modmult_1/xin[607] ) );
  DFF \modmult_1/xreg_reg[606]  ( .D(\modmult_1/xin[605] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[606]), .Q(\modmult_1/xin[606] ) );
  DFF \modmult_1/xreg_reg[605]  ( .D(\modmult_1/xin[604] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[605]), .Q(\modmult_1/xin[605] ) );
  DFF \modmult_1/xreg_reg[604]  ( .D(\modmult_1/xin[603] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[604]), .Q(\modmult_1/xin[604] ) );
  DFF \modmult_1/xreg_reg[603]  ( .D(\modmult_1/xin[602] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[603]), .Q(\modmult_1/xin[603] ) );
  DFF \modmult_1/xreg_reg[602]  ( .D(\modmult_1/xin[601] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[602]), .Q(\modmult_1/xin[602] ) );
  DFF \modmult_1/xreg_reg[601]  ( .D(\modmult_1/xin[600] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[601]), .Q(\modmult_1/xin[601] ) );
  DFF \modmult_1/xreg_reg[600]  ( .D(\modmult_1/xin[599] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[600]), .Q(\modmult_1/xin[600] ) );
  DFF \modmult_1/xreg_reg[599]  ( .D(\modmult_1/xin[598] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[599]), .Q(\modmult_1/xin[599] ) );
  DFF \modmult_1/xreg_reg[598]  ( .D(\modmult_1/xin[597] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[598]), .Q(\modmult_1/xin[598] ) );
  DFF \modmult_1/xreg_reg[597]  ( .D(\modmult_1/xin[596] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[597]), .Q(\modmult_1/xin[597] ) );
  DFF \modmult_1/xreg_reg[596]  ( .D(\modmult_1/xin[595] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[596]), .Q(\modmult_1/xin[596] ) );
  DFF \modmult_1/xreg_reg[595]  ( .D(\modmult_1/xin[594] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[595]), .Q(\modmult_1/xin[595] ) );
  DFF \modmult_1/xreg_reg[594]  ( .D(\modmult_1/xin[593] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[594]), .Q(\modmult_1/xin[594] ) );
  DFF \modmult_1/xreg_reg[593]  ( .D(\modmult_1/xin[592] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[593]), .Q(\modmult_1/xin[593] ) );
  DFF \modmult_1/xreg_reg[592]  ( .D(\modmult_1/xin[591] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[592]), .Q(\modmult_1/xin[592] ) );
  DFF \modmult_1/xreg_reg[591]  ( .D(\modmult_1/xin[590] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[591]), .Q(\modmult_1/xin[591] ) );
  DFF \modmult_1/xreg_reg[590]  ( .D(\modmult_1/xin[589] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[590]), .Q(\modmult_1/xin[590] ) );
  DFF \modmult_1/xreg_reg[589]  ( .D(\modmult_1/xin[588] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[589]), .Q(\modmult_1/xin[589] ) );
  DFF \modmult_1/xreg_reg[588]  ( .D(\modmult_1/xin[587] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[588]), .Q(\modmult_1/xin[588] ) );
  DFF \modmult_1/xreg_reg[587]  ( .D(\modmult_1/xin[586] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[587]), .Q(\modmult_1/xin[587] ) );
  DFF \modmult_1/xreg_reg[586]  ( .D(\modmult_1/xin[585] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[586]), .Q(\modmult_1/xin[586] ) );
  DFF \modmult_1/xreg_reg[585]  ( .D(\modmult_1/xin[584] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[585]), .Q(\modmult_1/xin[585] ) );
  DFF \modmult_1/xreg_reg[584]  ( .D(\modmult_1/xin[583] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[584]), .Q(\modmult_1/xin[584] ) );
  DFF \modmult_1/xreg_reg[583]  ( .D(\modmult_1/xin[582] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[583]), .Q(\modmult_1/xin[583] ) );
  DFF \modmult_1/xreg_reg[582]  ( .D(\modmult_1/xin[581] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[582]), .Q(\modmult_1/xin[582] ) );
  DFF \modmult_1/xreg_reg[581]  ( .D(\modmult_1/xin[580] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[581]), .Q(\modmult_1/xin[581] ) );
  DFF \modmult_1/xreg_reg[580]  ( .D(\modmult_1/xin[579] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[580]), .Q(\modmult_1/xin[580] ) );
  DFF \modmult_1/xreg_reg[579]  ( .D(\modmult_1/xin[578] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[579]), .Q(\modmult_1/xin[579] ) );
  DFF \modmult_1/xreg_reg[578]  ( .D(\modmult_1/xin[577] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[578]), .Q(\modmult_1/xin[578] ) );
  DFF \modmult_1/xreg_reg[577]  ( .D(\modmult_1/xin[576] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[577]), .Q(\modmult_1/xin[577] ) );
  DFF \modmult_1/xreg_reg[576]  ( .D(\modmult_1/xin[575] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[576]), .Q(\modmult_1/xin[576] ) );
  DFF \modmult_1/xreg_reg[575]  ( .D(\modmult_1/xin[574] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[575]), .Q(\modmult_1/xin[575] ) );
  DFF \modmult_1/xreg_reg[574]  ( .D(\modmult_1/xin[573] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[574]), .Q(\modmult_1/xin[574] ) );
  DFF \modmult_1/xreg_reg[573]  ( .D(\modmult_1/xin[572] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[573]), .Q(\modmult_1/xin[573] ) );
  DFF \modmult_1/xreg_reg[572]  ( .D(\modmult_1/xin[571] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[572]), .Q(\modmult_1/xin[572] ) );
  DFF \modmult_1/xreg_reg[571]  ( .D(\modmult_1/xin[570] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[571]), .Q(\modmult_1/xin[571] ) );
  DFF \modmult_1/xreg_reg[570]  ( .D(\modmult_1/xin[569] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[570]), .Q(\modmult_1/xin[570] ) );
  DFF \modmult_1/xreg_reg[569]  ( .D(\modmult_1/xin[568] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[569]), .Q(\modmult_1/xin[569] ) );
  DFF \modmult_1/xreg_reg[568]  ( .D(\modmult_1/xin[567] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[568]), .Q(\modmult_1/xin[568] ) );
  DFF \modmult_1/xreg_reg[567]  ( .D(\modmult_1/xin[566] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[567]), .Q(\modmult_1/xin[567] ) );
  DFF \modmult_1/xreg_reg[566]  ( .D(\modmult_1/xin[565] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[566]), .Q(\modmult_1/xin[566] ) );
  DFF \modmult_1/xreg_reg[565]  ( .D(\modmult_1/xin[564] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[565]), .Q(\modmult_1/xin[565] ) );
  DFF \modmult_1/xreg_reg[564]  ( .D(\modmult_1/xin[563] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[564]), .Q(\modmult_1/xin[564] ) );
  DFF \modmult_1/xreg_reg[563]  ( .D(\modmult_1/xin[562] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[563]), .Q(\modmult_1/xin[563] ) );
  DFF \modmult_1/xreg_reg[562]  ( .D(\modmult_1/xin[561] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[562]), .Q(\modmult_1/xin[562] ) );
  DFF \modmult_1/xreg_reg[561]  ( .D(\modmult_1/xin[560] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[561]), .Q(\modmult_1/xin[561] ) );
  DFF \modmult_1/xreg_reg[560]  ( .D(\modmult_1/xin[559] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[560]), .Q(\modmult_1/xin[560] ) );
  DFF \modmult_1/xreg_reg[559]  ( .D(\modmult_1/xin[558] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[559]), .Q(\modmult_1/xin[559] ) );
  DFF \modmult_1/xreg_reg[558]  ( .D(\modmult_1/xin[557] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[558]), .Q(\modmult_1/xin[558] ) );
  DFF \modmult_1/xreg_reg[557]  ( .D(\modmult_1/xin[556] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[557]), .Q(\modmult_1/xin[557] ) );
  DFF \modmult_1/xreg_reg[556]  ( .D(\modmult_1/xin[555] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[556]), .Q(\modmult_1/xin[556] ) );
  DFF \modmult_1/xreg_reg[555]  ( .D(\modmult_1/xin[554] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[555]), .Q(\modmult_1/xin[555] ) );
  DFF \modmult_1/xreg_reg[554]  ( .D(\modmult_1/xin[553] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[554]), .Q(\modmult_1/xin[554] ) );
  DFF \modmult_1/xreg_reg[553]  ( .D(\modmult_1/xin[552] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[553]), .Q(\modmult_1/xin[553] ) );
  DFF \modmult_1/xreg_reg[552]  ( .D(\modmult_1/xin[551] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[552]), .Q(\modmult_1/xin[552] ) );
  DFF \modmult_1/xreg_reg[551]  ( .D(\modmult_1/xin[550] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[551]), .Q(\modmult_1/xin[551] ) );
  DFF \modmult_1/xreg_reg[550]  ( .D(\modmult_1/xin[549] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[550]), .Q(\modmult_1/xin[550] ) );
  DFF \modmult_1/xreg_reg[549]  ( .D(\modmult_1/xin[548] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[549]), .Q(\modmult_1/xin[549] ) );
  DFF \modmult_1/xreg_reg[548]  ( .D(\modmult_1/xin[547] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[548]), .Q(\modmult_1/xin[548] ) );
  DFF \modmult_1/xreg_reg[547]  ( .D(\modmult_1/xin[546] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[547]), .Q(\modmult_1/xin[547] ) );
  DFF \modmult_1/xreg_reg[546]  ( .D(\modmult_1/xin[545] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[546]), .Q(\modmult_1/xin[546] ) );
  DFF \modmult_1/xreg_reg[545]  ( .D(\modmult_1/xin[544] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[545]), .Q(\modmult_1/xin[545] ) );
  DFF \modmult_1/xreg_reg[544]  ( .D(\modmult_1/xin[543] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[544]), .Q(\modmult_1/xin[544] ) );
  DFF \modmult_1/xreg_reg[543]  ( .D(\modmult_1/xin[542] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[543]), .Q(\modmult_1/xin[543] ) );
  DFF \modmult_1/xreg_reg[542]  ( .D(\modmult_1/xin[541] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[542]), .Q(\modmult_1/xin[542] ) );
  DFF \modmult_1/xreg_reg[541]  ( .D(\modmult_1/xin[540] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[541]), .Q(\modmult_1/xin[541] ) );
  DFF \modmult_1/xreg_reg[540]  ( .D(\modmult_1/xin[539] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[540]), .Q(\modmult_1/xin[540] ) );
  DFF \modmult_1/xreg_reg[539]  ( .D(\modmult_1/xin[538] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[539]), .Q(\modmult_1/xin[539] ) );
  DFF \modmult_1/xreg_reg[538]  ( .D(\modmult_1/xin[537] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[538]), .Q(\modmult_1/xin[538] ) );
  DFF \modmult_1/xreg_reg[537]  ( .D(\modmult_1/xin[536] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[537]), .Q(\modmult_1/xin[537] ) );
  DFF \modmult_1/xreg_reg[536]  ( .D(\modmult_1/xin[535] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[536]), .Q(\modmult_1/xin[536] ) );
  DFF \modmult_1/xreg_reg[535]  ( .D(\modmult_1/xin[534] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[535]), .Q(\modmult_1/xin[535] ) );
  DFF \modmult_1/xreg_reg[534]  ( .D(\modmult_1/xin[533] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[534]), .Q(\modmult_1/xin[534] ) );
  DFF \modmult_1/xreg_reg[533]  ( .D(\modmult_1/xin[532] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[533]), .Q(\modmult_1/xin[533] ) );
  DFF \modmult_1/xreg_reg[532]  ( .D(\modmult_1/xin[531] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[532]), .Q(\modmult_1/xin[532] ) );
  DFF \modmult_1/xreg_reg[531]  ( .D(\modmult_1/xin[530] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[531]), .Q(\modmult_1/xin[531] ) );
  DFF \modmult_1/xreg_reg[530]  ( .D(\modmult_1/xin[529] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[530]), .Q(\modmult_1/xin[530] ) );
  DFF \modmult_1/xreg_reg[529]  ( .D(\modmult_1/xin[528] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[529]), .Q(\modmult_1/xin[529] ) );
  DFF \modmult_1/xreg_reg[528]  ( .D(\modmult_1/xin[527] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[528]), .Q(\modmult_1/xin[528] ) );
  DFF \modmult_1/xreg_reg[527]  ( .D(\modmult_1/xin[526] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[527]), .Q(\modmult_1/xin[527] ) );
  DFF \modmult_1/xreg_reg[526]  ( .D(\modmult_1/xin[525] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[526]), .Q(\modmult_1/xin[526] ) );
  DFF \modmult_1/xreg_reg[525]  ( .D(\modmult_1/xin[524] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[525]), .Q(\modmult_1/xin[525] ) );
  DFF \modmult_1/xreg_reg[524]  ( .D(\modmult_1/xin[523] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[524]), .Q(\modmult_1/xin[524] ) );
  DFF \modmult_1/xreg_reg[523]  ( .D(\modmult_1/xin[522] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[523]), .Q(\modmult_1/xin[523] ) );
  DFF \modmult_1/xreg_reg[522]  ( .D(\modmult_1/xin[521] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[522]), .Q(\modmult_1/xin[522] ) );
  DFF \modmult_1/xreg_reg[521]  ( .D(\modmult_1/xin[520] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[521]), .Q(\modmult_1/xin[521] ) );
  DFF \modmult_1/xreg_reg[520]  ( .D(\modmult_1/xin[519] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[520]), .Q(\modmult_1/xin[520] ) );
  DFF \modmult_1/xreg_reg[519]  ( .D(\modmult_1/xin[518] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[519]), .Q(\modmult_1/xin[519] ) );
  DFF \modmult_1/xreg_reg[518]  ( .D(\modmult_1/xin[517] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[518]), .Q(\modmult_1/xin[518] ) );
  DFF \modmult_1/xreg_reg[517]  ( .D(\modmult_1/xin[516] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[517]), .Q(\modmult_1/xin[517] ) );
  DFF \modmult_1/xreg_reg[516]  ( .D(\modmult_1/xin[515] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[516]), .Q(\modmult_1/xin[516] ) );
  DFF \modmult_1/xreg_reg[515]  ( .D(\modmult_1/xin[514] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[515]), .Q(\modmult_1/xin[515] ) );
  DFF \modmult_1/xreg_reg[514]  ( .D(\modmult_1/xin[513] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[514]), .Q(\modmult_1/xin[514] ) );
  DFF \modmult_1/xreg_reg[513]  ( .D(\modmult_1/xin[512] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[513]), .Q(\modmult_1/xin[513] ) );
  DFF \modmult_1/xreg_reg[512]  ( .D(\modmult_1/xin[511] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[512]), .Q(\modmult_1/xin[512] ) );
  DFF \modmult_1/xreg_reg[511]  ( .D(\modmult_1/xin[510] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[511]), .Q(\modmult_1/xin[511] ) );
  DFF \modmult_1/xreg_reg[510]  ( .D(\modmult_1/xin[509] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[510]), .Q(\modmult_1/xin[510] ) );
  DFF \modmult_1/xreg_reg[509]  ( .D(\modmult_1/xin[508] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[509]), .Q(\modmult_1/xin[509] ) );
  DFF \modmult_1/xreg_reg[508]  ( .D(\modmult_1/xin[507] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[508]), .Q(\modmult_1/xin[508] ) );
  DFF \modmult_1/xreg_reg[507]  ( .D(\modmult_1/xin[506] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[507]), .Q(\modmult_1/xin[507] ) );
  DFF \modmult_1/xreg_reg[506]  ( .D(\modmult_1/xin[505] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[506]), .Q(\modmult_1/xin[506] ) );
  DFF \modmult_1/xreg_reg[505]  ( .D(\modmult_1/xin[504] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[505]), .Q(\modmult_1/xin[505] ) );
  DFF \modmult_1/xreg_reg[504]  ( .D(\modmult_1/xin[503] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[504]), .Q(\modmult_1/xin[504] ) );
  DFF \modmult_1/xreg_reg[503]  ( .D(\modmult_1/xin[502] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[503]), .Q(\modmult_1/xin[503] ) );
  DFF \modmult_1/xreg_reg[502]  ( .D(\modmult_1/xin[501] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[502]), .Q(\modmult_1/xin[502] ) );
  DFF \modmult_1/xreg_reg[501]  ( .D(\modmult_1/xin[500] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[501]), .Q(\modmult_1/xin[501] ) );
  DFF \modmult_1/xreg_reg[500]  ( .D(\modmult_1/xin[499] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[500]), .Q(\modmult_1/xin[500] ) );
  DFF \modmult_1/xreg_reg[499]  ( .D(\modmult_1/xin[498] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[499]), .Q(\modmult_1/xin[499] ) );
  DFF \modmult_1/xreg_reg[498]  ( .D(\modmult_1/xin[497] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[498]), .Q(\modmult_1/xin[498] ) );
  DFF \modmult_1/xreg_reg[497]  ( .D(\modmult_1/xin[496] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[497]), .Q(\modmult_1/xin[497] ) );
  DFF \modmult_1/xreg_reg[496]  ( .D(\modmult_1/xin[495] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[496]), .Q(\modmult_1/xin[496] ) );
  DFF \modmult_1/xreg_reg[495]  ( .D(\modmult_1/xin[494] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[495]), .Q(\modmult_1/xin[495] ) );
  DFF \modmult_1/xreg_reg[494]  ( .D(\modmult_1/xin[493] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[494]), .Q(\modmult_1/xin[494] ) );
  DFF \modmult_1/xreg_reg[493]  ( .D(\modmult_1/xin[492] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[493]), .Q(\modmult_1/xin[493] ) );
  DFF \modmult_1/xreg_reg[492]  ( .D(\modmult_1/xin[491] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[492]), .Q(\modmult_1/xin[492] ) );
  DFF \modmult_1/xreg_reg[491]  ( .D(\modmult_1/xin[490] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[491]), .Q(\modmult_1/xin[491] ) );
  DFF \modmult_1/xreg_reg[490]  ( .D(\modmult_1/xin[489] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[490]), .Q(\modmult_1/xin[490] ) );
  DFF \modmult_1/xreg_reg[489]  ( .D(\modmult_1/xin[488] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[489]), .Q(\modmult_1/xin[489] ) );
  DFF \modmult_1/xreg_reg[488]  ( .D(\modmult_1/xin[487] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[488]), .Q(\modmult_1/xin[488] ) );
  DFF \modmult_1/xreg_reg[487]  ( .D(\modmult_1/xin[486] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[487]), .Q(\modmult_1/xin[487] ) );
  DFF \modmult_1/xreg_reg[486]  ( .D(\modmult_1/xin[485] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[486]), .Q(\modmult_1/xin[486] ) );
  DFF \modmult_1/xreg_reg[485]  ( .D(\modmult_1/xin[484] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[485]), .Q(\modmult_1/xin[485] ) );
  DFF \modmult_1/xreg_reg[484]  ( .D(\modmult_1/xin[483] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[484]), .Q(\modmult_1/xin[484] ) );
  DFF \modmult_1/xreg_reg[483]  ( .D(\modmult_1/xin[482] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[483]), .Q(\modmult_1/xin[483] ) );
  DFF \modmult_1/xreg_reg[482]  ( .D(\modmult_1/xin[481] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[482]), .Q(\modmult_1/xin[482] ) );
  DFF \modmult_1/xreg_reg[481]  ( .D(\modmult_1/xin[480] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[481]), .Q(\modmult_1/xin[481] ) );
  DFF \modmult_1/xreg_reg[480]  ( .D(\modmult_1/xin[479] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[480]), .Q(\modmult_1/xin[480] ) );
  DFF \modmult_1/xreg_reg[479]  ( .D(\modmult_1/xin[478] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[479]), .Q(\modmult_1/xin[479] ) );
  DFF \modmult_1/xreg_reg[478]  ( .D(\modmult_1/xin[477] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[478]), .Q(\modmult_1/xin[478] ) );
  DFF \modmult_1/xreg_reg[477]  ( .D(\modmult_1/xin[476] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[477]), .Q(\modmult_1/xin[477] ) );
  DFF \modmult_1/xreg_reg[476]  ( .D(\modmult_1/xin[475] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[476]), .Q(\modmult_1/xin[476] ) );
  DFF \modmult_1/xreg_reg[475]  ( .D(\modmult_1/xin[474] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[475]), .Q(\modmult_1/xin[475] ) );
  DFF \modmult_1/xreg_reg[474]  ( .D(\modmult_1/xin[473] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[474]), .Q(\modmult_1/xin[474] ) );
  DFF \modmult_1/xreg_reg[473]  ( .D(\modmult_1/xin[472] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[473]), .Q(\modmult_1/xin[473] ) );
  DFF \modmult_1/xreg_reg[472]  ( .D(\modmult_1/xin[471] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[472]), .Q(\modmult_1/xin[472] ) );
  DFF \modmult_1/xreg_reg[471]  ( .D(\modmult_1/xin[470] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[471]), .Q(\modmult_1/xin[471] ) );
  DFF \modmult_1/xreg_reg[470]  ( .D(\modmult_1/xin[469] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[470]), .Q(\modmult_1/xin[470] ) );
  DFF \modmult_1/xreg_reg[469]  ( .D(\modmult_1/xin[468] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[469]), .Q(\modmult_1/xin[469] ) );
  DFF \modmult_1/xreg_reg[468]  ( .D(\modmult_1/xin[467] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[468]), .Q(\modmult_1/xin[468] ) );
  DFF \modmult_1/xreg_reg[467]  ( .D(\modmult_1/xin[466] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[467]), .Q(\modmult_1/xin[467] ) );
  DFF \modmult_1/xreg_reg[466]  ( .D(\modmult_1/xin[465] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[466]), .Q(\modmult_1/xin[466] ) );
  DFF \modmult_1/xreg_reg[465]  ( .D(\modmult_1/xin[464] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[465]), .Q(\modmult_1/xin[465] ) );
  DFF \modmult_1/xreg_reg[464]  ( .D(\modmult_1/xin[463] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[464]), .Q(\modmult_1/xin[464] ) );
  DFF \modmult_1/xreg_reg[463]  ( .D(\modmult_1/xin[462] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[463]), .Q(\modmult_1/xin[463] ) );
  DFF \modmult_1/xreg_reg[462]  ( .D(\modmult_1/xin[461] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[462]), .Q(\modmult_1/xin[462] ) );
  DFF \modmult_1/xreg_reg[461]  ( .D(\modmult_1/xin[460] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[461]), .Q(\modmult_1/xin[461] ) );
  DFF \modmult_1/xreg_reg[460]  ( .D(\modmult_1/xin[459] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[460]), .Q(\modmult_1/xin[460] ) );
  DFF \modmult_1/xreg_reg[459]  ( .D(\modmult_1/xin[458] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[459]), .Q(\modmult_1/xin[459] ) );
  DFF \modmult_1/xreg_reg[458]  ( .D(\modmult_1/xin[457] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[458]), .Q(\modmult_1/xin[458] ) );
  DFF \modmult_1/xreg_reg[457]  ( .D(\modmult_1/xin[456] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[457]), .Q(\modmult_1/xin[457] ) );
  DFF \modmult_1/xreg_reg[456]  ( .D(\modmult_1/xin[455] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[456]), .Q(\modmult_1/xin[456] ) );
  DFF \modmult_1/xreg_reg[455]  ( .D(\modmult_1/xin[454] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[455]), .Q(\modmult_1/xin[455] ) );
  DFF \modmult_1/xreg_reg[454]  ( .D(\modmult_1/xin[453] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[454]), .Q(\modmult_1/xin[454] ) );
  DFF \modmult_1/xreg_reg[453]  ( .D(\modmult_1/xin[452] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[453]), .Q(\modmult_1/xin[453] ) );
  DFF \modmult_1/xreg_reg[452]  ( .D(\modmult_1/xin[451] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[452]), .Q(\modmult_1/xin[452] ) );
  DFF \modmult_1/xreg_reg[451]  ( .D(\modmult_1/xin[450] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[451]), .Q(\modmult_1/xin[451] ) );
  DFF \modmult_1/xreg_reg[450]  ( .D(\modmult_1/xin[449] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[450]), .Q(\modmult_1/xin[450] ) );
  DFF \modmult_1/xreg_reg[449]  ( .D(\modmult_1/xin[448] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[449]), .Q(\modmult_1/xin[449] ) );
  DFF \modmult_1/xreg_reg[448]  ( .D(\modmult_1/xin[447] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[448]), .Q(\modmult_1/xin[448] ) );
  DFF \modmult_1/xreg_reg[447]  ( .D(\modmult_1/xin[446] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[447]), .Q(\modmult_1/xin[447] ) );
  DFF \modmult_1/xreg_reg[446]  ( .D(\modmult_1/xin[445] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[446]), .Q(\modmult_1/xin[446] ) );
  DFF \modmult_1/xreg_reg[445]  ( .D(\modmult_1/xin[444] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[445]), .Q(\modmult_1/xin[445] ) );
  DFF \modmult_1/xreg_reg[444]  ( .D(\modmult_1/xin[443] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[444]), .Q(\modmult_1/xin[444] ) );
  DFF \modmult_1/xreg_reg[443]  ( .D(\modmult_1/xin[442] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[443]), .Q(\modmult_1/xin[443] ) );
  DFF \modmult_1/xreg_reg[442]  ( .D(\modmult_1/xin[441] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[442]), .Q(\modmult_1/xin[442] ) );
  DFF \modmult_1/xreg_reg[441]  ( .D(\modmult_1/xin[440] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[441]), .Q(\modmult_1/xin[441] ) );
  DFF \modmult_1/xreg_reg[440]  ( .D(\modmult_1/xin[439] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[440]), .Q(\modmult_1/xin[440] ) );
  DFF \modmult_1/xreg_reg[439]  ( .D(\modmult_1/xin[438] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[439]), .Q(\modmult_1/xin[439] ) );
  DFF \modmult_1/xreg_reg[438]  ( .D(\modmult_1/xin[437] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[438]), .Q(\modmult_1/xin[438] ) );
  DFF \modmult_1/xreg_reg[437]  ( .D(\modmult_1/xin[436] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[437]), .Q(\modmult_1/xin[437] ) );
  DFF \modmult_1/xreg_reg[436]  ( .D(\modmult_1/xin[435] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[436]), .Q(\modmult_1/xin[436] ) );
  DFF \modmult_1/xreg_reg[435]  ( .D(\modmult_1/xin[434] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[435]), .Q(\modmult_1/xin[435] ) );
  DFF \modmult_1/xreg_reg[434]  ( .D(\modmult_1/xin[433] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[434]), .Q(\modmult_1/xin[434] ) );
  DFF \modmult_1/xreg_reg[433]  ( .D(\modmult_1/xin[432] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[433]), .Q(\modmult_1/xin[433] ) );
  DFF \modmult_1/xreg_reg[432]  ( .D(\modmult_1/xin[431] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[432]), .Q(\modmult_1/xin[432] ) );
  DFF \modmult_1/xreg_reg[431]  ( .D(\modmult_1/xin[430] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[431]), .Q(\modmult_1/xin[431] ) );
  DFF \modmult_1/xreg_reg[430]  ( .D(\modmult_1/xin[429] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[430]), .Q(\modmult_1/xin[430] ) );
  DFF \modmult_1/xreg_reg[429]  ( .D(\modmult_1/xin[428] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[429]), .Q(\modmult_1/xin[429] ) );
  DFF \modmult_1/xreg_reg[428]  ( .D(\modmult_1/xin[427] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[428]), .Q(\modmult_1/xin[428] ) );
  DFF \modmult_1/xreg_reg[427]  ( .D(\modmult_1/xin[426] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[427]), .Q(\modmult_1/xin[427] ) );
  DFF \modmult_1/xreg_reg[426]  ( .D(\modmult_1/xin[425] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[426]), .Q(\modmult_1/xin[426] ) );
  DFF \modmult_1/xreg_reg[425]  ( .D(\modmult_1/xin[424] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[425]), .Q(\modmult_1/xin[425] ) );
  DFF \modmult_1/xreg_reg[424]  ( .D(\modmult_1/xin[423] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[424]), .Q(\modmult_1/xin[424] ) );
  DFF \modmult_1/xreg_reg[423]  ( .D(\modmult_1/xin[422] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[423]), .Q(\modmult_1/xin[423] ) );
  DFF \modmult_1/xreg_reg[422]  ( .D(\modmult_1/xin[421] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[422]), .Q(\modmult_1/xin[422] ) );
  DFF \modmult_1/xreg_reg[421]  ( .D(\modmult_1/xin[420] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[421]), .Q(\modmult_1/xin[421] ) );
  DFF \modmult_1/xreg_reg[420]  ( .D(\modmult_1/xin[419] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[420]), .Q(\modmult_1/xin[420] ) );
  DFF \modmult_1/xreg_reg[419]  ( .D(\modmult_1/xin[418] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[419]), .Q(\modmult_1/xin[419] ) );
  DFF \modmult_1/xreg_reg[418]  ( .D(\modmult_1/xin[417] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[418]), .Q(\modmult_1/xin[418] ) );
  DFF \modmult_1/xreg_reg[417]  ( .D(\modmult_1/xin[416] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[417]), .Q(\modmult_1/xin[417] ) );
  DFF \modmult_1/xreg_reg[416]  ( .D(\modmult_1/xin[415] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[416]), .Q(\modmult_1/xin[416] ) );
  DFF \modmult_1/xreg_reg[415]  ( .D(\modmult_1/xin[414] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[415]), .Q(\modmult_1/xin[415] ) );
  DFF \modmult_1/xreg_reg[414]  ( .D(\modmult_1/xin[413] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[414]), .Q(\modmult_1/xin[414] ) );
  DFF \modmult_1/xreg_reg[413]  ( .D(\modmult_1/xin[412] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[413]), .Q(\modmult_1/xin[413] ) );
  DFF \modmult_1/xreg_reg[412]  ( .D(\modmult_1/xin[411] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[412]), .Q(\modmult_1/xin[412] ) );
  DFF \modmult_1/xreg_reg[411]  ( .D(\modmult_1/xin[410] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[411]), .Q(\modmult_1/xin[411] ) );
  DFF \modmult_1/xreg_reg[410]  ( .D(\modmult_1/xin[409] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[410]), .Q(\modmult_1/xin[410] ) );
  DFF \modmult_1/xreg_reg[409]  ( .D(\modmult_1/xin[408] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[409]), .Q(\modmult_1/xin[409] ) );
  DFF \modmult_1/xreg_reg[408]  ( .D(\modmult_1/xin[407] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[408]), .Q(\modmult_1/xin[408] ) );
  DFF \modmult_1/xreg_reg[407]  ( .D(\modmult_1/xin[406] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[407]), .Q(\modmult_1/xin[407] ) );
  DFF \modmult_1/xreg_reg[406]  ( .D(\modmult_1/xin[405] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[406]), .Q(\modmult_1/xin[406] ) );
  DFF \modmult_1/xreg_reg[405]  ( .D(\modmult_1/xin[404] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[405]), .Q(\modmult_1/xin[405] ) );
  DFF \modmult_1/xreg_reg[404]  ( .D(\modmult_1/xin[403] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[404]), .Q(\modmult_1/xin[404] ) );
  DFF \modmult_1/xreg_reg[403]  ( .D(\modmult_1/xin[402] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[403]), .Q(\modmult_1/xin[403] ) );
  DFF \modmult_1/xreg_reg[402]  ( .D(\modmult_1/xin[401] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[402]), .Q(\modmult_1/xin[402] ) );
  DFF \modmult_1/xreg_reg[401]  ( .D(\modmult_1/xin[400] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[401]), .Q(\modmult_1/xin[401] ) );
  DFF \modmult_1/xreg_reg[400]  ( .D(\modmult_1/xin[399] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[400]), .Q(\modmult_1/xin[400] ) );
  DFF \modmult_1/xreg_reg[399]  ( .D(\modmult_1/xin[398] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[399]), .Q(\modmult_1/xin[399] ) );
  DFF \modmult_1/xreg_reg[398]  ( .D(\modmult_1/xin[397] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[398]), .Q(\modmult_1/xin[398] ) );
  DFF \modmult_1/xreg_reg[397]  ( .D(\modmult_1/xin[396] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[397]), .Q(\modmult_1/xin[397] ) );
  DFF \modmult_1/xreg_reg[396]  ( .D(\modmult_1/xin[395] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[396]), .Q(\modmult_1/xin[396] ) );
  DFF \modmult_1/xreg_reg[395]  ( .D(\modmult_1/xin[394] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[395]), .Q(\modmult_1/xin[395] ) );
  DFF \modmult_1/xreg_reg[394]  ( .D(\modmult_1/xin[393] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[394]), .Q(\modmult_1/xin[394] ) );
  DFF \modmult_1/xreg_reg[393]  ( .D(\modmult_1/xin[392] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[393]), .Q(\modmult_1/xin[393] ) );
  DFF \modmult_1/xreg_reg[392]  ( .D(\modmult_1/xin[391] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[392]), .Q(\modmult_1/xin[392] ) );
  DFF \modmult_1/xreg_reg[391]  ( .D(\modmult_1/xin[390] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[391]), .Q(\modmult_1/xin[391] ) );
  DFF \modmult_1/xreg_reg[390]  ( .D(\modmult_1/xin[389] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[390]), .Q(\modmult_1/xin[390] ) );
  DFF \modmult_1/xreg_reg[389]  ( .D(\modmult_1/xin[388] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[389]), .Q(\modmult_1/xin[389] ) );
  DFF \modmult_1/xreg_reg[388]  ( .D(\modmult_1/xin[387] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[388]), .Q(\modmult_1/xin[388] ) );
  DFF \modmult_1/xreg_reg[387]  ( .D(\modmult_1/xin[386] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[387]), .Q(\modmult_1/xin[387] ) );
  DFF \modmult_1/xreg_reg[386]  ( .D(\modmult_1/xin[385] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[386]), .Q(\modmult_1/xin[386] ) );
  DFF \modmult_1/xreg_reg[385]  ( .D(\modmult_1/xin[384] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[385]), .Q(\modmult_1/xin[385] ) );
  DFF \modmult_1/xreg_reg[384]  ( .D(\modmult_1/xin[383] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[384]), .Q(\modmult_1/xin[384] ) );
  DFF \modmult_1/xreg_reg[383]  ( .D(\modmult_1/xin[382] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[383]), .Q(\modmult_1/xin[383] ) );
  DFF \modmult_1/xreg_reg[382]  ( .D(\modmult_1/xin[381] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[382]), .Q(\modmult_1/xin[382] ) );
  DFF \modmult_1/xreg_reg[381]  ( .D(\modmult_1/xin[380] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[381]), .Q(\modmult_1/xin[381] ) );
  DFF \modmult_1/xreg_reg[380]  ( .D(\modmult_1/xin[379] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[380]), .Q(\modmult_1/xin[380] ) );
  DFF \modmult_1/xreg_reg[379]  ( .D(\modmult_1/xin[378] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[379]), .Q(\modmult_1/xin[379] ) );
  DFF \modmult_1/xreg_reg[378]  ( .D(\modmult_1/xin[377] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[378]), .Q(\modmult_1/xin[378] ) );
  DFF \modmult_1/xreg_reg[377]  ( .D(\modmult_1/xin[376] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[377]), .Q(\modmult_1/xin[377] ) );
  DFF \modmult_1/xreg_reg[376]  ( .D(\modmult_1/xin[375] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[376]), .Q(\modmult_1/xin[376] ) );
  DFF \modmult_1/xreg_reg[375]  ( .D(\modmult_1/xin[374] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[375]), .Q(\modmult_1/xin[375] ) );
  DFF \modmult_1/xreg_reg[374]  ( .D(\modmult_1/xin[373] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[374]), .Q(\modmult_1/xin[374] ) );
  DFF \modmult_1/xreg_reg[373]  ( .D(\modmult_1/xin[372] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[373]), .Q(\modmult_1/xin[373] ) );
  DFF \modmult_1/xreg_reg[372]  ( .D(\modmult_1/xin[371] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[372]), .Q(\modmult_1/xin[372] ) );
  DFF \modmult_1/xreg_reg[371]  ( .D(\modmult_1/xin[370] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[371]), .Q(\modmult_1/xin[371] ) );
  DFF \modmult_1/xreg_reg[370]  ( .D(\modmult_1/xin[369] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[370]), .Q(\modmult_1/xin[370] ) );
  DFF \modmult_1/xreg_reg[369]  ( .D(\modmult_1/xin[368] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[369]), .Q(\modmult_1/xin[369] ) );
  DFF \modmult_1/xreg_reg[368]  ( .D(\modmult_1/xin[367] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[368]), .Q(\modmult_1/xin[368] ) );
  DFF \modmult_1/xreg_reg[367]  ( .D(\modmult_1/xin[366] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[367]), .Q(\modmult_1/xin[367] ) );
  DFF \modmult_1/xreg_reg[366]  ( .D(\modmult_1/xin[365] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[366]), .Q(\modmult_1/xin[366] ) );
  DFF \modmult_1/xreg_reg[365]  ( .D(\modmult_1/xin[364] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[365]), .Q(\modmult_1/xin[365] ) );
  DFF \modmult_1/xreg_reg[364]  ( .D(\modmult_1/xin[363] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[364]), .Q(\modmult_1/xin[364] ) );
  DFF \modmult_1/xreg_reg[363]  ( .D(\modmult_1/xin[362] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[363]), .Q(\modmult_1/xin[363] ) );
  DFF \modmult_1/xreg_reg[362]  ( .D(\modmult_1/xin[361] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[362]), .Q(\modmult_1/xin[362] ) );
  DFF \modmult_1/xreg_reg[361]  ( .D(\modmult_1/xin[360] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[361]), .Q(\modmult_1/xin[361] ) );
  DFF \modmult_1/xreg_reg[360]  ( .D(\modmult_1/xin[359] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[360]), .Q(\modmult_1/xin[360] ) );
  DFF \modmult_1/xreg_reg[359]  ( .D(\modmult_1/xin[358] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[359]), .Q(\modmult_1/xin[359] ) );
  DFF \modmult_1/xreg_reg[358]  ( .D(\modmult_1/xin[357] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[358]), .Q(\modmult_1/xin[358] ) );
  DFF \modmult_1/xreg_reg[357]  ( .D(\modmult_1/xin[356] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[357]), .Q(\modmult_1/xin[357] ) );
  DFF \modmult_1/xreg_reg[356]  ( .D(\modmult_1/xin[355] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[356]), .Q(\modmult_1/xin[356] ) );
  DFF \modmult_1/xreg_reg[355]  ( .D(\modmult_1/xin[354] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[355]), .Q(\modmult_1/xin[355] ) );
  DFF \modmult_1/xreg_reg[354]  ( .D(\modmult_1/xin[353] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[354]), .Q(\modmult_1/xin[354] ) );
  DFF \modmult_1/xreg_reg[353]  ( .D(\modmult_1/xin[352] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[353]), .Q(\modmult_1/xin[353] ) );
  DFF \modmult_1/xreg_reg[352]  ( .D(\modmult_1/xin[351] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[352]), .Q(\modmult_1/xin[352] ) );
  DFF \modmult_1/xreg_reg[351]  ( .D(\modmult_1/xin[350] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[351]), .Q(\modmult_1/xin[351] ) );
  DFF \modmult_1/xreg_reg[350]  ( .D(\modmult_1/xin[349] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[350]), .Q(\modmult_1/xin[350] ) );
  DFF \modmult_1/xreg_reg[349]  ( .D(\modmult_1/xin[348] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[349]), .Q(\modmult_1/xin[349] ) );
  DFF \modmult_1/xreg_reg[348]  ( .D(\modmult_1/xin[347] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[348]), .Q(\modmult_1/xin[348] ) );
  DFF \modmult_1/xreg_reg[347]  ( .D(\modmult_1/xin[346] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[347]), .Q(\modmult_1/xin[347] ) );
  DFF \modmult_1/xreg_reg[346]  ( .D(\modmult_1/xin[345] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[346]), .Q(\modmult_1/xin[346] ) );
  DFF \modmult_1/xreg_reg[345]  ( .D(\modmult_1/xin[344] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[345]), .Q(\modmult_1/xin[345] ) );
  DFF \modmult_1/xreg_reg[344]  ( .D(\modmult_1/xin[343] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[344]), .Q(\modmult_1/xin[344] ) );
  DFF \modmult_1/xreg_reg[343]  ( .D(\modmult_1/xin[342] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[343]), .Q(\modmult_1/xin[343] ) );
  DFF \modmult_1/xreg_reg[342]  ( .D(\modmult_1/xin[341] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[342]), .Q(\modmult_1/xin[342] ) );
  DFF \modmult_1/xreg_reg[341]  ( .D(\modmult_1/xin[340] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[341]), .Q(\modmult_1/xin[341] ) );
  DFF \modmult_1/xreg_reg[340]  ( .D(\modmult_1/xin[339] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[340]), .Q(\modmult_1/xin[340] ) );
  DFF \modmult_1/xreg_reg[339]  ( .D(\modmult_1/xin[338] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[339]), .Q(\modmult_1/xin[339] ) );
  DFF \modmult_1/xreg_reg[338]  ( .D(\modmult_1/xin[337] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[338]), .Q(\modmult_1/xin[338] ) );
  DFF \modmult_1/xreg_reg[337]  ( .D(\modmult_1/xin[336] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[337]), .Q(\modmult_1/xin[337] ) );
  DFF \modmult_1/xreg_reg[336]  ( .D(\modmult_1/xin[335] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[336]), .Q(\modmult_1/xin[336] ) );
  DFF \modmult_1/xreg_reg[335]  ( .D(\modmult_1/xin[334] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[335]), .Q(\modmult_1/xin[335] ) );
  DFF \modmult_1/xreg_reg[334]  ( .D(\modmult_1/xin[333] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[334]), .Q(\modmult_1/xin[334] ) );
  DFF \modmult_1/xreg_reg[333]  ( .D(\modmult_1/xin[332] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[333]), .Q(\modmult_1/xin[333] ) );
  DFF \modmult_1/xreg_reg[332]  ( .D(\modmult_1/xin[331] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[332]), .Q(\modmult_1/xin[332] ) );
  DFF \modmult_1/xreg_reg[331]  ( .D(\modmult_1/xin[330] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[331]), .Q(\modmult_1/xin[331] ) );
  DFF \modmult_1/xreg_reg[330]  ( .D(\modmult_1/xin[329] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[330]), .Q(\modmult_1/xin[330] ) );
  DFF \modmult_1/xreg_reg[329]  ( .D(\modmult_1/xin[328] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[329]), .Q(\modmult_1/xin[329] ) );
  DFF \modmult_1/xreg_reg[328]  ( .D(\modmult_1/xin[327] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[328]), .Q(\modmult_1/xin[328] ) );
  DFF \modmult_1/xreg_reg[327]  ( .D(\modmult_1/xin[326] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[327]), .Q(\modmult_1/xin[327] ) );
  DFF \modmult_1/xreg_reg[326]  ( .D(\modmult_1/xin[325] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[326]), .Q(\modmult_1/xin[326] ) );
  DFF \modmult_1/xreg_reg[325]  ( .D(\modmult_1/xin[324] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[325]), .Q(\modmult_1/xin[325] ) );
  DFF \modmult_1/xreg_reg[324]  ( .D(\modmult_1/xin[323] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[324]), .Q(\modmult_1/xin[324] ) );
  DFF \modmult_1/xreg_reg[323]  ( .D(\modmult_1/xin[322] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[323]), .Q(\modmult_1/xin[323] ) );
  DFF \modmult_1/xreg_reg[322]  ( .D(\modmult_1/xin[321] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[322]), .Q(\modmult_1/xin[322] ) );
  DFF \modmult_1/xreg_reg[321]  ( .D(\modmult_1/xin[320] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[321]), .Q(\modmult_1/xin[321] ) );
  DFF \modmult_1/xreg_reg[320]  ( .D(\modmult_1/xin[319] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[320]), .Q(\modmult_1/xin[320] ) );
  DFF \modmult_1/xreg_reg[319]  ( .D(\modmult_1/xin[318] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[319]), .Q(\modmult_1/xin[319] ) );
  DFF \modmult_1/xreg_reg[318]  ( .D(\modmult_1/xin[317] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[318]), .Q(\modmult_1/xin[318] ) );
  DFF \modmult_1/xreg_reg[317]  ( .D(\modmult_1/xin[316] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[317]), .Q(\modmult_1/xin[317] ) );
  DFF \modmult_1/xreg_reg[316]  ( .D(\modmult_1/xin[315] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[316]), .Q(\modmult_1/xin[316] ) );
  DFF \modmult_1/xreg_reg[315]  ( .D(\modmult_1/xin[314] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[315]), .Q(\modmult_1/xin[315] ) );
  DFF \modmult_1/xreg_reg[314]  ( .D(\modmult_1/xin[313] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[314]), .Q(\modmult_1/xin[314] ) );
  DFF \modmult_1/xreg_reg[313]  ( .D(\modmult_1/xin[312] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[313]), .Q(\modmult_1/xin[313] ) );
  DFF \modmult_1/xreg_reg[312]  ( .D(\modmult_1/xin[311] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[312]), .Q(\modmult_1/xin[312] ) );
  DFF \modmult_1/xreg_reg[311]  ( .D(\modmult_1/xin[310] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[311]), .Q(\modmult_1/xin[311] ) );
  DFF \modmult_1/xreg_reg[310]  ( .D(\modmult_1/xin[309] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[310]), .Q(\modmult_1/xin[310] ) );
  DFF \modmult_1/xreg_reg[309]  ( .D(\modmult_1/xin[308] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[309]), .Q(\modmult_1/xin[309] ) );
  DFF \modmult_1/xreg_reg[308]  ( .D(\modmult_1/xin[307] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[308]), .Q(\modmult_1/xin[308] ) );
  DFF \modmult_1/xreg_reg[307]  ( .D(\modmult_1/xin[306] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[307]), .Q(\modmult_1/xin[307] ) );
  DFF \modmult_1/xreg_reg[306]  ( .D(\modmult_1/xin[305] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[306]), .Q(\modmult_1/xin[306] ) );
  DFF \modmult_1/xreg_reg[305]  ( .D(\modmult_1/xin[304] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[305]), .Q(\modmult_1/xin[305] ) );
  DFF \modmult_1/xreg_reg[304]  ( .D(\modmult_1/xin[303] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[304]), .Q(\modmult_1/xin[304] ) );
  DFF \modmult_1/xreg_reg[303]  ( .D(\modmult_1/xin[302] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[303]), .Q(\modmult_1/xin[303] ) );
  DFF \modmult_1/xreg_reg[302]  ( .D(\modmult_1/xin[301] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[302]), .Q(\modmult_1/xin[302] ) );
  DFF \modmult_1/xreg_reg[301]  ( .D(\modmult_1/xin[300] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[301]), .Q(\modmult_1/xin[301] ) );
  DFF \modmult_1/xreg_reg[300]  ( .D(\modmult_1/xin[299] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[300]), .Q(\modmult_1/xin[300] ) );
  DFF \modmult_1/xreg_reg[299]  ( .D(\modmult_1/xin[298] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[299]), .Q(\modmult_1/xin[299] ) );
  DFF \modmult_1/xreg_reg[298]  ( .D(\modmult_1/xin[297] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[298]), .Q(\modmult_1/xin[298] ) );
  DFF \modmult_1/xreg_reg[297]  ( .D(\modmult_1/xin[296] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[297]), .Q(\modmult_1/xin[297] ) );
  DFF \modmult_1/xreg_reg[296]  ( .D(\modmult_1/xin[295] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[296]), .Q(\modmult_1/xin[296] ) );
  DFF \modmult_1/xreg_reg[295]  ( .D(\modmult_1/xin[294] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[295]), .Q(\modmult_1/xin[295] ) );
  DFF \modmult_1/xreg_reg[294]  ( .D(\modmult_1/xin[293] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[294]), .Q(\modmult_1/xin[294] ) );
  DFF \modmult_1/xreg_reg[293]  ( .D(\modmult_1/xin[292] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[293]), .Q(\modmult_1/xin[293] ) );
  DFF \modmult_1/xreg_reg[292]  ( .D(\modmult_1/xin[291] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[292]), .Q(\modmult_1/xin[292] ) );
  DFF \modmult_1/xreg_reg[291]  ( .D(\modmult_1/xin[290] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[291]), .Q(\modmult_1/xin[291] ) );
  DFF \modmult_1/xreg_reg[290]  ( .D(\modmult_1/xin[289] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[290]), .Q(\modmult_1/xin[290] ) );
  DFF \modmult_1/xreg_reg[289]  ( .D(\modmult_1/xin[288] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[289]), .Q(\modmult_1/xin[289] ) );
  DFF \modmult_1/xreg_reg[288]  ( .D(\modmult_1/xin[287] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[288]), .Q(\modmult_1/xin[288] ) );
  DFF \modmult_1/xreg_reg[287]  ( .D(\modmult_1/xin[286] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[287]), .Q(\modmult_1/xin[287] ) );
  DFF \modmult_1/xreg_reg[286]  ( .D(\modmult_1/xin[285] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[286]), .Q(\modmult_1/xin[286] ) );
  DFF \modmult_1/xreg_reg[285]  ( .D(\modmult_1/xin[284] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[285]), .Q(\modmult_1/xin[285] ) );
  DFF \modmult_1/xreg_reg[284]  ( .D(\modmult_1/xin[283] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[284]), .Q(\modmult_1/xin[284] ) );
  DFF \modmult_1/xreg_reg[283]  ( .D(\modmult_1/xin[282] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[283]), .Q(\modmult_1/xin[283] ) );
  DFF \modmult_1/xreg_reg[282]  ( .D(\modmult_1/xin[281] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[282]), .Q(\modmult_1/xin[282] ) );
  DFF \modmult_1/xreg_reg[281]  ( .D(\modmult_1/xin[280] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[281]), .Q(\modmult_1/xin[281] ) );
  DFF \modmult_1/xreg_reg[280]  ( .D(\modmult_1/xin[279] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[280]), .Q(\modmult_1/xin[280] ) );
  DFF \modmult_1/xreg_reg[279]  ( .D(\modmult_1/xin[278] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[279]), .Q(\modmult_1/xin[279] ) );
  DFF \modmult_1/xreg_reg[278]  ( .D(\modmult_1/xin[277] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[278]), .Q(\modmult_1/xin[278] ) );
  DFF \modmult_1/xreg_reg[277]  ( .D(\modmult_1/xin[276] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[277]), .Q(\modmult_1/xin[277] ) );
  DFF \modmult_1/xreg_reg[276]  ( .D(\modmult_1/xin[275] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[276]), .Q(\modmult_1/xin[276] ) );
  DFF \modmult_1/xreg_reg[275]  ( .D(\modmult_1/xin[274] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[275]), .Q(\modmult_1/xin[275] ) );
  DFF \modmult_1/xreg_reg[274]  ( .D(\modmult_1/xin[273] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[274]), .Q(\modmult_1/xin[274] ) );
  DFF \modmult_1/xreg_reg[273]  ( .D(\modmult_1/xin[272] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[273]), .Q(\modmult_1/xin[273] ) );
  DFF \modmult_1/xreg_reg[272]  ( .D(\modmult_1/xin[271] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[272]), .Q(\modmult_1/xin[272] ) );
  DFF \modmult_1/xreg_reg[271]  ( .D(\modmult_1/xin[270] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[271]), .Q(\modmult_1/xin[271] ) );
  DFF \modmult_1/xreg_reg[270]  ( .D(\modmult_1/xin[269] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[270]), .Q(\modmult_1/xin[270] ) );
  DFF \modmult_1/xreg_reg[269]  ( .D(\modmult_1/xin[268] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[269]), .Q(\modmult_1/xin[269] ) );
  DFF \modmult_1/xreg_reg[268]  ( .D(\modmult_1/xin[267] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[268]), .Q(\modmult_1/xin[268] ) );
  DFF \modmult_1/xreg_reg[267]  ( .D(\modmult_1/xin[266] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[267]), .Q(\modmult_1/xin[267] ) );
  DFF \modmult_1/xreg_reg[266]  ( .D(\modmult_1/xin[265] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[266]), .Q(\modmult_1/xin[266] ) );
  DFF \modmult_1/xreg_reg[265]  ( .D(\modmult_1/xin[264] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[265]), .Q(\modmult_1/xin[265] ) );
  DFF \modmult_1/xreg_reg[264]  ( .D(\modmult_1/xin[263] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[264]), .Q(\modmult_1/xin[264] ) );
  DFF \modmult_1/xreg_reg[263]  ( .D(\modmult_1/xin[262] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[263]), .Q(\modmult_1/xin[263] ) );
  DFF \modmult_1/xreg_reg[262]  ( .D(\modmult_1/xin[261] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[262]), .Q(\modmult_1/xin[262] ) );
  DFF \modmult_1/xreg_reg[261]  ( .D(\modmult_1/xin[260] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[261]), .Q(\modmult_1/xin[261] ) );
  DFF \modmult_1/xreg_reg[260]  ( .D(\modmult_1/xin[259] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[260]), .Q(\modmult_1/xin[260] ) );
  DFF \modmult_1/xreg_reg[259]  ( .D(\modmult_1/xin[258] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[259]), .Q(\modmult_1/xin[259] ) );
  DFF \modmult_1/xreg_reg[258]  ( .D(\modmult_1/xin[257] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[258]), .Q(\modmult_1/xin[258] ) );
  DFF \modmult_1/xreg_reg[257]  ( .D(\modmult_1/xin[256] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[257]), .Q(\modmult_1/xin[257] ) );
  DFF \modmult_1/xreg_reg[256]  ( .D(\modmult_1/xin[255] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[256]), .Q(\modmult_1/xin[256] ) );
  DFF \modmult_1/xreg_reg[255]  ( .D(\modmult_1/xin[254] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[255]), .Q(\modmult_1/xin[255] ) );
  DFF \modmult_1/xreg_reg[254]  ( .D(\modmult_1/xin[253] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[254]), .Q(\modmult_1/xin[254] ) );
  DFF \modmult_1/xreg_reg[253]  ( .D(\modmult_1/xin[252] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[253]), .Q(\modmult_1/xin[253] ) );
  DFF \modmult_1/xreg_reg[252]  ( .D(\modmult_1/xin[251] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[252]), .Q(\modmult_1/xin[252] ) );
  DFF \modmult_1/xreg_reg[251]  ( .D(\modmult_1/xin[250] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[251]), .Q(\modmult_1/xin[251] ) );
  DFF \modmult_1/xreg_reg[250]  ( .D(\modmult_1/xin[249] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[250]), .Q(\modmult_1/xin[250] ) );
  DFF \modmult_1/xreg_reg[249]  ( .D(\modmult_1/xin[248] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[249]), .Q(\modmult_1/xin[249] ) );
  DFF \modmult_1/xreg_reg[248]  ( .D(\modmult_1/xin[247] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[248]), .Q(\modmult_1/xin[248] ) );
  DFF \modmult_1/xreg_reg[247]  ( .D(\modmult_1/xin[246] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[247]), .Q(\modmult_1/xin[247] ) );
  DFF \modmult_1/xreg_reg[246]  ( .D(\modmult_1/xin[245] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[246]), .Q(\modmult_1/xin[246] ) );
  DFF \modmult_1/xreg_reg[245]  ( .D(\modmult_1/xin[244] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[245]), .Q(\modmult_1/xin[245] ) );
  DFF \modmult_1/xreg_reg[244]  ( .D(\modmult_1/xin[243] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[244]), .Q(\modmult_1/xin[244] ) );
  DFF \modmult_1/xreg_reg[243]  ( .D(\modmult_1/xin[242] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[243]), .Q(\modmult_1/xin[243] ) );
  DFF \modmult_1/xreg_reg[242]  ( .D(\modmult_1/xin[241] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[242]), .Q(\modmult_1/xin[242] ) );
  DFF \modmult_1/xreg_reg[241]  ( .D(\modmult_1/xin[240] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[241]), .Q(\modmult_1/xin[241] ) );
  DFF \modmult_1/xreg_reg[240]  ( .D(\modmult_1/xin[239] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[240]), .Q(\modmult_1/xin[240] ) );
  DFF \modmult_1/xreg_reg[239]  ( .D(\modmult_1/xin[238] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[239]), .Q(\modmult_1/xin[239] ) );
  DFF \modmult_1/xreg_reg[238]  ( .D(\modmult_1/xin[237] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[238]), .Q(\modmult_1/xin[238] ) );
  DFF \modmult_1/xreg_reg[237]  ( .D(\modmult_1/xin[236] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[237]), .Q(\modmult_1/xin[237] ) );
  DFF \modmult_1/xreg_reg[236]  ( .D(\modmult_1/xin[235] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[236]), .Q(\modmult_1/xin[236] ) );
  DFF \modmult_1/xreg_reg[235]  ( .D(\modmult_1/xin[234] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[235]), .Q(\modmult_1/xin[235] ) );
  DFF \modmult_1/xreg_reg[234]  ( .D(\modmult_1/xin[233] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[234]), .Q(\modmult_1/xin[234] ) );
  DFF \modmult_1/xreg_reg[233]  ( .D(\modmult_1/xin[232] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[233]), .Q(\modmult_1/xin[233] ) );
  DFF \modmult_1/xreg_reg[232]  ( .D(\modmult_1/xin[231] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[232]), .Q(\modmult_1/xin[232] ) );
  DFF \modmult_1/xreg_reg[231]  ( .D(\modmult_1/xin[230] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[231]), .Q(\modmult_1/xin[231] ) );
  DFF \modmult_1/xreg_reg[230]  ( .D(\modmult_1/xin[229] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[230]), .Q(\modmult_1/xin[230] ) );
  DFF \modmult_1/xreg_reg[229]  ( .D(\modmult_1/xin[228] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[229]), .Q(\modmult_1/xin[229] ) );
  DFF \modmult_1/xreg_reg[228]  ( .D(\modmult_1/xin[227] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[228]), .Q(\modmult_1/xin[228] ) );
  DFF \modmult_1/xreg_reg[227]  ( .D(\modmult_1/xin[226] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[227]), .Q(\modmult_1/xin[227] ) );
  DFF \modmult_1/xreg_reg[226]  ( .D(\modmult_1/xin[225] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[226]), .Q(\modmult_1/xin[226] ) );
  DFF \modmult_1/xreg_reg[225]  ( .D(\modmult_1/xin[224] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[225]), .Q(\modmult_1/xin[225] ) );
  DFF \modmult_1/xreg_reg[224]  ( .D(\modmult_1/xin[223] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[224]), .Q(\modmult_1/xin[224] ) );
  DFF \modmult_1/xreg_reg[223]  ( .D(\modmult_1/xin[222] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[223]), .Q(\modmult_1/xin[223] ) );
  DFF \modmult_1/xreg_reg[222]  ( .D(\modmult_1/xin[221] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[222]), .Q(\modmult_1/xin[222] ) );
  DFF \modmult_1/xreg_reg[221]  ( .D(\modmult_1/xin[220] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[221]), .Q(\modmult_1/xin[221] ) );
  DFF \modmult_1/xreg_reg[220]  ( .D(\modmult_1/xin[219] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[220]), .Q(\modmult_1/xin[220] ) );
  DFF \modmult_1/xreg_reg[219]  ( .D(\modmult_1/xin[218] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[219]), .Q(\modmult_1/xin[219] ) );
  DFF \modmult_1/xreg_reg[218]  ( .D(\modmult_1/xin[217] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[218]), .Q(\modmult_1/xin[218] ) );
  DFF \modmult_1/xreg_reg[217]  ( .D(\modmult_1/xin[216] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[217]), .Q(\modmult_1/xin[217] ) );
  DFF \modmult_1/xreg_reg[216]  ( .D(\modmult_1/xin[215] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[216]), .Q(\modmult_1/xin[216] ) );
  DFF \modmult_1/xreg_reg[215]  ( .D(\modmult_1/xin[214] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[215]), .Q(\modmult_1/xin[215] ) );
  DFF \modmult_1/xreg_reg[214]  ( .D(\modmult_1/xin[213] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[214]), .Q(\modmult_1/xin[214] ) );
  DFF \modmult_1/xreg_reg[213]  ( .D(\modmult_1/xin[212] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[213]), .Q(\modmult_1/xin[213] ) );
  DFF \modmult_1/xreg_reg[212]  ( .D(\modmult_1/xin[211] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[212]), .Q(\modmult_1/xin[212] ) );
  DFF \modmult_1/xreg_reg[211]  ( .D(\modmult_1/xin[210] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[211]), .Q(\modmult_1/xin[211] ) );
  DFF \modmult_1/xreg_reg[210]  ( .D(\modmult_1/xin[209] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[210]), .Q(\modmult_1/xin[210] ) );
  DFF \modmult_1/xreg_reg[209]  ( .D(\modmult_1/xin[208] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[209]), .Q(\modmult_1/xin[209] ) );
  DFF \modmult_1/xreg_reg[208]  ( .D(\modmult_1/xin[207] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[208]), .Q(\modmult_1/xin[208] ) );
  DFF \modmult_1/xreg_reg[207]  ( .D(\modmult_1/xin[206] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[207]), .Q(\modmult_1/xin[207] ) );
  DFF \modmult_1/xreg_reg[206]  ( .D(\modmult_1/xin[205] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[206]), .Q(\modmult_1/xin[206] ) );
  DFF \modmult_1/xreg_reg[205]  ( .D(\modmult_1/xin[204] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[205]), .Q(\modmult_1/xin[205] ) );
  DFF \modmult_1/xreg_reg[204]  ( .D(\modmult_1/xin[203] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[204]), .Q(\modmult_1/xin[204] ) );
  DFF \modmult_1/xreg_reg[203]  ( .D(\modmult_1/xin[202] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[203]), .Q(\modmult_1/xin[203] ) );
  DFF \modmult_1/xreg_reg[202]  ( .D(\modmult_1/xin[201] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[202]), .Q(\modmult_1/xin[202] ) );
  DFF \modmult_1/xreg_reg[201]  ( .D(\modmult_1/xin[200] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[201]), .Q(\modmult_1/xin[201] ) );
  DFF \modmult_1/xreg_reg[200]  ( .D(\modmult_1/xin[199] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[200]), .Q(\modmult_1/xin[200] ) );
  DFF \modmult_1/xreg_reg[199]  ( .D(\modmult_1/xin[198] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[199]), .Q(\modmult_1/xin[199] ) );
  DFF \modmult_1/xreg_reg[198]  ( .D(\modmult_1/xin[197] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[198]), .Q(\modmult_1/xin[198] ) );
  DFF \modmult_1/xreg_reg[197]  ( .D(\modmult_1/xin[196] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[197]), .Q(\modmult_1/xin[197] ) );
  DFF \modmult_1/xreg_reg[196]  ( .D(\modmult_1/xin[195] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[196]), .Q(\modmult_1/xin[196] ) );
  DFF \modmult_1/xreg_reg[195]  ( .D(\modmult_1/xin[194] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[195]), .Q(\modmult_1/xin[195] ) );
  DFF \modmult_1/xreg_reg[194]  ( .D(\modmult_1/xin[193] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[194]), .Q(\modmult_1/xin[194] ) );
  DFF \modmult_1/xreg_reg[193]  ( .D(\modmult_1/xin[192] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[193]), .Q(\modmult_1/xin[193] ) );
  DFF \modmult_1/xreg_reg[192]  ( .D(\modmult_1/xin[191] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[192]), .Q(\modmult_1/xin[192] ) );
  DFF \modmult_1/xreg_reg[191]  ( .D(\modmult_1/xin[190] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[191]), .Q(\modmult_1/xin[191] ) );
  DFF \modmult_1/xreg_reg[190]  ( .D(\modmult_1/xin[189] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[190]), .Q(\modmult_1/xin[190] ) );
  DFF \modmult_1/xreg_reg[189]  ( .D(\modmult_1/xin[188] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[189]), .Q(\modmult_1/xin[189] ) );
  DFF \modmult_1/xreg_reg[188]  ( .D(\modmult_1/xin[187] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[188]), .Q(\modmult_1/xin[188] ) );
  DFF \modmult_1/xreg_reg[187]  ( .D(\modmult_1/xin[186] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[187]), .Q(\modmult_1/xin[187] ) );
  DFF \modmult_1/xreg_reg[186]  ( .D(\modmult_1/xin[185] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[186]), .Q(\modmult_1/xin[186] ) );
  DFF \modmult_1/xreg_reg[185]  ( .D(\modmult_1/xin[184] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[185]), .Q(\modmult_1/xin[185] ) );
  DFF \modmult_1/xreg_reg[184]  ( .D(\modmult_1/xin[183] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[184]), .Q(\modmult_1/xin[184] ) );
  DFF \modmult_1/xreg_reg[183]  ( .D(\modmult_1/xin[182] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[183]), .Q(\modmult_1/xin[183] ) );
  DFF \modmult_1/xreg_reg[182]  ( .D(\modmult_1/xin[181] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[182]), .Q(\modmult_1/xin[182] ) );
  DFF \modmult_1/xreg_reg[181]  ( .D(\modmult_1/xin[180] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[181]), .Q(\modmult_1/xin[181] ) );
  DFF \modmult_1/xreg_reg[180]  ( .D(\modmult_1/xin[179] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[180]), .Q(\modmult_1/xin[180] ) );
  DFF \modmult_1/xreg_reg[179]  ( .D(\modmult_1/xin[178] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[179]), .Q(\modmult_1/xin[179] ) );
  DFF \modmult_1/xreg_reg[178]  ( .D(\modmult_1/xin[177] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[178]), .Q(\modmult_1/xin[178] ) );
  DFF \modmult_1/xreg_reg[177]  ( .D(\modmult_1/xin[176] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[177]), .Q(\modmult_1/xin[177] ) );
  DFF \modmult_1/xreg_reg[176]  ( .D(\modmult_1/xin[175] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[176]), .Q(\modmult_1/xin[176] ) );
  DFF \modmult_1/xreg_reg[175]  ( .D(\modmult_1/xin[174] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[175]), .Q(\modmult_1/xin[175] ) );
  DFF \modmult_1/xreg_reg[174]  ( .D(\modmult_1/xin[173] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[174]), .Q(\modmult_1/xin[174] ) );
  DFF \modmult_1/xreg_reg[173]  ( .D(\modmult_1/xin[172] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[173]), .Q(\modmult_1/xin[173] ) );
  DFF \modmult_1/xreg_reg[172]  ( .D(\modmult_1/xin[171] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[172]), .Q(\modmult_1/xin[172] ) );
  DFF \modmult_1/xreg_reg[171]  ( .D(\modmult_1/xin[170] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[171]), .Q(\modmult_1/xin[171] ) );
  DFF \modmult_1/xreg_reg[170]  ( .D(\modmult_1/xin[169] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[170]), .Q(\modmult_1/xin[170] ) );
  DFF \modmult_1/xreg_reg[169]  ( .D(\modmult_1/xin[168] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[169]), .Q(\modmult_1/xin[169] ) );
  DFF \modmult_1/xreg_reg[168]  ( .D(\modmult_1/xin[167] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[168]), .Q(\modmult_1/xin[168] ) );
  DFF \modmult_1/xreg_reg[167]  ( .D(\modmult_1/xin[166] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[167]), .Q(\modmult_1/xin[167] ) );
  DFF \modmult_1/xreg_reg[166]  ( .D(\modmult_1/xin[165] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[166]), .Q(\modmult_1/xin[166] ) );
  DFF \modmult_1/xreg_reg[165]  ( .D(\modmult_1/xin[164] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[165]), .Q(\modmult_1/xin[165] ) );
  DFF \modmult_1/xreg_reg[164]  ( .D(\modmult_1/xin[163] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[164]), .Q(\modmult_1/xin[164] ) );
  DFF \modmult_1/xreg_reg[163]  ( .D(\modmult_1/xin[162] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[163]), .Q(\modmult_1/xin[163] ) );
  DFF \modmult_1/xreg_reg[162]  ( .D(\modmult_1/xin[161] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[162]), .Q(\modmult_1/xin[162] ) );
  DFF \modmult_1/xreg_reg[161]  ( .D(\modmult_1/xin[160] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[161]), .Q(\modmult_1/xin[161] ) );
  DFF \modmult_1/xreg_reg[160]  ( .D(\modmult_1/xin[159] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[160]), .Q(\modmult_1/xin[160] ) );
  DFF \modmult_1/xreg_reg[159]  ( .D(\modmult_1/xin[158] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[159]), .Q(\modmult_1/xin[159] ) );
  DFF \modmult_1/xreg_reg[158]  ( .D(\modmult_1/xin[157] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[158]), .Q(\modmult_1/xin[158] ) );
  DFF \modmult_1/xreg_reg[157]  ( .D(\modmult_1/xin[156] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[157]), .Q(\modmult_1/xin[157] ) );
  DFF \modmult_1/xreg_reg[156]  ( .D(\modmult_1/xin[155] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[156]), .Q(\modmult_1/xin[156] ) );
  DFF \modmult_1/xreg_reg[155]  ( .D(\modmult_1/xin[154] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[155]), .Q(\modmult_1/xin[155] ) );
  DFF \modmult_1/xreg_reg[154]  ( .D(\modmult_1/xin[153] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[154]), .Q(\modmult_1/xin[154] ) );
  DFF \modmult_1/xreg_reg[153]  ( .D(\modmult_1/xin[152] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[153]), .Q(\modmult_1/xin[153] ) );
  DFF \modmult_1/xreg_reg[152]  ( .D(\modmult_1/xin[151] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[152]), .Q(\modmult_1/xin[152] ) );
  DFF \modmult_1/xreg_reg[151]  ( .D(\modmult_1/xin[150] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[151]), .Q(\modmult_1/xin[151] ) );
  DFF \modmult_1/xreg_reg[150]  ( .D(\modmult_1/xin[149] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[150]), .Q(\modmult_1/xin[150] ) );
  DFF \modmult_1/xreg_reg[149]  ( .D(\modmult_1/xin[148] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[149]), .Q(\modmult_1/xin[149] ) );
  DFF \modmult_1/xreg_reg[148]  ( .D(\modmult_1/xin[147] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[148]), .Q(\modmult_1/xin[148] ) );
  DFF \modmult_1/xreg_reg[147]  ( .D(\modmult_1/xin[146] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[147]), .Q(\modmult_1/xin[147] ) );
  DFF \modmult_1/xreg_reg[146]  ( .D(\modmult_1/xin[145] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[146]), .Q(\modmult_1/xin[146] ) );
  DFF \modmult_1/xreg_reg[145]  ( .D(\modmult_1/xin[144] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[145]), .Q(\modmult_1/xin[145] ) );
  DFF \modmult_1/xreg_reg[144]  ( .D(\modmult_1/xin[143] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[144]), .Q(\modmult_1/xin[144] ) );
  DFF \modmult_1/xreg_reg[143]  ( .D(\modmult_1/xin[142] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[143]), .Q(\modmult_1/xin[143] ) );
  DFF \modmult_1/xreg_reg[142]  ( .D(\modmult_1/xin[141] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[142]), .Q(\modmult_1/xin[142] ) );
  DFF \modmult_1/xreg_reg[141]  ( .D(\modmult_1/xin[140] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[141]), .Q(\modmult_1/xin[141] ) );
  DFF \modmult_1/xreg_reg[140]  ( .D(\modmult_1/xin[139] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[140]), .Q(\modmult_1/xin[140] ) );
  DFF \modmult_1/xreg_reg[139]  ( .D(\modmult_1/xin[138] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[139]), .Q(\modmult_1/xin[139] ) );
  DFF \modmult_1/xreg_reg[138]  ( .D(\modmult_1/xin[137] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[138]), .Q(\modmult_1/xin[138] ) );
  DFF \modmult_1/xreg_reg[137]  ( .D(\modmult_1/xin[136] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[137]), .Q(\modmult_1/xin[137] ) );
  DFF \modmult_1/xreg_reg[136]  ( .D(\modmult_1/xin[135] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[136]), .Q(\modmult_1/xin[136] ) );
  DFF \modmult_1/xreg_reg[135]  ( .D(\modmult_1/xin[134] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[135]), .Q(\modmult_1/xin[135] ) );
  DFF \modmult_1/xreg_reg[134]  ( .D(\modmult_1/xin[133] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[134]), .Q(\modmult_1/xin[134] ) );
  DFF \modmult_1/xreg_reg[133]  ( .D(\modmult_1/xin[132] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[133]), .Q(\modmult_1/xin[133] ) );
  DFF \modmult_1/xreg_reg[132]  ( .D(\modmult_1/xin[131] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[132]), .Q(\modmult_1/xin[132] ) );
  DFF \modmult_1/xreg_reg[131]  ( .D(\modmult_1/xin[130] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[131]), .Q(\modmult_1/xin[131] ) );
  DFF \modmult_1/xreg_reg[130]  ( .D(\modmult_1/xin[129] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[130]), .Q(\modmult_1/xin[130] ) );
  DFF \modmult_1/xreg_reg[129]  ( .D(\modmult_1/xin[128] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[129]), .Q(\modmult_1/xin[129] ) );
  DFF \modmult_1/xreg_reg[128]  ( .D(\modmult_1/xin[127] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[128]), .Q(\modmult_1/xin[128] ) );
  DFF \modmult_1/xreg_reg[127]  ( .D(\modmult_1/xin[126] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[127]), .Q(\modmult_1/xin[127] ) );
  DFF \modmult_1/xreg_reg[126]  ( .D(\modmult_1/xin[125] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[126]), .Q(\modmult_1/xin[126] ) );
  DFF \modmult_1/xreg_reg[125]  ( .D(\modmult_1/xin[124] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[125]), .Q(\modmult_1/xin[125] ) );
  DFF \modmult_1/xreg_reg[124]  ( .D(\modmult_1/xin[123] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[124]), .Q(\modmult_1/xin[124] ) );
  DFF \modmult_1/xreg_reg[123]  ( .D(\modmult_1/xin[122] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[123]), .Q(\modmult_1/xin[123] ) );
  DFF \modmult_1/xreg_reg[122]  ( .D(\modmult_1/xin[121] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[122]), .Q(\modmult_1/xin[122] ) );
  DFF \modmult_1/xreg_reg[121]  ( .D(\modmult_1/xin[120] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[121]), .Q(\modmult_1/xin[121] ) );
  DFF \modmult_1/xreg_reg[120]  ( .D(\modmult_1/xin[119] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[120]), .Q(\modmult_1/xin[120] ) );
  DFF \modmult_1/xreg_reg[119]  ( .D(\modmult_1/xin[118] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[119]), .Q(\modmult_1/xin[119] ) );
  DFF \modmult_1/xreg_reg[118]  ( .D(\modmult_1/xin[117] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[118]), .Q(\modmult_1/xin[118] ) );
  DFF \modmult_1/xreg_reg[117]  ( .D(\modmult_1/xin[116] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[117]), .Q(\modmult_1/xin[117] ) );
  DFF \modmult_1/xreg_reg[116]  ( .D(\modmult_1/xin[115] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[116]), .Q(\modmult_1/xin[116] ) );
  DFF \modmult_1/xreg_reg[115]  ( .D(\modmult_1/xin[114] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[115]), .Q(\modmult_1/xin[115] ) );
  DFF \modmult_1/xreg_reg[114]  ( .D(\modmult_1/xin[113] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[114]), .Q(\modmult_1/xin[114] ) );
  DFF \modmult_1/xreg_reg[113]  ( .D(\modmult_1/xin[112] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[113]), .Q(\modmult_1/xin[113] ) );
  DFF \modmult_1/xreg_reg[112]  ( .D(\modmult_1/xin[111] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[112]), .Q(\modmult_1/xin[112] ) );
  DFF \modmult_1/xreg_reg[111]  ( .D(\modmult_1/xin[110] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[111]), .Q(\modmult_1/xin[111] ) );
  DFF \modmult_1/xreg_reg[110]  ( .D(\modmult_1/xin[109] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[110]), .Q(\modmult_1/xin[110] ) );
  DFF \modmult_1/xreg_reg[109]  ( .D(\modmult_1/xin[108] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[109]), .Q(\modmult_1/xin[109] ) );
  DFF \modmult_1/xreg_reg[108]  ( .D(\modmult_1/xin[107] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[108]), .Q(\modmult_1/xin[108] ) );
  DFF \modmult_1/xreg_reg[107]  ( .D(\modmult_1/xin[106] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[107]), .Q(\modmult_1/xin[107] ) );
  DFF \modmult_1/xreg_reg[106]  ( .D(\modmult_1/xin[105] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[106]), .Q(\modmult_1/xin[106] ) );
  DFF \modmult_1/xreg_reg[105]  ( .D(\modmult_1/xin[104] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[105]), .Q(\modmult_1/xin[105] ) );
  DFF \modmult_1/xreg_reg[104]  ( .D(\modmult_1/xin[103] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[104]), .Q(\modmult_1/xin[104] ) );
  DFF \modmult_1/xreg_reg[103]  ( .D(\modmult_1/xin[102] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[103]), .Q(\modmult_1/xin[103] ) );
  DFF \modmult_1/xreg_reg[102]  ( .D(\modmult_1/xin[101] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[102]), .Q(\modmult_1/xin[102] ) );
  DFF \modmult_1/xreg_reg[101]  ( .D(\modmult_1/xin[100] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[101]), .Q(\modmult_1/xin[101] ) );
  DFF \modmult_1/xreg_reg[100]  ( .D(\modmult_1/xin[99] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[100]), .Q(\modmult_1/xin[100] ) );
  DFF \modmult_1/xreg_reg[99]  ( .D(\modmult_1/xin[98] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[99]), .Q(\modmult_1/xin[99] ) );
  DFF \modmult_1/xreg_reg[98]  ( .D(\modmult_1/xin[97] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[98]), .Q(\modmult_1/xin[98] ) );
  DFF \modmult_1/xreg_reg[97]  ( .D(\modmult_1/xin[96] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[97]), .Q(\modmult_1/xin[97] ) );
  DFF \modmult_1/xreg_reg[96]  ( .D(\modmult_1/xin[95] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[96]), .Q(\modmult_1/xin[96] ) );
  DFF \modmult_1/xreg_reg[95]  ( .D(\modmult_1/xin[94] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[95]), .Q(\modmult_1/xin[95] ) );
  DFF \modmult_1/xreg_reg[94]  ( .D(\modmult_1/xin[93] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[94]), .Q(\modmult_1/xin[94] ) );
  DFF \modmult_1/xreg_reg[93]  ( .D(\modmult_1/xin[92] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[93]), .Q(\modmult_1/xin[93] ) );
  DFF \modmult_1/xreg_reg[92]  ( .D(\modmult_1/xin[91] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[92]), .Q(\modmult_1/xin[92] ) );
  DFF \modmult_1/xreg_reg[91]  ( .D(\modmult_1/xin[90] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[91]), .Q(\modmult_1/xin[91] ) );
  DFF \modmult_1/xreg_reg[90]  ( .D(\modmult_1/xin[89] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[90]), .Q(\modmult_1/xin[90] ) );
  DFF \modmult_1/xreg_reg[89]  ( .D(\modmult_1/xin[88] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[89]), .Q(\modmult_1/xin[89] ) );
  DFF \modmult_1/xreg_reg[88]  ( .D(\modmult_1/xin[87] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[88]), .Q(\modmult_1/xin[88] ) );
  DFF \modmult_1/xreg_reg[87]  ( .D(\modmult_1/xin[86] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[87]), .Q(\modmult_1/xin[87] ) );
  DFF \modmult_1/xreg_reg[86]  ( .D(\modmult_1/xin[85] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[86]), .Q(\modmult_1/xin[86] ) );
  DFF \modmult_1/xreg_reg[85]  ( .D(\modmult_1/xin[84] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[85]), .Q(\modmult_1/xin[85] ) );
  DFF \modmult_1/xreg_reg[84]  ( .D(\modmult_1/xin[83] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[84]), .Q(\modmult_1/xin[84] ) );
  DFF \modmult_1/xreg_reg[83]  ( .D(\modmult_1/xin[82] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[83]), .Q(\modmult_1/xin[83] ) );
  DFF \modmult_1/xreg_reg[82]  ( .D(\modmult_1/xin[81] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[82]), .Q(\modmult_1/xin[82] ) );
  DFF \modmult_1/xreg_reg[81]  ( .D(\modmult_1/xin[80] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[81]), .Q(\modmult_1/xin[81] ) );
  DFF \modmult_1/xreg_reg[80]  ( .D(\modmult_1/xin[79] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[80]), .Q(\modmult_1/xin[80] ) );
  DFF \modmult_1/xreg_reg[79]  ( .D(\modmult_1/xin[78] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[79]), .Q(\modmult_1/xin[79] ) );
  DFF \modmult_1/xreg_reg[78]  ( .D(\modmult_1/xin[77] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[78]), .Q(\modmult_1/xin[78] ) );
  DFF \modmult_1/xreg_reg[77]  ( .D(\modmult_1/xin[76] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[77]), .Q(\modmult_1/xin[77] ) );
  DFF \modmult_1/xreg_reg[76]  ( .D(\modmult_1/xin[75] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[76]), .Q(\modmult_1/xin[76] ) );
  DFF \modmult_1/xreg_reg[75]  ( .D(\modmult_1/xin[74] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[75]), .Q(\modmult_1/xin[75] ) );
  DFF \modmult_1/xreg_reg[74]  ( .D(\modmult_1/xin[73] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[74]), .Q(\modmult_1/xin[74] ) );
  DFF \modmult_1/xreg_reg[73]  ( .D(\modmult_1/xin[72] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[73]), .Q(\modmult_1/xin[73] ) );
  DFF \modmult_1/xreg_reg[72]  ( .D(\modmult_1/xin[71] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[72]), .Q(\modmult_1/xin[72] ) );
  DFF \modmult_1/xreg_reg[71]  ( .D(\modmult_1/xin[70] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[71]), .Q(\modmult_1/xin[71] ) );
  DFF \modmult_1/xreg_reg[70]  ( .D(\modmult_1/xin[69] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[70]), .Q(\modmult_1/xin[70] ) );
  DFF \modmult_1/xreg_reg[69]  ( .D(\modmult_1/xin[68] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[69]), .Q(\modmult_1/xin[69] ) );
  DFF \modmult_1/xreg_reg[68]  ( .D(\modmult_1/xin[67] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[68]), .Q(\modmult_1/xin[68] ) );
  DFF \modmult_1/xreg_reg[67]  ( .D(\modmult_1/xin[66] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[67]), .Q(\modmult_1/xin[67] ) );
  DFF \modmult_1/xreg_reg[66]  ( .D(\modmult_1/xin[65] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[66]), .Q(\modmult_1/xin[66] ) );
  DFF \modmult_1/xreg_reg[65]  ( .D(\modmult_1/xin[64] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[65]), .Q(\modmult_1/xin[65] ) );
  DFF \modmult_1/xreg_reg[64]  ( .D(\modmult_1/xin[63] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[64]), .Q(\modmult_1/xin[64] ) );
  DFF \modmult_1/xreg_reg[63]  ( .D(\modmult_1/xin[62] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[63]), .Q(\modmult_1/xin[63] ) );
  DFF \modmult_1/xreg_reg[62]  ( .D(\modmult_1/xin[61] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[62]), .Q(\modmult_1/xin[62] ) );
  DFF \modmult_1/xreg_reg[61]  ( .D(\modmult_1/xin[60] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[61]), .Q(\modmult_1/xin[61] ) );
  DFF \modmult_1/xreg_reg[60]  ( .D(\modmult_1/xin[59] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[60]), .Q(\modmult_1/xin[60] ) );
  DFF \modmult_1/xreg_reg[59]  ( .D(\modmult_1/xin[58] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[59]), .Q(\modmult_1/xin[59] ) );
  DFF \modmult_1/xreg_reg[58]  ( .D(\modmult_1/xin[57] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[58]), .Q(\modmult_1/xin[58] ) );
  DFF \modmult_1/xreg_reg[57]  ( .D(\modmult_1/xin[56] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[57]), .Q(\modmult_1/xin[57] ) );
  DFF \modmult_1/xreg_reg[56]  ( .D(\modmult_1/xin[55] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[56]), .Q(\modmult_1/xin[56] ) );
  DFF \modmult_1/xreg_reg[55]  ( .D(\modmult_1/xin[54] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[55]), .Q(\modmult_1/xin[55] ) );
  DFF \modmult_1/xreg_reg[54]  ( .D(\modmult_1/xin[53] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[54]), .Q(\modmult_1/xin[54] ) );
  DFF \modmult_1/xreg_reg[53]  ( .D(\modmult_1/xin[52] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[53]), .Q(\modmult_1/xin[53] ) );
  DFF \modmult_1/xreg_reg[52]  ( .D(\modmult_1/xin[51] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[52]), .Q(\modmult_1/xin[52] ) );
  DFF \modmult_1/xreg_reg[51]  ( .D(\modmult_1/xin[50] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[51]), .Q(\modmult_1/xin[51] ) );
  DFF \modmult_1/xreg_reg[50]  ( .D(\modmult_1/xin[49] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[50]), .Q(\modmult_1/xin[50] ) );
  DFF \modmult_1/xreg_reg[49]  ( .D(\modmult_1/xin[48] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[49]), .Q(\modmult_1/xin[49] ) );
  DFF \modmult_1/xreg_reg[48]  ( .D(\modmult_1/xin[47] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[48]), .Q(\modmult_1/xin[48] ) );
  DFF \modmult_1/xreg_reg[47]  ( .D(\modmult_1/xin[46] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[47]), .Q(\modmult_1/xin[47] ) );
  DFF \modmult_1/xreg_reg[46]  ( .D(\modmult_1/xin[45] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[46]), .Q(\modmult_1/xin[46] ) );
  DFF \modmult_1/xreg_reg[45]  ( .D(\modmult_1/xin[44] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[45]), .Q(\modmult_1/xin[45] ) );
  DFF \modmult_1/xreg_reg[44]  ( .D(\modmult_1/xin[43] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[44]), .Q(\modmult_1/xin[44] ) );
  DFF \modmult_1/xreg_reg[43]  ( .D(\modmult_1/xin[42] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[43]), .Q(\modmult_1/xin[43] ) );
  DFF \modmult_1/xreg_reg[42]  ( .D(\modmult_1/xin[41] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[42]), .Q(\modmult_1/xin[42] ) );
  DFF \modmult_1/xreg_reg[41]  ( .D(\modmult_1/xin[40] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[41]), .Q(\modmult_1/xin[41] ) );
  DFF \modmult_1/xreg_reg[40]  ( .D(\modmult_1/xin[39] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[40]), .Q(\modmult_1/xin[40] ) );
  DFF \modmult_1/xreg_reg[39]  ( .D(\modmult_1/xin[38] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[39]), .Q(\modmult_1/xin[39] ) );
  DFF \modmult_1/xreg_reg[38]  ( .D(\modmult_1/xin[37] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[38]), .Q(\modmult_1/xin[38] ) );
  DFF \modmult_1/xreg_reg[37]  ( .D(\modmult_1/xin[36] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[37]), .Q(\modmult_1/xin[37] ) );
  DFF \modmult_1/xreg_reg[36]  ( .D(\modmult_1/xin[35] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[36]), .Q(\modmult_1/xin[36] ) );
  DFF \modmult_1/xreg_reg[35]  ( .D(\modmult_1/xin[34] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[35]), .Q(\modmult_1/xin[35] ) );
  DFF \modmult_1/xreg_reg[34]  ( .D(\modmult_1/xin[33] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[34]), .Q(\modmult_1/xin[34] ) );
  DFF \modmult_1/xreg_reg[33]  ( .D(\modmult_1/xin[32] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[33]), .Q(\modmult_1/xin[33] ) );
  DFF \modmult_1/xreg_reg[32]  ( .D(\modmult_1/xin[31] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[32]), .Q(\modmult_1/xin[32] ) );
  DFF \modmult_1/xreg_reg[31]  ( .D(\modmult_1/xin[30] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[31]), .Q(\modmult_1/xin[31] ) );
  DFF \modmult_1/xreg_reg[30]  ( .D(\modmult_1/xin[29] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[30]), .Q(\modmult_1/xin[30] ) );
  DFF \modmult_1/xreg_reg[29]  ( .D(\modmult_1/xin[28] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[29]), .Q(\modmult_1/xin[29] ) );
  DFF \modmult_1/xreg_reg[28]  ( .D(\modmult_1/xin[27] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[28]), .Q(\modmult_1/xin[28] ) );
  DFF \modmult_1/xreg_reg[27]  ( .D(\modmult_1/xin[26] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[27]), .Q(\modmult_1/xin[27] ) );
  DFF \modmult_1/xreg_reg[26]  ( .D(\modmult_1/xin[25] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[26]), .Q(\modmult_1/xin[26] ) );
  DFF \modmult_1/xreg_reg[25]  ( .D(\modmult_1/xin[24] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[25]), .Q(\modmult_1/xin[25] ) );
  DFF \modmult_1/xreg_reg[24]  ( .D(\modmult_1/xin[23] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[24]), .Q(\modmult_1/xin[24] ) );
  DFF \modmult_1/xreg_reg[23]  ( .D(\modmult_1/xin[22] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[23]), .Q(\modmult_1/xin[23] ) );
  DFF \modmult_1/xreg_reg[22]  ( .D(\modmult_1/xin[21] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[22]), .Q(\modmult_1/xin[22] ) );
  DFF \modmult_1/xreg_reg[21]  ( .D(\modmult_1/xin[20] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[21]), .Q(\modmult_1/xin[21] ) );
  DFF \modmult_1/xreg_reg[20]  ( .D(\modmult_1/xin[19] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[20]), .Q(\modmult_1/xin[20] ) );
  DFF \modmult_1/xreg_reg[19]  ( .D(\modmult_1/xin[18] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[19]), .Q(\modmult_1/xin[19] ) );
  DFF \modmult_1/xreg_reg[18]  ( .D(\modmult_1/xin[17] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[18]), .Q(\modmult_1/xin[18] ) );
  DFF \modmult_1/xreg_reg[17]  ( .D(\modmult_1/xin[16] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[17]), .Q(\modmult_1/xin[17] ) );
  DFF \modmult_1/xreg_reg[16]  ( .D(\modmult_1/xin[15] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[16]), .Q(\modmult_1/xin[16] ) );
  DFF \modmult_1/xreg_reg[15]  ( .D(\modmult_1/xin[14] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[15]), .Q(\modmult_1/xin[15] ) );
  DFF \modmult_1/xreg_reg[14]  ( .D(\modmult_1/xin[13] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[14]), .Q(\modmult_1/xin[14] ) );
  DFF \modmult_1/xreg_reg[13]  ( .D(\modmult_1/xin[12] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[13]), .Q(\modmult_1/xin[13] ) );
  DFF \modmult_1/xreg_reg[12]  ( .D(\modmult_1/xin[11] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[12]), .Q(\modmult_1/xin[12] ) );
  DFF \modmult_1/xreg_reg[11]  ( .D(\modmult_1/xin[10] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[11]), .Q(\modmult_1/xin[11] ) );
  DFF \modmult_1/xreg_reg[10]  ( .D(\modmult_1/xin[9] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[10]), .Q(\modmult_1/xin[10] ) );
  DFF \modmult_1/xreg_reg[9]  ( .D(\modmult_1/xin[8] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[9]), .Q(\modmult_1/xin[9] ) );
  DFF \modmult_1/xreg_reg[8]  ( .D(\modmult_1/xin[7] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[8]), .Q(\modmult_1/xin[8] ) );
  DFF \modmult_1/xreg_reg[7]  ( .D(\modmult_1/xin[6] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[7]), .Q(\modmult_1/xin[7] ) );
  DFF \modmult_1/xreg_reg[6]  ( .D(\modmult_1/xin[5] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[6]), .Q(\modmult_1/xin[6] ) );
  DFF \modmult_1/xreg_reg[5]  ( .D(\modmult_1/xin[4] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[5]), .Q(\modmult_1/xin[5] ) );
  DFF \modmult_1/xreg_reg[4]  ( .D(\modmult_1/xin[3] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[4]), .Q(\modmult_1/xin[4] ) );
  DFF \modmult_1/xreg_reg[3]  ( .D(\modmult_1/xin[2] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[3]), .Q(\modmult_1/xin[3] ) );
  DFF \modmult_1/xreg_reg[2]  ( .D(\modmult_1/xin[1] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[2]), .Q(\modmult_1/xin[2] ) );
  DFF \modmult_1/xreg_reg[1]  ( .D(\modmult_1/xin[0] ), .CLK(clk), .RST(
        start_in[0]), .I(creg[1]), .Q(\modmult_1/xin[1] ) );
  DFF \modmult_1/xreg_reg[0]  ( .D(1'b0), .CLK(clk), .RST(start_in[0]), .I(
        creg[0]), .Q(\modmult_1/xin[0] ) );
  XNOR U1036 ( .A(n1033), .B(n1034), .Z(o[9]) );
  AND U1037 ( .A(n1035), .B(n1036), .Z(n1033) );
  XOR U1038 ( .A(creg[9]), .B(mod_mult_o[9]), .Z(n1036) );
  XNOR U1039 ( .A(n1037), .B(n1038), .Z(o[99]) );
  AND U1040 ( .A(n1035), .B(n1039), .Z(n1037) );
  XOR U1041 ( .A(creg[99]), .B(mod_mult_o[99]), .Z(n1039) );
  XNOR U1042 ( .A(n1040), .B(n1041), .Z(o[999]) );
  AND U1043 ( .A(n1035), .B(n1042), .Z(n1040) );
  XOR U1044 ( .A(creg[999]), .B(mod_mult_o[999]), .Z(n1042) );
  XNOR U1045 ( .A(n1043), .B(n1044), .Z(o[998]) );
  AND U1046 ( .A(n1035), .B(n1045), .Z(n1043) );
  XOR U1047 ( .A(creg[998]), .B(mod_mult_o[998]), .Z(n1045) );
  XNOR U1048 ( .A(n1046), .B(n1047), .Z(o[997]) );
  AND U1049 ( .A(n1035), .B(n1048), .Z(n1046) );
  XOR U1050 ( .A(creg[997]), .B(mod_mult_o[997]), .Z(n1048) );
  XNOR U1051 ( .A(n1049), .B(n1050), .Z(o[996]) );
  AND U1052 ( .A(n1035), .B(n1051), .Z(n1049) );
  XOR U1053 ( .A(creg[996]), .B(mod_mult_o[996]), .Z(n1051) );
  XNOR U1054 ( .A(n1052), .B(n1053), .Z(o[995]) );
  AND U1055 ( .A(n1035), .B(n1054), .Z(n1052) );
  XOR U1056 ( .A(creg[995]), .B(mod_mult_o[995]), .Z(n1054) );
  XNOR U1057 ( .A(n1055), .B(n1056), .Z(o[994]) );
  AND U1058 ( .A(n1035), .B(n1057), .Z(n1055) );
  XOR U1059 ( .A(creg[994]), .B(mod_mult_o[994]), .Z(n1057) );
  XNOR U1060 ( .A(n1058), .B(n1059), .Z(o[993]) );
  AND U1061 ( .A(n1035), .B(n1060), .Z(n1058) );
  XOR U1062 ( .A(creg[993]), .B(mod_mult_o[993]), .Z(n1060) );
  XNOR U1063 ( .A(n1061), .B(n1062), .Z(o[992]) );
  AND U1064 ( .A(n1035), .B(n1063), .Z(n1061) );
  XOR U1065 ( .A(creg[992]), .B(mod_mult_o[992]), .Z(n1063) );
  XNOR U1066 ( .A(n1064), .B(n1065), .Z(o[991]) );
  AND U1067 ( .A(n1035), .B(n1066), .Z(n1064) );
  XOR U1068 ( .A(creg[991]), .B(mod_mult_o[991]), .Z(n1066) );
  XNOR U1069 ( .A(n1067), .B(n1068), .Z(o[990]) );
  AND U1070 ( .A(n1035), .B(n1069), .Z(n1067) );
  XOR U1071 ( .A(creg[990]), .B(mod_mult_o[990]), .Z(n1069) );
  XNOR U1072 ( .A(n1070), .B(n1071), .Z(o[98]) );
  AND U1073 ( .A(n1035), .B(n1072), .Z(n1070) );
  XOR U1074 ( .A(creg[98]), .B(mod_mult_o[98]), .Z(n1072) );
  XNOR U1075 ( .A(n1073), .B(n1074), .Z(o[989]) );
  AND U1076 ( .A(n1035), .B(n1075), .Z(n1073) );
  XOR U1077 ( .A(creg[989]), .B(mod_mult_o[989]), .Z(n1075) );
  XNOR U1078 ( .A(n1076), .B(n1077), .Z(o[988]) );
  AND U1079 ( .A(n1035), .B(n1078), .Z(n1076) );
  XOR U1080 ( .A(creg[988]), .B(mod_mult_o[988]), .Z(n1078) );
  XNOR U1081 ( .A(n1079), .B(n1080), .Z(o[987]) );
  AND U1082 ( .A(n1035), .B(n1081), .Z(n1079) );
  XOR U1083 ( .A(creg[987]), .B(mod_mult_o[987]), .Z(n1081) );
  XNOR U1084 ( .A(n1082), .B(n1083), .Z(o[986]) );
  AND U1085 ( .A(n1035), .B(n1084), .Z(n1082) );
  XOR U1086 ( .A(creg[986]), .B(mod_mult_o[986]), .Z(n1084) );
  XNOR U1087 ( .A(n1085), .B(n1086), .Z(o[985]) );
  AND U1088 ( .A(n1035), .B(n1087), .Z(n1085) );
  XOR U1089 ( .A(creg[985]), .B(mod_mult_o[985]), .Z(n1087) );
  XNOR U1090 ( .A(n1088), .B(n1089), .Z(o[984]) );
  AND U1091 ( .A(n1035), .B(n1090), .Z(n1088) );
  XOR U1092 ( .A(creg[984]), .B(mod_mult_o[984]), .Z(n1090) );
  XNOR U1093 ( .A(n1091), .B(n1092), .Z(o[983]) );
  AND U1094 ( .A(n1035), .B(n1093), .Z(n1091) );
  XOR U1095 ( .A(creg[983]), .B(mod_mult_o[983]), .Z(n1093) );
  XNOR U1096 ( .A(n1094), .B(n1095), .Z(o[982]) );
  AND U1097 ( .A(n1035), .B(n1096), .Z(n1094) );
  XOR U1098 ( .A(creg[982]), .B(mod_mult_o[982]), .Z(n1096) );
  XNOR U1099 ( .A(n1097), .B(n1098), .Z(o[981]) );
  AND U1100 ( .A(n1035), .B(n1099), .Z(n1097) );
  XOR U1101 ( .A(creg[981]), .B(mod_mult_o[981]), .Z(n1099) );
  XNOR U1102 ( .A(n1100), .B(n1101), .Z(o[980]) );
  AND U1103 ( .A(n1035), .B(n1102), .Z(n1100) );
  XOR U1104 ( .A(creg[980]), .B(mod_mult_o[980]), .Z(n1102) );
  XNOR U1105 ( .A(n1103), .B(n1104), .Z(o[97]) );
  AND U1106 ( .A(n1035), .B(n1105), .Z(n1103) );
  XOR U1107 ( .A(creg[97]), .B(mod_mult_o[97]), .Z(n1105) );
  XNOR U1108 ( .A(n1106), .B(n1107), .Z(o[979]) );
  AND U1109 ( .A(n1035), .B(n1108), .Z(n1106) );
  XOR U1110 ( .A(creg[979]), .B(mod_mult_o[979]), .Z(n1108) );
  XNOR U1111 ( .A(n1109), .B(n1110), .Z(o[978]) );
  AND U1112 ( .A(n1035), .B(n1111), .Z(n1109) );
  XOR U1113 ( .A(creg[978]), .B(mod_mult_o[978]), .Z(n1111) );
  XNOR U1114 ( .A(n1112), .B(n1113), .Z(o[977]) );
  AND U1115 ( .A(n1035), .B(n1114), .Z(n1112) );
  XOR U1116 ( .A(creg[977]), .B(mod_mult_o[977]), .Z(n1114) );
  XNOR U1117 ( .A(n1115), .B(n1116), .Z(o[976]) );
  AND U1118 ( .A(n1035), .B(n1117), .Z(n1115) );
  XOR U1119 ( .A(creg[976]), .B(mod_mult_o[976]), .Z(n1117) );
  XNOR U1120 ( .A(n1118), .B(n1119), .Z(o[975]) );
  AND U1121 ( .A(n1035), .B(n1120), .Z(n1118) );
  XOR U1122 ( .A(creg[975]), .B(mod_mult_o[975]), .Z(n1120) );
  XNOR U1123 ( .A(n1121), .B(n1122), .Z(o[974]) );
  AND U1124 ( .A(n1035), .B(n1123), .Z(n1121) );
  XOR U1125 ( .A(creg[974]), .B(mod_mult_o[974]), .Z(n1123) );
  XNOR U1126 ( .A(n1124), .B(n1125), .Z(o[973]) );
  AND U1127 ( .A(n1035), .B(n1126), .Z(n1124) );
  XOR U1128 ( .A(creg[973]), .B(mod_mult_o[973]), .Z(n1126) );
  XNOR U1129 ( .A(n1127), .B(n1128), .Z(o[972]) );
  AND U1130 ( .A(n1035), .B(n1129), .Z(n1127) );
  XOR U1131 ( .A(creg[972]), .B(mod_mult_o[972]), .Z(n1129) );
  XNOR U1132 ( .A(n1130), .B(n1131), .Z(o[971]) );
  AND U1133 ( .A(n1035), .B(n1132), .Z(n1130) );
  XOR U1134 ( .A(creg[971]), .B(mod_mult_o[971]), .Z(n1132) );
  XNOR U1135 ( .A(n1133), .B(n1134), .Z(o[970]) );
  AND U1136 ( .A(n1035), .B(n1135), .Z(n1133) );
  XOR U1137 ( .A(creg[970]), .B(mod_mult_o[970]), .Z(n1135) );
  XNOR U1138 ( .A(n1136), .B(n1137), .Z(o[96]) );
  AND U1139 ( .A(n1035), .B(n1138), .Z(n1136) );
  XOR U1140 ( .A(creg[96]), .B(mod_mult_o[96]), .Z(n1138) );
  XNOR U1141 ( .A(n1139), .B(n1140), .Z(o[969]) );
  AND U1142 ( .A(n1035), .B(n1141), .Z(n1139) );
  XOR U1143 ( .A(creg[969]), .B(mod_mult_o[969]), .Z(n1141) );
  XNOR U1144 ( .A(n1142), .B(n1143), .Z(o[968]) );
  AND U1145 ( .A(n1035), .B(n1144), .Z(n1142) );
  XOR U1146 ( .A(creg[968]), .B(mod_mult_o[968]), .Z(n1144) );
  XNOR U1147 ( .A(n1145), .B(n1146), .Z(o[967]) );
  AND U1148 ( .A(n1035), .B(n1147), .Z(n1145) );
  XOR U1149 ( .A(creg[967]), .B(mod_mult_o[967]), .Z(n1147) );
  XNOR U1150 ( .A(n1148), .B(n1149), .Z(o[966]) );
  AND U1151 ( .A(n1035), .B(n1150), .Z(n1148) );
  XOR U1152 ( .A(creg[966]), .B(mod_mult_o[966]), .Z(n1150) );
  XNOR U1153 ( .A(n1151), .B(n1152), .Z(o[965]) );
  AND U1154 ( .A(n1035), .B(n1153), .Z(n1151) );
  XOR U1155 ( .A(creg[965]), .B(mod_mult_o[965]), .Z(n1153) );
  XNOR U1156 ( .A(n1154), .B(n1155), .Z(o[964]) );
  AND U1157 ( .A(n1035), .B(n1156), .Z(n1154) );
  XOR U1158 ( .A(creg[964]), .B(mod_mult_o[964]), .Z(n1156) );
  XNOR U1159 ( .A(n1157), .B(n1158), .Z(o[963]) );
  AND U1160 ( .A(n1035), .B(n1159), .Z(n1157) );
  XOR U1161 ( .A(creg[963]), .B(mod_mult_o[963]), .Z(n1159) );
  XNOR U1162 ( .A(n1160), .B(n1161), .Z(o[962]) );
  AND U1163 ( .A(n1035), .B(n1162), .Z(n1160) );
  XOR U1164 ( .A(creg[962]), .B(mod_mult_o[962]), .Z(n1162) );
  XNOR U1165 ( .A(n1163), .B(n1164), .Z(o[961]) );
  AND U1166 ( .A(n1035), .B(n1165), .Z(n1163) );
  XOR U1167 ( .A(creg[961]), .B(mod_mult_o[961]), .Z(n1165) );
  XNOR U1168 ( .A(n1166), .B(n1167), .Z(o[960]) );
  AND U1169 ( .A(n1035), .B(n1168), .Z(n1166) );
  XOR U1170 ( .A(creg[960]), .B(mod_mult_o[960]), .Z(n1168) );
  XNOR U1171 ( .A(n1169), .B(n1170), .Z(o[95]) );
  AND U1172 ( .A(n1035), .B(n1171), .Z(n1169) );
  XOR U1173 ( .A(creg[95]), .B(mod_mult_o[95]), .Z(n1171) );
  XNOR U1174 ( .A(n1172), .B(n1173), .Z(o[959]) );
  AND U1175 ( .A(n1035), .B(n1174), .Z(n1172) );
  XOR U1176 ( .A(creg[959]), .B(mod_mult_o[959]), .Z(n1174) );
  XNOR U1177 ( .A(n1175), .B(n1176), .Z(o[958]) );
  AND U1178 ( .A(n1035), .B(n1177), .Z(n1175) );
  XOR U1179 ( .A(creg[958]), .B(mod_mult_o[958]), .Z(n1177) );
  XNOR U1180 ( .A(n1178), .B(n1179), .Z(o[957]) );
  AND U1181 ( .A(n1035), .B(n1180), .Z(n1178) );
  XOR U1182 ( .A(creg[957]), .B(mod_mult_o[957]), .Z(n1180) );
  XNOR U1183 ( .A(n1181), .B(n1182), .Z(o[956]) );
  AND U1184 ( .A(n1035), .B(n1183), .Z(n1181) );
  XOR U1185 ( .A(creg[956]), .B(mod_mult_o[956]), .Z(n1183) );
  XNOR U1186 ( .A(n1184), .B(n1185), .Z(o[955]) );
  AND U1187 ( .A(n1035), .B(n1186), .Z(n1184) );
  XOR U1188 ( .A(creg[955]), .B(mod_mult_o[955]), .Z(n1186) );
  XNOR U1189 ( .A(n1187), .B(n1188), .Z(o[954]) );
  AND U1190 ( .A(n1035), .B(n1189), .Z(n1187) );
  XOR U1191 ( .A(creg[954]), .B(mod_mult_o[954]), .Z(n1189) );
  XNOR U1192 ( .A(n1190), .B(n1191), .Z(o[953]) );
  AND U1193 ( .A(n1035), .B(n1192), .Z(n1190) );
  XOR U1194 ( .A(creg[953]), .B(mod_mult_o[953]), .Z(n1192) );
  XNOR U1195 ( .A(n1193), .B(n1194), .Z(o[952]) );
  AND U1196 ( .A(n1035), .B(n1195), .Z(n1193) );
  XOR U1197 ( .A(creg[952]), .B(mod_mult_o[952]), .Z(n1195) );
  XNOR U1198 ( .A(n1196), .B(n1197), .Z(o[951]) );
  AND U1199 ( .A(n1035), .B(n1198), .Z(n1196) );
  XOR U1200 ( .A(creg[951]), .B(mod_mult_o[951]), .Z(n1198) );
  XNOR U1201 ( .A(n1199), .B(n1200), .Z(o[950]) );
  AND U1202 ( .A(n1035), .B(n1201), .Z(n1199) );
  XOR U1203 ( .A(creg[950]), .B(mod_mult_o[950]), .Z(n1201) );
  XNOR U1204 ( .A(n1202), .B(n1203), .Z(o[94]) );
  AND U1205 ( .A(n1035), .B(n1204), .Z(n1202) );
  XOR U1206 ( .A(creg[94]), .B(mod_mult_o[94]), .Z(n1204) );
  XNOR U1207 ( .A(n1205), .B(n1206), .Z(o[949]) );
  AND U1208 ( .A(n1035), .B(n1207), .Z(n1205) );
  XOR U1209 ( .A(creg[949]), .B(mod_mult_o[949]), .Z(n1207) );
  XNOR U1210 ( .A(n1208), .B(n1209), .Z(o[948]) );
  AND U1211 ( .A(n1035), .B(n1210), .Z(n1208) );
  XOR U1212 ( .A(creg[948]), .B(mod_mult_o[948]), .Z(n1210) );
  XNOR U1213 ( .A(n1211), .B(n1212), .Z(o[947]) );
  AND U1214 ( .A(n1035), .B(n1213), .Z(n1211) );
  XOR U1215 ( .A(creg[947]), .B(mod_mult_o[947]), .Z(n1213) );
  XNOR U1216 ( .A(n1214), .B(n1215), .Z(o[946]) );
  AND U1217 ( .A(n1035), .B(n1216), .Z(n1214) );
  XOR U1218 ( .A(creg[946]), .B(mod_mult_o[946]), .Z(n1216) );
  XNOR U1219 ( .A(n1217), .B(n1218), .Z(o[945]) );
  AND U1220 ( .A(n1035), .B(n1219), .Z(n1217) );
  XOR U1221 ( .A(creg[945]), .B(mod_mult_o[945]), .Z(n1219) );
  XNOR U1222 ( .A(n1220), .B(n1221), .Z(o[944]) );
  AND U1223 ( .A(n1035), .B(n1222), .Z(n1220) );
  XOR U1224 ( .A(creg[944]), .B(mod_mult_o[944]), .Z(n1222) );
  XNOR U1225 ( .A(n1223), .B(n1224), .Z(o[943]) );
  AND U1226 ( .A(n1035), .B(n1225), .Z(n1223) );
  XOR U1227 ( .A(creg[943]), .B(mod_mult_o[943]), .Z(n1225) );
  XNOR U1228 ( .A(n1226), .B(n1227), .Z(o[942]) );
  AND U1229 ( .A(n1035), .B(n1228), .Z(n1226) );
  XOR U1230 ( .A(creg[942]), .B(mod_mult_o[942]), .Z(n1228) );
  XNOR U1231 ( .A(n1229), .B(n1230), .Z(o[941]) );
  AND U1232 ( .A(n1035), .B(n1231), .Z(n1229) );
  XOR U1233 ( .A(creg[941]), .B(mod_mult_o[941]), .Z(n1231) );
  XNOR U1234 ( .A(n1232), .B(n1233), .Z(o[940]) );
  AND U1235 ( .A(n1035), .B(n1234), .Z(n1232) );
  XOR U1236 ( .A(creg[940]), .B(mod_mult_o[940]), .Z(n1234) );
  XNOR U1237 ( .A(n1235), .B(n1236), .Z(o[93]) );
  AND U1238 ( .A(n1035), .B(n1237), .Z(n1235) );
  XOR U1239 ( .A(creg[93]), .B(mod_mult_o[93]), .Z(n1237) );
  XNOR U1240 ( .A(n1238), .B(n1239), .Z(o[939]) );
  AND U1241 ( .A(n1035), .B(n1240), .Z(n1238) );
  XOR U1242 ( .A(creg[939]), .B(mod_mult_o[939]), .Z(n1240) );
  XNOR U1243 ( .A(n1241), .B(n1242), .Z(o[938]) );
  AND U1244 ( .A(n1035), .B(n1243), .Z(n1241) );
  XOR U1245 ( .A(creg[938]), .B(mod_mult_o[938]), .Z(n1243) );
  XNOR U1246 ( .A(n1244), .B(n1245), .Z(o[937]) );
  AND U1247 ( .A(n1035), .B(n1246), .Z(n1244) );
  XOR U1248 ( .A(creg[937]), .B(mod_mult_o[937]), .Z(n1246) );
  XNOR U1249 ( .A(n1247), .B(n1248), .Z(o[936]) );
  AND U1250 ( .A(n1035), .B(n1249), .Z(n1247) );
  XOR U1251 ( .A(creg[936]), .B(mod_mult_o[936]), .Z(n1249) );
  XNOR U1252 ( .A(n1250), .B(n1251), .Z(o[935]) );
  AND U1253 ( .A(n1035), .B(n1252), .Z(n1250) );
  XOR U1254 ( .A(creg[935]), .B(mod_mult_o[935]), .Z(n1252) );
  XNOR U1255 ( .A(n1253), .B(n1254), .Z(o[934]) );
  AND U1256 ( .A(n1035), .B(n1255), .Z(n1253) );
  XOR U1257 ( .A(creg[934]), .B(mod_mult_o[934]), .Z(n1255) );
  XNOR U1258 ( .A(n1256), .B(n1257), .Z(o[933]) );
  AND U1259 ( .A(n1035), .B(n1258), .Z(n1256) );
  XOR U1260 ( .A(creg[933]), .B(mod_mult_o[933]), .Z(n1258) );
  XNOR U1261 ( .A(n1259), .B(n1260), .Z(o[932]) );
  AND U1262 ( .A(n1035), .B(n1261), .Z(n1259) );
  XOR U1263 ( .A(creg[932]), .B(mod_mult_o[932]), .Z(n1261) );
  XNOR U1264 ( .A(n1262), .B(n1263), .Z(o[931]) );
  AND U1265 ( .A(n1035), .B(n1264), .Z(n1262) );
  XOR U1266 ( .A(creg[931]), .B(mod_mult_o[931]), .Z(n1264) );
  XNOR U1267 ( .A(n1265), .B(n1266), .Z(o[930]) );
  AND U1268 ( .A(n1035), .B(n1267), .Z(n1265) );
  XOR U1269 ( .A(creg[930]), .B(mod_mult_o[930]), .Z(n1267) );
  XNOR U1270 ( .A(n1268), .B(n1269), .Z(o[92]) );
  AND U1271 ( .A(n1035), .B(n1270), .Z(n1268) );
  XOR U1272 ( .A(creg[92]), .B(mod_mult_o[92]), .Z(n1270) );
  XNOR U1273 ( .A(n1271), .B(n1272), .Z(o[929]) );
  AND U1274 ( .A(n1035), .B(n1273), .Z(n1271) );
  XOR U1275 ( .A(creg[929]), .B(mod_mult_o[929]), .Z(n1273) );
  XNOR U1276 ( .A(n1274), .B(n1275), .Z(o[928]) );
  AND U1277 ( .A(n1035), .B(n1276), .Z(n1274) );
  XOR U1278 ( .A(creg[928]), .B(mod_mult_o[928]), .Z(n1276) );
  XNOR U1279 ( .A(n1277), .B(n1278), .Z(o[927]) );
  AND U1280 ( .A(n1035), .B(n1279), .Z(n1277) );
  XOR U1281 ( .A(creg[927]), .B(mod_mult_o[927]), .Z(n1279) );
  XNOR U1282 ( .A(n1280), .B(n1281), .Z(o[926]) );
  AND U1283 ( .A(n1035), .B(n1282), .Z(n1280) );
  XOR U1284 ( .A(creg[926]), .B(mod_mult_o[926]), .Z(n1282) );
  XNOR U1285 ( .A(n1283), .B(n1284), .Z(o[925]) );
  AND U1286 ( .A(n1035), .B(n1285), .Z(n1283) );
  XOR U1287 ( .A(creg[925]), .B(mod_mult_o[925]), .Z(n1285) );
  XNOR U1288 ( .A(n1286), .B(n1287), .Z(o[924]) );
  AND U1289 ( .A(n1035), .B(n1288), .Z(n1286) );
  XOR U1290 ( .A(creg[924]), .B(mod_mult_o[924]), .Z(n1288) );
  XNOR U1291 ( .A(n1289), .B(n1290), .Z(o[923]) );
  AND U1292 ( .A(n1035), .B(n1291), .Z(n1289) );
  XOR U1293 ( .A(creg[923]), .B(mod_mult_o[923]), .Z(n1291) );
  XNOR U1294 ( .A(n1292), .B(n1293), .Z(o[922]) );
  AND U1295 ( .A(n1035), .B(n1294), .Z(n1292) );
  XOR U1296 ( .A(creg[922]), .B(mod_mult_o[922]), .Z(n1294) );
  XNOR U1297 ( .A(n1295), .B(n1296), .Z(o[921]) );
  AND U1298 ( .A(n1035), .B(n1297), .Z(n1295) );
  XOR U1299 ( .A(creg[921]), .B(mod_mult_o[921]), .Z(n1297) );
  XNOR U1300 ( .A(n1298), .B(n1299), .Z(o[920]) );
  AND U1301 ( .A(n1035), .B(n1300), .Z(n1298) );
  XOR U1302 ( .A(creg[920]), .B(mod_mult_o[920]), .Z(n1300) );
  XNOR U1303 ( .A(n1301), .B(n1302), .Z(o[91]) );
  AND U1304 ( .A(n1035), .B(n1303), .Z(n1301) );
  XOR U1305 ( .A(creg[91]), .B(mod_mult_o[91]), .Z(n1303) );
  XNOR U1306 ( .A(n1304), .B(n1305), .Z(o[919]) );
  AND U1307 ( .A(n1035), .B(n1306), .Z(n1304) );
  XOR U1308 ( .A(creg[919]), .B(mod_mult_o[919]), .Z(n1306) );
  XNOR U1309 ( .A(n1307), .B(n1308), .Z(o[918]) );
  AND U1310 ( .A(n1035), .B(n1309), .Z(n1307) );
  XOR U1311 ( .A(creg[918]), .B(mod_mult_o[918]), .Z(n1309) );
  XNOR U1312 ( .A(n1310), .B(n1311), .Z(o[917]) );
  AND U1313 ( .A(n1035), .B(n1312), .Z(n1310) );
  XOR U1314 ( .A(creg[917]), .B(mod_mult_o[917]), .Z(n1312) );
  XNOR U1315 ( .A(n1313), .B(n1314), .Z(o[916]) );
  AND U1316 ( .A(n1035), .B(n1315), .Z(n1313) );
  XOR U1317 ( .A(creg[916]), .B(mod_mult_o[916]), .Z(n1315) );
  XNOR U1318 ( .A(n1316), .B(n1317), .Z(o[915]) );
  AND U1319 ( .A(n1035), .B(n1318), .Z(n1316) );
  XOR U1320 ( .A(creg[915]), .B(mod_mult_o[915]), .Z(n1318) );
  XNOR U1321 ( .A(n1319), .B(n1320), .Z(o[914]) );
  AND U1322 ( .A(n1035), .B(n1321), .Z(n1319) );
  XOR U1323 ( .A(creg[914]), .B(mod_mult_o[914]), .Z(n1321) );
  XNOR U1324 ( .A(n1322), .B(n1323), .Z(o[913]) );
  AND U1325 ( .A(n1035), .B(n1324), .Z(n1322) );
  XOR U1326 ( .A(creg[913]), .B(mod_mult_o[913]), .Z(n1324) );
  XNOR U1327 ( .A(n1325), .B(n1326), .Z(o[912]) );
  AND U1328 ( .A(n1035), .B(n1327), .Z(n1325) );
  XOR U1329 ( .A(creg[912]), .B(mod_mult_o[912]), .Z(n1327) );
  XNOR U1330 ( .A(n1328), .B(n1329), .Z(o[911]) );
  AND U1331 ( .A(n1035), .B(n1330), .Z(n1328) );
  XOR U1332 ( .A(creg[911]), .B(mod_mult_o[911]), .Z(n1330) );
  XNOR U1333 ( .A(n1331), .B(n1332), .Z(o[910]) );
  AND U1334 ( .A(n1035), .B(n1333), .Z(n1331) );
  XOR U1335 ( .A(creg[910]), .B(mod_mult_o[910]), .Z(n1333) );
  XNOR U1336 ( .A(n1334), .B(n1335), .Z(o[90]) );
  AND U1337 ( .A(n1035), .B(n1336), .Z(n1334) );
  XOR U1338 ( .A(creg[90]), .B(mod_mult_o[90]), .Z(n1336) );
  XNOR U1339 ( .A(n1337), .B(n1338), .Z(o[909]) );
  AND U1340 ( .A(n1035), .B(n1339), .Z(n1337) );
  XOR U1341 ( .A(creg[909]), .B(mod_mult_o[909]), .Z(n1339) );
  XNOR U1342 ( .A(n1340), .B(n1341), .Z(o[908]) );
  AND U1343 ( .A(n1035), .B(n1342), .Z(n1340) );
  XOR U1344 ( .A(creg[908]), .B(mod_mult_o[908]), .Z(n1342) );
  XNOR U1345 ( .A(n1343), .B(n1344), .Z(o[907]) );
  AND U1346 ( .A(n1035), .B(n1345), .Z(n1343) );
  XOR U1347 ( .A(creg[907]), .B(mod_mult_o[907]), .Z(n1345) );
  XNOR U1348 ( .A(n1346), .B(n1347), .Z(o[906]) );
  AND U1349 ( .A(n1035), .B(n1348), .Z(n1346) );
  XOR U1350 ( .A(creg[906]), .B(mod_mult_o[906]), .Z(n1348) );
  XNOR U1351 ( .A(n1349), .B(n1350), .Z(o[905]) );
  AND U1352 ( .A(n1035), .B(n1351), .Z(n1349) );
  XOR U1353 ( .A(creg[905]), .B(mod_mult_o[905]), .Z(n1351) );
  XNOR U1354 ( .A(n1352), .B(n1353), .Z(o[904]) );
  AND U1355 ( .A(n1035), .B(n1354), .Z(n1352) );
  XOR U1356 ( .A(creg[904]), .B(mod_mult_o[904]), .Z(n1354) );
  XNOR U1357 ( .A(n1355), .B(n1356), .Z(o[903]) );
  AND U1358 ( .A(n1035), .B(n1357), .Z(n1355) );
  XOR U1359 ( .A(creg[903]), .B(mod_mult_o[903]), .Z(n1357) );
  XNOR U1360 ( .A(n1358), .B(n1359), .Z(o[902]) );
  AND U1361 ( .A(n1035), .B(n1360), .Z(n1358) );
  XOR U1362 ( .A(creg[902]), .B(mod_mult_o[902]), .Z(n1360) );
  XNOR U1363 ( .A(n1361), .B(n1362), .Z(o[901]) );
  AND U1364 ( .A(n1035), .B(n1363), .Z(n1361) );
  XOR U1365 ( .A(creg[901]), .B(mod_mult_o[901]), .Z(n1363) );
  XNOR U1366 ( .A(n1364), .B(n1365), .Z(o[900]) );
  AND U1367 ( .A(n1035), .B(n1366), .Z(n1364) );
  XOR U1368 ( .A(creg[900]), .B(mod_mult_o[900]), .Z(n1366) );
  XNOR U1369 ( .A(n1367), .B(n1368), .Z(o[8]) );
  AND U1370 ( .A(n1035), .B(n1369), .Z(n1367) );
  XOR U1371 ( .A(creg[8]), .B(mod_mult_o[8]), .Z(n1369) );
  XNOR U1372 ( .A(n1370), .B(n1371), .Z(o[89]) );
  AND U1373 ( .A(n1035), .B(n1372), .Z(n1370) );
  XOR U1374 ( .A(creg[89]), .B(mod_mult_o[89]), .Z(n1372) );
  XNOR U1375 ( .A(n1373), .B(n1374), .Z(o[899]) );
  AND U1376 ( .A(n1035), .B(n1375), .Z(n1373) );
  XOR U1377 ( .A(creg[899]), .B(mod_mult_o[899]), .Z(n1375) );
  XNOR U1378 ( .A(n1376), .B(n1377), .Z(o[898]) );
  AND U1379 ( .A(n1035), .B(n1378), .Z(n1376) );
  XOR U1380 ( .A(creg[898]), .B(mod_mult_o[898]), .Z(n1378) );
  XNOR U1381 ( .A(n1379), .B(n1380), .Z(o[897]) );
  AND U1382 ( .A(n1035), .B(n1381), .Z(n1379) );
  XOR U1383 ( .A(creg[897]), .B(mod_mult_o[897]), .Z(n1381) );
  XNOR U1384 ( .A(n1382), .B(n1383), .Z(o[896]) );
  AND U1385 ( .A(n1035), .B(n1384), .Z(n1382) );
  XOR U1386 ( .A(creg[896]), .B(mod_mult_o[896]), .Z(n1384) );
  XNOR U1387 ( .A(n1385), .B(n1386), .Z(o[895]) );
  AND U1388 ( .A(n1035), .B(n1387), .Z(n1385) );
  XOR U1389 ( .A(creg[895]), .B(mod_mult_o[895]), .Z(n1387) );
  XNOR U1390 ( .A(n1388), .B(n1389), .Z(o[894]) );
  AND U1391 ( .A(n1035), .B(n1390), .Z(n1388) );
  XOR U1392 ( .A(creg[894]), .B(mod_mult_o[894]), .Z(n1390) );
  XNOR U1393 ( .A(n1391), .B(n1392), .Z(o[893]) );
  AND U1394 ( .A(n1035), .B(n1393), .Z(n1391) );
  XOR U1395 ( .A(creg[893]), .B(mod_mult_o[893]), .Z(n1393) );
  XNOR U1396 ( .A(n1394), .B(n1395), .Z(o[892]) );
  AND U1397 ( .A(n1035), .B(n1396), .Z(n1394) );
  XOR U1398 ( .A(creg[892]), .B(mod_mult_o[892]), .Z(n1396) );
  XNOR U1399 ( .A(n1397), .B(n1398), .Z(o[891]) );
  AND U1400 ( .A(n1035), .B(n1399), .Z(n1397) );
  XOR U1401 ( .A(creg[891]), .B(mod_mult_o[891]), .Z(n1399) );
  XNOR U1402 ( .A(n1400), .B(n1401), .Z(o[890]) );
  AND U1403 ( .A(n1035), .B(n1402), .Z(n1400) );
  XOR U1404 ( .A(creg[890]), .B(mod_mult_o[890]), .Z(n1402) );
  XNOR U1405 ( .A(n1403), .B(n1404), .Z(o[88]) );
  AND U1406 ( .A(n1035), .B(n1405), .Z(n1403) );
  XOR U1407 ( .A(creg[88]), .B(mod_mult_o[88]), .Z(n1405) );
  XNOR U1408 ( .A(n1406), .B(n1407), .Z(o[889]) );
  AND U1409 ( .A(n1035), .B(n1408), .Z(n1406) );
  XOR U1410 ( .A(creg[889]), .B(mod_mult_o[889]), .Z(n1408) );
  XNOR U1411 ( .A(n1409), .B(n1410), .Z(o[888]) );
  AND U1412 ( .A(n1035), .B(n1411), .Z(n1409) );
  XOR U1413 ( .A(creg[888]), .B(mod_mult_o[888]), .Z(n1411) );
  XNOR U1414 ( .A(n1412), .B(n1413), .Z(o[887]) );
  AND U1415 ( .A(n1035), .B(n1414), .Z(n1412) );
  XOR U1416 ( .A(creg[887]), .B(mod_mult_o[887]), .Z(n1414) );
  XNOR U1417 ( .A(n1415), .B(n1416), .Z(o[886]) );
  AND U1418 ( .A(n1035), .B(n1417), .Z(n1415) );
  XOR U1419 ( .A(creg[886]), .B(mod_mult_o[886]), .Z(n1417) );
  XNOR U1420 ( .A(n1418), .B(n1419), .Z(o[885]) );
  AND U1421 ( .A(n1035), .B(n1420), .Z(n1418) );
  XOR U1422 ( .A(creg[885]), .B(mod_mult_o[885]), .Z(n1420) );
  XNOR U1423 ( .A(n1421), .B(n1422), .Z(o[884]) );
  AND U1424 ( .A(n1035), .B(n1423), .Z(n1421) );
  XOR U1425 ( .A(creg[884]), .B(mod_mult_o[884]), .Z(n1423) );
  XNOR U1426 ( .A(n1424), .B(n1425), .Z(o[883]) );
  AND U1427 ( .A(n1035), .B(n1426), .Z(n1424) );
  XOR U1428 ( .A(creg[883]), .B(mod_mult_o[883]), .Z(n1426) );
  XNOR U1429 ( .A(n1427), .B(n1428), .Z(o[882]) );
  AND U1430 ( .A(n1035), .B(n1429), .Z(n1427) );
  XOR U1431 ( .A(creg[882]), .B(mod_mult_o[882]), .Z(n1429) );
  XNOR U1432 ( .A(n1430), .B(n1431), .Z(o[881]) );
  AND U1433 ( .A(n1035), .B(n1432), .Z(n1430) );
  XOR U1434 ( .A(creg[881]), .B(mod_mult_o[881]), .Z(n1432) );
  XNOR U1435 ( .A(n1433), .B(n1434), .Z(o[880]) );
  AND U1436 ( .A(n1035), .B(n1435), .Z(n1433) );
  XOR U1437 ( .A(creg[880]), .B(mod_mult_o[880]), .Z(n1435) );
  XNOR U1438 ( .A(n1436), .B(n1437), .Z(o[87]) );
  AND U1439 ( .A(n1035), .B(n1438), .Z(n1436) );
  XOR U1440 ( .A(creg[87]), .B(mod_mult_o[87]), .Z(n1438) );
  XNOR U1441 ( .A(n1439), .B(n1440), .Z(o[879]) );
  AND U1442 ( .A(n1035), .B(n1441), .Z(n1439) );
  XOR U1443 ( .A(creg[879]), .B(mod_mult_o[879]), .Z(n1441) );
  XNOR U1444 ( .A(n1442), .B(n1443), .Z(o[878]) );
  AND U1445 ( .A(n1035), .B(n1444), .Z(n1442) );
  XOR U1446 ( .A(creg[878]), .B(mod_mult_o[878]), .Z(n1444) );
  XNOR U1447 ( .A(n1445), .B(n1446), .Z(o[877]) );
  AND U1448 ( .A(n1035), .B(n1447), .Z(n1445) );
  XOR U1449 ( .A(creg[877]), .B(mod_mult_o[877]), .Z(n1447) );
  XNOR U1450 ( .A(n1448), .B(n1449), .Z(o[876]) );
  AND U1451 ( .A(n1035), .B(n1450), .Z(n1448) );
  XOR U1452 ( .A(creg[876]), .B(mod_mult_o[876]), .Z(n1450) );
  XNOR U1453 ( .A(n1451), .B(n1452), .Z(o[875]) );
  AND U1454 ( .A(n1035), .B(n1453), .Z(n1451) );
  XOR U1455 ( .A(creg[875]), .B(mod_mult_o[875]), .Z(n1453) );
  XNOR U1456 ( .A(n1454), .B(n1455), .Z(o[874]) );
  AND U1457 ( .A(n1035), .B(n1456), .Z(n1454) );
  XOR U1458 ( .A(creg[874]), .B(mod_mult_o[874]), .Z(n1456) );
  XNOR U1459 ( .A(n1457), .B(n1458), .Z(o[873]) );
  AND U1460 ( .A(n1035), .B(n1459), .Z(n1457) );
  XOR U1461 ( .A(creg[873]), .B(mod_mult_o[873]), .Z(n1459) );
  XNOR U1462 ( .A(n1460), .B(n1461), .Z(o[872]) );
  AND U1463 ( .A(n1035), .B(n1462), .Z(n1460) );
  XOR U1464 ( .A(creg[872]), .B(mod_mult_o[872]), .Z(n1462) );
  XNOR U1465 ( .A(n1463), .B(n1464), .Z(o[871]) );
  AND U1466 ( .A(n1035), .B(n1465), .Z(n1463) );
  XOR U1467 ( .A(creg[871]), .B(mod_mult_o[871]), .Z(n1465) );
  XNOR U1468 ( .A(n1466), .B(n1467), .Z(o[870]) );
  AND U1469 ( .A(n1035), .B(n1468), .Z(n1466) );
  XOR U1470 ( .A(creg[870]), .B(mod_mult_o[870]), .Z(n1468) );
  XNOR U1471 ( .A(n1469), .B(n1470), .Z(o[86]) );
  AND U1472 ( .A(n1035), .B(n1471), .Z(n1469) );
  XOR U1473 ( .A(creg[86]), .B(mod_mult_o[86]), .Z(n1471) );
  XNOR U1474 ( .A(n1472), .B(n1473), .Z(o[869]) );
  AND U1475 ( .A(n1035), .B(n1474), .Z(n1472) );
  XOR U1476 ( .A(creg[869]), .B(mod_mult_o[869]), .Z(n1474) );
  XNOR U1477 ( .A(n1475), .B(n1476), .Z(o[868]) );
  AND U1478 ( .A(n1035), .B(n1477), .Z(n1475) );
  XOR U1479 ( .A(creg[868]), .B(mod_mult_o[868]), .Z(n1477) );
  XNOR U1480 ( .A(n1478), .B(n1479), .Z(o[867]) );
  AND U1481 ( .A(n1035), .B(n1480), .Z(n1478) );
  XOR U1482 ( .A(creg[867]), .B(mod_mult_o[867]), .Z(n1480) );
  XNOR U1483 ( .A(n1481), .B(n1482), .Z(o[866]) );
  AND U1484 ( .A(n1035), .B(n1483), .Z(n1481) );
  XOR U1485 ( .A(creg[866]), .B(mod_mult_o[866]), .Z(n1483) );
  XNOR U1486 ( .A(n1484), .B(n1485), .Z(o[865]) );
  AND U1487 ( .A(n1035), .B(n1486), .Z(n1484) );
  XOR U1488 ( .A(creg[865]), .B(mod_mult_o[865]), .Z(n1486) );
  XNOR U1489 ( .A(n1487), .B(n1488), .Z(o[864]) );
  AND U1490 ( .A(n1035), .B(n1489), .Z(n1487) );
  XOR U1491 ( .A(creg[864]), .B(mod_mult_o[864]), .Z(n1489) );
  XNOR U1492 ( .A(n1490), .B(n1491), .Z(o[863]) );
  AND U1493 ( .A(n1035), .B(n1492), .Z(n1490) );
  XOR U1494 ( .A(creg[863]), .B(mod_mult_o[863]), .Z(n1492) );
  XNOR U1495 ( .A(n1493), .B(n1494), .Z(o[862]) );
  AND U1496 ( .A(n1035), .B(n1495), .Z(n1493) );
  XOR U1497 ( .A(creg[862]), .B(mod_mult_o[862]), .Z(n1495) );
  XNOR U1498 ( .A(n1496), .B(n1497), .Z(o[861]) );
  AND U1499 ( .A(n1035), .B(n1498), .Z(n1496) );
  XOR U1500 ( .A(creg[861]), .B(mod_mult_o[861]), .Z(n1498) );
  XNOR U1501 ( .A(n1499), .B(n1500), .Z(o[860]) );
  AND U1502 ( .A(n1035), .B(n1501), .Z(n1499) );
  XOR U1503 ( .A(creg[860]), .B(mod_mult_o[860]), .Z(n1501) );
  XNOR U1504 ( .A(n1502), .B(n1503), .Z(o[85]) );
  AND U1505 ( .A(n1035), .B(n1504), .Z(n1502) );
  XOR U1506 ( .A(creg[85]), .B(mod_mult_o[85]), .Z(n1504) );
  XNOR U1507 ( .A(n1505), .B(n1506), .Z(o[859]) );
  AND U1508 ( .A(n1035), .B(n1507), .Z(n1505) );
  XOR U1509 ( .A(creg[859]), .B(mod_mult_o[859]), .Z(n1507) );
  XNOR U1510 ( .A(n1508), .B(n1509), .Z(o[858]) );
  AND U1511 ( .A(n1035), .B(n1510), .Z(n1508) );
  XOR U1512 ( .A(creg[858]), .B(mod_mult_o[858]), .Z(n1510) );
  XNOR U1513 ( .A(n1511), .B(n1512), .Z(o[857]) );
  AND U1514 ( .A(n1035), .B(n1513), .Z(n1511) );
  XOR U1515 ( .A(creg[857]), .B(mod_mult_o[857]), .Z(n1513) );
  XNOR U1516 ( .A(n1514), .B(n1515), .Z(o[856]) );
  AND U1517 ( .A(n1035), .B(n1516), .Z(n1514) );
  XOR U1518 ( .A(creg[856]), .B(mod_mult_o[856]), .Z(n1516) );
  XNOR U1519 ( .A(n1517), .B(n1518), .Z(o[855]) );
  AND U1520 ( .A(n1035), .B(n1519), .Z(n1517) );
  XOR U1521 ( .A(creg[855]), .B(mod_mult_o[855]), .Z(n1519) );
  XNOR U1522 ( .A(n1520), .B(n1521), .Z(o[854]) );
  AND U1523 ( .A(n1035), .B(n1522), .Z(n1520) );
  XOR U1524 ( .A(creg[854]), .B(mod_mult_o[854]), .Z(n1522) );
  XNOR U1525 ( .A(n1523), .B(n1524), .Z(o[853]) );
  AND U1526 ( .A(n1035), .B(n1525), .Z(n1523) );
  XOR U1527 ( .A(creg[853]), .B(mod_mult_o[853]), .Z(n1525) );
  XNOR U1528 ( .A(n1526), .B(n1527), .Z(o[852]) );
  AND U1529 ( .A(n1035), .B(n1528), .Z(n1526) );
  XOR U1530 ( .A(creg[852]), .B(mod_mult_o[852]), .Z(n1528) );
  XNOR U1531 ( .A(n1529), .B(n1530), .Z(o[851]) );
  AND U1532 ( .A(n1035), .B(n1531), .Z(n1529) );
  XOR U1533 ( .A(creg[851]), .B(mod_mult_o[851]), .Z(n1531) );
  XNOR U1534 ( .A(n1532), .B(n1533), .Z(o[850]) );
  AND U1535 ( .A(n1035), .B(n1534), .Z(n1532) );
  XOR U1536 ( .A(creg[850]), .B(mod_mult_o[850]), .Z(n1534) );
  XNOR U1537 ( .A(n1535), .B(n1536), .Z(o[84]) );
  AND U1538 ( .A(n1035), .B(n1537), .Z(n1535) );
  XOR U1539 ( .A(creg[84]), .B(mod_mult_o[84]), .Z(n1537) );
  XNOR U1540 ( .A(n1538), .B(n1539), .Z(o[849]) );
  AND U1541 ( .A(n1035), .B(n1540), .Z(n1538) );
  XOR U1542 ( .A(creg[849]), .B(mod_mult_o[849]), .Z(n1540) );
  XNOR U1543 ( .A(n1541), .B(n1542), .Z(o[848]) );
  AND U1544 ( .A(n1035), .B(n1543), .Z(n1541) );
  XOR U1545 ( .A(creg[848]), .B(mod_mult_o[848]), .Z(n1543) );
  XNOR U1546 ( .A(n1544), .B(n1545), .Z(o[847]) );
  AND U1547 ( .A(n1035), .B(n1546), .Z(n1544) );
  XOR U1548 ( .A(creg[847]), .B(mod_mult_o[847]), .Z(n1546) );
  XNOR U1549 ( .A(n1547), .B(n1548), .Z(o[846]) );
  AND U1550 ( .A(n1035), .B(n1549), .Z(n1547) );
  XOR U1551 ( .A(creg[846]), .B(mod_mult_o[846]), .Z(n1549) );
  XNOR U1552 ( .A(n1550), .B(n1551), .Z(o[845]) );
  AND U1553 ( .A(n1035), .B(n1552), .Z(n1550) );
  XOR U1554 ( .A(creg[845]), .B(mod_mult_o[845]), .Z(n1552) );
  XNOR U1555 ( .A(n1553), .B(n1554), .Z(o[844]) );
  AND U1556 ( .A(n1035), .B(n1555), .Z(n1553) );
  XOR U1557 ( .A(creg[844]), .B(mod_mult_o[844]), .Z(n1555) );
  XNOR U1558 ( .A(n1556), .B(n1557), .Z(o[843]) );
  AND U1559 ( .A(n1035), .B(n1558), .Z(n1556) );
  XOR U1560 ( .A(creg[843]), .B(mod_mult_o[843]), .Z(n1558) );
  XNOR U1561 ( .A(n1559), .B(n1560), .Z(o[842]) );
  AND U1562 ( .A(n1035), .B(n1561), .Z(n1559) );
  XOR U1563 ( .A(creg[842]), .B(mod_mult_o[842]), .Z(n1561) );
  XNOR U1564 ( .A(n1562), .B(n1563), .Z(o[841]) );
  AND U1565 ( .A(n1035), .B(n1564), .Z(n1562) );
  XOR U1566 ( .A(creg[841]), .B(mod_mult_o[841]), .Z(n1564) );
  XNOR U1567 ( .A(n1565), .B(n1566), .Z(o[840]) );
  AND U1568 ( .A(n1035), .B(n1567), .Z(n1565) );
  XOR U1569 ( .A(creg[840]), .B(mod_mult_o[840]), .Z(n1567) );
  XNOR U1570 ( .A(n1568), .B(n1569), .Z(o[83]) );
  AND U1571 ( .A(n1035), .B(n1570), .Z(n1568) );
  XOR U1572 ( .A(creg[83]), .B(mod_mult_o[83]), .Z(n1570) );
  XNOR U1573 ( .A(n1571), .B(n1572), .Z(o[839]) );
  AND U1574 ( .A(n1035), .B(n1573), .Z(n1571) );
  XOR U1575 ( .A(creg[839]), .B(mod_mult_o[839]), .Z(n1573) );
  XNOR U1576 ( .A(n1574), .B(n1575), .Z(o[838]) );
  AND U1577 ( .A(n1035), .B(n1576), .Z(n1574) );
  XOR U1578 ( .A(creg[838]), .B(mod_mult_o[838]), .Z(n1576) );
  XNOR U1579 ( .A(n1577), .B(n1578), .Z(o[837]) );
  AND U1580 ( .A(n1035), .B(n1579), .Z(n1577) );
  XOR U1581 ( .A(creg[837]), .B(mod_mult_o[837]), .Z(n1579) );
  XNOR U1582 ( .A(n1580), .B(n1581), .Z(o[836]) );
  AND U1583 ( .A(n1035), .B(n1582), .Z(n1580) );
  XOR U1584 ( .A(creg[836]), .B(mod_mult_o[836]), .Z(n1582) );
  XNOR U1585 ( .A(n1583), .B(n1584), .Z(o[835]) );
  AND U1586 ( .A(n1035), .B(n1585), .Z(n1583) );
  XOR U1587 ( .A(creg[835]), .B(mod_mult_o[835]), .Z(n1585) );
  XNOR U1588 ( .A(n1586), .B(n1587), .Z(o[834]) );
  AND U1589 ( .A(n1035), .B(n1588), .Z(n1586) );
  XOR U1590 ( .A(creg[834]), .B(mod_mult_o[834]), .Z(n1588) );
  XNOR U1591 ( .A(n1589), .B(n1590), .Z(o[833]) );
  AND U1592 ( .A(n1035), .B(n1591), .Z(n1589) );
  XOR U1593 ( .A(creg[833]), .B(mod_mult_o[833]), .Z(n1591) );
  XNOR U1594 ( .A(n1592), .B(n1593), .Z(o[832]) );
  AND U1595 ( .A(n1035), .B(n1594), .Z(n1592) );
  XOR U1596 ( .A(creg[832]), .B(mod_mult_o[832]), .Z(n1594) );
  XNOR U1597 ( .A(n1595), .B(n1596), .Z(o[831]) );
  AND U1598 ( .A(n1035), .B(n1597), .Z(n1595) );
  XOR U1599 ( .A(creg[831]), .B(mod_mult_o[831]), .Z(n1597) );
  XNOR U1600 ( .A(n1598), .B(n1599), .Z(o[830]) );
  AND U1601 ( .A(n1035), .B(n1600), .Z(n1598) );
  XOR U1602 ( .A(creg[830]), .B(mod_mult_o[830]), .Z(n1600) );
  XNOR U1603 ( .A(n1601), .B(n1602), .Z(o[82]) );
  AND U1604 ( .A(n1035), .B(n1603), .Z(n1601) );
  XOR U1605 ( .A(creg[82]), .B(mod_mult_o[82]), .Z(n1603) );
  XNOR U1606 ( .A(n1604), .B(n1605), .Z(o[829]) );
  AND U1607 ( .A(n1035), .B(n1606), .Z(n1604) );
  XOR U1608 ( .A(creg[829]), .B(mod_mult_o[829]), .Z(n1606) );
  XNOR U1609 ( .A(n1607), .B(n1608), .Z(o[828]) );
  AND U1610 ( .A(n1035), .B(n1609), .Z(n1607) );
  XOR U1611 ( .A(creg[828]), .B(mod_mult_o[828]), .Z(n1609) );
  XNOR U1612 ( .A(n1610), .B(n1611), .Z(o[827]) );
  AND U1613 ( .A(n1035), .B(n1612), .Z(n1610) );
  XOR U1614 ( .A(creg[827]), .B(mod_mult_o[827]), .Z(n1612) );
  XNOR U1615 ( .A(n1613), .B(n1614), .Z(o[826]) );
  AND U1616 ( .A(n1035), .B(n1615), .Z(n1613) );
  XOR U1617 ( .A(creg[826]), .B(mod_mult_o[826]), .Z(n1615) );
  XNOR U1618 ( .A(n1616), .B(n1617), .Z(o[825]) );
  AND U1619 ( .A(n1035), .B(n1618), .Z(n1616) );
  XOR U1620 ( .A(creg[825]), .B(mod_mult_o[825]), .Z(n1618) );
  XNOR U1621 ( .A(n1619), .B(n1620), .Z(o[824]) );
  AND U1622 ( .A(n1035), .B(n1621), .Z(n1619) );
  XOR U1623 ( .A(creg[824]), .B(mod_mult_o[824]), .Z(n1621) );
  XNOR U1624 ( .A(n1622), .B(n1623), .Z(o[823]) );
  AND U1625 ( .A(n1035), .B(n1624), .Z(n1622) );
  XOR U1626 ( .A(creg[823]), .B(mod_mult_o[823]), .Z(n1624) );
  XNOR U1627 ( .A(n1625), .B(n1626), .Z(o[822]) );
  AND U1628 ( .A(n1035), .B(n1627), .Z(n1625) );
  XOR U1629 ( .A(creg[822]), .B(mod_mult_o[822]), .Z(n1627) );
  XNOR U1630 ( .A(n1628), .B(n1629), .Z(o[821]) );
  AND U1631 ( .A(n1035), .B(n1630), .Z(n1628) );
  XOR U1632 ( .A(creg[821]), .B(mod_mult_o[821]), .Z(n1630) );
  XNOR U1633 ( .A(n1631), .B(n1632), .Z(o[820]) );
  AND U1634 ( .A(n1035), .B(n1633), .Z(n1631) );
  XOR U1635 ( .A(creg[820]), .B(mod_mult_o[820]), .Z(n1633) );
  XNOR U1636 ( .A(n1634), .B(n1635), .Z(o[81]) );
  AND U1637 ( .A(n1035), .B(n1636), .Z(n1634) );
  XOR U1638 ( .A(creg[81]), .B(mod_mult_o[81]), .Z(n1636) );
  XNOR U1639 ( .A(n1637), .B(n1638), .Z(o[819]) );
  AND U1640 ( .A(n1035), .B(n1639), .Z(n1637) );
  XOR U1641 ( .A(creg[819]), .B(mod_mult_o[819]), .Z(n1639) );
  XNOR U1642 ( .A(n1640), .B(n1641), .Z(o[818]) );
  AND U1643 ( .A(n1035), .B(n1642), .Z(n1640) );
  XOR U1644 ( .A(creg[818]), .B(mod_mult_o[818]), .Z(n1642) );
  XNOR U1645 ( .A(n1643), .B(n1644), .Z(o[817]) );
  AND U1646 ( .A(n1035), .B(n1645), .Z(n1643) );
  XOR U1647 ( .A(creg[817]), .B(mod_mult_o[817]), .Z(n1645) );
  XNOR U1648 ( .A(n1646), .B(n1647), .Z(o[816]) );
  AND U1649 ( .A(n1035), .B(n1648), .Z(n1646) );
  XOR U1650 ( .A(creg[816]), .B(mod_mult_o[816]), .Z(n1648) );
  XNOR U1651 ( .A(n1649), .B(n1650), .Z(o[815]) );
  AND U1652 ( .A(n1035), .B(n1651), .Z(n1649) );
  XOR U1653 ( .A(creg[815]), .B(mod_mult_o[815]), .Z(n1651) );
  XNOR U1654 ( .A(n1652), .B(n1653), .Z(o[814]) );
  AND U1655 ( .A(n1035), .B(n1654), .Z(n1652) );
  XOR U1656 ( .A(creg[814]), .B(mod_mult_o[814]), .Z(n1654) );
  XNOR U1657 ( .A(n1655), .B(n1656), .Z(o[813]) );
  AND U1658 ( .A(n1035), .B(n1657), .Z(n1655) );
  XOR U1659 ( .A(creg[813]), .B(mod_mult_o[813]), .Z(n1657) );
  XNOR U1660 ( .A(n1658), .B(n1659), .Z(o[812]) );
  AND U1661 ( .A(n1035), .B(n1660), .Z(n1658) );
  XOR U1662 ( .A(creg[812]), .B(mod_mult_o[812]), .Z(n1660) );
  XNOR U1663 ( .A(n1661), .B(n1662), .Z(o[811]) );
  AND U1664 ( .A(n1035), .B(n1663), .Z(n1661) );
  XOR U1665 ( .A(creg[811]), .B(mod_mult_o[811]), .Z(n1663) );
  XNOR U1666 ( .A(n1664), .B(n1665), .Z(o[810]) );
  AND U1667 ( .A(n1035), .B(n1666), .Z(n1664) );
  XOR U1668 ( .A(creg[810]), .B(mod_mult_o[810]), .Z(n1666) );
  XNOR U1669 ( .A(n1667), .B(n1668), .Z(o[80]) );
  AND U1670 ( .A(n1035), .B(n1669), .Z(n1667) );
  XOR U1671 ( .A(creg[80]), .B(mod_mult_o[80]), .Z(n1669) );
  XNOR U1672 ( .A(n1670), .B(n1671), .Z(o[809]) );
  AND U1673 ( .A(n1035), .B(n1672), .Z(n1670) );
  XOR U1674 ( .A(creg[809]), .B(mod_mult_o[809]), .Z(n1672) );
  XNOR U1675 ( .A(n1673), .B(n1674), .Z(o[808]) );
  AND U1676 ( .A(n1035), .B(n1675), .Z(n1673) );
  XOR U1677 ( .A(creg[808]), .B(mod_mult_o[808]), .Z(n1675) );
  XNOR U1678 ( .A(n1676), .B(n1677), .Z(o[807]) );
  AND U1679 ( .A(n1035), .B(n1678), .Z(n1676) );
  XOR U1680 ( .A(creg[807]), .B(mod_mult_o[807]), .Z(n1678) );
  XNOR U1681 ( .A(n1679), .B(n1680), .Z(o[806]) );
  AND U1682 ( .A(n1035), .B(n1681), .Z(n1679) );
  XOR U1683 ( .A(creg[806]), .B(mod_mult_o[806]), .Z(n1681) );
  XNOR U1684 ( .A(n1682), .B(n1683), .Z(o[805]) );
  AND U1685 ( .A(n1035), .B(n1684), .Z(n1682) );
  XOR U1686 ( .A(creg[805]), .B(mod_mult_o[805]), .Z(n1684) );
  XNOR U1687 ( .A(n1685), .B(n1686), .Z(o[804]) );
  AND U1688 ( .A(n1035), .B(n1687), .Z(n1685) );
  XOR U1689 ( .A(creg[804]), .B(mod_mult_o[804]), .Z(n1687) );
  XNOR U1690 ( .A(n1688), .B(n1689), .Z(o[803]) );
  AND U1691 ( .A(n1035), .B(n1690), .Z(n1688) );
  XOR U1692 ( .A(creg[803]), .B(mod_mult_o[803]), .Z(n1690) );
  XNOR U1693 ( .A(n1691), .B(n1692), .Z(o[802]) );
  AND U1694 ( .A(n1035), .B(n1693), .Z(n1691) );
  XOR U1695 ( .A(creg[802]), .B(mod_mult_o[802]), .Z(n1693) );
  XNOR U1696 ( .A(n1694), .B(n1695), .Z(o[801]) );
  AND U1697 ( .A(n1035), .B(n1696), .Z(n1694) );
  XOR U1698 ( .A(creg[801]), .B(mod_mult_o[801]), .Z(n1696) );
  XNOR U1699 ( .A(n1697), .B(n1698), .Z(o[800]) );
  AND U1700 ( .A(n1035), .B(n1699), .Z(n1697) );
  XOR U1701 ( .A(creg[800]), .B(mod_mult_o[800]), .Z(n1699) );
  XNOR U1702 ( .A(n1700), .B(n1701), .Z(o[7]) );
  AND U1703 ( .A(n1035), .B(n1702), .Z(n1700) );
  XOR U1704 ( .A(creg[7]), .B(mod_mult_o[7]), .Z(n1702) );
  XNOR U1705 ( .A(n1703), .B(n1704), .Z(o[79]) );
  AND U1706 ( .A(n1035), .B(n1705), .Z(n1703) );
  XOR U1707 ( .A(creg[79]), .B(mod_mult_o[79]), .Z(n1705) );
  XNOR U1708 ( .A(n1706), .B(n1707), .Z(o[799]) );
  AND U1709 ( .A(n1035), .B(n1708), .Z(n1706) );
  XOR U1710 ( .A(creg[799]), .B(mod_mult_o[799]), .Z(n1708) );
  XNOR U1711 ( .A(n1709), .B(n1710), .Z(o[798]) );
  AND U1712 ( .A(n1035), .B(n1711), .Z(n1709) );
  XOR U1713 ( .A(creg[798]), .B(mod_mult_o[798]), .Z(n1711) );
  XNOR U1714 ( .A(n1712), .B(n1713), .Z(o[797]) );
  AND U1715 ( .A(n1035), .B(n1714), .Z(n1712) );
  XOR U1716 ( .A(creg[797]), .B(mod_mult_o[797]), .Z(n1714) );
  XNOR U1717 ( .A(n1715), .B(n1716), .Z(o[796]) );
  AND U1718 ( .A(n1035), .B(n1717), .Z(n1715) );
  XOR U1719 ( .A(creg[796]), .B(mod_mult_o[796]), .Z(n1717) );
  XNOR U1720 ( .A(n1718), .B(n1719), .Z(o[795]) );
  AND U1721 ( .A(n1035), .B(n1720), .Z(n1718) );
  XOR U1722 ( .A(creg[795]), .B(mod_mult_o[795]), .Z(n1720) );
  XNOR U1723 ( .A(n1721), .B(n1722), .Z(o[794]) );
  AND U1724 ( .A(n1035), .B(n1723), .Z(n1721) );
  XOR U1725 ( .A(creg[794]), .B(mod_mult_o[794]), .Z(n1723) );
  XNOR U1726 ( .A(n1724), .B(n1725), .Z(o[793]) );
  AND U1727 ( .A(n1035), .B(n1726), .Z(n1724) );
  XOR U1728 ( .A(creg[793]), .B(mod_mult_o[793]), .Z(n1726) );
  XNOR U1729 ( .A(n1727), .B(n1728), .Z(o[792]) );
  AND U1730 ( .A(n1035), .B(n1729), .Z(n1727) );
  XOR U1731 ( .A(creg[792]), .B(mod_mult_o[792]), .Z(n1729) );
  XNOR U1732 ( .A(n1730), .B(n1731), .Z(o[791]) );
  AND U1733 ( .A(n1035), .B(n1732), .Z(n1730) );
  XOR U1734 ( .A(creg[791]), .B(mod_mult_o[791]), .Z(n1732) );
  XNOR U1735 ( .A(n1733), .B(n1734), .Z(o[790]) );
  AND U1736 ( .A(n1035), .B(n1735), .Z(n1733) );
  XOR U1737 ( .A(creg[790]), .B(mod_mult_o[790]), .Z(n1735) );
  XNOR U1738 ( .A(n1736), .B(n1737), .Z(o[78]) );
  AND U1739 ( .A(n1035), .B(n1738), .Z(n1736) );
  XOR U1740 ( .A(creg[78]), .B(mod_mult_o[78]), .Z(n1738) );
  XNOR U1741 ( .A(n1739), .B(n1740), .Z(o[789]) );
  AND U1742 ( .A(n1035), .B(n1741), .Z(n1739) );
  XOR U1743 ( .A(creg[789]), .B(mod_mult_o[789]), .Z(n1741) );
  XNOR U1744 ( .A(n1742), .B(n1743), .Z(o[788]) );
  AND U1745 ( .A(n1035), .B(n1744), .Z(n1742) );
  XOR U1746 ( .A(creg[788]), .B(mod_mult_o[788]), .Z(n1744) );
  XNOR U1747 ( .A(n1745), .B(n1746), .Z(o[787]) );
  AND U1748 ( .A(n1035), .B(n1747), .Z(n1745) );
  XOR U1749 ( .A(creg[787]), .B(mod_mult_o[787]), .Z(n1747) );
  XNOR U1750 ( .A(n1748), .B(n1749), .Z(o[786]) );
  AND U1751 ( .A(n1035), .B(n1750), .Z(n1748) );
  XOR U1752 ( .A(creg[786]), .B(mod_mult_o[786]), .Z(n1750) );
  XNOR U1753 ( .A(n1751), .B(n1752), .Z(o[785]) );
  AND U1754 ( .A(n1035), .B(n1753), .Z(n1751) );
  XOR U1755 ( .A(creg[785]), .B(mod_mult_o[785]), .Z(n1753) );
  XNOR U1756 ( .A(n1754), .B(n1755), .Z(o[784]) );
  AND U1757 ( .A(n1035), .B(n1756), .Z(n1754) );
  XOR U1758 ( .A(creg[784]), .B(mod_mult_o[784]), .Z(n1756) );
  XNOR U1759 ( .A(n1757), .B(n1758), .Z(o[783]) );
  AND U1760 ( .A(n1035), .B(n1759), .Z(n1757) );
  XOR U1761 ( .A(creg[783]), .B(mod_mult_o[783]), .Z(n1759) );
  XNOR U1762 ( .A(n1760), .B(n1761), .Z(o[782]) );
  AND U1763 ( .A(n1035), .B(n1762), .Z(n1760) );
  XOR U1764 ( .A(creg[782]), .B(mod_mult_o[782]), .Z(n1762) );
  XNOR U1765 ( .A(n1763), .B(n1764), .Z(o[781]) );
  AND U1766 ( .A(n1035), .B(n1765), .Z(n1763) );
  XOR U1767 ( .A(creg[781]), .B(mod_mult_o[781]), .Z(n1765) );
  XNOR U1768 ( .A(n1766), .B(n1767), .Z(o[780]) );
  AND U1769 ( .A(n1035), .B(n1768), .Z(n1766) );
  XOR U1770 ( .A(creg[780]), .B(mod_mult_o[780]), .Z(n1768) );
  XNOR U1771 ( .A(n1769), .B(n1770), .Z(o[77]) );
  AND U1772 ( .A(n1035), .B(n1771), .Z(n1769) );
  XOR U1773 ( .A(creg[77]), .B(mod_mult_o[77]), .Z(n1771) );
  XNOR U1774 ( .A(n1772), .B(n1773), .Z(o[779]) );
  AND U1775 ( .A(n1035), .B(n1774), .Z(n1772) );
  XOR U1776 ( .A(creg[779]), .B(mod_mult_o[779]), .Z(n1774) );
  XNOR U1777 ( .A(n1775), .B(n1776), .Z(o[778]) );
  AND U1778 ( .A(n1035), .B(n1777), .Z(n1775) );
  XOR U1779 ( .A(creg[778]), .B(mod_mult_o[778]), .Z(n1777) );
  XNOR U1780 ( .A(n1778), .B(n1779), .Z(o[777]) );
  AND U1781 ( .A(n1035), .B(n1780), .Z(n1778) );
  XOR U1782 ( .A(creg[777]), .B(mod_mult_o[777]), .Z(n1780) );
  XNOR U1783 ( .A(n1781), .B(n1782), .Z(o[776]) );
  AND U1784 ( .A(n1035), .B(n1783), .Z(n1781) );
  XOR U1785 ( .A(creg[776]), .B(mod_mult_o[776]), .Z(n1783) );
  XNOR U1786 ( .A(n1784), .B(n1785), .Z(o[775]) );
  AND U1787 ( .A(n1035), .B(n1786), .Z(n1784) );
  XOR U1788 ( .A(creg[775]), .B(mod_mult_o[775]), .Z(n1786) );
  XNOR U1789 ( .A(n1787), .B(n1788), .Z(o[774]) );
  AND U1790 ( .A(n1035), .B(n1789), .Z(n1787) );
  XOR U1791 ( .A(creg[774]), .B(mod_mult_o[774]), .Z(n1789) );
  XNOR U1792 ( .A(n1790), .B(n1791), .Z(o[773]) );
  AND U1793 ( .A(n1035), .B(n1792), .Z(n1790) );
  XOR U1794 ( .A(creg[773]), .B(mod_mult_o[773]), .Z(n1792) );
  XNOR U1795 ( .A(n1793), .B(n1794), .Z(o[772]) );
  AND U1796 ( .A(n1035), .B(n1795), .Z(n1793) );
  XOR U1797 ( .A(creg[772]), .B(mod_mult_o[772]), .Z(n1795) );
  XNOR U1798 ( .A(n1796), .B(n1797), .Z(o[771]) );
  AND U1799 ( .A(n1035), .B(n1798), .Z(n1796) );
  XOR U1800 ( .A(creg[771]), .B(mod_mult_o[771]), .Z(n1798) );
  XNOR U1801 ( .A(n1799), .B(n1800), .Z(o[770]) );
  AND U1802 ( .A(n1035), .B(n1801), .Z(n1799) );
  XOR U1803 ( .A(creg[770]), .B(mod_mult_o[770]), .Z(n1801) );
  XNOR U1804 ( .A(n1802), .B(n1803), .Z(o[76]) );
  AND U1805 ( .A(n1035), .B(n1804), .Z(n1802) );
  XOR U1806 ( .A(creg[76]), .B(mod_mult_o[76]), .Z(n1804) );
  XNOR U1807 ( .A(n1805), .B(n1806), .Z(o[769]) );
  AND U1808 ( .A(n1035), .B(n1807), .Z(n1805) );
  XOR U1809 ( .A(creg[769]), .B(mod_mult_o[769]), .Z(n1807) );
  XNOR U1810 ( .A(n1808), .B(n1809), .Z(o[768]) );
  AND U1811 ( .A(n1035), .B(n1810), .Z(n1808) );
  XOR U1812 ( .A(creg[768]), .B(mod_mult_o[768]), .Z(n1810) );
  XNOR U1813 ( .A(n1811), .B(n1812), .Z(o[767]) );
  AND U1814 ( .A(n1035), .B(n1813), .Z(n1811) );
  XOR U1815 ( .A(creg[767]), .B(mod_mult_o[767]), .Z(n1813) );
  XNOR U1816 ( .A(n1814), .B(n1815), .Z(o[766]) );
  AND U1817 ( .A(n1035), .B(n1816), .Z(n1814) );
  XOR U1818 ( .A(creg[766]), .B(mod_mult_o[766]), .Z(n1816) );
  XNOR U1819 ( .A(n1817), .B(n1818), .Z(o[765]) );
  AND U1820 ( .A(n1035), .B(n1819), .Z(n1817) );
  XOR U1821 ( .A(creg[765]), .B(mod_mult_o[765]), .Z(n1819) );
  XNOR U1822 ( .A(n1820), .B(n1821), .Z(o[764]) );
  AND U1823 ( .A(n1035), .B(n1822), .Z(n1820) );
  XOR U1824 ( .A(creg[764]), .B(mod_mult_o[764]), .Z(n1822) );
  XNOR U1825 ( .A(n1823), .B(n1824), .Z(o[763]) );
  AND U1826 ( .A(n1035), .B(n1825), .Z(n1823) );
  XOR U1827 ( .A(creg[763]), .B(mod_mult_o[763]), .Z(n1825) );
  XNOR U1828 ( .A(n1826), .B(n1827), .Z(o[762]) );
  AND U1829 ( .A(n1035), .B(n1828), .Z(n1826) );
  XOR U1830 ( .A(creg[762]), .B(mod_mult_o[762]), .Z(n1828) );
  XNOR U1831 ( .A(n1829), .B(n1830), .Z(o[761]) );
  AND U1832 ( .A(n1035), .B(n1831), .Z(n1829) );
  XOR U1833 ( .A(creg[761]), .B(mod_mult_o[761]), .Z(n1831) );
  XNOR U1834 ( .A(n1832), .B(n1833), .Z(o[760]) );
  AND U1835 ( .A(n1035), .B(n1834), .Z(n1832) );
  XOR U1836 ( .A(creg[760]), .B(mod_mult_o[760]), .Z(n1834) );
  XNOR U1837 ( .A(n1835), .B(n1836), .Z(o[75]) );
  AND U1838 ( .A(n1035), .B(n1837), .Z(n1835) );
  XOR U1839 ( .A(creg[75]), .B(mod_mult_o[75]), .Z(n1837) );
  XNOR U1840 ( .A(n1838), .B(n1839), .Z(o[759]) );
  AND U1841 ( .A(n1035), .B(n1840), .Z(n1838) );
  XOR U1842 ( .A(creg[759]), .B(mod_mult_o[759]), .Z(n1840) );
  XNOR U1843 ( .A(n1841), .B(n1842), .Z(o[758]) );
  AND U1844 ( .A(n1035), .B(n1843), .Z(n1841) );
  XOR U1845 ( .A(creg[758]), .B(mod_mult_o[758]), .Z(n1843) );
  XNOR U1846 ( .A(n1844), .B(n1845), .Z(o[757]) );
  AND U1847 ( .A(n1035), .B(n1846), .Z(n1844) );
  XOR U1848 ( .A(creg[757]), .B(mod_mult_o[757]), .Z(n1846) );
  XNOR U1849 ( .A(n1847), .B(n1848), .Z(o[756]) );
  AND U1850 ( .A(n1035), .B(n1849), .Z(n1847) );
  XOR U1851 ( .A(creg[756]), .B(mod_mult_o[756]), .Z(n1849) );
  XNOR U1852 ( .A(n1850), .B(n1851), .Z(o[755]) );
  AND U1853 ( .A(n1035), .B(n1852), .Z(n1850) );
  XOR U1854 ( .A(creg[755]), .B(mod_mult_o[755]), .Z(n1852) );
  XNOR U1855 ( .A(n1853), .B(n1854), .Z(o[754]) );
  AND U1856 ( .A(n1035), .B(n1855), .Z(n1853) );
  XOR U1857 ( .A(creg[754]), .B(mod_mult_o[754]), .Z(n1855) );
  XNOR U1858 ( .A(n1856), .B(n1857), .Z(o[753]) );
  AND U1859 ( .A(n1035), .B(n1858), .Z(n1856) );
  XOR U1860 ( .A(creg[753]), .B(mod_mult_o[753]), .Z(n1858) );
  XNOR U1861 ( .A(n1859), .B(n1860), .Z(o[752]) );
  AND U1862 ( .A(n1035), .B(n1861), .Z(n1859) );
  XOR U1863 ( .A(creg[752]), .B(mod_mult_o[752]), .Z(n1861) );
  XNOR U1864 ( .A(n1862), .B(n1863), .Z(o[751]) );
  AND U1865 ( .A(n1035), .B(n1864), .Z(n1862) );
  XOR U1866 ( .A(creg[751]), .B(mod_mult_o[751]), .Z(n1864) );
  XNOR U1867 ( .A(n1865), .B(n1866), .Z(o[750]) );
  AND U1868 ( .A(n1035), .B(n1867), .Z(n1865) );
  XOR U1869 ( .A(creg[750]), .B(mod_mult_o[750]), .Z(n1867) );
  XNOR U1870 ( .A(n1868), .B(n1869), .Z(o[74]) );
  AND U1871 ( .A(n1035), .B(n1870), .Z(n1868) );
  XOR U1872 ( .A(creg[74]), .B(mod_mult_o[74]), .Z(n1870) );
  XNOR U1873 ( .A(n1871), .B(n1872), .Z(o[749]) );
  AND U1874 ( .A(n1035), .B(n1873), .Z(n1871) );
  XOR U1875 ( .A(creg[749]), .B(mod_mult_o[749]), .Z(n1873) );
  XNOR U1876 ( .A(n1874), .B(n1875), .Z(o[748]) );
  AND U1877 ( .A(n1035), .B(n1876), .Z(n1874) );
  XOR U1878 ( .A(creg[748]), .B(mod_mult_o[748]), .Z(n1876) );
  XNOR U1879 ( .A(n1877), .B(n1878), .Z(o[747]) );
  AND U1880 ( .A(n1035), .B(n1879), .Z(n1877) );
  XOR U1881 ( .A(creg[747]), .B(mod_mult_o[747]), .Z(n1879) );
  XNOR U1882 ( .A(n1880), .B(n1881), .Z(o[746]) );
  AND U1883 ( .A(n1035), .B(n1882), .Z(n1880) );
  XOR U1884 ( .A(creg[746]), .B(mod_mult_o[746]), .Z(n1882) );
  XNOR U1885 ( .A(n1883), .B(n1884), .Z(o[745]) );
  AND U1886 ( .A(n1035), .B(n1885), .Z(n1883) );
  XOR U1887 ( .A(creg[745]), .B(mod_mult_o[745]), .Z(n1885) );
  XNOR U1888 ( .A(n1886), .B(n1887), .Z(o[744]) );
  AND U1889 ( .A(n1035), .B(n1888), .Z(n1886) );
  XOR U1890 ( .A(creg[744]), .B(mod_mult_o[744]), .Z(n1888) );
  XNOR U1891 ( .A(n1889), .B(n1890), .Z(o[743]) );
  AND U1892 ( .A(n1035), .B(n1891), .Z(n1889) );
  XOR U1893 ( .A(creg[743]), .B(mod_mult_o[743]), .Z(n1891) );
  XNOR U1894 ( .A(n1892), .B(n1893), .Z(o[742]) );
  AND U1895 ( .A(n1035), .B(n1894), .Z(n1892) );
  XOR U1896 ( .A(creg[742]), .B(mod_mult_o[742]), .Z(n1894) );
  XNOR U1897 ( .A(n1895), .B(n1896), .Z(o[741]) );
  AND U1898 ( .A(n1035), .B(n1897), .Z(n1895) );
  XOR U1899 ( .A(creg[741]), .B(mod_mult_o[741]), .Z(n1897) );
  XNOR U1900 ( .A(n1898), .B(n1899), .Z(o[740]) );
  AND U1901 ( .A(n1035), .B(n1900), .Z(n1898) );
  XOR U1902 ( .A(creg[740]), .B(mod_mult_o[740]), .Z(n1900) );
  XNOR U1903 ( .A(n1901), .B(n1902), .Z(o[73]) );
  AND U1904 ( .A(n1035), .B(n1903), .Z(n1901) );
  XOR U1905 ( .A(creg[73]), .B(mod_mult_o[73]), .Z(n1903) );
  XNOR U1906 ( .A(n1904), .B(n1905), .Z(o[739]) );
  AND U1907 ( .A(n1035), .B(n1906), .Z(n1904) );
  XOR U1908 ( .A(creg[739]), .B(mod_mult_o[739]), .Z(n1906) );
  XNOR U1909 ( .A(n1907), .B(n1908), .Z(o[738]) );
  AND U1910 ( .A(n1035), .B(n1909), .Z(n1907) );
  XOR U1911 ( .A(creg[738]), .B(mod_mult_o[738]), .Z(n1909) );
  XNOR U1912 ( .A(n1910), .B(n1911), .Z(o[737]) );
  AND U1913 ( .A(n1035), .B(n1912), .Z(n1910) );
  XOR U1914 ( .A(creg[737]), .B(mod_mult_o[737]), .Z(n1912) );
  XNOR U1915 ( .A(n1913), .B(n1914), .Z(o[736]) );
  AND U1916 ( .A(n1035), .B(n1915), .Z(n1913) );
  XOR U1917 ( .A(creg[736]), .B(mod_mult_o[736]), .Z(n1915) );
  XNOR U1918 ( .A(n1916), .B(n1917), .Z(o[735]) );
  AND U1919 ( .A(n1035), .B(n1918), .Z(n1916) );
  XOR U1920 ( .A(creg[735]), .B(mod_mult_o[735]), .Z(n1918) );
  XNOR U1921 ( .A(n1919), .B(n1920), .Z(o[734]) );
  AND U1922 ( .A(n1035), .B(n1921), .Z(n1919) );
  XOR U1923 ( .A(creg[734]), .B(mod_mult_o[734]), .Z(n1921) );
  XNOR U1924 ( .A(n1922), .B(n1923), .Z(o[733]) );
  AND U1925 ( .A(n1035), .B(n1924), .Z(n1922) );
  XOR U1926 ( .A(creg[733]), .B(mod_mult_o[733]), .Z(n1924) );
  XNOR U1927 ( .A(n1925), .B(n1926), .Z(o[732]) );
  AND U1928 ( .A(n1035), .B(n1927), .Z(n1925) );
  XOR U1929 ( .A(creg[732]), .B(mod_mult_o[732]), .Z(n1927) );
  XNOR U1930 ( .A(n1928), .B(n1929), .Z(o[731]) );
  AND U1931 ( .A(n1035), .B(n1930), .Z(n1928) );
  XOR U1932 ( .A(creg[731]), .B(mod_mult_o[731]), .Z(n1930) );
  XNOR U1933 ( .A(n1931), .B(n1932), .Z(o[730]) );
  AND U1934 ( .A(n1035), .B(n1933), .Z(n1931) );
  XOR U1935 ( .A(creg[730]), .B(mod_mult_o[730]), .Z(n1933) );
  XNOR U1936 ( .A(n1934), .B(n1935), .Z(o[72]) );
  AND U1937 ( .A(n1035), .B(n1936), .Z(n1934) );
  XOR U1938 ( .A(creg[72]), .B(mod_mult_o[72]), .Z(n1936) );
  XNOR U1939 ( .A(n1937), .B(n1938), .Z(o[729]) );
  AND U1940 ( .A(n1035), .B(n1939), .Z(n1937) );
  XOR U1941 ( .A(creg[729]), .B(mod_mult_o[729]), .Z(n1939) );
  XNOR U1942 ( .A(n1940), .B(n1941), .Z(o[728]) );
  AND U1943 ( .A(n1035), .B(n1942), .Z(n1940) );
  XOR U1944 ( .A(creg[728]), .B(mod_mult_o[728]), .Z(n1942) );
  XNOR U1945 ( .A(n1943), .B(n1944), .Z(o[727]) );
  AND U1946 ( .A(n1035), .B(n1945), .Z(n1943) );
  XOR U1947 ( .A(creg[727]), .B(mod_mult_o[727]), .Z(n1945) );
  XNOR U1948 ( .A(n1946), .B(n1947), .Z(o[726]) );
  AND U1949 ( .A(n1035), .B(n1948), .Z(n1946) );
  XOR U1950 ( .A(creg[726]), .B(mod_mult_o[726]), .Z(n1948) );
  XNOR U1951 ( .A(n1949), .B(n1950), .Z(o[725]) );
  AND U1952 ( .A(n1035), .B(n1951), .Z(n1949) );
  XOR U1953 ( .A(creg[725]), .B(mod_mult_o[725]), .Z(n1951) );
  XNOR U1954 ( .A(n1952), .B(n1953), .Z(o[724]) );
  AND U1955 ( .A(n1035), .B(n1954), .Z(n1952) );
  XOR U1956 ( .A(creg[724]), .B(mod_mult_o[724]), .Z(n1954) );
  XNOR U1957 ( .A(n1955), .B(n1956), .Z(o[723]) );
  AND U1958 ( .A(n1035), .B(n1957), .Z(n1955) );
  XOR U1959 ( .A(creg[723]), .B(mod_mult_o[723]), .Z(n1957) );
  XNOR U1960 ( .A(n1958), .B(n1959), .Z(o[722]) );
  AND U1961 ( .A(n1035), .B(n1960), .Z(n1958) );
  XOR U1962 ( .A(creg[722]), .B(mod_mult_o[722]), .Z(n1960) );
  XNOR U1963 ( .A(n1961), .B(n1962), .Z(o[721]) );
  AND U1964 ( .A(n1035), .B(n1963), .Z(n1961) );
  XOR U1965 ( .A(creg[721]), .B(mod_mult_o[721]), .Z(n1963) );
  XNOR U1966 ( .A(n1964), .B(n1965), .Z(o[720]) );
  AND U1967 ( .A(n1035), .B(n1966), .Z(n1964) );
  XOR U1968 ( .A(creg[720]), .B(mod_mult_o[720]), .Z(n1966) );
  XNOR U1969 ( .A(n1967), .B(n1968), .Z(o[71]) );
  AND U1970 ( .A(n1035), .B(n1969), .Z(n1967) );
  XOR U1971 ( .A(creg[71]), .B(mod_mult_o[71]), .Z(n1969) );
  XNOR U1972 ( .A(n1970), .B(n1971), .Z(o[719]) );
  AND U1973 ( .A(n1035), .B(n1972), .Z(n1970) );
  XOR U1974 ( .A(creg[719]), .B(mod_mult_o[719]), .Z(n1972) );
  XNOR U1975 ( .A(n1973), .B(n1974), .Z(o[718]) );
  AND U1976 ( .A(n1035), .B(n1975), .Z(n1973) );
  XOR U1977 ( .A(creg[718]), .B(mod_mult_o[718]), .Z(n1975) );
  XNOR U1978 ( .A(n1976), .B(n1977), .Z(o[717]) );
  AND U1979 ( .A(n1035), .B(n1978), .Z(n1976) );
  XOR U1980 ( .A(creg[717]), .B(mod_mult_o[717]), .Z(n1978) );
  XNOR U1981 ( .A(n1979), .B(n1980), .Z(o[716]) );
  AND U1982 ( .A(n1035), .B(n1981), .Z(n1979) );
  XOR U1983 ( .A(creg[716]), .B(mod_mult_o[716]), .Z(n1981) );
  XNOR U1984 ( .A(n1982), .B(n1983), .Z(o[715]) );
  AND U1985 ( .A(n1035), .B(n1984), .Z(n1982) );
  XOR U1986 ( .A(creg[715]), .B(mod_mult_o[715]), .Z(n1984) );
  XNOR U1987 ( .A(n1985), .B(n1986), .Z(o[714]) );
  AND U1988 ( .A(n1035), .B(n1987), .Z(n1985) );
  XOR U1989 ( .A(creg[714]), .B(mod_mult_o[714]), .Z(n1987) );
  XNOR U1990 ( .A(n1988), .B(n1989), .Z(o[713]) );
  AND U1991 ( .A(n1035), .B(n1990), .Z(n1988) );
  XOR U1992 ( .A(creg[713]), .B(mod_mult_o[713]), .Z(n1990) );
  XNOR U1993 ( .A(n1991), .B(n1992), .Z(o[712]) );
  AND U1994 ( .A(n1035), .B(n1993), .Z(n1991) );
  XOR U1995 ( .A(creg[712]), .B(mod_mult_o[712]), .Z(n1993) );
  XNOR U1996 ( .A(n1994), .B(n1995), .Z(o[711]) );
  AND U1997 ( .A(n1035), .B(n1996), .Z(n1994) );
  XOR U1998 ( .A(creg[711]), .B(mod_mult_o[711]), .Z(n1996) );
  XNOR U1999 ( .A(n1997), .B(n1998), .Z(o[710]) );
  AND U2000 ( .A(n1035), .B(n1999), .Z(n1997) );
  XOR U2001 ( .A(creg[710]), .B(mod_mult_o[710]), .Z(n1999) );
  XNOR U2002 ( .A(n2000), .B(n2001), .Z(o[70]) );
  AND U2003 ( .A(n1035), .B(n2002), .Z(n2000) );
  XOR U2004 ( .A(creg[70]), .B(mod_mult_o[70]), .Z(n2002) );
  XNOR U2005 ( .A(n2003), .B(n2004), .Z(o[709]) );
  AND U2006 ( .A(n1035), .B(n2005), .Z(n2003) );
  XOR U2007 ( .A(creg[709]), .B(mod_mult_o[709]), .Z(n2005) );
  XNOR U2008 ( .A(n2006), .B(n2007), .Z(o[708]) );
  AND U2009 ( .A(n1035), .B(n2008), .Z(n2006) );
  XOR U2010 ( .A(creg[708]), .B(mod_mult_o[708]), .Z(n2008) );
  XNOR U2011 ( .A(n2009), .B(n2010), .Z(o[707]) );
  AND U2012 ( .A(n1035), .B(n2011), .Z(n2009) );
  XOR U2013 ( .A(creg[707]), .B(mod_mult_o[707]), .Z(n2011) );
  XNOR U2014 ( .A(n2012), .B(n2013), .Z(o[706]) );
  AND U2015 ( .A(n1035), .B(n2014), .Z(n2012) );
  XOR U2016 ( .A(creg[706]), .B(mod_mult_o[706]), .Z(n2014) );
  XNOR U2017 ( .A(n2015), .B(n2016), .Z(o[705]) );
  AND U2018 ( .A(n1035), .B(n2017), .Z(n2015) );
  XOR U2019 ( .A(creg[705]), .B(mod_mult_o[705]), .Z(n2017) );
  XNOR U2020 ( .A(n2018), .B(n2019), .Z(o[704]) );
  AND U2021 ( .A(n1035), .B(n2020), .Z(n2018) );
  XOR U2022 ( .A(creg[704]), .B(mod_mult_o[704]), .Z(n2020) );
  XNOR U2023 ( .A(n2021), .B(n2022), .Z(o[703]) );
  AND U2024 ( .A(n1035), .B(n2023), .Z(n2021) );
  XOR U2025 ( .A(creg[703]), .B(mod_mult_o[703]), .Z(n2023) );
  XNOR U2026 ( .A(n2024), .B(n2025), .Z(o[702]) );
  AND U2027 ( .A(n1035), .B(n2026), .Z(n2024) );
  XOR U2028 ( .A(creg[702]), .B(mod_mult_o[702]), .Z(n2026) );
  XNOR U2029 ( .A(n2027), .B(n2028), .Z(o[701]) );
  AND U2030 ( .A(n1035), .B(n2029), .Z(n2027) );
  XOR U2031 ( .A(creg[701]), .B(mod_mult_o[701]), .Z(n2029) );
  XNOR U2032 ( .A(n2030), .B(n2031), .Z(o[700]) );
  AND U2033 ( .A(n1035), .B(n2032), .Z(n2030) );
  XOR U2034 ( .A(creg[700]), .B(mod_mult_o[700]), .Z(n2032) );
  XNOR U2035 ( .A(n2033), .B(n2034), .Z(o[6]) );
  AND U2036 ( .A(n1035), .B(n2035), .Z(n2033) );
  XOR U2037 ( .A(creg[6]), .B(mod_mult_o[6]), .Z(n2035) );
  XNOR U2038 ( .A(n2036), .B(n2037), .Z(o[69]) );
  AND U2039 ( .A(n1035), .B(n2038), .Z(n2036) );
  XOR U2040 ( .A(creg[69]), .B(mod_mult_o[69]), .Z(n2038) );
  XNOR U2041 ( .A(n2039), .B(n2040), .Z(o[699]) );
  AND U2042 ( .A(n1035), .B(n2041), .Z(n2039) );
  XOR U2043 ( .A(creg[699]), .B(mod_mult_o[699]), .Z(n2041) );
  XNOR U2044 ( .A(n2042), .B(n2043), .Z(o[698]) );
  AND U2045 ( .A(n1035), .B(n2044), .Z(n2042) );
  XOR U2046 ( .A(creg[698]), .B(mod_mult_o[698]), .Z(n2044) );
  XNOR U2047 ( .A(n2045), .B(n2046), .Z(o[697]) );
  AND U2048 ( .A(n1035), .B(n2047), .Z(n2045) );
  XOR U2049 ( .A(creg[697]), .B(mod_mult_o[697]), .Z(n2047) );
  XNOR U2050 ( .A(n2048), .B(n2049), .Z(o[696]) );
  AND U2051 ( .A(n1035), .B(n2050), .Z(n2048) );
  XOR U2052 ( .A(creg[696]), .B(mod_mult_o[696]), .Z(n2050) );
  XNOR U2053 ( .A(n2051), .B(n2052), .Z(o[695]) );
  AND U2054 ( .A(n1035), .B(n2053), .Z(n2051) );
  XOR U2055 ( .A(creg[695]), .B(mod_mult_o[695]), .Z(n2053) );
  XNOR U2056 ( .A(n2054), .B(n2055), .Z(o[694]) );
  AND U2057 ( .A(n1035), .B(n2056), .Z(n2054) );
  XOR U2058 ( .A(creg[694]), .B(mod_mult_o[694]), .Z(n2056) );
  XNOR U2059 ( .A(n2057), .B(n2058), .Z(o[693]) );
  AND U2060 ( .A(n1035), .B(n2059), .Z(n2057) );
  XOR U2061 ( .A(creg[693]), .B(mod_mult_o[693]), .Z(n2059) );
  XNOR U2062 ( .A(n2060), .B(n2061), .Z(o[692]) );
  AND U2063 ( .A(n1035), .B(n2062), .Z(n2060) );
  XOR U2064 ( .A(creg[692]), .B(mod_mult_o[692]), .Z(n2062) );
  XNOR U2065 ( .A(n2063), .B(n2064), .Z(o[691]) );
  AND U2066 ( .A(n1035), .B(n2065), .Z(n2063) );
  XOR U2067 ( .A(creg[691]), .B(mod_mult_o[691]), .Z(n2065) );
  XNOR U2068 ( .A(n2066), .B(n2067), .Z(o[690]) );
  AND U2069 ( .A(n1035), .B(n2068), .Z(n2066) );
  XOR U2070 ( .A(creg[690]), .B(mod_mult_o[690]), .Z(n2068) );
  XNOR U2071 ( .A(n2069), .B(n2070), .Z(o[68]) );
  AND U2072 ( .A(n1035), .B(n2071), .Z(n2069) );
  XOR U2073 ( .A(creg[68]), .B(mod_mult_o[68]), .Z(n2071) );
  XNOR U2074 ( .A(n2072), .B(n2073), .Z(o[689]) );
  AND U2075 ( .A(n1035), .B(n2074), .Z(n2072) );
  XOR U2076 ( .A(creg[689]), .B(mod_mult_o[689]), .Z(n2074) );
  XNOR U2077 ( .A(n2075), .B(n2076), .Z(o[688]) );
  AND U2078 ( .A(n1035), .B(n2077), .Z(n2075) );
  XOR U2079 ( .A(creg[688]), .B(mod_mult_o[688]), .Z(n2077) );
  XNOR U2080 ( .A(n2078), .B(n2079), .Z(o[687]) );
  AND U2081 ( .A(n1035), .B(n2080), .Z(n2078) );
  XOR U2082 ( .A(creg[687]), .B(mod_mult_o[687]), .Z(n2080) );
  XNOR U2083 ( .A(n2081), .B(n2082), .Z(o[686]) );
  AND U2084 ( .A(n1035), .B(n2083), .Z(n2081) );
  XOR U2085 ( .A(creg[686]), .B(mod_mult_o[686]), .Z(n2083) );
  XNOR U2086 ( .A(n2084), .B(n2085), .Z(o[685]) );
  AND U2087 ( .A(n1035), .B(n2086), .Z(n2084) );
  XOR U2088 ( .A(creg[685]), .B(mod_mult_o[685]), .Z(n2086) );
  XNOR U2089 ( .A(n2087), .B(n2088), .Z(o[684]) );
  AND U2090 ( .A(n1035), .B(n2089), .Z(n2087) );
  XOR U2091 ( .A(creg[684]), .B(mod_mult_o[684]), .Z(n2089) );
  XNOR U2092 ( .A(n2090), .B(n2091), .Z(o[683]) );
  AND U2093 ( .A(n1035), .B(n2092), .Z(n2090) );
  XOR U2094 ( .A(creg[683]), .B(mod_mult_o[683]), .Z(n2092) );
  XNOR U2095 ( .A(n2093), .B(n2094), .Z(o[682]) );
  AND U2096 ( .A(n1035), .B(n2095), .Z(n2093) );
  XOR U2097 ( .A(creg[682]), .B(mod_mult_o[682]), .Z(n2095) );
  XNOR U2098 ( .A(n2096), .B(n2097), .Z(o[681]) );
  AND U2099 ( .A(n1035), .B(n2098), .Z(n2096) );
  XOR U2100 ( .A(creg[681]), .B(mod_mult_o[681]), .Z(n2098) );
  XNOR U2101 ( .A(n2099), .B(n2100), .Z(o[680]) );
  AND U2102 ( .A(n1035), .B(n2101), .Z(n2099) );
  XOR U2103 ( .A(creg[680]), .B(mod_mult_o[680]), .Z(n2101) );
  XNOR U2104 ( .A(n2102), .B(n2103), .Z(o[67]) );
  AND U2105 ( .A(n1035), .B(n2104), .Z(n2102) );
  XOR U2106 ( .A(creg[67]), .B(mod_mult_o[67]), .Z(n2104) );
  XNOR U2107 ( .A(n2105), .B(n2106), .Z(o[679]) );
  AND U2108 ( .A(n1035), .B(n2107), .Z(n2105) );
  XOR U2109 ( .A(creg[679]), .B(mod_mult_o[679]), .Z(n2107) );
  XNOR U2110 ( .A(n2108), .B(n2109), .Z(o[678]) );
  AND U2111 ( .A(n1035), .B(n2110), .Z(n2108) );
  XOR U2112 ( .A(creg[678]), .B(mod_mult_o[678]), .Z(n2110) );
  XNOR U2113 ( .A(n2111), .B(n2112), .Z(o[677]) );
  AND U2114 ( .A(n1035), .B(n2113), .Z(n2111) );
  XOR U2115 ( .A(creg[677]), .B(mod_mult_o[677]), .Z(n2113) );
  XNOR U2116 ( .A(n2114), .B(n2115), .Z(o[676]) );
  AND U2117 ( .A(n1035), .B(n2116), .Z(n2114) );
  XOR U2118 ( .A(creg[676]), .B(mod_mult_o[676]), .Z(n2116) );
  XNOR U2119 ( .A(n2117), .B(n2118), .Z(o[675]) );
  AND U2120 ( .A(n1035), .B(n2119), .Z(n2117) );
  XOR U2121 ( .A(creg[675]), .B(mod_mult_o[675]), .Z(n2119) );
  XNOR U2122 ( .A(n2120), .B(n2121), .Z(o[674]) );
  AND U2123 ( .A(n1035), .B(n2122), .Z(n2120) );
  XOR U2124 ( .A(creg[674]), .B(mod_mult_o[674]), .Z(n2122) );
  XNOR U2125 ( .A(n2123), .B(n2124), .Z(o[673]) );
  AND U2126 ( .A(n1035), .B(n2125), .Z(n2123) );
  XOR U2127 ( .A(creg[673]), .B(mod_mult_o[673]), .Z(n2125) );
  XNOR U2128 ( .A(n2126), .B(n2127), .Z(o[672]) );
  AND U2129 ( .A(n1035), .B(n2128), .Z(n2126) );
  XOR U2130 ( .A(creg[672]), .B(mod_mult_o[672]), .Z(n2128) );
  XNOR U2131 ( .A(n2129), .B(n2130), .Z(o[671]) );
  AND U2132 ( .A(n1035), .B(n2131), .Z(n2129) );
  XOR U2133 ( .A(creg[671]), .B(mod_mult_o[671]), .Z(n2131) );
  XNOR U2134 ( .A(n2132), .B(n2133), .Z(o[670]) );
  AND U2135 ( .A(n1035), .B(n2134), .Z(n2132) );
  XOR U2136 ( .A(creg[670]), .B(mod_mult_o[670]), .Z(n2134) );
  XNOR U2137 ( .A(n2135), .B(n2136), .Z(o[66]) );
  AND U2138 ( .A(n1035), .B(n2137), .Z(n2135) );
  XOR U2139 ( .A(creg[66]), .B(mod_mult_o[66]), .Z(n2137) );
  XNOR U2140 ( .A(n2138), .B(n2139), .Z(o[669]) );
  AND U2141 ( .A(n1035), .B(n2140), .Z(n2138) );
  XOR U2142 ( .A(creg[669]), .B(mod_mult_o[669]), .Z(n2140) );
  XNOR U2143 ( .A(n2141), .B(n2142), .Z(o[668]) );
  AND U2144 ( .A(n1035), .B(n2143), .Z(n2141) );
  XOR U2145 ( .A(creg[668]), .B(mod_mult_o[668]), .Z(n2143) );
  XNOR U2146 ( .A(n2144), .B(n2145), .Z(o[667]) );
  AND U2147 ( .A(n1035), .B(n2146), .Z(n2144) );
  XOR U2148 ( .A(creg[667]), .B(mod_mult_o[667]), .Z(n2146) );
  XNOR U2149 ( .A(n2147), .B(n2148), .Z(o[666]) );
  AND U2150 ( .A(n1035), .B(n2149), .Z(n2147) );
  XOR U2151 ( .A(creg[666]), .B(mod_mult_o[666]), .Z(n2149) );
  XNOR U2152 ( .A(n2150), .B(n2151), .Z(o[665]) );
  AND U2153 ( .A(n1035), .B(n2152), .Z(n2150) );
  XOR U2154 ( .A(creg[665]), .B(mod_mult_o[665]), .Z(n2152) );
  XNOR U2155 ( .A(n2153), .B(n2154), .Z(o[664]) );
  AND U2156 ( .A(n1035), .B(n2155), .Z(n2153) );
  XOR U2157 ( .A(creg[664]), .B(mod_mult_o[664]), .Z(n2155) );
  XNOR U2158 ( .A(n2156), .B(n2157), .Z(o[663]) );
  AND U2159 ( .A(n1035), .B(n2158), .Z(n2156) );
  XOR U2160 ( .A(creg[663]), .B(mod_mult_o[663]), .Z(n2158) );
  XNOR U2161 ( .A(n2159), .B(n2160), .Z(o[662]) );
  AND U2162 ( .A(n1035), .B(n2161), .Z(n2159) );
  XOR U2163 ( .A(creg[662]), .B(mod_mult_o[662]), .Z(n2161) );
  XNOR U2164 ( .A(n2162), .B(n2163), .Z(o[661]) );
  AND U2165 ( .A(n1035), .B(n2164), .Z(n2162) );
  XOR U2166 ( .A(creg[661]), .B(mod_mult_o[661]), .Z(n2164) );
  XNOR U2167 ( .A(n2165), .B(n2166), .Z(o[660]) );
  AND U2168 ( .A(n1035), .B(n2167), .Z(n2165) );
  XOR U2169 ( .A(creg[660]), .B(mod_mult_o[660]), .Z(n2167) );
  XNOR U2170 ( .A(n2168), .B(n2169), .Z(o[65]) );
  AND U2171 ( .A(n1035), .B(n2170), .Z(n2168) );
  XOR U2172 ( .A(creg[65]), .B(mod_mult_o[65]), .Z(n2170) );
  XNOR U2173 ( .A(n2171), .B(n2172), .Z(o[659]) );
  AND U2174 ( .A(n1035), .B(n2173), .Z(n2171) );
  XOR U2175 ( .A(creg[659]), .B(mod_mult_o[659]), .Z(n2173) );
  XNOR U2176 ( .A(n2174), .B(n2175), .Z(o[658]) );
  AND U2177 ( .A(n1035), .B(n2176), .Z(n2174) );
  XOR U2178 ( .A(creg[658]), .B(mod_mult_o[658]), .Z(n2176) );
  XNOR U2179 ( .A(n2177), .B(n2178), .Z(o[657]) );
  AND U2180 ( .A(n1035), .B(n2179), .Z(n2177) );
  XOR U2181 ( .A(creg[657]), .B(mod_mult_o[657]), .Z(n2179) );
  XNOR U2182 ( .A(n2180), .B(n2181), .Z(o[656]) );
  AND U2183 ( .A(n1035), .B(n2182), .Z(n2180) );
  XOR U2184 ( .A(creg[656]), .B(mod_mult_o[656]), .Z(n2182) );
  XNOR U2185 ( .A(n2183), .B(n2184), .Z(o[655]) );
  AND U2186 ( .A(n1035), .B(n2185), .Z(n2183) );
  XOR U2187 ( .A(creg[655]), .B(mod_mult_o[655]), .Z(n2185) );
  XNOR U2188 ( .A(n2186), .B(n2187), .Z(o[654]) );
  AND U2189 ( .A(n1035), .B(n2188), .Z(n2186) );
  XOR U2190 ( .A(creg[654]), .B(mod_mult_o[654]), .Z(n2188) );
  XNOR U2191 ( .A(n2189), .B(n2190), .Z(o[653]) );
  AND U2192 ( .A(n1035), .B(n2191), .Z(n2189) );
  XOR U2193 ( .A(creg[653]), .B(mod_mult_o[653]), .Z(n2191) );
  XNOR U2194 ( .A(n2192), .B(n2193), .Z(o[652]) );
  AND U2195 ( .A(n1035), .B(n2194), .Z(n2192) );
  XOR U2196 ( .A(creg[652]), .B(mod_mult_o[652]), .Z(n2194) );
  XNOR U2197 ( .A(n2195), .B(n2196), .Z(o[651]) );
  AND U2198 ( .A(n1035), .B(n2197), .Z(n2195) );
  XOR U2199 ( .A(creg[651]), .B(mod_mult_o[651]), .Z(n2197) );
  XNOR U2200 ( .A(n2198), .B(n2199), .Z(o[650]) );
  AND U2201 ( .A(n1035), .B(n2200), .Z(n2198) );
  XOR U2202 ( .A(creg[650]), .B(mod_mult_o[650]), .Z(n2200) );
  XNOR U2203 ( .A(n2201), .B(n2202), .Z(o[64]) );
  AND U2204 ( .A(n1035), .B(n2203), .Z(n2201) );
  XOR U2205 ( .A(creg[64]), .B(mod_mult_o[64]), .Z(n2203) );
  XNOR U2206 ( .A(n2204), .B(n2205), .Z(o[649]) );
  AND U2207 ( .A(n1035), .B(n2206), .Z(n2204) );
  XOR U2208 ( .A(creg[649]), .B(mod_mult_o[649]), .Z(n2206) );
  XNOR U2209 ( .A(n2207), .B(n2208), .Z(o[648]) );
  AND U2210 ( .A(n1035), .B(n2209), .Z(n2207) );
  XOR U2211 ( .A(creg[648]), .B(mod_mult_o[648]), .Z(n2209) );
  XNOR U2212 ( .A(n2210), .B(n2211), .Z(o[647]) );
  AND U2213 ( .A(n1035), .B(n2212), .Z(n2210) );
  XOR U2214 ( .A(creg[647]), .B(mod_mult_o[647]), .Z(n2212) );
  XNOR U2215 ( .A(n2213), .B(n2214), .Z(o[646]) );
  AND U2216 ( .A(n1035), .B(n2215), .Z(n2213) );
  XOR U2217 ( .A(creg[646]), .B(mod_mult_o[646]), .Z(n2215) );
  XNOR U2218 ( .A(n2216), .B(n2217), .Z(o[645]) );
  AND U2219 ( .A(n1035), .B(n2218), .Z(n2216) );
  XOR U2220 ( .A(creg[645]), .B(mod_mult_o[645]), .Z(n2218) );
  XNOR U2221 ( .A(n2219), .B(n2220), .Z(o[644]) );
  AND U2222 ( .A(n1035), .B(n2221), .Z(n2219) );
  XOR U2223 ( .A(creg[644]), .B(mod_mult_o[644]), .Z(n2221) );
  XNOR U2224 ( .A(n2222), .B(n2223), .Z(o[643]) );
  AND U2225 ( .A(n1035), .B(n2224), .Z(n2222) );
  XOR U2226 ( .A(creg[643]), .B(mod_mult_o[643]), .Z(n2224) );
  XNOR U2227 ( .A(n2225), .B(n2226), .Z(o[642]) );
  AND U2228 ( .A(n1035), .B(n2227), .Z(n2225) );
  XOR U2229 ( .A(creg[642]), .B(mod_mult_o[642]), .Z(n2227) );
  XNOR U2230 ( .A(n2228), .B(n2229), .Z(o[641]) );
  AND U2231 ( .A(n1035), .B(n2230), .Z(n2228) );
  XOR U2232 ( .A(creg[641]), .B(mod_mult_o[641]), .Z(n2230) );
  XNOR U2233 ( .A(n2231), .B(n2232), .Z(o[640]) );
  AND U2234 ( .A(n1035), .B(n2233), .Z(n2231) );
  XOR U2235 ( .A(creg[640]), .B(mod_mult_o[640]), .Z(n2233) );
  XNOR U2236 ( .A(n2234), .B(n2235), .Z(o[63]) );
  AND U2237 ( .A(n1035), .B(n2236), .Z(n2234) );
  XOR U2238 ( .A(creg[63]), .B(mod_mult_o[63]), .Z(n2236) );
  XNOR U2239 ( .A(n2237), .B(n2238), .Z(o[639]) );
  AND U2240 ( .A(n1035), .B(n2239), .Z(n2237) );
  XOR U2241 ( .A(creg[639]), .B(mod_mult_o[639]), .Z(n2239) );
  XNOR U2242 ( .A(n2240), .B(n2241), .Z(o[638]) );
  AND U2243 ( .A(n1035), .B(n2242), .Z(n2240) );
  XOR U2244 ( .A(creg[638]), .B(mod_mult_o[638]), .Z(n2242) );
  XNOR U2245 ( .A(n2243), .B(n2244), .Z(o[637]) );
  AND U2246 ( .A(n1035), .B(n2245), .Z(n2243) );
  XOR U2247 ( .A(creg[637]), .B(mod_mult_o[637]), .Z(n2245) );
  XNOR U2248 ( .A(n2246), .B(n2247), .Z(o[636]) );
  AND U2249 ( .A(n1035), .B(n2248), .Z(n2246) );
  XOR U2250 ( .A(creg[636]), .B(mod_mult_o[636]), .Z(n2248) );
  XNOR U2251 ( .A(n2249), .B(n2250), .Z(o[635]) );
  AND U2252 ( .A(n1035), .B(n2251), .Z(n2249) );
  XOR U2253 ( .A(creg[635]), .B(mod_mult_o[635]), .Z(n2251) );
  XNOR U2254 ( .A(n2252), .B(n2253), .Z(o[634]) );
  AND U2255 ( .A(n1035), .B(n2254), .Z(n2252) );
  XOR U2256 ( .A(creg[634]), .B(mod_mult_o[634]), .Z(n2254) );
  XNOR U2257 ( .A(n2255), .B(n2256), .Z(o[633]) );
  AND U2258 ( .A(n1035), .B(n2257), .Z(n2255) );
  XOR U2259 ( .A(creg[633]), .B(mod_mult_o[633]), .Z(n2257) );
  XNOR U2260 ( .A(n2258), .B(n2259), .Z(o[632]) );
  AND U2261 ( .A(n1035), .B(n2260), .Z(n2258) );
  XOR U2262 ( .A(creg[632]), .B(mod_mult_o[632]), .Z(n2260) );
  XNOR U2263 ( .A(n2261), .B(n2262), .Z(o[631]) );
  AND U2264 ( .A(n1035), .B(n2263), .Z(n2261) );
  XOR U2265 ( .A(creg[631]), .B(mod_mult_o[631]), .Z(n2263) );
  XNOR U2266 ( .A(n2264), .B(n2265), .Z(o[630]) );
  AND U2267 ( .A(n1035), .B(n2266), .Z(n2264) );
  XOR U2268 ( .A(creg[630]), .B(mod_mult_o[630]), .Z(n2266) );
  XNOR U2269 ( .A(n2267), .B(n2268), .Z(o[62]) );
  AND U2270 ( .A(n1035), .B(n2269), .Z(n2267) );
  XOR U2271 ( .A(creg[62]), .B(mod_mult_o[62]), .Z(n2269) );
  XNOR U2272 ( .A(n2270), .B(n2271), .Z(o[629]) );
  AND U2273 ( .A(n1035), .B(n2272), .Z(n2270) );
  XOR U2274 ( .A(creg[629]), .B(mod_mult_o[629]), .Z(n2272) );
  XNOR U2275 ( .A(n2273), .B(n2274), .Z(o[628]) );
  AND U2276 ( .A(n1035), .B(n2275), .Z(n2273) );
  XOR U2277 ( .A(creg[628]), .B(mod_mult_o[628]), .Z(n2275) );
  XNOR U2278 ( .A(n2276), .B(n2277), .Z(o[627]) );
  AND U2279 ( .A(n1035), .B(n2278), .Z(n2276) );
  XOR U2280 ( .A(creg[627]), .B(mod_mult_o[627]), .Z(n2278) );
  XNOR U2281 ( .A(n2279), .B(n2280), .Z(o[626]) );
  AND U2282 ( .A(n1035), .B(n2281), .Z(n2279) );
  XOR U2283 ( .A(creg[626]), .B(mod_mult_o[626]), .Z(n2281) );
  XNOR U2284 ( .A(n2282), .B(n2283), .Z(o[625]) );
  AND U2285 ( .A(n1035), .B(n2284), .Z(n2282) );
  XOR U2286 ( .A(creg[625]), .B(mod_mult_o[625]), .Z(n2284) );
  XNOR U2287 ( .A(n2285), .B(n2286), .Z(o[624]) );
  AND U2288 ( .A(n1035), .B(n2287), .Z(n2285) );
  XOR U2289 ( .A(creg[624]), .B(mod_mult_o[624]), .Z(n2287) );
  XNOR U2290 ( .A(n2288), .B(n2289), .Z(o[623]) );
  AND U2291 ( .A(n1035), .B(n2290), .Z(n2288) );
  XOR U2292 ( .A(creg[623]), .B(mod_mult_o[623]), .Z(n2290) );
  XNOR U2293 ( .A(n2291), .B(n2292), .Z(o[622]) );
  AND U2294 ( .A(n1035), .B(n2293), .Z(n2291) );
  XOR U2295 ( .A(creg[622]), .B(mod_mult_o[622]), .Z(n2293) );
  XNOR U2296 ( .A(n2294), .B(n2295), .Z(o[621]) );
  AND U2297 ( .A(n1035), .B(n2296), .Z(n2294) );
  XOR U2298 ( .A(creg[621]), .B(mod_mult_o[621]), .Z(n2296) );
  XNOR U2299 ( .A(n2297), .B(n2298), .Z(o[620]) );
  AND U2300 ( .A(n1035), .B(n2299), .Z(n2297) );
  XOR U2301 ( .A(creg[620]), .B(mod_mult_o[620]), .Z(n2299) );
  XNOR U2302 ( .A(n2300), .B(n2301), .Z(o[61]) );
  AND U2303 ( .A(n1035), .B(n2302), .Z(n2300) );
  XOR U2304 ( .A(creg[61]), .B(mod_mult_o[61]), .Z(n2302) );
  XNOR U2305 ( .A(n2303), .B(n2304), .Z(o[619]) );
  AND U2306 ( .A(n1035), .B(n2305), .Z(n2303) );
  XOR U2307 ( .A(creg[619]), .B(mod_mult_o[619]), .Z(n2305) );
  XNOR U2308 ( .A(n2306), .B(n2307), .Z(o[618]) );
  AND U2309 ( .A(n1035), .B(n2308), .Z(n2306) );
  XOR U2310 ( .A(creg[618]), .B(mod_mult_o[618]), .Z(n2308) );
  XNOR U2311 ( .A(n2309), .B(n2310), .Z(o[617]) );
  AND U2312 ( .A(n1035), .B(n2311), .Z(n2309) );
  XOR U2313 ( .A(creg[617]), .B(mod_mult_o[617]), .Z(n2311) );
  XNOR U2314 ( .A(n2312), .B(n2313), .Z(o[616]) );
  AND U2315 ( .A(n1035), .B(n2314), .Z(n2312) );
  XOR U2316 ( .A(creg[616]), .B(mod_mult_o[616]), .Z(n2314) );
  XNOR U2317 ( .A(n2315), .B(n2316), .Z(o[615]) );
  AND U2318 ( .A(n1035), .B(n2317), .Z(n2315) );
  XOR U2319 ( .A(creg[615]), .B(mod_mult_o[615]), .Z(n2317) );
  XNOR U2320 ( .A(n2318), .B(n2319), .Z(o[614]) );
  AND U2321 ( .A(n1035), .B(n2320), .Z(n2318) );
  XOR U2322 ( .A(creg[614]), .B(mod_mult_o[614]), .Z(n2320) );
  XNOR U2323 ( .A(n2321), .B(n2322), .Z(o[613]) );
  AND U2324 ( .A(n1035), .B(n2323), .Z(n2321) );
  XOR U2325 ( .A(creg[613]), .B(mod_mult_o[613]), .Z(n2323) );
  XNOR U2326 ( .A(n2324), .B(n2325), .Z(o[612]) );
  AND U2327 ( .A(n1035), .B(n2326), .Z(n2324) );
  XOR U2328 ( .A(creg[612]), .B(mod_mult_o[612]), .Z(n2326) );
  XNOR U2329 ( .A(n2327), .B(n2328), .Z(o[611]) );
  AND U2330 ( .A(n1035), .B(n2329), .Z(n2327) );
  XOR U2331 ( .A(creg[611]), .B(mod_mult_o[611]), .Z(n2329) );
  XNOR U2332 ( .A(n2330), .B(n2331), .Z(o[610]) );
  AND U2333 ( .A(n1035), .B(n2332), .Z(n2330) );
  XOR U2334 ( .A(creg[610]), .B(mod_mult_o[610]), .Z(n2332) );
  XNOR U2335 ( .A(n2333), .B(n2334), .Z(o[60]) );
  AND U2336 ( .A(n1035), .B(n2335), .Z(n2333) );
  XOR U2337 ( .A(creg[60]), .B(mod_mult_o[60]), .Z(n2335) );
  XNOR U2338 ( .A(n2336), .B(n2337), .Z(o[609]) );
  AND U2339 ( .A(n1035), .B(n2338), .Z(n2336) );
  XOR U2340 ( .A(creg[609]), .B(mod_mult_o[609]), .Z(n2338) );
  XNOR U2341 ( .A(n2339), .B(n2340), .Z(o[608]) );
  AND U2342 ( .A(n1035), .B(n2341), .Z(n2339) );
  XOR U2343 ( .A(creg[608]), .B(mod_mult_o[608]), .Z(n2341) );
  XNOR U2344 ( .A(n2342), .B(n2343), .Z(o[607]) );
  AND U2345 ( .A(n1035), .B(n2344), .Z(n2342) );
  XOR U2346 ( .A(creg[607]), .B(mod_mult_o[607]), .Z(n2344) );
  XNOR U2347 ( .A(n2345), .B(n2346), .Z(o[606]) );
  AND U2348 ( .A(n1035), .B(n2347), .Z(n2345) );
  XOR U2349 ( .A(creg[606]), .B(mod_mult_o[606]), .Z(n2347) );
  XNOR U2350 ( .A(n2348), .B(n2349), .Z(o[605]) );
  AND U2351 ( .A(n1035), .B(n2350), .Z(n2348) );
  XOR U2352 ( .A(creg[605]), .B(mod_mult_o[605]), .Z(n2350) );
  XNOR U2353 ( .A(n2351), .B(n2352), .Z(o[604]) );
  AND U2354 ( .A(n1035), .B(n2353), .Z(n2351) );
  XOR U2355 ( .A(creg[604]), .B(mod_mult_o[604]), .Z(n2353) );
  XNOR U2356 ( .A(n2354), .B(n2355), .Z(o[603]) );
  AND U2357 ( .A(n1035), .B(n2356), .Z(n2354) );
  XOR U2358 ( .A(creg[603]), .B(mod_mult_o[603]), .Z(n2356) );
  XNOR U2359 ( .A(n2357), .B(n2358), .Z(o[602]) );
  AND U2360 ( .A(n1035), .B(n2359), .Z(n2357) );
  XOR U2361 ( .A(creg[602]), .B(mod_mult_o[602]), .Z(n2359) );
  XNOR U2362 ( .A(n2360), .B(n2361), .Z(o[601]) );
  AND U2363 ( .A(n1035), .B(n2362), .Z(n2360) );
  XOR U2364 ( .A(creg[601]), .B(mod_mult_o[601]), .Z(n2362) );
  XNOR U2365 ( .A(n2363), .B(n2364), .Z(o[600]) );
  AND U2366 ( .A(n1035), .B(n2365), .Z(n2363) );
  XOR U2367 ( .A(creg[600]), .B(mod_mult_o[600]), .Z(n2365) );
  XNOR U2368 ( .A(n2366), .B(n2367), .Z(o[5]) );
  AND U2369 ( .A(n1035), .B(n2368), .Z(n2366) );
  XOR U2370 ( .A(creg[5]), .B(mod_mult_o[5]), .Z(n2368) );
  XNOR U2371 ( .A(n2369), .B(n2370), .Z(o[59]) );
  AND U2372 ( .A(n1035), .B(n2371), .Z(n2369) );
  XOR U2373 ( .A(creg[59]), .B(mod_mult_o[59]), .Z(n2371) );
  XNOR U2374 ( .A(n2372), .B(n2373), .Z(o[599]) );
  AND U2375 ( .A(n1035), .B(n2374), .Z(n2372) );
  XOR U2376 ( .A(creg[599]), .B(mod_mult_o[599]), .Z(n2374) );
  XNOR U2377 ( .A(n2375), .B(n2376), .Z(o[598]) );
  AND U2378 ( .A(n1035), .B(n2377), .Z(n2375) );
  XOR U2379 ( .A(creg[598]), .B(mod_mult_o[598]), .Z(n2377) );
  XNOR U2380 ( .A(n2378), .B(n2379), .Z(o[597]) );
  AND U2381 ( .A(n1035), .B(n2380), .Z(n2378) );
  XOR U2382 ( .A(creg[597]), .B(mod_mult_o[597]), .Z(n2380) );
  XNOR U2383 ( .A(n2381), .B(n2382), .Z(o[596]) );
  AND U2384 ( .A(n1035), .B(n2383), .Z(n2381) );
  XOR U2385 ( .A(creg[596]), .B(mod_mult_o[596]), .Z(n2383) );
  XNOR U2386 ( .A(n2384), .B(n2385), .Z(o[595]) );
  AND U2387 ( .A(n1035), .B(n2386), .Z(n2384) );
  XOR U2388 ( .A(creg[595]), .B(mod_mult_o[595]), .Z(n2386) );
  XNOR U2389 ( .A(n2387), .B(n2388), .Z(o[594]) );
  AND U2390 ( .A(n1035), .B(n2389), .Z(n2387) );
  XOR U2391 ( .A(creg[594]), .B(mod_mult_o[594]), .Z(n2389) );
  XNOR U2392 ( .A(n2390), .B(n2391), .Z(o[593]) );
  AND U2393 ( .A(n1035), .B(n2392), .Z(n2390) );
  XOR U2394 ( .A(creg[593]), .B(mod_mult_o[593]), .Z(n2392) );
  XNOR U2395 ( .A(n2393), .B(n2394), .Z(o[592]) );
  AND U2396 ( .A(n1035), .B(n2395), .Z(n2393) );
  XOR U2397 ( .A(creg[592]), .B(mod_mult_o[592]), .Z(n2395) );
  XNOR U2398 ( .A(n2396), .B(n2397), .Z(o[591]) );
  AND U2399 ( .A(n1035), .B(n2398), .Z(n2396) );
  XOR U2400 ( .A(creg[591]), .B(mod_mult_o[591]), .Z(n2398) );
  XNOR U2401 ( .A(n2399), .B(n2400), .Z(o[590]) );
  AND U2402 ( .A(n1035), .B(n2401), .Z(n2399) );
  XOR U2403 ( .A(creg[590]), .B(mod_mult_o[590]), .Z(n2401) );
  XNOR U2404 ( .A(n2402), .B(n2403), .Z(o[58]) );
  AND U2405 ( .A(n1035), .B(n2404), .Z(n2402) );
  XOR U2406 ( .A(creg[58]), .B(mod_mult_o[58]), .Z(n2404) );
  XNOR U2407 ( .A(n2405), .B(n2406), .Z(o[589]) );
  AND U2408 ( .A(n1035), .B(n2407), .Z(n2405) );
  XOR U2409 ( .A(creg[589]), .B(mod_mult_o[589]), .Z(n2407) );
  XNOR U2410 ( .A(n2408), .B(n2409), .Z(o[588]) );
  AND U2411 ( .A(n1035), .B(n2410), .Z(n2408) );
  XOR U2412 ( .A(creg[588]), .B(mod_mult_o[588]), .Z(n2410) );
  XNOR U2413 ( .A(n2411), .B(n2412), .Z(o[587]) );
  AND U2414 ( .A(n1035), .B(n2413), .Z(n2411) );
  XOR U2415 ( .A(creg[587]), .B(mod_mult_o[587]), .Z(n2413) );
  XNOR U2416 ( .A(n2414), .B(n2415), .Z(o[586]) );
  AND U2417 ( .A(n1035), .B(n2416), .Z(n2414) );
  XOR U2418 ( .A(creg[586]), .B(mod_mult_o[586]), .Z(n2416) );
  XNOR U2419 ( .A(n2417), .B(n2418), .Z(o[585]) );
  AND U2420 ( .A(n1035), .B(n2419), .Z(n2417) );
  XOR U2421 ( .A(creg[585]), .B(mod_mult_o[585]), .Z(n2419) );
  XNOR U2422 ( .A(n2420), .B(n2421), .Z(o[584]) );
  AND U2423 ( .A(n1035), .B(n2422), .Z(n2420) );
  XOR U2424 ( .A(creg[584]), .B(mod_mult_o[584]), .Z(n2422) );
  XNOR U2425 ( .A(n2423), .B(n2424), .Z(o[583]) );
  AND U2426 ( .A(n1035), .B(n2425), .Z(n2423) );
  XOR U2427 ( .A(creg[583]), .B(mod_mult_o[583]), .Z(n2425) );
  XNOR U2428 ( .A(n2426), .B(n2427), .Z(o[582]) );
  AND U2429 ( .A(n1035), .B(n2428), .Z(n2426) );
  XOR U2430 ( .A(creg[582]), .B(mod_mult_o[582]), .Z(n2428) );
  XNOR U2431 ( .A(n2429), .B(n2430), .Z(o[581]) );
  AND U2432 ( .A(n1035), .B(n2431), .Z(n2429) );
  XOR U2433 ( .A(creg[581]), .B(mod_mult_o[581]), .Z(n2431) );
  XNOR U2434 ( .A(n2432), .B(n2433), .Z(o[580]) );
  AND U2435 ( .A(n1035), .B(n2434), .Z(n2432) );
  XOR U2436 ( .A(creg[580]), .B(mod_mult_o[580]), .Z(n2434) );
  XNOR U2437 ( .A(n2435), .B(n2436), .Z(o[57]) );
  AND U2438 ( .A(n1035), .B(n2437), .Z(n2435) );
  XOR U2439 ( .A(creg[57]), .B(mod_mult_o[57]), .Z(n2437) );
  XNOR U2440 ( .A(n2438), .B(n2439), .Z(o[579]) );
  AND U2441 ( .A(n1035), .B(n2440), .Z(n2438) );
  XOR U2442 ( .A(creg[579]), .B(mod_mult_o[579]), .Z(n2440) );
  XNOR U2443 ( .A(n2441), .B(n2442), .Z(o[578]) );
  AND U2444 ( .A(n1035), .B(n2443), .Z(n2441) );
  XOR U2445 ( .A(creg[578]), .B(mod_mult_o[578]), .Z(n2443) );
  XNOR U2446 ( .A(n2444), .B(n2445), .Z(o[577]) );
  AND U2447 ( .A(n1035), .B(n2446), .Z(n2444) );
  XOR U2448 ( .A(creg[577]), .B(mod_mult_o[577]), .Z(n2446) );
  XNOR U2449 ( .A(n2447), .B(n2448), .Z(o[576]) );
  AND U2450 ( .A(n1035), .B(n2449), .Z(n2447) );
  XOR U2451 ( .A(creg[576]), .B(mod_mult_o[576]), .Z(n2449) );
  XNOR U2452 ( .A(n2450), .B(n2451), .Z(o[575]) );
  AND U2453 ( .A(n1035), .B(n2452), .Z(n2450) );
  XOR U2454 ( .A(creg[575]), .B(mod_mult_o[575]), .Z(n2452) );
  XNOR U2455 ( .A(n2453), .B(n2454), .Z(o[574]) );
  AND U2456 ( .A(n1035), .B(n2455), .Z(n2453) );
  XOR U2457 ( .A(creg[574]), .B(mod_mult_o[574]), .Z(n2455) );
  XNOR U2458 ( .A(n2456), .B(n2457), .Z(o[573]) );
  AND U2459 ( .A(n1035), .B(n2458), .Z(n2456) );
  XOR U2460 ( .A(creg[573]), .B(mod_mult_o[573]), .Z(n2458) );
  XNOR U2461 ( .A(n2459), .B(n2460), .Z(o[572]) );
  AND U2462 ( .A(n1035), .B(n2461), .Z(n2459) );
  XOR U2463 ( .A(creg[572]), .B(mod_mult_o[572]), .Z(n2461) );
  XNOR U2464 ( .A(n2462), .B(n2463), .Z(o[571]) );
  AND U2465 ( .A(n1035), .B(n2464), .Z(n2462) );
  XOR U2466 ( .A(creg[571]), .B(mod_mult_o[571]), .Z(n2464) );
  XNOR U2467 ( .A(n2465), .B(n2466), .Z(o[570]) );
  AND U2468 ( .A(n1035), .B(n2467), .Z(n2465) );
  XOR U2469 ( .A(creg[570]), .B(mod_mult_o[570]), .Z(n2467) );
  XNOR U2470 ( .A(n2468), .B(n2469), .Z(o[56]) );
  AND U2471 ( .A(n1035), .B(n2470), .Z(n2468) );
  XOR U2472 ( .A(creg[56]), .B(mod_mult_o[56]), .Z(n2470) );
  XNOR U2473 ( .A(n2471), .B(n2472), .Z(o[569]) );
  AND U2474 ( .A(n1035), .B(n2473), .Z(n2471) );
  XOR U2475 ( .A(creg[569]), .B(mod_mult_o[569]), .Z(n2473) );
  XNOR U2476 ( .A(n2474), .B(n2475), .Z(o[568]) );
  AND U2477 ( .A(n1035), .B(n2476), .Z(n2474) );
  XOR U2478 ( .A(creg[568]), .B(mod_mult_o[568]), .Z(n2476) );
  XNOR U2479 ( .A(n2477), .B(n2478), .Z(o[567]) );
  AND U2480 ( .A(n1035), .B(n2479), .Z(n2477) );
  XOR U2481 ( .A(creg[567]), .B(mod_mult_o[567]), .Z(n2479) );
  XNOR U2482 ( .A(n2480), .B(n2481), .Z(o[566]) );
  AND U2483 ( .A(n1035), .B(n2482), .Z(n2480) );
  XOR U2484 ( .A(creg[566]), .B(mod_mult_o[566]), .Z(n2482) );
  XNOR U2485 ( .A(n2483), .B(n2484), .Z(o[565]) );
  AND U2486 ( .A(n1035), .B(n2485), .Z(n2483) );
  XOR U2487 ( .A(creg[565]), .B(mod_mult_o[565]), .Z(n2485) );
  XNOR U2488 ( .A(n2486), .B(n2487), .Z(o[564]) );
  AND U2489 ( .A(n1035), .B(n2488), .Z(n2486) );
  XOR U2490 ( .A(creg[564]), .B(mod_mult_o[564]), .Z(n2488) );
  XNOR U2491 ( .A(n2489), .B(n2490), .Z(o[563]) );
  AND U2492 ( .A(n1035), .B(n2491), .Z(n2489) );
  XOR U2493 ( .A(creg[563]), .B(mod_mult_o[563]), .Z(n2491) );
  XNOR U2494 ( .A(n2492), .B(n2493), .Z(o[562]) );
  AND U2495 ( .A(n1035), .B(n2494), .Z(n2492) );
  XOR U2496 ( .A(creg[562]), .B(mod_mult_o[562]), .Z(n2494) );
  XNOR U2497 ( .A(n2495), .B(n2496), .Z(o[561]) );
  AND U2498 ( .A(n1035), .B(n2497), .Z(n2495) );
  XOR U2499 ( .A(creg[561]), .B(mod_mult_o[561]), .Z(n2497) );
  XNOR U2500 ( .A(n2498), .B(n2499), .Z(o[560]) );
  AND U2501 ( .A(n1035), .B(n2500), .Z(n2498) );
  XOR U2502 ( .A(creg[560]), .B(mod_mult_o[560]), .Z(n2500) );
  XNOR U2503 ( .A(n2501), .B(n2502), .Z(o[55]) );
  AND U2504 ( .A(n1035), .B(n2503), .Z(n2501) );
  XOR U2505 ( .A(creg[55]), .B(mod_mult_o[55]), .Z(n2503) );
  XNOR U2506 ( .A(n2504), .B(n2505), .Z(o[559]) );
  AND U2507 ( .A(n1035), .B(n2506), .Z(n2504) );
  XOR U2508 ( .A(creg[559]), .B(mod_mult_o[559]), .Z(n2506) );
  XNOR U2509 ( .A(n2507), .B(n2508), .Z(o[558]) );
  AND U2510 ( .A(n1035), .B(n2509), .Z(n2507) );
  XOR U2511 ( .A(creg[558]), .B(mod_mult_o[558]), .Z(n2509) );
  XNOR U2512 ( .A(n2510), .B(n2511), .Z(o[557]) );
  AND U2513 ( .A(n1035), .B(n2512), .Z(n2510) );
  XOR U2514 ( .A(creg[557]), .B(mod_mult_o[557]), .Z(n2512) );
  XNOR U2515 ( .A(n2513), .B(n2514), .Z(o[556]) );
  AND U2516 ( .A(n1035), .B(n2515), .Z(n2513) );
  XOR U2517 ( .A(creg[556]), .B(mod_mult_o[556]), .Z(n2515) );
  XNOR U2518 ( .A(n2516), .B(n2517), .Z(o[555]) );
  AND U2519 ( .A(n1035), .B(n2518), .Z(n2516) );
  XOR U2520 ( .A(creg[555]), .B(mod_mult_o[555]), .Z(n2518) );
  XNOR U2521 ( .A(n2519), .B(n2520), .Z(o[554]) );
  AND U2522 ( .A(n1035), .B(n2521), .Z(n2519) );
  XOR U2523 ( .A(creg[554]), .B(mod_mult_o[554]), .Z(n2521) );
  XNOR U2524 ( .A(n2522), .B(n2523), .Z(o[553]) );
  AND U2525 ( .A(n1035), .B(n2524), .Z(n2522) );
  XOR U2526 ( .A(creg[553]), .B(mod_mult_o[553]), .Z(n2524) );
  XNOR U2527 ( .A(n2525), .B(n2526), .Z(o[552]) );
  AND U2528 ( .A(n1035), .B(n2527), .Z(n2525) );
  XOR U2529 ( .A(creg[552]), .B(mod_mult_o[552]), .Z(n2527) );
  XNOR U2530 ( .A(n2528), .B(n2529), .Z(o[551]) );
  AND U2531 ( .A(n1035), .B(n2530), .Z(n2528) );
  XOR U2532 ( .A(creg[551]), .B(mod_mult_o[551]), .Z(n2530) );
  XNOR U2533 ( .A(n2531), .B(n2532), .Z(o[550]) );
  AND U2534 ( .A(n1035), .B(n2533), .Z(n2531) );
  XOR U2535 ( .A(creg[550]), .B(mod_mult_o[550]), .Z(n2533) );
  XNOR U2536 ( .A(n2534), .B(n2535), .Z(o[54]) );
  AND U2537 ( .A(n1035), .B(n2536), .Z(n2534) );
  XOR U2538 ( .A(creg[54]), .B(mod_mult_o[54]), .Z(n2536) );
  XNOR U2539 ( .A(n2537), .B(n2538), .Z(o[549]) );
  AND U2540 ( .A(n1035), .B(n2539), .Z(n2537) );
  XOR U2541 ( .A(creg[549]), .B(mod_mult_o[549]), .Z(n2539) );
  XNOR U2542 ( .A(n2540), .B(n2541), .Z(o[548]) );
  AND U2543 ( .A(n1035), .B(n2542), .Z(n2540) );
  XOR U2544 ( .A(creg[548]), .B(mod_mult_o[548]), .Z(n2542) );
  XNOR U2545 ( .A(n2543), .B(n2544), .Z(o[547]) );
  AND U2546 ( .A(n1035), .B(n2545), .Z(n2543) );
  XOR U2547 ( .A(creg[547]), .B(mod_mult_o[547]), .Z(n2545) );
  XNOR U2548 ( .A(n2546), .B(n2547), .Z(o[546]) );
  AND U2549 ( .A(n1035), .B(n2548), .Z(n2546) );
  XOR U2550 ( .A(creg[546]), .B(mod_mult_o[546]), .Z(n2548) );
  XNOR U2551 ( .A(n2549), .B(n2550), .Z(o[545]) );
  AND U2552 ( .A(n1035), .B(n2551), .Z(n2549) );
  XOR U2553 ( .A(creg[545]), .B(mod_mult_o[545]), .Z(n2551) );
  XNOR U2554 ( .A(n2552), .B(n2553), .Z(o[544]) );
  AND U2555 ( .A(n1035), .B(n2554), .Z(n2552) );
  XOR U2556 ( .A(creg[544]), .B(mod_mult_o[544]), .Z(n2554) );
  XNOR U2557 ( .A(n2555), .B(n2556), .Z(o[543]) );
  AND U2558 ( .A(n1035), .B(n2557), .Z(n2555) );
  XOR U2559 ( .A(creg[543]), .B(mod_mult_o[543]), .Z(n2557) );
  XNOR U2560 ( .A(n2558), .B(n2559), .Z(o[542]) );
  AND U2561 ( .A(n1035), .B(n2560), .Z(n2558) );
  XOR U2562 ( .A(creg[542]), .B(mod_mult_o[542]), .Z(n2560) );
  XNOR U2563 ( .A(n2561), .B(n2562), .Z(o[541]) );
  AND U2564 ( .A(n1035), .B(n2563), .Z(n2561) );
  XOR U2565 ( .A(creg[541]), .B(mod_mult_o[541]), .Z(n2563) );
  XNOR U2566 ( .A(n2564), .B(n2565), .Z(o[540]) );
  AND U2567 ( .A(n1035), .B(n2566), .Z(n2564) );
  XOR U2568 ( .A(creg[540]), .B(mod_mult_o[540]), .Z(n2566) );
  XNOR U2569 ( .A(n2567), .B(n2568), .Z(o[53]) );
  AND U2570 ( .A(n1035), .B(n2569), .Z(n2567) );
  XOR U2571 ( .A(creg[53]), .B(mod_mult_o[53]), .Z(n2569) );
  XNOR U2572 ( .A(n2570), .B(n2571), .Z(o[539]) );
  AND U2573 ( .A(n1035), .B(n2572), .Z(n2570) );
  XOR U2574 ( .A(creg[539]), .B(mod_mult_o[539]), .Z(n2572) );
  XNOR U2575 ( .A(n2573), .B(n2574), .Z(o[538]) );
  AND U2576 ( .A(n1035), .B(n2575), .Z(n2573) );
  XOR U2577 ( .A(creg[538]), .B(mod_mult_o[538]), .Z(n2575) );
  XNOR U2578 ( .A(n2576), .B(n2577), .Z(o[537]) );
  AND U2579 ( .A(n1035), .B(n2578), .Z(n2576) );
  XOR U2580 ( .A(creg[537]), .B(mod_mult_o[537]), .Z(n2578) );
  XNOR U2581 ( .A(n2579), .B(n2580), .Z(o[536]) );
  AND U2582 ( .A(n1035), .B(n2581), .Z(n2579) );
  XOR U2583 ( .A(creg[536]), .B(mod_mult_o[536]), .Z(n2581) );
  XNOR U2584 ( .A(n2582), .B(n2583), .Z(o[535]) );
  AND U2585 ( .A(n1035), .B(n2584), .Z(n2582) );
  XOR U2586 ( .A(creg[535]), .B(mod_mult_o[535]), .Z(n2584) );
  XNOR U2587 ( .A(n2585), .B(n2586), .Z(o[534]) );
  AND U2588 ( .A(n1035), .B(n2587), .Z(n2585) );
  XOR U2589 ( .A(creg[534]), .B(mod_mult_o[534]), .Z(n2587) );
  XNOR U2590 ( .A(n2588), .B(n2589), .Z(o[533]) );
  AND U2591 ( .A(n1035), .B(n2590), .Z(n2588) );
  XOR U2592 ( .A(creg[533]), .B(mod_mult_o[533]), .Z(n2590) );
  XNOR U2593 ( .A(n2591), .B(n2592), .Z(o[532]) );
  AND U2594 ( .A(n1035), .B(n2593), .Z(n2591) );
  XOR U2595 ( .A(creg[532]), .B(mod_mult_o[532]), .Z(n2593) );
  XNOR U2596 ( .A(n2594), .B(n2595), .Z(o[531]) );
  AND U2597 ( .A(n1035), .B(n2596), .Z(n2594) );
  XOR U2598 ( .A(creg[531]), .B(mod_mult_o[531]), .Z(n2596) );
  XNOR U2599 ( .A(n2597), .B(n2598), .Z(o[530]) );
  AND U2600 ( .A(n1035), .B(n2599), .Z(n2597) );
  XOR U2601 ( .A(creg[530]), .B(mod_mult_o[530]), .Z(n2599) );
  XNOR U2602 ( .A(n2600), .B(n2601), .Z(o[52]) );
  AND U2603 ( .A(n1035), .B(n2602), .Z(n2600) );
  XOR U2604 ( .A(creg[52]), .B(mod_mult_o[52]), .Z(n2602) );
  XNOR U2605 ( .A(n2603), .B(n2604), .Z(o[529]) );
  AND U2606 ( .A(n1035), .B(n2605), .Z(n2603) );
  XOR U2607 ( .A(creg[529]), .B(mod_mult_o[529]), .Z(n2605) );
  XNOR U2608 ( .A(n2606), .B(n2607), .Z(o[528]) );
  AND U2609 ( .A(n1035), .B(n2608), .Z(n2606) );
  XOR U2610 ( .A(creg[528]), .B(mod_mult_o[528]), .Z(n2608) );
  XNOR U2611 ( .A(n2609), .B(n2610), .Z(o[527]) );
  AND U2612 ( .A(n1035), .B(n2611), .Z(n2609) );
  XOR U2613 ( .A(creg[527]), .B(mod_mult_o[527]), .Z(n2611) );
  XNOR U2614 ( .A(n2612), .B(n2613), .Z(o[526]) );
  AND U2615 ( .A(n1035), .B(n2614), .Z(n2612) );
  XOR U2616 ( .A(creg[526]), .B(mod_mult_o[526]), .Z(n2614) );
  XNOR U2617 ( .A(n2615), .B(n2616), .Z(o[525]) );
  AND U2618 ( .A(n1035), .B(n2617), .Z(n2615) );
  XOR U2619 ( .A(creg[525]), .B(mod_mult_o[525]), .Z(n2617) );
  XNOR U2620 ( .A(n2618), .B(n2619), .Z(o[524]) );
  AND U2621 ( .A(n1035), .B(n2620), .Z(n2618) );
  XOR U2622 ( .A(creg[524]), .B(mod_mult_o[524]), .Z(n2620) );
  XNOR U2623 ( .A(n2621), .B(n2622), .Z(o[523]) );
  AND U2624 ( .A(n1035), .B(n2623), .Z(n2621) );
  XOR U2625 ( .A(creg[523]), .B(mod_mult_o[523]), .Z(n2623) );
  XNOR U2626 ( .A(n2624), .B(n2625), .Z(o[522]) );
  AND U2627 ( .A(n1035), .B(n2626), .Z(n2624) );
  XOR U2628 ( .A(creg[522]), .B(mod_mult_o[522]), .Z(n2626) );
  XNOR U2629 ( .A(n2627), .B(n2628), .Z(o[521]) );
  AND U2630 ( .A(n1035), .B(n2629), .Z(n2627) );
  XOR U2631 ( .A(creg[521]), .B(mod_mult_o[521]), .Z(n2629) );
  XNOR U2632 ( .A(n2630), .B(n2631), .Z(o[520]) );
  AND U2633 ( .A(n1035), .B(n2632), .Z(n2630) );
  XOR U2634 ( .A(creg[520]), .B(mod_mult_o[520]), .Z(n2632) );
  XNOR U2635 ( .A(n2633), .B(n2634), .Z(o[51]) );
  AND U2636 ( .A(n1035), .B(n2635), .Z(n2633) );
  XOR U2637 ( .A(creg[51]), .B(mod_mult_o[51]), .Z(n2635) );
  XNOR U2638 ( .A(n2636), .B(n2637), .Z(o[519]) );
  AND U2639 ( .A(n1035), .B(n2638), .Z(n2636) );
  XOR U2640 ( .A(creg[519]), .B(mod_mult_o[519]), .Z(n2638) );
  XNOR U2641 ( .A(n2639), .B(n2640), .Z(o[518]) );
  AND U2642 ( .A(n1035), .B(n2641), .Z(n2639) );
  XOR U2643 ( .A(creg[518]), .B(mod_mult_o[518]), .Z(n2641) );
  XNOR U2644 ( .A(n2642), .B(n2643), .Z(o[517]) );
  AND U2645 ( .A(n1035), .B(n2644), .Z(n2642) );
  XOR U2646 ( .A(creg[517]), .B(mod_mult_o[517]), .Z(n2644) );
  XNOR U2647 ( .A(n2645), .B(n2646), .Z(o[516]) );
  AND U2648 ( .A(n1035), .B(n2647), .Z(n2645) );
  XOR U2649 ( .A(creg[516]), .B(mod_mult_o[516]), .Z(n2647) );
  XNOR U2650 ( .A(n2648), .B(n2649), .Z(o[515]) );
  AND U2651 ( .A(n1035), .B(n2650), .Z(n2648) );
  XOR U2652 ( .A(creg[515]), .B(mod_mult_o[515]), .Z(n2650) );
  XNOR U2653 ( .A(n2651), .B(n2652), .Z(o[514]) );
  AND U2654 ( .A(n1035), .B(n2653), .Z(n2651) );
  XOR U2655 ( .A(creg[514]), .B(mod_mult_o[514]), .Z(n2653) );
  XNOR U2656 ( .A(n2654), .B(n2655), .Z(o[513]) );
  AND U2657 ( .A(n1035), .B(n2656), .Z(n2654) );
  XOR U2658 ( .A(creg[513]), .B(mod_mult_o[513]), .Z(n2656) );
  XNOR U2659 ( .A(n2657), .B(n2658), .Z(o[512]) );
  AND U2660 ( .A(n1035), .B(n2659), .Z(n2657) );
  XOR U2661 ( .A(creg[512]), .B(mod_mult_o[512]), .Z(n2659) );
  XNOR U2662 ( .A(n2660), .B(n2661), .Z(o[511]) );
  AND U2663 ( .A(n1035), .B(n2662), .Z(n2660) );
  XOR U2664 ( .A(creg[511]), .B(mod_mult_o[511]), .Z(n2662) );
  XNOR U2665 ( .A(n2663), .B(n2664), .Z(o[510]) );
  AND U2666 ( .A(n1035), .B(n2665), .Z(n2663) );
  XOR U2667 ( .A(creg[510]), .B(mod_mult_o[510]), .Z(n2665) );
  XNOR U2668 ( .A(n2666), .B(n2667), .Z(o[50]) );
  AND U2669 ( .A(n1035), .B(n2668), .Z(n2666) );
  XOR U2670 ( .A(creg[50]), .B(mod_mult_o[50]), .Z(n2668) );
  XNOR U2671 ( .A(n2669), .B(n2670), .Z(o[509]) );
  AND U2672 ( .A(n1035), .B(n2671), .Z(n2669) );
  XOR U2673 ( .A(creg[509]), .B(mod_mult_o[509]), .Z(n2671) );
  XNOR U2674 ( .A(n2672), .B(n2673), .Z(o[508]) );
  AND U2675 ( .A(n1035), .B(n2674), .Z(n2672) );
  XOR U2676 ( .A(creg[508]), .B(mod_mult_o[508]), .Z(n2674) );
  XNOR U2677 ( .A(n2675), .B(n2676), .Z(o[507]) );
  AND U2678 ( .A(n1035), .B(n2677), .Z(n2675) );
  XOR U2679 ( .A(creg[507]), .B(mod_mult_o[507]), .Z(n2677) );
  XNOR U2680 ( .A(n2678), .B(n2679), .Z(o[506]) );
  AND U2681 ( .A(n1035), .B(n2680), .Z(n2678) );
  XOR U2682 ( .A(creg[506]), .B(mod_mult_o[506]), .Z(n2680) );
  XNOR U2683 ( .A(n2681), .B(n2682), .Z(o[505]) );
  AND U2684 ( .A(n1035), .B(n2683), .Z(n2681) );
  XOR U2685 ( .A(creg[505]), .B(mod_mult_o[505]), .Z(n2683) );
  XNOR U2686 ( .A(n2684), .B(n2685), .Z(o[504]) );
  AND U2687 ( .A(n1035), .B(n2686), .Z(n2684) );
  XOR U2688 ( .A(creg[504]), .B(mod_mult_o[504]), .Z(n2686) );
  XNOR U2689 ( .A(n2687), .B(n2688), .Z(o[503]) );
  AND U2690 ( .A(n1035), .B(n2689), .Z(n2687) );
  XOR U2691 ( .A(creg[503]), .B(mod_mult_o[503]), .Z(n2689) );
  XNOR U2692 ( .A(n2690), .B(n2691), .Z(o[502]) );
  AND U2693 ( .A(n1035), .B(n2692), .Z(n2690) );
  XOR U2694 ( .A(creg[502]), .B(mod_mult_o[502]), .Z(n2692) );
  XNOR U2695 ( .A(n2693), .B(n2694), .Z(o[501]) );
  AND U2696 ( .A(n1035), .B(n2695), .Z(n2693) );
  XOR U2697 ( .A(creg[501]), .B(mod_mult_o[501]), .Z(n2695) );
  XNOR U2698 ( .A(n2696), .B(n2697), .Z(o[500]) );
  AND U2699 ( .A(n1035), .B(n2698), .Z(n2696) );
  XOR U2700 ( .A(creg[500]), .B(mod_mult_o[500]), .Z(n2698) );
  XNOR U2701 ( .A(n2699), .B(n2700), .Z(o[4]) );
  AND U2702 ( .A(n1035), .B(n2701), .Z(n2699) );
  XOR U2703 ( .A(creg[4]), .B(mod_mult_o[4]), .Z(n2701) );
  XNOR U2704 ( .A(n2702), .B(n2703), .Z(o[49]) );
  AND U2705 ( .A(n1035), .B(n2704), .Z(n2702) );
  XOR U2706 ( .A(creg[49]), .B(mod_mult_o[49]), .Z(n2704) );
  XNOR U2707 ( .A(n2705), .B(n2706), .Z(o[499]) );
  AND U2708 ( .A(n1035), .B(n2707), .Z(n2705) );
  XOR U2709 ( .A(creg[499]), .B(mod_mult_o[499]), .Z(n2707) );
  XNOR U2710 ( .A(n2708), .B(n2709), .Z(o[498]) );
  AND U2711 ( .A(n1035), .B(n2710), .Z(n2708) );
  XOR U2712 ( .A(creg[498]), .B(mod_mult_o[498]), .Z(n2710) );
  XNOR U2713 ( .A(n2711), .B(n2712), .Z(o[497]) );
  AND U2714 ( .A(n1035), .B(n2713), .Z(n2711) );
  XOR U2715 ( .A(creg[497]), .B(mod_mult_o[497]), .Z(n2713) );
  XNOR U2716 ( .A(n2714), .B(n2715), .Z(o[496]) );
  AND U2717 ( .A(n1035), .B(n2716), .Z(n2714) );
  XOR U2718 ( .A(creg[496]), .B(mod_mult_o[496]), .Z(n2716) );
  XNOR U2719 ( .A(n2717), .B(n2718), .Z(o[495]) );
  AND U2720 ( .A(n1035), .B(n2719), .Z(n2717) );
  XOR U2721 ( .A(creg[495]), .B(mod_mult_o[495]), .Z(n2719) );
  XNOR U2722 ( .A(n2720), .B(n2721), .Z(o[494]) );
  AND U2723 ( .A(n1035), .B(n2722), .Z(n2720) );
  XOR U2724 ( .A(creg[494]), .B(mod_mult_o[494]), .Z(n2722) );
  XNOR U2725 ( .A(n2723), .B(n2724), .Z(o[493]) );
  AND U2726 ( .A(n1035), .B(n2725), .Z(n2723) );
  XOR U2727 ( .A(creg[493]), .B(mod_mult_o[493]), .Z(n2725) );
  XNOR U2728 ( .A(n2726), .B(n2727), .Z(o[492]) );
  AND U2729 ( .A(n1035), .B(n2728), .Z(n2726) );
  XOR U2730 ( .A(creg[492]), .B(mod_mult_o[492]), .Z(n2728) );
  XNOR U2731 ( .A(n2729), .B(n2730), .Z(o[491]) );
  AND U2732 ( .A(n1035), .B(n2731), .Z(n2729) );
  XOR U2733 ( .A(creg[491]), .B(mod_mult_o[491]), .Z(n2731) );
  XNOR U2734 ( .A(n2732), .B(n2733), .Z(o[490]) );
  AND U2735 ( .A(n1035), .B(n2734), .Z(n2732) );
  XOR U2736 ( .A(creg[490]), .B(mod_mult_o[490]), .Z(n2734) );
  XNOR U2737 ( .A(n2735), .B(n2736), .Z(o[48]) );
  AND U2738 ( .A(n1035), .B(n2737), .Z(n2735) );
  XOR U2739 ( .A(creg[48]), .B(mod_mult_o[48]), .Z(n2737) );
  XNOR U2740 ( .A(n2738), .B(n2739), .Z(o[489]) );
  AND U2741 ( .A(n1035), .B(n2740), .Z(n2738) );
  XOR U2742 ( .A(creg[489]), .B(mod_mult_o[489]), .Z(n2740) );
  XNOR U2743 ( .A(n2741), .B(n2742), .Z(o[488]) );
  AND U2744 ( .A(n1035), .B(n2743), .Z(n2741) );
  XOR U2745 ( .A(creg[488]), .B(mod_mult_o[488]), .Z(n2743) );
  XNOR U2746 ( .A(n2744), .B(n2745), .Z(o[487]) );
  AND U2747 ( .A(n1035), .B(n2746), .Z(n2744) );
  XOR U2748 ( .A(creg[487]), .B(mod_mult_o[487]), .Z(n2746) );
  XNOR U2749 ( .A(n2747), .B(n2748), .Z(o[486]) );
  AND U2750 ( .A(n1035), .B(n2749), .Z(n2747) );
  XOR U2751 ( .A(creg[486]), .B(mod_mult_o[486]), .Z(n2749) );
  XNOR U2752 ( .A(n2750), .B(n2751), .Z(o[485]) );
  AND U2753 ( .A(n1035), .B(n2752), .Z(n2750) );
  XOR U2754 ( .A(creg[485]), .B(mod_mult_o[485]), .Z(n2752) );
  XNOR U2755 ( .A(n2753), .B(n2754), .Z(o[484]) );
  AND U2756 ( .A(n1035), .B(n2755), .Z(n2753) );
  XOR U2757 ( .A(creg[484]), .B(mod_mult_o[484]), .Z(n2755) );
  XNOR U2758 ( .A(n2756), .B(n2757), .Z(o[483]) );
  AND U2759 ( .A(n1035), .B(n2758), .Z(n2756) );
  XOR U2760 ( .A(creg[483]), .B(mod_mult_o[483]), .Z(n2758) );
  XNOR U2761 ( .A(n2759), .B(n2760), .Z(o[482]) );
  AND U2762 ( .A(n1035), .B(n2761), .Z(n2759) );
  XOR U2763 ( .A(creg[482]), .B(mod_mult_o[482]), .Z(n2761) );
  XNOR U2764 ( .A(n2762), .B(n2763), .Z(o[481]) );
  AND U2765 ( .A(n1035), .B(n2764), .Z(n2762) );
  XOR U2766 ( .A(creg[481]), .B(mod_mult_o[481]), .Z(n2764) );
  XNOR U2767 ( .A(n2765), .B(n2766), .Z(o[480]) );
  AND U2768 ( .A(n1035), .B(n2767), .Z(n2765) );
  XOR U2769 ( .A(creg[480]), .B(mod_mult_o[480]), .Z(n2767) );
  XNOR U2770 ( .A(n2768), .B(n2769), .Z(o[47]) );
  AND U2771 ( .A(n1035), .B(n2770), .Z(n2768) );
  XOR U2772 ( .A(creg[47]), .B(mod_mult_o[47]), .Z(n2770) );
  XNOR U2773 ( .A(n2771), .B(n2772), .Z(o[479]) );
  AND U2774 ( .A(n1035), .B(n2773), .Z(n2771) );
  XOR U2775 ( .A(creg[479]), .B(mod_mult_o[479]), .Z(n2773) );
  XNOR U2776 ( .A(n2774), .B(n2775), .Z(o[478]) );
  AND U2777 ( .A(n1035), .B(n2776), .Z(n2774) );
  XOR U2778 ( .A(creg[478]), .B(mod_mult_o[478]), .Z(n2776) );
  XNOR U2779 ( .A(n2777), .B(n2778), .Z(o[477]) );
  AND U2780 ( .A(n1035), .B(n2779), .Z(n2777) );
  XOR U2781 ( .A(creg[477]), .B(mod_mult_o[477]), .Z(n2779) );
  XNOR U2782 ( .A(n2780), .B(n2781), .Z(o[476]) );
  AND U2783 ( .A(n1035), .B(n2782), .Z(n2780) );
  XOR U2784 ( .A(creg[476]), .B(mod_mult_o[476]), .Z(n2782) );
  XNOR U2785 ( .A(n2783), .B(n2784), .Z(o[475]) );
  AND U2786 ( .A(n1035), .B(n2785), .Z(n2783) );
  XOR U2787 ( .A(creg[475]), .B(mod_mult_o[475]), .Z(n2785) );
  XNOR U2788 ( .A(n2786), .B(n2787), .Z(o[474]) );
  AND U2789 ( .A(n1035), .B(n2788), .Z(n2786) );
  XOR U2790 ( .A(creg[474]), .B(mod_mult_o[474]), .Z(n2788) );
  XNOR U2791 ( .A(n2789), .B(n2790), .Z(o[473]) );
  AND U2792 ( .A(n1035), .B(n2791), .Z(n2789) );
  XOR U2793 ( .A(creg[473]), .B(mod_mult_o[473]), .Z(n2791) );
  XNOR U2794 ( .A(n2792), .B(n2793), .Z(o[472]) );
  AND U2795 ( .A(n1035), .B(n2794), .Z(n2792) );
  XOR U2796 ( .A(creg[472]), .B(mod_mult_o[472]), .Z(n2794) );
  XNOR U2797 ( .A(n2795), .B(n2796), .Z(o[471]) );
  AND U2798 ( .A(n1035), .B(n2797), .Z(n2795) );
  XOR U2799 ( .A(creg[471]), .B(mod_mult_o[471]), .Z(n2797) );
  XNOR U2800 ( .A(n2798), .B(n2799), .Z(o[470]) );
  AND U2801 ( .A(n1035), .B(n2800), .Z(n2798) );
  XOR U2802 ( .A(creg[470]), .B(mod_mult_o[470]), .Z(n2800) );
  XNOR U2803 ( .A(n2801), .B(n2802), .Z(o[46]) );
  AND U2804 ( .A(n1035), .B(n2803), .Z(n2801) );
  XOR U2805 ( .A(creg[46]), .B(mod_mult_o[46]), .Z(n2803) );
  XNOR U2806 ( .A(n2804), .B(n2805), .Z(o[469]) );
  AND U2807 ( .A(n1035), .B(n2806), .Z(n2804) );
  XOR U2808 ( .A(creg[469]), .B(mod_mult_o[469]), .Z(n2806) );
  XNOR U2809 ( .A(n2807), .B(n2808), .Z(o[468]) );
  AND U2810 ( .A(n1035), .B(n2809), .Z(n2807) );
  XOR U2811 ( .A(creg[468]), .B(mod_mult_o[468]), .Z(n2809) );
  XNOR U2812 ( .A(n2810), .B(n2811), .Z(o[467]) );
  AND U2813 ( .A(n1035), .B(n2812), .Z(n2810) );
  XOR U2814 ( .A(creg[467]), .B(mod_mult_o[467]), .Z(n2812) );
  XNOR U2815 ( .A(n2813), .B(n2814), .Z(o[466]) );
  AND U2816 ( .A(n1035), .B(n2815), .Z(n2813) );
  XOR U2817 ( .A(creg[466]), .B(mod_mult_o[466]), .Z(n2815) );
  XNOR U2818 ( .A(n2816), .B(n2817), .Z(o[465]) );
  AND U2819 ( .A(n1035), .B(n2818), .Z(n2816) );
  XOR U2820 ( .A(creg[465]), .B(mod_mult_o[465]), .Z(n2818) );
  XNOR U2821 ( .A(n2819), .B(n2820), .Z(o[464]) );
  AND U2822 ( .A(n1035), .B(n2821), .Z(n2819) );
  XOR U2823 ( .A(creg[464]), .B(mod_mult_o[464]), .Z(n2821) );
  XNOR U2824 ( .A(n2822), .B(n2823), .Z(o[463]) );
  AND U2825 ( .A(n1035), .B(n2824), .Z(n2822) );
  XOR U2826 ( .A(creg[463]), .B(mod_mult_o[463]), .Z(n2824) );
  XNOR U2827 ( .A(n2825), .B(n2826), .Z(o[462]) );
  AND U2828 ( .A(n1035), .B(n2827), .Z(n2825) );
  XOR U2829 ( .A(creg[462]), .B(mod_mult_o[462]), .Z(n2827) );
  XNOR U2830 ( .A(n2828), .B(n2829), .Z(o[461]) );
  AND U2831 ( .A(n1035), .B(n2830), .Z(n2828) );
  XOR U2832 ( .A(creg[461]), .B(mod_mult_o[461]), .Z(n2830) );
  XNOR U2833 ( .A(n2831), .B(n2832), .Z(o[460]) );
  AND U2834 ( .A(n1035), .B(n2833), .Z(n2831) );
  XOR U2835 ( .A(creg[460]), .B(mod_mult_o[460]), .Z(n2833) );
  XNOR U2836 ( .A(n2834), .B(n2835), .Z(o[45]) );
  AND U2837 ( .A(n1035), .B(n2836), .Z(n2834) );
  XOR U2838 ( .A(creg[45]), .B(mod_mult_o[45]), .Z(n2836) );
  XNOR U2839 ( .A(n2837), .B(n2838), .Z(o[459]) );
  AND U2840 ( .A(n1035), .B(n2839), .Z(n2837) );
  XOR U2841 ( .A(creg[459]), .B(mod_mult_o[459]), .Z(n2839) );
  XNOR U2842 ( .A(n2840), .B(n2841), .Z(o[458]) );
  AND U2843 ( .A(n1035), .B(n2842), .Z(n2840) );
  XOR U2844 ( .A(creg[458]), .B(mod_mult_o[458]), .Z(n2842) );
  XNOR U2845 ( .A(n2843), .B(n2844), .Z(o[457]) );
  AND U2846 ( .A(n1035), .B(n2845), .Z(n2843) );
  XOR U2847 ( .A(creg[457]), .B(mod_mult_o[457]), .Z(n2845) );
  XNOR U2848 ( .A(n2846), .B(n2847), .Z(o[456]) );
  AND U2849 ( .A(n1035), .B(n2848), .Z(n2846) );
  XOR U2850 ( .A(creg[456]), .B(mod_mult_o[456]), .Z(n2848) );
  XNOR U2851 ( .A(n2849), .B(n2850), .Z(o[455]) );
  AND U2852 ( .A(n1035), .B(n2851), .Z(n2849) );
  XOR U2853 ( .A(creg[455]), .B(mod_mult_o[455]), .Z(n2851) );
  XNOR U2854 ( .A(n2852), .B(n2853), .Z(o[454]) );
  AND U2855 ( .A(n1035), .B(n2854), .Z(n2852) );
  XOR U2856 ( .A(creg[454]), .B(mod_mult_o[454]), .Z(n2854) );
  XNOR U2857 ( .A(n2855), .B(n2856), .Z(o[453]) );
  AND U2858 ( .A(n1035), .B(n2857), .Z(n2855) );
  XOR U2859 ( .A(creg[453]), .B(mod_mult_o[453]), .Z(n2857) );
  XNOR U2860 ( .A(n2858), .B(n2859), .Z(o[452]) );
  AND U2861 ( .A(n1035), .B(n2860), .Z(n2858) );
  XOR U2862 ( .A(creg[452]), .B(mod_mult_o[452]), .Z(n2860) );
  XNOR U2863 ( .A(n2861), .B(n2862), .Z(o[451]) );
  AND U2864 ( .A(n1035), .B(n2863), .Z(n2861) );
  XOR U2865 ( .A(creg[451]), .B(mod_mult_o[451]), .Z(n2863) );
  XNOR U2866 ( .A(n2864), .B(n2865), .Z(o[450]) );
  AND U2867 ( .A(n1035), .B(n2866), .Z(n2864) );
  XOR U2868 ( .A(creg[450]), .B(mod_mult_o[450]), .Z(n2866) );
  XNOR U2869 ( .A(n2867), .B(n2868), .Z(o[44]) );
  AND U2870 ( .A(n1035), .B(n2869), .Z(n2867) );
  XOR U2871 ( .A(creg[44]), .B(mod_mult_o[44]), .Z(n2869) );
  XNOR U2872 ( .A(n2870), .B(n2871), .Z(o[449]) );
  AND U2873 ( .A(n1035), .B(n2872), .Z(n2870) );
  XOR U2874 ( .A(creg[449]), .B(mod_mult_o[449]), .Z(n2872) );
  XNOR U2875 ( .A(n2873), .B(n2874), .Z(o[448]) );
  AND U2876 ( .A(n1035), .B(n2875), .Z(n2873) );
  XOR U2877 ( .A(creg[448]), .B(mod_mult_o[448]), .Z(n2875) );
  XNOR U2878 ( .A(n2876), .B(n2877), .Z(o[447]) );
  AND U2879 ( .A(n1035), .B(n2878), .Z(n2876) );
  XOR U2880 ( .A(creg[447]), .B(mod_mult_o[447]), .Z(n2878) );
  XNOR U2881 ( .A(n2879), .B(n2880), .Z(o[446]) );
  AND U2882 ( .A(n1035), .B(n2881), .Z(n2879) );
  XOR U2883 ( .A(creg[446]), .B(mod_mult_o[446]), .Z(n2881) );
  XNOR U2884 ( .A(n2882), .B(n2883), .Z(o[445]) );
  AND U2885 ( .A(n1035), .B(n2884), .Z(n2882) );
  XOR U2886 ( .A(creg[445]), .B(mod_mult_o[445]), .Z(n2884) );
  XNOR U2887 ( .A(n2885), .B(n2886), .Z(o[444]) );
  AND U2888 ( .A(n1035), .B(n2887), .Z(n2885) );
  XOR U2889 ( .A(creg[444]), .B(mod_mult_o[444]), .Z(n2887) );
  XNOR U2890 ( .A(n2888), .B(n2889), .Z(o[443]) );
  AND U2891 ( .A(n1035), .B(n2890), .Z(n2888) );
  XOR U2892 ( .A(creg[443]), .B(mod_mult_o[443]), .Z(n2890) );
  XNOR U2893 ( .A(n2891), .B(n2892), .Z(o[442]) );
  AND U2894 ( .A(n1035), .B(n2893), .Z(n2891) );
  XOR U2895 ( .A(creg[442]), .B(mod_mult_o[442]), .Z(n2893) );
  XNOR U2896 ( .A(n2894), .B(n2895), .Z(o[441]) );
  AND U2897 ( .A(n1035), .B(n2896), .Z(n2894) );
  XOR U2898 ( .A(creg[441]), .B(mod_mult_o[441]), .Z(n2896) );
  XNOR U2899 ( .A(n2897), .B(n2898), .Z(o[440]) );
  AND U2900 ( .A(n1035), .B(n2899), .Z(n2897) );
  XOR U2901 ( .A(creg[440]), .B(mod_mult_o[440]), .Z(n2899) );
  XNOR U2902 ( .A(n2900), .B(n2901), .Z(o[43]) );
  AND U2903 ( .A(n1035), .B(n2902), .Z(n2900) );
  XOR U2904 ( .A(creg[43]), .B(mod_mult_o[43]), .Z(n2902) );
  XNOR U2905 ( .A(n2903), .B(n2904), .Z(o[439]) );
  AND U2906 ( .A(n1035), .B(n2905), .Z(n2903) );
  XOR U2907 ( .A(creg[439]), .B(mod_mult_o[439]), .Z(n2905) );
  XNOR U2908 ( .A(n2906), .B(n2907), .Z(o[438]) );
  AND U2909 ( .A(n1035), .B(n2908), .Z(n2906) );
  XOR U2910 ( .A(creg[438]), .B(mod_mult_o[438]), .Z(n2908) );
  XNOR U2911 ( .A(n2909), .B(n2910), .Z(o[437]) );
  AND U2912 ( .A(n1035), .B(n2911), .Z(n2909) );
  XOR U2913 ( .A(creg[437]), .B(mod_mult_o[437]), .Z(n2911) );
  XNOR U2914 ( .A(n2912), .B(n2913), .Z(o[436]) );
  AND U2915 ( .A(n1035), .B(n2914), .Z(n2912) );
  XOR U2916 ( .A(creg[436]), .B(mod_mult_o[436]), .Z(n2914) );
  XNOR U2917 ( .A(n2915), .B(n2916), .Z(o[435]) );
  AND U2918 ( .A(n1035), .B(n2917), .Z(n2915) );
  XOR U2919 ( .A(creg[435]), .B(mod_mult_o[435]), .Z(n2917) );
  XNOR U2920 ( .A(n2918), .B(n2919), .Z(o[434]) );
  AND U2921 ( .A(n1035), .B(n2920), .Z(n2918) );
  XOR U2922 ( .A(creg[434]), .B(mod_mult_o[434]), .Z(n2920) );
  XNOR U2923 ( .A(n2921), .B(n2922), .Z(o[433]) );
  AND U2924 ( .A(n1035), .B(n2923), .Z(n2921) );
  XOR U2925 ( .A(creg[433]), .B(mod_mult_o[433]), .Z(n2923) );
  XNOR U2926 ( .A(n2924), .B(n2925), .Z(o[432]) );
  AND U2927 ( .A(n1035), .B(n2926), .Z(n2924) );
  XOR U2928 ( .A(creg[432]), .B(mod_mult_o[432]), .Z(n2926) );
  XNOR U2929 ( .A(n2927), .B(n2928), .Z(o[431]) );
  AND U2930 ( .A(n1035), .B(n2929), .Z(n2927) );
  XOR U2931 ( .A(creg[431]), .B(mod_mult_o[431]), .Z(n2929) );
  XNOR U2932 ( .A(n2930), .B(n2931), .Z(o[430]) );
  AND U2933 ( .A(n1035), .B(n2932), .Z(n2930) );
  XOR U2934 ( .A(creg[430]), .B(mod_mult_o[430]), .Z(n2932) );
  XNOR U2935 ( .A(n2933), .B(n2934), .Z(o[42]) );
  AND U2936 ( .A(n1035), .B(n2935), .Z(n2933) );
  XOR U2937 ( .A(creg[42]), .B(mod_mult_o[42]), .Z(n2935) );
  XNOR U2938 ( .A(n2936), .B(n2937), .Z(o[429]) );
  AND U2939 ( .A(n1035), .B(n2938), .Z(n2936) );
  XOR U2940 ( .A(creg[429]), .B(mod_mult_o[429]), .Z(n2938) );
  XNOR U2941 ( .A(n2939), .B(n2940), .Z(o[428]) );
  AND U2942 ( .A(n1035), .B(n2941), .Z(n2939) );
  XOR U2943 ( .A(creg[428]), .B(mod_mult_o[428]), .Z(n2941) );
  XNOR U2944 ( .A(n2942), .B(n2943), .Z(o[427]) );
  AND U2945 ( .A(n1035), .B(n2944), .Z(n2942) );
  XOR U2946 ( .A(creg[427]), .B(mod_mult_o[427]), .Z(n2944) );
  XNOR U2947 ( .A(n2945), .B(n2946), .Z(o[426]) );
  AND U2948 ( .A(n1035), .B(n2947), .Z(n2945) );
  XOR U2949 ( .A(creg[426]), .B(mod_mult_o[426]), .Z(n2947) );
  XNOR U2950 ( .A(n2948), .B(n2949), .Z(o[425]) );
  AND U2951 ( .A(n1035), .B(n2950), .Z(n2948) );
  XOR U2952 ( .A(creg[425]), .B(mod_mult_o[425]), .Z(n2950) );
  XNOR U2953 ( .A(n2951), .B(n2952), .Z(o[424]) );
  AND U2954 ( .A(n1035), .B(n2953), .Z(n2951) );
  XOR U2955 ( .A(creg[424]), .B(mod_mult_o[424]), .Z(n2953) );
  XNOR U2956 ( .A(n2954), .B(n2955), .Z(o[423]) );
  AND U2957 ( .A(n1035), .B(n2956), .Z(n2954) );
  XOR U2958 ( .A(creg[423]), .B(mod_mult_o[423]), .Z(n2956) );
  XNOR U2959 ( .A(n2957), .B(n2958), .Z(o[422]) );
  AND U2960 ( .A(n1035), .B(n2959), .Z(n2957) );
  XOR U2961 ( .A(creg[422]), .B(mod_mult_o[422]), .Z(n2959) );
  XNOR U2962 ( .A(n2960), .B(n2961), .Z(o[421]) );
  AND U2963 ( .A(n1035), .B(n2962), .Z(n2960) );
  XOR U2964 ( .A(creg[421]), .B(mod_mult_o[421]), .Z(n2962) );
  XNOR U2965 ( .A(n2963), .B(n2964), .Z(o[420]) );
  AND U2966 ( .A(n1035), .B(n2965), .Z(n2963) );
  XOR U2967 ( .A(creg[420]), .B(mod_mult_o[420]), .Z(n2965) );
  XNOR U2968 ( .A(n2966), .B(n2967), .Z(o[41]) );
  AND U2969 ( .A(n1035), .B(n2968), .Z(n2966) );
  XOR U2970 ( .A(creg[41]), .B(mod_mult_o[41]), .Z(n2968) );
  XNOR U2971 ( .A(n2969), .B(n2970), .Z(o[419]) );
  AND U2972 ( .A(n1035), .B(n2971), .Z(n2969) );
  XOR U2973 ( .A(creg[419]), .B(mod_mult_o[419]), .Z(n2971) );
  XNOR U2974 ( .A(n2972), .B(n2973), .Z(o[418]) );
  AND U2975 ( .A(n1035), .B(n2974), .Z(n2972) );
  XOR U2976 ( .A(creg[418]), .B(mod_mult_o[418]), .Z(n2974) );
  XNOR U2977 ( .A(n2975), .B(n2976), .Z(o[417]) );
  AND U2978 ( .A(n1035), .B(n2977), .Z(n2975) );
  XOR U2979 ( .A(creg[417]), .B(mod_mult_o[417]), .Z(n2977) );
  XNOR U2980 ( .A(n2978), .B(n2979), .Z(o[416]) );
  AND U2981 ( .A(n1035), .B(n2980), .Z(n2978) );
  XOR U2982 ( .A(creg[416]), .B(mod_mult_o[416]), .Z(n2980) );
  XNOR U2983 ( .A(n2981), .B(n2982), .Z(o[415]) );
  AND U2984 ( .A(n1035), .B(n2983), .Z(n2981) );
  XOR U2985 ( .A(creg[415]), .B(mod_mult_o[415]), .Z(n2983) );
  XNOR U2986 ( .A(n2984), .B(n2985), .Z(o[414]) );
  AND U2987 ( .A(n1035), .B(n2986), .Z(n2984) );
  XOR U2988 ( .A(creg[414]), .B(mod_mult_o[414]), .Z(n2986) );
  XNOR U2989 ( .A(n2987), .B(n2988), .Z(o[413]) );
  AND U2990 ( .A(n1035), .B(n2989), .Z(n2987) );
  XOR U2991 ( .A(creg[413]), .B(mod_mult_o[413]), .Z(n2989) );
  XNOR U2992 ( .A(n2990), .B(n2991), .Z(o[412]) );
  AND U2993 ( .A(n1035), .B(n2992), .Z(n2990) );
  XOR U2994 ( .A(creg[412]), .B(mod_mult_o[412]), .Z(n2992) );
  XNOR U2995 ( .A(n2993), .B(n2994), .Z(o[411]) );
  AND U2996 ( .A(n1035), .B(n2995), .Z(n2993) );
  XOR U2997 ( .A(creg[411]), .B(mod_mult_o[411]), .Z(n2995) );
  XNOR U2998 ( .A(n2996), .B(n2997), .Z(o[410]) );
  AND U2999 ( .A(n1035), .B(n2998), .Z(n2996) );
  XOR U3000 ( .A(creg[410]), .B(mod_mult_o[410]), .Z(n2998) );
  XNOR U3001 ( .A(n2999), .B(n3000), .Z(o[40]) );
  AND U3002 ( .A(n1035), .B(n3001), .Z(n2999) );
  XOR U3003 ( .A(creg[40]), .B(mod_mult_o[40]), .Z(n3001) );
  XNOR U3004 ( .A(n3002), .B(n3003), .Z(o[409]) );
  AND U3005 ( .A(n1035), .B(n3004), .Z(n3002) );
  XOR U3006 ( .A(creg[409]), .B(mod_mult_o[409]), .Z(n3004) );
  XNOR U3007 ( .A(n3005), .B(n3006), .Z(o[408]) );
  AND U3008 ( .A(n1035), .B(n3007), .Z(n3005) );
  XOR U3009 ( .A(creg[408]), .B(mod_mult_o[408]), .Z(n3007) );
  XNOR U3010 ( .A(n3008), .B(n3009), .Z(o[407]) );
  AND U3011 ( .A(n1035), .B(n3010), .Z(n3008) );
  XOR U3012 ( .A(creg[407]), .B(mod_mult_o[407]), .Z(n3010) );
  XNOR U3013 ( .A(n3011), .B(n3012), .Z(o[406]) );
  AND U3014 ( .A(n1035), .B(n3013), .Z(n3011) );
  XOR U3015 ( .A(creg[406]), .B(mod_mult_o[406]), .Z(n3013) );
  XNOR U3016 ( .A(n3014), .B(n3015), .Z(o[405]) );
  AND U3017 ( .A(n1035), .B(n3016), .Z(n3014) );
  XOR U3018 ( .A(creg[405]), .B(mod_mult_o[405]), .Z(n3016) );
  XNOR U3019 ( .A(n3017), .B(n3018), .Z(o[404]) );
  AND U3020 ( .A(n1035), .B(n3019), .Z(n3017) );
  XOR U3021 ( .A(creg[404]), .B(mod_mult_o[404]), .Z(n3019) );
  XNOR U3022 ( .A(n3020), .B(n3021), .Z(o[403]) );
  AND U3023 ( .A(n1035), .B(n3022), .Z(n3020) );
  XOR U3024 ( .A(creg[403]), .B(mod_mult_o[403]), .Z(n3022) );
  XNOR U3025 ( .A(n3023), .B(n3024), .Z(o[402]) );
  AND U3026 ( .A(n1035), .B(n3025), .Z(n3023) );
  XOR U3027 ( .A(creg[402]), .B(mod_mult_o[402]), .Z(n3025) );
  XNOR U3028 ( .A(n3026), .B(n3027), .Z(o[401]) );
  AND U3029 ( .A(n1035), .B(n3028), .Z(n3026) );
  XOR U3030 ( .A(creg[401]), .B(mod_mult_o[401]), .Z(n3028) );
  XNOR U3031 ( .A(n3029), .B(n3030), .Z(o[400]) );
  AND U3032 ( .A(n1035), .B(n3031), .Z(n3029) );
  XOR U3033 ( .A(creg[400]), .B(mod_mult_o[400]), .Z(n3031) );
  XNOR U3034 ( .A(n3032), .B(n3033), .Z(o[3]) );
  AND U3035 ( .A(n1035), .B(n3034), .Z(n3032) );
  XOR U3036 ( .A(creg[3]), .B(mod_mult_o[3]), .Z(n3034) );
  XNOR U3037 ( .A(n3035), .B(n3036), .Z(o[39]) );
  AND U3038 ( .A(n1035), .B(n3037), .Z(n3035) );
  XOR U3039 ( .A(creg[39]), .B(mod_mult_o[39]), .Z(n3037) );
  XNOR U3040 ( .A(n3038), .B(n3039), .Z(o[399]) );
  AND U3041 ( .A(n1035), .B(n3040), .Z(n3038) );
  XOR U3042 ( .A(creg[399]), .B(mod_mult_o[399]), .Z(n3040) );
  XNOR U3043 ( .A(n3041), .B(n3042), .Z(o[398]) );
  AND U3044 ( .A(n1035), .B(n3043), .Z(n3041) );
  XOR U3045 ( .A(creg[398]), .B(mod_mult_o[398]), .Z(n3043) );
  XNOR U3046 ( .A(n3044), .B(n3045), .Z(o[397]) );
  AND U3047 ( .A(n1035), .B(n3046), .Z(n3044) );
  XOR U3048 ( .A(creg[397]), .B(mod_mult_o[397]), .Z(n3046) );
  XNOR U3049 ( .A(n3047), .B(n3048), .Z(o[396]) );
  AND U3050 ( .A(n1035), .B(n3049), .Z(n3047) );
  XOR U3051 ( .A(creg[396]), .B(mod_mult_o[396]), .Z(n3049) );
  XNOR U3052 ( .A(n3050), .B(n3051), .Z(o[395]) );
  AND U3053 ( .A(n1035), .B(n3052), .Z(n3050) );
  XOR U3054 ( .A(creg[395]), .B(mod_mult_o[395]), .Z(n3052) );
  XNOR U3055 ( .A(n3053), .B(n3054), .Z(o[394]) );
  AND U3056 ( .A(n1035), .B(n3055), .Z(n3053) );
  XOR U3057 ( .A(creg[394]), .B(mod_mult_o[394]), .Z(n3055) );
  XNOR U3058 ( .A(n3056), .B(n3057), .Z(o[393]) );
  AND U3059 ( .A(n1035), .B(n3058), .Z(n3056) );
  XOR U3060 ( .A(creg[393]), .B(mod_mult_o[393]), .Z(n3058) );
  XNOR U3061 ( .A(n3059), .B(n3060), .Z(o[392]) );
  AND U3062 ( .A(n1035), .B(n3061), .Z(n3059) );
  XOR U3063 ( .A(creg[392]), .B(mod_mult_o[392]), .Z(n3061) );
  XNOR U3064 ( .A(n3062), .B(n3063), .Z(o[391]) );
  AND U3065 ( .A(n1035), .B(n3064), .Z(n3062) );
  XOR U3066 ( .A(creg[391]), .B(mod_mult_o[391]), .Z(n3064) );
  XNOR U3067 ( .A(n3065), .B(n3066), .Z(o[390]) );
  AND U3068 ( .A(n1035), .B(n3067), .Z(n3065) );
  XOR U3069 ( .A(creg[390]), .B(mod_mult_o[390]), .Z(n3067) );
  XNOR U3070 ( .A(n3068), .B(n3069), .Z(o[38]) );
  AND U3071 ( .A(n1035), .B(n3070), .Z(n3068) );
  XOR U3072 ( .A(creg[38]), .B(mod_mult_o[38]), .Z(n3070) );
  XNOR U3073 ( .A(n3071), .B(n3072), .Z(o[389]) );
  AND U3074 ( .A(n1035), .B(n3073), .Z(n3071) );
  XOR U3075 ( .A(creg[389]), .B(mod_mult_o[389]), .Z(n3073) );
  XNOR U3076 ( .A(n3074), .B(n3075), .Z(o[388]) );
  AND U3077 ( .A(n1035), .B(n3076), .Z(n3074) );
  XOR U3078 ( .A(creg[388]), .B(mod_mult_o[388]), .Z(n3076) );
  XNOR U3079 ( .A(n3077), .B(n3078), .Z(o[387]) );
  AND U3080 ( .A(n1035), .B(n3079), .Z(n3077) );
  XOR U3081 ( .A(creg[387]), .B(mod_mult_o[387]), .Z(n3079) );
  XNOR U3082 ( .A(n3080), .B(n3081), .Z(o[386]) );
  AND U3083 ( .A(n1035), .B(n3082), .Z(n3080) );
  XOR U3084 ( .A(creg[386]), .B(mod_mult_o[386]), .Z(n3082) );
  XNOR U3085 ( .A(n3083), .B(n3084), .Z(o[385]) );
  AND U3086 ( .A(n1035), .B(n3085), .Z(n3083) );
  XOR U3087 ( .A(creg[385]), .B(mod_mult_o[385]), .Z(n3085) );
  XNOR U3088 ( .A(n3086), .B(n3087), .Z(o[384]) );
  AND U3089 ( .A(n1035), .B(n3088), .Z(n3086) );
  XOR U3090 ( .A(creg[384]), .B(mod_mult_o[384]), .Z(n3088) );
  XNOR U3091 ( .A(n3089), .B(n3090), .Z(o[383]) );
  AND U3092 ( .A(n1035), .B(n3091), .Z(n3089) );
  XOR U3093 ( .A(creg[383]), .B(mod_mult_o[383]), .Z(n3091) );
  XNOR U3094 ( .A(n3092), .B(n3093), .Z(o[382]) );
  AND U3095 ( .A(n1035), .B(n3094), .Z(n3092) );
  XOR U3096 ( .A(creg[382]), .B(mod_mult_o[382]), .Z(n3094) );
  XNOR U3097 ( .A(n3095), .B(n3096), .Z(o[381]) );
  AND U3098 ( .A(n1035), .B(n3097), .Z(n3095) );
  XOR U3099 ( .A(creg[381]), .B(mod_mult_o[381]), .Z(n3097) );
  XNOR U3100 ( .A(n3098), .B(n3099), .Z(o[380]) );
  AND U3101 ( .A(n1035), .B(n3100), .Z(n3098) );
  XOR U3102 ( .A(creg[380]), .B(mod_mult_o[380]), .Z(n3100) );
  XNOR U3103 ( .A(n3101), .B(n3102), .Z(o[37]) );
  AND U3104 ( .A(n1035), .B(n3103), .Z(n3101) );
  XOR U3105 ( .A(creg[37]), .B(mod_mult_o[37]), .Z(n3103) );
  XNOR U3106 ( .A(n3104), .B(n3105), .Z(o[379]) );
  AND U3107 ( .A(n1035), .B(n3106), .Z(n3104) );
  XOR U3108 ( .A(creg[379]), .B(mod_mult_o[379]), .Z(n3106) );
  XNOR U3109 ( .A(n3107), .B(n3108), .Z(o[378]) );
  AND U3110 ( .A(n1035), .B(n3109), .Z(n3107) );
  XOR U3111 ( .A(creg[378]), .B(mod_mult_o[378]), .Z(n3109) );
  XNOR U3112 ( .A(n3110), .B(n3111), .Z(o[377]) );
  AND U3113 ( .A(n1035), .B(n3112), .Z(n3110) );
  XOR U3114 ( .A(creg[377]), .B(mod_mult_o[377]), .Z(n3112) );
  XNOR U3115 ( .A(n3113), .B(n3114), .Z(o[376]) );
  AND U3116 ( .A(n1035), .B(n3115), .Z(n3113) );
  XOR U3117 ( .A(creg[376]), .B(mod_mult_o[376]), .Z(n3115) );
  XNOR U3118 ( .A(n3116), .B(n3117), .Z(o[375]) );
  AND U3119 ( .A(n1035), .B(n3118), .Z(n3116) );
  XOR U3120 ( .A(creg[375]), .B(mod_mult_o[375]), .Z(n3118) );
  XNOR U3121 ( .A(n3119), .B(n3120), .Z(o[374]) );
  AND U3122 ( .A(n1035), .B(n3121), .Z(n3119) );
  XOR U3123 ( .A(creg[374]), .B(mod_mult_o[374]), .Z(n3121) );
  XNOR U3124 ( .A(n3122), .B(n3123), .Z(o[373]) );
  AND U3125 ( .A(n1035), .B(n3124), .Z(n3122) );
  XOR U3126 ( .A(creg[373]), .B(mod_mult_o[373]), .Z(n3124) );
  XNOR U3127 ( .A(n3125), .B(n3126), .Z(o[372]) );
  AND U3128 ( .A(n1035), .B(n3127), .Z(n3125) );
  XOR U3129 ( .A(creg[372]), .B(mod_mult_o[372]), .Z(n3127) );
  XNOR U3130 ( .A(n3128), .B(n3129), .Z(o[371]) );
  AND U3131 ( .A(n1035), .B(n3130), .Z(n3128) );
  XOR U3132 ( .A(creg[371]), .B(mod_mult_o[371]), .Z(n3130) );
  XNOR U3133 ( .A(n3131), .B(n3132), .Z(o[370]) );
  AND U3134 ( .A(n1035), .B(n3133), .Z(n3131) );
  XOR U3135 ( .A(creg[370]), .B(mod_mult_o[370]), .Z(n3133) );
  XNOR U3136 ( .A(n3134), .B(n3135), .Z(o[36]) );
  AND U3137 ( .A(n1035), .B(n3136), .Z(n3134) );
  XOR U3138 ( .A(creg[36]), .B(mod_mult_o[36]), .Z(n3136) );
  XNOR U3139 ( .A(n3137), .B(n3138), .Z(o[369]) );
  AND U3140 ( .A(n1035), .B(n3139), .Z(n3137) );
  XOR U3141 ( .A(creg[369]), .B(mod_mult_o[369]), .Z(n3139) );
  XNOR U3142 ( .A(n3140), .B(n3141), .Z(o[368]) );
  AND U3143 ( .A(n1035), .B(n3142), .Z(n3140) );
  XOR U3144 ( .A(creg[368]), .B(mod_mult_o[368]), .Z(n3142) );
  XNOR U3145 ( .A(n3143), .B(n3144), .Z(o[367]) );
  AND U3146 ( .A(n1035), .B(n3145), .Z(n3143) );
  XOR U3147 ( .A(creg[367]), .B(mod_mult_o[367]), .Z(n3145) );
  XNOR U3148 ( .A(n3146), .B(n3147), .Z(o[366]) );
  AND U3149 ( .A(n1035), .B(n3148), .Z(n3146) );
  XOR U3150 ( .A(creg[366]), .B(mod_mult_o[366]), .Z(n3148) );
  XNOR U3151 ( .A(n3149), .B(n3150), .Z(o[365]) );
  AND U3152 ( .A(n1035), .B(n3151), .Z(n3149) );
  XOR U3153 ( .A(creg[365]), .B(mod_mult_o[365]), .Z(n3151) );
  XNOR U3154 ( .A(n3152), .B(n3153), .Z(o[364]) );
  AND U3155 ( .A(n1035), .B(n3154), .Z(n3152) );
  XOR U3156 ( .A(creg[364]), .B(mod_mult_o[364]), .Z(n3154) );
  XNOR U3157 ( .A(n3155), .B(n3156), .Z(o[363]) );
  AND U3158 ( .A(n1035), .B(n3157), .Z(n3155) );
  XOR U3159 ( .A(creg[363]), .B(mod_mult_o[363]), .Z(n3157) );
  XNOR U3160 ( .A(n3158), .B(n3159), .Z(o[362]) );
  AND U3161 ( .A(n1035), .B(n3160), .Z(n3158) );
  XOR U3162 ( .A(creg[362]), .B(mod_mult_o[362]), .Z(n3160) );
  XNOR U3163 ( .A(n3161), .B(n3162), .Z(o[361]) );
  AND U3164 ( .A(n1035), .B(n3163), .Z(n3161) );
  XOR U3165 ( .A(creg[361]), .B(mod_mult_o[361]), .Z(n3163) );
  XNOR U3166 ( .A(n3164), .B(n3165), .Z(o[360]) );
  AND U3167 ( .A(n1035), .B(n3166), .Z(n3164) );
  XOR U3168 ( .A(creg[360]), .B(mod_mult_o[360]), .Z(n3166) );
  XNOR U3169 ( .A(n3167), .B(n3168), .Z(o[35]) );
  AND U3170 ( .A(n1035), .B(n3169), .Z(n3167) );
  XOR U3171 ( .A(creg[35]), .B(mod_mult_o[35]), .Z(n3169) );
  XNOR U3172 ( .A(n3170), .B(n3171), .Z(o[359]) );
  AND U3173 ( .A(n1035), .B(n3172), .Z(n3170) );
  XOR U3174 ( .A(creg[359]), .B(mod_mult_o[359]), .Z(n3172) );
  XNOR U3175 ( .A(n3173), .B(n3174), .Z(o[358]) );
  AND U3176 ( .A(n1035), .B(n3175), .Z(n3173) );
  XOR U3177 ( .A(creg[358]), .B(mod_mult_o[358]), .Z(n3175) );
  XNOR U3178 ( .A(n3176), .B(n3177), .Z(o[357]) );
  AND U3179 ( .A(n1035), .B(n3178), .Z(n3176) );
  XOR U3180 ( .A(creg[357]), .B(mod_mult_o[357]), .Z(n3178) );
  XNOR U3181 ( .A(n3179), .B(n3180), .Z(o[356]) );
  AND U3182 ( .A(n1035), .B(n3181), .Z(n3179) );
  XOR U3183 ( .A(creg[356]), .B(mod_mult_o[356]), .Z(n3181) );
  XNOR U3184 ( .A(n3182), .B(n3183), .Z(o[355]) );
  AND U3185 ( .A(n1035), .B(n3184), .Z(n3182) );
  XOR U3186 ( .A(creg[355]), .B(mod_mult_o[355]), .Z(n3184) );
  XNOR U3187 ( .A(n3185), .B(n3186), .Z(o[354]) );
  AND U3188 ( .A(n1035), .B(n3187), .Z(n3185) );
  XOR U3189 ( .A(creg[354]), .B(mod_mult_o[354]), .Z(n3187) );
  XNOR U3190 ( .A(n3188), .B(n3189), .Z(o[353]) );
  AND U3191 ( .A(n1035), .B(n3190), .Z(n3188) );
  XOR U3192 ( .A(creg[353]), .B(mod_mult_o[353]), .Z(n3190) );
  XNOR U3193 ( .A(n3191), .B(n3192), .Z(o[352]) );
  AND U3194 ( .A(n1035), .B(n3193), .Z(n3191) );
  XOR U3195 ( .A(creg[352]), .B(mod_mult_o[352]), .Z(n3193) );
  XNOR U3196 ( .A(n3194), .B(n3195), .Z(o[351]) );
  AND U3197 ( .A(n1035), .B(n3196), .Z(n3194) );
  XOR U3198 ( .A(creg[351]), .B(mod_mult_o[351]), .Z(n3196) );
  XNOR U3199 ( .A(n3197), .B(n3198), .Z(o[350]) );
  AND U3200 ( .A(n1035), .B(n3199), .Z(n3197) );
  XOR U3201 ( .A(creg[350]), .B(mod_mult_o[350]), .Z(n3199) );
  XNOR U3202 ( .A(n3200), .B(n3201), .Z(o[34]) );
  AND U3203 ( .A(n1035), .B(n3202), .Z(n3200) );
  XOR U3204 ( .A(creg[34]), .B(mod_mult_o[34]), .Z(n3202) );
  XNOR U3205 ( .A(n3203), .B(n3204), .Z(o[349]) );
  AND U3206 ( .A(n1035), .B(n3205), .Z(n3203) );
  XOR U3207 ( .A(creg[349]), .B(mod_mult_o[349]), .Z(n3205) );
  XNOR U3208 ( .A(n3206), .B(n3207), .Z(o[348]) );
  AND U3209 ( .A(n1035), .B(n3208), .Z(n3206) );
  XOR U3210 ( .A(creg[348]), .B(mod_mult_o[348]), .Z(n3208) );
  XNOR U3211 ( .A(n3209), .B(n3210), .Z(o[347]) );
  AND U3212 ( .A(n1035), .B(n3211), .Z(n3209) );
  XOR U3213 ( .A(creg[347]), .B(mod_mult_o[347]), .Z(n3211) );
  XNOR U3214 ( .A(n3212), .B(n3213), .Z(o[346]) );
  AND U3215 ( .A(n1035), .B(n3214), .Z(n3212) );
  XOR U3216 ( .A(creg[346]), .B(mod_mult_o[346]), .Z(n3214) );
  XNOR U3217 ( .A(n3215), .B(n3216), .Z(o[345]) );
  AND U3218 ( .A(n1035), .B(n3217), .Z(n3215) );
  XOR U3219 ( .A(creg[345]), .B(mod_mult_o[345]), .Z(n3217) );
  XNOR U3220 ( .A(n3218), .B(n3219), .Z(o[344]) );
  AND U3221 ( .A(n1035), .B(n3220), .Z(n3218) );
  XOR U3222 ( .A(creg[344]), .B(mod_mult_o[344]), .Z(n3220) );
  XNOR U3223 ( .A(n3221), .B(n3222), .Z(o[343]) );
  AND U3224 ( .A(n1035), .B(n3223), .Z(n3221) );
  XOR U3225 ( .A(creg[343]), .B(mod_mult_o[343]), .Z(n3223) );
  XNOR U3226 ( .A(n3224), .B(n3225), .Z(o[342]) );
  AND U3227 ( .A(n1035), .B(n3226), .Z(n3224) );
  XOR U3228 ( .A(creg[342]), .B(mod_mult_o[342]), .Z(n3226) );
  XNOR U3229 ( .A(n3227), .B(n3228), .Z(o[341]) );
  AND U3230 ( .A(n1035), .B(n3229), .Z(n3227) );
  XOR U3231 ( .A(creg[341]), .B(mod_mult_o[341]), .Z(n3229) );
  XNOR U3232 ( .A(n3230), .B(n3231), .Z(o[340]) );
  AND U3233 ( .A(n1035), .B(n3232), .Z(n3230) );
  XOR U3234 ( .A(creg[340]), .B(mod_mult_o[340]), .Z(n3232) );
  XNOR U3235 ( .A(n3233), .B(n3234), .Z(o[33]) );
  AND U3236 ( .A(n1035), .B(n3235), .Z(n3233) );
  XOR U3237 ( .A(creg[33]), .B(mod_mult_o[33]), .Z(n3235) );
  XNOR U3238 ( .A(n3236), .B(n3237), .Z(o[339]) );
  AND U3239 ( .A(n1035), .B(n3238), .Z(n3236) );
  XOR U3240 ( .A(creg[339]), .B(mod_mult_o[339]), .Z(n3238) );
  XNOR U3241 ( .A(n3239), .B(n3240), .Z(o[338]) );
  AND U3242 ( .A(n1035), .B(n3241), .Z(n3239) );
  XOR U3243 ( .A(creg[338]), .B(mod_mult_o[338]), .Z(n3241) );
  XNOR U3244 ( .A(n3242), .B(n3243), .Z(o[337]) );
  AND U3245 ( .A(n1035), .B(n3244), .Z(n3242) );
  XOR U3246 ( .A(creg[337]), .B(mod_mult_o[337]), .Z(n3244) );
  XNOR U3247 ( .A(n3245), .B(n3246), .Z(o[336]) );
  AND U3248 ( .A(n1035), .B(n3247), .Z(n3245) );
  XOR U3249 ( .A(creg[336]), .B(mod_mult_o[336]), .Z(n3247) );
  XNOR U3250 ( .A(n3248), .B(n3249), .Z(o[335]) );
  AND U3251 ( .A(n1035), .B(n3250), .Z(n3248) );
  XOR U3252 ( .A(creg[335]), .B(mod_mult_o[335]), .Z(n3250) );
  XNOR U3253 ( .A(n3251), .B(n3252), .Z(o[334]) );
  AND U3254 ( .A(n1035), .B(n3253), .Z(n3251) );
  XOR U3255 ( .A(creg[334]), .B(mod_mult_o[334]), .Z(n3253) );
  XNOR U3256 ( .A(n3254), .B(n3255), .Z(o[333]) );
  AND U3257 ( .A(n1035), .B(n3256), .Z(n3254) );
  XOR U3258 ( .A(creg[333]), .B(mod_mult_o[333]), .Z(n3256) );
  XNOR U3259 ( .A(n3257), .B(n3258), .Z(o[332]) );
  AND U3260 ( .A(n1035), .B(n3259), .Z(n3257) );
  XOR U3261 ( .A(creg[332]), .B(mod_mult_o[332]), .Z(n3259) );
  XNOR U3262 ( .A(n3260), .B(n3261), .Z(o[331]) );
  AND U3263 ( .A(n1035), .B(n3262), .Z(n3260) );
  XOR U3264 ( .A(creg[331]), .B(mod_mult_o[331]), .Z(n3262) );
  XNOR U3265 ( .A(n3263), .B(n3264), .Z(o[330]) );
  AND U3266 ( .A(n1035), .B(n3265), .Z(n3263) );
  XOR U3267 ( .A(creg[330]), .B(mod_mult_o[330]), .Z(n3265) );
  XNOR U3268 ( .A(n3266), .B(n3267), .Z(o[32]) );
  AND U3269 ( .A(n1035), .B(n3268), .Z(n3266) );
  XOR U3270 ( .A(creg[32]), .B(mod_mult_o[32]), .Z(n3268) );
  XNOR U3271 ( .A(n3269), .B(n3270), .Z(o[329]) );
  AND U3272 ( .A(n1035), .B(n3271), .Z(n3269) );
  XOR U3273 ( .A(creg[329]), .B(mod_mult_o[329]), .Z(n3271) );
  XNOR U3274 ( .A(n3272), .B(n3273), .Z(o[328]) );
  AND U3275 ( .A(n1035), .B(n3274), .Z(n3272) );
  XOR U3276 ( .A(creg[328]), .B(mod_mult_o[328]), .Z(n3274) );
  XNOR U3277 ( .A(n3275), .B(n3276), .Z(o[327]) );
  AND U3278 ( .A(n1035), .B(n3277), .Z(n3275) );
  XOR U3279 ( .A(creg[327]), .B(mod_mult_o[327]), .Z(n3277) );
  XNOR U3280 ( .A(n3278), .B(n3279), .Z(o[326]) );
  AND U3281 ( .A(n1035), .B(n3280), .Z(n3278) );
  XOR U3282 ( .A(creg[326]), .B(mod_mult_o[326]), .Z(n3280) );
  XNOR U3283 ( .A(n3281), .B(n3282), .Z(o[325]) );
  AND U3284 ( .A(n1035), .B(n3283), .Z(n3281) );
  XOR U3285 ( .A(creg[325]), .B(mod_mult_o[325]), .Z(n3283) );
  XNOR U3286 ( .A(n3284), .B(n3285), .Z(o[324]) );
  AND U3287 ( .A(n1035), .B(n3286), .Z(n3284) );
  XOR U3288 ( .A(creg[324]), .B(mod_mult_o[324]), .Z(n3286) );
  XNOR U3289 ( .A(n3287), .B(n3288), .Z(o[323]) );
  AND U3290 ( .A(n1035), .B(n3289), .Z(n3287) );
  XOR U3291 ( .A(creg[323]), .B(mod_mult_o[323]), .Z(n3289) );
  XNOR U3292 ( .A(n3290), .B(n3291), .Z(o[322]) );
  AND U3293 ( .A(n1035), .B(n3292), .Z(n3290) );
  XOR U3294 ( .A(creg[322]), .B(mod_mult_o[322]), .Z(n3292) );
  XNOR U3295 ( .A(n3293), .B(n3294), .Z(o[321]) );
  AND U3296 ( .A(n1035), .B(n3295), .Z(n3293) );
  XOR U3297 ( .A(creg[321]), .B(mod_mult_o[321]), .Z(n3295) );
  XNOR U3298 ( .A(n3296), .B(n3297), .Z(o[320]) );
  AND U3299 ( .A(n1035), .B(n3298), .Z(n3296) );
  XOR U3300 ( .A(creg[320]), .B(mod_mult_o[320]), .Z(n3298) );
  XNOR U3301 ( .A(n3299), .B(n3300), .Z(o[31]) );
  AND U3302 ( .A(n1035), .B(n3301), .Z(n3299) );
  XOR U3303 ( .A(creg[31]), .B(mod_mult_o[31]), .Z(n3301) );
  XNOR U3304 ( .A(n3302), .B(n3303), .Z(o[319]) );
  AND U3305 ( .A(n1035), .B(n3304), .Z(n3302) );
  XOR U3306 ( .A(creg[319]), .B(mod_mult_o[319]), .Z(n3304) );
  XNOR U3307 ( .A(n3305), .B(n3306), .Z(o[318]) );
  AND U3308 ( .A(n1035), .B(n3307), .Z(n3305) );
  XOR U3309 ( .A(creg[318]), .B(mod_mult_o[318]), .Z(n3307) );
  XNOR U3310 ( .A(n3308), .B(n3309), .Z(o[317]) );
  AND U3311 ( .A(n1035), .B(n3310), .Z(n3308) );
  XOR U3312 ( .A(creg[317]), .B(mod_mult_o[317]), .Z(n3310) );
  XNOR U3313 ( .A(n3311), .B(n3312), .Z(o[316]) );
  AND U3314 ( .A(n1035), .B(n3313), .Z(n3311) );
  XOR U3315 ( .A(creg[316]), .B(mod_mult_o[316]), .Z(n3313) );
  XNOR U3316 ( .A(n3314), .B(n3315), .Z(o[315]) );
  AND U3317 ( .A(n1035), .B(n3316), .Z(n3314) );
  XOR U3318 ( .A(creg[315]), .B(mod_mult_o[315]), .Z(n3316) );
  XNOR U3319 ( .A(n3317), .B(n3318), .Z(o[314]) );
  AND U3320 ( .A(n1035), .B(n3319), .Z(n3317) );
  XOR U3321 ( .A(creg[314]), .B(mod_mult_o[314]), .Z(n3319) );
  XNOR U3322 ( .A(n3320), .B(n3321), .Z(o[313]) );
  AND U3323 ( .A(n1035), .B(n3322), .Z(n3320) );
  XOR U3324 ( .A(creg[313]), .B(mod_mult_o[313]), .Z(n3322) );
  XNOR U3325 ( .A(n3323), .B(n3324), .Z(o[312]) );
  AND U3326 ( .A(n1035), .B(n3325), .Z(n3323) );
  XOR U3327 ( .A(creg[312]), .B(mod_mult_o[312]), .Z(n3325) );
  XNOR U3328 ( .A(n3326), .B(n3327), .Z(o[311]) );
  AND U3329 ( .A(n1035), .B(n3328), .Z(n3326) );
  XOR U3330 ( .A(creg[311]), .B(mod_mult_o[311]), .Z(n3328) );
  XNOR U3331 ( .A(n3329), .B(n3330), .Z(o[310]) );
  AND U3332 ( .A(n1035), .B(n3331), .Z(n3329) );
  XOR U3333 ( .A(creg[310]), .B(mod_mult_o[310]), .Z(n3331) );
  XNOR U3334 ( .A(n3332), .B(n3333), .Z(o[30]) );
  AND U3335 ( .A(n1035), .B(n3334), .Z(n3332) );
  XOR U3336 ( .A(creg[30]), .B(mod_mult_o[30]), .Z(n3334) );
  XNOR U3337 ( .A(n3335), .B(n3336), .Z(o[309]) );
  AND U3338 ( .A(n1035), .B(n3337), .Z(n3335) );
  XOR U3339 ( .A(creg[309]), .B(mod_mult_o[309]), .Z(n3337) );
  XNOR U3340 ( .A(n3338), .B(n3339), .Z(o[308]) );
  AND U3341 ( .A(n1035), .B(n3340), .Z(n3338) );
  XOR U3342 ( .A(creg[308]), .B(mod_mult_o[308]), .Z(n3340) );
  XNOR U3343 ( .A(n3341), .B(n3342), .Z(o[307]) );
  AND U3344 ( .A(n1035), .B(n3343), .Z(n3341) );
  XOR U3345 ( .A(creg[307]), .B(mod_mult_o[307]), .Z(n3343) );
  XNOR U3346 ( .A(n3344), .B(n3345), .Z(o[306]) );
  AND U3347 ( .A(n1035), .B(n3346), .Z(n3344) );
  XOR U3348 ( .A(creg[306]), .B(mod_mult_o[306]), .Z(n3346) );
  XNOR U3349 ( .A(n3347), .B(n3348), .Z(o[305]) );
  AND U3350 ( .A(n1035), .B(n3349), .Z(n3347) );
  XOR U3351 ( .A(creg[305]), .B(mod_mult_o[305]), .Z(n3349) );
  XNOR U3352 ( .A(n3350), .B(n3351), .Z(o[304]) );
  AND U3353 ( .A(n1035), .B(n3352), .Z(n3350) );
  XOR U3354 ( .A(creg[304]), .B(mod_mult_o[304]), .Z(n3352) );
  XNOR U3355 ( .A(n3353), .B(n3354), .Z(o[303]) );
  AND U3356 ( .A(n1035), .B(n3355), .Z(n3353) );
  XOR U3357 ( .A(creg[303]), .B(mod_mult_o[303]), .Z(n3355) );
  XNOR U3358 ( .A(n3356), .B(n3357), .Z(o[302]) );
  AND U3359 ( .A(n1035), .B(n3358), .Z(n3356) );
  XOR U3360 ( .A(creg[302]), .B(mod_mult_o[302]), .Z(n3358) );
  XNOR U3361 ( .A(n3359), .B(n3360), .Z(o[301]) );
  AND U3362 ( .A(n1035), .B(n3361), .Z(n3359) );
  XOR U3363 ( .A(creg[301]), .B(mod_mult_o[301]), .Z(n3361) );
  XNOR U3364 ( .A(n3362), .B(n3363), .Z(o[300]) );
  AND U3365 ( .A(n1035), .B(n3364), .Z(n3362) );
  XOR U3366 ( .A(creg[300]), .B(mod_mult_o[300]), .Z(n3364) );
  XNOR U3367 ( .A(n3365), .B(n3366), .Z(o[2]) );
  AND U3368 ( .A(n1035), .B(n3367), .Z(n3365) );
  XOR U3369 ( .A(creg[2]), .B(mod_mult_o[2]), .Z(n3367) );
  XNOR U3370 ( .A(n3368), .B(n3369), .Z(o[29]) );
  AND U3371 ( .A(n1035), .B(n3370), .Z(n3368) );
  XOR U3372 ( .A(creg[29]), .B(mod_mult_o[29]), .Z(n3370) );
  XNOR U3373 ( .A(n3371), .B(n3372), .Z(o[299]) );
  AND U3374 ( .A(n1035), .B(n3373), .Z(n3371) );
  XOR U3375 ( .A(creg[299]), .B(mod_mult_o[299]), .Z(n3373) );
  XNOR U3376 ( .A(n3374), .B(n3375), .Z(o[298]) );
  AND U3377 ( .A(n1035), .B(n3376), .Z(n3374) );
  XOR U3378 ( .A(creg[298]), .B(mod_mult_o[298]), .Z(n3376) );
  XNOR U3379 ( .A(n3377), .B(n3378), .Z(o[297]) );
  AND U3380 ( .A(n1035), .B(n3379), .Z(n3377) );
  XOR U3381 ( .A(creg[297]), .B(mod_mult_o[297]), .Z(n3379) );
  XNOR U3382 ( .A(n3380), .B(n3381), .Z(o[296]) );
  AND U3383 ( .A(n1035), .B(n3382), .Z(n3380) );
  XOR U3384 ( .A(creg[296]), .B(mod_mult_o[296]), .Z(n3382) );
  XNOR U3385 ( .A(n3383), .B(n3384), .Z(o[295]) );
  AND U3386 ( .A(n1035), .B(n3385), .Z(n3383) );
  XOR U3387 ( .A(creg[295]), .B(mod_mult_o[295]), .Z(n3385) );
  XNOR U3388 ( .A(n3386), .B(n3387), .Z(o[294]) );
  AND U3389 ( .A(n1035), .B(n3388), .Z(n3386) );
  XOR U3390 ( .A(creg[294]), .B(mod_mult_o[294]), .Z(n3388) );
  XNOR U3391 ( .A(n3389), .B(n3390), .Z(o[293]) );
  AND U3392 ( .A(n1035), .B(n3391), .Z(n3389) );
  XOR U3393 ( .A(creg[293]), .B(mod_mult_o[293]), .Z(n3391) );
  XNOR U3394 ( .A(n3392), .B(n3393), .Z(o[292]) );
  AND U3395 ( .A(n1035), .B(n3394), .Z(n3392) );
  XOR U3396 ( .A(creg[292]), .B(mod_mult_o[292]), .Z(n3394) );
  XNOR U3397 ( .A(n3395), .B(n3396), .Z(o[291]) );
  AND U3398 ( .A(n1035), .B(n3397), .Z(n3395) );
  XOR U3399 ( .A(creg[291]), .B(mod_mult_o[291]), .Z(n3397) );
  XNOR U3400 ( .A(n3398), .B(n3399), .Z(o[290]) );
  AND U3401 ( .A(n1035), .B(n3400), .Z(n3398) );
  XOR U3402 ( .A(creg[290]), .B(mod_mult_o[290]), .Z(n3400) );
  XNOR U3403 ( .A(n3401), .B(n3402), .Z(o[28]) );
  AND U3404 ( .A(n1035), .B(n3403), .Z(n3401) );
  XOR U3405 ( .A(creg[28]), .B(mod_mult_o[28]), .Z(n3403) );
  XNOR U3406 ( .A(n3404), .B(n3405), .Z(o[289]) );
  AND U3407 ( .A(n1035), .B(n3406), .Z(n3404) );
  XOR U3408 ( .A(creg[289]), .B(mod_mult_o[289]), .Z(n3406) );
  XNOR U3409 ( .A(n3407), .B(n3408), .Z(o[288]) );
  AND U3410 ( .A(n1035), .B(n3409), .Z(n3407) );
  XOR U3411 ( .A(creg[288]), .B(mod_mult_o[288]), .Z(n3409) );
  XNOR U3412 ( .A(n3410), .B(n3411), .Z(o[287]) );
  AND U3413 ( .A(n1035), .B(n3412), .Z(n3410) );
  XOR U3414 ( .A(creg[287]), .B(mod_mult_o[287]), .Z(n3412) );
  XNOR U3415 ( .A(n3413), .B(n3414), .Z(o[286]) );
  AND U3416 ( .A(n1035), .B(n3415), .Z(n3413) );
  XOR U3417 ( .A(creg[286]), .B(mod_mult_o[286]), .Z(n3415) );
  XNOR U3418 ( .A(n3416), .B(n3417), .Z(o[285]) );
  AND U3419 ( .A(n1035), .B(n3418), .Z(n3416) );
  XOR U3420 ( .A(creg[285]), .B(mod_mult_o[285]), .Z(n3418) );
  XNOR U3421 ( .A(n3419), .B(n3420), .Z(o[284]) );
  AND U3422 ( .A(n1035), .B(n3421), .Z(n3419) );
  XOR U3423 ( .A(creg[284]), .B(mod_mult_o[284]), .Z(n3421) );
  XNOR U3424 ( .A(n3422), .B(n3423), .Z(o[283]) );
  AND U3425 ( .A(n1035), .B(n3424), .Z(n3422) );
  XOR U3426 ( .A(creg[283]), .B(mod_mult_o[283]), .Z(n3424) );
  XNOR U3427 ( .A(n3425), .B(n3426), .Z(o[282]) );
  AND U3428 ( .A(n1035), .B(n3427), .Z(n3425) );
  XOR U3429 ( .A(creg[282]), .B(mod_mult_o[282]), .Z(n3427) );
  XNOR U3430 ( .A(n3428), .B(n3429), .Z(o[281]) );
  AND U3431 ( .A(n1035), .B(n3430), .Z(n3428) );
  XOR U3432 ( .A(creg[281]), .B(mod_mult_o[281]), .Z(n3430) );
  XNOR U3433 ( .A(n3431), .B(n3432), .Z(o[280]) );
  AND U3434 ( .A(n1035), .B(n3433), .Z(n3431) );
  XOR U3435 ( .A(creg[280]), .B(mod_mult_o[280]), .Z(n3433) );
  XNOR U3436 ( .A(n3434), .B(n3435), .Z(o[27]) );
  AND U3437 ( .A(n1035), .B(n3436), .Z(n3434) );
  XOR U3438 ( .A(creg[27]), .B(mod_mult_o[27]), .Z(n3436) );
  XNOR U3439 ( .A(n3437), .B(n3438), .Z(o[279]) );
  AND U3440 ( .A(n1035), .B(n3439), .Z(n3437) );
  XOR U3441 ( .A(creg[279]), .B(mod_mult_o[279]), .Z(n3439) );
  XNOR U3442 ( .A(n3440), .B(n3441), .Z(o[278]) );
  AND U3443 ( .A(n1035), .B(n3442), .Z(n3440) );
  XOR U3444 ( .A(creg[278]), .B(mod_mult_o[278]), .Z(n3442) );
  XNOR U3445 ( .A(n3443), .B(n3444), .Z(o[277]) );
  AND U3446 ( .A(n1035), .B(n3445), .Z(n3443) );
  XOR U3447 ( .A(creg[277]), .B(mod_mult_o[277]), .Z(n3445) );
  XNOR U3448 ( .A(n3446), .B(n3447), .Z(o[276]) );
  AND U3449 ( .A(n1035), .B(n3448), .Z(n3446) );
  XOR U3450 ( .A(creg[276]), .B(mod_mult_o[276]), .Z(n3448) );
  XNOR U3451 ( .A(n3449), .B(n3450), .Z(o[275]) );
  AND U3452 ( .A(n1035), .B(n3451), .Z(n3449) );
  XOR U3453 ( .A(creg[275]), .B(mod_mult_o[275]), .Z(n3451) );
  XNOR U3454 ( .A(n3452), .B(n3453), .Z(o[274]) );
  AND U3455 ( .A(n1035), .B(n3454), .Z(n3452) );
  XOR U3456 ( .A(creg[274]), .B(mod_mult_o[274]), .Z(n3454) );
  XNOR U3457 ( .A(n3455), .B(n3456), .Z(o[273]) );
  AND U3458 ( .A(n1035), .B(n3457), .Z(n3455) );
  XOR U3459 ( .A(creg[273]), .B(mod_mult_o[273]), .Z(n3457) );
  XNOR U3460 ( .A(n3458), .B(n3459), .Z(o[272]) );
  AND U3461 ( .A(n1035), .B(n3460), .Z(n3458) );
  XOR U3462 ( .A(creg[272]), .B(mod_mult_o[272]), .Z(n3460) );
  XNOR U3463 ( .A(n3461), .B(n3462), .Z(o[271]) );
  AND U3464 ( .A(n1035), .B(n3463), .Z(n3461) );
  XOR U3465 ( .A(creg[271]), .B(mod_mult_o[271]), .Z(n3463) );
  XNOR U3466 ( .A(n3464), .B(n3465), .Z(o[270]) );
  AND U3467 ( .A(n1035), .B(n3466), .Z(n3464) );
  XOR U3468 ( .A(creg[270]), .B(mod_mult_o[270]), .Z(n3466) );
  XNOR U3469 ( .A(n3467), .B(n3468), .Z(o[26]) );
  AND U3470 ( .A(n1035), .B(n3469), .Z(n3467) );
  XOR U3471 ( .A(creg[26]), .B(mod_mult_o[26]), .Z(n3469) );
  XNOR U3472 ( .A(n3470), .B(n3471), .Z(o[269]) );
  AND U3473 ( .A(n1035), .B(n3472), .Z(n3470) );
  XOR U3474 ( .A(creg[269]), .B(mod_mult_o[269]), .Z(n3472) );
  XNOR U3475 ( .A(n3473), .B(n3474), .Z(o[268]) );
  AND U3476 ( .A(n1035), .B(n3475), .Z(n3473) );
  XOR U3477 ( .A(creg[268]), .B(mod_mult_o[268]), .Z(n3475) );
  XNOR U3478 ( .A(n3476), .B(n3477), .Z(o[267]) );
  AND U3479 ( .A(n1035), .B(n3478), .Z(n3476) );
  XOR U3480 ( .A(creg[267]), .B(mod_mult_o[267]), .Z(n3478) );
  XNOR U3481 ( .A(n3479), .B(n3480), .Z(o[266]) );
  AND U3482 ( .A(n1035), .B(n3481), .Z(n3479) );
  XOR U3483 ( .A(creg[266]), .B(mod_mult_o[266]), .Z(n3481) );
  XNOR U3484 ( .A(n3482), .B(n3483), .Z(o[265]) );
  AND U3485 ( .A(n1035), .B(n3484), .Z(n3482) );
  XOR U3486 ( .A(creg[265]), .B(mod_mult_o[265]), .Z(n3484) );
  XNOR U3487 ( .A(n3485), .B(n3486), .Z(o[264]) );
  AND U3488 ( .A(n1035), .B(n3487), .Z(n3485) );
  XOR U3489 ( .A(creg[264]), .B(mod_mult_o[264]), .Z(n3487) );
  XNOR U3490 ( .A(n3488), .B(n3489), .Z(o[263]) );
  AND U3491 ( .A(n1035), .B(n3490), .Z(n3488) );
  XOR U3492 ( .A(creg[263]), .B(mod_mult_o[263]), .Z(n3490) );
  XNOR U3493 ( .A(n3491), .B(n3492), .Z(o[262]) );
  AND U3494 ( .A(n1035), .B(n3493), .Z(n3491) );
  XOR U3495 ( .A(creg[262]), .B(mod_mult_o[262]), .Z(n3493) );
  XNOR U3496 ( .A(n3494), .B(n3495), .Z(o[261]) );
  AND U3497 ( .A(n1035), .B(n3496), .Z(n3494) );
  XOR U3498 ( .A(creg[261]), .B(mod_mult_o[261]), .Z(n3496) );
  XNOR U3499 ( .A(n3497), .B(n3498), .Z(o[260]) );
  AND U3500 ( .A(n1035), .B(n3499), .Z(n3497) );
  XOR U3501 ( .A(creg[260]), .B(mod_mult_o[260]), .Z(n3499) );
  XNOR U3502 ( .A(n3500), .B(n3501), .Z(o[25]) );
  AND U3503 ( .A(n1035), .B(n3502), .Z(n3500) );
  XOR U3504 ( .A(creg[25]), .B(mod_mult_o[25]), .Z(n3502) );
  XNOR U3505 ( .A(n3503), .B(n3504), .Z(o[259]) );
  AND U3506 ( .A(n1035), .B(n3505), .Z(n3503) );
  XOR U3507 ( .A(creg[259]), .B(mod_mult_o[259]), .Z(n3505) );
  XNOR U3508 ( .A(n3506), .B(n3507), .Z(o[258]) );
  AND U3509 ( .A(n1035), .B(n3508), .Z(n3506) );
  XOR U3510 ( .A(creg[258]), .B(mod_mult_o[258]), .Z(n3508) );
  XNOR U3511 ( .A(n3509), .B(n3510), .Z(o[257]) );
  AND U3512 ( .A(n1035), .B(n3511), .Z(n3509) );
  XOR U3513 ( .A(creg[257]), .B(mod_mult_o[257]), .Z(n3511) );
  XNOR U3514 ( .A(n3512), .B(n3513), .Z(o[256]) );
  AND U3515 ( .A(n1035), .B(n3514), .Z(n3512) );
  XOR U3516 ( .A(creg[256]), .B(mod_mult_o[256]), .Z(n3514) );
  XNOR U3517 ( .A(n3515), .B(n3516), .Z(o[255]) );
  AND U3518 ( .A(n1035), .B(n3517), .Z(n3515) );
  XOR U3519 ( .A(creg[255]), .B(mod_mult_o[255]), .Z(n3517) );
  XNOR U3520 ( .A(n3518), .B(n3519), .Z(o[254]) );
  AND U3521 ( .A(n1035), .B(n3520), .Z(n3518) );
  XOR U3522 ( .A(creg[254]), .B(mod_mult_o[254]), .Z(n3520) );
  XNOR U3523 ( .A(n3521), .B(n3522), .Z(o[253]) );
  AND U3524 ( .A(n1035), .B(n3523), .Z(n3521) );
  XOR U3525 ( .A(creg[253]), .B(mod_mult_o[253]), .Z(n3523) );
  XNOR U3526 ( .A(n3524), .B(n3525), .Z(o[252]) );
  AND U3527 ( .A(n1035), .B(n3526), .Z(n3524) );
  XOR U3528 ( .A(creg[252]), .B(mod_mult_o[252]), .Z(n3526) );
  XNOR U3529 ( .A(n3527), .B(n3528), .Z(o[251]) );
  AND U3530 ( .A(n1035), .B(n3529), .Z(n3527) );
  XOR U3531 ( .A(creg[251]), .B(mod_mult_o[251]), .Z(n3529) );
  XNOR U3532 ( .A(n3530), .B(n3531), .Z(o[250]) );
  AND U3533 ( .A(n1035), .B(n3532), .Z(n3530) );
  XOR U3534 ( .A(creg[250]), .B(mod_mult_o[250]), .Z(n3532) );
  XNOR U3535 ( .A(n3533), .B(n3534), .Z(o[24]) );
  AND U3536 ( .A(n1035), .B(n3535), .Z(n3533) );
  XOR U3537 ( .A(creg[24]), .B(mod_mult_o[24]), .Z(n3535) );
  XNOR U3538 ( .A(n3536), .B(n3537), .Z(o[249]) );
  AND U3539 ( .A(n1035), .B(n3538), .Z(n3536) );
  XOR U3540 ( .A(creg[249]), .B(mod_mult_o[249]), .Z(n3538) );
  XNOR U3541 ( .A(n3539), .B(n3540), .Z(o[248]) );
  AND U3542 ( .A(n1035), .B(n3541), .Z(n3539) );
  XOR U3543 ( .A(creg[248]), .B(mod_mult_o[248]), .Z(n3541) );
  XNOR U3544 ( .A(n3542), .B(n3543), .Z(o[247]) );
  AND U3545 ( .A(n1035), .B(n3544), .Z(n3542) );
  XOR U3546 ( .A(creg[247]), .B(mod_mult_o[247]), .Z(n3544) );
  XNOR U3547 ( .A(n3545), .B(n3546), .Z(o[246]) );
  AND U3548 ( .A(n1035), .B(n3547), .Z(n3545) );
  XOR U3549 ( .A(creg[246]), .B(mod_mult_o[246]), .Z(n3547) );
  XNOR U3550 ( .A(n3548), .B(n3549), .Z(o[245]) );
  AND U3551 ( .A(n1035), .B(n3550), .Z(n3548) );
  XOR U3552 ( .A(creg[245]), .B(mod_mult_o[245]), .Z(n3550) );
  XNOR U3553 ( .A(n3551), .B(n3552), .Z(o[244]) );
  AND U3554 ( .A(n1035), .B(n3553), .Z(n3551) );
  XOR U3555 ( .A(creg[244]), .B(mod_mult_o[244]), .Z(n3553) );
  XNOR U3556 ( .A(n3554), .B(n3555), .Z(o[243]) );
  AND U3557 ( .A(n1035), .B(n3556), .Z(n3554) );
  XOR U3558 ( .A(creg[243]), .B(mod_mult_o[243]), .Z(n3556) );
  XNOR U3559 ( .A(n3557), .B(n3558), .Z(o[242]) );
  AND U3560 ( .A(n1035), .B(n3559), .Z(n3557) );
  XOR U3561 ( .A(creg[242]), .B(mod_mult_o[242]), .Z(n3559) );
  XNOR U3562 ( .A(n3560), .B(n3561), .Z(o[241]) );
  AND U3563 ( .A(n1035), .B(n3562), .Z(n3560) );
  XOR U3564 ( .A(creg[241]), .B(mod_mult_o[241]), .Z(n3562) );
  XNOR U3565 ( .A(n3563), .B(n3564), .Z(o[240]) );
  AND U3566 ( .A(n1035), .B(n3565), .Z(n3563) );
  XOR U3567 ( .A(creg[240]), .B(mod_mult_o[240]), .Z(n3565) );
  XNOR U3568 ( .A(n3566), .B(n3567), .Z(o[23]) );
  AND U3569 ( .A(n1035), .B(n3568), .Z(n3566) );
  XOR U3570 ( .A(creg[23]), .B(mod_mult_o[23]), .Z(n3568) );
  XNOR U3571 ( .A(n3569), .B(n3570), .Z(o[239]) );
  AND U3572 ( .A(n1035), .B(n3571), .Z(n3569) );
  XOR U3573 ( .A(creg[239]), .B(mod_mult_o[239]), .Z(n3571) );
  XNOR U3574 ( .A(n3572), .B(n3573), .Z(o[238]) );
  AND U3575 ( .A(n1035), .B(n3574), .Z(n3572) );
  XOR U3576 ( .A(creg[238]), .B(mod_mult_o[238]), .Z(n3574) );
  XNOR U3577 ( .A(n3575), .B(n3576), .Z(o[237]) );
  AND U3578 ( .A(n1035), .B(n3577), .Z(n3575) );
  XOR U3579 ( .A(creg[237]), .B(mod_mult_o[237]), .Z(n3577) );
  XNOR U3580 ( .A(n3578), .B(n3579), .Z(o[236]) );
  AND U3581 ( .A(n1035), .B(n3580), .Z(n3578) );
  XOR U3582 ( .A(creg[236]), .B(mod_mult_o[236]), .Z(n3580) );
  XNOR U3583 ( .A(n3581), .B(n3582), .Z(o[235]) );
  AND U3584 ( .A(n1035), .B(n3583), .Z(n3581) );
  XOR U3585 ( .A(creg[235]), .B(mod_mult_o[235]), .Z(n3583) );
  XNOR U3586 ( .A(n3584), .B(n3585), .Z(o[234]) );
  AND U3587 ( .A(n1035), .B(n3586), .Z(n3584) );
  XOR U3588 ( .A(creg[234]), .B(mod_mult_o[234]), .Z(n3586) );
  XNOR U3589 ( .A(n3587), .B(n3588), .Z(o[233]) );
  AND U3590 ( .A(n1035), .B(n3589), .Z(n3587) );
  XOR U3591 ( .A(creg[233]), .B(mod_mult_o[233]), .Z(n3589) );
  XNOR U3592 ( .A(n3590), .B(n3591), .Z(o[232]) );
  AND U3593 ( .A(n1035), .B(n3592), .Z(n3590) );
  XOR U3594 ( .A(creg[232]), .B(mod_mult_o[232]), .Z(n3592) );
  XNOR U3595 ( .A(n3593), .B(n3594), .Z(o[231]) );
  AND U3596 ( .A(n1035), .B(n3595), .Z(n3593) );
  XOR U3597 ( .A(creg[231]), .B(mod_mult_o[231]), .Z(n3595) );
  XNOR U3598 ( .A(n3596), .B(n3597), .Z(o[230]) );
  AND U3599 ( .A(n1035), .B(n3598), .Z(n3596) );
  XOR U3600 ( .A(creg[230]), .B(mod_mult_o[230]), .Z(n3598) );
  XNOR U3601 ( .A(n3599), .B(n3600), .Z(o[22]) );
  AND U3602 ( .A(n1035), .B(n3601), .Z(n3599) );
  XOR U3603 ( .A(creg[22]), .B(mod_mult_o[22]), .Z(n3601) );
  XNOR U3604 ( .A(n3602), .B(n3603), .Z(o[229]) );
  AND U3605 ( .A(n1035), .B(n3604), .Z(n3602) );
  XOR U3606 ( .A(creg[229]), .B(mod_mult_o[229]), .Z(n3604) );
  XNOR U3607 ( .A(n3605), .B(n3606), .Z(o[228]) );
  AND U3608 ( .A(n1035), .B(n3607), .Z(n3605) );
  XOR U3609 ( .A(creg[228]), .B(mod_mult_o[228]), .Z(n3607) );
  XNOR U3610 ( .A(n3608), .B(n3609), .Z(o[227]) );
  AND U3611 ( .A(n1035), .B(n3610), .Z(n3608) );
  XOR U3612 ( .A(creg[227]), .B(mod_mult_o[227]), .Z(n3610) );
  XNOR U3613 ( .A(n3611), .B(n3612), .Z(o[226]) );
  AND U3614 ( .A(n1035), .B(n3613), .Z(n3611) );
  XOR U3615 ( .A(creg[226]), .B(mod_mult_o[226]), .Z(n3613) );
  XNOR U3616 ( .A(n3614), .B(n3615), .Z(o[225]) );
  AND U3617 ( .A(n1035), .B(n3616), .Z(n3614) );
  XOR U3618 ( .A(creg[225]), .B(mod_mult_o[225]), .Z(n3616) );
  XNOR U3619 ( .A(n3617), .B(n3618), .Z(o[224]) );
  AND U3620 ( .A(n1035), .B(n3619), .Z(n3617) );
  XOR U3621 ( .A(creg[224]), .B(mod_mult_o[224]), .Z(n3619) );
  XNOR U3622 ( .A(n3620), .B(n3621), .Z(o[223]) );
  AND U3623 ( .A(n1035), .B(n3622), .Z(n3620) );
  XOR U3624 ( .A(creg[223]), .B(mod_mult_o[223]), .Z(n3622) );
  XNOR U3625 ( .A(n3623), .B(n3624), .Z(o[222]) );
  AND U3626 ( .A(n1035), .B(n3625), .Z(n3623) );
  XOR U3627 ( .A(creg[222]), .B(mod_mult_o[222]), .Z(n3625) );
  XNOR U3628 ( .A(n3626), .B(n3627), .Z(o[221]) );
  AND U3629 ( .A(n1035), .B(n3628), .Z(n3626) );
  XOR U3630 ( .A(creg[221]), .B(mod_mult_o[221]), .Z(n3628) );
  XNOR U3631 ( .A(n3629), .B(n3630), .Z(o[220]) );
  AND U3632 ( .A(n1035), .B(n3631), .Z(n3629) );
  XOR U3633 ( .A(creg[220]), .B(mod_mult_o[220]), .Z(n3631) );
  XNOR U3634 ( .A(n3632), .B(n3633), .Z(o[21]) );
  AND U3635 ( .A(n1035), .B(n3634), .Z(n3632) );
  XOR U3636 ( .A(creg[21]), .B(mod_mult_o[21]), .Z(n3634) );
  XNOR U3637 ( .A(n3635), .B(n3636), .Z(o[219]) );
  AND U3638 ( .A(n1035), .B(n3637), .Z(n3635) );
  XOR U3639 ( .A(creg[219]), .B(mod_mult_o[219]), .Z(n3637) );
  XNOR U3640 ( .A(n3638), .B(n3639), .Z(o[218]) );
  AND U3641 ( .A(n1035), .B(n3640), .Z(n3638) );
  XOR U3642 ( .A(creg[218]), .B(mod_mult_o[218]), .Z(n3640) );
  XNOR U3643 ( .A(n3641), .B(n3642), .Z(o[217]) );
  AND U3644 ( .A(n1035), .B(n3643), .Z(n3641) );
  XOR U3645 ( .A(creg[217]), .B(mod_mult_o[217]), .Z(n3643) );
  XNOR U3646 ( .A(n3644), .B(n3645), .Z(o[216]) );
  AND U3647 ( .A(n1035), .B(n3646), .Z(n3644) );
  XOR U3648 ( .A(creg[216]), .B(mod_mult_o[216]), .Z(n3646) );
  XNOR U3649 ( .A(n3647), .B(n3648), .Z(o[215]) );
  AND U3650 ( .A(n1035), .B(n3649), .Z(n3647) );
  XOR U3651 ( .A(creg[215]), .B(mod_mult_o[215]), .Z(n3649) );
  XNOR U3652 ( .A(n3650), .B(n3651), .Z(o[214]) );
  AND U3653 ( .A(n1035), .B(n3652), .Z(n3650) );
  XOR U3654 ( .A(creg[214]), .B(mod_mult_o[214]), .Z(n3652) );
  XNOR U3655 ( .A(n3653), .B(n3654), .Z(o[213]) );
  AND U3656 ( .A(n1035), .B(n3655), .Z(n3653) );
  XOR U3657 ( .A(creg[213]), .B(mod_mult_o[213]), .Z(n3655) );
  XNOR U3658 ( .A(n3656), .B(n3657), .Z(o[212]) );
  AND U3659 ( .A(n1035), .B(n3658), .Z(n3656) );
  XOR U3660 ( .A(creg[212]), .B(mod_mult_o[212]), .Z(n3658) );
  XNOR U3661 ( .A(n3659), .B(n3660), .Z(o[211]) );
  AND U3662 ( .A(n1035), .B(n3661), .Z(n3659) );
  XOR U3663 ( .A(creg[211]), .B(mod_mult_o[211]), .Z(n3661) );
  XNOR U3664 ( .A(n3662), .B(n3663), .Z(o[210]) );
  AND U3665 ( .A(n1035), .B(n3664), .Z(n3662) );
  XOR U3666 ( .A(creg[210]), .B(mod_mult_o[210]), .Z(n3664) );
  XNOR U3667 ( .A(n3665), .B(n3666), .Z(o[20]) );
  AND U3668 ( .A(n1035), .B(n3667), .Z(n3665) );
  XOR U3669 ( .A(creg[20]), .B(mod_mult_o[20]), .Z(n3667) );
  XNOR U3670 ( .A(n3668), .B(n3669), .Z(o[209]) );
  AND U3671 ( .A(n1035), .B(n3670), .Z(n3668) );
  XOR U3672 ( .A(creg[209]), .B(mod_mult_o[209]), .Z(n3670) );
  XNOR U3673 ( .A(n3671), .B(n3672), .Z(o[208]) );
  AND U3674 ( .A(n1035), .B(n3673), .Z(n3671) );
  XOR U3675 ( .A(creg[208]), .B(mod_mult_o[208]), .Z(n3673) );
  XNOR U3676 ( .A(n3674), .B(n3675), .Z(o[207]) );
  AND U3677 ( .A(n1035), .B(n3676), .Z(n3674) );
  XOR U3678 ( .A(creg[207]), .B(mod_mult_o[207]), .Z(n3676) );
  XNOR U3679 ( .A(n3677), .B(n3678), .Z(o[206]) );
  AND U3680 ( .A(n1035), .B(n3679), .Z(n3677) );
  XOR U3681 ( .A(creg[206]), .B(mod_mult_o[206]), .Z(n3679) );
  XNOR U3682 ( .A(n3680), .B(n3681), .Z(o[205]) );
  AND U3683 ( .A(n1035), .B(n3682), .Z(n3680) );
  XOR U3684 ( .A(creg[205]), .B(mod_mult_o[205]), .Z(n3682) );
  XNOR U3685 ( .A(n3683), .B(n3684), .Z(o[204]) );
  AND U3686 ( .A(n1035), .B(n3685), .Z(n3683) );
  XOR U3687 ( .A(creg[204]), .B(mod_mult_o[204]), .Z(n3685) );
  XNOR U3688 ( .A(n3686), .B(n3687), .Z(o[203]) );
  AND U3689 ( .A(n1035), .B(n3688), .Z(n3686) );
  XOR U3690 ( .A(creg[203]), .B(mod_mult_o[203]), .Z(n3688) );
  XNOR U3691 ( .A(n3689), .B(n3690), .Z(o[202]) );
  AND U3692 ( .A(n1035), .B(n3691), .Z(n3689) );
  XOR U3693 ( .A(creg[202]), .B(mod_mult_o[202]), .Z(n3691) );
  XNOR U3694 ( .A(n3692), .B(n3693), .Z(o[201]) );
  AND U3695 ( .A(n1035), .B(n3694), .Z(n3692) );
  XOR U3696 ( .A(creg[201]), .B(mod_mult_o[201]), .Z(n3694) );
  XNOR U3697 ( .A(n3695), .B(n3696), .Z(o[200]) );
  AND U3698 ( .A(n1035), .B(n3697), .Z(n3695) );
  XOR U3699 ( .A(creg[200]), .B(mod_mult_o[200]), .Z(n3697) );
  XNOR U3700 ( .A(n3698), .B(n3699), .Z(o[1]) );
  AND U3701 ( .A(n1035), .B(n3700), .Z(n3698) );
  XOR U3702 ( .A(creg[1]), .B(mod_mult_o[1]), .Z(n3700) );
  XNOR U3703 ( .A(n3701), .B(n3702), .Z(o[19]) );
  AND U3704 ( .A(n1035), .B(n3703), .Z(n3701) );
  XOR U3705 ( .A(creg[19]), .B(mod_mult_o[19]), .Z(n3703) );
  XNOR U3706 ( .A(n3704), .B(n3705), .Z(o[199]) );
  AND U3707 ( .A(n1035), .B(n3706), .Z(n3704) );
  XOR U3708 ( .A(creg[199]), .B(mod_mult_o[199]), .Z(n3706) );
  XNOR U3709 ( .A(n3707), .B(n3708), .Z(o[198]) );
  AND U3710 ( .A(n1035), .B(n3709), .Z(n3707) );
  XOR U3711 ( .A(creg[198]), .B(mod_mult_o[198]), .Z(n3709) );
  XNOR U3712 ( .A(n3710), .B(n3711), .Z(o[197]) );
  AND U3713 ( .A(n1035), .B(n3712), .Z(n3710) );
  XOR U3714 ( .A(creg[197]), .B(mod_mult_o[197]), .Z(n3712) );
  XNOR U3715 ( .A(n3713), .B(n3714), .Z(o[196]) );
  AND U3716 ( .A(n1035), .B(n3715), .Z(n3713) );
  XOR U3717 ( .A(creg[196]), .B(mod_mult_o[196]), .Z(n3715) );
  XNOR U3718 ( .A(n3716), .B(n3717), .Z(o[195]) );
  AND U3719 ( .A(n1035), .B(n3718), .Z(n3716) );
  XOR U3720 ( .A(creg[195]), .B(mod_mult_o[195]), .Z(n3718) );
  XNOR U3721 ( .A(n3719), .B(n3720), .Z(o[194]) );
  AND U3722 ( .A(n1035), .B(n3721), .Z(n3719) );
  XOR U3723 ( .A(creg[194]), .B(mod_mult_o[194]), .Z(n3721) );
  XNOR U3724 ( .A(n3722), .B(n3723), .Z(o[193]) );
  AND U3725 ( .A(n1035), .B(n3724), .Z(n3722) );
  XOR U3726 ( .A(creg[193]), .B(mod_mult_o[193]), .Z(n3724) );
  XNOR U3727 ( .A(n3725), .B(n3726), .Z(o[192]) );
  AND U3728 ( .A(n1035), .B(n3727), .Z(n3725) );
  XOR U3729 ( .A(creg[192]), .B(mod_mult_o[192]), .Z(n3727) );
  XNOR U3730 ( .A(n3728), .B(n3729), .Z(o[191]) );
  AND U3731 ( .A(n1035), .B(n3730), .Z(n3728) );
  XOR U3732 ( .A(creg[191]), .B(mod_mult_o[191]), .Z(n3730) );
  XNOR U3733 ( .A(n3731), .B(n3732), .Z(o[190]) );
  AND U3734 ( .A(n1035), .B(n3733), .Z(n3731) );
  XOR U3735 ( .A(creg[190]), .B(mod_mult_o[190]), .Z(n3733) );
  XNOR U3736 ( .A(n3734), .B(n3735), .Z(o[18]) );
  AND U3737 ( .A(n1035), .B(n3736), .Z(n3734) );
  XOR U3738 ( .A(creg[18]), .B(mod_mult_o[18]), .Z(n3736) );
  XNOR U3739 ( .A(n3737), .B(n3738), .Z(o[189]) );
  AND U3740 ( .A(n1035), .B(n3739), .Z(n3737) );
  XOR U3741 ( .A(creg[189]), .B(mod_mult_o[189]), .Z(n3739) );
  XNOR U3742 ( .A(n3740), .B(n3741), .Z(o[188]) );
  AND U3743 ( .A(n1035), .B(n3742), .Z(n3740) );
  XOR U3744 ( .A(creg[188]), .B(mod_mult_o[188]), .Z(n3742) );
  XNOR U3745 ( .A(n3743), .B(n3744), .Z(o[187]) );
  AND U3746 ( .A(n1035), .B(n3745), .Z(n3743) );
  XOR U3747 ( .A(creg[187]), .B(mod_mult_o[187]), .Z(n3745) );
  XNOR U3748 ( .A(n3746), .B(n3747), .Z(o[186]) );
  AND U3749 ( .A(n1035), .B(n3748), .Z(n3746) );
  XOR U3750 ( .A(creg[186]), .B(mod_mult_o[186]), .Z(n3748) );
  XNOR U3751 ( .A(n3749), .B(n3750), .Z(o[185]) );
  AND U3752 ( .A(n1035), .B(n3751), .Z(n3749) );
  XOR U3753 ( .A(creg[185]), .B(mod_mult_o[185]), .Z(n3751) );
  XNOR U3754 ( .A(n3752), .B(n3753), .Z(o[184]) );
  AND U3755 ( .A(n1035), .B(n3754), .Z(n3752) );
  XOR U3756 ( .A(creg[184]), .B(mod_mult_o[184]), .Z(n3754) );
  XNOR U3757 ( .A(n3755), .B(n3756), .Z(o[183]) );
  AND U3758 ( .A(n1035), .B(n3757), .Z(n3755) );
  XOR U3759 ( .A(creg[183]), .B(mod_mult_o[183]), .Z(n3757) );
  XNOR U3760 ( .A(n3758), .B(n3759), .Z(o[182]) );
  AND U3761 ( .A(n1035), .B(n3760), .Z(n3758) );
  XOR U3762 ( .A(creg[182]), .B(mod_mult_o[182]), .Z(n3760) );
  XNOR U3763 ( .A(n3761), .B(n3762), .Z(o[181]) );
  AND U3764 ( .A(n1035), .B(n3763), .Z(n3761) );
  XOR U3765 ( .A(creg[181]), .B(mod_mult_o[181]), .Z(n3763) );
  XNOR U3766 ( .A(n3764), .B(n3765), .Z(o[180]) );
  AND U3767 ( .A(n1035), .B(n3766), .Z(n3764) );
  XOR U3768 ( .A(creg[180]), .B(mod_mult_o[180]), .Z(n3766) );
  XNOR U3769 ( .A(n3767), .B(n3768), .Z(o[17]) );
  AND U3770 ( .A(n1035), .B(n3769), .Z(n3767) );
  XOR U3771 ( .A(creg[17]), .B(mod_mult_o[17]), .Z(n3769) );
  XNOR U3772 ( .A(n3770), .B(n3771), .Z(o[179]) );
  AND U3773 ( .A(n1035), .B(n3772), .Z(n3770) );
  XOR U3774 ( .A(creg[179]), .B(mod_mult_o[179]), .Z(n3772) );
  XNOR U3775 ( .A(n3773), .B(n3774), .Z(o[178]) );
  AND U3776 ( .A(n1035), .B(n3775), .Z(n3773) );
  XOR U3777 ( .A(creg[178]), .B(mod_mult_o[178]), .Z(n3775) );
  XNOR U3778 ( .A(n3776), .B(n3777), .Z(o[177]) );
  AND U3779 ( .A(n1035), .B(n3778), .Z(n3776) );
  XOR U3780 ( .A(creg[177]), .B(mod_mult_o[177]), .Z(n3778) );
  XNOR U3781 ( .A(n3779), .B(n3780), .Z(o[176]) );
  AND U3782 ( .A(n1035), .B(n3781), .Z(n3779) );
  XOR U3783 ( .A(creg[176]), .B(mod_mult_o[176]), .Z(n3781) );
  XNOR U3784 ( .A(n3782), .B(n3783), .Z(o[175]) );
  AND U3785 ( .A(n1035), .B(n3784), .Z(n3782) );
  XOR U3786 ( .A(creg[175]), .B(mod_mult_o[175]), .Z(n3784) );
  XNOR U3787 ( .A(n3785), .B(n3786), .Z(o[174]) );
  AND U3788 ( .A(n1035), .B(n3787), .Z(n3785) );
  XOR U3789 ( .A(creg[174]), .B(mod_mult_o[174]), .Z(n3787) );
  XNOR U3790 ( .A(n3788), .B(n3789), .Z(o[173]) );
  AND U3791 ( .A(n1035), .B(n3790), .Z(n3788) );
  XOR U3792 ( .A(creg[173]), .B(mod_mult_o[173]), .Z(n3790) );
  XNOR U3793 ( .A(n3791), .B(n3792), .Z(o[172]) );
  AND U3794 ( .A(n1035), .B(n3793), .Z(n3791) );
  XOR U3795 ( .A(creg[172]), .B(mod_mult_o[172]), .Z(n3793) );
  XNOR U3796 ( .A(n3794), .B(n3795), .Z(o[171]) );
  AND U3797 ( .A(n1035), .B(n3796), .Z(n3794) );
  XOR U3798 ( .A(creg[171]), .B(mod_mult_o[171]), .Z(n3796) );
  XNOR U3799 ( .A(n3797), .B(n3798), .Z(o[170]) );
  AND U3800 ( .A(n1035), .B(n3799), .Z(n3797) );
  XOR U3801 ( .A(creg[170]), .B(mod_mult_o[170]), .Z(n3799) );
  XNOR U3802 ( .A(n3800), .B(n3801), .Z(o[16]) );
  AND U3803 ( .A(n1035), .B(n3802), .Z(n3800) );
  XOR U3804 ( .A(creg[16]), .B(mod_mult_o[16]), .Z(n3802) );
  XNOR U3805 ( .A(n3803), .B(n3804), .Z(o[169]) );
  AND U3806 ( .A(n1035), .B(n3805), .Z(n3803) );
  XOR U3807 ( .A(creg[169]), .B(mod_mult_o[169]), .Z(n3805) );
  XNOR U3808 ( .A(n3806), .B(n3807), .Z(o[168]) );
  AND U3809 ( .A(n1035), .B(n3808), .Z(n3806) );
  XOR U3810 ( .A(creg[168]), .B(mod_mult_o[168]), .Z(n3808) );
  XNOR U3811 ( .A(n3809), .B(n3810), .Z(o[167]) );
  AND U3812 ( .A(n1035), .B(n3811), .Z(n3809) );
  XOR U3813 ( .A(creg[167]), .B(mod_mult_o[167]), .Z(n3811) );
  XNOR U3814 ( .A(n3812), .B(n3813), .Z(o[166]) );
  AND U3815 ( .A(n1035), .B(n3814), .Z(n3812) );
  XOR U3816 ( .A(creg[166]), .B(mod_mult_o[166]), .Z(n3814) );
  XNOR U3817 ( .A(n3815), .B(n3816), .Z(o[165]) );
  AND U3818 ( .A(n1035), .B(n3817), .Z(n3815) );
  XOR U3819 ( .A(creg[165]), .B(mod_mult_o[165]), .Z(n3817) );
  XNOR U3820 ( .A(n3818), .B(n3819), .Z(o[164]) );
  AND U3821 ( .A(n1035), .B(n3820), .Z(n3818) );
  XOR U3822 ( .A(creg[164]), .B(mod_mult_o[164]), .Z(n3820) );
  XNOR U3823 ( .A(n3821), .B(n3822), .Z(o[163]) );
  AND U3824 ( .A(n1035), .B(n3823), .Z(n3821) );
  XOR U3825 ( .A(creg[163]), .B(mod_mult_o[163]), .Z(n3823) );
  XNOR U3826 ( .A(n3824), .B(n3825), .Z(o[162]) );
  AND U3827 ( .A(n1035), .B(n3826), .Z(n3824) );
  XOR U3828 ( .A(creg[162]), .B(mod_mult_o[162]), .Z(n3826) );
  XNOR U3829 ( .A(n3827), .B(n3828), .Z(o[161]) );
  AND U3830 ( .A(n1035), .B(n3829), .Z(n3827) );
  XOR U3831 ( .A(creg[161]), .B(mod_mult_o[161]), .Z(n3829) );
  XNOR U3832 ( .A(n3830), .B(n3831), .Z(o[160]) );
  AND U3833 ( .A(n1035), .B(n3832), .Z(n3830) );
  XOR U3834 ( .A(creg[160]), .B(mod_mult_o[160]), .Z(n3832) );
  XNOR U3835 ( .A(n3833), .B(n3834), .Z(o[15]) );
  AND U3836 ( .A(n1035), .B(n3835), .Z(n3833) );
  XOR U3837 ( .A(creg[15]), .B(mod_mult_o[15]), .Z(n3835) );
  XNOR U3838 ( .A(n3836), .B(n3837), .Z(o[159]) );
  AND U3839 ( .A(n1035), .B(n3838), .Z(n3836) );
  XOR U3840 ( .A(creg[159]), .B(mod_mult_o[159]), .Z(n3838) );
  XNOR U3841 ( .A(n3839), .B(n3840), .Z(o[158]) );
  AND U3842 ( .A(n1035), .B(n3841), .Z(n3839) );
  XOR U3843 ( .A(creg[158]), .B(mod_mult_o[158]), .Z(n3841) );
  XNOR U3844 ( .A(n3842), .B(n3843), .Z(o[157]) );
  AND U3845 ( .A(n1035), .B(n3844), .Z(n3842) );
  XOR U3846 ( .A(creg[157]), .B(mod_mult_o[157]), .Z(n3844) );
  XNOR U3847 ( .A(n3845), .B(n3846), .Z(o[156]) );
  AND U3848 ( .A(n1035), .B(n3847), .Z(n3845) );
  XOR U3849 ( .A(creg[156]), .B(mod_mult_o[156]), .Z(n3847) );
  XNOR U3850 ( .A(n3848), .B(n3849), .Z(o[155]) );
  AND U3851 ( .A(n1035), .B(n3850), .Z(n3848) );
  XOR U3852 ( .A(creg[155]), .B(mod_mult_o[155]), .Z(n3850) );
  XNOR U3853 ( .A(n3851), .B(n3852), .Z(o[154]) );
  AND U3854 ( .A(n1035), .B(n3853), .Z(n3851) );
  XOR U3855 ( .A(creg[154]), .B(mod_mult_o[154]), .Z(n3853) );
  XNOR U3856 ( .A(n3854), .B(n3855), .Z(o[153]) );
  AND U3857 ( .A(n1035), .B(n3856), .Z(n3854) );
  XOR U3858 ( .A(creg[153]), .B(mod_mult_o[153]), .Z(n3856) );
  XNOR U3859 ( .A(n3857), .B(n3858), .Z(o[152]) );
  AND U3860 ( .A(n1035), .B(n3859), .Z(n3857) );
  XOR U3861 ( .A(creg[152]), .B(mod_mult_o[152]), .Z(n3859) );
  XNOR U3862 ( .A(n3860), .B(n3861), .Z(o[151]) );
  AND U3863 ( .A(n1035), .B(n3862), .Z(n3860) );
  XOR U3864 ( .A(creg[151]), .B(mod_mult_o[151]), .Z(n3862) );
  XNOR U3865 ( .A(n3863), .B(n3864), .Z(o[150]) );
  AND U3866 ( .A(n1035), .B(n3865), .Z(n3863) );
  XOR U3867 ( .A(creg[150]), .B(mod_mult_o[150]), .Z(n3865) );
  XNOR U3868 ( .A(n3866), .B(n3867), .Z(o[14]) );
  AND U3869 ( .A(n1035), .B(n3868), .Z(n3866) );
  XOR U3870 ( .A(creg[14]), .B(mod_mult_o[14]), .Z(n3868) );
  XNOR U3871 ( .A(n3869), .B(n3870), .Z(o[149]) );
  AND U3872 ( .A(n1035), .B(n3871), .Z(n3869) );
  XOR U3873 ( .A(creg[149]), .B(mod_mult_o[149]), .Z(n3871) );
  XNOR U3874 ( .A(n3872), .B(n3873), .Z(o[148]) );
  AND U3875 ( .A(n1035), .B(n3874), .Z(n3872) );
  XOR U3876 ( .A(creg[148]), .B(mod_mult_o[148]), .Z(n3874) );
  XNOR U3877 ( .A(n3875), .B(n3876), .Z(o[147]) );
  AND U3878 ( .A(n1035), .B(n3877), .Z(n3875) );
  XOR U3879 ( .A(creg[147]), .B(mod_mult_o[147]), .Z(n3877) );
  XNOR U3880 ( .A(n3878), .B(n3879), .Z(o[146]) );
  AND U3881 ( .A(n1035), .B(n3880), .Z(n3878) );
  XOR U3882 ( .A(creg[146]), .B(mod_mult_o[146]), .Z(n3880) );
  XNOR U3883 ( .A(n3881), .B(n3882), .Z(o[145]) );
  AND U3884 ( .A(n1035), .B(n3883), .Z(n3881) );
  XOR U3885 ( .A(creg[145]), .B(mod_mult_o[145]), .Z(n3883) );
  XNOR U3886 ( .A(n3884), .B(n3885), .Z(o[144]) );
  AND U3887 ( .A(n1035), .B(n3886), .Z(n3884) );
  XOR U3888 ( .A(creg[144]), .B(mod_mult_o[144]), .Z(n3886) );
  XNOR U3889 ( .A(n3887), .B(n3888), .Z(o[143]) );
  AND U3890 ( .A(n1035), .B(n3889), .Z(n3887) );
  XOR U3891 ( .A(creg[143]), .B(mod_mult_o[143]), .Z(n3889) );
  XNOR U3892 ( .A(n3890), .B(n3891), .Z(o[142]) );
  AND U3893 ( .A(n1035), .B(n3892), .Z(n3890) );
  XOR U3894 ( .A(creg[142]), .B(mod_mult_o[142]), .Z(n3892) );
  XNOR U3895 ( .A(n3893), .B(n3894), .Z(o[141]) );
  AND U3896 ( .A(n1035), .B(n3895), .Z(n3893) );
  XOR U3897 ( .A(creg[141]), .B(mod_mult_o[141]), .Z(n3895) );
  XNOR U3898 ( .A(n3896), .B(n3897), .Z(o[140]) );
  AND U3899 ( .A(n1035), .B(n3898), .Z(n3896) );
  XOR U3900 ( .A(creg[140]), .B(mod_mult_o[140]), .Z(n3898) );
  XNOR U3901 ( .A(n3899), .B(n3900), .Z(o[13]) );
  AND U3902 ( .A(n1035), .B(n3901), .Z(n3899) );
  XOR U3903 ( .A(creg[13]), .B(mod_mult_o[13]), .Z(n3901) );
  XNOR U3904 ( .A(n3902), .B(n3903), .Z(o[139]) );
  AND U3905 ( .A(n1035), .B(n3904), .Z(n3902) );
  XOR U3906 ( .A(creg[139]), .B(mod_mult_o[139]), .Z(n3904) );
  XNOR U3907 ( .A(n3905), .B(n3906), .Z(o[138]) );
  AND U3908 ( .A(n1035), .B(n3907), .Z(n3905) );
  XOR U3909 ( .A(creg[138]), .B(mod_mult_o[138]), .Z(n3907) );
  XNOR U3910 ( .A(n3908), .B(n3909), .Z(o[137]) );
  AND U3911 ( .A(n1035), .B(n3910), .Z(n3908) );
  XOR U3912 ( .A(creg[137]), .B(mod_mult_o[137]), .Z(n3910) );
  XNOR U3913 ( .A(n3911), .B(n3912), .Z(o[136]) );
  AND U3914 ( .A(n1035), .B(n3913), .Z(n3911) );
  XOR U3915 ( .A(creg[136]), .B(mod_mult_o[136]), .Z(n3913) );
  XNOR U3916 ( .A(n3914), .B(n3915), .Z(o[135]) );
  AND U3917 ( .A(n1035), .B(n3916), .Z(n3914) );
  XOR U3918 ( .A(creg[135]), .B(mod_mult_o[135]), .Z(n3916) );
  XNOR U3919 ( .A(n3917), .B(n3918), .Z(o[134]) );
  AND U3920 ( .A(n1035), .B(n3919), .Z(n3917) );
  XOR U3921 ( .A(creg[134]), .B(mod_mult_o[134]), .Z(n3919) );
  XNOR U3922 ( .A(n3920), .B(n3921), .Z(o[133]) );
  AND U3923 ( .A(n1035), .B(n3922), .Z(n3920) );
  XOR U3924 ( .A(creg[133]), .B(mod_mult_o[133]), .Z(n3922) );
  XNOR U3925 ( .A(n3923), .B(n3924), .Z(o[132]) );
  AND U3926 ( .A(n1035), .B(n3925), .Z(n3923) );
  XOR U3927 ( .A(creg[132]), .B(mod_mult_o[132]), .Z(n3925) );
  XNOR U3928 ( .A(n3926), .B(n3927), .Z(o[131]) );
  AND U3929 ( .A(n1035), .B(n3928), .Z(n3926) );
  XOR U3930 ( .A(creg[131]), .B(mod_mult_o[131]), .Z(n3928) );
  XNOR U3931 ( .A(n3929), .B(n3930), .Z(o[130]) );
  AND U3932 ( .A(n1035), .B(n3931), .Z(n3929) );
  XOR U3933 ( .A(creg[130]), .B(mod_mult_o[130]), .Z(n3931) );
  XNOR U3934 ( .A(n3932), .B(n3933), .Z(o[12]) );
  AND U3935 ( .A(n1035), .B(n3934), .Z(n3932) );
  XOR U3936 ( .A(creg[12]), .B(mod_mult_o[12]), .Z(n3934) );
  XNOR U3937 ( .A(n3935), .B(n3936), .Z(o[129]) );
  AND U3938 ( .A(n1035), .B(n3937), .Z(n3935) );
  XOR U3939 ( .A(creg[129]), .B(mod_mult_o[129]), .Z(n3937) );
  XNOR U3940 ( .A(n3938), .B(n3939), .Z(o[128]) );
  AND U3941 ( .A(n1035), .B(n3940), .Z(n3938) );
  XOR U3942 ( .A(creg[128]), .B(mod_mult_o[128]), .Z(n3940) );
  XNOR U3943 ( .A(n3941), .B(n3942), .Z(o[127]) );
  AND U3944 ( .A(n1035), .B(n3943), .Z(n3941) );
  XOR U3945 ( .A(creg[127]), .B(mod_mult_o[127]), .Z(n3943) );
  XNOR U3946 ( .A(n3944), .B(n3945), .Z(o[126]) );
  AND U3947 ( .A(n1035), .B(n3946), .Z(n3944) );
  XOR U3948 ( .A(creg[126]), .B(mod_mult_o[126]), .Z(n3946) );
  XNOR U3949 ( .A(n3947), .B(n3948), .Z(o[125]) );
  AND U3950 ( .A(n1035), .B(n3949), .Z(n3947) );
  XOR U3951 ( .A(creg[125]), .B(mod_mult_o[125]), .Z(n3949) );
  XNOR U3952 ( .A(n3950), .B(n3951), .Z(o[124]) );
  AND U3953 ( .A(n1035), .B(n3952), .Z(n3950) );
  XOR U3954 ( .A(creg[124]), .B(mod_mult_o[124]), .Z(n3952) );
  XNOR U3955 ( .A(n3953), .B(n3954), .Z(o[123]) );
  AND U3956 ( .A(n1035), .B(n3955), .Z(n3953) );
  XOR U3957 ( .A(creg[123]), .B(mod_mult_o[123]), .Z(n3955) );
  XNOR U3958 ( .A(n3956), .B(n3957), .Z(o[122]) );
  AND U3959 ( .A(n1035), .B(n3958), .Z(n3956) );
  XOR U3960 ( .A(creg[122]), .B(mod_mult_o[122]), .Z(n3958) );
  XNOR U3961 ( .A(n3959), .B(n3960), .Z(o[121]) );
  AND U3962 ( .A(n1035), .B(n3961), .Z(n3959) );
  XOR U3963 ( .A(creg[121]), .B(mod_mult_o[121]), .Z(n3961) );
  XNOR U3964 ( .A(n3962), .B(n3963), .Z(o[120]) );
  AND U3965 ( .A(n1035), .B(n3964), .Z(n3962) );
  XOR U3966 ( .A(creg[120]), .B(mod_mult_o[120]), .Z(n3964) );
  XNOR U3967 ( .A(n3965), .B(n3966), .Z(o[11]) );
  AND U3968 ( .A(n1035), .B(n3967), .Z(n3965) );
  XOR U3969 ( .A(creg[11]), .B(mod_mult_o[11]), .Z(n3967) );
  XNOR U3970 ( .A(n3968), .B(n3969), .Z(o[119]) );
  AND U3971 ( .A(n1035), .B(n3970), .Z(n3968) );
  XOR U3972 ( .A(creg[119]), .B(mod_mult_o[119]), .Z(n3970) );
  XNOR U3973 ( .A(n3971), .B(n3972), .Z(o[118]) );
  AND U3974 ( .A(n1035), .B(n3973), .Z(n3971) );
  XOR U3975 ( .A(creg[118]), .B(mod_mult_o[118]), .Z(n3973) );
  XNOR U3976 ( .A(n3974), .B(n3975), .Z(o[117]) );
  AND U3977 ( .A(n1035), .B(n3976), .Z(n3974) );
  XOR U3978 ( .A(creg[117]), .B(mod_mult_o[117]), .Z(n3976) );
  XNOR U3979 ( .A(n3977), .B(n3978), .Z(o[116]) );
  AND U3980 ( .A(n1035), .B(n3979), .Z(n3977) );
  XOR U3981 ( .A(creg[116]), .B(mod_mult_o[116]), .Z(n3979) );
  XNOR U3982 ( .A(n3980), .B(n3981), .Z(o[115]) );
  AND U3983 ( .A(n1035), .B(n3982), .Z(n3980) );
  XOR U3984 ( .A(creg[115]), .B(mod_mult_o[115]), .Z(n3982) );
  XNOR U3985 ( .A(n3983), .B(n3984), .Z(o[114]) );
  AND U3986 ( .A(n1035), .B(n3985), .Z(n3983) );
  XOR U3987 ( .A(creg[114]), .B(mod_mult_o[114]), .Z(n3985) );
  XNOR U3988 ( .A(n3986), .B(n3987), .Z(o[113]) );
  AND U3989 ( .A(n1035), .B(n3988), .Z(n3986) );
  XOR U3990 ( .A(creg[113]), .B(mod_mult_o[113]), .Z(n3988) );
  XNOR U3991 ( .A(n3989), .B(n3990), .Z(o[112]) );
  AND U3992 ( .A(n1035), .B(n3991), .Z(n3989) );
  XOR U3993 ( .A(creg[112]), .B(mod_mult_o[112]), .Z(n3991) );
  XNOR U3994 ( .A(n3992), .B(n3993), .Z(o[111]) );
  AND U3995 ( .A(n1035), .B(n3994), .Z(n3992) );
  XOR U3996 ( .A(creg[111]), .B(mod_mult_o[111]), .Z(n3994) );
  XNOR U3997 ( .A(n3995), .B(n3996), .Z(o[110]) );
  AND U3998 ( .A(n1035), .B(n3997), .Z(n3995) );
  XOR U3999 ( .A(creg[110]), .B(mod_mult_o[110]), .Z(n3997) );
  XNOR U4000 ( .A(n3998), .B(n3999), .Z(o[10]) );
  AND U4001 ( .A(n1035), .B(n4000), .Z(n3998) );
  XOR U4002 ( .A(creg[10]), .B(mod_mult_o[10]), .Z(n4000) );
  XNOR U4003 ( .A(n4001), .B(n4002), .Z(o[109]) );
  AND U4004 ( .A(n1035), .B(n4003), .Z(n4001) );
  XOR U4005 ( .A(creg[109]), .B(mod_mult_o[109]), .Z(n4003) );
  XNOR U4006 ( .A(n4004), .B(n4005), .Z(o[108]) );
  AND U4007 ( .A(n1035), .B(n4006), .Z(n4004) );
  XOR U4008 ( .A(creg[108]), .B(mod_mult_o[108]), .Z(n4006) );
  XNOR U4009 ( .A(n4007), .B(n4008), .Z(o[107]) );
  AND U4010 ( .A(n1035), .B(n4009), .Z(n4007) );
  XOR U4011 ( .A(creg[107]), .B(mod_mult_o[107]), .Z(n4009) );
  XNOR U4012 ( .A(n4010), .B(n4011), .Z(o[106]) );
  AND U4013 ( .A(n1035), .B(n4012), .Z(n4010) );
  XOR U4014 ( .A(creg[106]), .B(mod_mult_o[106]), .Z(n4012) );
  XNOR U4015 ( .A(n4013), .B(n4014), .Z(o[105]) );
  AND U4016 ( .A(n1035), .B(n4015), .Z(n4013) );
  XOR U4017 ( .A(creg[105]), .B(mod_mult_o[105]), .Z(n4015) );
  XNOR U4018 ( .A(n4016), .B(n4017), .Z(o[104]) );
  AND U4019 ( .A(n1035), .B(n4018), .Z(n4016) );
  XOR U4020 ( .A(creg[104]), .B(mod_mult_o[104]), .Z(n4018) );
  XNOR U4021 ( .A(n4019), .B(n4020), .Z(o[103]) );
  AND U4022 ( .A(n1035), .B(n4021), .Z(n4019) );
  XOR U4023 ( .A(creg[103]), .B(mod_mult_o[103]), .Z(n4021) );
  XNOR U4024 ( .A(n4022), .B(n4023), .Z(o[102]) );
  AND U4025 ( .A(n1035), .B(n4024), .Z(n4022) );
  XOR U4026 ( .A(creg[102]), .B(mod_mult_o[102]), .Z(n4024) );
  XNOR U4027 ( .A(n4025), .B(n4026), .Z(o[1023]) );
  AND U4028 ( .A(n1035), .B(n4027), .Z(n4025) );
  XOR U4029 ( .A(creg[1023]), .B(mod_mult_o[1023]), .Z(n4027) );
  XNOR U4030 ( .A(n4028), .B(n4029), .Z(o[1022]) );
  AND U4031 ( .A(n1035), .B(n4030), .Z(n4028) );
  XOR U4032 ( .A(creg[1022]), .B(mod_mult_o[1022]), .Z(n4030) );
  XNOR U4033 ( .A(n4031), .B(n4032), .Z(o[1021]) );
  AND U4034 ( .A(n1035), .B(n4033), .Z(n4031) );
  XOR U4035 ( .A(creg[1021]), .B(mod_mult_o[1021]), .Z(n4033) );
  XNOR U4036 ( .A(n4034), .B(n4035), .Z(o[1020]) );
  AND U4037 ( .A(n1035), .B(n4036), .Z(n4034) );
  XOR U4038 ( .A(creg[1020]), .B(mod_mult_o[1020]), .Z(n4036) );
  XNOR U4039 ( .A(n4037), .B(n4038), .Z(o[101]) );
  AND U4040 ( .A(n1035), .B(n4039), .Z(n4037) );
  XOR U4041 ( .A(creg[101]), .B(mod_mult_o[101]), .Z(n4039) );
  XNOR U4042 ( .A(n4040), .B(n4041), .Z(o[1019]) );
  AND U4043 ( .A(n1035), .B(n4042), .Z(n4040) );
  XOR U4044 ( .A(creg[1019]), .B(mod_mult_o[1019]), .Z(n4042) );
  XNOR U4045 ( .A(n4043), .B(n4044), .Z(o[1018]) );
  AND U4046 ( .A(n1035), .B(n4045), .Z(n4043) );
  XOR U4047 ( .A(creg[1018]), .B(mod_mult_o[1018]), .Z(n4045) );
  XNOR U4048 ( .A(n4046), .B(n4047), .Z(o[1017]) );
  AND U4049 ( .A(n1035), .B(n4048), .Z(n4046) );
  XOR U4050 ( .A(creg[1017]), .B(mod_mult_o[1017]), .Z(n4048) );
  XNOR U4051 ( .A(n4049), .B(n4050), .Z(o[1016]) );
  AND U4052 ( .A(n1035), .B(n4051), .Z(n4049) );
  XOR U4053 ( .A(creg[1016]), .B(mod_mult_o[1016]), .Z(n4051) );
  XNOR U4054 ( .A(n4052), .B(n4053), .Z(o[1015]) );
  AND U4055 ( .A(n1035), .B(n4054), .Z(n4052) );
  XOR U4056 ( .A(creg[1015]), .B(mod_mult_o[1015]), .Z(n4054) );
  XNOR U4057 ( .A(n4055), .B(n4056), .Z(o[1014]) );
  AND U4058 ( .A(n1035), .B(n4057), .Z(n4055) );
  XOR U4059 ( .A(creg[1014]), .B(mod_mult_o[1014]), .Z(n4057) );
  XNOR U4060 ( .A(n4058), .B(n4059), .Z(o[1013]) );
  AND U4061 ( .A(n1035), .B(n4060), .Z(n4058) );
  XOR U4062 ( .A(creg[1013]), .B(mod_mult_o[1013]), .Z(n4060) );
  XNOR U4063 ( .A(n4061), .B(n4062), .Z(o[1012]) );
  AND U4064 ( .A(n1035), .B(n4063), .Z(n4061) );
  XOR U4065 ( .A(creg[1012]), .B(mod_mult_o[1012]), .Z(n4063) );
  XNOR U4066 ( .A(n4064), .B(n4065), .Z(o[1011]) );
  AND U4067 ( .A(n1035), .B(n4066), .Z(n4064) );
  XOR U4068 ( .A(creg[1011]), .B(mod_mult_o[1011]), .Z(n4066) );
  XNOR U4069 ( .A(n4067), .B(n4068), .Z(o[1010]) );
  AND U4070 ( .A(n1035), .B(n4069), .Z(n4067) );
  XOR U4071 ( .A(creg[1010]), .B(mod_mult_o[1010]), .Z(n4069) );
  XNOR U4072 ( .A(n4070), .B(n4071), .Z(o[100]) );
  AND U4073 ( .A(n1035), .B(n4072), .Z(n4070) );
  XOR U4074 ( .A(creg[100]), .B(mod_mult_o[100]), .Z(n4072) );
  XNOR U4075 ( .A(n4073), .B(n4074), .Z(o[1009]) );
  AND U4076 ( .A(n1035), .B(n4075), .Z(n4073) );
  XOR U4077 ( .A(creg[1009]), .B(mod_mult_o[1009]), .Z(n4075) );
  XNOR U4078 ( .A(n4076), .B(n4077), .Z(o[1008]) );
  AND U4079 ( .A(n1035), .B(n4078), .Z(n4076) );
  XOR U4080 ( .A(creg[1008]), .B(mod_mult_o[1008]), .Z(n4078) );
  XNOR U4081 ( .A(n4079), .B(n4080), .Z(o[1007]) );
  AND U4082 ( .A(n1035), .B(n4081), .Z(n4079) );
  XOR U4083 ( .A(creg[1007]), .B(mod_mult_o[1007]), .Z(n4081) );
  XNOR U4084 ( .A(n4082), .B(n4083), .Z(o[1006]) );
  AND U4085 ( .A(n1035), .B(n4084), .Z(n4082) );
  XOR U4086 ( .A(creg[1006]), .B(mod_mult_o[1006]), .Z(n4084) );
  XNOR U4087 ( .A(n4085), .B(n4086), .Z(o[1005]) );
  AND U4088 ( .A(n1035), .B(n4087), .Z(n4085) );
  XOR U4089 ( .A(creg[1005]), .B(mod_mult_o[1005]), .Z(n4087) );
  XNOR U4090 ( .A(n4088), .B(n4089), .Z(o[1004]) );
  AND U4091 ( .A(n1035), .B(n4090), .Z(n4088) );
  XOR U4092 ( .A(creg[1004]), .B(mod_mult_o[1004]), .Z(n4090) );
  XNOR U4093 ( .A(n4091), .B(n4092), .Z(o[1003]) );
  AND U4094 ( .A(n1035), .B(n4093), .Z(n4091) );
  XOR U4095 ( .A(creg[1003]), .B(mod_mult_o[1003]), .Z(n4093) );
  XNOR U4096 ( .A(n4094), .B(n4095), .Z(o[1002]) );
  AND U4097 ( .A(n1035), .B(n4096), .Z(n4094) );
  XOR U4098 ( .A(creg[1002]), .B(mod_mult_o[1002]), .Z(n4096) );
  XNOR U4099 ( .A(n4097), .B(n4098), .Z(o[1001]) );
  AND U4100 ( .A(n1035), .B(n4099), .Z(n4097) );
  XOR U4101 ( .A(creg[1001]), .B(mod_mult_o[1001]), .Z(n4099) );
  XNOR U4102 ( .A(n4100), .B(n4101), .Z(o[1000]) );
  AND U4103 ( .A(n1035), .B(n4102), .Z(n4100) );
  XOR U4104 ( .A(creg[1000]), .B(mod_mult_o[1000]), .Z(n4102) );
  XOR U4105 ( .A(n4103), .B(mod_mult_o[0]), .Z(o[0]) );
  AND U4106 ( .A(n1035), .B(n4104), .Z(n4103) );
  XOR U4107 ( .A(creg[0]), .B(mod_mult_o[0]), .Z(n4104) );
  NAND U4108 ( .A(n4105), .B(n4106), .Z(n1035) );
  NANDN U4109 ( .B(mul_pow), .A(first_one), .Z(n4106) );
  NAND U4110 ( .A(first_one), .B(ein[1023]), .Z(n4105) );
  XOR U4111 ( .A(start_in[1023]), .B(mul_pow), .Z(n8) );
  NANDN U4112 ( .B(first_one), .A(n4107), .Z(n6) );
  NAND U4113 ( .A(n4108), .B(start_in[1023]), .Z(n4107) );
  AND U4114 ( .A(ein[1023]), .B(mul_pow), .Z(n4108) );
  XNOR U4115 ( .A(n4109), .B(n4110), .Z(\modmult_1/zout[0][1024] ) );
  XOR U4116 ( .A(n4111), .B(n4112), .Z(n4110) );
  ANDN U4117 ( .A(n4113), .B(n4114), .Z(n4111) );
  XNOR U4118 ( .A(n4115), .B(n4116), .Z(n4113) );
  IV U4119 ( .A(n1034), .Z(mod_mult_o[9]) );
  XOR U4120 ( .A(n4117), .B(n4118), .Z(n1034) );
  IV U4121 ( .A(n1038), .Z(mod_mult_o[99]) );
  XOR U4122 ( .A(n4119), .B(n4120), .Z(n1038) );
  IV U4123 ( .A(n1041), .Z(mod_mult_o[999]) );
  XOR U4124 ( .A(n4121), .B(n4122), .Z(n1041) );
  IV U4125 ( .A(n1044), .Z(mod_mult_o[998]) );
  XOR U4126 ( .A(n4123), .B(n4124), .Z(n1044) );
  IV U4127 ( .A(n1047), .Z(mod_mult_o[997]) );
  XOR U4128 ( .A(n4125), .B(n4126), .Z(n1047) );
  IV U4129 ( .A(n1050), .Z(mod_mult_o[996]) );
  XOR U4130 ( .A(n4127), .B(n4128), .Z(n1050) );
  IV U4131 ( .A(n1053), .Z(mod_mult_o[995]) );
  XOR U4132 ( .A(n4129), .B(n4130), .Z(n1053) );
  IV U4133 ( .A(n1056), .Z(mod_mult_o[994]) );
  XOR U4134 ( .A(n4131), .B(n4132), .Z(n1056) );
  IV U4135 ( .A(n1059), .Z(mod_mult_o[993]) );
  XOR U4136 ( .A(n4133), .B(n4134), .Z(n1059) );
  IV U4137 ( .A(n1062), .Z(mod_mult_o[992]) );
  XOR U4138 ( .A(n4135), .B(n4136), .Z(n1062) );
  IV U4139 ( .A(n1065), .Z(mod_mult_o[991]) );
  XOR U4140 ( .A(n4137), .B(n4138), .Z(n1065) );
  IV U4141 ( .A(n1068), .Z(mod_mult_o[990]) );
  XOR U4142 ( .A(n4139), .B(n4140), .Z(n1068) );
  IV U4143 ( .A(n1071), .Z(mod_mult_o[98]) );
  XOR U4144 ( .A(n4141), .B(n4142), .Z(n1071) );
  IV U4145 ( .A(n1074), .Z(mod_mult_o[989]) );
  XOR U4146 ( .A(n4143), .B(n4144), .Z(n1074) );
  IV U4147 ( .A(n1077), .Z(mod_mult_o[988]) );
  XOR U4148 ( .A(n4145), .B(n4146), .Z(n1077) );
  IV U4149 ( .A(n1080), .Z(mod_mult_o[987]) );
  XOR U4150 ( .A(n4147), .B(n4148), .Z(n1080) );
  IV U4151 ( .A(n1083), .Z(mod_mult_o[986]) );
  XOR U4152 ( .A(n4149), .B(n4150), .Z(n1083) );
  IV U4153 ( .A(n1086), .Z(mod_mult_o[985]) );
  XOR U4154 ( .A(n4151), .B(n4152), .Z(n1086) );
  IV U4155 ( .A(n1089), .Z(mod_mult_o[984]) );
  XOR U4156 ( .A(n4153), .B(n4154), .Z(n1089) );
  IV U4157 ( .A(n1092), .Z(mod_mult_o[983]) );
  XOR U4158 ( .A(n4155), .B(n4156), .Z(n1092) );
  IV U4159 ( .A(n1095), .Z(mod_mult_o[982]) );
  XOR U4160 ( .A(n4157), .B(n4158), .Z(n1095) );
  IV U4161 ( .A(n1098), .Z(mod_mult_o[981]) );
  XOR U4162 ( .A(n4159), .B(n4160), .Z(n1098) );
  IV U4163 ( .A(n1101), .Z(mod_mult_o[980]) );
  XOR U4164 ( .A(n4161), .B(n4162), .Z(n1101) );
  IV U4165 ( .A(n1104), .Z(mod_mult_o[97]) );
  XOR U4166 ( .A(n4163), .B(n4164), .Z(n1104) );
  IV U4167 ( .A(n1107), .Z(mod_mult_o[979]) );
  XOR U4168 ( .A(n4165), .B(n4166), .Z(n1107) );
  IV U4169 ( .A(n1110), .Z(mod_mult_o[978]) );
  XOR U4170 ( .A(n4167), .B(n4168), .Z(n1110) );
  IV U4171 ( .A(n1113), .Z(mod_mult_o[977]) );
  XOR U4172 ( .A(n4169), .B(n4170), .Z(n1113) );
  IV U4173 ( .A(n1116), .Z(mod_mult_o[976]) );
  XOR U4174 ( .A(n4171), .B(n4172), .Z(n1116) );
  IV U4175 ( .A(n1119), .Z(mod_mult_o[975]) );
  XOR U4176 ( .A(n4173), .B(n4174), .Z(n1119) );
  IV U4177 ( .A(n1122), .Z(mod_mult_o[974]) );
  XOR U4178 ( .A(n4175), .B(n4176), .Z(n1122) );
  IV U4179 ( .A(n1125), .Z(mod_mult_o[973]) );
  XOR U4180 ( .A(n4177), .B(n4178), .Z(n1125) );
  IV U4181 ( .A(n1128), .Z(mod_mult_o[972]) );
  XOR U4182 ( .A(n4179), .B(n4180), .Z(n1128) );
  IV U4183 ( .A(n1131), .Z(mod_mult_o[971]) );
  XOR U4184 ( .A(n4181), .B(n4182), .Z(n1131) );
  IV U4185 ( .A(n1134), .Z(mod_mult_o[970]) );
  XOR U4186 ( .A(n4183), .B(n4184), .Z(n1134) );
  IV U4187 ( .A(n1137), .Z(mod_mult_o[96]) );
  XOR U4188 ( .A(n4185), .B(n4186), .Z(n1137) );
  IV U4189 ( .A(n1140), .Z(mod_mult_o[969]) );
  XOR U4190 ( .A(n4187), .B(n4188), .Z(n1140) );
  IV U4191 ( .A(n1143), .Z(mod_mult_o[968]) );
  XOR U4192 ( .A(n4189), .B(n4190), .Z(n1143) );
  IV U4193 ( .A(n1146), .Z(mod_mult_o[967]) );
  XOR U4194 ( .A(n4191), .B(n4192), .Z(n1146) );
  IV U4195 ( .A(n1149), .Z(mod_mult_o[966]) );
  XOR U4196 ( .A(n4193), .B(n4194), .Z(n1149) );
  IV U4197 ( .A(n1152), .Z(mod_mult_o[965]) );
  XOR U4198 ( .A(n4195), .B(n4196), .Z(n1152) );
  IV U4199 ( .A(n1155), .Z(mod_mult_o[964]) );
  XOR U4200 ( .A(n4197), .B(n4198), .Z(n1155) );
  IV U4201 ( .A(n1158), .Z(mod_mult_o[963]) );
  XOR U4202 ( .A(n4199), .B(n4200), .Z(n1158) );
  IV U4203 ( .A(n1161), .Z(mod_mult_o[962]) );
  XOR U4204 ( .A(n4201), .B(n4202), .Z(n1161) );
  IV U4205 ( .A(n1164), .Z(mod_mult_o[961]) );
  XOR U4206 ( .A(n4203), .B(n4204), .Z(n1164) );
  IV U4207 ( .A(n1167), .Z(mod_mult_o[960]) );
  XOR U4208 ( .A(n4205), .B(n4206), .Z(n1167) );
  IV U4209 ( .A(n1170), .Z(mod_mult_o[95]) );
  XOR U4210 ( .A(n4207), .B(n4208), .Z(n1170) );
  IV U4211 ( .A(n1173), .Z(mod_mult_o[959]) );
  XOR U4212 ( .A(n4209), .B(n4210), .Z(n1173) );
  IV U4213 ( .A(n1176), .Z(mod_mult_o[958]) );
  XOR U4214 ( .A(n4211), .B(n4212), .Z(n1176) );
  IV U4215 ( .A(n1179), .Z(mod_mult_o[957]) );
  XOR U4216 ( .A(n4213), .B(n4214), .Z(n1179) );
  IV U4217 ( .A(n1182), .Z(mod_mult_o[956]) );
  XOR U4218 ( .A(n4215), .B(n4216), .Z(n1182) );
  IV U4219 ( .A(n1185), .Z(mod_mult_o[955]) );
  XOR U4220 ( .A(n4217), .B(n4218), .Z(n1185) );
  IV U4221 ( .A(n1188), .Z(mod_mult_o[954]) );
  XOR U4222 ( .A(n4219), .B(n4220), .Z(n1188) );
  IV U4223 ( .A(n1191), .Z(mod_mult_o[953]) );
  XOR U4224 ( .A(n4221), .B(n4222), .Z(n1191) );
  IV U4225 ( .A(n1194), .Z(mod_mult_o[952]) );
  XOR U4226 ( .A(n4223), .B(n4224), .Z(n1194) );
  IV U4227 ( .A(n1197), .Z(mod_mult_o[951]) );
  XOR U4228 ( .A(n4225), .B(n4226), .Z(n1197) );
  IV U4229 ( .A(n1200), .Z(mod_mult_o[950]) );
  XOR U4230 ( .A(n4227), .B(n4228), .Z(n1200) );
  IV U4231 ( .A(n1203), .Z(mod_mult_o[94]) );
  XOR U4232 ( .A(n4229), .B(n4230), .Z(n1203) );
  IV U4233 ( .A(n1206), .Z(mod_mult_o[949]) );
  XOR U4234 ( .A(n4231), .B(n4232), .Z(n1206) );
  IV U4235 ( .A(n1209), .Z(mod_mult_o[948]) );
  XOR U4236 ( .A(n4233), .B(n4234), .Z(n1209) );
  IV U4237 ( .A(n1212), .Z(mod_mult_o[947]) );
  XOR U4238 ( .A(n4235), .B(n4236), .Z(n1212) );
  IV U4239 ( .A(n1215), .Z(mod_mult_o[946]) );
  XOR U4240 ( .A(n4237), .B(n4238), .Z(n1215) );
  IV U4241 ( .A(n1218), .Z(mod_mult_o[945]) );
  XOR U4242 ( .A(n4239), .B(n4240), .Z(n1218) );
  IV U4243 ( .A(n1221), .Z(mod_mult_o[944]) );
  XOR U4244 ( .A(n4241), .B(n4242), .Z(n1221) );
  IV U4245 ( .A(n1224), .Z(mod_mult_o[943]) );
  XOR U4246 ( .A(n4243), .B(n4244), .Z(n1224) );
  IV U4247 ( .A(n1227), .Z(mod_mult_o[942]) );
  XOR U4248 ( .A(n4245), .B(n4246), .Z(n1227) );
  IV U4249 ( .A(n1230), .Z(mod_mult_o[941]) );
  XOR U4250 ( .A(n4247), .B(n4248), .Z(n1230) );
  IV U4251 ( .A(n1233), .Z(mod_mult_o[940]) );
  XOR U4252 ( .A(n4249), .B(n4250), .Z(n1233) );
  IV U4253 ( .A(n1236), .Z(mod_mult_o[93]) );
  XOR U4254 ( .A(n4251), .B(n4252), .Z(n1236) );
  IV U4255 ( .A(n1239), .Z(mod_mult_o[939]) );
  XOR U4256 ( .A(n4253), .B(n4254), .Z(n1239) );
  IV U4257 ( .A(n1242), .Z(mod_mult_o[938]) );
  XOR U4258 ( .A(n4255), .B(n4256), .Z(n1242) );
  IV U4259 ( .A(n1245), .Z(mod_mult_o[937]) );
  XOR U4260 ( .A(n4257), .B(n4258), .Z(n1245) );
  IV U4261 ( .A(n1248), .Z(mod_mult_o[936]) );
  XOR U4262 ( .A(n4259), .B(n4260), .Z(n1248) );
  IV U4263 ( .A(n1251), .Z(mod_mult_o[935]) );
  XOR U4264 ( .A(n4261), .B(n4262), .Z(n1251) );
  IV U4265 ( .A(n1254), .Z(mod_mult_o[934]) );
  XOR U4266 ( .A(n4263), .B(n4264), .Z(n1254) );
  IV U4267 ( .A(n1257), .Z(mod_mult_o[933]) );
  XOR U4268 ( .A(n4265), .B(n4266), .Z(n1257) );
  IV U4269 ( .A(n1260), .Z(mod_mult_o[932]) );
  XOR U4270 ( .A(n4267), .B(n4268), .Z(n1260) );
  IV U4271 ( .A(n1263), .Z(mod_mult_o[931]) );
  XOR U4272 ( .A(n4269), .B(n4270), .Z(n1263) );
  IV U4273 ( .A(n1266), .Z(mod_mult_o[930]) );
  XOR U4274 ( .A(n4271), .B(n4272), .Z(n1266) );
  IV U4275 ( .A(n1269), .Z(mod_mult_o[92]) );
  XOR U4276 ( .A(n4273), .B(n4274), .Z(n1269) );
  IV U4277 ( .A(n1272), .Z(mod_mult_o[929]) );
  XOR U4278 ( .A(n4275), .B(n4276), .Z(n1272) );
  IV U4279 ( .A(n1275), .Z(mod_mult_o[928]) );
  XOR U4280 ( .A(n4277), .B(n4278), .Z(n1275) );
  IV U4281 ( .A(n1278), .Z(mod_mult_o[927]) );
  XOR U4282 ( .A(n4279), .B(n4280), .Z(n1278) );
  IV U4283 ( .A(n1281), .Z(mod_mult_o[926]) );
  XOR U4284 ( .A(n4281), .B(n4282), .Z(n1281) );
  IV U4285 ( .A(n1284), .Z(mod_mult_o[925]) );
  XOR U4286 ( .A(n4283), .B(n4284), .Z(n1284) );
  IV U4287 ( .A(n1287), .Z(mod_mult_o[924]) );
  XOR U4288 ( .A(n4285), .B(n4286), .Z(n1287) );
  IV U4289 ( .A(n1290), .Z(mod_mult_o[923]) );
  XOR U4290 ( .A(n4287), .B(n4288), .Z(n1290) );
  IV U4291 ( .A(n1293), .Z(mod_mult_o[922]) );
  XOR U4292 ( .A(n4289), .B(n4290), .Z(n1293) );
  IV U4293 ( .A(n1296), .Z(mod_mult_o[921]) );
  XOR U4294 ( .A(n4291), .B(n4292), .Z(n1296) );
  IV U4295 ( .A(n1299), .Z(mod_mult_o[920]) );
  XOR U4296 ( .A(n4293), .B(n4294), .Z(n1299) );
  IV U4297 ( .A(n1302), .Z(mod_mult_o[91]) );
  XOR U4298 ( .A(n4295), .B(n4296), .Z(n1302) );
  IV U4299 ( .A(n1305), .Z(mod_mult_o[919]) );
  XOR U4300 ( .A(n4297), .B(n4298), .Z(n1305) );
  IV U4301 ( .A(n1308), .Z(mod_mult_o[918]) );
  XOR U4302 ( .A(n4299), .B(n4300), .Z(n1308) );
  IV U4303 ( .A(n1311), .Z(mod_mult_o[917]) );
  XOR U4304 ( .A(n4301), .B(n4302), .Z(n1311) );
  IV U4305 ( .A(n1314), .Z(mod_mult_o[916]) );
  XOR U4306 ( .A(n4303), .B(n4304), .Z(n1314) );
  IV U4307 ( .A(n1317), .Z(mod_mult_o[915]) );
  XOR U4308 ( .A(n4305), .B(n4306), .Z(n1317) );
  IV U4309 ( .A(n1320), .Z(mod_mult_o[914]) );
  XOR U4310 ( .A(n4307), .B(n4308), .Z(n1320) );
  IV U4311 ( .A(n1323), .Z(mod_mult_o[913]) );
  XOR U4312 ( .A(n4309), .B(n4310), .Z(n1323) );
  IV U4313 ( .A(n1326), .Z(mod_mult_o[912]) );
  XOR U4314 ( .A(n4311), .B(n4312), .Z(n1326) );
  IV U4315 ( .A(n1329), .Z(mod_mult_o[911]) );
  XOR U4316 ( .A(n4313), .B(n4314), .Z(n1329) );
  IV U4317 ( .A(n1332), .Z(mod_mult_o[910]) );
  XOR U4318 ( .A(n4315), .B(n4316), .Z(n1332) );
  IV U4319 ( .A(n1335), .Z(mod_mult_o[90]) );
  XOR U4320 ( .A(n4317), .B(n4318), .Z(n1335) );
  IV U4321 ( .A(n1338), .Z(mod_mult_o[909]) );
  XOR U4322 ( .A(n4319), .B(n4320), .Z(n1338) );
  IV U4323 ( .A(n1341), .Z(mod_mult_o[908]) );
  XOR U4324 ( .A(n4321), .B(n4322), .Z(n1341) );
  IV U4325 ( .A(n1344), .Z(mod_mult_o[907]) );
  XOR U4326 ( .A(n4323), .B(n4324), .Z(n1344) );
  IV U4327 ( .A(n1347), .Z(mod_mult_o[906]) );
  XOR U4328 ( .A(n4325), .B(n4326), .Z(n1347) );
  IV U4329 ( .A(n1350), .Z(mod_mult_o[905]) );
  XOR U4330 ( .A(n4327), .B(n4328), .Z(n1350) );
  IV U4331 ( .A(n1353), .Z(mod_mult_o[904]) );
  XOR U4332 ( .A(n4329), .B(n4330), .Z(n1353) );
  IV U4333 ( .A(n1356), .Z(mod_mult_o[903]) );
  XOR U4334 ( .A(n4331), .B(n4332), .Z(n1356) );
  IV U4335 ( .A(n1359), .Z(mod_mult_o[902]) );
  XOR U4336 ( .A(n4333), .B(n4334), .Z(n1359) );
  IV U4337 ( .A(n1362), .Z(mod_mult_o[901]) );
  XOR U4338 ( .A(n4335), .B(n4336), .Z(n1362) );
  IV U4339 ( .A(n1365), .Z(mod_mult_o[900]) );
  XOR U4340 ( .A(n4337), .B(n4338), .Z(n1365) );
  IV U4341 ( .A(n1368), .Z(mod_mult_o[8]) );
  XOR U4342 ( .A(n4339), .B(n4340), .Z(n1368) );
  IV U4343 ( .A(n1371), .Z(mod_mult_o[89]) );
  XOR U4344 ( .A(n4341), .B(n4342), .Z(n1371) );
  IV U4345 ( .A(n1374), .Z(mod_mult_o[899]) );
  XOR U4346 ( .A(n4343), .B(n4344), .Z(n1374) );
  IV U4347 ( .A(n1377), .Z(mod_mult_o[898]) );
  XOR U4348 ( .A(n4345), .B(n4346), .Z(n1377) );
  IV U4349 ( .A(n1380), .Z(mod_mult_o[897]) );
  XOR U4350 ( .A(n4347), .B(n4348), .Z(n1380) );
  IV U4351 ( .A(n1383), .Z(mod_mult_o[896]) );
  XOR U4352 ( .A(n4349), .B(n4350), .Z(n1383) );
  IV U4353 ( .A(n1386), .Z(mod_mult_o[895]) );
  XOR U4354 ( .A(n4351), .B(n4352), .Z(n1386) );
  IV U4355 ( .A(n1389), .Z(mod_mult_o[894]) );
  XOR U4356 ( .A(n4353), .B(n4354), .Z(n1389) );
  IV U4357 ( .A(n1392), .Z(mod_mult_o[893]) );
  XOR U4358 ( .A(n4355), .B(n4356), .Z(n1392) );
  IV U4359 ( .A(n1395), .Z(mod_mult_o[892]) );
  XOR U4360 ( .A(n4357), .B(n4358), .Z(n1395) );
  IV U4361 ( .A(n1398), .Z(mod_mult_o[891]) );
  XOR U4362 ( .A(n4359), .B(n4360), .Z(n1398) );
  IV U4363 ( .A(n1401), .Z(mod_mult_o[890]) );
  XOR U4364 ( .A(n4361), .B(n4362), .Z(n1401) );
  IV U4365 ( .A(n1404), .Z(mod_mult_o[88]) );
  XOR U4366 ( .A(n4363), .B(n4364), .Z(n1404) );
  IV U4367 ( .A(n1407), .Z(mod_mult_o[889]) );
  XOR U4368 ( .A(n4365), .B(n4366), .Z(n1407) );
  IV U4369 ( .A(n1410), .Z(mod_mult_o[888]) );
  XOR U4370 ( .A(n4367), .B(n4368), .Z(n1410) );
  IV U4371 ( .A(n1413), .Z(mod_mult_o[887]) );
  XOR U4372 ( .A(n4369), .B(n4370), .Z(n1413) );
  IV U4373 ( .A(n1416), .Z(mod_mult_o[886]) );
  XOR U4374 ( .A(n4371), .B(n4372), .Z(n1416) );
  IV U4375 ( .A(n1419), .Z(mod_mult_o[885]) );
  XOR U4376 ( .A(n4373), .B(n4374), .Z(n1419) );
  IV U4377 ( .A(n1422), .Z(mod_mult_o[884]) );
  XOR U4378 ( .A(n4375), .B(n4376), .Z(n1422) );
  IV U4379 ( .A(n1425), .Z(mod_mult_o[883]) );
  XOR U4380 ( .A(n4377), .B(n4378), .Z(n1425) );
  IV U4381 ( .A(n1428), .Z(mod_mult_o[882]) );
  XOR U4382 ( .A(n4379), .B(n4380), .Z(n1428) );
  IV U4383 ( .A(n1431), .Z(mod_mult_o[881]) );
  XOR U4384 ( .A(n4381), .B(n4382), .Z(n1431) );
  IV U4385 ( .A(n1434), .Z(mod_mult_o[880]) );
  XOR U4386 ( .A(n4383), .B(n4384), .Z(n1434) );
  IV U4387 ( .A(n1437), .Z(mod_mult_o[87]) );
  XOR U4388 ( .A(n4385), .B(n4386), .Z(n1437) );
  IV U4389 ( .A(n1440), .Z(mod_mult_o[879]) );
  XOR U4390 ( .A(n4387), .B(n4388), .Z(n1440) );
  IV U4391 ( .A(n1443), .Z(mod_mult_o[878]) );
  XOR U4392 ( .A(n4389), .B(n4390), .Z(n1443) );
  IV U4393 ( .A(n1446), .Z(mod_mult_o[877]) );
  XOR U4394 ( .A(n4391), .B(n4392), .Z(n1446) );
  IV U4395 ( .A(n1449), .Z(mod_mult_o[876]) );
  XOR U4396 ( .A(n4393), .B(n4394), .Z(n1449) );
  IV U4397 ( .A(n1452), .Z(mod_mult_o[875]) );
  XOR U4398 ( .A(n4395), .B(n4396), .Z(n1452) );
  IV U4399 ( .A(n1455), .Z(mod_mult_o[874]) );
  XOR U4400 ( .A(n4397), .B(n4398), .Z(n1455) );
  IV U4401 ( .A(n1458), .Z(mod_mult_o[873]) );
  XOR U4402 ( .A(n4399), .B(n4400), .Z(n1458) );
  IV U4403 ( .A(n1461), .Z(mod_mult_o[872]) );
  XOR U4404 ( .A(n4401), .B(n4402), .Z(n1461) );
  IV U4405 ( .A(n1464), .Z(mod_mult_o[871]) );
  XOR U4406 ( .A(n4403), .B(n4404), .Z(n1464) );
  IV U4407 ( .A(n1467), .Z(mod_mult_o[870]) );
  XOR U4408 ( .A(n4405), .B(n4406), .Z(n1467) );
  IV U4409 ( .A(n1470), .Z(mod_mult_o[86]) );
  XOR U4410 ( .A(n4407), .B(n4408), .Z(n1470) );
  IV U4411 ( .A(n1473), .Z(mod_mult_o[869]) );
  XOR U4412 ( .A(n4409), .B(n4410), .Z(n1473) );
  IV U4413 ( .A(n1476), .Z(mod_mult_o[868]) );
  XOR U4414 ( .A(n4411), .B(n4412), .Z(n1476) );
  IV U4415 ( .A(n1479), .Z(mod_mult_o[867]) );
  XOR U4416 ( .A(n4413), .B(n4414), .Z(n1479) );
  IV U4417 ( .A(n1482), .Z(mod_mult_o[866]) );
  XOR U4418 ( .A(n4415), .B(n4416), .Z(n1482) );
  IV U4419 ( .A(n1485), .Z(mod_mult_o[865]) );
  XOR U4420 ( .A(n4417), .B(n4418), .Z(n1485) );
  IV U4421 ( .A(n1488), .Z(mod_mult_o[864]) );
  XOR U4422 ( .A(n4419), .B(n4420), .Z(n1488) );
  IV U4423 ( .A(n1491), .Z(mod_mult_o[863]) );
  XOR U4424 ( .A(n4421), .B(n4422), .Z(n1491) );
  IV U4425 ( .A(n1494), .Z(mod_mult_o[862]) );
  XOR U4426 ( .A(n4423), .B(n4424), .Z(n1494) );
  IV U4427 ( .A(n1497), .Z(mod_mult_o[861]) );
  XOR U4428 ( .A(n4425), .B(n4426), .Z(n1497) );
  IV U4429 ( .A(n1500), .Z(mod_mult_o[860]) );
  XOR U4430 ( .A(n4427), .B(n4428), .Z(n1500) );
  IV U4431 ( .A(n1503), .Z(mod_mult_o[85]) );
  XOR U4432 ( .A(n4429), .B(n4430), .Z(n1503) );
  IV U4433 ( .A(n1506), .Z(mod_mult_o[859]) );
  XOR U4434 ( .A(n4431), .B(n4432), .Z(n1506) );
  IV U4435 ( .A(n1509), .Z(mod_mult_o[858]) );
  XOR U4436 ( .A(n4433), .B(n4434), .Z(n1509) );
  IV U4437 ( .A(n1512), .Z(mod_mult_o[857]) );
  XOR U4438 ( .A(n4435), .B(n4436), .Z(n1512) );
  IV U4439 ( .A(n1515), .Z(mod_mult_o[856]) );
  XOR U4440 ( .A(n4437), .B(n4438), .Z(n1515) );
  IV U4441 ( .A(n1518), .Z(mod_mult_o[855]) );
  XOR U4442 ( .A(n4439), .B(n4440), .Z(n1518) );
  IV U4443 ( .A(n1521), .Z(mod_mult_o[854]) );
  XOR U4444 ( .A(n4441), .B(n4442), .Z(n1521) );
  IV U4445 ( .A(n1524), .Z(mod_mult_o[853]) );
  XOR U4446 ( .A(n4443), .B(n4444), .Z(n1524) );
  IV U4447 ( .A(n1527), .Z(mod_mult_o[852]) );
  XOR U4448 ( .A(n4445), .B(n4446), .Z(n1527) );
  IV U4449 ( .A(n1530), .Z(mod_mult_o[851]) );
  XOR U4450 ( .A(n4447), .B(n4448), .Z(n1530) );
  IV U4451 ( .A(n1533), .Z(mod_mult_o[850]) );
  XOR U4452 ( .A(n4449), .B(n4450), .Z(n1533) );
  IV U4453 ( .A(n1536), .Z(mod_mult_o[84]) );
  XOR U4454 ( .A(n4451), .B(n4452), .Z(n1536) );
  IV U4455 ( .A(n1539), .Z(mod_mult_o[849]) );
  XOR U4456 ( .A(n4453), .B(n4454), .Z(n1539) );
  IV U4457 ( .A(n1542), .Z(mod_mult_o[848]) );
  XOR U4458 ( .A(n4455), .B(n4456), .Z(n1542) );
  IV U4459 ( .A(n1545), .Z(mod_mult_o[847]) );
  XOR U4460 ( .A(n4457), .B(n4458), .Z(n1545) );
  IV U4461 ( .A(n1548), .Z(mod_mult_o[846]) );
  XOR U4462 ( .A(n4459), .B(n4460), .Z(n1548) );
  IV U4463 ( .A(n1551), .Z(mod_mult_o[845]) );
  XOR U4464 ( .A(n4461), .B(n4462), .Z(n1551) );
  IV U4465 ( .A(n1554), .Z(mod_mult_o[844]) );
  XOR U4466 ( .A(n4463), .B(n4464), .Z(n1554) );
  IV U4467 ( .A(n1557), .Z(mod_mult_o[843]) );
  XOR U4468 ( .A(n4465), .B(n4466), .Z(n1557) );
  IV U4469 ( .A(n1560), .Z(mod_mult_o[842]) );
  XOR U4470 ( .A(n4467), .B(n4468), .Z(n1560) );
  IV U4471 ( .A(n1563), .Z(mod_mult_o[841]) );
  XOR U4472 ( .A(n4469), .B(n4470), .Z(n1563) );
  IV U4473 ( .A(n1566), .Z(mod_mult_o[840]) );
  XOR U4474 ( .A(n4471), .B(n4472), .Z(n1566) );
  IV U4475 ( .A(n1569), .Z(mod_mult_o[83]) );
  XOR U4476 ( .A(n4473), .B(n4474), .Z(n1569) );
  IV U4477 ( .A(n1572), .Z(mod_mult_o[839]) );
  XOR U4478 ( .A(n4475), .B(n4476), .Z(n1572) );
  IV U4479 ( .A(n1575), .Z(mod_mult_o[838]) );
  XOR U4480 ( .A(n4477), .B(n4478), .Z(n1575) );
  IV U4481 ( .A(n1578), .Z(mod_mult_o[837]) );
  XOR U4482 ( .A(n4479), .B(n4480), .Z(n1578) );
  IV U4483 ( .A(n1581), .Z(mod_mult_o[836]) );
  XOR U4484 ( .A(n4481), .B(n4482), .Z(n1581) );
  IV U4485 ( .A(n1584), .Z(mod_mult_o[835]) );
  XOR U4486 ( .A(n4483), .B(n4484), .Z(n1584) );
  IV U4487 ( .A(n1587), .Z(mod_mult_o[834]) );
  XOR U4488 ( .A(n4485), .B(n4486), .Z(n1587) );
  IV U4489 ( .A(n1590), .Z(mod_mult_o[833]) );
  XOR U4490 ( .A(n4487), .B(n4488), .Z(n1590) );
  IV U4491 ( .A(n1593), .Z(mod_mult_o[832]) );
  XOR U4492 ( .A(n4489), .B(n4490), .Z(n1593) );
  IV U4493 ( .A(n1596), .Z(mod_mult_o[831]) );
  XOR U4494 ( .A(n4491), .B(n4492), .Z(n1596) );
  IV U4495 ( .A(n1599), .Z(mod_mult_o[830]) );
  XOR U4496 ( .A(n4493), .B(n4494), .Z(n1599) );
  IV U4497 ( .A(n1602), .Z(mod_mult_o[82]) );
  XOR U4498 ( .A(n4495), .B(n4496), .Z(n1602) );
  IV U4499 ( .A(n1605), .Z(mod_mult_o[829]) );
  XOR U4500 ( .A(n4497), .B(n4498), .Z(n1605) );
  IV U4501 ( .A(n1608), .Z(mod_mult_o[828]) );
  XOR U4502 ( .A(n4499), .B(n4500), .Z(n1608) );
  IV U4503 ( .A(n1611), .Z(mod_mult_o[827]) );
  XOR U4504 ( .A(n4501), .B(n4502), .Z(n1611) );
  IV U4505 ( .A(n1614), .Z(mod_mult_o[826]) );
  XOR U4506 ( .A(n4503), .B(n4504), .Z(n1614) );
  IV U4507 ( .A(n1617), .Z(mod_mult_o[825]) );
  XOR U4508 ( .A(n4505), .B(n4506), .Z(n1617) );
  IV U4509 ( .A(n1620), .Z(mod_mult_o[824]) );
  XOR U4510 ( .A(n4507), .B(n4508), .Z(n1620) );
  IV U4511 ( .A(n1623), .Z(mod_mult_o[823]) );
  XOR U4512 ( .A(n4509), .B(n4510), .Z(n1623) );
  IV U4513 ( .A(n1626), .Z(mod_mult_o[822]) );
  XOR U4514 ( .A(n4511), .B(n4512), .Z(n1626) );
  IV U4515 ( .A(n1629), .Z(mod_mult_o[821]) );
  XOR U4516 ( .A(n4513), .B(n4514), .Z(n1629) );
  IV U4517 ( .A(n1632), .Z(mod_mult_o[820]) );
  XOR U4518 ( .A(n4515), .B(n4516), .Z(n1632) );
  IV U4519 ( .A(n1635), .Z(mod_mult_o[81]) );
  XOR U4520 ( .A(n4517), .B(n4518), .Z(n1635) );
  IV U4521 ( .A(n1638), .Z(mod_mult_o[819]) );
  XOR U4522 ( .A(n4519), .B(n4520), .Z(n1638) );
  IV U4523 ( .A(n1641), .Z(mod_mult_o[818]) );
  XOR U4524 ( .A(n4521), .B(n4522), .Z(n1641) );
  IV U4525 ( .A(n1644), .Z(mod_mult_o[817]) );
  XOR U4526 ( .A(n4523), .B(n4524), .Z(n1644) );
  IV U4527 ( .A(n1647), .Z(mod_mult_o[816]) );
  XOR U4528 ( .A(n4525), .B(n4526), .Z(n1647) );
  IV U4529 ( .A(n1650), .Z(mod_mult_o[815]) );
  XOR U4530 ( .A(n4527), .B(n4528), .Z(n1650) );
  IV U4531 ( .A(n1653), .Z(mod_mult_o[814]) );
  XOR U4532 ( .A(n4529), .B(n4530), .Z(n1653) );
  IV U4533 ( .A(n1656), .Z(mod_mult_o[813]) );
  XOR U4534 ( .A(n4531), .B(n4532), .Z(n1656) );
  IV U4535 ( .A(n1659), .Z(mod_mult_o[812]) );
  XOR U4536 ( .A(n4533), .B(n4534), .Z(n1659) );
  IV U4537 ( .A(n1662), .Z(mod_mult_o[811]) );
  XOR U4538 ( .A(n4535), .B(n4536), .Z(n1662) );
  IV U4539 ( .A(n1665), .Z(mod_mult_o[810]) );
  XOR U4540 ( .A(n4537), .B(n4538), .Z(n1665) );
  IV U4541 ( .A(n1668), .Z(mod_mult_o[80]) );
  XOR U4542 ( .A(n4539), .B(n4540), .Z(n1668) );
  IV U4543 ( .A(n1671), .Z(mod_mult_o[809]) );
  XOR U4544 ( .A(n4541), .B(n4542), .Z(n1671) );
  IV U4545 ( .A(n1674), .Z(mod_mult_o[808]) );
  XOR U4546 ( .A(n4543), .B(n4544), .Z(n1674) );
  IV U4547 ( .A(n1677), .Z(mod_mult_o[807]) );
  XOR U4548 ( .A(n4545), .B(n4546), .Z(n1677) );
  IV U4549 ( .A(n1680), .Z(mod_mult_o[806]) );
  XOR U4550 ( .A(n4547), .B(n4548), .Z(n1680) );
  IV U4551 ( .A(n1683), .Z(mod_mult_o[805]) );
  XOR U4552 ( .A(n4549), .B(n4550), .Z(n1683) );
  IV U4553 ( .A(n1686), .Z(mod_mult_o[804]) );
  XOR U4554 ( .A(n4551), .B(n4552), .Z(n1686) );
  IV U4555 ( .A(n1689), .Z(mod_mult_o[803]) );
  XOR U4556 ( .A(n4553), .B(n4554), .Z(n1689) );
  IV U4557 ( .A(n1692), .Z(mod_mult_o[802]) );
  XOR U4558 ( .A(n4555), .B(n4556), .Z(n1692) );
  IV U4559 ( .A(n1695), .Z(mod_mult_o[801]) );
  XOR U4560 ( .A(n4557), .B(n4558), .Z(n1695) );
  IV U4561 ( .A(n1698), .Z(mod_mult_o[800]) );
  XOR U4562 ( .A(n4559), .B(n4560), .Z(n1698) );
  IV U4563 ( .A(n1701), .Z(mod_mult_o[7]) );
  XOR U4564 ( .A(n4561), .B(n4562), .Z(n1701) );
  IV U4565 ( .A(n1704), .Z(mod_mult_o[79]) );
  XOR U4566 ( .A(n4563), .B(n4564), .Z(n1704) );
  IV U4567 ( .A(n1707), .Z(mod_mult_o[799]) );
  XOR U4568 ( .A(n4565), .B(n4566), .Z(n1707) );
  IV U4569 ( .A(n1710), .Z(mod_mult_o[798]) );
  XOR U4570 ( .A(n4567), .B(n4568), .Z(n1710) );
  IV U4571 ( .A(n1713), .Z(mod_mult_o[797]) );
  XOR U4572 ( .A(n4569), .B(n4570), .Z(n1713) );
  IV U4573 ( .A(n1716), .Z(mod_mult_o[796]) );
  XOR U4574 ( .A(n4571), .B(n4572), .Z(n1716) );
  IV U4575 ( .A(n1719), .Z(mod_mult_o[795]) );
  XOR U4576 ( .A(n4573), .B(n4574), .Z(n1719) );
  IV U4577 ( .A(n1722), .Z(mod_mult_o[794]) );
  XOR U4578 ( .A(n4575), .B(n4576), .Z(n1722) );
  IV U4579 ( .A(n1725), .Z(mod_mult_o[793]) );
  XOR U4580 ( .A(n4577), .B(n4578), .Z(n1725) );
  IV U4581 ( .A(n1728), .Z(mod_mult_o[792]) );
  XOR U4582 ( .A(n4579), .B(n4580), .Z(n1728) );
  IV U4583 ( .A(n1731), .Z(mod_mult_o[791]) );
  XOR U4584 ( .A(n4581), .B(n4582), .Z(n1731) );
  IV U4585 ( .A(n1734), .Z(mod_mult_o[790]) );
  XOR U4586 ( .A(n4583), .B(n4584), .Z(n1734) );
  IV U4587 ( .A(n1737), .Z(mod_mult_o[78]) );
  XOR U4588 ( .A(n4585), .B(n4586), .Z(n1737) );
  IV U4589 ( .A(n1740), .Z(mod_mult_o[789]) );
  XOR U4590 ( .A(n4587), .B(n4588), .Z(n1740) );
  IV U4591 ( .A(n1743), .Z(mod_mult_o[788]) );
  XOR U4592 ( .A(n4589), .B(n4590), .Z(n1743) );
  IV U4593 ( .A(n1746), .Z(mod_mult_o[787]) );
  XOR U4594 ( .A(n4591), .B(n4592), .Z(n1746) );
  IV U4595 ( .A(n1749), .Z(mod_mult_o[786]) );
  XOR U4596 ( .A(n4593), .B(n4594), .Z(n1749) );
  IV U4597 ( .A(n1752), .Z(mod_mult_o[785]) );
  XOR U4598 ( .A(n4595), .B(n4596), .Z(n1752) );
  IV U4599 ( .A(n1755), .Z(mod_mult_o[784]) );
  XOR U4600 ( .A(n4597), .B(n4598), .Z(n1755) );
  IV U4601 ( .A(n1758), .Z(mod_mult_o[783]) );
  XOR U4602 ( .A(n4599), .B(n4600), .Z(n1758) );
  IV U4603 ( .A(n1761), .Z(mod_mult_o[782]) );
  XOR U4604 ( .A(n4601), .B(n4602), .Z(n1761) );
  IV U4605 ( .A(n1764), .Z(mod_mult_o[781]) );
  XOR U4606 ( .A(n4603), .B(n4604), .Z(n1764) );
  IV U4607 ( .A(n1767), .Z(mod_mult_o[780]) );
  XOR U4608 ( .A(n4605), .B(n4606), .Z(n1767) );
  IV U4609 ( .A(n1770), .Z(mod_mult_o[77]) );
  XOR U4610 ( .A(n4607), .B(n4608), .Z(n1770) );
  IV U4611 ( .A(n1773), .Z(mod_mult_o[779]) );
  XOR U4612 ( .A(n4609), .B(n4610), .Z(n1773) );
  IV U4613 ( .A(n1776), .Z(mod_mult_o[778]) );
  XOR U4614 ( .A(n4611), .B(n4612), .Z(n1776) );
  IV U4615 ( .A(n1779), .Z(mod_mult_o[777]) );
  XOR U4616 ( .A(n4613), .B(n4614), .Z(n1779) );
  IV U4617 ( .A(n1782), .Z(mod_mult_o[776]) );
  XOR U4618 ( .A(n4615), .B(n4616), .Z(n1782) );
  IV U4619 ( .A(n1785), .Z(mod_mult_o[775]) );
  XOR U4620 ( .A(n4617), .B(n4618), .Z(n1785) );
  IV U4621 ( .A(n1788), .Z(mod_mult_o[774]) );
  XOR U4622 ( .A(n4619), .B(n4620), .Z(n1788) );
  IV U4623 ( .A(n1791), .Z(mod_mult_o[773]) );
  XOR U4624 ( .A(n4621), .B(n4622), .Z(n1791) );
  IV U4625 ( .A(n1794), .Z(mod_mult_o[772]) );
  XOR U4626 ( .A(n4623), .B(n4624), .Z(n1794) );
  IV U4627 ( .A(n1797), .Z(mod_mult_o[771]) );
  XOR U4628 ( .A(n4625), .B(n4626), .Z(n1797) );
  IV U4629 ( .A(n1800), .Z(mod_mult_o[770]) );
  XOR U4630 ( .A(n4627), .B(n4628), .Z(n1800) );
  IV U4631 ( .A(n1803), .Z(mod_mult_o[76]) );
  XOR U4632 ( .A(n4629), .B(n4630), .Z(n1803) );
  IV U4633 ( .A(n1806), .Z(mod_mult_o[769]) );
  XOR U4634 ( .A(n4631), .B(n4632), .Z(n1806) );
  IV U4635 ( .A(n1809), .Z(mod_mult_o[768]) );
  XOR U4636 ( .A(n4633), .B(n4634), .Z(n1809) );
  IV U4637 ( .A(n1812), .Z(mod_mult_o[767]) );
  XOR U4638 ( .A(n4635), .B(n4636), .Z(n1812) );
  IV U4639 ( .A(n1815), .Z(mod_mult_o[766]) );
  XOR U4640 ( .A(n4637), .B(n4638), .Z(n1815) );
  IV U4641 ( .A(n1818), .Z(mod_mult_o[765]) );
  XOR U4642 ( .A(n4639), .B(n4640), .Z(n1818) );
  IV U4643 ( .A(n1821), .Z(mod_mult_o[764]) );
  XOR U4644 ( .A(n4641), .B(n4642), .Z(n1821) );
  IV U4645 ( .A(n1824), .Z(mod_mult_o[763]) );
  XOR U4646 ( .A(n4643), .B(n4644), .Z(n1824) );
  IV U4647 ( .A(n1827), .Z(mod_mult_o[762]) );
  XOR U4648 ( .A(n4645), .B(n4646), .Z(n1827) );
  IV U4649 ( .A(n1830), .Z(mod_mult_o[761]) );
  XOR U4650 ( .A(n4647), .B(n4648), .Z(n1830) );
  IV U4651 ( .A(n1833), .Z(mod_mult_o[760]) );
  XOR U4652 ( .A(n4649), .B(n4650), .Z(n1833) );
  IV U4653 ( .A(n1836), .Z(mod_mult_o[75]) );
  XOR U4654 ( .A(n4651), .B(n4652), .Z(n1836) );
  IV U4655 ( .A(n1839), .Z(mod_mult_o[759]) );
  XOR U4656 ( .A(n4653), .B(n4654), .Z(n1839) );
  IV U4657 ( .A(n1842), .Z(mod_mult_o[758]) );
  XOR U4658 ( .A(n4655), .B(n4656), .Z(n1842) );
  IV U4659 ( .A(n1845), .Z(mod_mult_o[757]) );
  XOR U4660 ( .A(n4657), .B(n4658), .Z(n1845) );
  IV U4661 ( .A(n1848), .Z(mod_mult_o[756]) );
  XOR U4662 ( .A(n4659), .B(n4660), .Z(n1848) );
  IV U4663 ( .A(n1851), .Z(mod_mult_o[755]) );
  XOR U4664 ( .A(n4661), .B(n4662), .Z(n1851) );
  IV U4665 ( .A(n1854), .Z(mod_mult_o[754]) );
  XOR U4666 ( .A(n4663), .B(n4664), .Z(n1854) );
  IV U4667 ( .A(n1857), .Z(mod_mult_o[753]) );
  XOR U4668 ( .A(n4665), .B(n4666), .Z(n1857) );
  IV U4669 ( .A(n1860), .Z(mod_mult_o[752]) );
  XOR U4670 ( .A(n4667), .B(n4668), .Z(n1860) );
  IV U4671 ( .A(n1863), .Z(mod_mult_o[751]) );
  XOR U4672 ( .A(n4669), .B(n4670), .Z(n1863) );
  IV U4673 ( .A(n1866), .Z(mod_mult_o[750]) );
  XOR U4674 ( .A(n4671), .B(n4672), .Z(n1866) );
  IV U4675 ( .A(n1869), .Z(mod_mult_o[74]) );
  XOR U4676 ( .A(n4673), .B(n4674), .Z(n1869) );
  IV U4677 ( .A(n1872), .Z(mod_mult_o[749]) );
  XOR U4678 ( .A(n4675), .B(n4676), .Z(n1872) );
  IV U4679 ( .A(n1875), .Z(mod_mult_o[748]) );
  XOR U4680 ( .A(n4677), .B(n4678), .Z(n1875) );
  IV U4681 ( .A(n1878), .Z(mod_mult_o[747]) );
  XOR U4682 ( .A(n4679), .B(n4680), .Z(n1878) );
  IV U4683 ( .A(n1881), .Z(mod_mult_o[746]) );
  XOR U4684 ( .A(n4681), .B(n4682), .Z(n1881) );
  IV U4685 ( .A(n1884), .Z(mod_mult_o[745]) );
  XOR U4686 ( .A(n4683), .B(n4684), .Z(n1884) );
  IV U4687 ( .A(n1887), .Z(mod_mult_o[744]) );
  XOR U4688 ( .A(n4685), .B(n4686), .Z(n1887) );
  IV U4689 ( .A(n1890), .Z(mod_mult_o[743]) );
  XOR U4690 ( .A(n4687), .B(n4688), .Z(n1890) );
  IV U4691 ( .A(n1893), .Z(mod_mult_o[742]) );
  XOR U4692 ( .A(n4689), .B(n4690), .Z(n1893) );
  IV U4693 ( .A(n1896), .Z(mod_mult_o[741]) );
  XOR U4694 ( .A(n4691), .B(n4692), .Z(n1896) );
  IV U4695 ( .A(n1899), .Z(mod_mult_o[740]) );
  XOR U4696 ( .A(n4693), .B(n4694), .Z(n1899) );
  IV U4697 ( .A(n1902), .Z(mod_mult_o[73]) );
  XOR U4698 ( .A(n4695), .B(n4696), .Z(n1902) );
  IV U4699 ( .A(n1905), .Z(mod_mult_o[739]) );
  XOR U4700 ( .A(n4697), .B(n4698), .Z(n1905) );
  IV U4701 ( .A(n1908), .Z(mod_mult_o[738]) );
  XOR U4702 ( .A(n4699), .B(n4700), .Z(n1908) );
  IV U4703 ( .A(n1911), .Z(mod_mult_o[737]) );
  XOR U4704 ( .A(n4701), .B(n4702), .Z(n1911) );
  IV U4705 ( .A(n1914), .Z(mod_mult_o[736]) );
  XOR U4706 ( .A(n4703), .B(n4704), .Z(n1914) );
  IV U4707 ( .A(n1917), .Z(mod_mult_o[735]) );
  XOR U4708 ( .A(n4705), .B(n4706), .Z(n1917) );
  IV U4709 ( .A(n1920), .Z(mod_mult_o[734]) );
  XOR U4710 ( .A(n4707), .B(n4708), .Z(n1920) );
  IV U4711 ( .A(n1923), .Z(mod_mult_o[733]) );
  XOR U4712 ( .A(n4709), .B(n4710), .Z(n1923) );
  IV U4713 ( .A(n1926), .Z(mod_mult_o[732]) );
  XOR U4714 ( .A(n4711), .B(n4712), .Z(n1926) );
  IV U4715 ( .A(n1929), .Z(mod_mult_o[731]) );
  XOR U4716 ( .A(n4713), .B(n4714), .Z(n1929) );
  IV U4717 ( .A(n1932), .Z(mod_mult_o[730]) );
  XOR U4718 ( .A(n4715), .B(n4716), .Z(n1932) );
  IV U4719 ( .A(n1935), .Z(mod_mult_o[72]) );
  XOR U4720 ( .A(n4717), .B(n4718), .Z(n1935) );
  IV U4721 ( .A(n1938), .Z(mod_mult_o[729]) );
  XOR U4722 ( .A(n4719), .B(n4720), .Z(n1938) );
  IV U4723 ( .A(n1941), .Z(mod_mult_o[728]) );
  XOR U4724 ( .A(n4721), .B(n4722), .Z(n1941) );
  IV U4725 ( .A(n1944), .Z(mod_mult_o[727]) );
  XOR U4726 ( .A(n4723), .B(n4724), .Z(n1944) );
  IV U4727 ( .A(n1947), .Z(mod_mult_o[726]) );
  XOR U4728 ( .A(n4725), .B(n4726), .Z(n1947) );
  IV U4729 ( .A(n1950), .Z(mod_mult_o[725]) );
  XOR U4730 ( .A(n4727), .B(n4728), .Z(n1950) );
  IV U4731 ( .A(n1953), .Z(mod_mult_o[724]) );
  XOR U4732 ( .A(n4729), .B(n4730), .Z(n1953) );
  IV U4733 ( .A(n1956), .Z(mod_mult_o[723]) );
  XOR U4734 ( .A(n4731), .B(n4732), .Z(n1956) );
  IV U4735 ( .A(n1959), .Z(mod_mult_o[722]) );
  XOR U4736 ( .A(n4733), .B(n4734), .Z(n1959) );
  IV U4737 ( .A(n1962), .Z(mod_mult_o[721]) );
  XOR U4738 ( .A(n4735), .B(n4736), .Z(n1962) );
  IV U4739 ( .A(n1965), .Z(mod_mult_o[720]) );
  XOR U4740 ( .A(n4737), .B(n4738), .Z(n1965) );
  IV U4741 ( .A(n1968), .Z(mod_mult_o[71]) );
  XOR U4742 ( .A(n4739), .B(n4740), .Z(n1968) );
  IV U4743 ( .A(n1971), .Z(mod_mult_o[719]) );
  XOR U4744 ( .A(n4741), .B(n4742), .Z(n1971) );
  IV U4745 ( .A(n1974), .Z(mod_mult_o[718]) );
  XOR U4746 ( .A(n4743), .B(n4744), .Z(n1974) );
  IV U4747 ( .A(n1977), .Z(mod_mult_o[717]) );
  XOR U4748 ( .A(n4745), .B(n4746), .Z(n1977) );
  IV U4749 ( .A(n1980), .Z(mod_mult_o[716]) );
  XOR U4750 ( .A(n4747), .B(n4748), .Z(n1980) );
  IV U4751 ( .A(n1983), .Z(mod_mult_o[715]) );
  XOR U4752 ( .A(n4749), .B(n4750), .Z(n1983) );
  IV U4753 ( .A(n1986), .Z(mod_mult_o[714]) );
  XOR U4754 ( .A(n4751), .B(n4752), .Z(n1986) );
  IV U4755 ( .A(n1989), .Z(mod_mult_o[713]) );
  XOR U4756 ( .A(n4753), .B(n4754), .Z(n1989) );
  IV U4757 ( .A(n1992), .Z(mod_mult_o[712]) );
  XOR U4758 ( .A(n4755), .B(n4756), .Z(n1992) );
  IV U4759 ( .A(n1995), .Z(mod_mult_o[711]) );
  XOR U4760 ( .A(n4757), .B(n4758), .Z(n1995) );
  IV U4761 ( .A(n1998), .Z(mod_mult_o[710]) );
  XOR U4762 ( .A(n4759), .B(n4760), .Z(n1998) );
  IV U4763 ( .A(n2001), .Z(mod_mult_o[70]) );
  XOR U4764 ( .A(n4761), .B(n4762), .Z(n2001) );
  IV U4765 ( .A(n2004), .Z(mod_mult_o[709]) );
  XOR U4766 ( .A(n4763), .B(n4764), .Z(n2004) );
  IV U4767 ( .A(n2007), .Z(mod_mult_o[708]) );
  XOR U4768 ( .A(n4765), .B(n4766), .Z(n2007) );
  IV U4769 ( .A(n2010), .Z(mod_mult_o[707]) );
  XOR U4770 ( .A(n4767), .B(n4768), .Z(n2010) );
  IV U4771 ( .A(n2013), .Z(mod_mult_o[706]) );
  XOR U4772 ( .A(n4769), .B(n4770), .Z(n2013) );
  IV U4773 ( .A(n2016), .Z(mod_mult_o[705]) );
  XOR U4774 ( .A(n4771), .B(n4772), .Z(n2016) );
  IV U4775 ( .A(n2019), .Z(mod_mult_o[704]) );
  XOR U4776 ( .A(n4773), .B(n4774), .Z(n2019) );
  IV U4777 ( .A(n2022), .Z(mod_mult_o[703]) );
  XOR U4778 ( .A(n4775), .B(n4776), .Z(n2022) );
  IV U4779 ( .A(n2025), .Z(mod_mult_o[702]) );
  XOR U4780 ( .A(n4777), .B(n4778), .Z(n2025) );
  IV U4781 ( .A(n2028), .Z(mod_mult_o[701]) );
  XOR U4782 ( .A(n4779), .B(n4780), .Z(n2028) );
  IV U4783 ( .A(n2031), .Z(mod_mult_o[700]) );
  XOR U4784 ( .A(n4781), .B(n4782), .Z(n2031) );
  IV U4785 ( .A(n2034), .Z(mod_mult_o[6]) );
  XOR U4786 ( .A(n4783), .B(n4784), .Z(n2034) );
  IV U4787 ( .A(n2037), .Z(mod_mult_o[69]) );
  XOR U4788 ( .A(n4785), .B(n4786), .Z(n2037) );
  IV U4789 ( .A(n2040), .Z(mod_mult_o[699]) );
  XOR U4790 ( .A(n4787), .B(n4788), .Z(n2040) );
  IV U4791 ( .A(n2043), .Z(mod_mult_o[698]) );
  XOR U4792 ( .A(n4789), .B(n4790), .Z(n2043) );
  IV U4793 ( .A(n2046), .Z(mod_mult_o[697]) );
  XOR U4794 ( .A(n4791), .B(n4792), .Z(n2046) );
  IV U4795 ( .A(n2049), .Z(mod_mult_o[696]) );
  XOR U4796 ( .A(n4793), .B(n4794), .Z(n2049) );
  IV U4797 ( .A(n2052), .Z(mod_mult_o[695]) );
  XOR U4798 ( .A(n4795), .B(n4796), .Z(n2052) );
  IV U4799 ( .A(n2055), .Z(mod_mult_o[694]) );
  XOR U4800 ( .A(n4797), .B(n4798), .Z(n2055) );
  IV U4801 ( .A(n2058), .Z(mod_mult_o[693]) );
  XOR U4802 ( .A(n4799), .B(n4800), .Z(n2058) );
  IV U4803 ( .A(n2061), .Z(mod_mult_o[692]) );
  XOR U4804 ( .A(n4801), .B(n4802), .Z(n2061) );
  IV U4805 ( .A(n2064), .Z(mod_mult_o[691]) );
  XOR U4806 ( .A(n4803), .B(n4804), .Z(n2064) );
  IV U4807 ( .A(n2067), .Z(mod_mult_o[690]) );
  XOR U4808 ( .A(n4805), .B(n4806), .Z(n2067) );
  IV U4809 ( .A(n2070), .Z(mod_mult_o[68]) );
  XOR U4810 ( .A(n4807), .B(n4808), .Z(n2070) );
  IV U4811 ( .A(n2073), .Z(mod_mult_o[689]) );
  XOR U4812 ( .A(n4809), .B(n4810), .Z(n2073) );
  IV U4813 ( .A(n2076), .Z(mod_mult_o[688]) );
  XOR U4814 ( .A(n4811), .B(n4812), .Z(n2076) );
  IV U4815 ( .A(n2079), .Z(mod_mult_o[687]) );
  XOR U4816 ( .A(n4813), .B(n4814), .Z(n2079) );
  IV U4817 ( .A(n2082), .Z(mod_mult_o[686]) );
  XOR U4818 ( .A(n4815), .B(n4816), .Z(n2082) );
  IV U4819 ( .A(n2085), .Z(mod_mult_o[685]) );
  XOR U4820 ( .A(n4817), .B(n4818), .Z(n2085) );
  IV U4821 ( .A(n2088), .Z(mod_mult_o[684]) );
  XOR U4822 ( .A(n4819), .B(n4820), .Z(n2088) );
  IV U4823 ( .A(n2091), .Z(mod_mult_o[683]) );
  XOR U4824 ( .A(n4821), .B(n4822), .Z(n2091) );
  IV U4825 ( .A(n2094), .Z(mod_mult_o[682]) );
  XOR U4826 ( .A(n4823), .B(n4824), .Z(n2094) );
  IV U4827 ( .A(n2097), .Z(mod_mult_o[681]) );
  XOR U4828 ( .A(n4825), .B(n4826), .Z(n2097) );
  IV U4829 ( .A(n2100), .Z(mod_mult_o[680]) );
  XOR U4830 ( .A(n4827), .B(n4828), .Z(n2100) );
  IV U4831 ( .A(n2103), .Z(mod_mult_o[67]) );
  XOR U4832 ( .A(n4829), .B(n4830), .Z(n2103) );
  IV U4833 ( .A(n2106), .Z(mod_mult_o[679]) );
  XOR U4834 ( .A(n4831), .B(n4832), .Z(n2106) );
  IV U4835 ( .A(n2109), .Z(mod_mult_o[678]) );
  XOR U4836 ( .A(n4833), .B(n4834), .Z(n2109) );
  IV U4837 ( .A(n2112), .Z(mod_mult_o[677]) );
  XOR U4838 ( .A(n4835), .B(n4836), .Z(n2112) );
  IV U4839 ( .A(n2115), .Z(mod_mult_o[676]) );
  XOR U4840 ( .A(n4837), .B(n4838), .Z(n2115) );
  IV U4841 ( .A(n2118), .Z(mod_mult_o[675]) );
  XOR U4842 ( .A(n4839), .B(n4840), .Z(n2118) );
  IV U4843 ( .A(n2121), .Z(mod_mult_o[674]) );
  XOR U4844 ( .A(n4841), .B(n4842), .Z(n2121) );
  IV U4845 ( .A(n2124), .Z(mod_mult_o[673]) );
  XOR U4846 ( .A(n4843), .B(n4844), .Z(n2124) );
  IV U4847 ( .A(n2127), .Z(mod_mult_o[672]) );
  XOR U4848 ( .A(n4845), .B(n4846), .Z(n2127) );
  IV U4849 ( .A(n2130), .Z(mod_mult_o[671]) );
  XOR U4850 ( .A(n4847), .B(n4848), .Z(n2130) );
  IV U4851 ( .A(n2133), .Z(mod_mult_o[670]) );
  XOR U4852 ( .A(n4849), .B(n4850), .Z(n2133) );
  IV U4853 ( .A(n2136), .Z(mod_mult_o[66]) );
  XOR U4854 ( .A(n4851), .B(n4852), .Z(n2136) );
  IV U4855 ( .A(n2139), .Z(mod_mult_o[669]) );
  XOR U4856 ( .A(n4853), .B(n4854), .Z(n2139) );
  IV U4857 ( .A(n2142), .Z(mod_mult_o[668]) );
  XOR U4858 ( .A(n4855), .B(n4856), .Z(n2142) );
  IV U4859 ( .A(n2145), .Z(mod_mult_o[667]) );
  XOR U4860 ( .A(n4857), .B(n4858), .Z(n2145) );
  IV U4861 ( .A(n2148), .Z(mod_mult_o[666]) );
  XOR U4862 ( .A(n4859), .B(n4860), .Z(n2148) );
  IV U4863 ( .A(n2151), .Z(mod_mult_o[665]) );
  XOR U4864 ( .A(n4861), .B(n4862), .Z(n2151) );
  IV U4865 ( .A(n2154), .Z(mod_mult_o[664]) );
  XOR U4866 ( .A(n4863), .B(n4864), .Z(n2154) );
  IV U4867 ( .A(n2157), .Z(mod_mult_o[663]) );
  XOR U4868 ( .A(n4865), .B(n4866), .Z(n2157) );
  IV U4869 ( .A(n2160), .Z(mod_mult_o[662]) );
  XOR U4870 ( .A(n4867), .B(n4868), .Z(n2160) );
  IV U4871 ( .A(n2163), .Z(mod_mult_o[661]) );
  XOR U4872 ( .A(n4869), .B(n4870), .Z(n2163) );
  IV U4873 ( .A(n2166), .Z(mod_mult_o[660]) );
  XOR U4874 ( .A(n4871), .B(n4872), .Z(n2166) );
  IV U4875 ( .A(n2169), .Z(mod_mult_o[65]) );
  XOR U4876 ( .A(n4873), .B(n4874), .Z(n2169) );
  IV U4877 ( .A(n2172), .Z(mod_mult_o[659]) );
  XOR U4878 ( .A(n4875), .B(n4876), .Z(n2172) );
  IV U4879 ( .A(n2175), .Z(mod_mult_o[658]) );
  XOR U4880 ( .A(n4877), .B(n4878), .Z(n2175) );
  IV U4881 ( .A(n2178), .Z(mod_mult_o[657]) );
  XOR U4882 ( .A(n4879), .B(n4880), .Z(n2178) );
  IV U4883 ( .A(n2181), .Z(mod_mult_o[656]) );
  XOR U4884 ( .A(n4881), .B(n4882), .Z(n2181) );
  IV U4885 ( .A(n2184), .Z(mod_mult_o[655]) );
  XOR U4886 ( .A(n4883), .B(n4884), .Z(n2184) );
  IV U4887 ( .A(n2187), .Z(mod_mult_o[654]) );
  XOR U4888 ( .A(n4885), .B(n4886), .Z(n2187) );
  IV U4889 ( .A(n2190), .Z(mod_mult_o[653]) );
  XOR U4890 ( .A(n4887), .B(n4888), .Z(n2190) );
  IV U4891 ( .A(n2193), .Z(mod_mult_o[652]) );
  XOR U4892 ( .A(n4889), .B(n4890), .Z(n2193) );
  IV U4893 ( .A(n2196), .Z(mod_mult_o[651]) );
  XOR U4894 ( .A(n4891), .B(n4892), .Z(n2196) );
  IV U4895 ( .A(n2199), .Z(mod_mult_o[650]) );
  XOR U4896 ( .A(n4893), .B(n4894), .Z(n2199) );
  IV U4897 ( .A(n2202), .Z(mod_mult_o[64]) );
  XOR U4898 ( .A(n4895), .B(n4896), .Z(n2202) );
  IV U4899 ( .A(n2205), .Z(mod_mult_o[649]) );
  XOR U4900 ( .A(n4897), .B(n4898), .Z(n2205) );
  IV U4901 ( .A(n2208), .Z(mod_mult_o[648]) );
  XOR U4902 ( .A(n4899), .B(n4900), .Z(n2208) );
  IV U4903 ( .A(n2211), .Z(mod_mult_o[647]) );
  XOR U4904 ( .A(n4901), .B(n4902), .Z(n2211) );
  IV U4905 ( .A(n2214), .Z(mod_mult_o[646]) );
  XOR U4906 ( .A(n4903), .B(n4904), .Z(n2214) );
  IV U4907 ( .A(n2217), .Z(mod_mult_o[645]) );
  XOR U4908 ( .A(n4905), .B(n4906), .Z(n2217) );
  IV U4909 ( .A(n2220), .Z(mod_mult_o[644]) );
  XOR U4910 ( .A(n4907), .B(n4908), .Z(n2220) );
  IV U4911 ( .A(n2223), .Z(mod_mult_o[643]) );
  XOR U4912 ( .A(n4909), .B(n4910), .Z(n2223) );
  IV U4913 ( .A(n2226), .Z(mod_mult_o[642]) );
  XOR U4914 ( .A(n4911), .B(n4912), .Z(n2226) );
  IV U4915 ( .A(n2229), .Z(mod_mult_o[641]) );
  XOR U4916 ( .A(n4913), .B(n4914), .Z(n2229) );
  IV U4917 ( .A(n2232), .Z(mod_mult_o[640]) );
  XOR U4918 ( .A(n4915), .B(n4916), .Z(n2232) );
  IV U4919 ( .A(n2235), .Z(mod_mult_o[63]) );
  XOR U4920 ( .A(n4917), .B(n4918), .Z(n2235) );
  IV U4921 ( .A(n2238), .Z(mod_mult_o[639]) );
  XOR U4922 ( .A(n4919), .B(n4920), .Z(n2238) );
  IV U4923 ( .A(n2241), .Z(mod_mult_o[638]) );
  XOR U4924 ( .A(n4921), .B(n4922), .Z(n2241) );
  IV U4925 ( .A(n2244), .Z(mod_mult_o[637]) );
  XOR U4926 ( .A(n4923), .B(n4924), .Z(n2244) );
  IV U4927 ( .A(n2247), .Z(mod_mult_o[636]) );
  XOR U4928 ( .A(n4925), .B(n4926), .Z(n2247) );
  IV U4929 ( .A(n2250), .Z(mod_mult_o[635]) );
  XOR U4930 ( .A(n4927), .B(n4928), .Z(n2250) );
  IV U4931 ( .A(n2253), .Z(mod_mult_o[634]) );
  XOR U4932 ( .A(n4929), .B(n4930), .Z(n2253) );
  IV U4933 ( .A(n2256), .Z(mod_mult_o[633]) );
  XOR U4934 ( .A(n4931), .B(n4932), .Z(n2256) );
  IV U4935 ( .A(n2259), .Z(mod_mult_o[632]) );
  XOR U4936 ( .A(n4933), .B(n4934), .Z(n2259) );
  IV U4937 ( .A(n2262), .Z(mod_mult_o[631]) );
  XOR U4938 ( .A(n4935), .B(n4936), .Z(n2262) );
  IV U4939 ( .A(n2265), .Z(mod_mult_o[630]) );
  XOR U4940 ( .A(n4937), .B(n4938), .Z(n2265) );
  IV U4941 ( .A(n2268), .Z(mod_mult_o[62]) );
  XOR U4942 ( .A(n4939), .B(n4940), .Z(n2268) );
  IV U4943 ( .A(n2271), .Z(mod_mult_o[629]) );
  XOR U4944 ( .A(n4941), .B(n4942), .Z(n2271) );
  IV U4945 ( .A(n2274), .Z(mod_mult_o[628]) );
  XOR U4946 ( .A(n4943), .B(n4944), .Z(n2274) );
  IV U4947 ( .A(n2277), .Z(mod_mult_o[627]) );
  XOR U4948 ( .A(n4945), .B(n4946), .Z(n2277) );
  IV U4949 ( .A(n2280), .Z(mod_mult_o[626]) );
  XOR U4950 ( .A(n4947), .B(n4948), .Z(n2280) );
  IV U4951 ( .A(n2283), .Z(mod_mult_o[625]) );
  XOR U4952 ( .A(n4949), .B(n4950), .Z(n2283) );
  IV U4953 ( .A(n2286), .Z(mod_mult_o[624]) );
  XOR U4954 ( .A(n4951), .B(n4952), .Z(n2286) );
  IV U4955 ( .A(n2289), .Z(mod_mult_o[623]) );
  XOR U4956 ( .A(n4953), .B(n4954), .Z(n2289) );
  IV U4957 ( .A(n2292), .Z(mod_mult_o[622]) );
  XOR U4958 ( .A(n4955), .B(n4956), .Z(n2292) );
  IV U4959 ( .A(n2295), .Z(mod_mult_o[621]) );
  XOR U4960 ( .A(n4957), .B(n4958), .Z(n2295) );
  IV U4961 ( .A(n2298), .Z(mod_mult_o[620]) );
  XOR U4962 ( .A(n4959), .B(n4960), .Z(n2298) );
  IV U4963 ( .A(n2301), .Z(mod_mult_o[61]) );
  XOR U4964 ( .A(n4961), .B(n4962), .Z(n2301) );
  IV U4965 ( .A(n2304), .Z(mod_mult_o[619]) );
  XOR U4966 ( .A(n4963), .B(n4964), .Z(n2304) );
  IV U4967 ( .A(n2307), .Z(mod_mult_o[618]) );
  XOR U4968 ( .A(n4965), .B(n4966), .Z(n2307) );
  IV U4969 ( .A(n2310), .Z(mod_mult_o[617]) );
  XOR U4970 ( .A(n4967), .B(n4968), .Z(n2310) );
  IV U4971 ( .A(n2313), .Z(mod_mult_o[616]) );
  XOR U4972 ( .A(n4969), .B(n4970), .Z(n2313) );
  IV U4973 ( .A(n2316), .Z(mod_mult_o[615]) );
  XOR U4974 ( .A(n4971), .B(n4972), .Z(n2316) );
  IV U4975 ( .A(n2319), .Z(mod_mult_o[614]) );
  XOR U4976 ( .A(n4973), .B(n4974), .Z(n2319) );
  IV U4977 ( .A(n2322), .Z(mod_mult_o[613]) );
  XOR U4978 ( .A(n4975), .B(n4976), .Z(n2322) );
  IV U4979 ( .A(n2325), .Z(mod_mult_o[612]) );
  XOR U4980 ( .A(n4977), .B(n4978), .Z(n2325) );
  IV U4981 ( .A(n2328), .Z(mod_mult_o[611]) );
  XOR U4982 ( .A(n4979), .B(n4980), .Z(n2328) );
  IV U4983 ( .A(n2331), .Z(mod_mult_o[610]) );
  XOR U4984 ( .A(n4981), .B(n4982), .Z(n2331) );
  IV U4985 ( .A(n2334), .Z(mod_mult_o[60]) );
  XOR U4986 ( .A(n4983), .B(n4984), .Z(n2334) );
  IV U4987 ( .A(n2337), .Z(mod_mult_o[609]) );
  XOR U4988 ( .A(n4985), .B(n4986), .Z(n2337) );
  IV U4989 ( .A(n2340), .Z(mod_mult_o[608]) );
  XOR U4990 ( .A(n4987), .B(n4988), .Z(n2340) );
  IV U4991 ( .A(n2343), .Z(mod_mult_o[607]) );
  XOR U4992 ( .A(n4989), .B(n4990), .Z(n2343) );
  IV U4993 ( .A(n2346), .Z(mod_mult_o[606]) );
  XOR U4994 ( .A(n4991), .B(n4992), .Z(n2346) );
  IV U4995 ( .A(n2349), .Z(mod_mult_o[605]) );
  XOR U4996 ( .A(n4993), .B(n4994), .Z(n2349) );
  IV U4997 ( .A(n2352), .Z(mod_mult_o[604]) );
  XOR U4998 ( .A(n4995), .B(n4996), .Z(n2352) );
  IV U4999 ( .A(n2355), .Z(mod_mult_o[603]) );
  XOR U5000 ( .A(n4997), .B(n4998), .Z(n2355) );
  IV U5001 ( .A(n2358), .Z(mod_mult_o[602]) );
  XOR U5002 ( .A(n4999), .B(n5000), .Z(n2358) );
  IV U5003 ( .A(n2361), .Z(mod_mult_o[601]) );
  XOR U5004 ( .A(n5001), .B(n5002), .Z(n2361) );
  IV U5005 ( .A(n2364), .Z(mod_mult_o[600]) );
  XOR U5006 ( .A(n5003), .B(n5004), .Z(n2364) );
  IV U5007 ( .A(n2367), .Z(mod_mult_o[5]) );
  XOR U5008 ( .A(n5005), .B(n5006), .Z(n2367) );
  IV U5009 ( .A(n2370), .Z(mod_mult_o[59]) );
  XOR U5010 ( .A(n5007), .B(n5008), .Z(n2370) );
  IV U5011 ( .A(n2373), .Z(mod_mult_o[599]) );
  XOR U5012 ( .A(n5009), .B(n5010), .Z(n2373) );
  IV U5013 ( .A(n2376), .Z(mod_mult_o[598]) );
  XOR U5014 ( .A(n5011), .B(n5012), .Z(n2376) );
  IV U5015 ( .A(n2379), .Z(mod_mult_o[597]) );
  XOR U5016 ( .A(n5013), .B(n5014), .Z(n2379) );
  IV U5017 ( .A(n2382), .Z(mod_mult_o[596]) );
  XOR U5018 ( .A(n5015), .B(n5016), .Z(n2382) );
  IV U5019 ( .A(n2385), .Z(mod_mult_o[595]) );
  XOR U5020 ( .A(n5017), .B(n5018), .Z(n2385) );
  IV U5021 ( .A(n2388), .Z(mod_mult_o[594]) );
  XOR U5022 ( .A(n5019), .B(n5020), .Z(n2388) );
  IV U5023 ( .A(n2391), .Z(mod_mult_o[593]) );
  XOR U5024 ( .A(n5021), .B(n5022), .Z(n2391) );
  IV U5025 ( .A(n2394), .Z(mod_mult_o[592]) );
  XOR U5026 ( .A(n5023), .B(n5024), .Z(n2394) );
  IV U5027 ( .A(n2397), .Z(mod_mult_o[591]) );
  XOR U5028 ( .A(n5025), .B(n5026), .Z(n2397) );
  IV U5029 ( .A(n2400), .Z(mod_mult_o[590]) );
  XOR U5030 ( .A(n5027), .B(n5028), .Z(n2400) );
  IV U5031 ( .A(n2403), .Z(mod_mult_o[58]) );
  XOR U5032 ( .A(n5029), .B(n5030), .Z(n2403) );
  IV U5033 ( .A(n2406), .Z(mod_mult_o[589]) );
  XOR U5034 ( .A(n5031), .B(n5032), .Z(n2406) );
  IV U5035 ( .A(n2409), .Z(mod_mult_o[588]) );
  XOR U5036 ( .A(n5033), .B(n5034), .Z(n2409) );
  IV U5037 ( .A(n2412), .Z(mod_mult_o[587]) );
  XOR U5038 ( .A(n5035), .B(n5036), .Z(n2412) );
  IV U5039 ( .A(n2415), .Z(mod_mult_o[586]) );
  XOR U5040 ( .A(n5037), .B(n5038), .Z(n2415) );
  IV U5041 ( .A(n2418), .Z(mod_mult_o[585]) );
  XOR U5042 ( .A(n5039), .B(n5040), .Z(n2418) );
  IV U5043 ( .A(n2421), .Z(mod_mult_o[584]) );
  XOR U5044 ( .A(n5041), .B(n5042), .Z(n2421) );
  IV U5045 ( .A(n2424), .Z(mod_mult_o[583]) );
  XOR U5046 ( .A(n5043), .B(n5044), .Z(n2424) );
  IV U5047 ( .A(n2427), .Z(mod_mult_o[582]) );
  XOR U5048 ( .A(n5045), .B(n5046), .Z(n2427) );
  IV U5049 ( .A(n2430), .Z(mod_mult_o[581]) );
  XOR U5050 ( .A(n5047), .B(n5048), .Z(n2430) );
  IV U5051 ( .A(n2433), .Z(mod_mult_o[580]) );
  XOR U5052 ( .A(n5049), .B(n5050), .Z(n2433) );
  IV U5053 ( .A(n2436), .Z(mod_mult_o[57]) );
  XOR U5054 ( .A(n5051), .B(n5052), .Z(n2436) );
  IV U5055 ( .A(n2439), .Z(mod_mult_o[579]) );
  XOR U5056 ( .A(n5053), .B(n5054), .Z(n2439) );
  IV U5057 ( .A(n2442), .Z(mod_mult_o[578]) );
  XOR U5058 ( .A(n5055), .B(n5056), .Z(n2442) );
  IV U5059 ( .A(n2445), .Z(mod_mult_o[577]) );
  XOR U5060 ( .A(n5057), .B(n5058), .Z(n2445) );
  IV U5061 ( .A(n2448), .Z(mod_mult_o[576]) );
  XOR U5062 ( .A(n5059), .B(n5060), .Z(n2448) );
  IV U5063 ( .A(n2451), .Z(mod_mult_o[575]) );
  XOR U5064 ( .A(n5061), .B(n5062), .Z(n2451) );
  IV U5065 ( .A(n2454), .Z(mod_mult_o[574]) );
  XOR U5066 ( .A(n5063), .B(n5064), .Z(n2454) );
  IV U5067 ( .A(n2457), .Z(mod_mult_o[573]) );
  XOR U5068 ( .A(n5065), .B(n5066), .Z(n2457) );
  IV U5069 ( .A(n2460), .Z(mod_mult_o[572]) );
  XOR U5070 ( .A(n5067), .B(n5068), .Z(n2460) );
  IV U5071 ( .A(n2463), .Z(mod_mult_o[571]) );
  XOR U5072 ( .A(n5069), .B(n5070), .Z(n2463) );
  IV U5073 ( .A(n2466), .Z(mod_mult_o[570]) );
  XOR U5074 ( .A(n5071), .B(n5072), .Z(n2466) );
  IV U5075 ( .A(n2469), .Z(mod_mult_o[56]) );
  XOR U5076 ( .A(n5073), .B(n5074), .Z(n2469) );
  IV U5077 ( .A(n2472), .Z(mod_mult_o[569]) );
  XOR U5078 ( .A(n5075), .B(n5076), .Z(n2472) );
  IV U5079 ( .A(n2475), .Z(mod_mult_o[568]) );
  XOR U5080 ( .A(n5077), .B(n5078), .Z(n2475) );
  IV U5081 ( .A(n2478), .Z(mod_mult_o[567]) );
  XOR U5082 ( .A(n5079), .B(n5080), .Z(n2478) );
  IV U5083 ( .A(n2481), .Z(mod_mult_o[566]) );
  XOR U5084 ( .A(n5081), .B(n5082), .Z(n2481) );
  IV U5085 ( .A(n2484), .Z(mod_mult_o[565]) );
  XOR U5086 ( .A(n5083), .B(n5084), .Z(n2484) );
  IV U5087 ( .A(n2487), .Z(mod_mult_o[564]) );
  XOR U5088 ( .A(n5085), .B(n5086), .Z(n2487) );
  IV U5089 ( .A(n2490), .Z(mod_mult_o[563]) );
  XOR U5090 ( .A(n5087), .B(n5088), .Z(n2490) );
  IV U5091 ( .A(n2493), .Z(mod_mult_o[562]) );
  XOR U5092 ( .A(n5089), .B(n5090), .Z(n2493) );
  IV U5093 ( .A(n2496), .Z(mod_mult_o[561]) );
  XOR U5094 ( .A(n5091), .B(n5092), .Z(n2496) );
  IV U5095 ( .A(n2499), .Z(mod_mult_o[560]) );
  XOR U5096 ( .A(n5093), .B(n5094), .Z(n2499) );
  IV U5097 ( .A(n2502), .Z(mod_mult_o[55]) );
  XOR U5098 ( .A(n5095), .B(n5096), .Z(n2502) );
  IV U5099 ( .A(n2505), .Z(mod_mult_o[559]) );
  XOR U5100 ( .A(n5097), .B(n5098), .Z(n2505) );
  IV U5101 ( .A(n2508), .Z(mod_mult_o[558]) );
  XOR U5102 ( .A(n5099), .B(n5100), .Z(n2508) );
  IV U5103 ( .A(n2511), .Z(mod_mult_o[557]) );
  XOR U5104 ( .A(n5101), .B(n5102), .Z(n2511) );
  IV U5105 ( .A(n2514), .Z(mod_mult_o[556]) );
  XOR U5106 ( .A(n5103), .B(n5104), .Z(n2514) );
  IV U5107 ( .A(n2517), .Z(mod_mult_o[555]) );
  XOR U5108 ( .A(n5105), .B(n5106), .Z(n2517) );
  IV U5109 ( .A(n2520), .Z(mod_mult_o[554]) );
  XOR U5110 ( .A(n5107), .B(n5108), .Z(n2520) );
  IV U5111 ( .A(n2523), .Z(mod_mult_o[553]) );
  XOR U5112 ( .A(n5109), .B(n5110), .Z(n2523) );
  IV U5113 ( .A(n2526), .Z(mod_mult_o[552]) );
  XOR U5114 ( .A(n5111), .B(n5112), .Z(n2526) );
  IV U5115 ( .A(n2529), .Z(mod_mult_o[551]) );
  XOR U5116 ( .A(n5113), .B(n5114), .Z(n2529) );
  IV U5117 ( .A(n2532), .Z(mod_mult_o[550]) );
  XOR U5118 ( .A(n5115), .B(n5116), .Z(n2532) );
  IV U5119 ( .A(n2535), .Z(mod_mult_o[54]) );
  XOR U5120 ( .A(n5117), .B(n5118), .Z(n2535) );
  IV U5121 ( .A(n2538), .Z(mod_mult_o[549]) );
  XOR U5122 ( .A(n5119), .B(n5120), .Z(n2538) );
  IV U5123 ( .A(n2541), .Z(mod_mult_o[548]) );
  XOR U5124 ( .A(n5121), .B(n5122), .Z(n2541) );
  IV U5125 ( .A(n2544), .Z(mod_mult_o[547]) );
  XOR U5126 ( .A(n5123), .B(n5124), .Z(n2544) );
  IV U5127 ( .A(n2547), .Z(mod_mult_o[546]) );
  XOR U5128 ( .A(n5125), .B(n5126), .Z(n2547) );
  IV U5129 ( .A(n2550), .Z(mod_mult_o[545]) );
  XOR U5130 ( .A(n5127), .B(n5128), .Z(n2550) );
  IV U5131 ( .A(n2553), .Z(mod_mult_o[544]) );
  XOR U5132 ( .A(n5129), .B(n5130), .Z(n2553) );
  IV U5133 ( .A(n2556), .Z(mod_mult_o[543]) );
  XOR U5134 ( .A(n5131), .B(n5132), .Z(n2556) );
  IV U5135 ( .A(n2559), .Z(mod_mult_o[542]) );
  XOR U5136 ( .A(n5133), .B(n5134), .Z(n2559) );
  IV U5137 ( .A(n2562), .Z(mod_mult_o[541]) );
  XOR U5138 ( .A(n5135), .B(n5136), .Z(n2562) );
  IV U5139 ( .A(n2565), .Z(mod_mult_o[540]) );
  XOR U5140 ( .A(n5137), .B(n5138), .Z(n2565) );
  IV U5141 ( .A(n2568), .Z(mod_mult_o[53]) );
  XOR U5142 ( .A(n5139), .B(n5140), .Z(n2568) );
  IV U5143 ( .A(n2571), .Z(mod_mult_o[539]) );
  XOR U5144 ( .A(n5141), .B(n5142), .Z(n2571) );
  IV U5145 ( .A(n2574), .Z(mod_mult_o[538]) );
  XOR U5146 ( .A(n5143), .B(n5144), .Z(n2574) );
  IV U5147 ( .A(n2577), .Z(mod_mult_o[537]) );
  XOR U5148 ( .A(n5145), .B(n5146), .Z(n2577) );
  IV U5149 ( .A(n2580), .Z(mod_mult_o[536]) );
  XOR U5150 ( .A(n5147), .B(n5148), .Z(n2580) );
  IV U5151 ( .A(n2583), .Z(mod_mult_o[535]) );
  XOR U5152 ( .A(n5149), .B(n5150), .Z(n2583) );
  IV U5153 ( .A(n2586), .Z(mod_mult_o[534]) );
  XOR U5154 ( .A(n5151), .B(n5152), .Z(n2586) );
  IV U5155 ( .A(n2589), .Z(mod_mult_o[533]) );
  XOR U5156 ( .A(n5153), .B(n5154), .Z(n2589) );
  IV U5157 ( .A(n2592), .Z(mod_mult_o[532]) );
  XOR U5158 ( .A(n5155), .B(n5156), .Z(n2592) );
  IV U5159 ( .A(n2595), .Z(mod_mult_o[531]) );
  XOR U5160 ( .A(n5157), .B(n5158), .Z(n2595) );
  IV U5161 ( .A(n2598), .Z(mod_mult_o[530]) );
  XOR U5162 ( .A(n5159), .B(n5160), .Z(n2598) );
  IV U5163 ( .A(n2601), .Z(mod_mult_o[52]) );
  XOR U5164 ( .A(n5161), .B(n5162), .Z(n2601) );
  IV U5165 ( .A(n2604), .Z(mod_mult_o[529]) );
  XOR U5166 ( .A(n5163), .B(n5164), .Z(n2604) );
  IV U5167 ( .A(n2607), .Z(mod_mult_o[528]) );
  XOR U5168 ( .A(n5165), .B(n5166), .Z(n2607) );
  IV U5169 ( .A(n2610), .Z(mod_mult_o[527]) );
  XOR U5170 ( .A(n5167), .B(n5168), .Z(n2610) );
  IV U5171 ( .A(n2613), .Z(mod_mult_o[526]) );
  XOR U5172 ( .A(n5169), .B(n5170), .Z(n2613) );
  IV U5173 ( .A(n2616), .Z(mod_mult_o[525]) );
  XOR U5174 ( .A(n5171), .B(n5172), .Z(n2616) );
  IV U5175 ( .A(n2619), .Z(mod_mult_o[524]) );
  XOR U5176 ( .A(n5173), .B(n5174), .Z(n2619) );
  IV U5177 ( .A(n2622), .Z(mod_mult_o[523]) );
  XOR U5178 ( .A(n5175), .B(n5176), .Z(n2622) );
  IV U5179 ( .A(n2625), .Z(mod_mult_o[522]) );
  XOR U5180 ( .A(n5177), .B(n5178), .Z(n2625) );
  IV U5181 ( .A(n2628), .Z(mod_mult_o[521]) );
  XOR U5182 ( .A(n5179), .B(n5180), .Z(n2628) );
  IV U5183 ( .A(n2631), .Z(mod_mult_o[520]) );
  XOR U5184 ( .A(n5181), .B(n5182), .Z(n2631) );
  IV U5185 ( .A(n2634), .Z(mod_mult_o[51]) );
  XOR U5186 ( .A(n5183), .B(n5184), .Z(n2634) );
  IV U5187 ( .A(n2637), .Z(mod_mult_o[519]) );
  XOR U5188 ( .A(n5185), .B(n5186), .Z(n2637) );
  IV U5189 ( .A(n2640), .Z(mod_mult_o[518]) );
  XOR U5190 ( .A(n5187), .B(n5188), .Z(n2640) );
  IV U5191 ( .A(n2643), .Z(mod_mult_o[517]) );
  XOR U5192 ( .A(n5189), .B(n5190), .Z(n2643) );
  IV U5193 ( .A(n2646), .Z(mod_mult_o[516]) );
  XOR U5194 ( .A(n5191), .B(n5192), .Z(n2646) );
  IV U5195 ( .A(n2649), .Z(mod_mult_o[515]) );
  XOR U5196 ( .A(n5193), .B(n5194), .Z(n2649) );
  IV U5197 ( .A(n2652), .Z(mod_mult_o[514]) );
  XOR U5198 ( .A(n5195), .B(n5196), .Z(n2652) );
  IV U5199 ( .A(n2655), .Z(mod_mult_o[513]) );
  XOR U5200 ( .A(n5197), .B(n5198), .Z(n2655) );
  IV U5201 ( .A(n2658), .Z(mod_mult_o[512]) );
  XOR U5202 ( .A(n5199), .B(n5200), .Z(n2658) );
  IV U5203 ( .A(n2661), .Z(mod_mult_o[511]) );
  XOR U5204 ( .A(n5201), .B(n5202), .Z(n2661) );
  IV U5205 ( .A(n2664), .Z(mod_mult_o[510]) );
  XOR U5206 ( .A(n5203), .B(n5204), .Z(n2664) );
  IV U5207 ( .A(n2667), .Z(mod_mult_o[50]) );
  XOR U5208 ( .A(n5205), .B(n5206), .Z(n2667) );
  IV U5209 ( .A(n2670), .Z(mod_mult_o[509]) );
  XOR U5210 ( .A(n5207), .B(n5208), .Z(n2670) );
  IV U5211 ( .A(n2673), .Z(mod_mult_o[508]) );
  XOR U5212 ( .A(n5209), .B(n5210), .Z(n2673) );
  IV U5213 ( .A(n2676), .Z(mod_mult_o[507]) );
  XOR U5214 ( .A(n5211), .B(n5212), .Z(n2676) );
  IV U5215 ( .A(n2679), .Z(mod_mult_o[506]) );
  XOR U5216 ( .A(n5213), .B(n5214), .Z(n2679) );
  IV U5217 ( .A(n2682), .Z(mod_mult_o[505]) );
  XOR U5218 ( .A(n5215), .B(n5216), .Z(n2682) );
  IV U5219 ( .A(n2685), .Z(mod_mult_o[504]) );
  XOR U5220 ( .A(n5217), .B(n5218), .Z(n2685) );
  IV U5221 ( .A(n2688), .Z(mod_mult_o[503]) );
  XOR U5222 ( .A(n5219), .B(n5220), .Z(n2688) );
  IV U5223 ( .A(n2691), .Z(mod_mult_o[502]) );
  XOR U5224 ( .A(n5221), .B(n5222), .Z(n2691) );
  IV U5225 ( .A(n2694), .Z(mod_mult_o[501]) );
  XOR U5226 ( .A(n5223), .B(n5224), .Z(n2694) );
  IV U5227 ( .A(n2697), .Z(mod_mult_o[500]) );
  XOR U5228 ( .A(n5225), .B(n5226), .Z(n2697) );
  IV U5229 ( .A(n2700), .Z(mod_mult_o[4]) );
  XOR U5230 ( .A(n5227), .B(n5228), .Z(n2700) );
  IV U5231 ( .A(n2703), .Z(mod_mult_o[49]) );
  XOR U5232 ( .A(n5229), .B(n5230), .Z(n2703) );
  IV U5233 ( .A(n2706), .Z(mod_mult_o[499]) );
  XOR U5234 ( .A(n5231), .B(n5232), .Z(n2706) );
  IV U5235 ( .A(n2709), .Z(mod_mult_o[498]) );
  XOR U5236 ( .A(n5233), .B(n5234), .Z(n2709) );
  IV U5237 ( .A(n2712), .Z(mod_mult_o[497]) );
  XOR U5238 ( .A(n5235), .B(n5236), .Z(n2712) );
  IV U5239 ( .A(n2715), .Z(mod_mult_o[496]) );
  XOR U5240 ( .A(n5237), .B(n5238), .Z(n2715) );
  IV U5241 ( .A(n2718), .Z(mod_mult_o[495]) );
  XOR U5242 ( .A(n5239), .B(n5240), .Z(n2718) );
  IV U5243 ( .A(n2721), .Z(mod_mult_o[494]) );
  XOR U5244 ( .A(n5241), .B(n5242), .Z(n2721) );
  IV U5245 ( .A(n2724), .Z(mod_mult_o[493]) );
  XOR U5246 ( .A(n5243), .B(n5244), .Z(n2724) );
  IV U5247 ( .A(n2727), .Z(mod_mult_o[492]) );
  XOR U5248 ( .A(n5245), .B(n5246), .Z(n2727) );
  IV U5249 ( .A(n2730), .Z(mod_mult_o[491]) );
  XOR U5250 ( .A(n5247), .B(n5248), .Z(n2730) );
  IV U5251 ( .A(n2733), .Z(mod_mult_o[490]) );
  XOR U5252 ( .A(n5249), .B(n5250), .Z(n2733) );
  IV U5253 ( .A(n2736), .Z(mod_mult_o[48]) );
  XOR U5254 ( .A(n5251), .B(n5252), .Z(n2736) );
  IV U5255 ( .A(n2739), .Z(mod_mult_o[489]) );
  XOR U5256 ( .A(n5253), .B(n5254), .Z(n2739) );
  IV U5257 ( .A(n2742), .Z(mod_mult_o[488]) );
  XOR U5258 ( .A(n5255), .B(n5256), .Z(n2742) );
  IV U5259 ( .A(n2745), .Z(mod_mult_o[487]) );
  XOR U5260 ( .A(n5257), .B(n5258), .Z(n2745) );
  IV U5261 ( .A(n2748), .Z(mod_mult_o[486]) );
  XOR U5262 ( .A(n5259), .B(n5260), .Z(n2748) );
  IV U5263 ( .A(n2751), .Z(mod_mult_o[485]) );
  XOR U5264 ( .A(n5261), .B(n5262), .Z(n2751) );
  IV U5265 ( .A(n2754), .Z(mod_mult_o[484]) );
  XOR U5266 ( .A(n5263), .B(n5264), .Z(n2754) );
  IV U5267 ( .A(n2757), .Z(mod_mult_o[483]) );
  XOR U5268 ( .A(n5265), .B(n5266), .Z(n2757) );
  IV U5269 ( .A(n2760), .Z(mod_mult_o[482]) );
  XOR U5270 ( .A(n5267), .B(n5268), .Z(n2760) );
  IV U5271 ( .A(n2763), .Z(mod_mult_o[481]) );
  XOR U5272 ( .A(n5269), .B(n5270), .Z(n2763) );
  IV U5273 ( .A(n2766), .Z(mod_mult_o[480]) );
  XOR U5274 ( .A(n5271), .B(n5272), .Z(n2766) );
  IV U5275 ( .A(n2769), .Z(mod_mult_o[47]) );
  XOR U5276 ( .A(n5273), .B(n5274), .Z(n2769) );
  IV U5277 ( .A(n2772), .Z(mod_mult_o[479]) );
  XOR U5278 ( .A(n5275), .B(n5276), .Z(n2772) );
  IV U5279 ( .A(n2775), .Z(mod_mult_o[478]) );
  XOR U5280 ( .A(n5277), .B(n5278), .Z(n2775) );
  IV U5281 ( .A(n2778), .Z(mod_mult_o[477]) );
  XOR U5282 ( .A(n5279), .B(n5280), .Z(n2778) );
  IV U5283 ( .A(n2781), .Z(mod_mult_o[476]) );
  XOR U5284 ( .A(n5281), .B(n5282), .Z(n2781) );
  IV U5285 ( .A(n2784), .Z(mod_mult_o[475]) );
  XOR U5286 ( .A(n5283), .B(n5284), .Z(n2784) );
  IV U5287 ( .A(n2787), .Z(mod_mult_o[474]) );
  XOR U5288 ( .A(n5285), .B(n5286), .Z(n2787) );
  IV U5289 ( .A(n2790), .Z(mod_mult_o[473]) );
  XOR U5290 ( .A(n5287), .B(n5288), .Z(n2790) );
  IV U5291 ( .A(n2793), .Z(mod_mult_o[472]) );
  XOR U5292 ( .A(n5289), .B(n5290), .Z(n2793) );
  IV U5293 ( .A(n2796), .Z(mod_mult_o[471]) );
  XOR U5294 ( .A(n5291), .B(n5292), .Z(n2796) );
  IV U5295 ( .A(n2799), .Z(mod_mult_o[470]) );
  XOR U5296 ( .A(n5293), .B(n5294), .Z(n2799) );
  IV U5297 ( .A(n2802), .Z(mod_mult_o[46]) );
  XOR U5298 ( .A(n5295), .B(n5296), .Z(n2802) );
  IV U5299 ( .A(n2805), .Z(mod_mult_o[469]) );
  XOR U5300 ( .A(n5297), .B(n5298), .Z(n2805) );
  IV U5301 ( .A(n2808), .Z(mod_mult_o[468]) );
  XOR U5302 ( .A(n5299), .B(n5300), .Z(n2808) );
  IV U5303 ( .A(n2811), .Z(mod_mult_o[467]) );
  XOR U5304 ( .A(n5301), .B(n5302), .Z(n2811) );
  IV U5305 ( .A(n2814), .Z(mod_mult_o[466]) );
  XOR U5306 ( .A(n5303), .B(n5304), .Z(n2814) );
  IV U5307 ( .A(n2817), .Z(mod_mult_o[465]) );
  XOR U5308 ( .A(n5305), .B(n5306), .Z(n2817) );
  IV U5309 ( .A(n2820), .Z(mod_mult_o[464]) );
  XOR U5310 ( .A(n5307), .B(n5308), .Z(n2820) );
  IV U5311 ( .A(n2823), .Z(mod_mult_o[463]) );
  XOR U5312 ( .A(n5309), .B(n5310), .Z(n2823) );
  IV U5313 ( .A(n2826), .Z(mod_mult_o[462]) );
  XOR U5314 ( .A(n5311), .B(n5312), .Z(n2826) );
  IV U5315 ( .A(n2829), .Z(mod_mult_o[461]) );
  XOR U5316 ( .A(n5313), .B(n5314), .Z(n2829) );
  IV U5317 ( .A(n2832), .Z(mod_mult_o[460]) );
  XOR U5318 ( .A(n5315), .B(n5316), .Z(n2832) );
  IV U5319 ( .A(n2835), .Z(mod_mult_o[45]) );
  XOR U5320 ( .A(n5317), .B(n5318), .Z(n2835) );
  IV U5321 ( .A(n2838), .Z(mod_mult_o[459]) );
  XOR U5322 ( .A(n5319), .B(n5320), .Z(n2838) );
  IV U5323 ( .A(n2841), .Z(mod_mult_o[458]) );
  XOR U5324 ( .A(n5321), .B(n5322), .Z(n2841) );
  IV U5325 ( .A(n2844), .Z(mod_mult_o[457]) );
  XOR U5326 ( .A(n5323), .B(n5324), .Z(n2844) );
  IV U5327 ( .A(n2847), .Z(mod_mult_o[456]) );
  XOR U5328 ( .A(n5325), .B(n5326), .Z(n2847) );
  IV U5329 ( .A(n2850), .Z(mod_mult_o[455]) );
  XOR U5330 ( .A(n5327), .B(n5328), .Z(n2850) );
  IV U5331 ( .A(n2853), .Z(mod_mult_o[454]) );
  XOR U5332 ( .A(n5329), .B(n5330), .Z(n2853) );
  IV U5333 ( .A(n2856), .Z(mod_mult_o[453]) );
  XOR U5334 ( .A(n5331), .B(n5332), .Z(n2856) );
  IV U5335 ( .A(n2859), .Z(mod_mult_o[452]) );
  XOR U5336 ( .A(n5333), .B(n5334), .Z(n2859) );
  IV U5337 ( .A(n2862), .Z(mod_mult_o[451]) );
  XOR U5338 ( .A(n5335), .B(n5336), .Z(n2862) );
  IV U5339 ( .A(n2865), .Z(mod_mult_o[450]) );
  XOR U5340 ( .A(n5337), .B(n5338), .Z(n2865) );
  IV U5341 ( .A(n2868), .Z(mod_mult_o[44]) );
  XOR U5342 ( .A(n5339), .B(n5340), .Z(n2868) );
  IV U5343 ( .A(n2871), .Z(mod_mult_o[449]) );
  XOR U5344 ( .A(n5341), .B(n5342), .Z(n2871) );
  IV U5345 ( .A(n2874), .Z(mod_mult_o[448]) );
  XOR U5346 ( .A(n5343), .B(n5344), .Z(n2874) );
  IV U5347 ( .A(n2877), .Z(mod_mult_o[447]) );
  XOR U5348 ( .A(n5345), .B(n5346), .Z(n2877) );
  IV U5349 ( .A(n2880), .Z(mod_mult_o[446]) );
  XOR U5350 ( .A(n5347), .B(n5348), .Z(n2880) );
  IV U5351 ( .A(n2883), .Z(mod_mult_o[445]) );
  XOR U5352 ( .A(n5349), .B(n5350), .Z(n2883) );
  IV U5353 ( .A(n2886), .Z(mod_mult_o[444]) );
  XOR U5354 ( .A(n5351), .B(n5352), .Z(n2886) );
  IV U5355 ( .A(n2889), .Z(mod_mult_o[443]) );
  XOR U5356 ( .A(n5353), .B(n5354), .Z(n2889) );
  IV U5357 ( .A(n2892), .Z(mod_mult_o[442]) );
  XOR U5358 ( .A(n5355), .B(n5356), .Z(n2892) );
  IV U5359 ( .A(n2895), .Z(mod_mult_o[441]) );
  XOR U5360 ( .A(n5357), .B(n5358), .Z(n2895) );
  IV U5361 ( .A(n2898), .Z(mod_mult_o[440]) );
  XOR U5362 ( .A(n5359), .B(n5360), .Z(n2898) );
  IV U5363 ( .A(n2901), .Z(mod_mult_o[43]) );
  XOR U5364 ( .A(n5361), .B(n5362), .Z(n2901) );
  IV U5365 ( .A(n2904), .Z(mod_mult_o[439]) );
  XOR U5366 ( .A(n5363), .B(n5364), .Z(n2904) );
  IV U5367 ( .A(n2907), .Z(mod_mult_o[438]) );
  XOR U5368 ( .A(n5365), .B(n5366), .Z(n2907) );
  IV U5369 ( .A(n2910), .Z(mod_mult_o[437]) );
  XOR U5370 ( .A(n5367), .B(n5368), .Z(n2910) );
  IV U5371 ( .A(n2913), .Z(mod_mult_o[436]) );
  XOR U5372 ( .A(n5369), .B(n5370), .Z(n2913) );
  IV U5373 ( .A(n2916), .Z(mod_mult_o[435]) );
  XOR U5374 ( .A(n5371), .B(n5372), .Z(n2916) );
  IV U5375 ( .A(n2919), .Z(mod_mult_o[434]) );
  XOR U5376 ( .A(n5373), .B(n5374), .Z(n2919) );
  IV U5377 ( .A(n2922), .Z(mod_mult_o[433]) );
  XOR U5378 ( .A(n5375), .B(n5376), .Z(n2922) );
  IV U5379 ( .A(n2925), .Z(mod_mult_o[432]) );
  XOR U5380 ( .A(n5377), .B(n5378), .Z(n2925) );
  IV U5381 ( .A(n2928), .Z(mod_mult_o[431]) );
  XOR U5382 ( .A(n5379), .B(n5380), .Z(n2928) );
  IV U5383 ( .A(n2931), .Z(mod_mult_o[430]) );
  XOR U5384 ( .A(n5381), .B(n5382), .Z(n2931) );
  IV U5385 ( .A(n2934), .Z(mod_mult_o[42]) );
  XOR U5386 ( .A(n5383), .B(n5384), .Z(n2934) );
  IV U5387 ( .A(n2937), .Z(mod_mult_o[429]) );
  XOR U5388 ( .A(n5385), .B(n5386), .Z(n2937) );
  IV U5389 ( .A(n2940), .Z(mod_mult_o[428]) );
  XOR U5390 ( .A(n5387), .B(n5388), .Z(n2940) );
  IV U5391 ( .A(n2943), .Z(mod_mult_o[427]) );
  XOR U5392 ( .A(n5389), .B(n5390), .Z(n2943) );
  IV U5393 ( .A(n2946), .Z(mod_mult_o[426]) );
  XOR U5394 ( .A(n5391), .B(n5392), .Z(n2946) );
  IV U5395 ( .A(n2949), .Z(mod_mult_o[425]) );
  XOR U5396 ( .A(n5393), .B(n5394), .Z(n2949) );
  IV U5397 ( .A(n2952), .Z(mod_mult_o[424]) );
  XOR U5398 ( .A(n5395), .B(n5396), .Z(n2952) );
  IV U5399 ( .A(n2955), .Z(mod_mult_o[423]) );
  XOR U5400 ( .A(n5397), .B(n5398), .Z(n2955) );
  IV U5401 ( .A(n2958), .Z(mod_mult_o[422]) );
  XOR U5402 ( .A(n5399), .B(n5400), .Z(n2958) );
  IV U5403 ( .A(n2961), .Z(mod_mult_o[421]) );
  XOR U5404 ( .A(n5401), .B(n5402), .Z(n2961) );
  IV U5405 ( .A(n2964), .Z(mod_mult_o[420]) );
  XOR U5406 ( .A(n5403), .B(n5404), .Z(n2964) );
  IV U5407 ( .A(n2967), .Z(mod_mult_o[41]) );
  XOR U5408 ( .A(n5405), .B(n5406), .Z(n2967) );
  IV U5409 ( .A(n2970), .Z(mod_mult_o[419]) );
  XOR U5410 ( .A(n5407), .B(n5408), .Z(n2970) );
  IV U5411 ( .A(n2973), .Z(mod_mult_o[418]) );
  XOR U5412 ( .A(n5409), .B(n5410), .Z(n2973) );
  IV U5413 ( .A(n2976), .Z(mod_mult_o[417]) );
  XOR U5414 ( .A(n5411), .B(n5412), .Z(n2976) );
  IV U5415 ( .A(n2979), .Z(mod_mult_o[416]) );
  XOR U5416 ( .A(n5413), .B(n5414), .Z(n2979) );
  IV U5417 ( .A(n2982), .Z(mod_mult_o[415]) );
  XOR U5418 ( .A(n5415), .B(n5416), .Z(n2982) );
  IV U5419 ( .A(n2985), .Z(mod_mult_o[414]) );
  XOR U5420 ( .A(n5417), .B(n5418), .Z(n2985) );
  IV U5421 ( .A(n2988), .Z(mod_mult_o[413]) );
  XOR U5422 ( .A(n5419), .B(n5420), .Z(n2988) );
  IV U5423 ( .A(n2991), .Z(mod_mult_o[412]) );
  XOR U5424 ( .A(n5421), .B(n5422), .Z(n2991) );
  IV U5425 ( .A(n2994), .Z(mod_mult_o[411]) );
  XOR U5426 ( .A(n5423), .B(n5424), .Z(n2994) );
  IV U5427 ( .A(n2997), .Z(mod_mult_o[410]) );
  XOR U5428 ( .A(n5425), .B(n5426), .Z(n2997) );
  IV U5429 ( .A(n3000), .Z(mod_mult_o[40]) );
  XOR U5430 ( .A(n5427), .B(n5428), .Z(n3000) );
  IV U5431 ( .A(n3003), .Z(mod_mult_o[409]) );
  XOR U5432 ( .A(n5429), .B(n5430), .Z(n3003) );
  IV U5433 ( .A(n3006), .Z(mod_mult_o[408]) );
  XOR U5434 ( .A(n5431), .B(n5432), .Z(n3006) );
  IV U5435 ( .A(n3009), .Z(mod_mult_o[407]) );
  XOR U5436 ( .A(n5433), .B(n5434), .Z(n3009) );
  IV U5437 ( .A(n3012), .Z(mod_mult_o[406]) );
  XOR U5438 ( .A(n5435), .B(n5436), .Z(n3012) );
  IV U5439 ( .A(n3015), .Z(mod_mult_o[405]) );
  XOR U5440 ( .A(n5437), .B(n5438), .Z(n3015) );
  IV U5441 ( .A(n3018), .Z(mod_mult_o[404]) );
  XOR U5442 ( .A(n5439), .B(n5440), .Z(n3018) );
  IV U5443 ( .A(n3021), .Z(mod_mult_o[403]) );
  XOR U5444 ( .A(n5441), .B(n5442), .Z(n3021) );
  IV U5445 ( .A(n3024), .Z(mod_mult_o[402]) );
  XOR U5446 ( .A(n5443), .B(n5444), .Z(n3024) );
  IV U5447 ( .A(n3027), .Z(mod_mult_o[401]) );
  XOR U5448 ( .A(n5445), .B(n5446), .Z(n3027) );
  IV U5449 ( .A(n3030), .Z(mod_mult_o[400]) );
  XOR U5450 ( .A(n5447), .B(n5448), .Z(n3030) );
  IV U5451 ( .A(n3033), .Z(mod_mult_o[3]) );
  XOR U5452 ( .A(n5449), .B(n5450), .Z(n3033) );
  IV U5453 ( .A(n3036), .Z(mod_mult_o[39]) );
  XOR U5454 ( .A(n5451), .B(n5452), .Z(n3036) );
  IV U5455 ( .A(n3039), .Z(mod_mult_o[399]) );
  XOR U5456 ( .A(n5453), .B(n5454), .Z(n3039) );
  IV U5457 ( .A(n3042), .Z(mod_mult_o[398]) );
  XOR U5458 ( .A(n5455), .B(n5456), .Z(n3042) );
  IV U5459 ( .A(n3045), .Z(mod_mult_o[397]) );
  XOR U5460 ( .A(n5457), .B(n5458), .Z(n3045) );
  IV U5461 ( .A(n3048), .Z(mod_mult_o[396]) );
  XOR U5462 ( .A(n5459), .B(n5460), .Z(n3048) );
  IV U5463 ( .A(n3051), .Z(mod_mult_o[395]) );
  XOR U5464 ( .A(n5461), .B(n5462), .Z(n3051) );
  IV U5465 ( .A(n3054), .Z(mod_mult_o[394]) );
  XOR U5466 ( .A(n5463), .B(n5464), .Z(n3054) );
  IV U5467 ( .A(n3057), .Z(mod_mult_o[393]) );
  XOR U5468 ( .A(n5465), .B(n5466), .Z(n3057) );
  IV U5469 ( .A(n3060), .Z(mod_mult_o[392]) );
  XOR U5470 ( .A(n5467), .B(n5468), .Z(n3060) );
  IV U5471 ( .A(n3063), .Z(mod_mult_o[391]) );
  XOR U5472 ( .A(n5469), .B(n5470), .Z(n3063) );
  IV U5473 ( .A(n3066), .Z(mod_mult_o[390]) );
  XOR U5474 ( .A(n5471), .B(n5472), .Z(n3066) );
  IV U5475 ( .A(n3069), .Z(mod_mult_o[38]) );
  XOR U5476 ( .A(n5473), .B(n5474), .Z(n3069) );
  IV U5477 ( .A(n3072), .Z(mod_mult_o[389]) );
  XOR U5478 ( .A(n5475), .B(n5476), .Z(n3072) );
  IV U5479 ( .A(n3075), .Z(mod_mult_o[388]) );
  XOR U5480 ( .A(n5477), .B(n5478), .Z(n3075) );
  IV U5481 ( .A(n3078), .Z(mod_mult_o[387]) );
  XOR U5482 ( .A(n5479), .B(n5480), .Z(n3078) );
  IV U5483 ( .A(n3081), .Z(mod_mult_o[386]) );
  XOR U5484 ( .A(n5481), .B(n5482), .Z(n3081) );
  IV U5485 ( .A(n3084), .Z(mod_mult_o[385]) );
  XOR U5486 ( .A(n5483), .B(n5484), .Z(n3084) );
  IV U5487 ( .A(n3087), .Z(mod_mult_o[384]) );
  XOR U5488 ( .A(n5485), .B(n5486), .Z(n3087) );
  IV U5489 ( .A(n3090), .Z(mod_mult_o[383]) );
  XOR U5490 ( .A(n5487), .B(n5488), .Z(n3090) );
  IV U5491 ( .A(n3093), .Z(mod_mult_o[382]) );
  XOR U5492 ( .A(n5489), .B(n5490), .Z(n3093) );
  IV U5493 ( .A(n3096), .Z(mod_mult_o[381]) );
  XOR U5494 ( .A(n5491), .B(n5492), .Z(n3096) );
  IV U5495 ( .A(n3099), .Z(mod_mult_o[380]) );
  XOR U5496 ( .A(n5493), .B(n5494), .Z(n3099) );
  IV U5497 ( .A(n3102), .Z(mod_mult_o[37]) );
  XOR U5498 ( .A(n5495), .B(n5496), .Z(n3102) );
  IV U5499 ( .A(n3105), .Z(mod_mult_o[379]) );
  XOR U5500 ( .A(n5497), .B(n5498), .Z(n3105) );
  IV U5501 ( .A(n3108), .Z(mod_mult_o[378]) );
  XOR U5502 ( .A(n5499), .B(n5500), .Z(n3108) );
  IV U5503 ( .A(n3111), .Z(mod_mult_o[377]) );
  XOR U5504 ( .A(n5501), .B(n5502), .Z(n3111) );
  IV U5505 ( .A(n3114), .Z(mod_mult_o[376]) );
  XOR U5506 ( .A(n5503), .B(n5504), .Z(n3114) );
  IV U5507 ( .A(n3117), .Z(mod_mult_o[375]) );
  XOR U5508 ( .A(n5505), .B(n5506), .Z(n3117) );
  IV U5509 ( .A(n3120), .Z(mod_mult_o[374]) );
  XOR U5510 ( .A(n5507), .B(n5508), .Z(n3120) );
  IV U5511 ( .A(n3123), .Z(mod_mult_o[373]) );
  XOR U5512 ( .A(n5509), .B(n5510), .Z(n3123) );
  IV U5513 ( .A(n3126), .Z(mod_mult_o[372]) );
  XOR U5514 ( .A(n5511), .B(n5512), .Z(n3126) );
  IV U5515 ( .A(n3129), .Z(mod_mult_o[371]) );
  XOR U5516 ( .A(n5513), .B(n5514), .Z(n3129) );
  IV U5517 ( .A(n3132), .Z(mod_mult_o[370]) );
  XOR U5518 ( .A(n5515), .B(n5516), .Z(n3132) );
  IV U5519 ( .A(n3135), .Z(mod_mult_o[36]) );
  XOR U5520 ( .A(n5517), .B(n5518), .Z(n3135) );
  IV U5521 ( .A(n3138), .Z(mod_mult_o[369]) );
  XOR U5522 ( .A(n5519), .B(n5520), .Z(n3138) );
  IV U5523 ( .A(n3141), .Z(mod_mult_o[368]) );
  XOR U5524 ( .A(n5521), .B(n5522), .Z(n3141) );
  IV U5525 ( .A(n3144), .Z(mod_mult_o[367]) );
  XOR U5526 ( .A(n5523), .B(n5524), .Z(n3144) );
  IV U5527 ( .A(n3147), .Z(mod_mult_o[366]) );
  XOR U5528 ( .A(n5525), .B(n5526), .Z(n3147) );
  IV U5529 ( .A(n3150), .Z(mod_mult_o[365]) );
  XOR U5530 ( .A(n5527), .B(n5528), .Z(n3150) );
  IV U5531 ( .A(n3153), .Z(mod_mult_o[364]) );
  XOR U5532 ( .A(n5529), .B(n5530), .Z(n3153) );
  IV U5533 ( .A(n3156), .Z(mod_mult_o[363]) );
  XOR U5534 ( .A(n5531), .B(n5532), .Z(n3156) );
  IV U5535 ( .A(n3159), .Z(mod_mult_o[362]) );
  XOR U5536 ( .A(n5533), .B(n5534), .Z(n3159) );
  IV U5537 ( .A(n3162), .Z(mod_mult_o[361]) );
  XOR U5538 ( .A(n5535), .B(n5536), .Z(n3162) );
  IV U5539 ( .A(n3165), .Z(mod_mult_o[360]) );
  XOR U5540 ( .A(n5537), .B(n5538), .Z(n3165) );
  IV U5541 ( .A(n3168), .Z(mod_mult_o[35]) );
  XOR U5542 ( .A(n5539), .B(n5540), .Z(n3168) );
  IV U5543 ( .A(n3171), .Z(mod_mult_o[359]) );
  XOR U5544 ( .A(n5541), .B(n5542), .Z(n3171) );
  IV U5545 ( .A(n3174), .Z(mod_mult_o[358]) );
  XOR U5546 ( .A(n5543), .B(n5544), .Z(n3174) );
  IV U5547 ( .A(n3177), .Z(mod_mult_o[357]) );
  XOR U5548 ( .A(n5545), .B(n5546), .Z(n3177) );
  IV U5549 ( .A(n3180), .Z(mod_mult_o[356]) );
  XOR U5550 ( .A(n5547), .B(n5548), .Z(n3180) );
  IV U5551 ( .A(n3183), .Z(mod_mult_o[355]) );
  XOR U5552 ( .A(n5549), .B(n5550), .Z(n3183) );
  IV U5553 ( .A(n3186), .Z(mod_mult_o[354]) );
  XOR U5554 ( .A(n5551), .B(n5552), .Z(n3186) );
  IV U5555 ( .A(n3189), .Z(mod_mult_o[353]) );
  XOR U5556 ( .A(n5553), .B(n5554), .Z(n3189) );
  IV U5557 ( .A(n3192), .Z(mod_mult_o[352]) );
  XOR U5558 ( .A(n5555), .B(n5556), .Z(n3192) );
  IV U5559 ( .A(n3195), .Z(mod_mult_o[351]) );
  XOR U5560 ( .A(n5557), .B(n5558), .Z(n3195) );
  IV U5561 ( .A(n3198), .Z(mod_mult_o[350]) );
  XOR U5562 ( .A(n5559), .B(n5560), .Z(n3198) );
  IV U5563 ( .A(n3201), .Z(mod_mult_o[34]) );
  XOR U5564 ( .A(n5561), .B(n5562), .Z(n3201) );
  IV U5565 ( .A(n3204), .Z(mod_mult_o[349]) );
  XOR U5566 ( .A(n5563), .B(n5564), .Z(n3204) );
  IV U5567 ( .A(n3207), .Z(mod_mult_o[348]) );
  XOR U5568 ( .A(n5565), .B(n5566), .Z(n3207) );
  IV U5569 ( .A(n3210), .Z(mod_mult_o[347]) );
  XOR U5570 ( .A(n5567), .B(n5568), .Z(n3210) );
  IV U5571 ( .A(n3213), .Z(mod_mult_o[346]) );
  XOR U5572 ( .A(n5569), .B(n5570), .Z(n3213) );
  IV U5573 ( .A(n3216), .Z(mod_mult_o[345]) );
  XOR U5574 ( .A(n5571), .B(n5572), .Z(n3216) );
  IV U5575 ( .A(n3219), .Z(mod_mult_o[344]) );
  XOR U5576 ( .A(n5573), .B(n5574), .Z(n3219) );
  IV U5577 ( .A(n3222), .Z(mod_mult_o[343]) );
  XOR U5578 ( .A(n5575), .B(n5576), .Z(n3222) );
  IV U5579 ( .A(n3225), .Z(mod_mult_o[342]) );
  XOR U5580 ( .A(n5577), .B(n5578), .Z(n3225) );
  IV U5581 ( .A(n3228), .Z(mod_mult_o[341]) );
  XOR U5582 ( .A(n5579), .B(n5580), .Z(n3228) );
  IV U5583 ( .A(n3231), .Z(mod_mult_o[340]) );
  XOR U5584 ( .A(n5581), .B(n5582), .Z(n3231) );
  IV U5585 ( .A(n3234), .Z(mod_mult_o[33]) );
  XOR U5586 ( .A(n5583), .B(n5584), .Z(n3234) );
  IV U5587 ( .A(n3237), .Z(mod_mult_o[339]) );
  XOR U5588 ( .A(n5585), .B(n5586), .Z(n3237) );
  IV U5589 ( .A(n3240), .Z(mod_mult_o[338]) );
  XOR U5590 ( .A(n5587), .B(n5588), .Z(n3240) );
  IV U5591 ( .A(n3243), .Z(mod_mult_o[337]) );
  XOR U5592 ( .A(n5589), .B(n5590), .Z(n3243) );
  IV U5593 ( .A(n3246), .Z(mod_mult_o[336]) );
  XOR U5594 ( .A(n5591), .B(n5592), .Z(n3246) );
  IV U5595 ( .A(n3249), .Z(mod_mult_o[335]) );
  XOR U5596 ( .A(n5593), .B(n5594), .Z(n3249) );
  IV U5597 ( .A(n3252), .Z(mod_mult_o[334]) );
  XOR U5598 ( .A(n5595), .B(n5596), .Z(n3252) );
  IV U5599 ( .A(n3255), .Z(mod_mult_o[333]) );
  XOR U5600 ( .A(n5597), .B(n5598), .Z(n3255) );
  IV U5601 ( .A(n3258), .Z(mod_mult_o[332]) );
  XOR U5602 ( .A(n5599), .B(n5600), .Z(n3258) );
  IV U5603 ( .A(n3261), .Z(mod_mult_o[331]) );
  XOR U5604 ( .A(n5601), .B(n5602), .Z(n3261) );
  IV U5605 ( .A(n3264), .Z(mod_mult_o[330]) );
  XOR U5606 ( .A(n5603), .B(n5604), .Z(n3264) );
  IV U5607 ( .A(n3267), .Z(mod_mult_o[32]) );
  XOR U5608 ( .A(n5605), .B(n5606), .Z(n3267) );
  IV U5609 ( .A(n3270), .Z(mod_mult_o[329]) );
  XOR U5610 ( .A(n5607), .B(n5608), .Z(n3270) );
  IV U5611 ( .A(n3273), .Z(mod_mult_o[328]) );
  XOR U5612 ( .A(n5609), .B(n5610), .Z(n3273) );
  IV U5613 ( .A(n3276), .Z(mod_mult_o[327]) );
  XOR U5614 ( .A(n5611), .B(n5612), .Z(n3276) );
  IV U5615 ( .A(n3279), .Z(mod_mult_o[326]) );
  XOR U5616 ( .A(n5613), .B(n5614), .Z(n3279) );
  IV U5617 ( .A(n3282), .Z(mod_mult_o[325]) );
  XOR U5618 ( .A(n5615), .B(n5616), .Z(n3282) );
  IV U5619 ( .A(n3285), .Z(mod_mult_o[324]) );
  XOR U5620 ( .A(n5617), .B(n5618), .Z(n3285) );
  IV U5621 ( .A(n3288), .Z(mod_mult_o[323]) );
  XOR U5622 ( .A(n5619), .B(n5620), .Z(n3288) );
  IV U5623 ( .A(n3291), .Z(mod_mult_o[322]) );
  XOR U5624 ( .A(n5621), .B(n5622), .Z(n3291) );
  IV U5625 ( .A(n3294), .Z(mod_mult_o[321]) );
  XOR U5626 ( .A(n5623), .B(n5624), .Z(n3294) );
  IV U5627 ( .A(n3297), .Z(mod_mult_o[320]) );
  XOR U5628 ( .A(n5625), .B(n5626), .Z(n3297) );
  IV U5629 ( .A(n3300), .Z(mod_mult_o[31]) );
  XOR U5630 ( .A(n5627), .B(n5628), .Z(n3300) );
  IV U5631 ( .A(n3303), .Z(mod_mult_o[319]) );
  XOR U5632 ( .A(n5629), .B(n5630), .Z(n3303) );
  IV U5633 ( .A(n3306), .Z(mod_mult_o[318]) );
  XOR U5634 ( .A(n5631), .B(n5632), .Z(n3306) );
  IV U5635 ( .A(n3309), .Z(mod_mult_o[317]) );
  XOR U5636 ( .A(n5633), .B(n5634), .Z(n3309) );
  IV U5637 ( .A(n3312), .Z(mod_mult_o[316]) );
  XOR U5638 ( .A(n5635), .B(n5636), .Z(n3312) );
  IV U5639 ( .A(n3315), .Z(mod_mult_o[315]) );
  XOR U5640 ( .A(n5637), .B(n5638), .Z(n3315) );
  IV U5641 ( .A(n3318), .Z(mod_mult_o[314]) );
  XOR U5642 ( .A(n5639), .B(n5640), .Z(n3318) );
  IV U5643 ( .A(n3321), .Z(mod_mult_o[313]) );
  XOR U5644 ( .A(n5641), .B(n5642), .Z(n3321) );
  IV U5645 ( .A(n3324), .Z(mod_mult_o[312]) );
  XOR U5646 ( .A(n5643), .B(n5644), .Z(n3324) );
  IV U5647 ( .A(n3327), .Z(mod_mult_o[311]) );
  XOR U5648 ( .A(n5645), .B(n5646), .Z(n3327) );
  IV U5649 ( .A(n3330), .Z(mod_mult_o[310]) );
  XOR U5650 ( .A(n5647), .B(n5648), .Z(n3330) );
  IV U5651 ( .A(n3333), .Z(mod_mult_o[30]) );
  XOR U5652 ( .A(n5649), .B(n5650), .Z(n3333) );
  IV U5653 ( .A(n3336), .Z(mod_mult_o[309]) );
  XOR U5654 ( .A(n5651), .B(n5652), .Z(n3336) );
  IV U5655 ( .A(n3339), .Z(mod_mult_o[308]) );
  XOR U5656 ( .A(n5653), .B(n5654), .Z(n3339) );
  IV U5657 ( .A(n3342), .Z(mod_mult_o[307]) );
  XOR U5658 ( .A(n5655), .B(n5656), .Z(n3342) );
  IV U5659 ( .A(n3345), .Z(mod_mult_o[306]) );
  XOR U5660 ( .A(n5657), .B(n5658), .Z(n3345) );
  IV U5661 ( .A(n3348), .Z(mod_mult_o[305]) );
  XOR U5662 ( .A(n5659), .B(n5660), .Z(n3348) );
  IV U5663 ( .A(n3351), .Z(mod_mult_o[304]) );
  XOR U5664 ( .A(n5661), .B(n5662), .Z(n3351) );
  IV U5665 ( .A(n3354), .Z(mod_mult_o[303]) );
  XOR U5666 ( .A(n5663), .B(n5664), .Z(n3354) );
  IV U5667 ( .A(n3357), .Z(mod_mult_o[302]) );
  XOR U5668 ( .A(n5665), .B(n5666), .Z(n3357) );
  IV U5669 ( .A(n3360), .Z(mod_mult_o[301]) );
  XOR U5670 ( .A(n5667), .B(n5668), .Z(n3360) );
  IV U5671 ( .A(n3363), .Z(mod_mult_o[300]) );
  XOR U5672 ( .A(n5669), .B(n5670), .Z(n3363) );
  IV U5673 ( .A(n3366), .Z(mod_mult_o[2]) );
  XOR U5674 ( .A(n5671), .B(n5672), .Z(n3366) );
  IV U5675 ( .A(n3369), .Z(mod_mult_o[29]) );
  XOR U5676 ( .A(n5673), .B(n5674), .Z(n3369) );
  IV U5677 ( .A(n3372), .Z(mod_mult_o[299]) );
  XOR U5678 ( .A(n5675), .B(n5676), .Z(n3372) );
  IV U5679 ( .A(n3375), .Z(mod_mult_o[298]) );
  XOR U5680 ( .A(n5677), .B(n5678), .Z(n3375) );
  IV U5681 ( .A(n3378), .Z(mod_mult_o[297]) );
  XOR U5682 ( .A(n5679), .B(n5680), .Z(n3378) );
  IV U5683 ( .A(n3381), .Z(mod_mult_o[296]) );
  XOR U5684 ( .A(n5681), .B(n5682), .Z(n3381) );
  IV U5685 ( .A(n3384), .Z(mod_mult_o[295]) );
  XOR U5686 ( .A(n5683), .B(n5684), .Z(n3384) );
  IV U5687 ( .A(n3387), .Z(mod_mult_o[294]) );
  XOR U5688 ( .A(n5685), .B(n5686), .Z(n3387) );
  IV U5689 ( .A(n3390), .Z(mod_mult_o[293]) );
  XOR U5690 ( .A(n5687), .B(n5688), .Z(n3390) );
  IV U5691 ( .A(n3393), .Z(mod_mult_o[292]) );
  XOR U5692 ( .A(n5689), .B(n5690), .Z(n3393) );
  IV U5693 ( .A(n3396), .Z(mod_mult_o[291]) );
  XOR U5694 ( .A(n5691), .B(n5692), .Z(n3396) );
  IV U5695 ( .A(n3399), .Z(mod_mult_o[290]) );
  XOR U5696 ( .A(n5693), .B(n5694), .Z(n3399) );
  IV U5697 ( .A(n3402), .Z(mod_mult_o[28]) );
  XOR U5698 ( .A(n5695), .B(n5696), .Z(n3402) );
  IV U5699 ( .A(n3405), .Z(mod_mult_o[289]) );
  XOR U5700 ( .A(n5697), .B(n5698), .Z(n3405) );
  IV U5701 ( .A(n3408), .Z(mod_mult_o[288]) );
  XOR U5702 ( .A(n5699), .B(n5700), .Z(n3408) );
  IV U5703 ( .A(n3411), .Z(mod_mult_o[287]) );
  XOR U5704 ( .A(n5701), .B(n5702), .Z(n3411) );
  IV U5705 ( .A(n3414), .Z(mod_mult_o[286]) );
  XOR U5706 ( .A(n5703), .B(n5704), .Z(n3414) );
  IV U5707 ( .A(n3417), .Z(mod_mult_o[285]) );
  XOR U5708 ( .A(n5705), .B(n5706), .Z(n3417) );
  IV U5709 ( .A(n3420), .Z(mod_mult_o[284]) );
  XOR U5710 ( .A(n5707), .B(n5708), .Z(n3420) );
  IV U5711 ( .A(n3423), .Z(mod_mult_o[283]) );
  XOR U5712 ( .A(n5709), .B(n5710), .Z(n3423) );
  IV U5713 ( .A(n3426), .Z(mod_mult_o[282]) );
  XOR U5714 ( .A(n5711), .B(n5712), .Z(n3426) );
  IV U5715 ( .A(n3429), .Z(mod_mult_o[281]) );
  XOR U5716 ( .A(n5713), .B(n5714), .Z(n3429) );
  IV U5717 ( .A(n3432), .Z(mod_mult_o[280]) );
  XOR U5718 ( .A(n5715), .B(n5716), .Z(n3432) );
  IV U5719 ( .A(n3435), .Z(mod_mult_o[27]) );
  XOR U5720 ( .A(n5717), .B(n5718), .Z(n3435) );
  IV U5721 ( .A(n3438), .Z(mod_mult_o[279]) );
  XOR U5722 ( .A(n5719), .B(n5720), .Z(n3438) );
  IV U5723 ( .A(n3441), .Z(mod_mult_o[278]) );
  XOR U5724 ( .A(n5721), .B(n5722), .Z(n3441) );
  IV U5725 ( .A(n3444), .Z(mod_mult_o[277]) );
  XOR U5726 ( .A(n5723), .B(n5724), .Z(n3444) );
  IV U5727 ( .A(n3447), .Z(mod_mult_o[276]) );
  XOR U5728 ( .A(n5725), .B(n5726), .Z(n3447) );
  IV U5729 ( .A(n3450), .Z(mod_mult_o[275]) );
  XOR U5730 ( .A(n5727), .B(n5728), .Z(n3450) );
  IV U5731 ( .A(n3453), .Z(mod_mult_o[274]) );
  XOR U5732 ( .A(n5729), .B(n5730), .Z(n3453) );
  IV U5733 ( .A(n3456), .Z(mod_mult_o[273]) );
  XOR U5734 ( .A(n5731), .B(n5732), .Z(n3456) );
  IV U5735 ( .A(n3459), .Z(mod_mult_o[272]) );
  XOR U5736 ( .A(n5733), .B(n5734), .Z(n3459) );
  IV U5737 ( .A(n3462), .Z(mod_mult_o[271]) );
  XOR U5738 ( .A(n5735), .B(n5736), .Z(n3462) );
  IV U5739 ( .A(n3465), .Z(mod_mult_o[270]) );
  XOR U5740 ( .A(n5737), .B(n5738), .Z(n3465) );
  IV U5741 ( .A(n3468), .Z(mod_mult_o[26]) );
  XOR U5742 ( .A(n5739), .B(n5740), .Z(n3468) );
  IV U5743 ( .A(n3471), .Z(mod_mult_o[269]) );
  XOR U5744 ( .A(n5741), .B(n5742), .Z(n3471) );
  IV U5745 ( .A(n3474), .Z(mod_mult_o[268]) );
  XOR U5746 ( .A(n5743), .B(n5744), .Z(n3474) );
  IV U5747 ( .A(n3477), .Z(mod_mult_o[267]) );
  XOR U5748 ( .A(n5745), .B(n5746), .Z(n3477) );
  IV U5749 ( .A(n3480), .Z(mod_mult_o[266]) );
  XOR U5750 ( .A(n5747), .B(n5748), .Z(n3480) );
  IV U5751 ( .A(n3483), .Z(mod_mult_o[265]) );
  XOR U5752 ( .A(n5749), .B(n5750), .Z(n3483) );
  IV U5753 ( .A(n3486), .Z(mod_mult_o[264]) );
  XOR U5754 ( .A(n5751), .B(n5752), .Z(n3486) );
  IV U5755 ( .A(n3489), .Z(mod_mult_o[263]) );
  XOR U5756 ( .A(n5753), .B(n5754), .Z(n3489) );
  IV U5757 ( .A(n3492), .Z(mod_mult_o[262]) );
  XOR U5758 ( .A(n5755), .B(n5756), .Z(n3492) );
  IV U5759 ( .A(n3495), .Z(mod_mult_o[261]) );
  XOR U5760 ( .A(n5757), .B(n5758), .Z(n3495) );
  IV U5761 ( .A(n3498), .Z(mod_mult_o[260]) );
  XOR U5762 ( .A(n5759), .B(n5760), .Z(n3498) );
  IV U5763 ( .A(n3501), .Z(mod_mult_o[25]) );
  XOR U5764 ( .A(n5761), .B(n5762), .Z(n3501) );
  IV U5765 ( .A(n3504), .Z(mod_mult_o[259]) );
  XOR U5766 ( .A(n5763), .B(n5764), .Z(n3504) );
  IV U5767 ( .A(n3507), .Z(mod_mult_o[258]) );
  XOR U5768 ( .A(n5765), .B(n5766), .Z(n3507) );
  IV U5769 ( .A(n3510), .Z(mod_mult_o[257]) );
  XOR U5770 ( .A(n5767), .B(n5768), .Z(n3510) );
  IV U5771 ( .A(n3513), .Z(mod_mult_o[256]) );
  XOR U5772 ( .A(n5769), .B(n5770), .Z(n3513) );
  IV U5773 ( .A(n3516), .Z(mod_mult_o[255]) );
  XOR U5774 ( .A(n5771), .B(n5772), .Z(n3516) );
  IV U5775 ( .A(n3519), .Z(mod_mult_o[254]) );
  XOR U5776 ( .A(n5773), .B(n5774), .Z(n3519) );
  IV U5777 ( .A(n3522), .Z(mod_mult_o[253]) );
  XOR U5778 ( .A(n5775), .B(n5776), .Z(n3522) );
  IV U5779 ( .A(n3525), .Z(mod_mult_o[252]) );
  XOR U5780 ( .A(n5777), .B(n5778), .Z(n3525) );
  IV U5781 ( .A(n3528), .Z(mod_mult_o[251]) );
  XOR U5782 ( .A(n5779), .B(n5780), .Z(n3528) );
  IV U5783 ( .A(n3531), .Z(mod_mult_o[250]) );
  XOR U5784 ( .A(n5781), .B(n5782), .Z(n3531) );
  IV U5785 ( .A(n3534), .Z(mod_mult_o[24]) );
  XOR U5786 ( .A(n5783), .B(n5784), .Z(n3534) );
  IV U5787 ( .A(n3537), .Z(mod_mult_o[249]) );
  XOR U5788 ( .A(n5785), .B(n5786), .Z(n3537) );
  IV U5789 ( .A(n3540), .Z(mod_mult_o[248]) );
  XOR U5790 ( .A(n5787), .B(n5788), .Z(n3540) );
  IV U5791 ( .A(n3543), .Z(mod_mult_o[247]) );
  XOR U5792 ( .A(n5789), .B(n5790), .Z(n3543) );
  IV U5793 ( .A(n3546), .Z(mod_mult_o[246]) );
  XOR U5794 ( .A(n5791), .B(n5792), .Z(n3546) );
  IV U5795 ( .A(n3549), .Z(mod_mult_o[245]) );
  XOR U5796 ( .A(n5793), .B(n5794), .Z(n3549) );
  IV U5797 ( .A(n3552), .Z(mod_mult_o[244]) );
  XOR U5798 ( .A(n5795), .B(n5796), .Z(n3552) );
  IV U5799 ( .A(n3555), .Z(mod_mult_o[243]) );
  XOR U5800 ( .A(n5797), .B(n5798), .Z(n3555) );
  IV U5801 ( .A(n3558), .Z(mod_mult_o[242]) );
  XOR U5802 ( .A(n5799), .B(n5800), .Z(n3558) );
  IV U5803 ( .A(n3561), .Z(mod_mult_o[241]) );
  XOR U5804 ( .A(n5801), .B(n5802), .Z(n3561) );
  IV U5805 ( .A(n3564), .Z(mod_mult_o[240]) );
  XOR U5806 ( .A(n5803), .B(n5804), .Z(n3564) );
  IV U5807 ( .A(n3567), .Z(mod_mult_o[23]) );
  XOR U5808 ( .A(n5805), .B(n5806), .Z(n3567) );
  IV U5809 ( .A(n3570), .Z(mod_mult_o[239]) );
  XOR U5810 ( .A(n5807), .B(n5808), .Z(n3570) );
  IV U5811 ( .A(n3573), .Z(mod_mult_o[238]) );
  XOR U5812 ( .A(n5809), .B(n5810), .Z(n3573) );
  IV U5813 ( .A(n3576), .Z(mod_mult_o[237]) );
  XOR U5814 ( .A(n5811), .B(n5812), .Z(n3576) );
  IV U5815 ( .A(n3579), .Z(mod_mult_o[236]) );
  XOR U5816 ( .A(n5813), .B(n5814), .Z(n3579) );
  IV U5817 ( .A(n3582), .Z(mod_mult_o[235]) );
  XOR U5818 ( .A(n5815), .B(n5816), .Z(n3582) );
  IV U5819 ( .A(n3585), .Z(mod_mult_o[234]) );
  XOR U5820 ( .A(n5817), .B(n5818), .Z(n3585) );
  IV U5821 ( .A(n3588), .Z(mod_mult_o[233]) );
  XOR U5822 ( .A(n5819), .B(n5820), .Z(n3588) );
  IV U5823 ( .A(n3591), .Z(mod_mult_o[232]) );
  XOR U5824 ( .A(n5821), .B(n5822), .Z(n3591) );
  IV U5825 ( .A(n3594), .Z(mod_mult_o[231]) );
  XOR U5826 ( .A(n5823), .B(n5824), .Z(n3594) );
  IV U5827 ( .A(n3597), .Z(mod_mult_o[230]) );
  XOR U5828 ( .A(n5825), .B(n5826), .Z(n3597) );
  IV U5829 ( .A(n3600), .Z(mod_mult_o[22]) );
  XOR U5830 ( .A(n5827), .B(n5828), .Z(n3600) );
  IV U5831 ( .A(n3603), .Z(mod_mult_o[229]) );
  XOR U5832 ( .A(n5829), .B(n5830), .Z(n3603) );
  IV U5833 ( .A(n3606), .Z(mod_mult_o[228]) );
  XOR U5834 ( .A(n5831), .B(n5832), .Z(n3606) );
  IV U5835 ( .A(n3609), .Z(mod_mult_o[227]) );
  XOR U5836 ( .A(n5833), .B(n5834), .Z(n3609) );
  IV U5837 ( .A(n3612), .Z(mod_mult_o[226]) );
  XOR U5838 ( .A(n5835), .B(n5836), .Z(n3612) );
  IV U5839 ( .A(n3615), .Z(mod_mult_o[225]) );
  XOR U5840 ( .A(n5837), .B(n5838), .Z(n3615) );
  IV U5841 ( .A(n3618), .Z(mod_mult_o[224]) );
  XOR U5842 ( .A(n5839), .B(n5840), .Z(n3618) );
  IV U5843 ( .A(n3621), .Z(mod_mult_o[223]) );
  XOR U5844 ( .A(n5841), .B(n5842), .Z(n3621) );
  IV U5845 ( .A(n3624), .Z(mod_mult_o[222]) );
  XOR U5846 ( .A(n5843), .B(n5844), .Z(n3624) );
  IV U5847 ( .A(n3627), .Z(mod_mult_o[221]) );
  XOR U5848 ( .A(n5845), .B(n5846), .Z(n3627) );
  IV U5849 ( .A(n3630), .Z(mod_mult_o[220]) );
  XOR U5850 ( .A(n5847), .B(n5848), .Z(n3630) );
  IV U5851 ( .A(n3633), .Z(mod_mult_o[21]) );
  XOR U5852 ( .A(n5849), .B(n5850), .Z(n3633) );
  IV U5853 ( .A(n3636), .Z(mod_mult_o[219]) );
  XOR U5854 ( .A(n5851), .B(n5852), .Z(n3636) );
  IV U5855 ( .A(n3639), .Z(mod_mult_o[218]) );
  XOR U5856 ( .A(n5853), .B(n5854), .Z(n3639) );
  IV U5857 ( .A(n3642), .Z(mod_mult_o[217]) );
  XOR U5858 ( .A(n5855), .B(n5856), .Z(n3642) );
  IV U5859 ( .A(n3645), .Z(mod_mult_o[216]) );
  XOR U5860 ( .A(n5857), .B(n5858), .Z(n3645) );
  IV U5861 ( .A(n3648), .Z(mod_mult_o[215]) );
  XOR U5862 ( .A(n5859), .B(n5860), .Z(n3648) );
  IV U5863 ( .A(n3651), .Z(mod_mult_o[214]) );
  XOR U5864 ( .A(n5861), .B(n5862), .Z(n3651) );
  IV U5865 ( .A(n3654), .Z(mod_mult_o[213]) );
  XOR U5866 ( .A(n5863), .B(n5864), .Z(n3654) );
  IV U5867 ( .A(n3657), .Z(mod_mult_o[212]) );
  XOR U5868 ( .A(n5865), .B(n5866), .Z(n3657) );
  IV U5869 ( .A(n3660), .Z(mod_mult_o[211]) );
  XOR U5870 ( .A(n5867), .B(n5868), .Z(n3660) );
  IV U5871 ( .A(n3663), .Z(mod_mult_o[210]) );
  XOR U5872 ( .A(n5869), .B(n5870), .Z(n3663) );
  IV U5873 ( .A(n3666), .Z(mod_mult_o[20]) );
  XOR U5874 ( .A(n5871), .B(n5872), .Z(n3666) );
  IV U5875 ( .A(n3669), .Z(mod_mult_o[209]) );
  XOR U5876 ( .A(n5873), .B(n5874), .Z(n3669) );
  IV U5877 ( .A(n3672), .Z(mod_mult_o[208]) );
  XOR U5878 ( .A(n5875), .B(n5876), .Z(n3672) );
  IV U5879 ( .A(n3675), .Z(mod_mult_o[207]) );
  XOR U5880 ( .A(n5877), .B(n5878), .Z(n3675) );
  IV U5881 ( .A(n3678), .Z(mod_mult_o[206]) );
  XOR U5882 ( .A(n5879), .B(n5880), .Z(n3678) );
  IV U5883 ( .A(n3681), .Z(mod_mult_o[205]) );
  XOR U5884 ( .A(n5881), .B(n5882), .Z(n3681) );
  IV U5885 ( .A(n3684), .Z(mod_mult_o[204]) );
  XOR U5886 ( .A(n5883), .B(n5884), .Z(n3684) );
  IV U5887 ( .A(n3687), .Z(mod_mult_o[203]) );
  XOR U5888 ( .A(n5885), .B(n5886), .Z(n3687) );
  IV U5889 ( .A(n3690), .Z(mod_mult_o[202]) );
  XOR U5890 ( .A(n5887), .B(n5888), .Z(n3690) );
  IV U5891 ( .A(n3693), .Z(mod_mult_o[201]) );
  XOR U5892 ( .A(n5889), .B(n5890), .Z(n3693) );
  IV U5893 ( .A(n3696), .Z(mod_mult_o[200]) );
  XOR U5894 ( .A(n5891), .B(n5892), .Z(n3696) );
  IV U5895 ( .A(n3699), .Z(mod_mult_o[1]) );
  XOR U5896 ( .A(n5893), .B(n5894), .Z(n3699) );
  IV U5897 ( .A(n3702), .Z(mod_mult_o[19]) );
  XOR U5898 ( .A(n5895), .B(n5896), .Z(n3702) );
  IV U5899 ( .A(n3705), .Z(mod_mult_o[199]) );
  XOR U5900 ( .A(n5897), .B(n5898), .Z(n3705) );
  IV U5901 ( .A(n3708), .Z(mod_mult_o[198]) );
  XOR U5902 ( .A(n5899), .B(n5900), .Z(n3708) );
  IV U5903 ( .A(n3711), .Z(mod_mult_o[197]) );
  XOR U5904 ( .A(n5901), .B(n5902), .Z(n3711) );
  IV U5905 ( .A(n3714), .Z(mod_mult_o[196]) );
  XOR U5906 ( .A(n5903), .B(n5904), .Z(n3714) );
  IV U5907 ( .A(n3717), .Z(mod_mult_o[195]) );
  XOR U5908 ( .A(n5905), .B(n5906), .Z(n3717) );
  IV U5909 ( .A(n3720), .Z(mod_mult_o[194]) );
  XOR U5910 ( .A(n5907), .B(n5908), .Z(n3720) );
  IV U5911 ( .A(n3723), .Z(mod_mult_o[193]) );
  XOR U5912 ( .A(n5909), .B(n5910), .Z(n3723) );
  IV U5913 ( .A(n3726), .Z(mod_mult_o[192]) );
  XOR U5914 ( .A(n5911), .B(n5912), .Z(n3726) );
  IV U5915 ( .A(n3729), .Z(mod_mult_o[191]) );
  XOR U5916 ( .A(n5913), .B(n5914), .Z(n3729) );
  IV U5917 ( .A(n3732), .Z(mod_mult_o[190]) );
  XOR U5918 ( .A(n5915), .B(n5916), .Z(n3732) );
  IV U5919 ( .A(n3735), .Z(mod_mult_o[18]) );
  XOR U5920 ( .A(n5917), .B(n5918), .Z(n3735) );
  IV U5921 ( .A(n3738), .Z(mod_mult_o[189]) );
  XOR U5922 ( .A(n5919), .B(n5920), .Z(n3738) );
  IV U5923 ( .A(n3741), .Z(mod_mult_o[188]) );
  XOR U5924 ( .A(n5921), .B(n5922), .Z(n3741) );
  IV U5925 ( .A(n3744), .Z(mod_mult_o[187]) );
  XOR U5926 ( .A(n5923), .B(n5924), .Z(n3744) );
  IV U5927 ( .A(n3747), .Z(mod_mult_o[186]) );
  XOR U5928 ( .A(n5925), .B(n5926), .Z(n3747) );
  IV U5929 ( .A(n3750), .Z(mod_mult_o[185]) );
  XOR U5930 ( .A(n5927), .B(n5928), .Z(n3750) );
  IV U5931 ( .A(n3753), .Z(mod_mult_o[184]) );
  XOR U5932 ( .A(n5929), .B(n5930), .Z(n3753) );
  IV U5933 ( .A(n3756), .Z(mod_mult_o[183]) );
  XOR U5934 ( .A(n5931), .B(n5932), .Z(n3756) );
  IV U5935 ( .A(n3759), .Z(mod_mult_o[182]) );
  XOR U5936 ( .A(n5933), .B(n5934), .Z(n3759) );
  IV U5937 ( .A(n3762), .Z(mod_mult_o[181]) );
  XOR U5938 ( .A(n5935), .B(n5936), .Z(n3762) );
  IV U5939 ( .A(n3765), .Z(mod_mult_o[180]) );
  XOR U5940 ( .A(n5937), .B(n5938), .Z(n3765) );
  IV U5941 ( .A(n3768), .Z(mod_mult_o[17]) );
  XOR U5942 ( .A(n5939), .B(n5940), .Z(n3768) );
  IV U5943 ( .A(n3771), .Z(mod_mult_o[179]) );
  XOR U5944 ( .A(n5941), .B(n5942), .Z(n3771) );
  IV U5945 ( .A(n3774), .Z(mod_mult_o[178]) );
  XOR U5946 ( .A(n5943), .B(n5944), .Z(n3774) );
  IV U5947 ( .A(n3777), .Z(mod_mult_o[177]) );
  XOR U5948 ( .A(n5945), .B(n5946), .Z(n3777) );
  IV U5949 ( .A(n3780), .Z(mod_mult_o[176]) );
  XOR U5950 ( .A(n5947), .B(n5948), .Z(n3780) );
  IV U5951 ( .A(n3783), .Z(mod_mult_o[175]) );
  XOR U5952 ( .A(n5949), .B(n5950), .Z(n3783) );
  IV U5953 ( .A(n3786), .Z(mod_mult_o[174]) );
  XOR U5954 ( .A(n5951), .B(n5952), .Z(n3786) );
  IV U5955 ( .A(n3789), .Z(mod_mult_o[173]) );
  XOR U5956 ( .A(n5953), .B(n5954), .Z(n3789) );
  IV U5957 ( .A(n3792), .Z(mod_mult_o[172]) );
  XOR U5958 ( .A(n5955), .B(n5956), .Z(n3792) );
  IV U5959 ( .A(n3795), .Z(mod_mult_o[171]) );
  XOR U5960 ( .A(n5957), .B(n5958), .Z(n3795) );
  IV U5961 ( .A(n3798), .Z(mod_mult_o[170]) );
  XOR U5962 ( .A(n5959), .B(n5960), .Z(n3798) );
  IV U5963 ( .A(n3801), .Z(mod_mult_o[16]) );
  XOR U5964 ( .A(n5961), .B(n5962), .Z(n3801) );
  IV U5965 ( .A(n3804), .Z(mod_mult_o[169]) );
  XOR U5966 ( .A(n5963), .B(n5964), .Z(n3804) );
  IV U5967 ( .A(n3807), .Z(mod_mult_o[168]) );
  XOR U5968 ( .A(n5965), .B(n5966), .Z(n3807) );
  IV U5969 ( .A(n3810), .Z(mod_mult_o[167]) );
  XOR U5970 ( .A(n5967), .B(n5968), .Z(n3810) );
  IV U5971 ( .A(n3813), .Z(mod_mult_o[166]) );
  XOR U5972 ( .A(n5969), .B(n5970), .Z(n3813) );
  IV U5973 ( .A(n3816), .Z(mod_mult_o[165]) );
  XOR U5974 ( .A(n5971), .B(n5972), .Z(n3816) );
  IV U5975 ( .A(n3819), .Z(mod_mult_o[164]) );
  XOR U5976 ( .A(n5973), .B(n5974), .Z(n3819) );
  IV U5977 ( .A(n3822), .Z(mod_mult_o[163]) );
  XOR U5978 ( .A(n5975), .B(n5976), .Z(n3822) );
  IV U5979 ( .A(n3825), .Z(mod_mult_o[162]) );
  XOR U5980 ( .A(n5977), .B(n5978), .Z(n3825) );
  IV U5981 ( .A(n3828), .Z(mod_mult_o[161]) );
  XOR U5982 ( .A(n5979), .B(n5980), .Z(n3828) );
  IV U5983 ( .A(n3831), .Z(mod_mult_o[160]) );
  XOR U5984 ( .A(n5981), .B(n5982), .Z(n3831) );
  IV U5985 ( .A(n3834), .Z(mod_mult_o[15]) );
  XOR U5986 ( .A(n5983), .B(n5984), .Z(n3834) );
  IV U5987 ( .A(n3837), .Z(mod_mult_o[159]) );
  XOR U5988 ( .A(n5985), .B(n5986), .Z(n3837) );
  IV U5989 ( .A(n3840), .Z(mod_mult_o[158]) );
  XOR U5990 ( .A(n5987), .B(n5988), .Z(n3840) );
  IV U5991 ( .A(n3843), .Z(mod_mult_o[157]) );
  XOR U5992 ( .A(n5989), .B(n5990), .Z(n3843) );
  IV U5993 ( .A(n3846), .Z(mod_mult_o[156]) );
  XOR U5994 ( .A(n5991), .B(n5992), .Z(n3846) );
  IV U5995 ( .A(n3849), .Z(mod_mult_o[155]) );
  XOR U5996 ( .A(n5993), .B(n5994), .Z(n3849) );
  IV U5997 ( .A(n3852), .Z(mod_mult_o[154]) );
  XOR U5998 ( .A(n5995), .B(n5996), .Z(n3852) );
  IV U5999 ( .A(n3855), .Z(mod_mult_o[153]) );
  XOR U6000 ( .A(n5997), .B(n5998), .Z(n3855) );
  IV U6001 ( .A(n3858), .Z(mod_mult_o[152]) );
  XOR U6002 ( .A(n5999), .B(n6000), .Z(n3858) );
  IV U6003 ( .A(n3861), .Z(mod_mult_o[151]) );
  XOR U6004 ( .A(n6001), .B(n6002), .Z(n3861) );
  IV U6005 ( .A(n3864), .Z(mod_mult_o[150]) );
  XOR U6006 ( .A(n6003), .B(n6004), .Z(n3864) );
  IV U6007 ( .A(n3867), .Z(mod_mult_o[14]) );
  XOR U6008 ( .A(n6005), .B(n6006), .Z(n3867) );
  IV U6009 ( .A(n3870), .Z(mod_mult_o[149]) );
  XOR U6010 ( .A(n6007), .B(n6008), .Z(n3870) );
  IV U6011 ( .A(n3873), .Z(mod_mult_o[148]) );
  XOR U6012 ( .A(n6009), .B(n6010), .Z(n3873) );
  IV U6013 ( .A(n3876), .Z(mod_mult_o[147]) );
  XOR U6014 ( .A(n6011), .B(n6012), .Z(n3876) );
  IV U6015 ( .A(n3879), .Z(mod_mult_o[146]) );
  XOR U6016 ( .A(n6013), .B(n6014), .Z(n3879) );
  IV U6017 ( .A(n3882), .Z(mod_mult_o[145]) );
  XOR U6018 ( .A(n6015), .B(n6016), .Z(n3882) );
  IV U6019 ( .A(n3885), .Z(mod_mult_o[144]) );
  XOR U6020 ( .A(n6017), .B(n6018), .Z(n3885) );
  IV U6021 ( .A(n3888), .Z(mod_mult_o[143]) );
  XOR U6022 ( .A(n6019), .B(n6020), .Z(n3888) );
  IV U6023 ( .A(n3891), .Z(mod_mult_o[142]) );
  XOR U6024 ( .A(n6021), .B(n6022), .Z(n3891) );
  IV U6025 ( .A(n3894), .Z(mod_mult_o[141]) );
  XOR U6026 ( .A(n6023), .B(n6024), .Z(n3894) );
  IV U6027 ( .A(n3897), .Z(mod_mult_o[140]) );
  XOR U6028 ( .A(n6025), .B(n6026), .Z(n3897) );
  IV U6029 ( .A(n3900), .Z(mod_mult_o[13]) );
  XOR U6030 ( .A(n6027), .B(n6028), .Z(n3900) );
  IV U6031 ( .A(n3903), .Z(mod_mult_o[139]) );
  XOR U6032 ( .A(n6029), .B(n6030), .Z(n3903) );
  IV U6033 ( .A(n3906), .Z(mod_mult_o[138]) );
  XOR U6034 ( .A(n6031), .B(n6032), .Z(n3906) );
  IV U6035 ( .A(n3909), .Z(mod_mult_o[137]) );
  XOR U6036 ( .A(n6033), .B(n6034), .Z(n3909) );
  IV U6037 ( .A(n3912), .Z(mod_mult_o[136]) );
  XOR U6038 ( .A(n6035), .B(n6036), .Z(n3912) );
  IV U6039 ( .A(n3915), .Z(mod_mult_o[135]) );
  XOR U6040 ( .A(n6037), .B(n6038), .Z(n3915) );
  IV U6041 ( .A(n3918), .Z(mod_mult_o[134]) );
  XOR U6042 ( .A(n6039), .B(n6040), .Z(n3918) );
  IV U6043 ( .A(n3921), .Z(mod_mult_o[133]) );
  XOR U6044 ( .A(n6041), .B(n6042), .Z(n3921) );
  IV U6045 ( .A(n3924), .Z(mod_mult_o[132]) );
  XOR U6046 ( .A(n6043), .B(n6044), .Z(n3924) );
  IV U6047 ( .A(n3927), .Z(mod_mult_o[131]) );
  XOR U6048 ( .A(n6045), .B(n6046), .Z(n3927) );
  IV U6049 ( .A(n3930), .Z(mod_mult_o[130]) );
  XOR U6050 ( .A(n6047), .B(n6048), .Z(n3930) );
  IV U6051 ( .A(n3933), .Z(mod_mult_o[12]) );
  XOR U6052 ( .A(n6049), .B(n6050), .Z(n3933) );
  IV U6053 ( .A(n3936), .Z(mod_mult_o[129]) );
  XOR U6054 ( .A(n6051), .B(n6052), .Z(n3936) );
  IV U6055 ( .A(n3939), .Z(mod_mult_o[128]) );
  XOR U6056 ( .A(n6053), .B(n6054), .Z(n3939) );
  IV U6057 ( .A(n3942), .Z(mod_mult_o[127]) );
  XOR U6058 ( .A(n6055), .B(n6056), .Z(n3942) );
  IV U6059 ( .A(n3945), .Z(mod_mult_o[126]) );
  XOR U6060 ( .A(n6057), .B(n6058), .Z(n3945) );
  IV U6061 ( .A(n3948), .Z(mod_mult_o[125]) );
  XOR U6062 ( .A(n6059), .B(n6060), .Z(n3948) );
  IV U6063 ( .A(n3951), .Z(mod_mult_o[124]) );
  XOR U6064 ( .A(n6061), .B(n6062), .Z(n3951) );
  IV U6065 ( .A(n3954), .Z(mod_mult_o[123]) );
  XOR U6066 ( .A(n6063), .B(n6064), .Z(n3954) );
  IV U6067 ( .A(n3957), .Z(mod_mult_o[122]) );
  XOR U6068 ( .A(n6065), .B(n6066), .Z(n3957) );
  IV U6069 ( .A(n3960), .Z(mod_mult_o[121]) );
  XOR U6070 ( .A(n6067), .B(n6068), .Z(n3960) );
  IV U6071 ( .A(n3963), .Z(mod_mult_o[120]) );
  XOR U6072 ( .A(n6069), .B(n6070), .Z(n3963) );
  IV U6073 ( .A(n3966), .Z(mod_mult_o[11]) );
  XOR U6074 ( .A(n6071), .B(n6072), .Z(n3966) );
  IV U6075 ( .A(n3969), .Z(mod_mult_o[119]) );
  XOR U6076 ( .A(n6073), .B(n6074), .Z(n3969) );
  IV U6077 ( .A(n3972), .Z(mod_mult_o[118]) );
  XOR U6078 ( .A(n6075), .B(n6076), .Z(n3972) );
  IV U6079 ( .A(n3975), .Z(mod_mult_o[117]) );
  XOR U6080 ( .A(n6077), .B(n6078), .Z(n3975) );
  IV U6081 ( .A(n3978), .Z(mod_mult_o[116]) );
  XOR U6082 ( .A(n6079), .B(n6080), .Z(n3978) );
  IV U6083 ( .A(n3981), .Z(mod_mult_o[115]) );
  XOR U6084 ( .A(n6081), .B(n6082), .Z(n3981) );
  IV U6085 ( .A(n3984), .Z(mod_mult_o[114]) );
  XOR U6086 ( .A(n6083), .B(n6084), .Z(n3984) );
  IV U6087 ( .A(n3987), .Z(mod_mult_o[113]) );
  XOR U6088 ( .A(n6085), .B(n6086), .Z(n3987) );
  IV U6089 ( .A(n3990), .Z(mod_mult_o[112]) );
  XOR U6090 ( .A(n6087), .B(n6088), .Z(n3990) );
  IV U6091 ( .A(n3993), .Z(mod_mult_o[111]) );
  XOR U6092 ( .A(n6089), .B(n6090), .Z(n3993) );
  IV U6093 ( .A(n3996), .Z(mod_mult_o[110]) );
  XOR U6094 ( .A(n6091), .B(n6092), .Z(n3996) );
  IV U6095 ( .A(n3999), .Z(mod_mult_o[10]) );
  XOR U6096 ( .A(n6093), .B(n6094), .Z(n3999) );
  IV U6097 ( .A(n4002), .Z(mod_mult_o[109]) );
  XOR U6098 ( .A(n6095), .B(n6096), .Z(n4002) );
  IV U6099 ( .A(n4005), .Z(mod_mult_o[108]) );
  XOR U6100 ( .A(n6097), .B(n6098), .Z(n4005) );
  IV U6101 ( .A(n4008), .Z(mod_mult_o[107]) );
  XOR U6102 ( .A(n6099), .B(n6100), .Z(n4008) );
  IV U6103 ( .A(n4011), .Z(mod_mult_o[106]) );
  XOR U6104 ( .A(n6101), .B(n6102), .Z(n4011) );
  IV U6105 ( .A(n4014), .Z(mod_mult_o[105]) );
  XOR U6106 ( .A(n6103), .B(n6104), .Z(n4014) );
  IV U6107 ( .A(n4017), .Z(mod_mult_o[104]) );
  XOR U6108 ( .A(n6105), .B(n6106), .Z(n4017) );
  IV U6109 ( .A(n4020), .Z(mod_mult_o[103]) );
  XOR U6110 ( .A(n6107), .B(n6108), .Z(n4020) );
  IV U6111 ( .A(n4023), .Z(mod_mult_o[102]) );
  XOR U6112 ( .A(n6109), .B(n6110), .Z(n4023) );
  IV U6113 ( .A(n4026), .Z(mod_mult_o[1023]) );
  XOR U6114 ( .A(n4114), .B(n4115), .Z(n4026) );
  NAND U6115 ( .A(n6111), .B(e_input[1023]), .Z(n4115) );
  NAND U6116 ( .A(n6112), .B(e_input[1023]), .Z(n6111) );
  XOR U6117 ( .A(n4109), .B(n6113), .Z(n4114) );
  IV U6118 ( .A(n4116), .Z(n4109) );
  XOR U6119 ( .A(n6114), .B(n6115), .Z(n4116) );
  ANDN U6120 ( .A(n6116), .B(n6117), .Z(n6115) );
  XNOR U6121 ( .A(n6118), .B(n6114), .Z(n6116) );
  IV U6122 ( .A(n4029), .Z(mod_mult_o[1022]) );
  XOR U6123 ( .A(n6117), .B(n6118), .Z(n4029) );
  NAND U6124 ( .A(n6119), .B(e_input[1022]), .Z(n6118) );
  NAND U6125 ( .A(n6112), .B(e_input[1022]), .Z(n6119) );
  XOR U6126 ( .A(n6120), .B(n6121), .Z(n6117) );
  IV U6127 ( .A(n6114), .Z(n6120) );
  XOR U6128 ( .A(n6122), .B(n6123), .Z(n6114) );
  ANDN U6129 ( .A(n6124), .B(n6125), .Z(n6123) );
  XNOR U6130 ( .A(n6126), .B(n6122), .Z(n6124) );
  IV U6131 ( .A(n4032), .Z(mod_mult_o[1021]) );
  XOR U6132 ( .A(n6125), .B(n6126), .Z(n4032) );
  NAND U6133 ( .A(n6127), .B(e_input[1021]), .Z(n6126) );
  NAND U6134 ( .A(n6112), .B(e_input[1021]), .Z(n6127) );
  XOR U6135 ( .A(n6128), .B(n6129), .Z(n6125) );
  IV U6136 ( .A(n6122), .Z(n6128) );
  XOR U6137 ( .A(n6130), .B(n6131), .Z(n6122) );
  ANDN U6138 ( .A(n6132), .B(n6133), .Z(n6131) );
  XNOR U6139 ( .A(n6134), .B(n6130), .Z(n6132) );
  IV U6140 ( .A(n4035), .Z(mod_mult_o[1020]) );
  XOR U6141 ( .A(n6133), .B(n6134), .Z(n4035) );
  NAND U6142 ( .A(n6135), .B(e_input[1020]), .Z(n6134) );
  NAND U6143 ( .A(n6112), .B(e_input[1020]), .Z(n6135) );
  XOR U6144 ( .A(n6136), .B(n6137), .Z(n6133) );
  IV U6145 ( .A(n6130), .Z(n6136) );
  XOR U6146 ( .A(n6138), .B(n6139), .Z(n6130) );
  ANDN U6147 ( .A(n6140), .B(n6141), .Z(n6139) );
  XNOR U6148 ( .A(n6142), .B(n6138), .Z(n6140) );
  IV U6149 ( .A(n4038), .Z(mod_mult_o[101]) );
  XOR U6150 ( .A(n6143), .B(n6144), .Z(n4038) );
  IV U6151 ( .A(n4041), .Z(mod_mult_o[1019]) );
  XOR U6152 ( .A(n6141), .B(n6142), .Z(n4041) );
  NAND U6153 ( .A(n6145), .B(e_input[1019]), .Z(n6142) );
  NAND U6154 ( .A(n6112), .B(e_input[1019]), .Z(n6145) );
  XOR U6155 ( .A(n6146), .B(n6147), .Z(n6141) );
  IV U6156 ( .A(n6138), .Z(n6146) );
  XOR U6157 ( .A(n6148), .B(n6149), .Z(n6138) );
  ANDN U6158 ( .A(n6150), .B(n6151), .Z(n6149) );
  XNOR U6159 ( .A(n6152), .B(n6148), .Z(n6150) );
  IV U6160 ( .A(n4044), .Z(mod_mult_o[1018]) );
  XOR U6161 ( .A(n6151), .B(n6152), .Z(n4044) );
  NAND U6162 ( .A(n6153), .B(e_input[1018]), .Z(n6152) );
  NAND U6163 ( .A(n6112), .B(e_input[1018]), .Z(n6153) );
  XOR U6164 ( .A(n6154), .B(n6155), .Z(n6151) );
  IV U6165 ( .A(n6148), .Z(n6154) );
  XOR U6166 ( .A(n6156), .B(n6157), .Z(n6148) );
  ANDN U6167 ( .A(n6158), .B(n6159), .Z(n6157) );
  XNOR U6168 ( .A(n6160), .B(n6156), .Z(n6158) );
  IV U6169 ( .A(n4047), .Z(mod_mult_o[1017]) );
  XOR U6170 ( .A(n6159), .B(n6160), .Z(n4047) );
  NAND U6171 ( .A(n6161), .B(e_input[1017]), .Z(n6160) );
  NAND U6172 ( .A(n6112), .B(e_input[1017]), .Z(n6161) );
  XOR U6173 ( .A(n6162), .B(n6163), .Z(n6159) );
  IV U6174 ( .A(n6156), .Z(n6162) );
  XOR U6175 ( .A(n6164), .B(n6165), .Z(n6156) );
  ANDN U6176 ( .A(n6166), .B(n6167), .Z(n6165) );
  XNOR U6177 ( .A(n6168), .B(n6164), .Z(n6166) );
  IV U6178 ( .A(n4050), .Z(mod_mult_o[1016]) );
  XOR U6179 ( .A(n6167), .B(n6168), .Z(n4050) );
  NAND U6180 ( .A(n6169), .B(e_input[1016]), .Z(n6168) );
  NAND U6181 ( .A(n6112), .B(e_input[1016]), .Z(n6169) );
  XOR U6182 ( .A(n6170), .B(n6171), .Z(n6167) );
  IV U6183 ( .A(n6164), .Z(n6170) );
  XOR U6184 ( .A(n6172), .B(n6173), .Z(n6164) );
  ANDN U6185 ( .A(n6174), .B(n6175), .Z(n6173) );
  XNOR U6186 ( .A(n6176), .B(n6172), .Z(n6174) );
  IV U6187 ( .A(n4053), .Z(mod_mult_o[1015]) );
  XOR U6188 ( .A(n6175), .B(n6176), .Z(n4053) );
  NAND U6189 ( .A(n6177), .B(e_input[1015]), .Z(n6176) );
  NAND U6190 ( .A(n6112), .B(e_input[1015]), .Z(n6177) );
  XOR U6191 ( .A(n6178), .B(n6179), .Z(n6175) );
  IV U6192 ( .A(n6172), .Z(n6178) );
  XOR U6193 ( .A(n6180), .B(n6181), .Z(n6172) );
  ANDN U6194 ( .A(n6182), .B(n6183), .Z(n6181) );
  XNOR U6195 ( .A(n6184), .B(n6180), .Z(n6182) );
  IV U6196 ( .A(n4056), .Z(mod_mult_o[1014]) );
  XOR U6197 ( .A(n6183), .B(n6184), .Z(n4056) );
  NAND U6198 ( .A(n6185), .B(e_input[1014]), .Z(n6184) );
  NAND U6199 ( .A(n6112), .B(e_input[1014]), .Z(n6185) );
  XOR U6200 ( .A(n6186), .B(n6187), .Z(n6183) );
  IV U6201 ( .A(n6180), .Z(n6186) );
  XOR U6202 ( .A(n6188), .B(n6189), .Z(n6180) );
  ANDN U6203 ( .A(n6190), .B(n6191), .Z(n6189) );
  XNOR U6204 ( .A(n6192), .B(n6188), .Z(n6190) );
  IV U6205 ( .A(n4059), .Z(mod_mult_o[1013]) );
  XOR U6206 ( .A(n6191), .B(n6192), .Z(n4059) );
  NAND U6207 ( .A(n6193), .B(e_input[1013]), .Z(n6192) );
  NAND U6208 ( .A(n6112), .B(e_input[1013]), .Z(n6193) );
  XOR U6209 ( .A(n6194), .B(n6195), .Z(n6191) );
  IV U6210 ( .A(n6188), .Z(n6194) );
  XOR U6211 ( .A(n6196), .B(n6197), .Z(n6188) );
  ANDN U6212 ( .A(n6198), .B(n6199), .Z(n6197) );
  XNOR U6213 ( .A(n6200), .B(n6196), .Z(n6198) );
  IV U6214 ( .A(n4062), .Z(mod_mult_o[1012]) );
  XOR U6215 ( .A(n6199), .B(n6200), .Z(n4062) );
  NAND U6216 ( .A(n6201), .B(e_input[1012]), .Z(n6200) );
  NAND U6217 ( .A(n6112), .B(e_input[1012]), .Z(n6201) );
  XOR U6218 ( .A(n6202), .B(n6203), .Z(n6199) );
  IV U6219 ( .A(n6196), .Z(n6202) );
  XOR U6220 ( .A(n6204), .B(n6205), .Z(n6196) );
  ANDN U6221 ( .A(n6206), .B(n6207), .Z(n6205) );
  XNOR U6222 ( .A(n6208), .B(n6204), .Z(n6206) );
  IV U6223 ( .A(n4065), .Z(mod_mult_o[1011]) );
  XOR U6224 ( .A(n6207), .B(n6208), .Z(n4065) );
  NAND U6225 ( .A(n6209), .B(e_input[1011]), .Z(n6208) );
  NAND U6226 ( .A(n6112), .B(e_input[1011]), .Z(n6209) );
  XOR U6227 ( .A(n6210), .B(n6211), .Z(n6207) );
  IV U6228 ( .A(n6204), .Z(n6210) );
  XOR U6229 ( .A(n6212), .B(n6213), .Z(n6204) );
  ANDN U6230 ( .A(n6214), .B(n6215), .Z(n6213) );
  XNOR U6231 ( .A(n6216), .B(n6212), .Z(n6214) );
  IV U6232 ( .A(n4068), .Z(mod_mult_o[1010]) );
  XOR U6233 ( .A(n6215), .B(n6216), .Z(n4068) );
  NAND U6234 ( .A(n6217), .B(e_input[1010]), .Z(n6216) );
  NAND U6235 ( .A(n6112), .B(e_input[1010]), .Z(n6217) );
  XOR U6236 ( .A(n6218), .B(n6219), .Z(n6215) );
  IV U6237 ( .A(n6212), .Z(n6218) );
  XOR U6238 ( .A(n6220), .B(n6221), .Z(n6212) );
  ANDN U6239 ( .A(n6222), .B(n6223), .Z(n6221) );
  XNOR U6240 ( .A(n6224), .B(n6220), .Z(n6222) );
  IV U6241 ( .A(n4071), .Z(mod_mult_o[100]) );
  XOR U6242 ( .A(n6225), .B(n6226), .Z(n4071) );
  IV U6243 ( .A(n4074), .Z(mod_mult_o[1009]) );
  XOR U6244 ( .A(n6223), .B(n6224), .Z(n4074) );
  NAND U6245 ( .A(n6227), .B(e_input[1009]), .Z(n6224) );
  NAND U6246 ( .A(n6112), .B(e_input[1009]), .Z(n6227) );
  XOR U6247 ( .A(n6228), .B(n6229), .Z(n6223) );
  IV U6248 ( .A(n6220), .Z(n6228) );
  XOR U6249 ( .A(n6230), .B(n6231), .Z(n6220) );
  ANDN U6250 ( .A(n6232), .B(n6233), .Z(n6231) );
  XNOR U6251 ( .A(n6234), .B(n6230), .Z(n6232) );
  IV U6252 ( .A(n4077), .Z(mod_mult_o[1008]) );
  XOR U6253 ( .A(n6233), .B(n6234), .Z(n4077) );
  NAND U6254 ( .A(n6235), .B(e_input[1008]), .Z(n6234) );
  NAND U6255 ( .A(n6112), .B(e_input[1008]), .Z(n6235) );
  XOR U6256 ( .A(n6236), .B(n6237), .Z(n6233) );
  IV U6257 ( .A(n6230), .Z(n6236) );
  XOR U6258 ( .A(n6238), .B(n6239), .Z(n6230) );
  ANDN U6259 ( .A(n6240), .B(n6241), .Z(n6239) );
  XNOR U6260 ( .A(n6242), .B(n6238), .Z(n6240) );
  IV U6261 ( .A(n4080), .Z(mod_mult_o[1007]) );
  XOR U6262 ( .A(n6241), .B(n6242), .Z(n4080) );
  NAND U6263 ( .A(n6243), .B(e_input[1007]), .Z(n6242) );
  NAND U6264 ( .A(n6112), .B(e_input[1007]), .Z(n6243) );
  XOR U6265 ( .A(n6244), .B(n6245), .Z(n6241) );
  IV U6266 ( .A(n6238), .Z(n6244) );
  XOR U6267 ( .A(n6246), .B(n6247), .Z(n6238) );
  ANDN U6268 ( .A(n6248), .B(n6249), .Z(n6247) );
  XNOR U6269 ( .A(n6250), .B(n6246), .Z(n6248) );
  IV U6270 ( .A(n4083), .Z(mod_mult_o[1006]) );
  XOR U6271 ( .A(n6249), .B(n6250), .Z(n4083) );
  NAND U6272 ( .A(n6251), .B(e_input[1006]), .Z(n6250) );
  NAND U6273 ( .A(n6112), .B(e_input[1006]), .Z(n6251) );
  XOR U6274 ( .A(n6252), .B(n6253), .Z(n6249) );
  IV U6275 ( .A(n6246), .Z(n6252) );
  XOR U6276 ( .A(n6254), .B(n6255), .Z(n6246) );
  ANDN U6277 ( .A(n6256), .B(n6257), .Z(n6255) );
  XNOR U6278 ( .A(n6258), .B(n6254), .Z(n6256) );
  IV U6279 ( .A(n4086), .Z(mod_mult_o[1005]) );
  XOR U6280 ( .A(n6257), .B(n6258), .Z(n4086) );
  NAND U6281 ( .A(n6259), .B(e_input[1005]), .Z(n6258) );
  NAND U6282 ( .A(n6112), .B(e_input[1005]), .Z(n6259) );
  XOR U6283 ( .A(n6260), .B(n6261), .Z(n6257) );
  IV U6284 ( .A(n6254), .Z(n6260) );
  XOR U6285 ( .A(n6262), .B(n6263), .Z(n6254) );
  ANDN U6286 ( .A(n6264), .B(n6265), .Z(n6263) );
  XNOR U6287 ( .A(n6266), .B(n6262), .Z(n6264) );
  IV U6288 ( .A(n4089), .Z(mod_mult_o[1004]) );
  XOR U6289 ( .A(n6265), .B(n6266), .Z(n4089) );
  NAND U6290 ( .A(n6267), .B(e_input[1004]), .Z(n6266) );
  NAND U6291 ( .A(n6112), .B(e_input[1004]), .Z(n6267) );
  XOR U6292 ( .A(n6268), .B(n6269), .Z(n6265) );
  IV U6293 ( .A(n6262), .Z(n6268) );
  XOR U6294 ( .A(n6270), .B(n6271), .Z(n6262) );
  ANDN U6295 ( .A(n6272), .B(n6273), .Z(n6271) );
  XNOR U6296 ( .A(n6274), .B(n6270), .Z(n6272) );
  IV U6297 ( .A(n4092), .Z(mod_mult_o[1003]) );
  XOR U6298 ( .A(n6273), .B(n6274), .Z(n4092) );
  NAND U6299 ( .A(n6275), .B(e_input[1003]), .Z(n6274) );
  NAND U6300 ( .A(n6112), .B(e_input[1003]), .Z(n6275) );
  XOR U6301 ( .A(n6276), .B(n6277), .Z(n6273) );
  IV U6302 ( .A(n6270), .Z(n6276) );
  XOR U6303 ( .A(n6278), .B(n6279), .Z(n6270) );
  ANDN U6304 ( .A(n6280), .B(n6281), .Z(n6279) );
  XNOR U6305 ( .A(n6282), .B(n6278), .Z(n6280) );
  IV U6306 ( .A(n4095), .Z(mod_mult_o[1002]) );
  XOR U6307 ( .A(n6281), .B(n6282), .Z(n4095) );
  NAND U6308 ( .A(n6283), .B(e_input[1002]), .Z(n6282) );
  NAND U6309 ( .A(n6112), .B(e_input[1002]), .Z(n6283) );
  XOR U6310 ( .A(n6284), .B(n6285), .Z(n6281) );
  IV U6311 ( .A(n6278), .Z(n6284) );
  XOR U6312 ( .A(n6286), .B(n6287), .Z(n6278) );
  ANDN U6313 ( .A(n6288), .B(n6289), .Z(n6287) );
  XNOR U6314 ( .A(n6290), .B(n6286), .Z(n6288) );
  IV U6315 ( .A(n4098), .Z(mod_mult_o[1001]) );
  XOR U6316 ( .A(n6289), .B(n6290), .Z(n4098) );
  NAND U6317 ( .A(n6291), .B(e_input[1001]), .Z(n6290) );
  NAND U6318 ( .A(n6112), .B(e_input[1001]), .Z(n6291) );
  XOR U6319 ( .A(n6292), .B(n6293), .Z(n6289) );
  IV U6320 ( .A(n6286), .Z(n6292) );
  XOR U6321 ( .A(n6294), .B(n6295), .Z(n6286) );
  ANDN U6322 ( .A(n6296), .B(n6297), .Z(n6295) );
  XNOR U6323 ( .A(n6298), .B(n6294), .Z(n6296) );
  IV U6324 ( .A(n4101), .Z(mod_mult_o[1000]) );
  XOR U6325 ( .A(n6297), .B(n6298), .Z(n4101) );
  NAND U6326 ( .A(n6299), .B(e_input[1000]), .Z(n6298) );
  NAND U6327 ( .A(n6112), .B(e_input[1000]), .Z(n6299) );
  XOR U6328 ( .A(n6300), .B(n6301), .Z(n6297) );
  IV U6329 ( .A(n6294), .Z(n6300) );
  XOR U6330 ( .A(n6302), .B(n6303), .Z(n6294) );
  ANDN U6331 ( .A(n6304), .B(n4121), .Z(n6303) );
  XOR U6332 ( .A(n6305), .B(n6306), .Z(n4121) );
  IV U6333 ( .A(n6302), .Z(n6305) );
  XNOR U6334 ( .A(n4122), .B(n6302), .Z(n6304) );
  NAND U6335 ( .A(n6307), .B(e_input[999]), .Z(n4122) );
  NAND U6336 ( .A(n6112), .B(e_input[999]), .Z(n6307) );
  XOR U6337 ( .A(n6308), .B(n6309), .Z(n6302) );
  ANDN U6338 ( .A(n6310), .B(n4123), .Z(n6309) );
  XOR U6339 ( .A(n6311), .B(n6312), .Z(n4123) );
  IV U6340 ( .A(n6308), .Z(n6311) );
  XNOR U6341 ( .A(n4124), .B(n6308), .Z(n6310) );
  NAND U6342 ( .A(n6313), .B(e_input[998]), .Z(n4124) );
  NAND U6343 ( .A(n6112), .B(e_input[998]), .Z(n6313) );
  XOR U6344 ( .A(n6314), .B(n6315), .Z(n6308) );
  ANDN U6345 ( .A(n6316), .B(n4125), .Z(n6315) );
  XOR U6346 ( .A(n6317), .B(n6318), .Z(n4125) );
  IV U6347 ( .A(n6314), .Z(n6317) );
  XNOR U6348 ( .A(n4126), .B(n6314), .Z(n6316) );
  NAND U6349 ( .A(n6319), .B(e_input[997]), .Z(n4126) );
  NAND U6350 ( .A(n6112), .B(e_input[997]), .Z(n6319) );
  XOR U6351 ( .A(n6320), .B(n6321), .Z(n6314) );
  ANDN U6352 ( .A(n6322), .B(n4127), .Z(n6321) );
  XOR U6353 ( .A(n6323), .B(n6324), .Z(n4127) );
  IV U6354 ( .A(n6320), .Z(n6323) );
  XNOR U6355 ( .A(n4128), .B(n6320), .Z(n6322) );
  NAND U6356 ( .A(n6325), .B(e_input[996]), .Z(n4128) );
  NAND U6357 ( .A(n6112), .B(e_input[996]), .Z(n6325) );
  XOR U6358 ( .A(n6326), .B(n6327), .Z(n6320) );
  ANDN U6359 ( .A(n6328), .B(n4129), .Z(n6327) );
  XOR U6360 ( .A(n6329), .B(n6330), .Z(n4129) );
  IV U6361 ( .A(n6326), .Z(n6329) );
  XNOR U6362 ( .A(n4130), .B(n6326), .Z(n6328) );
  NAND U6363 ( .A(n6331), .B(e_input[995]), .Z(n4130) );
  NAND U6364 ( .A(n6112), .B(e_input[995]), .Z(n6331) );
  XOR U6365 ( .A(n6332), .B(n6333), .Z(n6326) );
  ANDN U6366 ( .A(n6334), .B(n4131), .Z(n6333) );
  XOR U6367 ( .A(n6335), .B(n6336), .Z(n4131) );
  IV U6368 ( .A(n6332), .Z(n6335) );
  XNOR U6369 ( .A(n4132), .B(n6332), .Z(n6334) );
  NAND U6370 ( .A(n6337), .B(e_input[994]), .Z(n4132) );
  NAND U6371 ( .A(n6112), .B(e_input[994]), .Z(n6337) );
  XOR U6372 ( .A(n6338), .B(n6339), .Z(n6332) );
  ANDN U6373 ( .A(n6340), .B(n4133), .Z(n6339) );
  XOR U6374 ( .A(n6341), .B(n6342), .Z(n4133) );
  IV U6375 ( .A(n6338), .Z(n6341) );
  XNOR U6376 ( .A(n4134), .B(n6338), .Z(n6340) );
  NAND U6377 ( .A(n6343), .B(e_input[993]), .Z(n4134) );
  NAND U6378 ( .A(n6112), .B(e_input[993]), .Z(n6343) );
  XOR U6379 ( .A(n6344), .B(n6345), .Z(n6338) );
  ANDN U6380 ( .A(n6346), .B(n4135), .Z(n6345) );
  XOR U6381 ( .A(n6347), .B(n6348), .Z(n4135) );
  IV U6382 ( .A(n6344), .Z(n6347) );
  XNOR U6383 ( .A(n4136), .B(n6344), .Z(n6346) );
  NAND U6384 ( .A(n6349), .B(e_input[992]), .Z(n4136) );
  NAND U6385 ( .A(n6112), .B(e_input[992]), .Z(n6349) );
  XOR U6386 ( .A(n6350), .B(n6351), .Z(n6344) );
  ANDN U6387 ( .A(n6352), .B(n4137), .Z(n6351) );
  XOR U6388 ( .A(n6353), .B(n6354), .Z(n4137) );
  IV U6389 ( .A(n6350), .Z(n6353) );
  XNOR U6390 ( .A(n4138), .B(n6350), .Z(n6352) );
  NAND U6391 ( .A(n6355), .B(e_input[991]), .Z(n4138) );
  NAND U6392 ( .A(n6112), .B(e_input[991]), .Z(n6355) );
  XOR U6393 ( .A(n6356), .B(n6357), .Z(n6350) );
  ANDN U6394 ( .A(n6358), .B(n4139), .Z(n6357) );
  XOR U6395 ( .A(n6359), .B(n6360), .Z(n4139) );
  IV U6396 ( .A(n6356), .Z(n6359) );
  XNOR U6397 ( .A(n4140), .B(n6356), .Z(n6358) );
  NAND U6398 ( .A(n6361), .B(e_input[990]), .Z(n4140) );
  NAND U6399 ( .A(n6112), .B(e_input[990]), .Z(n6361) );
  XOR U6400 ( .A(n6362), .B(n6363), .Z(n6356) );
  ANDN U6401 ( .A(n6364), .B(n4143), .Z(n6363) );
  XOR U6402 ( .A(n6365), .B(n6366), .Z(n4143) );
  IV U6403 ( .A(n6362), .Z(n6365) );
  XNOR U6404 ( .A(n4144), .B(n6362), .Z(n6364) );
  NAND U6405 ( .A(n6367), .B(e_input[989]), .Z(n4144) );
  NAND U6406 ( .A(n6112), .B(e_input[989]), .Z(n6367) );
  XOR U6407 ( .A(n6368), .B(n6369), .Z(n6362) );
  ANDN U6408 ( .A(n6370), .B(n4145), .Z(n6369) );
  XOR U6409 ( .A(n6371), .B(n6372), .Z(n4145) );
  IV U6410 ( .A(n6368), .Z(n6371) );
  XNOR U6411 ( .A(n4146), .B(n6368), .Z(n6370) );
  NAND U6412 ( .A(n6373), .B(e_input[988]), .Z(n4146) );
  NAND U6413 ( .A(n6112), .B(e_input[988]), .Z(n6373) );
  XOR U6414 ( .A(n6374), .B(n6375), .Z(n6368) );
  ANDN U6415 ( .A(n6376), .B(n4147), .Z(n6375) );
  XOR U6416 ( .A(n6377), .B(n6378), .Z(n4147) );
  IV U6417 ( .A(n6374), .Z(n6377) );
  XNOR U6418 ( .A(n4148), .B(n6374), .Z(n6376) );
  NAND U6419 ( .A(n6379), .B(e_input[987]), .Z(n4148) );
  NAND U6420 ( .A(n6112), .B(e_input[987]), .Z(n6379) );
  XOR U6421 ( .A(n6380), .B(n6381), .Z(n6374) );
  ANDN U6422 ( .A(n6382), .B(n4149), .Z(n6381) );
  XOR U6423 ( .A(n6383), .B(n6384), .Z(n4149) );
  IV U6424 ( .A(n6380), .Z(n6383) );
  XNOR U6425 ( .A(n4150), .B(n6380), .Z(n6382) );
  NAND U6426 ( .A(n6385), .B(e_input[986]), .Z(n4150) );
  NAND U6427 ( .A(n6112), .B(e_input[986]), .Z(n6385) );
  XOR U6428 ( .A(n6386), .B(n6387), .Z(n6380) );
  ANDN U6429 ( .A(n6388), .B(n4151), .Z(n6387) );
  XOR U6430 ( .A(n6389), .B(n6390), .Z(n4151) );
  IV U6431 ( .A(n6386), .Z(n6389) );
  XNOR U6432 ( .A(n4152), .B(n6386), .Z(n6388) );
  NAND U6433 ( .A(n6391), .B(e_input[985]), .Z(n4152) );
  NAND U6434 ( .A(n6112), .B(e_input[985]), .Z(n6391) );
  XOR U6435 ( .A(n6392), .B(n6393), .Z(n6386) );
  ANDN U6436 ( .A(n6394), .B(n4153), .Z(n6393) );
  XOR U6437 ( .A(n6395), .B(n6396), .Z(n4153) );
  IV U6438 ( .A(n6392), .Z(n6395) );
  XNOR U6439 ( .A(n4154), .B(n6392), .Z(n6394) );
  NAND U6440 ( .A(n6397), .B(e_input[984]), .Z(n4154) );
  NAND U6441 ( .A(n6112), .B(e_input[984]), .Z(n6397) );
  XOR U6442 ( .A(n6398), .B(n6399), .Z(n6392) );
  ANDN U6443 ( .A(n6400), .B(n4155), .Z(n6399) );
  XOR U6444 ( .A(n6401), .B(n6402), .Z(n4155) );
  IV U6445 ( .A(n6398), .Z(n6401) );
  XNOR U6446 ( .A(n4156), .B(n6398), .Z(n6400) );
  NAND U6447 ( .A(n6403), .B(e_input[983]), .Z(n4156) );
  NAND U6448 ( .A(n6112), .B(e_input[983]), .Z(n6403) );
  XOR U6449 ( .A(n6404), .B(n6405), .Z(n6398) );
  ANDN U6450 ( .A(n6406), .B(n4157), .Z(n6405) );
  XOR U6451 ( .A(n6407), .B(n6408), .Z(n4157) );
  IV U6452 ( .A(n6404), .Z(n6407) );
  XNOR U6453 ( .A(n4158), .B(n6404), .Z(n6406) );
  NAND U6454 ( .A(n6409), .B(e_input[982]), .Z(n4158) );
  NAND U6455 ( .A(n6112), .B(e_input[982]), .Z(n6409) );
  XOR U6456 ( .A(n6410), .B(n6411), .Z(n6404) );
  ANDN U6457 ( .A(n6412), .B(n4159), .Z(n6411) );
  XOR U6458 ( .A(n6413), .B(n6414), .Z(n4159) );
  IV U6459 ( .A(n6410), .Z(n6413) );
  XNOR U6460 ( .A(n4160), .B(n6410), .Z(n6412) );
  NAND U6461 ( .A(n6415), .B(e_input[981]), .Z(n4160) );
  NAND U6462 ( .A(n6112), .B(e_input[981]), .Z(n6415) );
  XOR U6463 ( .A(n6416), .B(n6417), .Z(n6410) );
  ANDN U6464 ( .A(n6418), .B(n4161), .Z(n6417) );
  XOR U6465 ( .A(n6419), .B(n6420), .Z(n4161) );
  IV U6466 ( .A(n6416), .Z(n6419) );
  XNOR U6467 ( .A(n4162), .B(n6416), .Z(n6418) );
  NAND U6468 ( .A(n6421), .B(e_input[980]), .Z(n4162) );
  NAND U6469 ( .A(n6112), .B(e_input[980]), .Z(n6421) );
  XOR U6470 ( .A(n6422), .B(n6423), .Z(n6416) );
  ANDN U6471 ( .A(n6424), .B(n4165), .Z(n6423) );
  XOR U6472 ( .A(n6425), .B(n6426), .Z(n4165) );
  IV U6473 ( .A(n6422), .Z(n6425) );
  XNOR U6474 ( .A(n4166), .B(n6422), .Z(n6424) );
  NAND U6475 ( .A(n6427), .B(e_input[979]), .Z(n4166) );
  NAND U6476 ( .A(n6112), .B(e_input[979]), .Z(n6427) );
  XOR U6477 ( .A(n6428), .B(n6429), .Z(n6422) );
  ANDN U6478 ( .A(n6430), .B(n4167), .Z(n6429) );
  XOR U6479 ( .A(n6431), .B(n6432), .Z(n4167) );
  IV U6480 ( .A(n6428), .Z(n6431) );
  XNOR U6481 ( .A(n4168), .B(n6428), .Z(n6430) );
  NAND U6482 ( .A(n6433), .B(e_input[978]), .Z(n4168) );
  NAND U6483 ( .A(n6112), .B(e_input[978]), .Z(n6433) );
  XOR U6484 ( .A(n6434), .B(n6435), .Z(n6428) );
  ANDN U6485 ( .A(n6436), .B(n4169), .Z(n6435) );
  XOR U6486 ( .A(n6437), .B(n6438), .Z(n4169) );
  IV U6487 ( .A(n6434), .Z(n6437) );
  XNOR U6488 ( .A(n4170), .B(n6434), .Z(n6436) );
  NAND U6489 ( .A(n6439), .B(e_input[977]), .Z(n4170) );
  NAND U6490 ( .A(n6112), .B(e_input[977]), .Z(n6439) );
  XOR U6491 ( .A(n6440), .B(n6441), .Z(n6434) );
  ANDN U6492 ( .A(n6442), .B(n4171), .Z(n6441) );
  XOR U6493 ( .A(n6443), .B(n6444), .Z(n4171) );
  IV U6494 ( .A(n6440), .Z(n6443) );
  XNOR U6495 ( .A(n4172), .B(n6440), .Z(n6442) );
  NAND U6496 ( .A(n6445), .B(e_input[976]), .Z(n4172) );
  NAND U6497 ( .A(n6112), .B(e_input[976]), .Z(n6445) );
  XOR U6498 ( .A(n6446), .B(n6447), .Z(n6440) );
  ANDN U6499 ( .A(n6448), .B(n4173), .Z(n6447) );
  XOR U6500 ( .A(n6449), .B(n6450), .Z(n4173) );
  IV U6501 ( .A(n6446), .Z(n6449) );
  XNOR U6502 ( .A(n4174), .B(n6446), .Z(n6448) );
  NAND U6503 ( .A(n6451), .B(e_input[975]), .Z(n4174) );
  NAND U6504 ( .A(n6112), .B(e_input[975]), .Z(n6451) );
  XOR U6505 ( .A(n6452), .B(n6453), .Z(n6446) );
  ANDN U6506 ( .A(n6454), .B(n4175), .Z(n6453) );
  XOR U6507 ( .A(n6455), .B(n6456), .Z(n4175) );
  IV U6508 ( .A(n6452), .Z(n6455) );
  XNOR U6509 ( .A(n4176), .B(n6452), .Z(n6454) );
  NAND U6510 ( .A(n6457), .B(e_input[974]), .Z(n4176) );
  NAND U6511 ( .A(n6112), .B(e_input[974]), .Z(n6457) );
  XOR U6512 ( .A(n6458), .B(n6459), .Z(n6452) );
  ANDN U6513 ( .A(n6460), .B(n4177), .Z(n6459) );
  XOR U6514 ( .A(n6461), .B(n6462), .Z(n4177) );
  IV U6515 ( .A(n6458), .Z(n6461) );
  XNOR U6516 ( .A(n4178), .B(n6458), .Z(n6460) );
  NAND U6517 ( .A(n6463), .B(e_input[973]), .Z(n4178) );
  NAND U6518 ( .A(n6112), .B(e_input[973]), .Z(n6463) );
  XOR U6519 ( .A(n6464), .B(n6465), .Z(n6458) );
  ANDN U6520 ( .A(n6466), .B(n4179), .Z(n6465) );
  XOR U6521 ( .A(n6467), .B(n6468), .Z(n4179) );
  IV U6522 ( .A(n6464), .Z(n6467) );
  XNOR U6523 ( .A(n4180), .B(n6464), .Z(n6466) );
  NAND U6524 ( .A(n6469), .B(e_input[972]), .Z(n4180) );
  NAND U6525 ( .A(n6112), .B(e_input[972]), .Z(n6469) );
  XOR U6526 ( .A(n6470), .B(n6471), .Z(n6464) );
  ANDN U6527 ( .A(n6472), .B(n4181), .Z(n6471) );
  XOR U6528 ( .A(n6473), .B(n6474), .Z(n4181) );
  IV U6529 ( .A(n6470), .Z(n6473) );
  XNOR U6530 ( .A(n4182), .B(n6470), .Z(n6472) );
  NAND U6531 ( .A(n6475), .B(e_input[971]), .Z(n4182) );
  NAND U6532 ( .A(n6112), .B(e_input[971]), .Z(n6475) );
  XOR U6533 ( .A(n6476), .B(n6477), .Z(n6470) );
  ANDN U6534 ( .A(n6478), .B(n4183), .Z(n6477) );
  XOR U6535 ( .A(n6479), .B(n6480), .Z(n4183) );
  IV U6536 ( .A(n6476), .Z(n6479) );
  XNOR U6537 ( .A(n4184), .B(n6476), .Z(n6478) );
  NAND U6538 ( .A(n6481), .B(e_input[970]), .Z(n4184) );
  NAND U6539 ( .A(n6112), .B(e_input[970]), .Z(n6481) );
  XOR U6540 ( .A(n6482), .B(n6483), .Z(n6476) );
  ANDN U6541 ( .A(n6484), .B(n4187), .Z(n6483) );
  XOR U6542 ( .A(n6485), .B(n6486), .Z(n4187) );
  IV U6543 ( .A(n6482), .Z(n6485) );
  XNOR U6544 ( .A(n4188), .B(n6482), .Z(n6484) );
  NAND U6545 ( .A(n6487), .B(e_input[969]), .Z(n4188) );
  NAND U6546 ( .A(n6112), .B(e_input[969]), .Z(n6487) );
  XOR U6547 ( .A(n6488), .B(n6489), .Z(n6482) );
  ANDN U6548 ( .A(n6490), .B(n4189), .Z(n6489) );
  XOR U6549 ( .A(n6491), .B(n6492), .Z(n4189) );
  IV U6550 ( .A(n6488), .Z(n6491) );
  XNOR U6551 ( .A(n4190), .B(n6488), .Z(n6490) );
  NAND U6552 ( .A(n6493), .B(e_input[968]), .Z(n4190) );
  NAND U6553 ( .A(n6112), .B(e_input[968]), .Z(n6493) );
  XOR U6554 ( .A(n6494), .B(n6495), .Z(n6488) );
  ANDN U6555 ( .A(n6496), .B(n4191), .Z(n6495) );
  XOR U6556 ( .A(n6497), .B(n6498), .Z(n4191) );
  IV U6557 ( .A(n6494), .Z(n6497) );
  XNOR U6558 ( .A(n4192), .B(n6494), .Z(n6496) );
  NAND U6559 ( .A(n6499), .B(e_input[967]), .Z(n4192) );
  NAND U6560 ( .A(n6112), .B(e_input[967]), .Z(n6499) );
  XOR U6561 ( .A(n6500), .B(n6501), .Z(n6494) );
  ANDN U6562 ( .A(n6502), .B(n4193), .Z(n6501) );
  XOR U6563 ( .A(n6503), .B(n6504), .Z(n4193) );
  IV U6564 ( .A(n6500), .Z(n6503) );
  XNOR U6565 ( .A(n4194), .B(n6500), .Z(n6502) );
  NAND U6566 ( .A(n6505), .B(e_input[966]), .Z(n4194) );
  NAND U6567 ( .A(n6112), .B(e_input[966]), .Z(n6505) );
  XOR U6568 ( .A(n6506), .B(n6507), .Z(n6500) );
  ANDN U6569 ( .A(n6508), .B(n4195), .Z(n6507) );
  XOR U6570 ( .A(n6509), .B(n6510), .Z(n4195) );
  IV U6571 ( .A(n6506), .Z(n6509) );
  XNOR U6572 ( .A(n4196), .B(n6506), .Z(n6508) );
  NAND U6573 ( .A(n6511), .B(e_input[965]), .Z(n4196) );
  NAND U6574 ( .A(n6112), .B(e_input[965]), .Z(n6511) );
  XOR U6575 ( .A(n6512), .B(n6513), .Z(n6506) );
  ANDN U6576 ( .A(n6514), .B(n4197), .Z(n6513) );
  XOR U6577 ( .A(n6515), .B(n6516), .Z(n4197) );
  IV U6578 ( .A(n6512), .Z(n6515) );
  XNOR U6579 ( .A(n4198), .B(n6512), .Z(n6514) );
  NAND U6580 ( .A(n6517), .B(e_input[964]), .Z(n4198) );
  NAND U6581 ( .A(n6112), .B(e_input[964]), .Z(n6517) );
  XOR U6582 ( .A(n6518), .B(n6519), .Z(n6512) );
  ANDN U6583 ( .A(n6520), .B(n4199), .Z(n6519) );
  XOR U6584 ( .A(n6521), .B(n6522), .Z(n4199) );
  IV U6585 ( .A(n6518), .Z(n6521) );
  XNOR U6586 ( .A(n4200), .B(n6518), .Z(n6520) );
  NAND U6587 ( .A(n6523), .B(e_input[963]), .Z(n4200) );
  NAND U6588 ( .A(n6112), .B(e_input[963]), .Z(n6523) );
  XOR U6589 ( .A(n6524), .B(n6525), .Z(n6518) );
  ANDN U6590 ( .A(n6526), .B(n4201), .Z(n6525) );
  XOR U6591 ( .A(n6527), .B(n6528), .Z(n4201) );
  IV U6592 ( .A(n6524), .Z(n6527) );
  XNOR U6593 ( .A(n4202), .B(n6524), .Z(n6526) );
  NAND U6594 ( .A(n6529), .B(e_input[962]), .Z(n4202) );
  NAND U6595 ( .A(n6112), .B(e_input[962]), .Z(n6529) );
  XOR U6596 ( .A(n6530), .B(n6531), .Z(n6524) );
  ANDN U6597 ( .A(n6532), .B(n4203), .Z(n6531) );
  XOR U6598 ( .A(n6533), .B(n6534), .Z(n4203) );
  IV U6599 ( .A(n6530), .Z(n6533) );
  XNOR U6600 ( .A(n4204), .B(n6530), .Z(n6532) );
  NAND U6601 ( .A(n6535), .B(e_input[961]), .Z(n4204) );
  NAND U6602 ( .A(n6112), .B(e_input[961]), .Z(n6535) );
  XOR U6603 ( .A(n6536), .B(n6537), .Z(n6530) );
  ANDN U6604 ( .A(n6538), .B(n4205), .Z(n6537) );
  XOR U6605 ( .A(n6539), .B(n6540), .Z(n4205) );
  IV U6606 ( .A(n6536), .Z(n6539) );
  XNOR U6607 ( .A(n4206), .B(n6536), .Z(n6538) );
  NAND U6608 ( .A(n6541), .B(e_input[960]), .Z(n4206) );
  NAND U6609 ( .A(n6112), .B(e_input[960]), .Z(n6541) );
  XOR U6610 ( .A(n6542), .B(n6543), .Z(n6536) );
  ANDN U6611 ( .A(n6544), .B(n4209), .Z(n6543) );
  XOR U6612 ( .A(n6545), .B(n6546), .Z(n4209) );
  IV U6613 ( .A(n6542), .Z(n6545) );
  XNOR U6614 ( .A(n4210), .B(n6542), .Z(n6544) );
  NAND U6615 ( .A(n6547), .B(e_input[959]), .Z(n4210) );
  NAND U6616 ( .A(n6112), .B(e_input[959]), .Z(n6547) );
  XOR U6617 ( .A(n6548), .B(n6549), .Z(n6542) );
  ANDN U6618 ( .A(n6550), .B(n4211), .Z(n6549) );
  XOR U6619 ( .A(n6551), .B(n6552), .Z(n4211) );
  IV U6620 ( .A(n6548), .Z(n6551) );
  XNOR U6621 ( .A(n4212), .B(n6548), .Z(n6550) );
  NAND U6622 ( .A(n6553), .B(e_input[958]), .Z(n4212) );
  NAND U6623 ( .A(n6112), .B(e_input[958]), .Z(n6553) );
  XOR U6624 ( .A(n6554), .B(n6555), .Z(n6548) );
  ANDN U6625 ( .A(n6556), .B(n4213), .Z(n6555) );
  XOR U6626 ( .A(n6557), .B(n6558), .Z(n4213) );
  IV U6627 ( .A(n6554), .Z(n6557) );
  XNOR U6628 ( .A(n4214), .B(n6554), .Z(n6556) );
  NAND U6629 ( .A(n6559), .B(e_input[957]), .Z(n4214) );
  NAND U6630 ( .A(n6112), .B(e_input[957]), .Z(n6559) );
  XOR U6631 ( .A(n6560), .B(n6561), .Z(n6554) );
  ANDN U6632 ( .A(n6562), .B(n4215), .Z(n6561) );
  XOR U6633 ( .A(n6563), .B(n6564), .Z(n4215) );
  IV U6634 ( .A(n6560), .Z(n6563) );
  XNOR U6635 ( .A(n4216), .B(n6560), .Z(n6562) );
  NAND U6636 ( .A(n6565), .B(e_input[956]), .Z(n4216) );
  NAND U6637 ( .A(n6112), .B(e_input[956]), .Z(n6565) );
  XOR U6638 ( .A(n6566), .B(n6567), .Z(n6560) );
  ANDN U6639 ( .A(n6568), .B(n4217), .Z(n6567) );
  XOR U6640 ( .A(n6569), .B(n6570), .Z(n4217) );
  IV U6641 ( .A(n6566), .Z(n6569) );
  XNOR U6642 ( .A(n4218), .B(n6566), .Z(n6568) );
  NAND U6643 ( .A(n6571), .B(e_input[955]), .Z(n4218) );
  NAND U6644 ( .A(n6112), .B(e_input[955]), .Z(n6571) );
  XOR U6645 ( .A(n6572), .B(n6573), .Z(n6566) );
  ANDN U6646 ( .A(n6574), .B(n4219), .Z(n6573) );
  XOR U6647 ( .A(n6575), .B(n6576), .Z(n4219) );
  IV U6648 ( .A(n6572), .Z(n6575) );
  XNOR U6649 ( .A(n4220), .B(n6572), .Z(n6574) );
  NAND U6650 ( .A(n6577), .B(e_input[954]), .Z(n4220) );
  NAND U6651 ( .A(n6112), .B(e_input[954]), .Z(n6577) );
  XOR U6652 ( .A(n6578), .B(n6579), .Z(n6572) );
  ANDN U6653 ( .A(n6580), .B(n4221), .Z(n6579) );
  XOR U6654 ( .A(n6581), .B(n6582), .Z(n4221) );
  IV U6655 ( .A(n6578), .Z(n6581) );
  XNOR U6656 ( .A(n4222), .B(n6578), .Z(n6580) );
  NAND U6657 ( .A(n6583), .B(e_input[953]), .Z(n4222) );
  NAND U6658 ( .A(n6112), .B(e_input[953]), .Z(n6583) );
  XOR U6659 ( .A(n6584), .B(n6585), .Z(n6578) );
  ANDN U6660 ( .A(n6586), .B(n4223), .Z(n6585) );
  XOR U6661 ( .A(n6587), .B(n6588), .Z(n4223) );
  IV U6662 ( .A(n6584), .Z(n6587) );
  XNOR U6663 ( .A(n4224), .B(n6584), .Z(n6586) );
  NAND U6664 ( .A(n6589), .B(e_input[952]), .Z(n4224) );
  NAND U6665 ( .A(n6112), .B(e_input[952]), .Z(n6589) );
  XOR U6666 ( .A(n6590), .B(n6591), .Z(n6584) );
  ANDN U6667 ( .A(n6592), .B(n4225), .Z(n6591) );
  XOR U6668 ( .A(n6593), .B(n6594), .Z(n4225) );
  IV U6669 ( .A(n6590), .Z(n6593) );
  XNOR U6670 ( .A(n4226), .B(n6590), .Z(n6592) );
  NAND U6671 ( .A(n6595), .B(e_input[951]), .Z(n4226) );
  NAND U6672 ( .A(n6112), .B(e_input[951]), .Z(n6595) );
  XOR U6673 ( .A(n6596), .B(n6597), .Z(n6590) );
  ANDN U6674 ( .A(n6598), .B(n4227), .Z(n6597) );
  XOR U6675 ( .A(n6599), .B(n6600), .Z(n4227) );
  IV U6676 ( .A(n6596), .Z(n6599) );
  XNOR U6677 ( .A(n4228), .B(n6596), .Z(n6598) );
  NAND U6678 ( .A(n6601), .B(e_input[950]), .Z(n4228) );
  NAND U6679 ( .A(n6112), .B(e_input[950]), .Z(n6601) );
  XOR U6680 ( .A(n6602), .B(n6603), .Z(n6596) );
  ANDN U6681 ( .A(n6604), .B(n4231), .Z(n6603) );
  XOR U6682 ( .A(n6605), .B(n6606), .Z(n4231) );
  IV U6683 ( .A(n6602), .Z(n6605) );
  XNOR U6684 ( .A(n4232), .B(n6602), .Z(n6604) );
  NAND U6685 ( .A(n6607), .B(e_input[949]), .Z(n4232) );
  NAND U6686 ( .A(n6112), .B(e_input[949]), .Z(n6607) );
  XOR U6687 ( .A(n6608), .B(n6609), .Z(n6602) );
  ANDN U6688 ( .A(n6610), .B(n4233), .Z(n6609) );
  XOR U6689 ( .A(n6611), .B(n6612), .Z(n4233) );
  IV U6690 ( .A(n6608), .Z(n6611) );
  XNOR U6691 ( .A(n4234), .B(n6608), .Z(n6610) );
  NAND U6692 ( .A(n6613), .B(e_input[948]), .Z(n4234) );
  NAND U6693 ( .A(n6112), .B(e_input[948]), .Z(n6613) );
  XOR U6694 ( .A(n6614), .B(n6615), .Z(n6608) );
  ANDN U6695 ( .A(n6616), .B(n4235), .Z(n6615) );
  XOR U6696 ( .A(n6617), .B(n6618), .Z(n4235) );
  IV U6697 ( .A(n6614), .Z(n6617) );
  XNOR U6698 ( .A(n4236), .B(n6614), .Z(n6616) );
  NAND U6699 ( .A(n6619), .B(e_input[947]), .Z(n4236) );
  NAND U6700 ( .A(n6112), .B(e_input[947]), .Z(n6619) );
  XOR U6701 ( .A(n6620), .B(n6621), .Z(n6614) );
  ANDN U6702 ( .A(n6622), .B(n4237), .Z(n6621) );
  XOR U6703 ( .A(n6623), .B(n6624), .Z(n4237) );
  IV U6704 ( .A(n6620), .Z(n6623) );
  XNOR U6705 ( .A(n4238), .B(n6620), .Z(n6622) );
  NAND U6706 ( .A(n6625), .B(e_input[946]), .Z(n4238) );
  NAND U6707 ( .A(n6112), .B(e_input[946]), .Z(n6625) );
  XOR U6708 ( .A(n6626), .B(n6627), .Z(n6620) );
  ANDN U6709 ( .A(n6628), .B(n4239), .Z(n6627) );
  XOR U6710 ( .A(n6629), .B(n6630), .Z(n4239) );
  IV U6711 ( .A(n6626), .Z(n6629) );
  XNOR U6712 ( .A(n4240), .B(n6626), .Z(n6628) );
  NAND U6713 ( .A(n6631), .B(e_input[945]), .Z(n4240) );
  NAND U6714 ( .A(n6112), .B(e_input[945]), .Z(n6631) );
  XOR U6715 ( .A(n6632), .B(n6633), .Z(n6626) );
  ANDN U6716 ( .A(n6634), .B(n4241), .Z(n6633) );
  XOR U6717 ( .A(n6635), .B(n6636), .Z(n4241) );
  IV U6718 ( .A(n6632), .Z(n6635) );
  XNOR U6719 ( .A(n4242), .B(n6632), .Z(n6634) );
  NAND U6720 ( .A(n6637), .B(e_input[944]), .Z(n4242) );
  NAND U6721 ( .A(n6112), .B(e_input[944]), .Z(n6637) );
  XOR U6722 ( .A(n6638), .B(n6639), .Z(n6632) );
  ANDN U6723 ( .A(n6640), .B(n4243), .Z(n6639) );
  XOR U6724 ( .A(n6641), .B(n6642), .Z(n4243) );
  IV U6725 ( .A(n6638), .Z(n6641) );
  XNOR U6726 ( .A(n4244), .B(n6638), .Z(n6640) );
  NAND U6727 ( .A(n6643), .B(e_input[943]), .Z(n4244) );
  NAND U6728 ( .A(n6112), .B(e_input[943]), .Z(n6643) );
  XOR U6729 ( .A(n6644), .B(n6645), .Z(n6638) );
  ANDN U6730 ( .A(n6646), .B(n4245), .Z(n6645) );
  XOR U6731 ( .A(n6647), .B(n6648), .Z(n4245) );
  IV U6732 ( .A(n6644), .Z(n6647) );
  XNOR U6733 ( .A(n4246), .B(n6644), .Z(n6646) );
  NAND U6734 ( .A(n6649), .B(e_input[942]), .Z(n4246) );
  NAND U6735 ( .A(n6112), .B(e_input[942]), .Z(n6649) );
  XOR U6736 ( .A(n6650), .B(n6651), .Z(n6644) );
  ANDN U6737 ( .A(n6652), .B(n4247), .Z(n6651) );
  XOR U6738 ( .A(n6653), .B(n6654), .Z(n4247) );
  IV U6739 ( .A(n6650), .Z(n6653) );
  XNOR U6740 ( .A(n4248), .B(n6650), .Z(n6652) );
  NAND U6741 ( .A(n6655), .B(e_input[941]), .Z(n4248) );
  NAND U6742 ( .A(n6112), .B(e_input[941]), .Z(n6655) );
  XOR U6743 ( .A(n6656), .B(n6657), .Z(n6650) );
  ANDN U6744 ( .A(n6658), .B(n4249), .Z(n6657) );
  XOR U6745 ( .A(n6659), .B(n6660), .Z(n4249) );
  IV U6746 ( .A(n6656), .Z(n6659) );
  XNOR U6747 ( .A(n4250), .B(n6656), .Z(n6658) );
  NAND U6748 ( .A(n6661), .B(e_input[940]), .Z(n4250) );
  NAND U6749 ( .A(n6112), .B(e_input[940]), .Z(n6661) );
  XOR U6750 ( .A(n6662), .B(n6663), .Z(n6656) );
  ANDN U6751 ( .A(n6664), .B(n4253), .Z(n6663) );
  XOR U6752 ( .A(n6665), .B(n6666), .Z(n4253) );
  IV U6753 ( .A(n6662), .Z(n6665) );
  XNOR U6754 ( .A(n4254), .B(n6662), .Z(n6664) );
  NAND U6755 ( .A(n6667), .B(e_input[939]), .Z(n4254) );
  NAND U6756 ( .A(n6112), .B(e_input[939]), .Z(n6667) );
  XOR U6757 ( .A(n6668), .B(n6669), .Z(n6662) );
  ANDN U6758 ( .A(n6670), .B(n4255), .Z(n6669) );
  XOR U6759 ( .A(n6671), .B(n6672), .Z(n4255) );
  IV U6760 ( .A(n6668), .Z(n6671) );
  XNOR U6761 ( .A(n4256), .B(n6668), .Z(n6670) );
  NAND U6762 ( .A(n6673), .B(e_input[938]), .Z(n4256) );
  NAND U6763 ( .A(n6112), .B(e_input[938]), .Z(n6673) );
  XOR U6764 ( .A(n6674), .B(n6675), .Z(n6668) );
  ANDN U6765 ( .A(n6676), .B(n4257), .Z(n6675) );
  XOR U6766 ( .A(n6677), .B(n6678), .Z(n4257) );
  IV U6767 ( .A(n6674), .Z(n6677) );
  XNOR U6768 ( .A(n4258), .B(n6674), .Z(n6676) );
  NAND U6769 ( .A(n6679), .B(e_input[937]), .Z(n4258) );
  NAND U6770 ( .A(n6112), .B(e_input[937]), .Z(n6679) );
  XOR U6771 ( .A(n6680), .B(n6681), .Z(n6674) );
  ANDN U6772 ( .A(n6682), .B(n4259), .Z(n6681) );
  XOR U6773 ( .A(n6683), .B(n6684), .Z(n4259) );
  IV U6774 ( .A(n6680), .Z(n6683) );
  XNOR U6775 ( .A(n4260), .B(n6680), .Z(n6682) );
  NAND U6776 ( .A(n6685), .B(e_input[936]), .Z(n4260) );
  NAND U6777 ( .A(n6112), .B(e_input[936]), .Z(n6685) );
  XOR U6778 ( .A(n6686), .B(n6687), .Z(n6680) );
  ANDN U6779 ( .A(n6688), .B(n4261), .Z(n6687) );
  XOR U6780 ( .A(n6689), .B(n6690), .Z(n4261) );
  IV U6781 ( .A(n6686), .Z(n6689) );
  XNOR U6782 ( .A(n4262), .B(n6686), .Z(n6688) );
  NAND U6783 ( .A(n6691), .B(e_input[935]), .Z(n4262) );
  NAND U6784 ( .A(n6112), .B(e_input[935]), .Z(n6691) );
  XOR U6785 ( .A(n6692), .B(n6693), .Z(n6686) );
  ANDN U6786 ( .A(n6694), .B(n4263), .Z(n6693) );
  XOR U6787 ( .A(n6695), .B(n6696), .Z(n4263) );
  IV U6788 ( .A(n6692), .Z(n6695) );
  XNOR U6789 ( .A(n4264), .B(n6692), .Z(n6694) );
  NAND U6790 ( .A(n6697), .B(e_input[934]), .Z(n4264) );
  NAND U6791 ( .A(n6112), .B(e_input[934]), .Z(n6697) );
  XOR U6792 ( .A(n6698), .B(n6699), .Z(n6692) );
  ANDN U6793 ( .A(n6700), .B(n4265), .Z(n6699) );
  XOR U6794 ( .A(n6701), .B(n6702), .Z(n4265) );
  IV U6795 ( .A(n6698), .Z(n6701) );
  XNOR U6796 ( .A(n4266), .B(n6698), .Z(n6700) );
  NAND U6797 ( .A(n6703), .B(e_input[933]), .Z(n4266) );
  NAND U6798 ( .A(n6112), .B(e_input[933]), .Z(n6703) );
  XOR U6799 ( .A(n6704), .B(n6705), .Z(n6698) );
  ANDN U6800 ( .A(n6706), .B(n4267), .Z(n6705) );
  XOR U6801 ( .A(n6707), .B(n6708), .Z(n4267) );
  IV U6802 ( .A(n6704), .Z(n6707) );
  XNOR U6803 ( .A(n4268), .B(n6704), .Z(n6706) );
  NAND U6804 ( .A(n6709), .B(e_input[932]), .Z(n4268) );
  NAND U6805 ( .A(n6112), .B(e_input[932]), .Z(n6709) );
  XOR U6806 ( .A(n6710), .B(n6711), .Z(n6704) );
  ANDN U6807 ( .A(n6712), .B(n4269), .Z(n6711) );
  XOR U6808 ( .A(n6713), .B(n6714), .Z(n4269) );
  IV U6809 ( .A(n6710), .Z(n6713) );
  XNOR U6810 ( .A(n4270), .B(n6710), .Z(n6712) );
  NAND U6811 ( .A(n6715), .B(e_input[931]), .Z(n4270) );
  NAND U6812 ( .A(n6112), .B(e_input[931]), .Z(n6715) );
  XOR U6813 ( .A(n6716), .B(n6717), .Z(n6710) );
  ANDN U6814 ( .A(n6718), .B(n4271), .Z(n6717) );
  XOR U6815 ( .A(n6719), .B(n6720), .Z(n4271) );
  IV U6816 ( .A(n6716), .Z(n6719) );
  XNOR U6817 ( .A(n4272), .B(n6716), .Z(n6718) );
  NAND U6818 ( .A(n6721), .B(e_input[930]), .Z(n4272) );
  NAND U6819 ( .A(n6112), .B(e_input[930]), .Z(n6721) );
  XOR U6820 ( .A(n6722), .B(n6723), .Z(n6716) );
  ANDN U6821 ( .A(n6724), .B(n4275), .Z(n6723) );
  XOR U6822 ( .A(n6725), .B(n6726), .Z(n4275) );
  IV U6823 ( .A(n6722), .Z(n6725) );
  XNOR U6824 ( .A(n4276), .B(n6722), .Z(n6724) );
  NAND U6825 ( .A(n6727), .B(e_input[929]), .Z(n4276) );
  NAND U6826 ( .A(n6112), .B(e_input[929]), .Z(n6727) );
  XOR U6827 ( .A(n6728), .B(n6729), .Z(n6722) );
  ANDN U6828 ( .A(n6730), .B(n4277), .Z(n6729) );
  XOR U6829 ( .A(n6731), .B(n6732), .Z(n4277) );
  IV U6830 ( .A(n6728), .Z(n6731) );
  XNOR U6831 ( .A(n4278), .B(n6728), .Z(n6730) );
  NAND U6832 ( .A(n6733), .B(e_input[928]), .Z(n4278) );
  NAND U6833 ( .A(n6112), .B(e_input[928]), .Z(n6733) );
  XOR U6834 ( .A(n6734), .B(n6735), .Z(n6728) );
  ANDN U6835 ( .A(n6736), .B(n4279), .Z(n6735) );
  XOR U6836 ( .A(n6737), .B(n6738), .Z(n4279) );
  IV U6837 ( .A(n6734), .Z(n6737) );
  XNOR U6838 ( .A(n4280), .B(n6734), .Z(n6736) );
  NAND U6839 ( .A(n6739), .B(e_input[927]), .Z(n4280) );
  NAND U6840 ( .A(n6112), .B(e_input[927]), .Z(n6739) );
  XOR U6841 ( .A(n6740), .B(n6741), .Z(n6734) );
  ANDN U6842 ( .A(n6742), .B(n4281), .Z(n6741) );
  XOR U6843 ( .A(n6743), .B(n6744), .Z(n4281) );
  IV U6844 ( .A(n6740), .Z(n6743) );
  XNOR U6845 ( .A(n4282), .B(n6740), .Z(n6742) );
  NAND U6846 ( .A(n6745), .B(e_input[926]), .Z(n4282) );
  NAND U6847 ( .A(n6112), .B(e_input[926]), .Z(n6745) );
  XOR U6848 ( .A(n6746), .B(n6747), .Z(n6740) );
  ANDN U6849 ( .A(n6748), .B(n4283), .Z(n6747) );
  XOR U6850 ( .A(n6749), .B(n6750), .Z(n4283) );
  IV U6851 ( .A(n6746), .Z(n6749) );
  XNOR U6852 ( .A(n4284), .B(n6746), .Z(n6748) );
  NAND U6853 ( .A(n6751), .B(e_input[925]), .Z(n4284) );
  NAND U6854 ( .A(n6112), .B(e_input[925]), .Z(n6751) );
  XOR U6855 ( .A(n6752), .B(n6753), .Z(n6746) );
  ANDN U6856 ( .A(n6754), .B(n4285), .Z(n6753) );
  XOR U6857 ( .A(n6755), .B(n6756), .Z(n4285) );
  IV U6858 ( .A(n6752), .Z(n6755) );
  XNOR U6859 ( .A(n4286), .B(n6752), .Z(n6754) );
  NAND U6860 ( .A(n6757), .B(e_input[924]), .Z(n4286) );
  NAND U6861 ( .A(n6112), .B(e_input[924]), .Z(n6757) );
  XOR U6862 ( .A(n6758), .B(n6759), .Z(n6752) );
  ANDN U6863 ( .A(n6760), .B(n4287), .Z(n6759) );
  XOR U6864 ( .A(n6761), .B(n6762), .Z(n4287) );
  IV U6865 ( .A(n6758), .Z(n6761) );
  XNOR U6866 ( .A(n4288), .B(n6758), .Z(n6760) );
  NAND U6867 ( .A(n6763), .B(e_input[923]), .Z(n4288) );
  NAND U6868 ( .A(n6112), .B(e_input[923]), .Z(n6763) );
  XOR U6869 ( .A(n6764), .B(n6765), .Z(n6758) );
  ANDN U6870 ( .A(n6766), .B(n4289), .Z(n6765) );
  XOR U6871 ( .A(n6767), .B(n6768), .Z(n4289) );
  IV U6872 ( .A(n6764), .Z(n6767) );
  XNOR U6873 ( .A(n4290), .B(n6764), .Z(n6766) );
  NAND U6874 ( .A(n6769), .B(e_input[922]), .Z(n4290) );
  NAND U6875 ( .A(n6112), .B(e_input[922]), .Z(n6769) );
  XOR U6876 ( .A(n6770), .B(n6771), .Z(n6764) );
  ANDN U6877 ( .A(n6772), .B(n4291), .Z(n6771) );
  XOR U6878 ( .A(n6773), .B(n6774), .Z(n4291) );
  IV U6879 ( .A(n6770), .Z(n6773) );
  XNOR U6880 ( .A(n4292), .B(n6770), .Z(n6772) );
  NAND U6881 ( .A(n6775), .B(e_input[921]), .Z(n4292) );
  NAND U6882 ( .A(n6112), .B(e_input[921]), .Z(n6775) );
  XOR U6883 ( .A(n6776), .B(n6777), .Z(n6770) );
  ANDN U6884 ( .A(n6778), .B(n4293), .Z(n6777) );
  XOR U6885 ( .A(n6779), .B(n6780), .Z(n4293) );
  IV U6886 ( .A(n6776), .Z(n6779) );
  XNOR U6887 ( .A(n4294), .B(n6776), .Z(n6778) );
  NAND U6888 ( .A(n6781), .B(e_input[920]), .Z(n4294) );
  NAND U6889 ( .A(n6112), .B(e_input[920]), .Z(n6781) );
  XOR U6890 ( .A(n6782), .B(n6783), .Z(n6776) );
  ANDN U6891 ( .A(n6784), .B(n4297), .Z(n6783) );
  XOR U6892 ( .A(n6785), .B(n6786), .Z(n4297) );
  IV U6893 ( .A(n6782), .Z(n6785) );
  XNOR U6894 ( .A(n4298), .B(n6782), .Z(n6784) );
  NAND U6895 ( .A(n6787), .B(e_input[919]), .Z(n4298) );
  NAND U6896 ( .A(n6112), .B(e_input[919]), .Z(n6787) );
  XOR U6897 ( .A(n6788), .B(n6789), .Z(n6782) );
  ANDN U6898 ( .A(n6790), .B(n4299), .Z(n6789) );
  XOR U6899 ( .A(n6791), .B(n6792), .Z(n4299) );
  IV U6900 ( .A(n6788), .Z(n6791) );
  XNOR U6901 ( .A(n4300), .B(n6788), .Z(n6790) );
  NAND U6902 ( .A(n6793), .B(e_input[918]), .Z(n4300) );
  NAND U6903 ( .A(n6112), .B(e_input[918]), .Z(n6793) );
  XOR U6904 ( .A(n6794), .B(n6795), .Z(n6788) );
  ANDN U6905 ( .A(n6796), .B(n4301), .Z(n6795) );
  XOR U6906 ( .A(n6797), .B(n6798), .Z(n4301) );
  IV U6907 ( .A(n6794), .Z(n6797) );
  XNOR U6908 ( .A(n4302), .B(n6794), .Z(n6796) );
  NAND U6909 ( .A(n6799), .B(e_input[917]), .Z(n4302) );
  NAND U6910 ( .A(n6112), .B(e_input[917]), .Z(n6799) );
  XOR U6911 ( .A(n6800), .B(n6801), .Z(n6794) );
  ANDN U6912 ( .A(n6802), .B(n4303), .Z(n6801) );
  XOR U6913 ( .A(n6803), .B(n6804), .Z(n4303) );
  IV U6914 ( .A(n6800), .Z(n6803) );
  XNOR U6915 ( .A(n4304), .B(n6800), .Z(n6802) );
  NAND U6916 ( .A(n6805), .B(e_input[916]), .Z(n4304) );
  NAND U6917 ( .A(n6112), .B(e_input[916]), .Z(n6805) );
  XOR U6918 ( .A(n6806), .B(n6807), .Z(n6800) );
  ANDN U6919 ( .A(n6808), .B(n4305), .Z(n6807) );
  XOR U6920 ( .A(n6809), .B(n6810), .Z(n4305) );
  IV U6921 ( .A(n6806), .Z(n6809) );
  XNOR U6922 ( .A(n4306), .B(n6806), .Z(n6808) );
  NAND U6923 ( .A(n6811), .B(e_input[915]), .Z(n4306) );
  NAND U6924 ( .A(n6112), .B(e_input[915]), .Z(n6811) );
  XOR U6925 ( .A(n6812), .B(n6813), .Z(n6806) );
  ANDN U6926 ( .A(n6814), .B(n4307), .Z(n6813) );
  XOR U6927 ( .A(n6815), .B(n6816), .Z(n4307) );
  IV U6928 ( .A(n6812), .Z(n6815) );
  XNOR U6929 ( .A(n4308), .B(n6812), .Z(n6814) );
  NAND U6930 ( .A(n6817), .B(e_input[914]), .Z(n4308) );
  NAND U6931 ( .A(n6112), .B(e_input[914]), .Z(n6817) );
  XOR U6932 ( .A(n6818), .B(n6819), .Z(n6812) );
  ANDN U6933 ( .A(n6820), .B(n4309), .Z(n6819) );
  XOR U6934 ( .A(n6821), .B(n6822), .Z(n4309) );
  IV U6935 ( .A(n6818), .Z(n6821) );
  XNOR U6936 ( .A(n4310), .B(n6818), .Z(n6820) );
  NAND U6937 ( .A(n6823), .B(e_input[913]), .Z(n4310) );
  NAND U6938 ( .A(n6112), .B(e_input[913]), .Z(n6823) );
  XOR U6939 ( .A(n6824), .B(n6825), .Z(n6818) );
  ANDN U6940 ( .A(n6826), .B(n4311), .Z(n6825) );
  XOR U6941 ( .A(n6827), .B(n6828), .Z(n4311) );
  IV U6942 ( .A(n6824), .Z(n6827) );
  XNOR U6943 ( .A(n4312), .B(n6824), .Z(n6826) );
  NAND U6944 ( .A(n6829), .B(e_input[912]), .Z(n4312) );
  NAND U6945 ( .A(n6112), .B(e_input[912]), .Z(n6829) );
  XOR U6946 ( .A(n6830), .B(n6831), .Z(n6824) );
  ANDN U6947 ( .A(n6832), .B(n4313), .Z(n6831) );
  XOR U6948 ( .A(n6833), .B(n6834), .Z(n4313) );
  IV U6949 ( .A(n6830), .Z(n6833) );
  XNOR U6950 ( .A(n4314), .B(n6830), .Z(n6832) );
  NAND U6951 ( .A(n6835), .B(e_input[911]), .Z(n4314) );
  NAND U6952 ( .A(n6112), .B(e_input[911]), .Z(n6835) );
  XOR U6953 ( .A(n6836), .B(n6837), .Z(n6830) );
  ANDN U6954 ( .A(n6838), .B(n4315), .Z(n6837) );
  XOR U6955 ( .A(n6839), .B(n6840), .Z(n4315) );
  IV U6956 ( .A(n6836), .Z(n6839) );
  XNOR U6957 ( .A(n4316), .B(n6836), .Z(n6838) );
  NAND U6958 ( .A(n6841), .B(e_input[910]), .Z(n4316) );
  NAND U6959 ( .A(n6112), .B(e_input[910]), .Z(n6841) );
  XOR U6960 ( .A(n6842), .B(n6843), .Z(n6836) );
  ANDN U6961 ( .A(n6844), .B(n4319), .Z(n6843) );
  XOR U6962 ( .A(n6845), .B(n6846), .Z(n4319) );
  IV U6963 ( .A(n6842), .Z(n6845) );
  XNOR U6964 ( .A(n4320), .B(n6842), .Z(n6844) );
  NAND U6965 ( .A(n6847), .B(e_input[909]), .Z(n4320) );
  NAND U6966 ( .A(n6112), .B(e_input[909]), .Z(n6847) );
  XOR U6967 ( .A(n6848), .B(n6849), .Z(n6842) );
  ANDN U6968 ( .A(n6850), .B(n4321), .Z(n6849) );
  XOR U6969 ( .A(n6851), .B(n6852), .Z(n4321) );
  IV U6970 ( .A(n6848), .Z(n6851) );
  XNOR U6971 ( .A(n4322), .B(n6848), .Z(n6850) );
  NAND U6972 ( .A(n6853), .B(e_input[908]), .Z(n4322) );
  NAND U6973 ( .A(n6112), .B(e_input[908]), .Z(n6853) );
  XOR U6974 ( .A(n6854), .B(n6855), .Z(n6848) );
  ANDN U6975 ( .A(n6856), .B(n4323), .Z(n6855) );
  XOR U6976 ( .A(n6857), .B(n6858), .Z(n4323) );
  IV U6977 ( .A(n6854), .Z(n6857) );
  XNOR U6978 ( .A(n4324), .B(n6854), .Z(n6856) );
  NAND U6979 ( .A(n6859), .B(e_input[907]), .Z(n4324) );
  NAND U6980 ( .A(n6112), .B(e_input[907]), .Z(n6859) );
  XOR U6981 ( .A(n6860), .B(n6861), .Z(n6854) );
  ANDN U6982 ( .A(n6862), .B(n4325), .Z(n6861) );
  XOR U6983 ( .A(n6863), .B(n6864), .Z(n4325) );
  IV U6984 ( .A(n6860), .Z(n6863) );
  XNOR U6985 ( .A(n4326), .B(n6860), .Z(n6862) );
  NAND U6986 ( .A(n6865), .B(e_input[906]), .Z(n4326) );
  NAND U6987 ( .A(n6112), .B(e_input[906]), .Z(n6865) );
  XOR U6988 ( .A(n6866), .B(n6867), .Z(n6860) );
  ANDN U6989 ( .A(n6868), .B(n4327), .Z(n6867) );
  XOR U6990 ( .A(n6869), .B(n6870), .Z(n4327) );
  IV U6991 ( .A(n6866), .Z(n6869) );
  XNOR U6992 ( .A(n4328), .B(n6866), .Z(n6868) );
  NAND U6993 ( .A(n6871), .B(e_input[905]), .Z(n4328) );
  NAND U6994 ( .A(n6112), .B(e_input[905]), .Z(n6871) );
  XOR U6995 ( .A(n6872), .B(n6873), .Z(n6866) );
  ANDN U6996 ( .A(n6874), .B(n4329), .Z(n6873) );
  XOR U6997 ( .A(n6875), .B(n6876), .Z(n4329) );
  IV U6998 ( .A(n6872), .Z(n6875) );
  XNOR U6999 ( .A(n4330), .B(n6872), .Z(n6874) );
  NAND U7000 ( .A(n6877), .B(e_input[904]), .Z(n4330) );
  NAND U7001 ( .A(n6112), .B(e_input[904]), .Z(n6877) );
  XOR U7002 ( .A(n6878), .B(n6879), .Z(n6872) );
  ANDN U7003 ( .A(n6880), .B(n4331), .Z(n6879) );
  XOR U7004 ( .A(n6881), .B(n6882), .Z(n4331) );
  IV U7005 ( .A(n6878), .Z(n6881) );
  XNOR U7006 ( .A(n4332), .B(n6878), .Z(n6880) );
  NAND U7007 ( .A(n6883), .B(e_input[903]), .Z(n4332) );
  NAND U7008 ( .A(n6112), .B(e_input[903]), .Z(n6883) );
  XOR U7009 ( .A(n6884), .B(n6885), .Z(n6878) );
  ANDN U7010 ( .A(n6886), .B(n4333), .Z(n6885) );
  XOR U7011 ( .A(n6887), .B(n6888), .Z(n4333) );
  IV U7012 ( .A(n6884), .Z(n6887) );
  XNOR U7013 ( .A(n4334), .B(n6884), .Z(n6886) );
  NAND U7014 ( .A(n6889), .B(e_input[902]), .Z(n4334) );
  NAND U7015 ( .A(n6112), .B(e_input[902]), .Z(n6889) );
  XOR U7016 ( .A(n6890), .B(n6891), .Z(n6884) );
  ANDN U7017 ( .A(n6892), .B(n4335), .Z(n6891) );
  XOR U7018 ( .A(n6893), .B(n6894), .Z(n4335) );
  IV U7019 ( .A(n6890), .Z(n6893) );
  XNOR U7020 ( .A(n4336), .B(n6890), .Z(n6892) );
  NAND U7021 ( .A(n6895), .B(e_input[901]), .Z(n4336) );
  NAND U7022 ( .A(n6112), .B(e_input[901]), .Z(n6895) );
  XOR U7023 ( .A(n6896), .B(n6897), .Z(n6890) );
  ANDN U7024 ( .A(n6898), .B(n4337), .Z(n6897) );
  XOR U7025 ( .A(n6899), .B(n6900), .Z(n4337) );
  IV U7026 ( .A(n6896), .Z(n6899) );
  XNOR U7027 ( .A(n4338), .B(n6896), .Z(n6898) );
  NAND U7028 ( .A(n6901), .B(e_input[900]), .Z(n4338) );
  NAND U7029 ( .A(n6112), .B(e_input[900]), .Z(n6901) );
  XOR U7030 ( .A(n6902), .B(n6903), .Z(n6896) );
  ANDN U7031 ( .A(n6904), .B(n4343), .Z(n6903) );
  XOR U7032 ( .A(n6905), .B(n6906), .Z(n4343) );
  IV U7033 ( .A(n6902), .Z(n6905) );
  XNOR U7034 ( .A(n4344), .B(n6902), .Z(n6904) );
  NAND U7035 ( .A(n6907), .B(e_input[899]), .Z(n4344) );
  NAND U7036 ( .A(n6112), .B(e_input[899]), .Z(n6907) );
  XOR U7037 ( .A(n6908), .B(n6909), .Z(n6902) );
  ANDN U7038 ( .A(n6910), .B(n4345), .Z(n6909) );
  XOR U7039 ( .A(n6911), .B(n6912), .Z(n4345) );
  IV U7040 ( .A(n6908), .Z(n6911) );
  XNOR U7041 ( .A(n4346), .B(n6908), .Z(n6910) );
  NAND U7042 ( .A(n6913), .B(e_input[898]), .Z(n4346) );
  NAND U7043 ( .A(n6112), .B(e_input[898]), .Z(n6913) );
  XOR U7044 ( .A(n6914), .B(n6915), .Z(n6908) );
  ANDN U7045 ( .A(n6916), .B(n4347), .Z(n6915) );
  XOR U7046 ( .A(n6917), .B(n6918), .Z(n4347) );
  IV U7047 ( .A(n6914), .Z(n6917) );
  XNOR U7048 ( .A(n4348), .B(n6914), .Z(n6916) );
  NAND U7049 ( .A(n6919), .B(e_input[897]), .Z(n4348) );
  NAND U7050 ( .A(n6112), .B(e_input[897]), .Z(n6919) );
  XOR U7051 ( .A(n6920), .B(n6921), .Z(n6914) );
  ANDN U7052 ( .A(n6922), .B(n4349), .Z(n6921) );
  XOR U7053 ( .A(n6923), .B(n6924), .Z(n4349) );
  IV U7054 ( .A(n6920), .Z(n6923) );
  XNOR U7055 ( .A(n4350), .B(n6920), .Z(n6922) );
  NAND U7056 ( .A(n6925), .B(e_input[896]), .Z(n4350) );
  NAND U7057 ( .A(n6112), .B(e_input[896]), .Z(n6925) );
  XOR U7058 ( .A(n6926), .B(n6927), .Z(n6920) );
  ANDN U7059 ( .A(n6928), .B(n4351), .Z(n6927) );
  XOR U7060 ( .A(n6929), .B(n6930), .Z(n4351) );
  IV U7061 ( .A(n6926), .Z(n6929) );
  XNOR U7062 ( .A(n4352), .B(n6926), .Z(n6928) );
  NAND U7063 ( .A(n6931), .B(e_input[895]), .Z(n4352) );
  NAND U7064 ( .A(n6112), .B(e_input[895]), .Z(n6931) );
  XOR U7065 ( .A(n6932), .B(n6933), .Z(n6926) );
  ANDN U7066 ( .A(n6934), .B(n4353), .Z(n6933) );
  XOR U7067 ( .A(n6935), .B(n6936), .Z(n4353) );
  IV U7068 ( .A(n6932), .Z(n6935) );
  XNOR U7069 ( .A(n4354), .B(n6932), .Z(n6934) );
  NAND U7070 ( .A(n6937), .B(e_input[894]), .Z(n4354) );
  NAND U7071 ( .A(n6112), .B(e_input[894]), .Z(n6937) );
  XOR U7072 ( .A(n6938), .B(n6939), .Z(n6932) );
  ANDN U7073 ( .A(n6940), .B(n4355), .Z(n6939) );
  XOR U7074 ( .A(n6941), .B(n6942), .Z(n4355) );
  IV U7075 ( .A(n6938), .Z(n6941) );
  XNOR U7076 ( .A(n4356), .B(n6938), .Z(n6940) );
  NAND U7077 ( .A(n6943), .B(e_input[893]), .Z(n4356) );
  NAND U7078 ( .A(n6112), .B(e_input[893]), .Z(n6943) );
  XOR U7079 ( .A(n6944), .B(n6945), .Z(n6938) );
  ANDN U7080 ( .A(n6946), .B(n4357), .Z(n6945) );
  XOR U7081 ( .A(n6947), .B(n6948), .Z(n4357) );
  IV U7082 ( .A(n6944), .Z(n6947) );
  XNOR U7083 ( .A(n4358), .B(n6944), .Z(n6946) );
  NAND U7084 ( .A(n6949), .B(e_input[892]), .Z(n4358) );
  NAND U7085 ( .A(n6112), .B(e_input[892]), .Z(n6949) );
  XOR U7086 ( .A(n6950), .B(n6951), .Z(n6944) );
  ANDN U7087 ( .A(n6952), .B(n4359), .Z(n6951) );
  XOR U7088 ( .A(n6953), .B(n6954), .Z(n4359) );
  IV U7089 ( .A(n6950), .Z(n6953) );
  XNOR U7090 ( .A(n4360), .B(n6950), .Z(n6952) );
  NAND U7091 ( .A(n6955), .B(e_input[891]), .Z(n4360) );
  NAND U7092 ( .A(n6112), .B(e_input[891]), .Z(n6955) );
  XOR U7093 ( .A(n6956), .B(n6957), .Z(n6950) );
  ANDN U7094 ( .A(n6958), .B(n4361), .Z(n6957) );
  XOR U7095 ( .A(n6959), .B(n6960), .Z(n4361) );
  IV U7096 ( .A(n6956), .Z(n6959) );
  XNOR U7097 ( .A(n4362), .B(n6956), .Z(n6958) );
  NAND U7098 ( .A(n6961), .B(e_input[890]), .Z(n4362) );
  NAND U7099 ( .A(n6112), .B(e_input[890]), .Z(n6961) );
  XOR U7100 ( .A(n6962), .B(n6963), .Z(n6956) );
  ANDN U7101 ( .A(n6964), .B(n4365), .Z(n6963) );
  XOR U7102 ( .A(n6965), .B(n6966), .Z(n4365) );
  IV U7103 ( .A(n6962), .Z(n6965) );
  XNOR U7104 ( .A(n4366), .B(n6962), .Z(n6964) );
  NAND U7105 ( .A(n6967), .B(e_input[889]), .Z(n4366) );
  NAND U7106 ( .A(n6112), .B(e_input[889]), .Z(n6967) );
  XOR U7107 ( .A(n6968), .B(n6969), .Z(n6962) );
  ANDN U7108 ( .A(n6970), .B(n4367), .Z(n6969) );
  XOR U7109 ( .A(n6971), .B(n6972), .Z(n4367) );
  IV U7110 ( .A(n6968), .Z(n6971) );
  XNOR U7111 ( .A(n4368), .B(n6968), .Z(n6970) );
  NAND U7112 ( .A(n6973), .B(e_input[888]), .Z(n4368) );
  NAND U7113 ( .A(n6112), .B(e_input[888]), .Z(n6973) );
  XOR U7114 ( .A(n6974), .B(n6975), .Z(n6968) );
  ANDN U7115 ( .A(n6976), .B(n4369), .Z(n6975) );
  XOR U7116 ( .A(n6977), .B(n6978), .Z(n4369) );
  IV U7117 ( .A(n6974), .Z(n6977) );
  XNOR U7118 ( .A(n4370), .B(n6974), .Z(n6976) );
  NAND U7119 ( .A(n6979), .B(e_input[887]), .Z(n4370) );
  NAND U7120 ( .A(n6112), .B(e_input[887]), .Z(n6979) );
  XOR U7121 ( .A(n6980), .B(n6981), .Z(n6974) );
  ANDN U7122 ( .A(n6982), .B(n4371), .Z(n6981) );
  XOR U7123 ( .A(n6983), .B(n6984), .Z(n4371) );
  IV U7124 ( .A(n6980), .Z(n6983) );
  XNOR U7125 ( .A(n4372), .B(n6980), .Z(n6982) );
  NAND U7126 ( .A(n6985), .B(e_input[886]), .Z(n4372) );
  NAND U7127 ( .A(n6112), .B(e_input[886]), .Z(n6985) );
  XOR U7128 ( .A(n6986), .B(n6987), .Z(n6980) );
  ANDN U7129 ( .A(n6988), .B(n4373), .Z(n6987) );
  XOR U7130 ( .A(n6989), .B(n6990), .Z(n4373) );
  IV U7131 ( .A(n6986), .Z(n6989) );
  XNOR U7132 ( .A(n4374), .B(n6986), .Z(n6988) );
  NAND U7133 ( .A(n6991), .B(e_input[885]), .Z(n4374) );
  NAND U7134 ( .A(n6112), .B(e_input[885]), .Z(n6991) );
  XOR U7135 ( .A(n6992), .B(n6993), .Z(n6986) );
  ANDN U7136 ( .A(n6994), .B(n4375), .Z(n6993) );
  XOR U7137 ( .A(n6995), .B(n6996), .Z(n4375) );
  IV U7138 ( .A(n6992), .Z(n6995) );
  XNOR U7139 ( .A(n4376), .B(n6992), .Z(n6994) );
  NAND U7140 ( .A(n6997), .B(e_input[884]), .Z(n4376) );
  NAND U7141 ( .A(n6112), .B(e_input[884]), .Z(n6997) );
  XOR U7142 ( .A(n6998), .B(n6999), .Z(n6992) );
  ANDN U7143 ( .A(n7000), .B(n4377), .Z(n6999) );
  XOR U7144 ( .A(n7001), .B(n7002), .Z(n4377) );
  IV U7145 ( .A(n6998), .Z(n7001) );
  XNOR U7146 ( .A(n4378), .B(n6998), .Z(n7000) );
  NAND U7147 ( .A(n7003), .B(e_input[883]), .Z(n4378) );
  NAND U7148 ( .A(n6112), .B(e_input[883]), .Z(n7003) );
  XOR U7149 ( .A(n7004), .B(n7005), .Z(n6998) );
  ANDN U7150 ( .A(n7006), .B(n4379), .Z(n7005) );
  XOR U7151 ( .A(n7007), .B(n7008), .Z(n4379) );
  IV U7152 ( .A(n7004), .Z(n7007) );
  XNOR U7153 ( .A(n4380), .B(n7004), .Z(n7006) );
  NAND U7154 ( .A(n7009), .B(e_input[882]), .Z(n4380) );
  NAND U7155 ( .A(n6112), .B(e_input[882]), .Z(n7009) );
  XOR U7156 ( .A(n7010), .B(n7011), .Z(n7004) );
  ANDN U7157 ( .A(n7012), .B(n4381), .Z(n7011) );
  XOR U7158 ( .A(n7013), .B(n7014), .Z(n4381) );
  IV U7159 ( .A(n7010), .Z(n7013) );
  XNOR U7160 ( .A(n4382), .B(n7010), .Z(n7012) );
  NAND U7161 ( .A(n7015), .B(e_input[881]), .Z(n4382) );
  NAND U7162 ( .A(n6112), .B(e_input[881]), .Z(n7015) );
  XOR U7163 ( .A(n7016), .B(n7017), .Z(n7010) );
  ANDN U7164 ( .A(n7018), .B(n4383), .Z(n7017) );
  XOR U7165 ( .A(n7019), .B(n7020), .Z(n4383) );
  IV U7166 ( .A(n7016), .Z(n7019) );
  XNOR U7167 ( .A(n4384), .B(n7016), .Z(n7018) );
  NAND U7168 ( .A(n7021), .B(e_input[880]), .Z(n4384) );
  NAND U7169 ( .A(n6112), .B(e_input[880]), .Z(n7021) );
  XOR U7170 ( .A(n7022), .B(n7023), .Z(n7016) );
  ANDN U7171 ( .A(n7024), .B(n4387), .Z(n7023) );
  XOR U7172 ( .A(n7025), .B(n7026), .Z(n4387) );
  IV U7173 ( .A(n7022), .Z(n7025) );
  XNOR U7174 ( .A(n4388), .B(n7022), .Z(n7024) );
  NAND U7175 ( .A(n7027), .B(e_input[879]), .Z(n4388) );
  NAND U7176 ( .A(n6112), .B(e_input[879]), .Z(n7027) );
  XOR U7177 ( .A(n7028), .B(n7029), .Z(n7022) );
  ANDN U7178 ( .A(n7030), .B(n4389), .Z(n7029) );
  XOR U7179 ( .A(n7031), .B(n7032), .Z(n4389) );
  IV U7180 ( .A(n7028), .Z(n7031) );
  XNOR U7181 ( .A(n4390), .B(n7028), .Z(n7030) );
  NAND U7182 ( .A(n7033), .B(e_input[878]), .Z(n4390) );
  NAND U7183 ( .A(n6112), .B(e_input[878]), .Z(n7033) );
  XOR U7184 ( .A(n7034), .B(n7035), .Z(n7028) );
  ANDN U7185 ( .A(n7036), .B(n4391), .Z(n7035) );
  XOR U7186 ( .A(n7037), .B(n7038), .Z(n4391) );
  IV U7187 ( .A(n7034), .Z(n7037) );
  XNOR U7188 ( .A(n4392), .B(n7034), .Z(n7036) );
  NAND U7189 ( .A(n7039), .B(e_input[877]), .Z(n4392) );
  NAND U7190 ( .A(n6112), .B(e_input[877]), .Z(n7039) );
  XOR U7191 ( .A(n7040), .B(n7041), .Z(n7034) );
  ANDN U7192 ( .A(n7042), .B(n4393), .Z(n7041) );
  XOR U7193 ( .A(n7043), .B(n7044), .Z(n4393) );
  IV U7194 ( .A(n7040), .Z(n7043) );
  XNOR U7195 ( .A(n4394), .B(n7040), .Z(n7042) );
  NAND U7196 ( .A(n7045), .B(e_input[876]), .Z(n4394) );
  NAND U7197 ( .A(n6112), .B(e_input[876]), .Z(n7045) );
  XOR U7198 ( .A(n7046), .B(n7047), .Z(n7040) );
  ANDN U7199 ( .A(n7048), .B(n4395), .Z(n7047) );
  XOR U7200 ( .A(n7049), .B(n7050), .Z(n4395) );
  IV U7201 ( .A(n7046), .Z(n7049) );
  XNOR U7202 ( .A(n4396), .B(n7046), .Z(n7048) );
  NAND U7203 ( .A(n7051), .B(e_input[875]), .Z(n4396) );
  NAND U7204 ( .A(n6112), .B(e_input[875]), .Z(n7051) );
  XOR U7205 ( .A(n7052), .B(n7053), .Z(n7046) );
  ANDN U7206 ( .A(n7054), .B(n4397), .Z(n7053) );
  XOR U7207 ( .A(n7055), .B(n7056), .Z(n4397) );
  IV U7208 ( .A(n7052), .Z(n7055) );
  XNOR U7209 ( .A(n4398), .B(n7052), .Z(n7054) );
  NAND U7210 ( .A(n7057), .B(e_input[874]), .Z(n4398) );
  NAND U7211 ( .A(n6112), .B(e_input[874]), .Z(n7057) );
  XOR U7212 ( .A(n7058), .B(n7059), .Z(n7052) );
  ANDN U7213 ( .A(n7060), .B(n4399), .Z(n7059) );
  XOR U7214 ( .A(n7061), .B(n7062), .Z(n4399) );
  IV U7215 ( .A(n7058), .Z(n7061) );
  XNOR U7216 ( .A(n4400), .B(n7058), .Z(n7060) );
  NAND U7217 ( .A(n7063), .B(e_input[873]), .Z(n4400) );
  NAND U7218 ( .A(n6112), .B(e_input[873]), .Z(n7063) );
  XOR U7219 ( .A(n7064), .B(n7065), .Z(n7058) );
  ANDN U7220 ( .A(n7066), .B(n4401), .Z(n7065) );
  XOR U7221 ( .A(n7067), .B(n7068), .Z(n4401) );
  IV U7222 ( .A(n7064), .Z(n7067) );
  XNOR U7223 ( .A(n4402), .B(n7064), .Z(n7066) );
  NAND U7224 ( .A(n7069), .B(e_input[872]), .Z(n4402) );
  NAND U7225 ( .A(n6112), .B(e_input[872]), .Z(n7069) );
  XOR U7226 ( .A(n7070), .B(n7071), .Z(n7064) );
  ANDN U7227 ( .A(n7072), .B(n4403), .Z(n7071) );
  XOR U7228 ( .A(n7073), .B(n7074), .Z(n4403) );
  IV U7229 ( .A(n7070), .Z(n7073) );
  XNOR U7230 ( .A(n4404), .B(n7070), .Z(n7072) );
  NAND U7231 ( .A(n7075), .B(e_input[871]), .Z(n4404) );
  NAND U7232 ( .A(n6112), .B(e_input[871]), .Z(n7075) );
  XOR U7233 ( .A(n7076), .B(n7077), .Z(n7070) );
  ANDN U7234 ( .A(n7078), .B(n4405), .Z(n7077) );
  XOR U7235 ( .A(n7079), .B(n7080), .Z(n4405) );
  IV U7236 ( .A(n7076), .Z(n7079) );
  XNOR U7237 ( .A(n4406), .B(n7076), .Z(n7078) );
  NAND U7238 ( .A(n7081), .B(e_input[870]), .Z(n4406) );
  NAND U7239 ( .A(n6112), .B(e_input[870]), .Z(n7081) );
  XOR U7240 ( .A(n7082), .B(n7083), .Z(n7076) );
  ANDN U7241 ( .A(n7084), .B(n4409), .Z(n7083) );
  XOR U7242 ( .A(n7085), .B(n7086), .Z(n4409) );
  IV U7243 ( .A(n7082), .Z(n7085) );
  XNOR U7244 ( .A(n4410), .B(n7082), .Z(n7084) );
  NAND U7245 ( .A(n7087), .B(e_input[869]), .Z(n4410) );
  NAND U7246 ( .A(n6112), .B(e_input[869]), .Z(n7087) );
  XOR U7247 ( .A(n7088), .B(n7089), .Z(n7082) );
  ANDN U7248 ( .A(n7090), .B(n4411), .Z(n7089) );
  XOR U7249 ( .A(n7091), .B(n7092), .Z(n4411) );
  IV U7250 ( .A(n7088), .Z(n7091) );
  XNOR U7251 ( .A(n4412), .B(n7088), .Z(n7090) );
  NAND U7252 ( .A(n7093), .B(e_input[868]), .Z(n4412) );
  NAND U7253 ( .A(n6112), .B(e_input[868]), .Z(n7093) );
  XOR U7254 ( .A(n7094), .B(n7095), .Z(n7088) );
  ANDN U7255 ( .A(n7096), .B(n4413), .Z(n7095) );
  XOR U7256 ( .A(n7097), .B(n7098), .Z(n4413) );
  IV U7257 ( .A(n7094), .Z(n7097) );
  XNOR U7258 ( .A(n4414), .B(n7094), .Z(n7096) );
  NAND U7259 ( .A(n7099), .B(e_input[867]), .Z(n4414) );
  NAND U7260 ( .A(n6112), .B(e_input[867]), .Z(n7099) );
  XOR U7261 ( .A(n7100), .B(n7101), .Z(n7094) );
  ANDN U7262 ( .A(n7102), .B(n4415), .Z(n7101) );
  XOR U7263 ( .A(n7103), .B(n7104), .Z(n4415) );
  IV U7264 ( .A(n7100), .Z(n7103) );
  XNOR U7265 ( .A(n4416), .B(n7100), .Z(n7102) );
  NAND U7266 ( .A(n7105), .B(e_input[866]), .Z(n4416) );
  NAND U7267 ( .A(n6112), .B(e_input[866]), .Z(n7105) );
  XOR U7268 ( .A(n7106), .B(n7107), .Z(n7100) );
  ANDN U7269 ( .A(n7108), .B(n4417), .Z(n7107) );
  XOR U7270 ( .A(n7109), .B(n7110), .Z(n4417) );
  IV U7271 ( .A(n7106), .Z(n7109) );
  XNOR U7272 ( .A(n4418), .B(n7106), .Z(n7108) );
  NAND U7273 ( .A(n7111), .B(e_input[865]), .Z(n4418) );
  NAND U7274 ( .A(n6112), .B(e_input[865]), .Z(n7111) );
  XOR U7275 ( .A(n7112), .B(n7113), .Z(n7106) );
  ANDN U7276 ( .A(n7114), .B(n4419), .Z(n7113) );
  XOR U7277 ( .A(n7115), .B(n7116), .Z(n4419) );
  IV U7278 ( .A(n7112), .Z(n7115) );
  XNOR U7279 ( .A(n4420), .B(n7112), .Z(n7114) );
  NAND U7280 ( .A(n7117), .B(e_input[864]), .Z(n4420) );
  NAND U7281 ( .A(n6112), .B(e_input[864]), .Z(n7117) );
  XOR U7282 ( .A(n7118), .B(n7119), .Z(n7112) );
  ANDN U7283 ( .A(n7120), .B(n4421), .Z(n7119) );
  XOR U7284 ( .A(n7121), .B(n7122), .Z(n4421) );
  IV U7285 ( .A(n7118), .Z(n7121) );
  XNOR U7286 ( .A(n4422), .B(n7118), .Z(n7120) );
  NAND U7287 ( .A(n7123), .B(e_input[863]), .Z(n4422) );
  NAND U7288 ( .A(n6112), .B(e_input[863]), .Z(n7123) );
  XOR U7289 ( .A(n7124), .B(n7125), .Z(n7118) );
  ANDN U7290 ( .A(n7126), .B(n4423), .Z(n7125) );
  XOR U7291 ( .A(n7127), .B(n7128), .Z(n4423) );
  IV U7292 ( .A(n7124), .Z(n7127) );
  XNOR U7293 ( .A(n4424), .B(n7124), .Z(n7126) );
  NAND U7294 ( .A(n7129), .B(e_input[862]), .Z(n4424) );
  NAND U7295 ( .A(n6112), .B(e_input[862]), .Z(n7129) );
  XOR U7296 ( .A(n7130), .B(n7131), .Z(n7124) );
  ANDN U7297 ( .A(n7132), .B(n4425), .Z(n7131) );
  XOR U7298 ( .A(n7133), .B(n7134), .Z(n4425) );
  IV U7299 ( .A(n7130), .Z(n7133) );
  XNOR U7300 ( .A(n4426), .B(n7130), .Z(n7132) );
  NAND U7301 ( .A(n7135), .B(e_input[861]), .Z(n4426) );
  NAND U7302 ( .A(n6112), .B(e_input[861]), .Z(n7135) );
  XOR U7303 ( .A(n7136), .B(n7137), .Z(n7130) );
  ANDN U7304 ( .A(n7138), .B(n4427), .Z(n7137) );
  XOR U7305 ( .A(n7139), .B(n7140), .Z(n4427) );
  IV U7306 ( .A(n7136), .Z(n7139) );
  XNOR U7307 ( .A(n4428), .B(n7136), .Z(n7138) );
  NAND U7308 ( .A(n7141), .B(e_input[860]), .Z(n4428) );
  NAND U7309 ( .A(n6112), .B(e_input[860]), .Z(n7141) );
  XOR U7310 ( .A(n7142), .B(n7143), .Z(n7136) );
  ANDN U7311 ( .A(n7144), .B(n4431), .Z(n7143) );
  XOR U7312 ( .A(n7145), .B(n7146), .Z(n4431) );
  IV U7313 ( .A(n7142), .Z(n7145) );
  XNOR U7314 ( .A(n4432), .B(n7142), .Z(n7144) );
  NAND U7315 ( .A(n7147), .B(e_input[859]), .Z(n4432) );
  NAND U7316 ( .A(n6112), .B(e_input[859]), .Z(n7147) );
  XOR U7317 ( .A(n7148), .B(n7149), .Z(n7142) );
  ANDN U7318 ( .A(n7150), .B(n4433), .Z(n7149) );
  XOR U7319 ( .A(n7151), .B(n7152), .Z(n4433) );
  IV U7320 ( .A(n7148), .Z(n7151) );
  XNOR U7321 ( .A(n4434), .B(n7148), .Z(n7150) );
  NAND U7322 ( .A(n7153), .B(e_input[858]), .Z(n4434) );
  NAND U7323 ( .A(n6112), .B(e_input[858]), .Z(n7153) );
  XOR U7324 ( .A(n7154), .B(n7155), .Z(n7148) );
  ANDN U7325 ( .A(n7156), .B(n4435), .Z(n7155) );
  XOR U7326 ( .A(n7157), .B(n7158), .Z(n4435) );
  IV U7327 ( .A(n7154), .Z(n7157) );
  XNOR U7328 ( .A(n4436), .B(n7154), .Z(n7156) );
  NAND U7329 ( .A(n7159), .B(e_input[857]), .Z(n4436) );
  NAND U7330 ( .A(n6112), .B(e_input[857]), .Z(n7159) );
  XOR U7331 ( .A(n7160), .B(n7161), .Z(n7154) );
  ANDN U7332 ( .A(n7162), .B(n4437), .Z(n7161) );
  XOR U7333 ( .A(n7163), .B(n7164), .Z(n4437) );
  IV U7334 ( .A(n7160), .Z(n7163) );
  XNOR U7335 ( .A(n4438), .B(n7160), .Z(n7162) );
  NAND U7336 ( .A(n7165), .B(e_input[856]), .Z(n4438) );
  NAND U7337 ( .A(n6112), .B(e_input[856]), .Z(n7165) );
  XOR U7338 ( .A(n7166), .B(n7167), .Z(n7160) );
  ANDN U7339 ( .A(n7168), .B(n4439), .Z(n7167) );
  XOR U7340 ( .A(n7169), .B(n7170), .Z(n4439) );
  IV U7341 ( .A(n7166), .Z(n7169) );
  XNOR U7342 ( .A(n4440), .B(n7166), .Z(n7168) );
  NAND U7343 ( .A(n7171), .B(e_input[855]), .Z(n4440) );
  NAND U7344 ( .A(n6112), .B(e_input[855]), .Z(n7171) );
  XOR U7345 ( .A(n7172), .B(n7173), .Z(n7166) );
  ANDN U7346 ( .A(n7174), .B(n4441), .Z(n7173) );
  XOR U7347 ( .A(n7175), .B(n7176), .Z(n4441) );
  IV U7348 ( .A(n7172), .Z(n7175) );
  XNOR U7349 ( .A(n4442), .B(n7172), .Z(n7174) );
  NAND U7350 ( .A(n7177), .B(e_input[854]), .Z(n4442) );
  NAND U7351 ( .A(n6112), .B(e_input[854]), .Z(n7177) );
  XOR U7352 ( .A(n7178), .B(n7179), .Z(n7172) );
  ANDN U7353 ( .A(n7180), .B(n4443), .Z(n7179) );
  XOR U7354 ( .A(n7181), .B(n7182), .Z(n4443) );
  IV U7355 ( .A(n7178), .Z(n7181) );
  XNOR U7356 ( .A(n4444), .B(n7178), .Z(n7180) );
  NAND U7357 ( .A(n7183), .B(e_input[853]), .Z(n4444) );
  NAND U7358 ( .A(n6112), .B(e_input[853]), .Z(n7183) );
  XOR U7359 ( .A(n7184), .B(n7185), .Z(n7178) );
  ANDN U7360 ( .A(n7186), .B(n4445), .Z(n7185) );
  XOR U7361 ( .A(n7187), .B(n7188), .Z(n4445) );
  IV U7362 ( .A(n7184), .Z(n7187) );
  XNOR U7363 ( .A(n4446), .B(n7184), .Z(n7186) );
  NAND U7364 ( .A(n7189), .B(e_input[852]), .Z(n4446) );
  NAND U7365 ( .A(n6112), .B(e_input[852]), .Z(n7189) );
  XOR U7366 ( .A(n7190), .B(n7191), .Z(n7184) );
  ANDN U7367 ( .A(n7192), .B(n4447), .Z(n7191) );
  XOR U7368 ( .A(n7193), .B(n7194), .Z(n4447) );
  IV U7369 ( .A(n7190), .Z(n7193) );
  XNOR U7370 ( .A(n4448), .B(n7190), .Z(n7192) );
  NAND U7371 ( .A(n7195), .B(e_input[851]), .Z(n4448) );
  NAND U7372 ( .A(n6112), .B(e_input[851]), .Z(n7195) );
  XOR U7373 ( .A(n7196), .B(n7197), .Z(n7190) );
  ANDN U7374 ( .A(n7198), .B(n4449), .Z(n7197) );
  XOR U7375 ( .A(n7199), .B(n7200), .Z(n4449) );
  IV U7376 ( .A(n7196), .Z(n7199) );
  XNOR U7377 ( .A(n4450), .B(n7196), .Z(n7198) );
  NAND U7378 ( .A(n7201), .B(e_input[850]), .Z(n4450) );
  NAND U7379 ( .A(n6112), .B(e_input[850]), .Z(n7201) );
  XOR U7380 ( .A(n7202), .B(n7203), .Z(n7196) );
  ANDN U7381 ( .A(n7204), .B(n4453), .Z(n7203) );
  XOR U7382 ( .A(n7205), .B(n7206), .Z(n4453) );
  IV U7383 ( .A(n7202), .Z(n7205) );
  XNOR U7384 ( .A(n4454), .B(n7202), .Z(n7204) );
  NAND U7385 ( .A(n7207), .B(e_input[849]), .Z(n4454) );
  NAND U7386 ( .A(n6112), .B(e_input[849]), .Z(n7207) );
  XOR U7387 ( .A(n7208), .B(n7209), .Z(n7202) );
  ANDN U7388 ( .A(n7210), .B(n4455), .Z(n7209) );
  XOR U7389 ( .A(n7211), .B(n7212), .Z(n4455) );
  IV U7390 ( .A(n7208), .Z(n7211) );
  XNOR U7391 ( .A(n4456), .B(n7208), .Z(n7210) );
  NAND U7392 ( .A(n7213), .B(e_input[848]), .Z(n4456) );
  NAND U7393 ( .A(n6112), .B(e_input[848]), .Z(n7213) );
  XOR U7394 ( .A(n7214), .B(n7215), .Z(n7208) );
  ANDN U7395 ( .A(n7216), .B(n4457), .Z(n7215) );
  XOR U7396 ( .A(n7217), .B(n7218), .Z(n4457) );
  IV U7397 ( .A(n7214), .Z(n7217) );
  XNOR U7398 ( .A(n4458), .B(n7214), .Z(n7216) );
  NAND U7399 ( .A(n7219), .B(e_input[847]), .Z(n4458) );
  NAND U7400 ( .A(n6112), .B(e_input[847]), .Z(n7219) );
  XOR U7401 ( .A(n7220), .B(n7221), .Z(n7214) );
  ANDN U7402 ( .A(n7222), .B(n4459), .Z(n7221) );
  XOR U7403 ( .A(n7223), .B(n7224), .Z(n4459) );
  IV U7404 ( .A(n7220), .Z(n7223) );
  XNOR U7405 ( .A(n4460), .B(n7220), .Z(n7222) );
  NAND U7406 ( .A(n7225), .B(e_input[846]), .Z(n4460) );
  NAND U7407 ( .A(n6112), .B(e_input[846]), .Z(n7225) );
  XOR U7408 ( .A(n7226), .B(n7227), .Z(n7220) );
  ANDN U7409 ( .A(n7228), .B(n4461), .Z(n7227) );
  XOR U7410 ( .A(n7229), .B(n7230), .Z(n4461) );
  IV U7411 ( .A(n7226), .Z(n7229) );
  XNOR U7412 ( .A(n4462), .B(n7226), .Z(n7228) );
  NAND U7413 ( .A(n7231), .B(e_input[845]), .Z(n4462) );
  NAND U7414 ( .A(n6112), .B(e_input[845]), .Z(n7231) );
  XOR U7415 ( .A(n7232), .B(n7233), .Z(n7226) );
  ANDN U7416 ( .A(n7234), .B(n4463), .Z(n7233) );
  XOR U7417 ( .A(n7235), .B(n7236), .Z(n4463) );
  IV U7418 ( .A(n7232), .Z(n7235) );
  XNOR U7419 ( .A(n4464), .B(n7232), .Z(n7234) );
  NAND U7420 ( .A(n7237), .B(e_input[844]), .Z(n4464) );
  NAND U7421 ( .A(n6112), .B(e_input[844]), .Z(n7237) );
  XOR U7422 ( .A(n7238), .B(n7239), .Z(n7232) );
  ANDN U7423 ( .A(n7240), .B(n4465), .Z(n7239) );
  XOR U7424 ( .A(n7241), .B(n7242), .Z(n4465) );
  IV U7425 ( .A(n7238), .Z(n7241) );
  XNOR U7426 ( .A(n4466), .B(n7238), .Z(n7240) );
  NAND U7427 ( .A(n7243), .B(e_input[843]), .Z(n4466) );
  NAND U7428 ( .A(n6112), .B(e_input[843]), .Z(n7243) );
  XOR U7429 ( .A(n7244), .B(n7245), .Z(n7238) );
  ANDN U7430 ( .A(n7246), .B(n4467), .Z(n7245) );
  XOR U7431 ( .A(n7247), .B(n7248), .Z(n4467) );
  IV U7432 ( .A(n7244), .Z(n7247) );
  XNOR U7433 ( .A(n4468), .B(n7244), .Z(n7246) );
  NAND U7434 ( .A(n7249), .B(e_input[842]), .Z(n4468) );
  NAND U7435 ( .A(n6112), .B(e_input[842]), .Z(n7249) );
  XOR U7436 ( .A(n7250), .B(n7251), .Z(n7244) );
  ANDN U7437 ( .A(n7252), .B(n4469), .Z(n7251) );
  XOR U7438 ( .A(n7253), .B(n7254), .Z(n4469) );
  IV U7439 ( .A(n7250), .Z(n7253) );
  XNOR U7440 ( .A(n4470), .B(n7250), .Z(n7252) );
  NAND U7441 ( .A(n7255), .B(e_input[841]), .Z(n4470) );
  NAND U7442 ( .A(n6112), .B(e_input[841]), .Z(n7255) );
  XOR U7443 ( .A(n7256), .B(n7257), .Z(n7250) );
  ANDN U7444 ( .A(n7258), .B(n4471), .Z(n7257) );
  XOR U7445 ( .A(n7259), .B(n7260), .Z(n4471) );
  IV U7446 ( .A(n7256), .Z(n7259) );
  XNOR U7447 ( .A(n4472), .B(n7256), .Z(n7258) );
  NAND U7448 ( .A(n7261), .B(e_input[840]), .Z(n4472) );
  NAND U7449 ( .A(n6112), .B(e_input[840]), .Z(n7261) );
  XOR U7450 ( .A(n7262), .B(n7263), .Z(n7256) );
  ANDN U7451 ( .A(n7264), .B(n4475), .Z(n7263) );
  XOR U7452 ( .A(n7265), .B(n7266), .Z(n4475) );
  IV U7453 ( .A(n7262), .Z(n7265) );
  XNOR U7454 ( .A(n4476), .B(n7262), .Z(n7264) );
  NAND U7455 ( .A(n7267), .B(e_input[839]), .Z(n4476) );
  NAND U7456 ( .A(n6112), .B(e_input[839]), .Z(n7267) );
  XOR U7457 ( .A(n7268), .B(n7269), .Z(n7262) );
  ANDN U7458 ( .A(n7270), .B(n4477), .Z(n7269) );
  XOR U7459 ( .A(n7271), .B(n7272), .Z(n4477) );
  IV U7460 ( .A(n7268), .Z(n7271) );
  XNOR U7461 ( .A(n4478), .B(n7268), .Z(n7270) );
  NAND U7462 ( .A(n7273), .B(e_input[838]), .Z(n4478) );
  NAND U7463 ( .A(n6112), .B(e_input[838]), .Z(n7273) );
  XOR U7464 ( .A(n7274), .B(n7275), .Z(n7268) );
  ANDN U7465 ( .A(n7276), .B(n4479), .Z(n7275) );
  XOR U7466 ( .A(n7277), .B(n7278), .Z(n4479) );
  IV U7467 ( .A(n7274), .Z(n7277) );
  XNOR U7468 ( .A(n4480), .B(n7274), .Z(n7276) );
  NAND U7469 ( .A(n7279), .B(e_input[837]), .Z(n4480) );
  NAND U7470 ( .A(n6112), .B(e_input[837]), .Z(n7279) );
  XOR U7471 ( .A(n7280), .B(n7281), .Z(n7274) );
  ANDN U7472 ( .A(n7282), .B(n4481), .Z(n7281) );
  XOR U7473 ( .A(n7283), .B(n7284), .Z(n4481) );
  IV U7474 ( .A(n7280), .Z(n7283) );
  XNOR U7475 ( .A(n4482), .B(n7280), .Z(n7282) );
  NAND U7476 ( .A(n7285), .B(e_input[836]), .Z(n4482) );
  NAND U7477 ( .A(n6112), .B(e_input[836]), .Z(n7285) );
  XOR U7478 ( .A(n7286), .B(n7287), .Z(n7280) );
  ANDN U7479 ( .A(n7288), .B(n4483), .Z(n7287) );
  XOR U7480 ( .A(n7289), .B(n7290), .Z(n4483) );
  IV U7481 ( .A(n7286), .Z(n7289) );
  XNOR U7482 ( .A(n4484), .B(n7286), .Z(n7288) );
  NAND U7483 ( .A(n7291), .B(e_input[835]), .Z(n4484) );
  NAND U7484 ( .A(n6112), .B(e_input[835]), .Z(n7291) );
  XOR U7485 ( .A(n7292), .B(n7293), .Z(n7286) );
  ANDN U7486 ( .A(n7294), .B(n4485), .Z(n7293) );
  XOR U7487 ( .A(n7295), .B(n7296), .Z(n4485) );
  IV U7488 ( .A(n7292), .Z(n7295) );
  XNOR U7489 ( .A(n4486), .B(n7292), .Z(n7294) );
  NAND U7490 ( .A(n7297), .B(e_input[834]), .Z(n4486) );
  NAND U7491 ( .A(n6112), .B(e_input[834]), .Z(n7297) );
  XOR U7492 ( .A(n7298), .B(n7299), .Z(n7292) );
  ANDN U7493 ( .A(n7300), .B(n4487), .Z(n7299) );
  XOR U7494 ( .A(n7301), .B(n7302), .Z(n4487) );
  IV U7495 ( .A(n7298), .Z(n7301) );
  XNOR U7496 ( .A(n4488), .B(n7298), .Z(n7300) );
  NAND U7497 ( .A(n7303), .B(e_input[833]), .Z(n4488) );
  NAND U7498 ( .A(n6112), .B(e_input[833]), .Z(n7303) );
  XOR U7499 ( .A(n7304), .B(n7305), .Z(n7298) );
  ANDN U7500 ( .A(n7306), .B(n4489), .Z(n7305) );
  XOR U7501 ( .A(n7307), .B(n7308), .Z(n4489) );
  IV U7502 ( .A(n7304), .Z(n7307) );
  XNOR U7503 ( .A(n4490), .B(n7304), .Z(n7306) );
  NAND U7504 ( .A(n7309), .B(e_input[832]), .Z(n4490) );
  NAND U7505 ( .A(n6112), .B(e_input[832]), .Z(n7309) );
  XOR U7506 ( .A(n7310), .B(n7311), .Z(n7304) );
  ANDN U7507 ( .A(n7312), .B(n4491), .Z(n7311) );
  XOR U7508 ( .A(n7313), .B(n7314), .Z(n4491) );
  IV U7509 ( .A(n7310), .Z(n7313) );
  XNOR U7510 ( .A(n4492), .B(n7310), .Z(n7312) );
  NAND U7511 ( .A(n7315), .B(e_input[831]), .Z(n4492) );
  NAND U7512 ( .A(n6112), .B(e_input[831]), .Z(n7315) );
  XOR U7513 ( .A(n7316), .B(n7317), .Z(n7310) );
  ANDN U7514 ( .A(n7318), .B(n4493), .Z(n7317) );
  XOR U7515 ( .A(n7319), .B(n7320), .Z(n4493) );
  IV U7516 ( .A(n7316), .Z(n7319) );
  XNOR U7517 ( .A(n4494), .B(n7316), .Z(n7318) );
  NAND U7518 ( .A(n7321), .B(e_input[830]), .Z(n4494) );
  NAND U7519 ( .A(n6112), .B(e_input[830]), .Z(n7321) );
  XOR U7520 ( .A(n7322), .B(n7323), .Z(n7316) );
  ANDN U7521 ( .A(n7324), .B(n4497), .Z(n7323) );
  XOR U7522 ( .A(n7325), .B(n7326), .Z(n4497) );
  IV U7523 ( .A(n7322), .Z(n7325) );
  XNOR U7524 ( .A(n4498), .B(n7322), .Z(n7324) );
  NAND U7525 ( .A(n7327), .B(e_input[829]), .Z(n4498) );
  NAND U7526 ( .A(n6112), .B(e_input[829]), .Z(n7327) );
  XOR U7527 ( .A(n7328), .B(n7329), .Z(n7322) );
  ANDN U7528 ( .A(n7330), .B(n4499), .Z(n7329) );
  XOR U7529 ( .A(n7331), .B(n7332), .Z(n4499) );
  IV U7530 ( .A(n7328), .Z(n7331) );
  XNOR U7531 ( .A(n4500), .B(n7328), .Z(n7330) );
  NAND U7532 ( .A(n7333), .B(e_input[828]), .Z(n4500) );
  NAND U7533 ( .A(n6112), .B(e_input[828]), .Z(n7333) );
  XOR U7534 ( .A(n7334), .B(n7335), .Z(n7328) );
  ANDN U7535 ( .A(n7336), .B(n4501), .Z(n7335) );
  XOR U7536 ( .A(n7337), .B(n7338), .Z(n4501) );
  IV U7537 ( .A(n7334), .Z(n7337) );
  XNOR U7538 ( .A(n4502), .B(n7334), .Z(n7336) );
  NAND U7539 ( .A(n7339), .B(e_input[827]), .Z(n4502) );
  NAND U7540 ( .A(n6112), .B(e_input[827]), .Z(n7339) );
  XOR U7541 ( .A(n7340), .B(n7341), .Z(n7334) );
  ANDN U7542 ( .A(n7342), .B(n4503), .Z(n7341) );
  XOR U7543 ( .A(n7343), .B(n7344), .Z(n4503) );
  IV U7544 ( .A(n7340), .Z(n7343) );
  XNOR U7545 ( .A(n4504), .B(n7340), .Z(n7342) );
  NAND U7546 ( .A(n7345), .B(e_input[826]), .Z(n4504) );
  NAND U7547 ( .A(n6112), .B(e_input[826]), .Z(n7345) );
  XOR U7548 ( .A(n7346), .B(n7347), .Z(n7340) );
  ANDN U7549 ( .A(n7348), .B(n4505), .Z(n7347) );
  XOR U7550 ( .A(n7349), .B(n7350), .Z(n4505) );
  IV U7551 ( .A(n7346), .Z(n7349) );
  XNOR U7552 ( .A(n4506), .B(n7346), .Z(n7348) );
  NAND U7553 ( .A(n7351), .B(e_input[825]), .Z(n4506) );
  NAND U7554 ( .A(n6112), .B(e_input[825]), .Z(n7351) );
  XOR U7555 ( .A(n7352), .B(n7353), .Z(n7346) );
  ANDN U7556 ( .A(n7354), .B(n4507), .Z(n7353) );
  XOR U7557 ( .A(n7355), .B(n7356), .Z(n4507) );
  IV U7558 ( .A(n7352), .Z(n7355) );
  XNOR U7559 ( .A(n4508), .B(n7352), .Z(n7354) );
  NAND U7560 ( .A(n7357), .B(e_input[824]), .Z(n4508) );
  NAND U7561 ( .A(n6112), .B(e_input[824]), .Z(n7357) );
  XOR U7562 ( .A(n7358), .B(n7359), .Z(n7352) );
  ANDN U7563 ( .A(n7360), .B(n4509), .Z(n7359) );
  XOR U7564 ( .A(n7361), .B(n7362), .Z(n4509) );
  IV U7565 ( .A(n7358), .Z(n7361) );
  XNOR U7566 ( .A(n4510), .B(n7358), .Z(n7360) );
  NAND U7567 ( .A(n7363), .B(e_input[823]), .Z(n4510) );
  NAND U7568 ( .A(n6112), .B(e_input[823]), .Z(n7363) );
  XOR U7569 ( .A(n7364), .B(n7365), .Z(n7358) );
  ANDN U7570 ( .A(n7366), .B(n4511), .Z(n7365) );
  XOR U7571 ( .A(n7367), .B(n7368), .Z(n4511) );
  IV U7572 ( .A(n7364), .Z(n7367) );
  XNOR U7573 ( .A(n4512), .B(n7364), .Z(n7366) );
  NAND U7574 ( .A(n7369), .B(e_input[822]), .Z(n4512) );
  NAND U7575 ( .A(n6112), .B(e_input[822]), .Z(n7369) );
  XOR U7576 ( .A(n7370), .B(n7371), .Z(n7364) );
  ANDN U7577 ( .A(n7372), .B(n4513), .Z(n7371) );
  XOR U7578 ( .A(n7373), .B(n7374), .Z(n4513) );
  IV U7579 ( .A(n7370), .Z(n7373) );
  XNOR U7580 ( .A(n4514), .B(n7370), .Z(n7372) );
  NAND U7581 ( .A(n7375), .B(e_input[821]), .Z(n4514) );
  NAND U7582 ( .A(n6112), .B(e_input[821]), .Z(n7375) );
  XOR U7583 ( .A(n7376), .B(n7377), .Z(n7370) );
  ANDN U7584 ( .A(n7378), .B(n4515), .Z(n7377) );
  XOR U7585 ( .A(n7379), .B(n7380), .Z(n4515) );
  IV U7586 ( .A(n7376), .Z(n7379) );
  XNOR U7587 ( .A(n4516), .B(n7376), .Z(n7378) );
  NAND U7588 ( .A(n7381), .B(e_input[820]), .Z(n4516) );
  NAND U7589 ( .A(n6112), .B(e_input[820]), .Z(n7381) );
  XOR U7590 ( .A(n7382), .B(n7383), .Z(n7376) );
  ANDN U7591 ( .A(n7384), .B(n4519), .Z(n7383) );
  XOR U7592 ( .A(n7385), .B(n7386), .Z(n4519) );
  IV U7593 ( .A(n7382), .Z(n7385) );
  XNOR U7594 ( .A(n4520), .B(n7382), .Z(n7384) );
  NAND U7595 ( .A(n7387), .B(e_input[819]), .Z(n4520) );
  NAND U7596 ( .A(n6112), .B(e_input[819]), .Z(n7387) );
  XOR U7597 ( .A(n7388), .B(n7389), .Z(n7382) );
  ANDN U7598 ( .A(n7390), .B(n4521), .Z(n7389) );
  XOR U7599 ( .A(n7391), .B(n7392), .Z(n4521) );
  IV U7600 ( .A(n7388), .Z(n7391) );
  XNOR U7601 ( .A(n4522), .B(n7388), .Z(n7390) );
  NAND U7602 ( .A(n7393), .B(e_input[818]), .Z(n4522) );
  NAND U7603 ( .A(n6112), .B(e_input[818]), .Z(n7393) );
  XOR U7604 ( .A(n7394), .B(n7395), .Z(n7388) );
  ANDN U7605 ( .A(n7396), .B(n4523), .Z(n7395) );
  XOR U7606 ( .A(n7397), .B(n7398), .Z(n4523) );
  IV U7607 ( .A(n7394), .Z(n7397) );
  XNOR U7608 ( .A(n4524), .B(n7394), .Z(n7396) );
  NAND U7609 ( .A(n7399), .B(e_input[817]), .Z(n4524) );
  NAND U7610 ( .A(n6112), .B(e_input[817]), .Z(n7399) );
  XOR U7611 ( .A(n7400), .B(n7401), .Z(n7394) );
  ANDN U7612 ( .A(n7402), .B(n4525), .Z(n7401) );
  XOR U7613 ( .A(n7403), .B(n7404), .Z(n4525) );
  IV U7614 ( .A(n7400), .Z(n7403) );
  XNOR U7615 ( .A(n4526), .B(n7400), .Z(n7402) );
  NAND U7616 ( .A(n7405), .B(e_input[816]), .Z(n4526) );
  NAND U7617 ( .A(n6112), .B(e_input[816]), .Z(n7405) );
  XOR U7618 ( .A(n7406), .B(n7407), .Z(n7400) );
  ANDN U7619 ( .A(n7408), .B(n4527), .Z(n7407) );
  XOR U7620 ( .A(n7409), .B(n7410), .Z(n4527) );
  IV U7621 ( .A(n7406), .Z(n7409) );
  XNOR U7622 ( .A(n4528), .B(n7406), .Z(n7408) );
  NAND U7623 ( .A(n7411), .B(e_input[815]), .Z(n4528) );
  NAND U7624 ( .A(n6112), .B(e_input[815]), .Z(n7411) );
  XOR U7625 ( .A(n7412), .B(n7413), .Z(n7406) );
  ANDN U7626 ( .A(n7414), .B(n4529), .Z(n7413) );
  XOR U7627 ( .A(n7415), .B(n7416), .Z(n4529) );
  IV U7628 ( .A(n7412), .Z(n7415) );
  XNOR U7629 ( .A(n4530), .B(n7412), .Z(n7414) );
  NAND U7630 ( .A(n7417), .B(e_input[814]), .Z(n4530) );
  NAND U7631 ( .A(n6112), .B(e_input[814]), .Z(n7417) );
  XOR U7632 ( .A(n7418), .B(n7419), .Z(n7412) );
  ANDN U7633 ( .A(n7420), .B(n4531), .Z(n7419) );
  XOR U7634 ( .A(n7421), .B(n7422), .Z(n4531) );
  IV U7635 ( .A(n7418), .Z(n7421) );
  XNOR U7636 ( .A(n4532), .B(n7418), .Z(n7420) );
  NAND U7637 ( .A(n7423), .B(e_input[813]), .Z(n4532) );
  NAND U7638 ( .A(n6112), .B(e_input[813]), .Z(n7423) );
  XOR U7639 ( .A(n7424), .B(n7425), .Z(n7418) );
  ANDN U7640 ( .A(n7426), .B(n4533), .Z(n7425) );
  XOR U7641 ( .A(n7427), .B(n7428), .Z(n4533) );
  IV U7642 ( .A(n7424), .Z(n7427) );
  XNOR U7643 ( .A(n4534), .B(n7424), .Z(n7426) );
  NAND U7644 ( .A(n7429), .B(e_input[812]), .Z(n4534) );
  NAND U7645 ( .A(n6112), .B(e_input[812]), .Z(n7429) );
  XOR U7646 ( .A(n7430), .B(n7431), .Z(n7424) );
  ANDN U7647 ( .A(n7432), .B(n4535), .Z(n7431) );
  XOR U7648 ( .A(n7433), .B(n7434), .Z(n4535) );
  IV U7649 ( .A(n7430), .Z(n7433) );
  XNOR U7650 ( .A(n4536), .B(n7430), .Z(n7432) );
  NAND U7651 ( .A(n7435), .B(e_input[811]), .Z(n4536) );
  NAND U7652 ( .A(n6112), .B(e_input[811]), .Z(n7435) );
  XOR U7653 ( .A(n7436), .B(n7437), .Z(n7430) );
  ANDN U7654 ( .A(n7438), .B(n4537), .Z(n7437) );
  XOR U7655 ( .A(n7439), .B(n7440), .Z(n4537) );
  IV U7656 ( .A(n7436), .Z(n7439) );
  XNOR U7657 ( .A(n4538), .B(n7436), .Z(n7438) );
  NAND U7658 ( .A(n7441), .B(e_input[810]), .Z(n4538) );
  NAND U7659 ( .A(n6112), .B(e_input[810]), .Z(n7441) );
  XOR U7660 ( .A(n7442), .B(n7443), .Z(n7436) );
  ANDN U7661 ( .A(n7444), .B(n4541), .Z(n7443) );
  XOR U7662 ( .A(n7445), .B(n7446), .Z(n4541) );
  IV U7663 ( .A(n7442), .Z(n7445) );
  XNOR U7664 ( .A(n4542), .B(n7442), .Z(n7444) );
  NAND U7665 ( .A(n7447), .B(e_input[809]), .Z(n4542) );
  NAND U7666 ( .A(n6112), .B(e_input[809]), .Z(n7447) );
  XOR U7667 ( .A(n7448), .B(n7449), .Z(n7442) );
  ANDN U7668 ( .A(n7450), .B(n4543), .Z(n7449) );
  XOR U7669 ( .A(n7451), .B(n7452), .Z(n4543) );
  IV U7670 ( .A(n7448), .Z(n7451) );
  XNOR U7671 ( .A(n4544), .B(n7448), .Z(n7450) );
  NAND U7672 ( .A(n7453), .B(e_input[808]), .Z(n4544) );
  NAND U7673 ( .A(n6112), .B(e_input[808]), .Z(n7453) );
  XOR U7674 ( .A(n7454), .B(n7455), .Z(n7448) );
  ANDN U7675 ( .A(n7456), .B(n4545), .Z(n7455) );
  XOR U7676 ( .A(n7457), .B(n7458), .Z(n4545) );
  IV U7677 ( .A(n7454), .Z(n7457) );
  XNOR U7678 ( .A(n4546), .B(n7454), .Z(n7456) );
  NAND U7679 ( .A(n7459), .B(e_input[807]), .Z(n4546) );
  NAND U7680 ( .A(n6112), .B(e_input[807]), .Z(n7459) );
  XOR U7681 ( .A(n7460), .B(n7461), .Z(n7454) );
  ANDN U7682 ( .A(n7462), .B(n4547), .Z(n7461) );
  XOR U7683 ( .A(n7463), .B(n7464), .Z(n4547) );
  IV U7684 ( .A(n7460), .Z(n7463) );
  XNOR U7685 ( .A(n4548), .B(n7460), .Z(n7462) );
  NAND U7686 ( .A(n7465), .B(e_input[806]), .Z(n4548) );
  NAND U7687 ( .A(n6112), .B(e_input[806]), .Z(n7465) );
  XOR U7688 ( .A(n7466), .B(n7467), .Z(n7460) );
  ANDN U7689 ( .A(n7468), .B(n4549), .Z(n7467) );
  XOR U7690 ( .A(n7469), .B(n7470), .Z(n4549) );
  IV U7691 ( .A(n7466), .Z(n7469) );
  XNOR U7692 ( .A(n4550), .B(n7466), .Z(n7468) );
  NAND U7693 ( .A(n7471), .B(e_input[805]), .Z(n4550) );
  NAND U7694 ( .A(n6112), .B(e_input[805]), .Z(n7471) );
  XOR U7695 ( .A(n7472), .B(n7473), .Z(n7466) );
  ANDN U7696 ( .A(n7474), .B(n4551), .Z(n7473) );
  XOR U7697 ( .A(n7475), .B(n7476), .Z(n4551) );
  IV U7698 ( .A(n7472), .Z(n7475) );
  XNOR U7699 ( .A(n4552), .B(n7472), .Z(n7474) );
  NAND U7700 ( .A(n7477), .B(e_input[804]), .Z(n4552) );
  NAND U7701 ( .A(n6112), .B(e_input[804]), .Z(n7477) );
  XOR U7702 ( .A(n7478), .B(n7479), .Z(n7472) );
  ANDN U7703 ( .A(n7480), .B(n4553), .Z(n7479) );
  XOR U7704 ( .A(n7481), .B(n7482), .Z(n4553) );
  IV U7705 ( .A(n7478), .Z(n7481) );
  XNOR U7706 ( .A(n4554), .B(n7478), .Z(n7480) );
  NAND U7707 ( .A(n7483), .B(e_input[803]), .Z(n4554) );
  NAND U7708 ( .A(n6112), .B(e_input[803]), .Z(n7483) );
  XOR U7709 ( .A(n7484), .B(n7485), .Z(n7478) );
  ANDN U7710 ( .A(n7486), .B(n4555), .Z(n7485) );
  XOR U7711 ( .A(n7487), .B(n7488), .Z(n4555) );
  IV U7712 ( .A(n7484), .Z(n7487) );
  XNOR U7713 ( .A(n4556), .B(n7484), .Z(n7486) );
  NAND U7714 ( .A(n7489), .B(e_input[802]), .Z(n4556) );
  NAND U7715 ( .A(n6112), .B(e_input[802]), .Z(n7489) );
  XOR U7716 ( .A(n7490), .B(n7491), .Z(n7484) );
  ANDN U7717 ( .A(n7492), .B(n4557), .Z(n7491) );
  XOR U7718 ( .A(n7493), .B(n7494), .Z(n4557) );
  IV U7719 ( .A(n7490), .Z(n7493) );
  XNOR U7720 ( .A(n4558), .B(n7490), .Z(n7492) );
  NAND U7721 ( .A(n7495), .B(e_input[801]), .Z(n4558) );
  NAND U7722 ( .A(n6112), .B(e_input[801]), .Z(n7495) );
  XOR U7723 ( .A(n7496), .B(n7497), .Z(n7490) );
  ANDN U7724 ( .A(n7498), .B(n4559), .Z(n7497) );
  XOR U7725 ( .A(n7499), .B(n7500), .Z(n4559) );
  IV U7726 ( .A(n7496), .Z(n7499) );
  XNOR U7727 ( .A(n4560), .B(n7496), .Z(n7498) );
  NAND U7728 ( .A(n7501), .B(e_input[800]), .Z(n4560) );
  NAND U7729 ( .A(n6112), .B(e_input[800]), .Z(n7501) );
  XOR U7730 ( .A(n7502), .B(n7503), .Z(n7496) );
  ANDN U7731 ( .A(n7504), .B(n4565), .Z(n7503) );
  XOR U7732 ( .A(n7505), .B(n7506), .Z(n4565) );
  IV U7733 ( .A(n7502), .Z(n7505) );
  XNOR U7734 ( .A(n4566), .B(n7502), .Z(n7504) );
  NAND U7735 ( .A(n7507), .B(e_input[799]), .Z(n4566) );
  NAND U7736 ( .A(n6112), .B(e_input[799]), .Z(n7507) );
  XOR U7737 ( .A(n7508), .B(n7509), .Z(n7502) );
  ANDN U7738 ( .A(n7510), .B(n4567), .Z(n7509) );
  XOR U7739 ( .A(n7511), .B(n7512), .Z(n4567) );
  IV U7740 ( .A(n7508), .Z(n7511) );
  XNOR U7741 ( .A(n4568), .B(n7508), .Z(n7510) );
  NAND U7742 ( .A(n7513), .B(e_input[798]), .Z(n4568) );
  NAND U7743 ( .A(n6112), .B(e_input[798]), .Z(n7513) );
  XOR U7744 ( .A(n7514), .B(n7515), .Z(n7508) );
  ANDN U7745 ( .A(n7516), .B(n4569), .Z(n7515) );
  XOR U7746 ( .A(n7517), .B(n7518), .Z(n4569) );
  IV U7747 ( .A(n7514), .Z(n7517) );
  XNOR U7748 ( .A(n4570), .B(n7514), .Z(n7516) );
  NAND U7749 ( .A(n7519), .B(e_input[797]), .Z(n4570) );
  NAND U7750 ( .A(n6112), .B(e_input[797]), .Z(n7519) );
  XOR U7751 ( .A(n7520), .B(n7521), .Z(n7514) );
  ANDN U7752 ( .A(n7522), .B(n4571), .Z(n7521) );
  XOR U7753 ( .A(n7523), .B(n7524), .Z(n4571) );
  IV U7754 ( .A(n7520), .Z(n7523) );
  XNOR U7755 ( .A(n4572), .B(n7520), .Z(n7522) );
  NAND U7756 ( .A(n7525), .B(e_input[796]), .Z(n4572) );
  NAND U7757 ( .A(n6112), .B(e_input[796]), .Z(n7525) );
  XOR U7758 ( .A(n7526), .B(n7527), .Z(n7520) );
  ANDN U7759 ( .A(n7528), .B(n4573), .Z(n7527) );
  XOR U7760 ( .A(n7529), .B(n7530), .Z(n4573) );
  IV U7761 ( .A(n7526), .Z(n7529) );
  XNOR U7762 ( .A(n4574), .B(n7526), .Z(n7528) );
  NAND U7763 ( .A(n7531), .B(e_input[795]), .Z(n4574) );
  NAND U7764 ( .A(n6112), .B(e_input[795]), .Z(n7531) );
  XOR U7765 ( .A(n7532), .B(n7533), .Z(n7526) );
  ANDN U7766 ( .A(n7534), .B(n4575), .Z(n7533) );
  XOR U7767 ( .A(n7535), .B(n7536), .Z(n4575) );
  IV U7768 ( .A(n7532), .Z(n7535) );
  XNOR U7769 ( .A(n4576), .B(n7532), .Z(n7534) );
  NAND U7770 ( .A(n7537), .B(e_input[794]), .Z(n4576) );
  NAND U7771 ( .A(n6112), .B(e_input[794]), .Z(n7537) );
  XOR U7772 ( .A(n7538), .B(n7539), .Z(n7532) );
  ANDN U7773 ( .A(n7540), .B(n4577), .Z(n7539) );
  XOR U7774 ( .A(n7541), .B(n7542), .Z(n4577) );
  IV U7775 ( .A(n7538), .Z(n7541) );
  XNOR U7776 ( .A(n4578), .B(n7538), .Z(n7540) );
  NAND U7777 ( .A(n7543), .B(e_input[793]), .Z(n4578) );
  NAND U7778 ( .A(n6112), .B(e_input[793]), .Z(n7543) );
  XOR U7779 ( .A(n7544), .B(n7545), .Z(n7538) );
  ANDN U7780 ( .A(n7546), .B(n4579), .Z(n7545) );
  XOR U7781 ( .A(n7547), .B(n7548), .Z(n4579) );
  IV U7782 ( .A(n7544), .Z(n7547) );
  XNOR U7783 ( .A(n4580), .B(n7544), .Z(n7546) );
  NAND U7784 ( .A(n7549), .B(e_input[792]), .Z(n4580) );
  NAND U7785 ( .A(n6112), .B(e_input[792]), .Z(n7549) );
  XOR U7786 ( .A(n7550), .B(n7551), .Z(n7544) );
  ANDN U7787 ( .A(n7552), .B(n4581), .Z(n7551) );
  XOR U7788 ( .A(n7553), .B(n7554), .Z(n4581) );
  IV U7789 ( .A(n7550), .Z(n7553) );
  XNOR U7790 ( .A(n4582), .B(n7550), .Z(n7552) );
  NAND U7791 ( .A(n7555), .B(e_input[791]), .Z(n4582) );
  NAND U7792 ( .A(n6112), .B(e_input[791]), .Z(n7555) );
  XOR U7793 ( .A(n7556), .B(n7557), .Z(n7550) );
  ANDN U7794 ( .A(n7558), .B(n4583), .Z(n7557) );
  XOR U7795 ( .A(n7559), .B(n7560), .Z(n4583) );
  IV U7796 ( .A(n7556), .Z(n7559) );
  XNOR U7797 ( .A(n4584), .B(n7556), .Z(n7558) );
  NAND U7798 ( .A(n7561), .B(e_input[790]), .Z(n4584) );
  NAND U7799 ( .A(n6112), .B(e_input[790]), .Z(n7561) );
  XOR U7800 ( .A(n7562), .B(n7563), .Z(n7556) );
  ANDN U7801 ( .A(n7564), .B(n4587), .Z(n7563) );
  XOR U7802 ( .A(n7565), .B(n7566), .Z(n4587) );
  IV U7803 ( .A(n7562), .Z(n7565) );
  XNOR U7804 ( .A(n4588), .B(n7562), .Z(n7564) );
  NAND U7805 ( .A(n7567), .B(e_input[789]), .Z(n4588) );
  NAND U7806 ( .A(n6112), .B(e_input[789]), .Z(n7567) );
  XOR U7807 ( .A(n7568), .B(n7569), .Z(n7562) );
  ANDN U7808 ( .A(n7570), .B(n4589), .Z(n7569) );
  XOR U7809 ( .A(n7571), .B(n7572), .Z(n4589) );
  IV U7810 ( .A(n7568), .Z(n7571) );
  XNOR U7811 ( .A(n4590), .B(n7568), .Z(n7570) );
  NAND U7812 ( .A(n7573), .B(e_input[788]), .Z(n4590) );
  NAND U7813 ( .A(n6112), .B(e_input[788]), .Z(n7573) );
  XOR U7814 ( .A(n7574), .B(n7575), .Z(n7568) );
  ANDN U7815 ( .A(n7576), .B(n4591), .Z(n7575) );
  XOR U7816 ( .A(n7577), .B(n7578), .Z(n4591) );
  IV U7817 ( .A(n7574), .Z(n7577) );
  XNOR U7818 ( .A(n4592), .B(n7574), .Z(n7576) );
  NAND U7819 ( .A(n7579), .B(e_input[787]), .Z(n4592) );
  NAND U7820 ( .A(n6112), .B(e_input[787]), .Z(n7579) );
  XOR U7821 ( .A(n7580), .B(n7581), .Z(n7574) );
  ANDN U7822 ( .A(n7582), .B(n4593), .Z(n7581) );
  XOR U7823 ( .A(n7583), .B(n7584), .Z(n4593) );
  IV U7824 ( .A(n7580), .Z(n7583) );
  XNOR U7825 ( .A(n4594), .B(n7580), .Z(n7582) );
  NAND U7826 ( .A(n7585), .B(e_input[786]), .Z(n4594) );
  NAND U7827 ( .A(n6112), .B(e_input[786]), .Z(n7585) );
  XOR U7828 ( .A(n7586), .B(n7587), .Z(n7580) );
  ANDN U7829 ( .A(n7588), .B(n4595), .Z(n7587) );
  XOR U7830 ( .A(n7589), .B(n7590), .Z(n4595) );
  IV U7831 ( .A(n7586), .Z(n7589) );
  XNOR U7832 ( .A(n4596), .B(n7586), .Z(n7588) );
  NAND U7833 ( .A(n7591), .B(e_input[785]), .Z(n4596) );
  NAND U7834 ( .A(n6112), .B(e_input[785]), .Z(n7591) );
  XOR U7835 ( .A(n7592), .B(n7593), .Z(n7586) );
  ANDN U7836 ( .A(n7594), .B(n4597), .Z(n7593) );
  XOR U7837 ( .A(n7595), .B(n7596), .Z(n4597) );
  IV U7838 ( .A(n7592), .Z(n7595) );
  XNOR U7839 ( .A(n4598), .B(n7592), .Z(n7594) );
  NAND U7840 ( .A(n7597), .B(e_input[784]), .Z(n4598) );
  NAND U7841 ( .A(n6112), .B(e_input[784]), .Z(n7597) );
  XOR U7842 ( .A(n7598), .B(n7599), .Z(n7592) );
  ANDN U7843 ( .A(n7600), .B(n4599), .Z(n7599) );
  XOR U7844 ( .A(n7601), .B(n7602), .Z(n4599) );
  IV U7845 ( .A(n7598), .Z(n7601) );
  XNOR U7846 ( .A(n4600), .B(n7598), .Z(n7600) );
  NAND U7847 ( .A(n7603), .B(e_input[783]), .Z(n4600) );
  NAND U7848 ( .A(n6112), .B(e_input[783]), .Z(n7603) );
  XOR U7849 ( .A(n7604), .B(n7605), .Z(n7598) );
  ANDN U7850 ( .A(n7606), .B(n4601), .Z(n7605) );
  XOR U7851 ( .A(n7607), .B(n7608), .Z(n4601) );
  IV U7852 ( .A(n7604), .Z(n7607) );
  XNOR U7853 ( .A(n4602), .B(n7604), .Z(n7606) );
  NAND U7854 ( .A(n7609), .B(e_input[782]), .Z(n4602) );
  NAND U7855 ( .A(n6112), .B(e_input[782]), .Z(n7609) );
  XOR U7856 ( .A(n7610), .B(n7611), .Z(n7604) );
  ANDN U7857 ( .A(n7612), .B(n4603), .Z(n7611) );
  XOR U7858 ( .A(n7613), .B(n7614), .Z(n4603) );
  IV U7859 ( .A(n7610), .Z(n7613) );
  XNOR U7860 ( .A(n4604), .B(n7610), .Z(n7612) );
  NAND U7861 ( .A(n7615), .B(e_input[781]), .Z(n4604) );
  NAND U7862 ( .A(n6112), .B(e_input[781]), .Z(n7615) );
  XOR U7863 ( .A(n7616), .B(n7617), .Z(n7610) );
  ANDN U7864 ( .A(n7618), .B(n4605), .Z(n7617) );
  XOR U7865 ( .A(n7619), .B(n7620), .Z(n4605) );
  IV U7866 ( .A(n7616), .Z(n7619) );
  XNOR U7867 ( .A(n4606), .B(n7616), .Z(n7618) );
  NAND U7868 ( .A(n7621), .B(e_input[780]), .Z(n4606) );
  NAND U7869 ( .A(n6112), .B(e_input[780]), .Z(n7621) );
  XOR U7870 ( .A(n7622), .B(n7623), .Z(n7616) );
  ANDN U7871 ( .A(n7624), .B(n4609), .Z(n7623) );
  XOR U7872 ( .A(n7625), .B(n7626), .Z(n4609) );
  IV U7873 ( .A(n7622), .Z(n7625) );
  XNOR U7874 ( .A(n4610), .B(n7622), .Z(n7624) );
  NAND U7875 ( .A(n7627), .B(e_input[779]), .Z(n4610) );
  NAND U7876 ( .A(n6112), .B(e_input[779]), .Z(n7627) );
  XOR U7877 ( .A(n7628), .B(n7629), .Z(n7622) );
  ANDN U7878 ( .A(n7630), .B(n4611), .Z(n7629) );
  XOR U7879 ( .A(n7631), .B(n7632), .Z(n4611) );
  IV U7880 ( .A(n7628), .Z(n7631) );
  XNOR U7881 ( .A(n4612), .B(n7628), .Z(n7630) );
  NAND U7882 ( .A(n7633), .B(e_input[778]), .Z(n4612) );
  NAND U7883 ( .A(n6112), .B(e_input[778]), .Z(n7633) );
  XOR U7884 ( .A(n7634), .B(n7635), .Z(n7628) );
  ANDN U7885 ( .A(n7636), .B(n4613), .Z(n7635) );
  XOR U7886 ( .A(n7637), .B(n7638), .Z(n4613) );
  IV U7887 ( .A(n7634), .Z(n7637) );
  XNOR U7888 ( .A(n4614), .B(n7634), .Z(n7636) );
  NAND U7889 ( .A(n7639), .B(e_input[777]), .Z(n4614) );
  NAND U7890 ( .A(n6112), .B(e_input[777]), .Z(n7639) );
  XOR U7891 ( .A(n7640), .B(n7641), .Z(n7634) );
  ANDN U7892 ( .A(n7642), .B(n4615), .Z(n7641) );
  XOR U7893 ( .A(n7643), .B(n7644), .Z(n4615) );
  IV U7894 ( .A(n7640), .Z(n7643) );
  XNOR U7895 ( .A(n4616), .B(n7640), .Z(n7642) );
  NAND U7896 ( .A(n7645), .B(e_input[776]), .Z(n4616) );
  NAND U7897 ( .A(n6112), .B(e_input[776]), .Z(n7645) );
  XOR U7898 ( .A(n7646), .B(n7647), .Z(n7640) );
  ANDN U7899 ( .A(n7648), .B(n4617), .Z(n7647) );
  XOR U7900 ( .A(n7649), .B(n7650), .Z(n4617) );
  IV U7901 ( .A(n7646), .Z(n7649) );
  XNOR U7902 ( .A(n4618), .B(n7646), .Z(n7648) );
  NAND U7903 ( .A(n7651), .B(e_input[775]), .Z(n4618) );
  NAND U7904 ( .A(n6112), .B(e_input[775]), .Z(n7651) );
  XOR U7905 ( .A(n7652), .B(n7653), .Z(n7646) );
  ANDN U7906 ( .A(n7654), .B(n4619), .Z(n7653) );
  XOR U7907 ( .A(n7655), .B(n7656), .Z(n4619) );
  IV U7908 ( .A(n7652), .Z(n7655) );
  XNOR U7909 ( .A(n4620), .B(n7652), .Z(n7654) );
  NAND U7910 ( .A(n7657), .B(e_input[774]), .Z(n4620) );
  NAND U7911 ( .A(n6112), .B(e_input[774]), .Z(n7657) );
  XOR U7912 ( .A(n7658), .B(n7659), .Z(n7652) );
  ANDN U7913 ( .A(n7660), .B(n4621), .Z(n7659) );
  XOR U7914 ( .A(n7661), .B(n7662), .Z(n4621) );
  IV U7915 ( .A(n7658), .Z(n7661) );
  XNOR U7916 ( .A(n4622), .B(n7658), .Z(n7660) );
  NAND U7917 ( .A(n7663), .B(e_input[773]), .Z(n4622) );
  NAND U7918 ( .A(n6112), .B(e_input[773]), .Z(n7663) );
  XOR U7919 ( .A(n7664), .B(n7665), .Z(n7658) );
  ANDN U7920 ( .A(n7666), .B(n4623), .Z(n7665) );
  XOR U7921 ( .A(n7667), .B(n7668), .Z(n4623) );
  IV U7922 ( .A(n7664), .Z(n7667) );
  XNOR U7923 ( .A(n4624), .B(n7664), .Z(n7666) );
  NAND U7924 ( .A(n7669), .B(e_input[772]), .Z(n4624) );
  NAND U7925 ( .A(n6112), .B(e_input[772]), .Z(n7669) );
  XOR U7926 ( .A(n7670), .B(n7671), .Z(n7664) );
  ANDN U7927 ( .A(n7672), .B(n4625), .Z(n7671) );
  XOR U7928 ( .A(n7673), .B(n7674), .Z(n4625) );
  IV U7929 ( .A(n7670), .Z(n7673) );
  XNOR U7930 ( .A(n4626), .B(n7670), .Z(n7672) );
  NAND U7931 ( .A(n7675), .B(e_input[771]), .Z(n4626) );
  NAND U7932 ( .A(n6112), .B(e_input[771]), .Z(n7675) );
  XOR U7933 ( .A(n7676), .B(n7677), .Z(n7670) );
  ANDN U7934 ( .A(n7678), .B(n4627), .Z(n7677) );
  XOR U7935 ( .A(n7679), .B(n7680), .Z(n4627) );
  IV U7936 ( .A(n7676), .Z(n7679) );
  XNOR U7937 ( .A(n4628), .B(n7676), .Z(n7678) );
  NAND U7938 ( .A(n7681), .B(e_input[770]), .Z(n4628) );
  NAND U7939 ( .A(n6112), .B(e_input[770]), .Z(n7681) );
  XOR U7940 ( .A(n7682), .B(n7683), .Z(n7676) );
  ANDN U7941 ( .A(n7684), .B(n4631), .Z(n7683) );
  XOR U7942 ( .A(n7685), .B(n7686), .Z(n4631) );
  IV U7943 ( .A(n7682), .Z(n7685) );
  XNOR U7944 ( .A(n4632), .B(n7682), .Z(n7684) );
  NAND U7945 ( .A(n7687), .B(e_input[769]), .Z(n4632) );
  NAND U7946 ( .A(n6112), .B(e_input[769]), .Z(n7687) );
  XOR U7947 ( .A(n7688), .B(n7689), .Z(n7682) );
  ANDN U7948 ( .A(n7690), .B(n4633), .Z(n7689) );
  XOR U7949 ( .A(n7691), .B(n7692), .Z(n4633) );
  IV U7950 ( .A(n7688), .Z(n7691) );
  XNOR U7951 ( .A(n4634), .B(n7688), .Z(n7690) );
  NAND U7952 ( .A(n7693), .B(e_input[768]), .Z(n4634) );
  NAND U7953 ( .A(n6112), .B(e_input[768]), .Z(n7693) );
  XOR U7954 ( .A(n7694), .B(n7695), .Z(n7688) );
  ANDN U7955 ( .A(n7696), .B(n4635), .Z(n7695) );
  XOR U7956 ( .A(n7697), .B(n7698), .Z(n4635) );
  IV U7957 ( .A(n7694), .Z(n7697) );
  XNOR U7958 ( .A(n4636), .B(n7694), .Z(n7696) );
  NAND U7959 ( .A(n7699), .B(e_input[767]), .Z(n4636) );
  NAND U7960 ( .A(n6112), .B(e_input[767]), .Z(n7699) );
  XOR U7961 ( .A(n7700), .B(n7701), .Z(n7694) );
  ANDN U7962 ( .A(n7702), .B(n4637), .Z(n7701) );
  XOR U7963 ( .A(n7703), .B(n7704), .Z(n4637) );
  IV U7964 ( .A(n7700), .Z(n7703) );
  XNOR U7965 ( .A(n4638), .B(n7700), .Z(n7702) );
  NAND U7966 ( .A(n7705), .B(e_input[766]), .Z(n4638) );
  NAND U7967 ( .A(n6112), .B(e_input[766]), .Z(n7705) );
  XOR U7968 ( .A(n7706), .B(n7707), .Z(n7700) );
  ANDN U7969 ( .A(n7708), .B(n4639), .Z(n7707) );
  XOR U7970 ( .A(n7709), .B(n7710), .Z(n4639) );
  IV U7971 ( .A(n7706), .Z(n7709) );
  XNOR U7972 ( .A(n4640), .B(n7706), .Z(n7708) );
  NAND U7973 ( .A(n7711), .B(e_input[765]), .Z(n4640) );
  NAND U7974 ( .A(n6112), .B(e_input[765]), .Z(n7711) );
  XOR U7975 ( .A(n7712), .B(n7713), .Z(n7706) );
  ANDN U7976 ( .A(n7714), .B(n4641), .Z(n7713) );
  XOR U7977 ( .A(n7715), .B(n7716), .Z(n4641) );
  IV U7978 ( .A(n7712), .Z(n7715) );
  XNOR U7979 ( .A(n4642), .B(n7712), .Z(n7714) );
  NAND U7980 ( .A(n7717), .B(e_input[764]), .Z(n4642) );
  NAND U7981 ( .A(n6112), .B(e_input[764]), .Z(n7717) );
  XOR U7982 ( .A(n7718), .B(n7719), .Z(n7712) );
  ANDN U7983 ( .A(n7720), .B(n4643), .Z(n7719) );
  XOR U7984 ( .A(n7721), .B(n7722), .Z(n4643) );
  IV U7985 ( .A(n7718), .Z(n7721) );
  XNOR U7986 ( .A(n4644), .B(n7718), .Z(n7720) );
  NAND U7987 ( .A(n7723), .B(e_input[763]), .Z(n4644) );
  NAND U7988 ( .A(n6112), .B(e_input[763]), .Z(n7723) );
  XOR U7989 ( .A(n7724), .B(n7725), .Z(n7718) );
  ANDN U7990 ( .A(n7726), .B(n4645), .Z(n7725) );
  XOR U7991 ( .A(n7727), .B(n7728), .Z(n4645) );
  IV U7992 ( .A(n7724), .Z(n7727) );
  XNOR U7993 ( .A(n4646), .B(n7724), .Z(n7726) );
  NAND U7994 ( .A(n7729), .B(e_input[762]), .Z(n4646) );
  NAND U7995 ( .A(n6112), .B(e_input[762]), .Z(n7729) );
  XOR U7996 ( .A(n7730), .B(n7731), .Z(n7724) );
  ANDN U7997 ( .A(n7732), .B(n4647), .Z(n7731) );
  XOR U7998 ( .A(n7733), .B(n7734), .Z(n4647) );
  IV U7999 ( .A(n7730), .Z(n7733) );
  XNOR U8000 ( .A(n4648), .B(n7730), .Z(n7732) );
  NAND U8001 ( .A(n7735), .B(e_input[761]), .Z(n4648) );
  NAND U8002 ( .A(n6112), .B(e_input[761]), .Z(n7735) );
  XOR U8003 ( .A(n7736), .B(n7737), .Z(n7730) );
  ANDN U8004 ( .A(n7738), .B(n4649), .Z(n7737) );
  XOR U8005 ( .A(n7739), .B(n7740), .Z(n4649) );
  IV U8006 ( .A(n7736), .Z(n7739) );
  XNOR U8007 ( .A(n4650), .B(n7736), .Z(n7738) );
  NAND U8008 ( .A(n7741), .B(e_input[760]), .Z(n4650) );
  NAND U8009 ( .A(n6112), .B(e_input[760]), .Z(n7741) );
  XOR U8010 ( .A(n7742), .B(n7743), .Z(n7736) );
  ANDN U8011 ( .A(n7744), .B(n4653), .Z(n7743) );
  XOR U8012 ( .A(n7745), .B(n7746), .Z(n4653) );
  IV U8013 ( .A(n7742), .Z(n7745) );
  XNOR U8014 ( .A(n4654), .B(n7742), .Z(n7744) );
  NAND U8015 ( .A(n7747), .B(e_input[759]), .Z(n4654) );
  NAND U8016 ( .A(n6112), .B(e_input[759]), .Z(n7747) );
  XOR U8017 ( .A(n7748), .B(n7749), .Z(n7742) );
  ANDN U8018 ( .A(n7750), .B(n4655), .Z(n7749) );
  XOR U8019 ( .A(n7751), .B(n7752), .Z(n4655) );
  IV U8020 ( .A(n7748), .Z(n7751) );
  XNOR U8021 ( .A(n4656), .B(n7748), .Z(n7750) );
  NAND U8022 ( .A(n7753), .B(e_input[758]), .Z(n4656) );
  NAND U8023 ( .A(n6112), .B(e_input[758]), .Z(n7753) );
  XOR U8024 ( .A(n7754), .B(n7755), .Z(n7748) );
  ANDN U8025 ( .A(n7756), .B(n4657), .Z(n7755) );
  XOR U8026 ( .A(n7757), .B(n7758), .Z(n4657) );
  IV U8027 ( .A(n7754), .Z(n7757) );
  XNOR U8028 ( .A(n4658), .B(n7754), .Z(n7756) );
  NAND U8029 ( .A(n7759), .B(e_input[757]), .Z(n4658) );
  NAND U8030 ( .A(n6112), .B(e_input[757]), .Z(n7759) );
  XOR U8031 ( .A(n7760), .B(n7761), .Z(n7754) );
  ANDN U8032 ( .A(n7762), .B(n4659), .Z(n7761) );
  XOR U8033 ( .A(n7763), .B(n7764), .Z(n4659) );
  IV U8034 ( .A(n7760), .Z(n7763) );
  XNOR U8035 ( .A(n4660), .B(n7760), .Z(n7762) );
  NAND U8036 ( .A(n7765), .B(e_input[756]), .Z(n4660) );
  NAND U8037 ( .A(n6112), .B(e_input[756]), .Z(n7765) );
  XOR U8038 ( .A(n7766), .B(n7767), .Z(n7760) );
  ANDN U8039 ( .A(n7768), .B(n4661), .Z(n7767) );
  XOR U8040 ( .A(n7769), .B(n7770), .Z(n4661) );
  IV U8041 ( .A(n7766), .Z(n7769) );
  XNOR U8042 ( .A(n4662), .B(n7766), .Z(n7768) );
  NAND U8043 ( .A(n7771), .B(e_input[755]), .Z(n4662) );
  NAND U8044 ( .A(n6112), .B(e_input[755]), .Z(n7771) );
  XOR U8045 ( .A(n7772), .B(n7773), .Z(n7766) );
  ANDN U8046 ( .A(n7774), .B(n4663), .Z(n7773) );
  XOR U8047 ( .A(n7775), .B(n7776), .Z(n4663) );
  IV U8048 ( .A(n7772), .Z(n7775) );
  XNOR U8049 ( .A(n4664), .B(n7772), .Z(n7774) );
  NAND U8050 ( .A(n7777), .B(e_input[754]), .Z(n4664) );
  NAND U8051 ( .A(n6112), .B(e_input[754]), .Z(n7777) );
  XOR U8052 ( .A(n7778), .B(n7779), .Z(n7772) );
  ANDN U8053 ( .A(n7780), .B(n4665), .Z(n7779) );
  XOR U8054 ( .A(n7781), .B(n7782), .Z(n4665) );
  IV U8055 ( .A(n7778), .Z(n7781) );
  XNOR U8056 ( .A(n4666), .B(n7778), .Z(n7780) );
  NAND U8057 ( .A(n7783), .B(e_input[753]), .Z(n4666) );
  NAND U8058 ( .A(n6112), .B(e_input[753]), .Z(n7783) );
  XOR U8059 ( .A(n7784), .B(n7785), .Z(n7778) );
  ANDN U8060 ( .A(n7786), .B(n4667), .Z(n7785) );
  XOR U8061 ( .A(n7787), .B(n7788), .Z(n4667) );
  IV U8062 ( .A(n7784), .Z(n7787) );
  XNOR U8063 ( .A(n4668), .B(n7784), .Z(n7786) );
  NAND U8064 ( .A(n7789), .B(e_input[752]), .Z(n4668) );
  NAND U8065 ( .A(n6112), .B(e_input[752]), .Z(n7789) );
  XOR U8066 ( .A(n7790), .B(n7791), .Z(n7784) );
  ANDN U8067 ( .A(n7792), .B(n4669), .Z(n7791) );
  XOR U8068 ( .A(n7793), .B(n7794), .Z(n4669) );
  IV U8069 ( .A(n7790), .Z(n7793) );
  XNOR U8070 ( .A(n4670), .B(n7790), .Z(n7792) );
  NAND U8071 ( .A(n7795), .B(e_input[751]), .Z(n4670) );
  NAND U8072 ( .A(n6112), .B(e_input[751]), .Z(n7795) );
  XOR U8073 ( .A(n7796), .B(n7797), .Z(n7790) );
  ANDN U8074 ( .A(n7798), .B(n4671), .Z(n7797) );
  XOR U8075 ( .A(n7799), .B(n7800), .Z(n4671) );
  IV U8076 ( .A(n7796), .Z(n7799) );
  XNOR U8077 ( .A(n4672), .B(n7796), .Z(n7798) );
  NAND U8078 ( .A(n7801), .B(e_input[750]), .Z(n4672) );
  NAND U8079 ( .A(n6112), .B(e_input[750]), .Z(n7801) );
  XOR U8080 ( .A(n7802), .B(n7803), .Z(n7796) );
  ANDN U8081 ( .A(n7804), .B(n4675), .Z(n7803) );
  XOR U8082 ( .A(n7805), .B(n7806), .Z(n4675) );
  IV U8083 ( .A(n7802), .Z(n7805) );
  XNOR U8084 ( .A(n4676), .B(n7802), .Z(n7804) );
  NAND U8085 ( .A(n7807), .B(e_input[749]), .Z(n4676) );
  NAND U8086 ( .A(n6112), .B(e_input[749]), .Z(n7807) );
  XOR U8087 ( .A(n7808), .B(n7809), .Z(n7802) );
  ANDN U8088 ( .A(n7810), .B(n4677), .Z(n7809) );
  XOR U8089 ( .A(n7811), .B(n7812), .Z(n4677) );
  IV U8090 ( .A(n7808), .Z(n7811) );
  XNOR U8091 ( .A(n4678), .B(n7808), .Z(n7810) );
  NAND U8092 ( .A(n7813), .B(e_input[748]), .Z(n4678) );
  NAND U8093 ( .A(n6112), .B(e_input[748]), .Z(n7813) );
  XOR U8094 ( .A(n7814), .B(n7815), .Z(n7808) );
  ANDN U8095 ( .A(n7816), .B(n4679), .Z(n7815) );
  XOR U8096 ( .A(n7817), .B(n7818), .Z(n4679) );
  IV U8097 ( .A(n7814), .Z(n7817) );
  XNOR U8098 ( .A(n4680), .B(n7814), .Z(n7816) );
  NAND U8099 ( .A(n7819), .B(e_input[747]), .Z(n4680) );
  NAND U8100 ( .A(n6112), .B(e_input[747]), .Z(n7819) );
  XOR U8101 ( .A(n7820), .B(n7821), .Z(n7814) );
  ANDN U8102 ( .A(n7822), .B(n4681), .Z(n7821) );
  XOR U8103 ( .A(n7823), .B(n7824), .Z(n4681) );
  IV U8104 ( .A(n7820), .Z(n7823) );
  XNOR U8105 ( .A(n4682), .B(n7820), .Z(n7822) );
  NAND U8106 ( .A(n7825), .B(e_input[746]), .Z(n4682) );
  NAND U8107 ( .A(n6112), .B(e_input[746]), .Z(n7825) );
  XOR U8108 ( .A(n7826), .B(n7827), .Z(n7820) );
  ANDN U8109 ( .A(n7828), .B(n4683), .Z(n7827) );
  XOR U8110 ( .A(n7829), .B(n7830), .Z(n4683) );
  IV U8111 ( .A(n7826), .Z(n7829) );
  XNOR U8112 ( .A(n4684), .B(n7826), .Z(n7828) );
  NAND U8113 ( .A(n7831), .B(e_input[745]), .Z(n4684) );
  NAND U8114 ( .A(n6112), .B(e_input[745]), .Z(n7831) );
  XOR U8115 ( .A(n7832), .B(n7833), .Z(n7826) );
  ANDN U8116 ( .A(n7834), .B(n4685), .Z(n7833) );
  XOR U8117 ( .A(n7835), .B(n7836), .Z(n4685) );
  IV U8118 ( .A(n7832), .Z(n7835) );
  XNOR U8119 ( .A(n4686), .B(n7832), .Z(n7834) );
  NAND U8120 ( .A(n7837), .B(e_input[744]), .Z(n4686) );
  NAND U8121 ( .A(n6112), .B(e_input[744]), .Z(n7837) );
  XOR U8122 ( .A(n7838), .B(n7839), .Z(n7832) );
  ANDN U8123 ( .A(n7840), .B(n4687), .Z(n7839) );
  XOR U8124 ( .A(n7841), .B(n7842), .Z(n4687) );
  IV U8125 ( .A(n7838), .Z(n7841) );
  XNOR U8126 ( .A(n4688), .B(n7838), .Z(n7840) );
  NAND U8127 ( .A(n7843), .B(e_input[743]), .Z(n4688) );
  NAND U8128 ( .A(n6112), .B(e_input[743]), .Z(n7843) );
  XOR U8129 ( .A(n7844), .B(n7845), .Z(n7838) );
  ANDN U8130 ( .A(n7846), .B(n4689), .Z(n7845) );
  XOR U8131 ( .A(n7847), .B(n7848), .Z(n4689) );
  IV U8132 ( .A(n7844), .Z(n7847) );
  XNOR U8133 ( .A(n4690), .B(n7844), .Z(n7846) );
  NAND U8134 ( .A(n7849), .B(e_input[742]), .Z(n4690) );
  NAND U8135 ( .A(n6112), .B(e_input[742]), .Z(n7849) );
  XOR U8136 ( .A(n7850), .B(n7851), .Z(n7844) );
  ANDN U8137 ( .A(n7852), .B(n4691), .Z(n7851) );
  XOR U8138 ( .A(n7853), .B(n7854), .Z(n4691) );
  IV U8139 ( .A(n7850), .Z(n7853) );
  XNOR U8140 ( .A(n4692), .B(n7850), .Z(n7852) );
  NAND U8141 ( .A(n7855), .B(e_input[741]), .Z(n4692) );
  NAND U8142 ( .A(n6112), .B(e_input[741]), .Z(n7855) );
  XOR U8143 ( .A(n7856), .B(n7857), .Z(n7850) );
  ANDN U8144 ( .A(n7858), .B(n4693), .Z(n7857) );
  XOR U8145 ( .A(n7859), .B(n7860), .Z(n4693) );
  IV U8146 ( .A(n7856), .Z(n7859) );
  XNOR U8147 ( .A(n4694), .B(n7856), .Z(n7858) );
  NAND U8148 ( .A(n7861), .B(e_input[740]), .Z(n4694) );
  NAND U8149 ( .A(n6112), .B(e_input[740]), .Z(n7861) );
  XOR U8150 ( .A(n7862), .B(n7863), .Z(n7856) );
  ANDN U8151 ( .A(n7864), .B(n4697), .Z(n7863) );
  XOR U8152 ( .A(n7865), .B(n7866), .Z(n4697) );
  IV U8153 ( .A(n7862), .Z(n7865) );
  XNOR U8154 ( .A(n4698), .B(n7862), .Z(n7864) );
  NAND U8155 ( .A(n7867), .B(e_input[739]), .Z(n4698) );
  NAND U8156 ( .A(n6112), .B(e_input[739]), .Z(n7867) );
  XOR U8157 ( .A(n7868), .B(n7869), .Z(n7862) );
  ANDN U8158 ( .A(n7870), .B(n4699), .Z(n7869) );
  XOR U8159 ( .A(n7871), .B(n7872), .Z(n4699) );
  IV U8160 ( .A(n7868), .Z(n7871) );
  XNOR U8161 ( .A(n4700), .B(n7868), .Z(n7870) );
  NAND U8162 ( .A(n7873), .B(e_input[738]), .Z(n4700) );
  NAND U8163 ( .A(n6112), .B(e_input[738]), .Z(n7873) );
  XOR U8164 ( .A(n7874), .B(n7875), .Z(n7868) );
  ANDN U8165 ( .A(n7876), .B(n4701), .Z(n7875) );
  XOR U8166 ( .A(n7877), .B(n7878), .Z(n4701) );
  IV U8167 ( .A(n7874), .Z(n7877) );
  XNOR U8168 ( .A(n4702), .B(n7874), .Z(n7876) );
  NAND U8169 ( .A(n7879), .B(e_input[737]), .Z(n4702) );
  NAND U8170 ( .A(n6112), .B(e_input[737]), .Z(n7879) );
  XOR U8171 ( .A(n7880), .B(n7881), .Z(n7874) );
  ANDN U8172 ( .A(n7882), .B(n4703), .Z(n7881) );
  XOR U8173 ( .A(n7883), .B(n7884), .Z(n4703) );
  IV U8174 ( .A(n7880), .Z(n7883) );
  XNOR U8175 ( .A(n4704), .B(n7880), .Z(n7882) );
  NAND U8176 ( .A(n7885), .B(e_input[736]), .Z(n4704) );
  NAND U8177 ( .A(n6112), .B(e_input[736]), .Z(n7885) );
  XOR U8178 ( .A(n7886), .B(n7887), .Z(n7880) );
  ANDN U8179 ( .A(n7888), .B(n4705), .Z(n7887) );
  XOR U8180 ( .A(n7889), .B(n7890), .Z(n4705) );
  IV U8181 ( .A(n7886), .Z(n7889) );
  XNOR U8182 ( .A(n4706), .B(n7886), .Z(n7888) );
  NAND U8183 ( .A(n7891), .B(e_input[735]), .Z(n4706) );
  NAND U8184 ( .A(n6112), .B(e_input[735]), .Z(n7891) );
  XOR U8185 ( .A(n7892), .B(n7893), .Z(n7886) );
  ANDN U8186 ( .A(n7894), .B(n4707), .Z(n7893) );
  XOR U8187 ( .A(n7895), .B(n7896), .Z(n4707) );
  IV U8188 ( .A(n7892), .Z(n7895) );
  XNOR U8189 ( .A(n4708), .B(n7892), .Z(n7894) );
  NAND U8190 ( .A(n7897), .B(e_input[734]), .Z(n4708) );
  NAND U8191 ( .A(n6112), .B(e_input[734]), .Z(n7897) );
  XOR U8192 ( .A(n7898), .B(n7899), .Z(n7892) );
  ANDN U8193 ( .A(n7900), .B(n4709), .Z(n7899) );
  XOR U8194 ( .A(n7901), .B(n7902), .Z(n4709) );
  IV U8195 ( .A(n7898), .Z(n7901) );
  XNOR U8196 ( .A(n4710), .B(n7898), .Z(n7900) );
  NAND U8197 ( .A(n7903), .B(e_input[733]), .Z(n4710) );
  NAND U8198 ( .A(n6112), .B(e_input[733]), .Z(n7903) );
  XOR U8199 ( .A(n7904), .B(n7905), .Z(n7898) );
  ANDN U8200 ( .A(n7906), .B(n4711), .Z(n7905) );
  XOR U8201 ( .A(n7907), .B(n7908), .Z(n4711) );
  IV U8202 ( .A(n7904), .Z(n7907) );
  XNOR U8203 ( .A(n4712), .B(n7904), .Z(n7906) );
  NAND U8204 ( .A(n7909), .B(e_input[732]), .Z(n4712) );
  NAND U8205 ( .A(n6112), .B(e_input[732]), .Z(n7909) );
  XOR U8206 ( .A(n7910), .B(n7911), .Z(n7904) );
  ANDN U8207 ( .A(n7912), .B(n4713), .Z(n7911) );
  XOR U8208 ( .A(n7913), .B(n7914), .Z(n4713) );
  IV U8209 ( .A(n7910), .Z(n7913) );
  XNOR U8210 ( .A(n4714), .B(n7910), .Z(n7912) );
  NAND U8211 ( .A(n7915), .B(e_input[731]), .Z(n4714) );
  NAND U8212 ( .A(n6112), .B(e_input[731]), .Z(n7915) );
  XOR U8213 ( .A(n7916), .B(n7917), .Z(n7910) );
  ANDN U8214 ( .A(n7918), .B(n4715), .Z(n7917) );
  XOR U8215 ( .A(n7919), .B(n7920), .Z(n4715) );
  IV U8216 ( .A(n7916), .Z(n7919) );
  XNOR U8217 ( .A(n4716), .B(n7916), .Z(n7918) );
  NAND U8218 ( .A(n7921), .B(e_input[730]), .Z(n4716) );
  NAND U8219 ( .A(n6112), .B(e_input[730]), .Z(n7921) );
  XOR U8220 ( .A(n7922), .B(n7923), .Z(n7916) );
  ANDN U8221 ( .A(n7924), .B(n4719), .Z(n7923) );
  XOR U8222 ( .A(n7925), .B(n7926), .Z(n4719) );
  IV U8223 ( .A(n7922), .Z(n7925) );
  XNOR U8224 ( .A(n4720), .B(n7922), .Z(n7924) );
  NAND U8225 ( .A(n7927), .B(e_input[729]), .Z(n4720) );
  NAND U8226 ( .A(n6112), .B(e_input[729]), .Z(n7927) );
  XOR U8227 ( .A(n7928), .B(n7929), .Z(n7922) );
  ANDN U8228 ( .A(n7930), .B(n4721), .Z(n7929) );
  XOR U8229 ( .A(n7931), .B(n7932), .Z(n4721) );
  IV U8230 ( .A(n7928), .Z(n7931) );
  XNOR U8231 ( .A(n4722), .B(n7928), .Z(n7930) );
  NAND U8232 ( .A(n7933), .B(e_input[728]), .Z(n4722) );
  NAND U8233 ( .A(n6112), .B(e_input[728]), .Z(n7933) );
  XOR U8234 ( .A(n7934), .B(n7935), .Z(n7928) );
  ANDN U8235 ( .A(n7936), .B(n4723), .Z(n7935) );
  XOR U8236 ( .A(n7937), .B(n7938), .Z(n4723) );
  IV U8237 ( .A(n7934), .Z(n7937) );
  XNOR U8238 ( .A(n4724), .B(n7934), .Z(n7936) );
  NAND U8239 ( .A(n7939), .B(e_input[727]), .Z(n4724) );
  NAND U8240 ( .A(n6112), .B(e_input[727]), .Z(n7939) );
  XOR U8241 ( .A(n7940), .B(n7941), .Z(n7934) );
  ANDN U8242 ( .A(n7942), .B(n4725), .Z(n7941) );
  XOR U8243 ( .A(n7943), .B(n7944), .Z(n4725) );
  IV U8244 ( .A(n7940), .Z(n7943) );
  XNOR U8245 ( .A(n4726), .B(n7940), .Z(n7942) );
  NAND U8246 ( .A(n7945), .B(e_input[726]), .Z(n4726) );
  NAND U8247 ( .A(n6112), .B(e_input[726]), .Z(n7945) );
  XOR U8248 ( .A(n7946), .B(n7947), .Z(n7940) );
  ANDN U8249 ( .A(n7948), .B(n4727), .Z(n7947) );
  XOR U8250 ( .A(n7949), .B(n7950), .Z(n4727) );
  IV U8251 ( .A(n7946), .Z(n7949) );
  XNOR U8252 ( .A(n4728), .B(n7946), .Z(n7948) );
  NAND U8253 ( .A(n7951), .B(e_input[725]), .Z(n4728) );
  NAND U8254 ( .A(n6112), .B(e_input[725]), .Z(n7951) );
  XOR U8255 ( .A(n7952), .B(n7953), .Z(n7946) );
  ANDN U8256 ( .A(n7954), .B(n4729), .Z(n7953) );
  XOR U8257 ( .A(n7955), .B(n7956), .Z(n4729) );
  IV U8258 ( .A(n7952), .Z(n7955) );
  XNOR U8259 ( .A(n4730), .B(n7952), .Z(n7954) );
  NAND U8260 ( .A(n7957), .B(e_input[724]), .Z(n4730) );
  NAND U8261 ( .A(n6112), .B(e_input[724]), .Z(n7957) );
  XOR U8262 ( .A(n7958), .B(n7959), .Z(n7952) );
  ANDN U8263 ( .A(n7960), .B(n4731), .Z(n7959) );
  XOR U8264 ( .A(n7961), .B(n7962), .Z(n4731) );
  IV U8265 ( .A(n7958), .Z(n7961) );
  XNOR U8266 ( .A(n4732), .B(n7958), .Z(n7960) );
  NAND U8267 ( .A(n7963), .B(e_input[723]), .Z(n4732) );
  NAND U8268 ( .A(n6112), .B(e_input[723]), .Z(n7963) );
  XOR U8269 ( .A(n7964), .B(n7965), .Z(n7958) );
  ANDN U8270 ( .A(n7966), .B(n4733), .Z(n7965) );
  XOR U8271 ( .A(n7967), .B(n7968), .Z(n4733) );
  IV U8272 ( .A(n7964), .Z(n7967) );
  XNOR U8273 ( .A(n4734), .B(n7964), .Z(n7966) );
  NAND U8274 ( .A(n7969), .B(e_input[722]), .Z(n4734) );
  NAND U8275 ( .A(n6112), .B(e_input[722]), .Z(n7969) );
  XOR U8276 ( .A(n7970), .B(n7971), .Z(n7964) );
  ANDN U8277 ( .A(n7972), .B(n4735), .Z(n7971) );
  XOR U8278 ( .A(n7973), .B(n7974), .Z(n4735) );
  IV U8279 ( .A(n7970), .Z(n7973) );
  XNOR U8280 ( .A(n4736), .B(n7970), .Z(n7972) );
  NAND U8281 ( .A(n7975), .B(e_input[721]), .Z(n4736) );
  NAND U8282 ( .A(n6112), .B(e_input[721]), .Z(n7975) );
  XOR U8283 ( .A(n7976), .B(n7977), .Z(n7970) );
  ANDN U8284 ( .A(n7978), .B(n4737), .Z(n7977) );
  XOR U8285 ( .A(n7979), .B(n7980), .Z(n4737) );
  IV U8286 ( .A(n7976), .Z(n7979) );
  XNOR U8287 ( .A(n4738), .B(n7976), .Z(n7978) );
  NAND U8288 ( .A(n7981), .B(e_input[720]), .Z(n4738) );
  NAND U8289 ( .A(n6112), .B(e_input[720]), .Z(n7981) );
  XOR U8290 ( .A(n7982), .B(n7983), .Z(n7976) );
  ANDN U8291 ( .A(n7984), .B(n4741), .Z(n7983) );
  XOR U8292 ( .A(n7985), .B(n7986), .Z(n4741) );
  IV U8293 ( .A(n7982), .Z(n7985) );
  XNOR U8294 ( .A(n4742), .B(n7982), .Z(n7984) );
  NAND U8295 ( .A(n7987), .B(e_input[719]), .Z(n4742) );
  NAND U8296 ( .A(n6112), .B(e_input[719]), .Z(n7987) );
  XOR U8297 ( .A(n7988), .B(n7989), .Z(n7982) );
  ANDN U8298 ( .A(n7990), .B(n4743), .Z(n7989) );
  XOR U8299 ( .A(n7991), .B(n7992), .Z(n4743) );
  IV U8300 ( .A(n7988), .Z(n7991) );
  XNOR U8301 ( .A(n4744), .B(n7988), .Z(n7990) );
  NAND U8302 ( .A(n7993), .B(e_input[718]), .Z(n4744) );
  NAND U8303 ( .A(n6112), .B(e_input[718]), .Z(n7993) );
  XOR U8304 ( .A(n7994), .B(n7995), .Z(n7988) );
  ANDN U8305 ( .A(n7996), .B(n4745), .Z(n7995) );
  XOR U8306 ( .A(n7997), .B(n7998), .Z(n4745) );
  IV U8307 ( .A(n7994), .Z(n7997) );
  XNOR U8308 ( .A(n4746), .B(n7994), .Z(n7996) );
  NAND U8309 ( .A(n7999), .B(e_input[717]), .Z(n4746) );
  NAND U8310 ( .A(n6112), .B(e_input[717]), .Z(n7999) );
  XOR U8311 ( .A(n8000), .B(n8001), .Z(n7994) );
  ANDN U8312 ( .A(n8002), .B(n4747), .Z(n8001) );
  XOR U8313 ( .A(n8003), .B(n8004), .Z(n4747) );
  IV U8314 ( .A(n8000), .Z(n8003) );
  XNOR U8315 ( .A(n4748), .B(n8000), .Z(n8002) );
  NAND U8316 ( .A(n8005), .B(e_input[716]), .Z(n4748) );
  NAND U8317 ( .A(n6112), .B(e_input[716]), .Z(n8005) );
  XOR U8318 ( .A(n8006), .B(n8007), .Z(n8000) );
  ANDN U8319 ( .A(n8008), .B(n4749), .Z(n8007) );
  XOR U8320 ( .A(n8009), .B(n8010), .Z(n4749) );
  IV U8321 ( .A(n8006), .Z(n8009) );
  XNOR U8322 ( .A(n4750), .B(n8006), .Z(n8008) );
  NAND U8323 ( .A(n8011), .B(e_input[715]), .Z(n4750) );
  NAND U8324 ( .A(n6112), .B(e_input[715]), .Z(n8011) );
  XOR U8325 ( .A(n8012), .B(n8013), .Z(n8006) );
  ANDN U8326 ( .A(n8014), .B(n4751), .Z(n8013) );
  XOR U8327 ( .A(n8015), .B(n8016), .Z(n4751) );
  IV U8328 ( .A(n8012), .Z(n8015) );
  XNOR U8329 ( .A(n4752), .B(n8012), .Z(n8014) );
  NAND U8330 ( .A(n8017), .B(e_input[714]), .Z(n4752) );
  NAND U8331 ( .A(n6112), .B(e_input[714]), .Z(n8017) );
  XOR U8332 ( .A(n8018), .B(n8019), .Z(n8012) );
  ANDN U8333 ( .A(n8020), .B(n4753), .Z(n8019) );
  XOR U8334 ( .A(n8021), .B(n8022), .Z(n4753) );
  IV U8335 ( .A(n8018), .Z(n8021) );
  XNOR U8336 ( .A(n4754), .B(n8018), .Z(n8020) );
  NAND U8337 ( .A(n8023), .B(e_input[713]), .Z(n4754) );
  NAND U8338 ( .A(n6112), .B(e_input[713]), .Z(n8023) );
  XOR U8339 ( .A(n8024), .B(n8025), .Z(n8018) );
  ANDN U8340 ( .A(n8026), .B(n4755), .Z(n8025) );
  XOR U8341 ( .A(n8027), .B(n8028), .Z(n4755) );
  IV U8342 ( .A(n8024), .Z(n8027) );
  XNOR U8343 ( .A(n4756), .B(n8024), .Z(n8026) );
  NAND U8344 ( .A(n8029), .B(e_input[712]), .Z(n4756) );
  NAND U8345 ( .A(n6112), .B(e_input[712]), .Z(n8029) );
  XOR U8346 ( .A(n8030), .B(n8031), .Z(n8024) );
  ANDN U8347 ( .A(n8032), .B(n4757), .Z(n8031) );
  XOR U8348 ( .A(n8033), .B(n8034), .Z(n4757) );
  IV U8349 ( .A(n8030), .Z(n8033) );
  XNOR U8350 ( .A(n4758), .B(n8030), .Z(n8032) );
  NAND U8351 ( .A(n8035), .B(e_input[711]), .Z(n4758) );
  NAND U8352 ( .A(n6112), .B(e_input[711]), .Z(n8035) );
  XOR U8353 ( .A(n8036), .B(n8037), .Z(n8030) );
  ANDN U8354 ( .A(n8038), .B(n4759), .Z(n8037) );
  XOR U8355 ( .A(n8039), .B(n8040), .Z(n4759) );
  IV U8356 ( .A(n8036), .Z(n8039) );
  XNOR U8357 ( .A(n4760), .B(n8036), .Z(n8038) );
  NAND U8358 ( .A(n8041), .B(e_input[710]), .Z(n4760) );
  NAND U8359 ( .A(n6112), .B(e_input[710]), .Z(n8041) );
  XOR U8360 ( .A(n8042), .B(n8043), .Z(n8036) );
  ANDN U8361 ( .A(n8044), .B(n4763), .Z(n8043) );
  XOR U8362 ( .A(n8045), .B(n8046), .Z(n4763) );
  IV U8363 ( .A(n8042), .Z(n8045) );
  XNOR U8364 ( .A(n4764), .B(n8042), .Z(n8044) );
  NAND U8365 ( .A(n8047), .B(e_input[709]), .Z(n4764) );
  NAND U8366 ( .A(n6112), .B(e_input[709]), .Z(n8047) );
  XOR U8367 ( .A(n8048), .B(n8049), .Z(n8042) );
  ANDN U8368 ( .A(n8050), .B(n4765), .Z(n8049) );
  XOR U8369 ( .A(n8051), .B(n8052), .Z(n4765) );
  IV U8370 ( .A(n8048), .Z(n8051) );
  XNOR U8371 ( .A(n4766), .B(n8048), .Z(n8050) );
  NAND U8372 ( .A(n8053), .B(e_input[708]), .Z(n4766) );
  NAND U8373 ( .A(n6112), .B(e_input[708]), .Z(n8053) );
  XOR U8374 ( .A(n8054), .B(n8055), .Z(n8048) );
  ANDN U8375 ( .A(n8056), .B(n4767), .Z(n8055) );
  XOR U8376 ( .A(n8057), .B(n8058), .Z(n4767) );
  IV U8377 ( .A(n8054), .Z(n8057) );
  XNOR U8378 ( .A(n4768), .B(n8054), .Z(n8056) );
  NAND U8379 ( .A(n8059), .B(e_input[707]), .Z(n4768) );
  NAND U8380 ( .A(n6112), .B(e_input[707]), .Z(n8059) );
  XOR U8381 ( .A(n8060), .B(n8061), .Z(n8054) );
  ANDN U8382 ( .A(n8062), .B(n4769), .Z(n8061) );
  XOR U8383 ( .A(n8063), .B(n8064), .Z(n4769) );
  IV U8384 ( .A(n8060), .Z(n8063) );
  XNOR U8385 ( .A(n4770), .B(n8060), .Z(n8062) );
  NAND U8386 ( .A(n8065), .B(e_input[706]), .Z(n4770) );
  NAND U8387 ( .A(n6112), .B(e_input[706]), .Z(n8065) );
  XOR U8388 ( .A(n8066), .B(n8067), .Z(n8060) );
  ANDN U8389 ( .A(n8068), .B(n4771), .Z(n8067) );
  XOR U8390 ( .A(n8069), .B(n8070), .Z(n4771) );
  IV U8391 ( .A(n8066), .Z(n8069) );
  XNOR U8392 ( .A(n4772), .B(n8066), .Z(n8068) );
  NAND U8393 ( .A(n8071), .B(e_input[705]), .Z(n4772) );
  NAND U8394 ( .A(n6112), .B(e_input[705]), .Z(n8071) );
  XOR U8395 ( .A(n8072), .B(n8073), .Z(n8066) );
  ANDN U8396 ( .A(n8074), .B(n4773), .Z(n8073) );
  XOR U8397 ( .A(n8075), .B(n8076), .Z(n4773) );
  IV U8398 ( .A(n8072), .Z(n8075) );
  XNOR U8399 ( .A(n4774), .B(n8072), .Z(n8074) );
  NAND U8400 ( .A(n8077), .B(e_input[704]), .Z(n4774) );
  NAND U8401 ( .A(n6112), .B(e_input[704]), .Z(n8077) );
  XOR U8402 ( .A(n8078), .B(n8079), .Z(n8072) );
  ANDN U8403 ( .A(n8080), .B(n4775), .Z(n8079) );
  XOR U8404 ( .A(n8081), .B(n8082), .Z(n4775) );
  IV U8405 ( .A(n8078), .Z(n8081) );
  XNOR U8406 ( .A(n4776), .B(n8078), .Z(n8080) );
  NAND U8407 ( .A(n8083), .B(e_input[703]), .Z(n4776) );
  NAND U8408 ( .A(n6112), .B(e_input[703]), .Z(n8083) );
  XOR U8409 ( .A(n8084), .B(n8085), .Z(n8078) );
  ANDN U8410 ( .A(n8086), .B(n4777), .Z(n8085) );
  XOR U8411 ( .A(n8087), .B(n8088), .Z(n4777) );
  IV U8412 ( .A(n8084), .Z(n8087) );
  XNOR U8413 ( .A(n4778), .B(n8084), .Z(n8086) );
  NAND U8414 ( .A(n8089), .B(e_input[702]), .Z(n4778) );
  NAND U8415 ( .A(n6112), .B(e_input[702]), .Z(n8089) );
  XOR U8416 ( .A(n8090), .B(n8091), .Z(n8084) );
  ANDN U8417 ( .A(n8092), .B(n4779), .Z(n8091) );
  XOR U8418 ( .A(n8093), .B(n8094), .Z(n4779) );
  IV U8419 ( .A(n8090), .Z(n8093) );
  XNOR U8420 ( .A(n4780), .B(n8090), .Z(n8092) );
  NAND U8421 ( .A(n8095), .B(e_input[701]), .Z(n4780) );
  NAND U8422 ( .A(n6112), .B(e_input[701]), .Z(n8095) );
  XOR U8423 ( .A(n8096), .B(n8097), .Z(n8090) );
  ANDN U8424 ( .A(n8098), .B(n4781), .Z(n8097) );
  XOR U8425 ( .A(n8099), .B(n8100), .Z(n4781) );
  IV U8426 ( .A(n8096), .Z(n8099) );
  XNOR U8427 ( .A(n4782), .B(n8096), .Z(n8098) );
  NAND U8428 ( .A(n8101), .B(e_input[700]), .Z(n4782) );
  NAND U8429 ( .A(n6112), .B(e_input[700]), .Z(n8101) );
  XOR U8430 ( .A(n8102), .B(n8103), .Z(n8096) );
  ANDN U8431 ( .A(n8104), .B(n4787), .Z(n8103) );
  XOR U8432 ( .A(n8105), .B(n8106), .Z(n4787) );
  IV U8433 ( .A(n8102), .Z(n8105) );
  XNOR U8434 ( .A(n4788), .B(n8102), .Z(n8104) );
  NAND U8435 ( .A(n8107), .B(e_input[699]), .Z(n4788) );
  NAND U8436 ( .A(n6112), .B(e_input[699]), .Z(n8107) );
  XOR U8437 ( .A(n8108), .B(n8109), .Z(n8102) );
  ANDN U8438 ( .A(n8110), .B(n4789), .Z(n8109) );
  XOR U8439 ( .A(n8111), .B(n8112), .Z(n4789) );
  IV U8440 ( .A(n8108), .Z(n8111) );
  XNOR U8441 ( .A(n4790), .B(n8108), .Z(n8110) );
  NAND U8442 ( .A(n8113), .B(e_input[698]), .Z(n4790) );
  NAND U8443 ( .A(n6112), .B(e_input[698]), .Z(n8113) );
  XOR U8444 ( .A(n8114), .B(n8115), .Z(n8108) );
  ANDN U8445 ( .A(n8116), .B(n4791), .Z(n8115) );
  XOR U8446 ( .A(n8117), .B(n8118), .Z(n4791) );
  IV U8447 ( .A(n8114), .Z(n8117) );
  XNOR U8448 ( .A(n4792), .B(n8114), .Z(n8116) );
  NAND U8449 ( .A(n8119), .B(e_input[697]), .Z(n4792) );
  NAND U8450 ( .A(n6112), .B(e_input[697]), .Z(n8119) );
  XOR U8451 ( .A(n8120), .B(n8121), .Z(n8114) );
  ANDN U8452 ( .A(n8122), .B(n4793), .Z(n8121) );
  XOR U8453 ( .A(n8123), .B(n8124), .Z(n4793) );
  IV U8454 ( .A(n8120), .Z(n8123) );
  XNOR U8455 ( .A(n4794), .B(n8120), .Z(n8122) );
  NAND U8456 ( .A(n8125), .B(e_input[696]), .Z(n4794) );
  NAND U8457 ( .A(n6112), .B(e_input[696]), .Z(n8125) );
  XOR U8458 ( .A(n8126), .B(n8127), .Z(n8120) );
  ANDN U8459 ( .A(n8128), .B(n4795), .Z(n8127) );
  XOR U8460 ( .A(n8129), .B(n8130), .Z(n4795) );
  IV U8461 ( .A(n8126), .Z(n8129) );
  XNOR U8462 ( .A(n4796), .B(n8126), .Z(n8128) );
  NAND U8463 ( .A(n8131), .B(e_input[695]), .Z(n4796) );
  NAND U8464 ( .A(n6112), .B(e_input[695]), .Z(n8131) );
  XOR U8465 ( .A(n8132), .B(n8133), .Z(n8126) );
  ANDN U8466 ( .A(n8134), .B(n4797), .Z(n8133) );
  XOR U8467 ( .A(n8135), .B(n8136), .Z(n4797) );
  IV U8468 ( .A(n8132), .Z(n8135) );
  XNOR U8469 ( .A(n4798), .B(n8132), .Z(n8134) );
  NAND U8470 ( .A(n8137), .B(e_input[694]), .Z(n4798) );
  NAND U8471 ( .A(n6112), .B(e_input[694]), .Z(n8137) );
  XOR U8472 ( .A(n8138), .B(n8139), .Z(n8132) );
  ANDN U8473 ( .A(n8140), .B(n4799), .Z(n8139) );
  XOR U8474 ( .A(n8141), .B(n8142), .Z(n4799) );
  IV U8475 ( .A(n8138), .Z(n8141) );
  XNOR U8476 ( .A(n4800), .B(n8138), .Z(n8140) );
  NAND U8477 ( .A(n8143), .B(e_input[693]), .Z(n4800) );
  NAND U8478 ( .A(n6112), .B(e_input[693]), .Z(n8143) );
  XOR U8479 ( .A(n8144), .B(n8145), .Z(n8138) );
  ANDN U8480 ( .A(n8146), .B(n4801), .Z(n8145) );
  XOR U8481 ( .A(n8147), .B(n8148), .Z(n4801) );
  IV U8482 ( .A(n8144), .Z(n8147) );
  XNOR U8483 ( .A(n4802), .B(n8144), .Z(n8146) );
  NAND U8484 ( .A(n8149), .B(e_input[692]), .Z(n4802) );
  NAND U8485 ( .A(n6112), .B(e_input[692]), .Z(n8149) );
  XOR U8486 ( .A(n8150), .B(n8151), .Z(n8144) );
  ANDN U8487 ( .A(n8152), .B(n4803), .Z(n8151) );
  XOR U8488 ( .A(n8153), .B(n8154), .Z(n4803) );
  IV U8489 ( .A(n8150), .Z(n8153) );
  XNOR U8490 ( .A(n4804), .B(n8150), .Z(n8152) );
  NAND U8491 ( .A(n8155), .B(e_input[691]), .Z(n4804) );
  NAND U8492 ( .A(n6112), .B(e_input[691]), .Z(n8155) );
  XOR U8493 ( .A(n8156), .B(n8157), .Z(n8150) );
  ANDN U8494 ( .A(n8158), .B(n4805), .Z(n8157) );
  XOR U8495 ( .A(n8159), .B(n8160), .Z(n4805) );
  IV U8496 ( .A(n8156), .Z(n8159) );
  XNOR U8497 ( .A(n4806), .B(n8156), .Z(n8158) );
  NAND U8498 ( .A(n8161), .B(e_input[690]), .Z(n4806) );
  NAND U8499 ( .A(n6112), .B(e_input[690]), .Z(n8161) );
  XOR U8500 ( .A(n8162), .B(n8163), .Z(n8156) );
  ANDN U8501 ( .A(n8164), .B(n4809), .Z(n8163) );
  XOR U8502 ( .A(n8165), .B(n8166), .Z(n4809) );
  IV U8503 ( .A(n8162), .Z(n8165) );
  XNOR U8504 ( .A(n4810), .B(n8162), .Z(n8164) );
  NAND U8505 ( .A(n8167), .B(e_input[689]), .Z(n4810) );
  NAND U8506 ( .A(n6112), .B(e_input[689]), .Z(n8167) );
  XOR U8507 ( .A(n8168), .B(n8169), .Z(n8162) );
  ANDN U8508 ( .A(n8170), .B(n4811), .Z(n8169) );
  XOR U8509 ( .A(n8171), .B(n8172), .Z(n4811) );
  IV U8510 ( .A(n8168), .Z(n8171) );
  XNOR U8511 ( .A(n4812), .B(n8168), .Z(n8170) );
  NAND U8512 ( .A(n8173), .B(e_input[688]), .Z(n4812) );
  NAND U8513 ( .A(n6112), .B(e_input[688]), .Z(n8173) );
  XOR U8514 ( .A(n8174), .B(n8175), .Z(n8168) );
  ANDN U8515 ( .A(n8176), .B(n4813), .Z(n8175) );
  XOR U8516 ( .A(n8177), .B(n8178), .Z(n4813) );
  IV U8517 ( .A(n8174), .Z(n8177) );
  XNOR U8518 ( .A(n4814), .B(n8174), .Z(n8176) );
  NAND U8519 ( .A(n8179), .B(e_input[687]), .Z(n4814) );
  NAND U8520 ( .A(n6112), .B(e_input[687]), .Z(n8179) );
  XOR U8521 ( .A(n8180), .B(n8181), .Z(n8174) );
  ANDN U8522 ( .A(n8182), .B(n4815), .Z(n8181) );
  XOR U8523 ( .A(n8183), .B(n8184), .Z(n4815) );
  IV U8524 ( .A(n8180), .Z(n8183) );
  XNOR U8525 ( .A(n4816), .B(n8180), .Z(n8182) );
  NAND U8526 ( .A(n8185), .B(e_input[686]), .Z(n4816) );
  NAND U8527 ( .A(n6112), .B(e_input[686]), .Z(n8185) );
  XOR U8528 ( .A(n8186), .B(n8187), .Z(n8180) );
  ANDN U8529 ( .A(n8188), .B(n4817), .Z(n8187) );
  XOR U8530 ( .A(n8189), .B(n8190), .Z(n4817) );
  IV U8531 ( .A(n8186), .Z(n8189) );
  XNOR U8532 ( .A(n4818), .B(n8186), .Z(n8188) );
  NAND U8533 ( .A(n8191), .B(e_input[685]), .Z(n4818) );
  NAND U8534 ( .A(n6112), .B(e_input[685]), .Z(n8191) );
  XOR U8535 ( .A(n8192), .B(n8193), .Z(n8186) );
  ANDN U8536 ( .A(n8194), .B(n4819), .Z(n8193) );
  XOR U8537 ( .A(n8195), .B(n8196), .Z(n4819) );
  IV U8538 ( .A(n8192), .Z(n8195) );
  XNOR U8539 ( .A(n4820), .B(n8192), .Z(n8194) );
  NAND U8540 ( .A(n8197), .B(e_input[684]), .Z(n4820) );
  NAND U8541 ( .A(n6112), .B(e_input[684]), .Z(n8197) );
  XOR U8542 ( .A(n8198), .B(n8199), .Z(n8192) );
  ANDN U8543 ( .A(n8200), .B(n4821), .Z(n8199) );
  XOR U8544 ( .A(n8201), .B(n8202), .Z(n4821) );
  IV U8545 ( .A(n8198), .Z(n8201) );
  XNOR U8546 ( .A(n4822), .B(n8198), .Z(n8200) );
  NAND U8547 ( .A(n8203), .B(e_input[683]), .Z(n4822) );
  NAND U8548 ( .A(n6112), .B(e_input[683]), .Z(n8203) );
  XOR U8549 ( .A(n8204), .B(n8205), .Z(n8198) );
  ANDN U8550 ( .A(n8206), .B(n4823), .Z(n8205) );
  XOR U8551 ( .A(n8207), .B(n8208), .Z(n4823) );
  IV U8552 ( .A(n8204), .Z(n8207) );
  XNOR U8553 ( .A(n4824), .B(n8204), .Z(n8206) );
  NAND U8554 ( .A(n8209), .B(e_input[682]), .Z(n4824) );
  NAND U8555 ( .A(n6112), .B(e_input[682]), .Z(n8209) );
  XOR U8556 ( .A(n8210), .B(n8211), .Z(n8204) );
  ANDN U8557 ( .A(n8212), .B(n4825), .Z(n8211) );
  XOR U8558 ( .A(n8213), .B(n8214), .Z(n4825) );
  IV U8559 ( .A(n8210), .Z(n8213) );
  XNOR U8560 ( .A(n4826), .B(n8210), .Z(n8212) );
  NAND U8561 ( .A(n8215), .B(e_input[681]), .Z(n4826) );
  NAND U8562 ( .A(n6112), .B(e_input[681]), .Z(n8215) );
  XOR U8563 ( .A(n8216), .B(n8217), .Z(n8210) );
  ANDN U8564 ( .A(n8218), .B(n4827), .Z(n8217) );
  XOR U8565 ( .A(n8219), .B(n8220), .Z(n4827) );
  IV U8566 ( .A(n8216), .Z(n8219) );
  XNOR U8567 ( .A(n4828), .B(n8216), .Z(n8218) );
  NAND U8568 ( .A(n8221), .B(e_input[680]), .Z(n4828) );
  NAND U8569 ( .A(n6112), .B(e_input[680]), .Z(n8221) );
  XOR U8570 ( .A(n8222), .B(n8223), .Z(n8216) );
  ANDN U8571 ( .A(n8224), .B(n4831), .Z(n8223) );
  XOR U8572 ( .A(n8225), .B(n8226), .Z(n4831) );
  IV U8573 ( .A(n8222), .Z(n8225) );
  XNOR U8574 ( .A(n4832), .B(n8222), .Z(n8224) );
  NAND U8575 ( .A(n8227), .B(e_input[679]), .Z(n4832) );
  NAND U8576 ( .A(n6112), .B(e_input[679]), .Z(n8227) );
  XOR U8577 ( .A(n8228), .B(n8229), .Z(n8222) );
  ANDN U8578 ( .A(n8230), .B(n4833), .Z(n8229) );
  XOR U8579 ( .A(n8231), .B(n8232), .Z(n4833) );
  IV U8580 ( .A(n8228), .Z(n8231) );
  XNOR U8581 ( .A(n4834), .B(n8228), .Z(n8230) );
  NAND U8582 ( .A(n8233), .B(e_input[678]), .Z(n4834) );
  NAND U8583 ( .A(n6112), .B(e_input[678]), .Z(n8233) );
  XOR U8584 ( .A(n8234), .B(n8235), .Z(n8228) );
  ANDN U8585 ( .A(n8236), .B(n4835), .Z(n8235) );
  XOR U8586 ( .A(n8237), .B(n8238), .Z(n4835) );
  IV U8587 ( .A(n8234), .Z(n8237) );
  XNOR U8588 ( .A(n4836), .B(n8234), .Z(n8236) );
  NAND U8589 ( .A(n8239), .B(e_input[677]), .Z(n4836) );
  NAND U8590 ( .A(n6112), .B(e_input[677]), .Z(n8239) );
  XOR U8591 ( .A(n8240), .B(n8241), .Z(n8234) );
  ANDN U8592 ( .A(n8242), .B(n4837), .Z(n8241) );
  XOR U8593 ( .A(n8243), .B(n8244), .Z(n4837) );
  IV U8594 ( .A(n8240), .Z(n8243) );
  XNOR U8595 ( .A(n4838), .B(n8240), .Z(n8242) );
  NAND U8596 ( .A(n8245), .B(e_input[676]), .Z(n4838) );
  NAND U8597 ( .A(n6112), .B(e_input[676]), .Z(n8245) );
  XOR U8598 ( .A(n8246), .B(n8247), .Z(n8240) );
  ANDN U8599 ( .A(n8248), .B(n4839), .Z(n8247) );
  XOR U8600 ( .A(n8249), .B(n8250), .Z(n4839) );
  IV U8601 ( .A(n8246), .Z(n8249) );
  XNOR U8602 ( .A(n4840), .B(n8246), .Z(n8248) );
  NAND U8603 ( .A(n8251), .B(e_input[675]), .Z(n4840) );
  NAND U8604 ( .A(n6112), .B(e_input[675]), .Z(n8251) );
  XOR U8605 ( .A(n8252), .B(n8253), .Z(n8246) );
  ANDN U8606 ( .A(n8254), .B(n4841), .Z(n8253) );
  XOR U8607 ( .A(n8255), .B(n8256), .Z(n4841) );
  IV U8608 ( .A(n8252), .Z(n8255) );
  XNOR U8609 ( .A(n4842), .B(n8252), .Z(n8254) );
  NAND U8610 ( .A(n8257), .B(e_input[674]), .Z(n4842) );
  NAND U8611 ( .A(n6112), .B(e_input[674]), .Z(n8257) );
  XOR U8612 ( .A(n8258), .B(n8259), .Z(n8252) );
  ANDN U8613 ( .A(n8260), .B(n4843), .Z(n8259) );
  XOR U8614 ( .A(n8261), .B(n8262), .Z(n4843) );
  IV U8615 ( .A(n8258), .Z(n8261) );
  XNOR U8616 ( .A(n4844), .B(n8258), .Z(n8260) );
  NAND U8617 ( .A(n8263), .B(e_input[673]), .Z(n4844) );
  NAND U8618 ( .A(n6112), .B(e_input[673]), .Z(n8263) );
  XOR U8619 ( .A(n8264), .B(n8265), .Z(n8258) );
  ANDN U8620 ( .A(n8266), .B(n4845), .Z(n8265) );
  XOR U8621 ( .A(n8267), .B(n8268), .Z(n4845) );
  IV U8622 ( .A(n8264), .Z(n8267) );
  XNOR U8623 ( .A(n4846), .B(n8264), .Z(n8266) );
  NAND U8624 ( .A(n8269), .B(e_input[672]), .Z(n4846) );
  NAND U8625 ( .A(n6112), .B(e_input[672]), .Z(n8269) );
  XOR U8626 ( .A(n8270), .B(n8271), .Z(n8264) );
  ANDN U8627 ( .A(n8272), .B(n4847), .Z(n8271) );
  XOR U8628 ( .A(n8273), .B(n8274), .Z(n4847) );
  IV U8629 ( .A(n8270), .Z(n8273) );
  XNOR U8630 ( .A(n4848), .B(n8270), .Z(n8272) );
  NAND U8631 ( .A(n8275), .B(e_input[671]), .Z(n4848) );
  NAND U8632 ( .A(n6112), .B(e_input[671]), .Z(n8275) );
  XOR U8633 ( .A(n8276), .B(n8277), .Z(n8270) );
  ANDN U8634 ( .A(n8278), .B(n4849), .Z(n8277) );
  XOR U8635 ( .A(n8279), .B(n8280), .Z(n4849) );
  IV U8636 ( .A(n8276), .Z(n8279) );
  XNOR U8637 ( .A(n4850), .B(n8276), .Z(n8278) );
  NAND U8638 ( .A(n8281), .B(e_input[670]), .Z(n4850) );
  NAND U8639 ( .A(n6112), .B(e_input[670]), .Z(n8281) );
  XOR U8640 ( .A(n8282), .B(n8283), .Z(n8276) );
  ANDN U8641 ( .A(n8284), .B(n4853), .Z(n8283) );
  XOR U8642 ( .A(n8285), .B(n8286), .Z(n4853) );
  IV U8643 ( .A(n8282), .Z(n8285) );
  XNOR U8644 ( .A(n4854), .B(n8282), .Z(n8284) );
  NAND U8645 ( .A(n8287), .B(e_input[669]), .Z(n4854) );
  NAND U8646 ( .A(n6112), .B(e_input[669]), .Z(n8287) );
  XOR U8647 ( .A(n8288), .B(n8289), .Z(n8282) );
  ANDN U8648 ( .A(n8290), .B(n4855), .Z(n8289) );
  XOR U8649 ( .A(n8291), .B(n8292), .Z(n4855) );
  IV U8650 ( .A(n8288), .Z(n8291) );
  XNOR U8651 ( .A(n4856), .B(n8288), .Z(n8290) );
  NAND U8652 ( .A(n8293), .B(e_input[668]), .Z(n4856) );
  NAND U8653 ( .A(n6112), .B(e_input[668]), .Z(n8293) );
  XOR U8654 ( .A(n8294), .B(n8295), .Z(n8288) );
  ANDN U8655 ( .A(n8296), .B(n4857), .Z(n8295) );
  XOR U8656 ( .A(n8297), .B(n8298), .Z(n4857) );
  IV U8657 ( .A(n8294), .Z(n8297) );
  XNOR U8658 ( .A(n4858), .B(n8294), .Z(n8296) );
  NAND U8659 ( .A(n8299), .B(e_input[667]), .Z(n4858) );
  NAND U8660 ( .A(n6112), .B(e_input[667]), .Z(n8299) );
  XOR U8661 ( .A(n8300), .B(n8301), .Z(n8294) );
  ANDN U8662 ( .A(n8302), .B(n4859), .Z(n8301) );
  XOR U8663 ( .A(n8303), .B(n8304), .Z(n4859) );
  IV U8664 ( .A(n8300), .Z(n8303) );
  XNOR U8665 ( .A(n4860), .B(n8300), .Z(n8302) );
  NAND U8666 ( .A(n8305), .B(e_input[666]), .Z(n4860) );
  NAND U8667 ( .A(n6112), .B(e_input[666]), .Z(n8305) );
  XOR U8668 ( .A(n8306), .B(n8307), .Z(n8300) );
  ANDN U8669 ( .A(n8308), .B(n4861), .Z(n8307) );
  XOR U8670 ( .A(n8309), .B(n8310), .Z(n4861) );
  IV U8671 ( .A(n8306), .Z(n8309) );
  XNOR U8672 ( .A(n4862), .B(n8306), .Z(n8308) );
  NAND U8673 ( .A(n8311), .B(e_input[665]), .Z(n4862) );
  NAND U8674 ( .A(n6112), .B(e_input[665]), .Z(n8311) );
  XOR U8675 ( .A(n8312), .B(n8313), .Z(n8306) );
  ANDN U8676 ( .A(n8314), .B(n4863), .Z(n8313) );
  XOR U8677 ( .A(n8315), .B(n8316), .Z(n4863) );
  IV U8678 ( .A(n8312), .Z(n8315) );
  XNOR U8679 ( .A(n4864), .B(n8312), .Z(n8314) );
  NAND U8680 ( .A(n8317), .B(e_input[664]), .Z(n4864) );
  NAND U8681 ( .A(n6112), .B(e_input[664]), .Z(n8317) );
  XOR U8682 ( .A(n8318), .B(n8319), .Z(n8312) );
  ANDN U8683 ( .A(n8320), .B(n4865), .Z(n8319) );
  XOR U8684 ( .A(n8321), .B(n8322), .Z(n4865) );
  IV U8685 ( .A(n8318), .Z(n8321) );
  XNOR U8686 ( .A(n4866), .B(n8318), .Z(n8320) );
  NAND U8687 ( .A(n8323), .B(e_input[663]), .Z(n4866) );
  NAND U8688 ( .A(n6112), .B(e_input[663]), .Z(n8323) );
  XOR U8689 ( .A(n8324), .B(n8325), .Z(n8318) );
  ANDN U8690 ( .A(n8326), .B(n4867), .Z(n8325) );
  XOR U8691 ( .A(n8327), .B(n8328), .Z(n4867) );
  IV U8692 ( .A(n8324), .Z(n8327) );
  XNOR U8693 ( .A(n4868), .B(n8324), .Z(n8326) );
  NAND U8694 ( .A(n8329), .B(e_input[662]), .Z(n4868) );
  NAND U8695 ( .A(n6112), .B(e_input[662]), .Z(n8329) );
  XOR U8696 ( .A(n8330), .B(n8331), .Z(n8324) );
  ANDN U8697 ( .A(n8332), .B(n4869), .Z(n8331) );
  XOR U8698 ( .A(n8333), .B(n8334), .Z(n4869) );
  IV U8699 ( .A(n8330), .Z(n8333) );
  XNOR U8700 ( .A(n4870), .B(n8330), .Z(n8332) );
  NAND U8701 ( .A(n8335), .B(e_input[661]), .Z(n4870) );
  NAND U8702 ( .A(n6112), .B(e_input[661]), .Z(n8335) );
  XOR U8703 ( .A(n8336), .B(n8337), .Z(n8330) );
  ANDN U8704 ( .A(n8338), .B(n4871), .Z(n8337) );
  XOR U8705 ( .A(n8339), .B(n8340), .Z(n4871) );
  IV U8706 ( .A(n8336), .Z(n8339) );
  XNOR U8707 ( .A(n4872), .B(n8336), .Z(n8338) );
  NAND U8708 ( .A(n8341), .B(e_input[660]), .Z(n4872) );
  NAND U8709 ( .A(n6112), .B(e_input[660]), .Z(n8341) );
  XOR U8710 ( .A(n8342), .B(n8343), .Z(n8336) );
  ANDN U8711 ( .A(n8344), .B(n4875), .Z(n8343) );
  XOR U8712 ( .A(n8345), .B(n8346), .Z(n4875) );
  IV U8713 ( .A(n8342), .Z(n8345) );
  XNOR U8714 ( .A(n4876), .B(n8342), .Z(n8344) );
  NAND U8715 ( .A(n8347), .B(e_input[659]), .Z(n4876) );
  NAND U8716 ( .A(n6112), .B(e_input[659]), .Z(n8347) );
  XOR U8717 ( .A(n8348), .B(n8349), .Z(n8342) );
  ANDN U8718 ( .A(n8350), .B(n4877), .Z(n8349) );
  XOR U8719 ( .A(n8351), .B(n8352), .Z(n4877) );
  IV U8720 ( .A(n8348), .Z(n8351) );
  XNOR U8721 ( .A(n4878), .B(n8348), .Z(n8350) );
  NAND U8722 ( .A(n8353), .B(e_input[658]), .Z(n4878) );
  NAND U8723 ( .A(n6112), .B(e_input[658]), .Z(n8353) );
  XOR U8724 ( .A(n8354), .B(n8355), .Z(n8348) );
  ANDN U8725 ( .A(n8356), .B(n4879), .Z(n8355) );
  XOR U8726 ( .A(n8357), .B(n8358), .Z(n4879) );
  IV U8727 ( .A(n8354), .Z(n8357) );
  XNOR U8728 ( .A(n4880), .B(n8354), .Z(n8356) );
  NAND U8729 ( .A(n8359), .B(e_input[657]), .Z(n4880) );
  NAND U8730 ( .A(n6112), .B(e_input[657]), .Z(n8359) );
  XOR U8731 ( .A(n8360), .B(n8361), .Z(n8354) );
  ANDN U8732 ( .A(n8362), .B(n4881), .Z(n8361) );
  XOR U8733 ( .A(n8363), .B(n8364), .Z(n4881) );
  IV U8734 ( .A(n8360), .Z(n8363) );
  XNOR U8735 ( .A(n4882), .B(n8360), .Z(n8362) );
  NAND U8736 ( .A(n8365), .B(e_input[656]), .Z(n4882) );
  NAND U8737 ( .A(n6112), .B(e_input[656]), .Z(n8365) );
  XOR U8738 ( .A(n8366), .B(n8367), .Z(n8360) );
  ANDN U8739 ( .A(n8368), .B(n4883), .Z(n8367) );
  XOR U8740 ( .A(n8369), .B(n8370), .Z(n4883) );
  IV U8741 ( .A(n8366), .Z(n8369) );
  XNOR U8742 ( .A(n4884), .B(n8366), .Z(n8368) );
  NAND U8743 ( .A(n8371), .B(e_input[655]), .Z(n4884) );
  NAND U8744 ( .A(n6112), .B(e_input[655]), .Z(n8371) );
  XOR U8745 ( .A(n8372), .B(n8373), .Z(n8366) );
  ANDN U8746 ( .A(n8374), .B(n4885), .Z(n8373) );
  XOR U8747 ( .A(n8375), .B(n8376), .Z(n4885) );
  IV U8748 ( .A(n8372), .Z(n8375) );
  XNOR U8749 ( .A(n4886), .B(n8372), .Z(n8374) );
  NAND U8750 ( .A(n8377), .B(e_input[654]), .Z(n4886) );
  NAND U8751 ( .A(n6112), .B(e_input[654]), .Z(n8377) );
  XOR U8752 ( .A(n8378), .B(n8379), .Z(n8372) );
  ANDN U8753 ( .A(n8380), .B(n4887), .Z(n8379) );
  XOR U8754 ( .A(n8381), .B(n8382), .Z(n4887) );
  IV U8755 ( .A(n8378), .Z(n8381) );
  XNOR U8756 ( .A(n4888), .B(n8378), .Z(n8380) );
  NAND U8757 ( .A(n8383), .B(e_input[653]), .Z(n4888) );
  NAND U8758 ( .A(n6112), .B(e_input[653]), .Z(n8383) );
  XOR U8759 ( .A(n8384), .B(n8385), .Z(n8378) );
  ANDN U8760 ( .A(n8386), .B(n4889), .Z(n8385) );
  XOR U8761 ( .A(n8387), .B(n8388), .Z(n4889) );
  IV U8762 ( .A(n8384), .Z(n8387) );
  XNOR U8763 ( .A(n4890), .B(n8384), .Z(n8386) );
  NAND U8764 ( .A(n8389), .B(e_input[652]), .Z(n4890) );
  NAND U8765 ( .A(n6112), .B(e_input[652]), .Z(n8389) );
  XOR U8766 ( .A(n8390), .B(n8391), .Z(n8384) );
  ANDN U8767 ( .A(n8392), .B(n4891), .Z(n8391) );
  XOR U8768 ( .A(n8393), .B(n8394), .Z(n4891) );
  IV U8769 ( .A(n8390), .Z(n8393) );
  XNOR U8770 ( .A(n4892), .B(n8390), .Z(n8392) );
  NAND U8771 ( .A(n8395), .B(e_input[651]), .Z(n4892) );
  NAND U8772 ( .A(n6112), .B(e_input[651]), .Z(n8395) );
  XOR U8773 ( .A(n8396), .B(n8397), .Z(n8390) );
  ANDN U8774 ( .A(n8398), .B(n4893), .Z(n8397) );
  XOR U8775 ( .A(n8399), .B(n8400), .Z(n4893) );
  IV U8776 ( .A(n8396), .Z(n8399) );
  XNOR U8777 ( .A(n4894), .B(n8396), .Z(n8398) );
  NAND U8778 ( .A(n8401), .B(e_input[650]), .Z(n4894) );
  NAND U8779 ( .A(n6112), .B(e_input[650]), .Z(n8401) );
  XOR U8780 ( .A(n8402), .B(n8403), .Z(n8396) );
  ANDN U8781 ( .A(n8404), .B(n4897), .Z(n8403) );
  XOR U8782 ( .A(n8405), .B(n8406), .Z(n4897) );
  IV U8783 ( .A(n8402), .Z(n8405) );
  XNOR U8784 ( .A(n4898), .B(n8402), .Z(n8404) );
  NAND U8785 ( .A(n8407), .B(e_input[649]), .Z(n4898) );
  NAND U8786 ( .A(n6112), .B(e_input[649]), .Z(n8407) );
  XOR U8787 ( .A(n8408), .B(n8409), .Z(n8402) );
  ANDN U8788 ( .A(n8410), .B(n4899), .Z(n8409) );
  XOR U8789 ( .A(n8411), .B(n8412), .Z(n4899) );
  IV U8790 ( .A(n8408), .Z(n8411) );
  XNOR U8791 ( .A(n4900), .B(n8408), .Z(n8410) );
  NAND U8792 ( .A(n8413), .B(e_input[648]), .Z(n4900) );
  NAND U8793 ( .A(n6112), .B(e_input[648]), .Z(n8413) );
  XOR U8794 ( .A(n8414), .B(n8415), .Z(n8408) );
  ANDN U8795 ( .A(n8416), .B(n4901), .Z(n8415) );
  XOR U8796 ( .A(n8417), .B(n8418), .Z(n4901) );
  IV U8797 ( .A(n8414), .Z(n8417) );
  XNOR U8798 ( .A(n4902), .B(n8414), .Z(n8416) );
  NAND U8799 ( .A(n8419), .B(e_input[647]), .Z(n4902) );
  NAND U8800 ( .A(n6112), .B(e_input[647]), .Z(n8419) );
  XOR U8801 ( .A(n8420), .B(n8421), .Z(n8414) );
  ANDN U8802 ( .A(n8422), .B(n4903), .Z(n8421) );
  XOR U8803 ( .A(n8423), .B(n8424), .Z(n4903) );
  IV U8804 ( .A(n8420), .Z(n8423) );
  XNOR U8805 ( .A(n4904), .B(n8420), .Z(n8422) );
  NAND U8806 ( .A(n8425), .B(e_input[646]), .Z(n4904) );
  NAND U8807 ( .A(n6112), .B(e_input[646]), .Z(n8425) );
  XOR U8808 ( .A(n8426), .B(n8427), .Z(n8420) );
  ANDN U8809 ( .A(n8428), .B(n4905), .Z(n8427) );
  XOR U8810 ( .A(n8429), .B(n8430), .Z(n4905) );
  IV U8811 ( .A(n8426), .Z(n8429) );
  XNOR U8812 ( .A(n4906), .B(n8426), .Z(n8428) );
  NAND U8813 ( .A(n8431), .B(e_input[645]), .Z(n4906) );
  NAND U8814 ( .A(n6112), .B(e_input[645]), .Z(n8431) );
  XOR U8815 ( .A(n8432), .B(n8433), .Z(n8426) );
  ANDN U8816 ( .A(n8434), .B(n4907), .Z(n8433) );
  XOR U8817 ( .A(n8435), .B(n8436), .Z(n4907) );
  IV U8818 ( .A(n8432), .Z(n8435) );
  XNOR U8819 ( .A(n4908), .B(n8432), .Z(n8434) );
  NAND U8820 ( .A(n8437), .B(e_input[644]), .Z(n4908) );
  NAND U8821 ( .A(n6112), .B(e_input[644]), .Z(n8437) );
  XOR U8822 ( .A(n8438), .B(n8439), .Z(n8432) );
  ANDN U8823 ( .A(n8440), .B(n4909), .Z(n8439) );
  XOR U8824 ( .A(n8441), .B(n8442), .Z(n4909) );
  IV U8825 ( .A(n8438), .Z(n8441) );
  XNOR U8826 ( .A(n4910), .B(n8438), .Z(n8440) );
  NAND U8827 ( .A(n8443), .B(e_input[643]), .Z(n4910) );
  NAND U8828 ( .A(n6112), .B(e_input[643]), .Z(n8443) );
  XOR U8829 ( .A(n8444), .B(n8445), .Z(n8438) );
  ANDN U8830 ( .A(n8446), .B(n4911), .Z(n8445) );
  XOR U8831 ( .A(n8447), .B(n8448), .Z(n4911) );
  IV U8832 ( .A(n8444), .Z(n8447) );
  XNOR U8833 ( .A(n4912), .B(n8444), .Z(n8446) );
  NAND U8834 ( .A(n8449), .B(e_input[642]), .Z(n4912) );
  NAND U8835 ( .A(n6112), .B(e_input[642]), .Z(n8449) );
  XOR U8836 ( .A(n8450), .B(n8451), .Z(n8444) );
  ANDN U8837 ( .A(n8452), .B(n4913), .Z(n8451) );
  XOR U8838 ( .A(n8453), .B(n8454), .Z(n4913) );
  IV U8839 ( .A(n8450), .Z(n8453) );
  XNOR U8840 ( .A(n4914), .B(n8450), .Z(n8452) );
  NAND U8841 ( .A(n8455), .B(e_input[641]), .Z(n4914) );
  NAND U8842 ( .A(n6112), .B(e_input[641]), .Z(n8455) );
  XOR U8843 ( .A(n8456), .B(n8457), .Z(n8450) );
  ANDN U8844 ( .A(n8458), .B(n4915), .Z(n8457) );
  XOR U8845 ( .A(n8459), .B(n8460), .Z(n4915) );
  IV U8846 ( .A(n8456), .Z(n8459) );
  XNOR U8847 ( .A(n4916), .B(n8456), .Z(n8458) );
  NAND U8848 ( .A(n8461), .B(e_input[640]), .Z(n4916) );
  NAND U8849 ( .A(n6112), .B(e_input[640]), .Z(n8461) );
  XOR U8850 ( .A(n8462), .B(n8463), .Z(n8456) );
  ANDN U8851 ( .A(n8464), .B(n4919), .Z(n8463) );
  XOR U8852 ( .A(n8465), .B(n8466), .Z(n4919) );
  IV U8853 ( .A(n8462), .Z(n8465) );
  XNOR U8854 ( .A(n4920), .B(n8462), .Z(n8464) );
  NAND U8855 ( .A(n8467), .B(e_input[639]), .Z(n4920) );
  NAND U8856 ( .A(n6112), .B(e_input[639]), .Z(n8467) );
  XOR U8857 ( .A(n8468), .B(n8469), .Z(n8462) );
  ANDN U8858 ( .A(n8470), .B(n4921), .Z(n8469) );
  XOR U8859 ( .A(n8471), .B(n8472), .Z(n4921) );
  IV U8860 ( .A(n8468), .Z(n8471) );
  XNOR U8861 ( .A(n4922), .B(n8468), .Z(n8470) );
  NAND U8862 ( .A(n8473), .B(e_input[638]), .Z(n4922) );
  NAND U8863 ( .A(n6112), .B(e_input[638]), .Z(n8473) );
  XOR U8864 ( .A(n8474), .B(n8475), .Z(n8468) );
  ANDN U8865 ( .A(n8476), .B(n4923), .Z(n8475) );
  XOR U8866 ( .A(n8477), .B(n8478), .Z(n4923) );
  IV U8867 ( .A(n8474), .Z(n8477) );
  XNOR U8868 ( .A(n4924), .B(n8474), .Z(n8476) );
  NAND U8869 ( .A(n8479), .B(e_input[637]), .Z(n4924) );
  NAND U8870 ( .A(n6112), .B(e_input[637]), .Z(n8479) );
  XOR U8871 ( .A(n8480), .B(n8481), .Z(n8474) );
  ANDN U8872 ( .A(n8482), .B(n4925), .Z(n8481) );
  XOR U8873 ( .A(n8483), .B(n8484), .Z(n4925) );
  IV U8874 ( .A(n8480), .Z(n8483) );
  XNOR U8875 ( .A(n4926), .B(n8480), .Z(n8482) );
  NAND U8876 ( .A(n8485), .B(e_input[636]), .Z(n4926) );
  NAND U8877 ( .A(n6112), .B(e_input[636]), .Z(n8485) );
  XOR U8878 ( .A(n8486), .B(n8487), .Z(n8480) );
  ANDN U8879 ( .A(n8488), .B(n4927), .Z(n8487) );
  XOR U8880 ( .A(n8489), .B(n8490), .Z(n4927) );
  IV U8881 ( .A(n8486), .Z(n8489) );
  XNOR U8882 ( .A(n4928), .B(n8486), .Z(n8488) );
  NAND U8883 ( .A(n8491), .B(e_input[635]), .Z(n4928) );
  NAND U8884 ( .A(n6112), .B(e_input[635]), .Z(n8491) );
  XOR U8885 ( .A(n8492), .B(n8493), .Z(n8486) );
  ANDN U8886 ( .A(n8494), .B(n4929), .Z(n8493) );
  XOR U8887 ( .A(n8495), .B(n8496), .Z(n4929) );
  IV U8888 ( .A(n8492), .Z(n8495) );
  XNOR U8889 ( .A(n4930), .B(n8492), .Z(n8494) );
  NAND U8890 ( .A(n8497), .B(e_input[634]), .Z(n4930) );
  NAND U8891 ( .A(n6112), .B(e_input[634]), .Z(n8497) );
  XOR U8892 ( .A(n8498), .B(n8499), .Z(n8492) );
  ANDN U8893 ( .A(n8500), .B(n4931), .Z(n8499) );
  XOR U8894 ( .A(n8501), .B(n8502), .Z(n4931) );
  IV U8895 ( .A(n8498), .Z(n8501) );
  XNOR U8896 ( .A(n4932), .B(n8498), .Z(n8500) );
  NAND U8897 ( .A(n8503), .B(e_input[633]), .Z(n4932) );
  NAND U8898 ( .A(n6112), .B(e_input[633]), .Z(n8503) );
  XOR U8899 ( .A(n8504), .B(n8505), .Z(n8498) );
  ANDN U8900 ( .A(n8506), .B(n4933), .Z(n8505) );
  XOR U8901 ( .A(n8507), .B(n8508), .Z(n4933) );
  IV U8902 ( .A(n8504), .Z(n8507) );
  XNOR U8903 ( .A(n4934), .B(n8504), .Z(n8506) );
  NAND U8904 ( .A(n8509), .B(e_input[632]), .Z(n4934) );
  NAND U8905 ( .A(n6112), .B(e_input[632]), .Z(n8509) );
  XOR U8906 ( .A(n8510), .B(n8511), .Z(n8504) );
  ANDN U8907 ( .A(n8512), .B(n4935), .Z(n8511) );
  XOR U8908 ( .A(n8513), .B(n8514), .Z(n4935) );
  IV U8909 ( .A(n8510), .Z(n8513) );
  XNOR U8910 ( .A(n4936), .B(n8510), .Z(n8512) );
  NAND U8911 ( .A(n8515), .B(e_input[631]), .Z(n4936) );
  NAND U8912 ( .A(n6112), .B(e_input[631]), .Z(n8515) );
  XOR U8913 ( .A(n8516), .B(n8517), .Z(n8510) );
  ANDN U8914 ( .A(n8518), .B(n4937), .Z(n8517) );
  XOR U8915 ( .A(n8519), .B(n8520), .Z(n4937) );
  IV U8916 ( .A(n8516), .Z(n8519) );
  XNOR U8917 ( .A(n4938), .B(n8516), .Z(n8518) );
  NAND U8918 ( .A(n8521), .B(e_input[630]), .Z(n4938) );
  NAND U8919 ( .A(n6112), .B(e_input[630]), .Z(n8521) );
  XOR U8920 ( .A(n8522), .B(n8523), .Z(n8516) );
  ANDN U8921 ( .A(n8524), .B(n4941), .Z(n8523) );
  XOR U8922 ( .A(n8525), .B(n8526), .Z(n4941) );
  IV U8923 ( .A(n8522), .Z(n8525) );
  XNOR U8924 ( .A(n4942), .B(n8522), .Z(n8524) );
  NAND U8925 ( .A(n8527), .B(e_input[629]), .Z(n4942) );
  NAND U8926 ( .A(n6112), .B(e_input[629]), .Z(n8527) );
  XOR U8927 ( .A(n8528), .B(n8529), .Z(n8522) );
  ANDN U8928 ( .A(n8530), .B(n4943), .Z(n8529) );
  XOR U8929 ( .A(n8531), .B(n8532), .Z(n4943) );
  IV U8930 ( .A(n8528), .Z(n8531) );
  XNOR U8931 ( .A(n4944), .B(n8528), .Z(n8530) );
  NAND U8932 ( .A(n8533), .B(e_input[628]), .Z(n4944) );
  NAND U8933 ( .A(n6112), .B(e_input[628]), .Z(n8533) );
  XOR U8934 ( .A(n8534), .B(n8535), .Z(n8528) );
  ANDN U8935 ( .A(n8536), .B(n4945), .Z(n8535) );
  XOR U8936 ( .A(n8537), .B(n8538), .Z(n4945) );
  IV U8937 ( .A(n8534), .Z(n8537) );
  XNOR U8938 ( .A(n4946), .B(n8534), .Z(n8536) );
  NAND U8939 ( .A(n8539), .B(e_input[627]), .Z(n4946) );
  NAND U8940 ( .A(n6112), .B(e_input[627]), .Z(n8539) );
  XOR U8941 ( .A(n8540), .B(n8541), .Z(n8534) );
  ANDN U8942 ( .A(n8542), .B(n4947), .Z(n8541) );
  XOR U8943 ( .A(n8543), .B(n8544), .Z(n4947) );
  IV U8944 ( .A(n8540), .Z(n8543) );
  XNOR U8945 ( .A(n4948), .B(n8540), .Z(n8542) );
  NAND U8946 ( .A(n8545), .B(e_input[626]), .Z(n4948) );
  NAND U8947 ( .A(n6112), .B(e_input[626]), .Z(n8545) );
  XOR U8948 ( .A(n8546), .B(n8547), .Z(n8540) );
  ANDN U8949 ( .A(n8548), .B(n4949), .Z(n8547) );
  XOR U8950 ( .A(n8549), .B(n8550), .Z(n4949) );
  IV U8951 ( .A(n8546), .Z(n8549) );
  XNOR U8952 ( .A(n4950), .B(n8546), .Z(n8548) );
  NAND U8953 ( .A(n8551), .B(e_input[625]), .Z(n4950) );
  NAND U8954 ( .A(n6112), .B(e_input[625]), .Z(n8551) );
  XOR U8955 ( .A(n8552), .B(n8553), .Z(n8546) );
  ANDN U8956 ( .A(n8554), .B(n4951), .Z(n8553) );
  XOR U8957 ( .A(n8555), .B(n8556), .Z(n4951) );
  IV U8958 ( .A(n8552), .Z(n8555) );
  XNOR U8959 ( .A(n4952), .B(n8552), .Z(n8554) );
  NAND U8960 ( .A(n8557), .B(e_input[624]), .Z(n4952) );
  NAND U8961 ( .A(n6112), .B(e_input[624]), .Z(n8557) );
  XOR U8962 ( .A(n8558), .B(n8559), .Z(n8552) );
  ANDN U8963 ( .A(n8560), .B(n4953), .Z(n8559) );
  XOR U8964 ( .A(n8561), .B(n8562), .Z(n4953) );
  IV U8965 ( .A(n8558), .Z(n8561) );
  XNOR U8966 ( .A(n4954), .B(n8558), .Z(n8560) );
  NAND U8967 ( .A(n8563), .B(e_input[623]), .Z(n4954) );
  NAND U8968 ( .A(n6112), .B(e_input[623]), .Z(n8563) );
  XOR U8969 ( .A(n8564), .B(n8565), .Z(n8558) );
  ANDN U8970 ( .A(n8566), .B(n4955), .Z(n8565) );
  XOR U8971 ( .A(n8567), .B(n8568), .Z(n4955) );
  IV U8972 ( .A(n8564), .Z(n8567) );
  XNOR U8973 ( .A(n4956), .B(n8564), .Z(n8566) );
  NAND U8974 ( .A(n8569), .B(e_input[622]), .Z(n4956) );
  NAND U8975 ( .A(n6112), .B(e_input[622]), .Z(n8569) );
  XOR U8976 ( .A(n8570), .B(n8571), .Z(n8564) );
  ANDN U8977 ( .A(n8572), .B(n4957), .Z(n8571) );
  XOR U8978 ( .A(n8573), .B(n8574), .Z(n4957) );
  IV U8979 ( .A(n8570), .Z(n8573) );
  XNOR U8980 ( .A(n4958), .B(n8570), .Z(n8572) );
  NAND U8981 ( .A(n8575), .B(e_input[621]), .Z(n4958) );
  NAND U8982 ( .A(n6112), .B(e_input[621]), .Z(n8575) );
  XOR U8983 ( .A(n8576), .B(n8577), .Z(n8570) );
  ANDN U8984 ( .A(n8578), .B(n4959), .Z(n8577) );
  XOR U8985 ( .A(n8579), .B(n8580), .Z(n4959) );
  IV U8986 ( .A(n8576), .Z(n8579) );
  XNOR U8987 ( .A(n4960), .B(n8576), .Z(n8578) );
  NAND U8988 ( .A(n8581), .B(e_input[620]), .Z(n4960) );
  NAND U8989 ( .A(n6112), .B(e_input[620]), .Z(n8581) );
  XOR U8990 ( .A(n8582), .B(n8583), .Z(n8576) );
  ANDN U8991 ( .A(n8584), .B(n4963), .Z(n8583) );
  XOR U8992 ( .A(n8585), .B(n8586), .Z(n4963) );
  IV U8993 ( .A(n8582), .Z(n8585) );
  XNOR U8994 ( .A(n4964), .B(n8582), .Z(n8584) );
  NAND U8995 ( .A(n8587), .B(e_input[619]), .Z(n4964) );
  NAND U8996 ( .A(n6112), .B(e_input[619]), .Z(n8587) );
  XOR U8997 ( .A(n8588), .B(n8589), .Z(n8582) );
  ANDN U8998 ( .A(n8590), .B(n4965), .Z(n8589) );
  XOR U8999 ( .A(n8591), .B(n8592), .Z(n4965) );
  IV U9000 ( .A(n8588), .Z(n8591) );
  XNOR U9001 ( .A(n4966), .B(n8588), .Z(n8590) );
  NAND U9002 ( .A(n8593), .B(e_input[618]), .Z(n4966) );
  NAND U9003 ( .A(n6112), .B(e_input[618]), .Z(n8593) );
  XOR U9004 ( .A(n8594), .B(n8595), .Z(n8588) );
  ANDN U9005 ( .A(n8596), .B(n4967), .Z(n8595) );
  XOR U9006 ( .A(n8597), .B(n8598), .Z(n4967) );
  IV U9007 ( .A(n8594), .Z(n8597) );
  XNOR U9008 ( .A(n4968), .B(n8594), .Z(n8596) );
  NAND U9009 ( .A(n8599), .B(e_input[617]), .Z(n4968) );
  NAND U9010 ( .A(n6112), .B(e_input[617]), .Z(n8599) );
  XOR U9011 ( .A(n8600), .B(n8601), .Z(n8594) );
  ANDN U9012 ( .A(n8602), .B(n4969), .Z(n8601) );
  XOR U9013 ( .A(n8603), .B(n8604), .Z(n4969) );
  IV U9014 ( .A(n8600), .Z(n8603) );
  XNOR U9015 ( .A(n4970), .B(n8600), .Z(n8602) );
  NAND U9016 ( .A(n8605), .B(e_input[616]), .Z(n4970) );
  NAND U9017 ( .A(n6112), .B(e_input[616]), .Z(n8605) );
  XOR U9018 ( .A(n8606), .B(n8607), .Z(n8600) );
  ANDN U9019 ( .A(n8608), .B(n4971), .Z(n8607) );
  XOR U9020 ( .A(n8609), .B(n8610), .Z(n4971) );
  IV U9021 ( .A(n8606), .Z(n8609) );
  XNOR U9022 ( .A(n4972), .B(n8606), .Z(n8608) );
  NAND U9023 ( .A(n8611), .B(e_input[615]), .Z(n4972) );
  NAND U9024 ( .A(n6112), .B(e_input[615]), .Z(n8611) );
  XOR U9025 ( .A(n8612), .B(n8613), .Z(n8606) );
  ANDN U9026 ( .A(n8614), .B(n4973), .Z(n8613) );
  XOR U9027 ( .A(n8615), .B(n8616), .Z(n4973) );
  IV U9028 ( .A(n8612), .Z(n8615) );
  XNOR U9029 ( .A(n4974), .B(n8612), .Z(n8614) );
  NAND U9030 ( .A(n8617), .B(e_input[614]), .Z(n4974) );
  NAND U9031 ( .A(n6112), .B(e_input[614]), .Z(n8617) );
  XOR U9032 ( .A(n8618), .B(n8619), .Z(n8612) );
  ANDN U9033 ( .A(n8620), .B(n4975), .Z(n8619) );
  XOR U9034 ( .A(n8621), .B(n8622), .Z(n4975) );
  IV U9035 ( .A(n8618), .Z(n8621) );
  XNOR U9036 ( .A(n4976), .B(n8618), .Z(n8620) );
  NAND U9037 ( .A(n8623), .B(e_input[613]), .Z(n4976) );
  NAND U9038 ( .A(n6112), .B(e_input[613]), .Z(n8623) );
  XOR U9039 ( .A(n8624), .B(n8625), .Z(n8618) );
  ANDN U9040 ( .A(n8626), .B(n4977), .Z(n8625) );
  XOR U9041 ( .A(n8627), .B(n8628), .Z(n4977) );
  IV U9042 ( .A(n8624), .Z(n8627) );
  XNOR U9043 ( .A(n4978), .B(n8624), .Z(n8626) );
  NAND U9044 ( .A(n8629), .B(e_input[612]), .Z(n4978) );
  NAND U9045 ( .A(n6112), .B(e_input[612]), .Z(n8629) );
  XOR U9046 ( .A(n8630), .B(n8631), .Z(n8624) );
  ANDN U9047 ( .A(n8632), .B(n4979), .Z(n8631) );
  XOR U9048 ( .A(n8633), .B(n8634), .Z(n4979) );
  IV U9049 ( .A(n8630), .Z(n8633) );
  XNOR U9050 ( .A(n4980), .B(n8630), .Z(n8632) );
  NAND U9051 ( .A(n8635), .B(e_input[611]), .Z(n4980) );
  NAND U9052 ( .A(n6112), .B(e_input[611]), .Z(n8635) );
  XOR U9053 ( .A(n8636), .B(n8637), .Z(n8630) );
  ANDN U9054 ( .A(n8638), .B(n4981), .Z(n8637) );
  XOR U9055 ( .A(n8639), .B(n8640), .Z(n4981) );
  IV U9056 ( .A(n8636), .Z(n8639) );
  XNOR U9057 ( .A(n4982), .B(n8636), .Z(n8638) );
  NAND U9058 ( .A(n8641), .B(e_input[610]), .Z(n4982) );
  NAND U9059 ( .A(n6112), .B(e_input[610]), .Z(n8641) );
  XOR U9060 ( .A(n8642), .B(n8643), .Z(n8636) );
  ANDN U9061 ( .A(n8644), .B(n4985), .Z(n8643) );
  XOR U9062 ( .A(n8645), .B(n8646), .Z(n4985) );
  IV U9063 ( .A(n8642), .Z(n8645) );
  XNOR U9064 ( .A(n4986), .B(n8642), .Z(n8644) );
  NAND U9065 ( .A(n8647), .B(e_input[609]), .Z(n4986) );
  NAND U9066 ( .A(n6112), .B(e_input[609]), .Z(n8647) );
  XOR U9067 ( .A(n8648), .B(n8649), .Z(n8642) );
  ANDN U9068 ( .A(n8650), .B(n4987), .Z(n8649) );
  XOR U9069 ( .A(n8651), .B(n8652), .Z(n4987) );
  IV U9070 ( .A(n8648), .Z(n8651) );
  XNOR U9071 ( .A(n4988), .B(n8648), .Z(n8650) );
  NAND U9072 ( .A(n8653), .B(e_input[608]), .Z(n4988) );
  NAND U9073 ( .A(n6112), .B(e_input[608]), .Z(n8653) );
  XOR U9074 ( .A(n8654), .B(n8655), .Z(n8648) );
  ANDN U9075 ( .A(n8656), .B(n4989), .Z(n8655) );
  XOR U9076 ( .A(n8657), .B(n8658), .Z(n4989) );
  IV U9077 ( .A(n8654), .Z(n8657) );
  XNOR U9078 ( .A(n4990), .B(n8654), .Z(n8656) );
  NAND U9079 ( .A(n8659), .B(e_input[607]), .Z(n4990) );
  NAND U9080 ( .A(n6112), .B(e_input[607]), .Z(n8659) );
  XOR U9081 ( .A(n8660), .B(n8661), .Z(n8654) );
  ANDN U9082 ( .A(n8662), .B(n4991), .Z(n8661) );
  XOR U9083 ( .A(n8663), .B(n8664), .Z(n4991) );
  IV U9084 ( .A(n8660), .Z(n8663) );
  XNOR U9085 ( .A(n4992), .B(n8660), .Z(n8662) );
  NAND U9086 ( .A(n8665), .B(e_input[606]), .Z(n4992) );
  NAND U9087 ( .A(n6112), .B(e_input[606]), .Z(n8665) );
  XOR U9088 ( .A(n8666), .B(n8667), .Z(n8660) );
  ANDN U9089 ( .A(n8668), .B(n4993), .Z(n8667) );
  XOR U9090 ( .A(n8669), .B(n8670), .Z(n4993) );
  IV U9091 ( .A(n8666), .Z(n8669) );
  XNOR U9092 ( .A(n4994), .B(n8666), .Z(n8668) );
  NAND U9093 ( .A(n8671), .B(e_input[605]), .Z(n4994) );
  NAND U9094 ( .A(n6112), .B(e_input[605]), .Z(n8671) );
  XOR U9095 ( .A(n8672), .B(n8673), .Z(n8666) );
  ANDN U9096 ( .A(n8674), .B(n4995), .Z(n8673) );
  XOR U9097 ( .A(n8675), .B(n8676), .Z(n4995) );
  IV U9098 ( .A(n8672), .Z(n8675) );
  XNOR U9099 ( .A(n4996), .B(n8672), .Z(n8674) );
  NAND U9100 ( .A(n8677), .B(e_input[604]), .Z(n4996) );
  NAND U9101 ( .A(n6112), .B(e_input[604]), .Z(n8677) );
  XOR U9102 ( .A(n8678), .B(n8679), .Z(n8672) );
  ANDN U9103 ( .A(n8680), .B(n4997), .Z(n8679) );
  XOR U9104 ( .A(n8681), .B(n8682), .Z(n4997) );
  IV U9105 ( .A(n8678), .Z(n8681) );
  XNOR U9106 ( .A(n4998), .B(n8678), .Z(n8680) );
  NAND U9107 ( .A(n8683), .B(e_input[603]), .Z(n4998) );
  NAND U9108 ( .A(n6112), .B(e_input[603]), .Z(n8683) );
  XOR U9109 ( .A(n8684), .B(n8685), .Z(n8678) );
  ANDN U9110 ( .A(n8686), .B(n4999), .Z(n8685) );
  XOR U9111 ( .A(n8687), .B(n8688), .Z(n4999) );
  IV U9112 ( .A(n8684), .Z(n8687) );
  XNOR U9113 ( .A(n5000), .B(n8684), .Z(n8686) );
  NAND U9114 ( .A(n8689), .B(e_input[602]), .Z(n5000) );
  NAND U9115 ( .A(n6112), .B(e_input[602]), .Z(n8689) );
  XOR U9116 ( .A(n8690), .B(n8691), .Z(n8684) );
  ANDN U9117 ( .A(n8692), .B(n5001), .Z(n8691) );
  XOR U9118 ( .A(n8693), .B(n8694), .Z(n5001) );
  IV U9119 ( .A(n8690), .Z(n8693) );
  XNOR U9120 ( .A(n5002), .B(n8690), .Z(n8692) );
  NAND U9121 ( .A(n8695), .B(e_input[601]), .Z(n5002) );
  NAND U9122 ( .A(n6112), .B(e_input[601]), .Z(n8695) );
  XOR U9123 ( .A(n8696), .B(n8697), .Z(n8690) );
  ANDN U9124 ( .A(n8698), .B(n5003), .Z(n8697) );
  XOR U9125 ( .A(n8699), .B(n8700), .Z(n5003) );
  IV U9126 ( .A(n8696), .Z(n8699) );
  XNOR U9127 ( .A(n5004), .B(n8696), .Z(n8698) );
  NAND U9128 ( .A(n8701), .B(e_input[600]), .Z(n5004) );
  NAND U9129 ( .A(n6112), .B(e_input[600]), .Z(n8701) );
  XOR U9130 ( .A(n8702), .B(n8703), .Z(n8696) );
  ANDN U9131 ( .A(n8704), .B(n5009), .Z(n8703) );
  XOR U9132 ( .A(n8705), .B(n8706), .Z(n5009) );
  IV U9133 ( .A(n8702), .Z(n8705) );
  XNOR U9134 ( .A(n5010), .B(n8702), .Z(n8704) );
  NAND U9135 ( .A(n8707), .B(e_input[599]), .Z(n5010) );
  NAND U9136 ( .A(n6112), .B(e_input[599]), .Z(n8707) );
  XOR U9137 ( .A(n8708), .B(n8709), .Z(n8702) );
  ANDN U9138 ( .A(n8710), .B(n5011), .Z(n8709) );
  XOR U9139 ( .A(n8711), .B(n8712), .Z(n5011) );
  IV U9140 ( .A(n8708), .Z(n8711) );
  XNOR U9141 ( .A(n5012), .B(n8708), .Z(n8710) );
  NAND U9142 ( .A(n8713), .B(e_input[598]), .Z(n5012) );
  NAND U9143 ( .A(n6112), .B(e_input[598]), .Z(n8713) );
  XOR U9144 ( .A(n8714), .B(n8715), .Z(n8708) );
  ANDN U9145 ( .A(n8716), .B(n5013), .Z(n8715) );
  XOR U9146 ( .A(n8717), .B(n8718), .Z(n5013) );
  IV U9147 ( .A(n8714), .Z(n8717) );
  XNOR U9148 ( .A(n5014), .B(n8714), .Z(n8716) );
  NAND U9149 ( .A(n8719), .B(e_input[597]), .Z(n5014) );
  NAND U9150 ( .A(n6112), .B(e_input[597]), .Z(n8719) );
  XOR U9151 ( .A(n8720), .B(n8721), .Z(n8714) );
  ANDN U9152 ( .A(n8722), .B(n5015), .Z(n8721) );
  XOR U9153 ( .A(n8723), .B(n8724), .Z(n5015) );
  IV U9154 ( .A(n8720), .Z(n8723) );
  XNOR U9155 ( .A(n5016), .B(n8720), .Z(n8722) );
  NAND U9156 ( .A(n8725), .B(e_input[596]), .Z(n5016) );
  NAND U9157 ( .A(n6112), .B(e_input[596]), .Z(n8725) );
  XOR U9158 ( .A(n8726), .B(n8727), .Z(n8720) );
  ANDN U9159 ( .A(n8728), .B(n5017), .Z(n8727) );
  XOR U9160 ( .A(n8729), .B(n8730), .Z(n5017) );
  IV U9161 ( .A(n8726), .Z(n8729) );
  XNOR U9162 ( .A(n5018), .B(n8726), .Z(n8728) );
  NAND U9163 ( .A(n8731), .B(e_input[595]), .Z(n5018) );
  NAND U9164 ( .A(n6112), .B(e_input[595]), .Z(n8731) );
  XOR U9165 ( .A(n8732), .B(n8733), .Z(n8726) );
  ANDN U9166 ( .A(n8734), .B(n5019), .Z(n8733) );
  XOR U9167 ( .A(n8735), .B(n8736), .Z(n5019) );
  IV U9168 ( .A(n8732), .Z(n8735) );
  XNOR U9169 ( .A(n5020), .B(n8732), .Z(n8734) );
  NAND U9170 ( .A(n8737), .B(e_input[594]), .Z(n5020) );
  NAND U9171 ( .A(n6112), .B(e_input[594]), .Z(n8737) );
  XOR U9172 ( .A(n8738), .B(n8739), .Z(n8732) );
  ANDN U9173 ( .A(n8740), .B(n5021), .Z(n8739) );
  XOR U9174 ( .A(n8741), .B(n8742), .Z(n5021) );
  IV U9175 ( .A(n8738), .Z(n8741) );
  XNOR U9176 ( .A(n5022), .B(n8738), .Z(n8740) );
  NAND U9177 ( .A(n8743), .B(e_input[593]), .Z(n5022) );
  NAND U9178 ( .A(n6112), .B(e_input[593]), .Z(n8743) );
  XOR U9179 ( .A(n8744), .B(n8745), .Z(n8738) );
  ANDN U9180 ( .A(n8746), .B(n5023), .Z(n8745) );
  XOR U9181 ( .A(n8747), .B(n8748), .Z(n5023) );
  IV U9182 ( .A(n8744), .Z(n8747) );
  XNOR U9183 ( .A(n5024), .B(n8744), .Z(n8746) );
  NAND U9184 ( .A(n8749), .B(e_input[592]), .Z(n5024) );
  NAND U9185 ( .A(n6112), .B(e_input[592]), .Z(n8749) );
  XOR U9186 ( .A(n8750), .B(n8751), .Z(n8744) );
  ANDN U9187 ( .A(n8752), .B(n5025), .Z(n8751) );
  XOR U9188 ( .A(n8753), .B(n8754), .Z(n5025) );
  IV U9189 ( .A(n8750), .Z(n8753) );
  XNOR U9190 ( .A(n5026), .B(n8750), .Z(n8752) );
  NAND U9191 ( .A(n8755), .B(e_input[591]), .Z(n5026) );
  NAND U9192 ( .A(n6112), .B(e_input[591]), .Z(n8755) );
  XOR U9193 ( .A(n8756), .B(n8757), .Z(n8750) );
  ANDN U9194 ( .A(n8758), .B(n5027), .Z(n8757) );
  XOR U9195 ( .A(n8759), .B(n8760), .Z(n5027) );
  IV U9196 ( .A(n8756), .Z(n8759) );
  XNOR U9197 ( .A(n5028), .B(n8756), .Z(n8758) );
  NAND U9198 ( .A(n8761), .B(e_input[590]), .Z(n5028) );
  NAND U9199 ( .A(n6112), .B(e_input[590]), .Z(n8761) );
  XOR U9200 ( .A(n8762), .B(n8763), .Z(n8756) );
  ANDN U9201 ( .A(n8764), .B(n5031), .Z(n8763) );
  XOR U9202 ( .A(n8765), .B(n8766), .Z(n5031) );
  IV U9203 ( .A(n8762), .Z(n8765) );
  XNOR U9204 ( .A(n5032), .B(n8762), .Z(n8764) );
  NAND U9205 ( .A(n8767), .B(e_input[589]), .Z(n5032) );
  NAND U9206 ( .A(n6112), .B(e_input[589]), .Z(n8767) );
  XOR U9207 ( .A(n8768), .B(n8769), .Z(n8762) );
  ANDN U9208 ( .A(n8770), .B(n5033), .Z(n8769) );
  XOR U9209 ( .A(n8771), .B(n8772), .Z(n5033) );
  IV U9210 ( .A(n8768), .Z(n8771) );
  XNOR U9211 ( .A(n5034), .B(n8768), .Z(n8770) );
  NAND U9212 ( .A(n8773), .B(e_input[588]), .Z(n5034) );
  NAND U9213 ( .A(n6112), .B(e_input[588]), .Z(n8773) );
  XOR U9214 ( .A(n8774), .B(n8775), .Z(n8768) );
  ANDN U9215 ( .A(n8776), .B(n5035), .Z(n8775) );
  XOR U9216 ( .A(n8777), .B(n8778), .Z(n5035) );
  IV U9217 ( .A(n8774), .Z(n8777) );
  XNOR U9218 ( .A(n5036), .B(n8774), .Z(n8776) );
  NAND U9219 ( .A(n8779), .B(e_input[587]), .Z(n5036) );
  NAND U9220 ( .A(n6112), .B(e_input[587]), .Z(n8779) );
  XOR U9221 ( .A(n8780), .B(n8781), .Z(n8774) );
  ANDN U9222 ( .A(n8782), .B(n5037), .Z(n8781) );
  XOR U9223 ( .A(n8783), .B(n8784), .Z(n5037) );
  IV U9224 ( .A(n8780), .Z(n8783) );
  XNOR U9225 ( .A(n5038), .B(n8780), .Z(n8782) );
  NAND U9226 ( .A(n8785), .B(e_input[586]), .Z(n5038) );
  NAND U9227 ( .A(n6112), .B(e_input[586]), .Z(n8785) );
  XOR U9228 ( .A(n8786), .B(n8787), .Z(n8780) );
  ANDN U9229 ( .A(n8788), .B(n5039), .Z(n8787) );
  XOR U9230 ( .A(n8789), .B(n8790), .Z(n5039) );
  IV U9231 ( .A(n8786), .Z(n8789) );
  XNOR U9232 ( .A(n5040), .B(n8786), .Z(n8788) );
  NAND U9233 ( .A(n8791), .B(e_input[585]), .Z(n5040) );
  NAND U9234 ( .A(n6112), .B(e_input[585]), .Z(n8791) );
  XOR U9235 ( .A(n8792), .B(n8793), .Z(n8786) );
  ANDN U9236 ( .A(n8794), .B(n5041), .Z(n8793) );
  XOR U9237 ( .A(n8795), .B(n8796), .Z(n5041) );
  IV U9238 ( .A(n8792), .Z(n8795) );
  XNOR U9239 ( .A(n5042), .B(n8792), .Z(n8794) );
  NAND U9240 ( .A(n8797), .B(e_input[584]), .Z(n5042) );
  NAND U9241 ( .A(n6112), .B(e_input[584]), .Z(n8797) );
  XOR U9242 ( .A(n8798), .B(n8799), .Z(n8792) );
  ANDN U9243 ( .A(n8800), .B(n5043), .Z(n8799) );
  XOR U9244 ( .A(n8801), .B(n8802), .Z(n5043) );
  IV U9245 ( .A(n8798), .Z(n8801) );
  XNOR U9246 ( .A(n5044), .B(n8798), .Z(n8800) );
  NAND U9247 ( .A(n8803), .B(e_input[583]), .Z(n5044) );
  NAND U9248 ( .A(n6112), .B(e_input[583]), .Z(n8803) );
  XOR U9249 ( .A(n8804), .B(n8805), .Z(n8798) );
  ANDN U9250 ( .A(n8806), .B(n5045), .Z(n8805) );
  XOR U9251 ( .A(n8807), .B(n8808), .Z(n5045) );
  IV U9252 ( .A(n8804), .Z(n8807) );
  XNOR U9253 ( .A(n5046), .B(n8804), .Z(n8806) );
  NAND U9254 ( .A(n8809), .B(e_input[582]), .Z(n5046) );
  NAND U9255 ( .A(n6112), .B(e_input[582]), .Z(n8809) );
  XOR U9256 ( .A(n8810), .B(n8811), .Z(n8804) );
  ANDN U9257 ( .A(n8812), .B(n5047), .Z(n8811) );
  XOR U9258 ( .A(n8813), .B(n8814), .Z(n5047) );
  IV U9259 ( .A(n8810), .Z(n8813) );
  XNOR U9260 ( .A(n5048), .B(n8810), .Z(n8812) );
  NAND U9261 ( .A(n8815), .B(e_input[581]), .Z(n5048) );
  NAND U9262 ( .A(n6112), .B(e_input[581]), .Z(n8815) );
  XOR U9263 ( .A(n8816), .B(n8817), .Z(n8810) );
  ANDN U9264 ( .A(n8818), .B(n5049), .Z(n8817) );
  XOR U9265 ( .A(n8819), .B(n8820), .Z(n5049) );
  IV U9266 ( .A(n8816), .Z(n8819) );
  XNOR U9267 ( .A(n5050), .B(n8816), .Z(n8818) );
  NAND U9268 ( .A(n8821), .B(e_input[580]), .Z(n5050) );
  NAND U9269 ( .A(n6112), .B(e_input[580]), .Z(n8821) );
  XOR U9270 ( .A(n8822), .B(n8823), .Z(n8816) );
  ANDN U9271 ( .A(n8824), .B(n5053), .Z(n8823) );
  XOR U9272 ( .A(n8825), .B(n8826), .Z(n5053) );
  IV U9273 ( .A(n8822), .Z(n8825) );
  XNOR U9274 ( .A(n5054), .B(n8822), .Z(n8824) );
  NAND U9275 ( .A(n8827), .B(e_input[579]), .Z(n5054) );
  NAND U9276 ( .A(n6112), .B(e_input[579]), .Z(n8827) );
  XOR U9277 ( .A(n8828), .B(n8829), .Z(n8822) );
  ANDN U9278 ( .A(n8830), .B(n5055), .Z(n8829) );
  XOR U9279 ( .A(n8831), .B(n8832), .Z(n5055) );
  IV U9280 ( .A(n8828), .Z(n8831) );
  XNOR U9281 ( .A(n5056), .B(n8828), .Z(n8830) );
  NAND U9282 ( .A(n8833), .B(e_input[578]), .Z(n5056) );
  NAND U9283 ( .A(n6112), .B(e_input[578]), .Z(n8833) );
  XOR U9284 ( .A(n8834), .B(n8835), .Z(n8828) );
  ANDN U9285 ( .A(n8836), .B(n5057), .Z(n8835) );
  XOR U9286 ( .A(n8837), .B(n8838), .Z(n5057) );
  IV U9287 ( .A(n8834), .Z(n8837) );
  XNOR U9288 ( .A(n5058), .B(n8834), .Z(n8836) );
  NAND U9289 ( .A(n8839), .B(e_input[577]), .Z(n5058) );
  NAND U9290 ( .A(n6112), .B(e_input[577]), .Z(n8839) );
  XOR U9291 ( .A(n8840), .B(n8841), .Z(n8834) );
  ANDN U9292 ( .A(n8842), .B(n5059), .Z(n8841) );
  XOR U9293 ( .A(n8843), .B(n8844), .Z(n5059) );
  IV U9294 ( .A(n8840), .Z(n8843) );
  XNOR U9295 ( .A(n5060), .B(n8840), .Z(n8842) );
  NAND U9296 ( .A(n8845), .B(e_input[576]), .Z(n5060) );
  NAND U9297 ( .A(n6112), .B(e_input[576]), .Z(n8845) );
  XOR U9298 ( .A(n8846), .B(n8847), .Z(n8840) );
  ANDN U9299 ( .A(n8848), .B(n5061), .Z(n8847) );
  XOR U9300 ( .A(n8849), .B(n8850), .Z(n5061) );
  IV U9301 ( .A(n8846), .Z(n8849) );
  XNOR U9302 ( .A(n5062), .B(n8846), .Z(n8848) );
  NAND U9303 ( .A(n8851), .B(e_input[575]), .Z(n5062) );
  NAND U9304 ( .A(n6112), .B(e_input[575]), .Z(n8851) );
  XOR U9305 ( .A(n8852), .B(n8853), .Z(n8846) );
  ANDN U9306 ( .A(n8854), .B(n5063), .Z(n8853) );
  XOR U9307 ( .A(n8855), .B(n8856), .Z(n5063) );
  IV U9308 ( .A(n8852), .Z(n8855) );
  XNOR U9309 ( .A(n5064), .B(n8852), .Z(n8854) );
  NAND U9310 ( .A(n8857), .B(e_input[574]), .Z(n5064) );
  NAND U9311 ( .A(n6112), .B(e_input[574]), .Z(n8857) );
  XOR U9312 ( .A(n8858), .B(n8859), .Z(n8852) );
  ANDN U9313 ( .A(n8860), .B(n5065), .Z(n8859) );
  XOR U9314 ( .A(n8861), .B(n8862), .Z(n5065) );
  IV U9315 ( .A(n8858), .Z(n8861) );
  XNOR U9316 ( .A(n5066), .B(n8858), .Z(n8860) );
  NAND U9317 ( .A(n8863), .B(e_input[573]), .Z(n5066) );
  NAND U9318 ( .A(n6112), .B(e_input[573]), .Z(n8863) );
  XOR U9319 ( .A(n8864), .B(n8865), .Z(n8858) );
  ANDN U9320 ( .A(n8866), .B(n5067), .Z(n8865) );
  XOR U9321 ( .A(n8867), .B(n8868), .Z(n5067) );
  IV U9322 ( .A(n8864), .Z(n8867) );
  XNOR U9323 ( .A(n5068), .B(n8864), .Z(n8866) );
  NAND U9324 ( .A(n8869), .B(e_input[572]), .Z(n5068) );
  NAND U9325 ( .A(n6112), .B(e_input[572]), .Z(n8869) );
  XOR U9326 ( .A(n8870), .B(n8871), .Z(n8864) );
  ANDN U9327 ( .A(n8872), .B(n5069), .Z(n8871) );
  XOR U9328 ( .A(n8873), .B(n8874), .Z(n5069) );
  IV U9329 ( .A(n8870), .Z(n8873) );
  XNOR U9330 ( .A(n5070), .B(n8870), .Z(n8872) );
  NAND U9331 ( .A(n8875), .B(e_input[571]), .Z(n5070) );
  NAND U9332 ( .A(n6112), .B(e_input[571]), .Z(n8875) );
  XOR U9333 ( .A(n8876), .B(n8877), .Z(n8870) );
  ANDN U9334 ( .A(n8878), .B(n5071), .Z(n8877) );
  XOR U9335 ( .A(n8879), .B(n8880), .Z(n5071) );
  IV U9336 ( .A(n8876), .Z(n8879) );
  XNOR U9337 ( .A(n5072), .B(n8876), .Z(n8878) );
  NAND U9338 ( .A(n8881), .B(e_input[570]), .Z(n5072) );
  NAND U9339 ( .A(n6112), .B(e_input[570]), .Z(n8881) );
  XOR U9340 ( .A(n8882), .B(n8883), .Z(n8876) );
  ANDN U9341 ( .A(n8884), .B(n5075), .Z(n8883) );
  XOR U9342 ( .A(n8885), .B(n8886), .Z(n5075) );
  IV U9343 ( .A(n8882), .Z(n8885) );
  XNOR U9344 ( .A(n5076), .B(n8882), .Z(n8884) );
  NAND U9345 ( .A(n8887), .B(e_input[569]), .Z(n5076) );
  NAND U9346 ( .A(n6112), .B(e_input[569]), .Z(n8887) );
  XOR U9347 ( .A(n8888), .B(n8889), .Z(n8882) );
  ANDN U9348 ( .A(n8890), .B(n5077), .Z(n8889) );
  XOR U9349 ( .A(n8891), .B(n8892), .Z(n5077) );
  IV U9350 ( .A(n8888), .Z(n8891) );
  XNOR U9351 ( .A(n5078), .B(n8888), .Z(n8890) );
  NAND U9352 ( .A(n8893), .B(e_input[568]), .Z(n5078) );
  NAND U9353 ( .A(n6112), .B(e_input[568]), .Z(n8893) );
  XOR U9354 ( .A(n8894), .B(n8895), .Z(n8888) );
  ANDN U9355 ( .A(n8896), .B(n5079), .Z(n8895) );
  XOR U9356 ( .A(n8897), .B(n8898), .Z(n5079) );
  IV U9357 ( .A(n8894), .Z(n8897) );
  XNOR U9358 ( .A(n5080), .B(n8894), .Z(n8896) );
  NAND U9359 ( .A(n8899), .B(e_input[567]), .Z(n5080) );
  NAND U9360 ( .A(n6112), .B(e_input[567]), .Z(n8899) );
  XOR U9361 ( .A(n8900), .B(n8901), .Z(n8894) );
  ANDN U9362 ( .A(n8902), .B(n5081), .Z(n8901) );
  XOR U9363 ( .A(n8903), .B(n8904), .Z(n5081) );
  IV U9364 ( .A(n8900), .Z(n8903) );
  XNOR U9365 ( .A(n5082), .B(n8900), .Z(n8902) );
  NAND U9366 ( .A(n8905), .B(e_input[566]), .Z(n5082) );
  NAND U9367 ( .A(n6112), .B(e_input[566]), .Z(n8905) );
  XOR U9368 ( .A(n8906), .B(n8907), .Z(n8900) );
  ANDN U9369 ( .A(n8908), .B(n5083), .Z(n8907) );
  XOR U9370 ( .A(n8909), .B(n8910), .Z(n5083) );
  IV U9371 ( .A(n8906), .Z(n8909) );
  XNOR U9372 ( .A(n5084), .B(n8906), .Z(n8908) );
  NAND U9373 ( .A(n8911), .B(e_input[565]), .Z(n5084) );
  NAND U9374 ( .A(n6112), .B(e_input[565]), .Z(n8911) );
  XOR U9375 ( .A(n8912), .B(n8913), .Z(n8906) );
  ANDN U9376 ( .A(n8914), .B(n5085), .Z(n8913) );
  XOR U9377 ( .A(n8915), .B(n8916), .Z(n5085) );
  IV U9378 ( .A(n8912), .Z(n8915) );
  XNOR U9379 ( .A(n5086), .B(n8912), .Z(n8914) );
  NAND U9380 ( .A(n8917), .B(e_input[564]), .Z(n5086) );
  NAND U9381 ( .A(n6112), .B(e_input[564]), .Z(n8917) );
  XOR U9382 ( .A(n8918), .B(n8919), .Z(n8912) );
  ANDN U9383 ( .A(n8920), .B(n5087), .Z(n8919) );
  XOR U9384 ( .A(n8921), .B(n8922), .Z(n5087) );
  IV U9385 ( .A(n8918), .Z(n8921) );
  XNOR U9386 ( .A(n5088), .B(n8918), .Z(n8920) );
  NAND U9387 ( .A(n8923), .B(e_input[563]), .Z(n5088) );
  NAND U9388 ( .A(n6112), .B(e_input[563]), .Z(n8923) );
  XOR U9389 ( .A(n8924), .B(n8925), .Z(n8918) );
  ANDN U9390 ( .A(n8926), .B(n5089), .Z(n8925) );
  XOR U9391 ( .A(n8927), .B(n8928), .Z(n5089) );
  IV U9392 ( .A(n8924), .Z(n8927) );
  XNOR U9393 ( .A(n5090), .B(n8924), .Z(n8926) );
  NAND U9394 ( .A(n8929), .B(e_input[562]), .Z(n5090) );
  NAND U9395 ( .A(n6112), .B(e_input[562]), .Z(n8929) );
  XOR U9396 ( .A(n8930), .B(n8931), .Z(n8924) );
  ANDN U9397 ( .A(n8932), .B(n5091), .Z(n8931) );
  XOR U9398 ( .A(n8933), .B(n8934), .Z(n5091) );
  IV U9399 ( .A(n8930), .Z(n8933) );
  XNOR U9400 ( .A(n5092), .B(n8930), .Z(n8932) );
  NAND U9401 ( .A(n8935), .B(e_input[561]), .Z(n5092) );
  NAND U9402 ( .A(n6112), .B(e_input[561]), .Z(n8935) );
  XOR U9403 ( .A(n8936), .B(n8937), .Z(n8930) );
  ANDN U9404 ( .A(n8938), .B(n5093), .Z(n8937) );
  XOR U9405 ( .A(n8939), .B(n8940), .Z(n5093) );
  IV U9406 ( .A(n8936), .Z(n8939) );
  XNOR U9407 ( .A(n5094), .B(n8936), .Z(n8938) );
  NAND U9408 ( .A(n8941), .B(e_input[560]), .Z(n5094) );
  NAND U9409 ( .A(n6112), .B(e_input[560]), .Z(n8941) );
  XOR U9410 ( .A(n8942), .B(n8943), .Z(n8936) );
  ANDN U9411 ( .A(n8944), .B(n5097), .Z(n8943) );
  XOR U9412 ( .A(n8945), .B(n8946), .Z(n5097) );
  IV U9413 ( .A(n8942), .Z(n8945) );
  XNOR U9414 ( .A(n5098), .B(n8942), .Z(n8944) );
  NAND U9415 ( .A(n8947), .B(e_input[559]), .Z(n5098) );
  NAND U9416 ( .A(n6112), .B(e_input[559]), .Z(n8947) );
  XOR U9417 ( .A(n8948), .B(n8949), .Z(n8942) );
  ANDN U9418 ( .A(n8950), .B(n5099), .Z(n8949) );
  XOR U9419 ( .A(n8951), .B(n8952), .Z(n5099) );
  IV U9420 ( .A(n8948), .Z(n8951) );
  XNOR U9421 ( .A(n5100), .B(n8948), .Z(n8950) );
  NAND U9422 ( .A(n8953), .B(e_input[558]), .Z(n5100) );
  NAND U9423 ( .A(n6112), .B(e_input[558]), .Z(n8953) );
  XOR U9424 ( .A(n8954), .B(n8955), .Z(n8948) );
  ANDN U9425 ( .A(n8956), .B(n5101), .Z(n8955) );
  XOR U9426 ( .A(n8957), .B(n8958), .Z(n5101) );
  IV U9427 ( .A(n8954), .Z(n8957) );
  XNOR U9428 ( .A(n5102), .B(n8954), .Z(n8956) );
  NAND U9429 ( .A(n8959), .B(e_input[557]), .Z(n5102) );
  NAND U9430 ( .A(n6112), .B(e_input[557]), .Z(n8959) );
  XOR U9431 ( .A(n8960), .B(n8961), .Z(n8954) );
  ANDN U9432 ( .A(n8962), .B(n5103), .Z(n8961) );
  XOR U9433 ( .A(n8963), .B(n8964), .Z(n5103) );
  IV U9434 ( .A(n8960), .Z(n8963) );
  XNOR U9435 ( .A(n5104), .B(n8960), .Z(n8962) );
  NAND U9436 ( .A(n8965), .B(e_input[556]), .Z(n5104) );
  NAND U9437 ( .A(n6112), .B(e_input[556]), .Z(n8965) );
  XOR U9438 ( .A(n8966), .B(n8967), .Z(n8960) );
  ANDN U9439 ( .A(n8968), .B(n5105), .Z(n8967) );
  XOR U9440 ( .A(n8969), .B(n8970), .Z(n5105) );
  IV U9441 ( .A(n8966), .Z(n8969) );
  XNOR U9442 ( .A(n5106), .B(n8966), .Z(n8968) );
  NAND U9443 ( .A(n8971), .B(e_input[555]), .Z(n5106) );
  NAND U9444 ( .A(n6112), .B(e_input[555]), .Z(n8971) );
  XOR U9445 ( .A(n8972), .B(n8973), .Z(n8966) );
  ANDN U9446 ( .A(n8974), .B(n5107), .Z(n8973) );
  XOR U9447 ( .A(n8975), .B(n8976), .Z(n5107) );
  IV U9448 ( .A(n8972), .Z(n8975) );
  XNOR U9449 ( .A(n5108), .B(n8972), .Z(n8974) );
  NAND U9450 ( .A(n8977), .B(e_input[554]), .Z(n5108) );
  NAND U9451 ( .A(n6112), .B(e_input[554]), .Z(n8977) );
  XOR U9452 ( .A(n8978), .B(n8979), .Z(n8972) );
  ANDN U9453 ( .A(n8980), .B(n5109), .Z(n8979) );
  XOR U9454 ( .A(n8981), .B(n8982), .Z(n5109) );
  IV U9455 ( .A(n8978), .Z(n8981) );
  XNOR U9456 ( .A(n5110), .B(n8978), .Z(n8980) );
  NAND U9457 ( .A(n8983), .B(e_input[553]), .Z(n5110) );
  NAND U9458 ( .A(n6112), .B(e_input[553]), .Z(n8983) );
  XOR U9459 ( .A(n8984), .B(n8985), .Z(n8978) );
  ANDN U9460 ( .A(n8986), .B(n5111), .Z(n8985) );
  XOR U9461 ( .A(n8987), .B(n8988), .Z(n5111) );
  IV U9462 ( .A(n8984), .Z(n8987) );
  XNOR U9463 ( .A(n5112), .B(n8984), .Z(n8986) );
  NAND U9464 ( .A(n8989), .B(e_input[552]), .Z(n5112) );
  NAND U9465 ( .A(n6112), .B(e_input[552]), .Z(n8989) );
  XOR U9466 ( .A(n8990), .B(n8991), .Z(n8984) );
  ANDN U9467 ( .A(n8992), .B(n5113), .Z(n8991) );
  XOR U9468 ( .A(n8993), .B(n8994), .Z(n5113) );
  IV U9469 ( .A(n8990), .Z(n8993) );
  XNOR U9470 ( .A(n5114), .B(n8990), .Z(n8992) );
  NAND U9471 ( .A(n8995), .B(e_input[551]), .Z(n5114) );
  NAND U9472 ( .A(n6112), .B(e_input[551]), .Z(n8995) );
  XOR U9473 ( .A(n8996), .B(n8997), .Z(n8990) );
  ANDN U9474 ( .A(n8998), .B(n5115), .Z(n8997) );
  XOR U9475 ( .A(n8999), .B(n9000), .Z(n5115) );
  IV U9476 ( .A(n8996), .Z(n8999) );
  XNOR U9477 ( .A(n5116), .B(n8996), .Z(n8998) );
  NAND U9478 ( .A(n9001), .B(e_input[550]), .Z(n5116) );
  NAND U9479 ( .A(n6112), .B(e_input[550]), .Z(n9001) );
  XOR U9480 ( .A(n9002), .B(n9003), .Z(n8996) );
  ANDN U9481 ( .A(n9004), .B(n5119), .Z(n9003) );
  XOR U9482 ( .A(n9005), .B(n9006), .Z(n5119) );
  IV U9483 ( .A(n9002), .Z(n9005) );
  XNOR U9484 ( .A(n5120), .B(n9002), .Z(n9004) );
  NAND U9485 ( .A(n9007), .B(e_input[549]), .Z(n5120) );
  NAND U9486 ( .A(n6112), .B(e_input[549]), .Z(n9007) );
  XOR U9487 ( .A(n9008), .B(n9009), .Z(n9002) );
  ANDN U9488 ( .A(n9010), .B(n5121), .Z(n9009) );
  XOR U9489 ( .A(n9011), .B(n9012), .Z(n5121) );
  IV U9490 ( .A(n9008), .Z(n9011) );
  XNOR U9491 ( .A(n5122), .B(n9008), .Z(n9010) );
  NAND U9492 ( .A(n9013), .B(e_input[548]), .Z(n5122) );
  NAND U9493 ( .A(n6112), .B(e_input[548]), .Z(n9013) );
  XOR U9494 ( .A(n9014), .B(n9015), .Z(n9008) );
  ANDN U9495 ( .A(n9016), .B(n5123), .Z(n9015) );
  XOR U9496 ( .A(n9017), .B(n9018), .Z(n5123) );
  IV U9497 ( .A(n9014), .Z(n9017) );
  XNOR U9498 ( .A(n5124), .B(n9014), .Z(n9016) );
  NAND U9499 ( .A(n9019), .B(e_input[547]), .Z(n5124) );
  NAND U9500 ( .A(n6112), .B(e_input[547]), .Z(n9019) );
  XOR U9501 ( .A(n9020), .B(n9021), .Z(n9014) );
  ANDN U9502 ( .A(n9022), .B(n5125), .Z(n9021) );
  XOR U9503 ( .A(n9023), .B(n9024), .Z(n5125) );
  IV U9504 ( .A(n9020), .Z(n9023) );
  XNOR U9505 ( .A(n5126), .B(n9020), .Z(n9022) );
  NAND U9506 ( .A(n9025), .B(e_input[546]), .Z(n5126) );
  NAND U9507 ( .A(n6112), .B(e_input[546]), .Z(n9025) );
  XOR U9508 ( .A(n9026), .B(n9027), .Z(n9020) );
  ANDN U9509 ( .A(n9028), .B(n5127), .Z(n9027) );
  XOR U9510 ( .A(n9029), .B(n9030), .Z(n5127) );
  IV U9511 ( .A(n9026), .Z(n9029) );
  XNOR U9512 ( .A(n5128), .B(n9026), .Z(n9028) );
  NAND U9513 ( .A(n9031), .B(e_input[545]), .Z(n5128) );
  NAND U9514 ( .A(n6112), .B(e_input[545]), .Z(n9031) );
  XOR U9515 ( .A(n9032), .B(n9033), .Z(n9026) );
  ANDN U9516 ( .A(n9034), .B(n5129), .Z(n9033) );
  XOR U9517 ( .A(n9035), .B(n9036), .Z(n5129) );
  IV U9518 ( .A(n9032), .Z(n9035) );
  XNOR U9519 ( .A(n5130), .B(n9032), .Z(n9034) );
  NAND U9520 ( .A(n9037), .B(e_input[544]), .Z(n5130) );
  NAND U9521 ( .A(n6112), .B(e_input[544]), .Z(n9037) );
  XOR U9522 ( .A(n9038), .B(n9039), .Z(n9032) );
  ANDN U9523 ( .A(n9040), .B(n5131), .Z(n9039) );
  XOR U9524 ( .A(n9041), .B(n9042), .Z(n5131) );
  IV U9525 ( .A(n9038), .Z(n9041) );
  XNOR U9526 ( .A(n5132), .B(n9038), .Z(n9040) );
  NAND U9527 ( .A(n9043), .B(e_input[543]), .Z(n5132) );
  NAND U9528 ( .A(n6112), .B(e_input[543]), .Z(n9043) );
  XOR U9529 ( .A(n9044), .B(n9045), .Z(n9038) );
  ANDN U9530 ( .A(n9046), .B(n5133), .Z(n9045) );
  XOR U9531 ( .A(n9047), .B(n9048), .Z(n5133) );
  IV U9532 ( .A(n9044), .Z(n9047) );
  XNOR U9533 ( .A(n5134), .B(n9044), .Z(n9046) );
  NAND U9534 ( .A(n9049), .B(e_input[542]), .Z(n5134) );
  NAND U9535 ( .A(n6112), .B(e_input[542]), .Z(n9049) );
  XOR U9536 ( .A(n9050), .B(n9051), .Z(n9044) );
  ANDN U9537 ( .A(n9052), .B(n5135), .Z(n9051) );
  XOR U9538 ( .A(n9053), .B(n9054), .Z(n5135) );
  IV U9539 ( .A(n9050), .Z(n9053) );
  XNOR U9540 ( .A(n5136), .B(n9050), .Z(n9052) );
  NAND U9541 ( .A(n9055), .B(e_input[541]), .Z(n5136) );
  NAND U9542 ( .A(n6112), .B(e_input[541]), .Z(n9055) );
  XOR U9543 ( .A(n9056), .B(n9057), .Z(n9050) );
  ANDN U9544 ( .A(n9058), .B(n5137), .Z(n9057) );
  XOR U9545 ( .A(n9059), .B(n9060), .Z(n5137) );
  IV U9546 ( .A(n9056), .Z(n9059) );
  XNOR U9547 ( .A(n5138), .B(n9056), .Z(n9058) );
  NAND U9548 ( .A(n9061), .B(e_input[540]), .Z(n5138) );
  NAND U9549 ( .A(n6112), .B(e_input[540]), .Z(n9061) );
  XOR U9550 ( .A(n9062), .B(n9063), .Z(n9056) );
  ANDN U9551 ( .A(n9064), .B(n5141), .Z(n9063) );
  XOR U9552 ( .A(n9065), .B(n9066), .Z(n5141) );
  IV U9553 ( .A(n9062), .Z(n9065) );
  XNOR U9554 ( .A(n5142), .B(n9062), .Z(n9064) );
  NAND U9555 ( .A(n9067), .B(e_input[539]), .Z(n5142) );
  NAND U9556 ( .A(n6112), .B(e_input[539]), .Z(n9067) );
  XOR U9557 ( .A(n9068), .B(n9069), .Z(n9062) );
  ANDN U9558 ( .A(n9070), .B(n5143), .Z(n9069) );
  XOR U9559 ( .A(n9071), .B(n9072), .Z(n5143) );
  IV U9560 ( .A(n9068), .Z(n9071) );
  XNOR U9561 ( .A(n5144), .B(n9068), .Z(n9070) );
  NAND U9562 ( .A(n9073), .B(e_input[538]), .Z(n5144) );
  NAND U9563 ( .A(n6112), .B(e_input[538]), .Z(n9073) );
  XOR U9564 ( .A(n9074), .B(n9075), .Z(n9068) );
  ANDN U9565 ( .A(n9076), .B(n5145), .Z(n9075) );
  XOR U9566 ( .A(n9077), .B(n9078), .Z(n5145) );
  IV U9567 ( .A(n9074), .Z(n9077) );
  XNOR U9568 ( .A(n5146), .B(n9074), .Z(n9076) );
  NAND U9569 ( .A(n9079), .B(e_input[537]), .Z(n5146) );
  NAND U9570 ( .A(n6112), .B(e_input[537]), .Z(n9079) );
  XOR U9571 ( .A(n9080), .B(n9081), .Z(n9074) );
  ANDN U9572 ( .A(n9082), .B(n5147), .Z(n9081) );
  XOR U9573 ( .A(n9083), .B(n9084), .Z(n5147) );
  IV U9574 ( .A(n9080), .Z(n9083) );
  XNOR U9575 ( .A(n5148), .B(n9080), .Z(n9082) );
  NAND U9576 ( .A(n9085), .B(e_input[536]), .Z(n5148) );
  NAND U9577 ( .A(n6112), .B(e_input[536]), .Z(n9085) );
  XOR U9578 ( .A(n9086), .B(n9087), .Z(n9080) );
  ANDN U9579 ( .A(n9088), .B(n5149), .Z(n9087) );
  XOR U9580 ( .A(n9089), .B(n9090), .Z(n5149) );
  IV U9581 ( .A(n9086), .Z(n9089) );
  XNOR U9582 ( .A(n5150), .B(n9086), .Z(n9088) );
  NAND U9583 ( .A(n9091), .B(e_input[535]), .Z(n5150) );
  NAND U9584 ( .A(n6112), .B(e_input[535]), .Z(n9091) );
  XOR U9585 ( .A(n9092), .B(n9093), .Z(n9086) );
  ANDN U9586 ( .A(n9094), .B(n5151), .Z(n9093) );
  XOR U9587 ( .A(n9095), .B(n9096), .Z(n5151) );
  IV U9588 ( .A(n9092), .Z(n9095) );
  XNOR U9589 ( .A(n5152), .B(n9092), .Z(n9094) );
  NAND U9590 ( .A(n9097), .B(e_input[534]), .Z(n5152) );
  NAND U9591 ( .A(n6112), .B(e_input[534]), .Z(n9097) );
  XOR U9592 ( .A(n9098), .B(n9099), .Z(n9092) );
  ANDN U9593 ( .A(n9100), .B(n5153), .Z(n9099) );
  XOR U9594 ( .A(n9101), .B(n9102), .Z(n5153) );
  IV U9595 ( .A(n9098), .Z(n9101) );
  XNOR U9596 ( .A(n5154), .B(n9098), .Z(n9100) );
  NAND U9597 ( .A(n9103), .B(e_input[533]), .Z(n5154) );
  NAND U9598 ( .A(n6112), .B(e_input[533]), .Z(n9103) );
  XOR U9599 ( .A(n9104), .B(n9105), .Z(n9098) );
  ANDN U9600 ( .A(n9106), .B(n5155), .Z(n9105) );
  XOR U9601 ( .A(n9107), .B(n9108), .Z(n5155) );
  IV U9602 ( .A(n9104), .Z(n9107) );
  XNOR U9603 ( .A(n5156), .B(n9104), .Z(n9106) );
  NAND U9604 ( .A(n9109), .B(e_input[532]), .Z(n5156) );
  NAND U9605 ( .A(n6112), .B(e_input[532]), .Z(n9109) );
  XOR U9606 ( .A(n9110), .B(n9111), .Z(n9104) );
  ANDN U9607 ( .A(n9112), .B(n5157), .Z(n9111) );
  XOR U9608 ( .A(n9113), .B(n9114), .Z(n5157) );
  IV U9609 ( .A(n9110), .Z(n9113) );
  XNOR U9610 ( .A(n5158), .B(n9110), .Z(n9112) );
  NAND U9611 ( .A(n9115), .B(e_input[531]), .Z(n5158) );
  NAND U9612 ( .A(n6112), .B(e_input[531]), .Z(n9115) );
  XOR U9613 ( .A(n9116), .B(n9117), .Z(n9110) );
  ANDN U9614 ( .A(n9118), .B(n5159), .Z(n9117) );
  XOR U9615 ( .A(n9119), .B(n9120), .Z(n5159) );
  IV U9616 ( .A(n9116), .Z(n9119) );
  XNOR U9617 ( .A(n5160), .B(n9116), .Z(n9118) );
  NAND U9618 ( .A(n9121), .B(e_input[530]), .Z(n5160) );
  NAND U9619 ( .A(n6112), .B(e_input[530]), .Z(n9121) );
  XOR U9620 ( .A(n9122), .B(n9123), .Z(n9116) );
  ANDN U9621 ( .A(n9124), .B(n5163), .Z(n9123) );
  XOR U9622 ( .A(n9125), .B(n9126), .Z(n5163) );
  IV U9623 ( .A(n9122), .Z(n9125) );
  XNOR U9624 ( .A(n5164), .B(n9122), .Z(n9124) );
  NAND U9625 ( .A(n9127), .B(e_input[529]), .Z(n5164) );
  NAND U9626 ( .A(n6112), .B(e_input[529]), .Z(n9127) );
  XOR U9627 ( .A(n9128), .B(n9129), .Z(n9122) );
  ANDN U9628 ( .A(n9130), .B(n5165), .Z(n9129) );
  XOR U9629 ( .A(n9131), .B(n9132), .Z(n5165) );
  IV U9630 ( .A(n9128), .Z(n9131) );
  XNOR U9631 ( .A(n5166), .B(n9128), .Z(n9130) );
  NAND U9632 ( .A(n9133), .B(e_input[528]), .Z(n5166) );
  NAND U9633 ( .A(n6112), .B(e_input[528]), .Z(n9133) );
  XOR U9634 ( .A(n9134), .B(n9135), .Z(n9128) );
  ANDN U9635 ( .A(n9136), .B(n5167), .Z(n9135) );
  XOR U9636 ( .A(n9137), .B(n9138), .Z(n5167) );
  IV U9637 ( .A(n9134), .Z(n9137) );
  XNOR U9638 ( .A(n5168), .B(n9134), .Z(n9136) );
  NAND U9639 ( .A(n9139), .B(e_input[527]), .Z(n5168) );
  NAND U9640 ( .A(n6112), .B(e_input[527]), .Z(n9139) );
  XOR U9641 ( .A(n9140), .B(n9141), .Z(n9134) );
  ANDN U9642 ( .A(n9142), .B(n5169), .Z(n9141) );
  XOR U9643 ( .A(n9143), .B(n9144), .Z(n5169) );
  IV U9644 ( .A(n9140), .Z(n9143) );
  XNOR U9645 ( .A(n5170), .B(n9140), .Z(n9142) );
  NAND U9646 ( .A(n9145), .B(e_input[526]), .Z(n5170) );
  NAND U9647 ( .A(n6112), .B(e_input[526]), .Z(n9145) );
  XOR U9648 ( .A(n9146), .B(n9147), .Z(n9140) );
  ANDN U9649 ( .A(n9148), .B(n5171), .Z(n9147) );
  XOR U9650 ( .A(n9149), .B(n9150), .Z(n5171) );
  IV U9651 ( .A(n9146), .Z(n9149) );
  XNOR U9652 ( .A(n5172), .B(n9146), .Z(n9148) );
  NAND U9653 ( .A(n9151), .B(e_input[525]), .Z(n5172) );
  NAND U9654 ( .A(n6112), .B(e_input[525]), .Z(n9151) );
  XOR U9655 ( .A(n9152), .B(n9153), .Z(n9146) );
  ANDN U9656 ( .A(n9154), .B(n5173), .Z(n9153) );
  XOR U9657 ( .A(n9155), .B(n9156), .Z(n5173) );
  IV U9658 ( .A(n9152), .Z(n9155) );
  XNOR U9659 ( .A(n5174), .B(n9152), .Z(n9154) );
  NAND U9660 ( .A(n9157), .B(e_input[524]), .Z(n5174) );
  NAND U9661 ( .A(n6112), .B(e_input[524]), .Z(n9157) );
  XOR U9662 ( .A(n9158), .B(n9159), .Z(n9152) );
  ANDN U9663 ( .A(n9160), .B(n5175), .Z(n9159) );
  XOR U9664 ( .A(n9161), .B(n9162), .Z(n5175) );
  IV U9665 ( .A(n9158), .Z(n9161) );
  XNOR U9666 ( .A(n5176), .B(n9158), .Z(n9160) );
  NAND U9667 ( .A(n9163), .B(e_input[523]), .Z(n5176) );
  NAND U9668 ( .A(n6112), .B(e_input[523]), .Z(n9163) );
  XOR U9669 ( .A(n9164), .B(n9165), .Z(n9158) );
  ANDN U9670 ( .A(n9166), .B(n5177), .Z(n9165) );
  XOR U9671 ( .A(n9167), .B(n9168), .Z(n5177) );
  IV U9672 ( .A(n9164), .Z(n9167) );
  XNOR U9673 ( .A(n5178), .B(n9164), .Z(n9166) );
  NAND U9674 ( .A(n9169), .B(e_input[522]), .Z(n5178) );
  NAND U9675 ( .A(n6112), .B(e_input[522]), .Z(n9169) );
  XOR U9676 ( .A(n9170), .B(n9171), .Z(n9164) );
  ANDN U9677 ( .A(n9172), .B(n5179), .Z(n9171) );
  XOR U9678 ( .A(n9173), .B(n9174), .Z(n5179) );
  IV U9679 ( .A(n9170), .Z(n9173) );
  XNOR U9680 ( .A(n5180), .B(n9170), .Z(n9172) );
  NAND U9681 ( .A(n9175), .B(e_input[521]), .Z(n5180) );
  NAND U9682 ( .A(n6112), .B(e_input[521]), .Z(n9175) );
  XOR U9683 ( .A(n9176), .B(n9177), .Z(n9170) );
  ANDN U9684 ( .A(n9178), .B(n5181), .Z(n9177) );
  XOR U9685 ( .A(n9179), .B(n9180), .Z(n5181) );
  IV U9686 ( .A(n9176), .Z(n9179) );
  XNOR U9687 ( .A(n5182), .B(n9176), .Z(n9178) );
  NAND U9688 ( .A(n9181), .B(e_input[520]), .Z(n5182) );
  NAND U9689 ( .A(n6112), .B(e_input[520]), .Z(n9181) );
  XOR U9690 ( .A(n9182), .B(n9183), .Z(n9176) );
  ANDN U9691 ( .A(n9184), .B(n5185), .Z(n9183) );
  XOR U9692 ( .A(n9185), .B(n9186), .Z(n5185) );
  IV U9693 ( .A(n9182), .Z(n9185) );
  XNOR U9694 ( .A(n5186), .B(n9182), .Z(n9184) );
  NAND U9695 ( .A(n9187), .B(e_input[519]), .Z(n5186) );
  NAND U9696 ( .A(n6112), .B(e_input[519]), .Z(n9187) );
  XOR U9697 ( .A(n9188), .B(n9189), .Z(n9182) );
  ANDN U9698 ( .A(n9190), .B(n5187), .Z(n9189) );
  XOR U9699 ( .A(n9191), .B(n9192), .Z(n5187) );
  IV U9700 ( .A(n9188), .Z(n9191) );
  XNOR U9701 ( .A(n5188), .B(n9188), .Z(n9190) );
  NAND U9702 ( .A(n9193), .B(e_input[518]), .Z(n5188) );
  NAND U9703 ( .A(n6112), .B(e_input[518]), .Z(n9193) );
  XOR U9704 ( .A(n9194), .B(n9195), .Z(n9188) );
  ANDN U9705 ( .A(n9196), .B(n5189), .Z(n9195) );
  XOR U9706 ( .A(n9197), .B(n9198), .Z(n5189) );
  IV U9707 ( .A(n9194), .Z(n9197) );
  XNOR U9708 ( .A(n5190), .B(n9194), .Z(n9196) );
  NAND U9709 ( .A(n9199), .B(e_input[517]), .Z(n5190) );
  NAND U9710 ( .A(n6112), .B(e_input[517]), .Z(n9199) );
  XOR U9711 ( .A(n9200), .B(n9201), .Z(n9194) );
  ANDN U9712 ( .A(n9202), .B(n5191), .Z(n9201) );
  XOR U9713 ( .A(n9203), .B(n9204), .Z(n5191) );
  IV U9714 ( .A(n9200), .Z(n9203) );
  XNOR U9715 ( .A(n5192), .B(n9200), .Z(n9202) );
  NAND U9716 ( .A(n9205), .B(e_input[516]), .Z(n5192) );
  NAND U9717 ( .A(n6112), .B(e_input[516]), .Z(n9205) );
  XOR U9718 ( .A(n9206), .B(n9207), .Z(n9200) );
  ANDN U9719 ( .A(n9208), .B(n5193), .Z(n9207) );
  XOR U9720 ( .A(n9209), .B(n9210), .Z(n5193) );
  IV U9721 ( .A(n9206), .Z(n9209) );
  XNOR U9722 ( .A(n5194), .B(n9206), .Z(n9208) );
  NAND U9723 ( .A(n9211), .B(e_input[515]), .Z(n5194) );
  NAND U9724 ( .A(n6112), .B(e_input[515]), .Z(n9211) );
  XOR U9725 ( .A(n9212), .B(n9213), .Z(n9206) );
  ANDN U9726 ( .A(n9214), .B(n5195), .Z(n9213) );
  XOR U9727 ( .A(n9215), .B(n9216), .Z(n5195) );
  IV U9728 ( .A(n9212), .Z(n9215) );
  XNOR U9729 ( .A(n5196), .B(n9212), .Z(n9214) );
  NAND U9730 ( .A(n9217), .B(e_input[514]), .Z(n5196) );
  NAND U9731 ( .A(n6112), .B(e_input[514]), .Z(n9217) );
  XOR U9732 ( .A(n9218), .B(n9219), .Z(n9212) );
  ANDN U9733 ( .A(n9220), .B(n5197), .Z(n9219) );
  XOR U9734 ( .A(n9221), .B(n9222), .Z(n5197) );
  IV U9735 ( .A(n9218), .Z(n9221) );
  XNOR U9736 ( .A(n5198), .B(n9218), .Z(n9220) );
  NAND U9737 ( .A(n9223), .B(e_input[513]), .Z(n5198) );
  NAND U9738 ( .A(n6112), .B(e_input[513]), .Z(n9223) );
  XOR U9739 ( .A(n9224), .B(n9225), .Z(n9218) );
  ANDN U9740 ( .A(n9226), .B(n5199), .Z(n9225) );
  XOR U9741 ( .A(n9227), .B(n9228), .Z(n5199) );
  IV U9742 ( .A(n9224), .Z(n9227) );
  XNOR U9743 ( .A(n5200), .B(n9224), .Z(n9226) );
  NAND U9744 ( .A(n9229), .B(e_input[512]), .Z(n5200) );
  NAND U9745 ( .A(n6112), .B(e_input[512]), .Z(n9229) );
  XOR U9746 ( .A(n9230), .B(n9231), .Z(n9224) );
  ANDN U9747 ( .A(n9232), .B(n5201), .Z(n9231) );
  XOR U9748 ( .A(n9233), .B(n9234), .Z(n5201) );
  IV U9749 ( .A(n9230), .Z(n9233) );
  XNOR U9750 ( .A(n5202), .B(n9230), .Z(n9232) );
  NAND U9751 ( .A(n9235), .B(e_input[511]), .Z(n5202) );
  NAND U9752 ( .A(n6112), .B(e_input[511]), .Z(n9235) );
  XOR U9753 ( .A(n9236), .B(n9237), .Z(n9230) );
  ANDN U9754 ( .A(n9238), .B(n5203), .Z(n9237) );
  XOR U9755 ( .A(n9239), .B(n9240), .Z(n5203) );
  IV U9756 ( .A(n9236), .Z(n9239) );
  XNOR U9757 ( .A(n5204), .B(n9236), .Z(n9238) );
  NAND U9758 ( .A(n9241), .B(e_input[510]), .Z(n5204) );
  NAND U9759 ( .A(n6112), .B(e_input[510]), .Z(n9241) );
  XOR U9760 ( .A(n9242), .B(n9243), .Z(n9236) );
  ANDN U9761 ( .A(n9244), .B(n5207), .Z(n9243) );
  XOR U9762 ( .A(n9245), .B(n9246), .Z(n5207) );
  IV U9763 ( .A(n9242), .Z(n9245) );
  XNOR U9764 ( .A(n5208), .B(n9242), .Z(n9244) );
  NAND U9765 ( .A(n9247), .B(e_input[509]), .Z(n5208) );
  NAND U9766 ( .A(n6112), .B(e_input[509]), .Z(n9247) );
  XOR U9767 ( .A(n9248), .B(n9249), .Z(n9242) );
  ANDN U9768 ( .A(n9250), .B(n5209), .Z(n9249) );
  XOR U9769 ( .A(n9251), .B(n9252), .Z(n5209) );
  IV U9770 ( .A(n9248), .Z(n9251) );
  XNOR U9771 ( .A(n5210), .B(n9248), .Z(n9250) );
  NAND U9772 ( .A(n9253), .B(e_input[508]), .Z(n5210) );
  NAND U9773 ( .A(n6112), .B(e_input[508]), .Z(n9253) );
  XOR U9774 ( .A(n9254), .B(n9255), .Z(n9248) );
  ANDN U9775 ( .A(n9256), .B(n5211), .Z(n9255) );
  XOR U9776 ( .A(n9257), .B(n9258), .Z(n5211) );
  IV U9777 ( .A(n9254), .Z(n9257) );
  XNOR U9778 ( .A(n5212), .B(n9254), .Z(n9256) );
  NAND U9779 ( .A(n9259), .B(e_input[507]), .Z(n5212) );
  NAND U9780 ( .A(n6112), .B(e_input[507]), .Z(n9259) );
  XOR U9781 ( .A(n9260), .B(n9261), .Z(n9254) );
  ANDN U9782 ( .A(n9262), .B(n5213), .Z(n9261) );
  XOR U9783 ( .A(n9263), .B(n9264), .Z(n5213) );
  IV U9784 ( .A(n9260), .Z(n9263) );
  XNOR U9785 ( .A(n5214), .B(n9260), .Z(n9262) );
  NAND U9786 ( .A(n9265), .B(e_input[506]), .Z(n5214) );
  NAND U9787 ( .A(n6112), .B(e_input[506]), .Z(n9265) );
  XOR U9788 ( .A(n9266), .B(n9267), .Z(n9260) );
  ANDN U9789 ( .A(n9268), .B(n5215), .Z(n9267) );
  XOR U9790 ( .A(n9269), .B(n9270), .Z(n5215) );
  IV U9791 ( .A(n9266), .Z(n9269) );
  XNOR U9792 ( .A(n5216), .B(n9266), .Z(n9268) );
  NAND U9793 ( .A(n9271), .B(e_input[505]), .Z(n5216) );
  NAND U9794 ( .A(n6112), .B(e_input[505]), .Z(n9271) );
  XOR U9795 ( .A(n9272), .B(n9273), .Z(n9266) );
  ANDN U9796 ( .A(n9274), .B(n5217), .Z(n9273) );
  XOR U9797 ( .A(n9275), .B(n9276), .Z(n5217) );
  IV U9798 ( .A(n9272), .Z(n9275) );
  XNOR U9799 ( .A(n5218), .B(n9272), .Z(n9274) );
  NAND U9800 ( .A(n9277), .B(e_input[504]), .Z(n5218) );
  NAND U9801 ( .A(n6112), .B(e_input[504]), .Z(n9277) );
  XOR U9802 ( .A(n9278), .B(n9279), .Z(n9272) );
  ANDN U9803 ( .A(n9280), .B(n5219), .Z(n9279) );
  XOR U9804 ( .A(n9281), .B(n9282), .Z(n5219) );
  IV U9805 ( .A(n9278), .Z(n9281) );
  XNOR U9806 ( .A(n5220), .B(n9278), .Z(n9280) );
  NAND U9807 ( .A(n9283), .B(e_input[503]), .Z(n5220) );
  NAND U9808 ( .A(n6112), .B(e_input[503]), .Z(n9283) );
  XOR U9809 ( .A(n9284), .B(n9285), .Z(n9278) );
  ANDN U9810 ( .A(n9286), .B(n5221), .Z(n9285) );
  XOR U9811 ( .A(n9287), .B(n9288), .Z(n5221) );
  IV U9812 ( .A(n9284), .Z(n9287) );
  XNOR U9813 ( .A(n5222), .B(n9284), .Z(n9286) );
  NAND U9814 ( .A(n9289), .B(e_input[502]), .Z(n5222) );
  NAND U9815 ( .A(n6112), .B(e_input[502]), .Z(n9289) );
  XOR U9816 ( .A(n9290), .B(n9291), .Z(n9284) );
  ANDN U9817 ( .A(n9292), .B(n5223), .Z(n9291) );
  XOR U9818 ( .A(n9293), .B(n9294), .Z(n5223) );
  IV U9819 ( .A(n9290), .Z(n9293) );
  XNOR U9820 ( .A(n5224), .B(n9290), .Z(n9292) );
  NAND U9821 ( .A(n9295), .B(e_input[501]), .Z(n5224) );
  NAND U9822 ( .A(n6112), .B(e_input[501]), .Z(n9295) );
  XOR U9823 ( .A(n9296), .B(n9297), .Z(n9290) );
  ANDN U9824 ( .A(n9298), .B(n5225), .Z(n9297) );
  XOR U9825 ( .A(n9299), .B(n9300), .Z(n5225) );
  IV U9826 ( .A(n9296), .Z(n9299) );
  XNOR U9827 ( .A(n5226), .B(n9296), .Z(n9298) );
  NAND U9828 ( .A(n9301), .B(e_input[500]), .Z(n5226) );
  NAND U9829 ( .A(n6112), .B(e_input[500]), .Z(n9301) );
  XOR U9830 ( .A(n9302), .B(n9303), .Z(n9296) );
  ANDN U9831 ( .A(n9304), .B(n5231), .Z(n9303) );
  XOR U9832 ( .A(n9305), .B(n9306), .Z(n5231) );
  IV U9833 ( .A(n9302), .Z(n9305) );
  XNOR U9834 ( .A(n5232), .B(n9302), .Z(n9304) );
  NAND U9835 ( .A(n9307), .B(e_input[499]), .Z(n5232) );
  NAND U9836 ( .A(n6112), .B(e_input[499]), .Z(n9307) );
  XOR U9837 ( .A(n9308), .B(n9309), .Z(n9302) );
  ANDN U9838 ( .A(n9310), .B(n5233), .Z(n9309) );
  XOR U9839 ( .A(n9311), .B(n9312), .Z(n5233) );
  IV U9840 ( .A(n9308), .Z(n9311) );
  XNOR U9841 ( .A(n5234), .B(n9308), .Z(n9310) );
  NAND U9842 ( .A(n9313), .B(e_input[498]), .Z(n5234) );
  NAND U9843 ( .A(n6112), .B(e_input[498]), .Z(n9313) );
  XOR U9844 ( .A(n9314), .B(n9315), .Z(n9308) );
  ANDN U9845 ( .A(n9316), .B(n5235), .Z(n9315) );
  XOR U9846 ( .A(n9317), .B(n9318), .Z(n5235) );
  IV U9847 ( .A(n9314), .Z(n9317) );
  XNOR U9848 ( .A(n5236), .B(n9314), .Z(n9316) );
  NAND U9849 ( .A(n9319), .B(e_input[497]), .Z(n5236) );
  NAND U9850 ( .A(n6112), .B(e_input[497]), .Z(n9319) );
  XOR U9851 ( .A(n9320), .B(n9321), .Z(n9314) );
  ANDN U9852 ( .A(n9322), .B(n5237), .Z(n9321) );
  XOR U9853 ( .A(n9323), .B(n9324), .Z(n5237) );
  IV U9854 ( .A(n9320), .Z(n9323) );
  XNOR U9855 ( .A(n5238), .B(n9320), .Z(n9322) );
  NAND U9856 ( .A(n9325), .B(e_input[496]), .Z(n5238) );
  NAND U9857 ( .A(n6112), .B(e_input[496]), .Z(n9325) );
  XOR U9858 ( .A(n9326), .B(n9327), .Z(n9320) );
  ANDN U9859 ( .A(n9328), .B(n5239), .Z(n9327) );
  XOR U9860 ( .A(n9329), .B(n9330), .Z(n5239) );
  IV U9861 ( .A(n9326), .Z(n9329) );
  XNOR U9862 ( .A(n5240), .B(n9326), .Z(n9328) );
  NAND U9863 ( .A(n9331), .B(e_input[495]), .Z(n5240) );
  NAND U9864 ( .A(n6112), .B(e_input[495]), .Z(n9331) );
  XOR U9865 ( .A(n9332), .B(n9333), .Z(n9326) );
  ANDN U9866 ( .A(n9334), .B(n5241), .Z(n9333) );
  XOR U9867 ( .A(n9335), .B(n9336), .Z(n5241) );
  IV U9868 ( .A(n9332), .Z(n9335) );
  XNOR U9869 ( .A(n5242), .B(n9332), .Z(n9334) );
  NAND U9870 ( .A(n9337), .B(e_input[494]), .Z(n5242) );
  NAND U9871 ( .A(n6112), .B(e_input[494]), .Z(n9337) );
  XOR U9872 ( .A(n9338), .B(n9339), .Z(n9332) );
  ANDN U9873 ( .A(n9340), .B(n5243), .Z(n9339) );
  XOR U9874 ( .A(n9341), .B(n9342), .Z(n5243) );
  IV U9875 ( .A(n9338), .Z(n9341) );
  XNOR U9876 ( .A(n5244), .B(n9338), .Z(n9340) );
  NAND U9877 ( .A(n9343), .B(e_input[493]), .Z(n5244) );
  NAND U9878 ( .A(n6112), .B(e_input[493]), .Z(n9343) );
  XOR U9879 ( .A(n9344), .B(n9345), .Z(n9338) );
  ANDN U9880 ( .A(n9346), .B(n5245), .Z(n9345) );
  XOR U9881 ( .A(n9347), .B(n9348), .Z(n5245) );
  IV U9882 ( .A(n9344), .Z(n9347) );
  XNOR U9883 ( .A(n5246), .B(n9344), .Z(n9346) );
  NAND U9884 ( .A(n9349), .B(e_input[492]), .Z(n5246) );
  NAND U9885 ( .A(n6112), .B(e_input[492]), .Z(n9349) );
  XOR U9886 ( .A(n9350), .B(n9351), .Z(n9344) );
  ANDN U9887 ( .A(n9352), .B(n5247), .Z(n9351) );
  XOR U9888 ( .A(n9353), .B(n9354), .Z(n5247) );
  IV U9889 ( .A(n9350), .Z(n9353) );
  XNOR U9890 ( .A(n5248), .B(n9350), .Z(n9352) );
  NAND U9891 ( .A(n9355), .B(e_input[491]), .Z(n5248) );
  NAND U9892 ( .A(n6112), .B(e_input[491]), .Z(n9355) );
  XOR U9893 ( .A(n9356), .B(n9357), .Z(n9350) );
  ANDN U9894 ( .A(n9358), .B(n5249), .Z(n9357) );
  XOR U9895 ( .A(n9359), .B(n9360), .Z(n5249) );
  IV U9896 ( .A(n9356), .Z(n9359) );
  XNOR U9897 ( .A(n5250), .B(n9356), .Z(n9358) );
  NAND U9898 ( .A(n9361), .B(e_input[490]), .Z(n5250) );
  NAND U9899 ( .A(n6112), .B(e_input[490]), .Z(n9361) );
  XOR U9900 ( .A(n9362), .B(n9363), .Z(n9356) );
  ANDN U9901 ( .A(n9364), .B(n5253), .Z(n9363) );
  XOR U9902 ( .A(n9365), .B(n9366), .Z(n5253) );
  IV U9903 ( .A(n9362), .Z(n9365) );
  XNOR U9904 ( .A(n5254), .B(n9362), .Z(n9364) );
  NAND U9905 ( .A(n9367), .B(e_input[489]), .Z(n5254) );
  NAND U9906 ( .A(n6112), .B(e_input[489]), .Z(n9367) );
  XOR U9907 ( .A(n9368), .B(n9369), .Z(n9362) );
  ANDN U9908 ( .A(n9370), .B(n5255), .Z(n9369) );
  XOR U9909 ( .A(n9371), .B(n9372), .Z(n5255) );
  IV U9910 ( .A(n9368), .Z(n9371) );
  XNOR U9911 ( .A(n5256), .B(n9368), .Z(n9370) );
  NAND U9912 ( .A(n9373), .B(e_input[488]), .Z(n5256) );
  NAND U9913 ( .A(n6112), .B(e_input[488]), .Z(n9373) );
  XOR U9914 ( .A(n9374), .B(n9375), .Z(n9368) );
  ANDN U9915 ( .A(n9376), .B(n5257), .Z(n9375) );
  XOR U9916 ( .A(n9377), .B(n9378), .Z(n5257) );
  IV U9917 ( .A(n9374), .Z(n9377) );
  XNOR U9918 ( .A(n5258), .B(n9374), .Z(n9376) );
  NAND U9919 ( .A(n9379), .B(e_input[487]), .Z(n5258) );
  NAND U9920 ( .A(n6112), .B(e_input[487]), .Z(n9379) );
  XOR U9921 ( .A(n9380), .B(n9381), .Z(n9374) );
  ANDN U9922 ( .A(n9382), .B(n5259), .Z(n9381) );
  XOR U9923 ( .A(n9383), .B(n9384), .Z(n5259) );
  IV U9924 ( .A(n9380), .Z(n9383) );
  XNOR U9925 ( .A(n5260), .B(n9380), .Z(n9382) );
  NAND U9926 ( .A(n9385), .B(e_input[486]), .Z(n5260) );
  NAND U9927 ( .A(n6112), .B(e_input[486]), .Z(n9385) );
  XOR U9928 ( .A(n9386), .B(n9387), .Z(n9380) );
  ANDN U9929 ( .A(n9388), .B(n5261), .Z(n9387) );
  XOR U9930 ( .A(n9389), .B(n9390), .Z(n5261) );
  IV U9931 ( .A(n9386), .Z(n9389) );
  XNOR U9932 ( .A(n5262), .B(n9386), .Z(n9388) );
  NAND U9933 ( .A(n9391), .B(e_input[485]), .Z(n5262) );
  NAND U9934 ( .A(n6112), .B(e_input[485]), .Z(n9391) );
  XOR U9935 ( .A(n9392), .B(n9393), .Z(n9386) );
  ANDN U9936 ( .A(n9394), .B(n5263), .Z(n9393) );
  XOR U9937 ( .A(n9395), .B(n9396), .Z(n5263) );
  IV U9938 ( .A(n9392), .Z(n9395) );
  XNOR U9939 ( .A(n5264), .B(n9392), .Z(n9394) );
  NAND U9940 ( .A(n9397), .B(e_input[484]), .Z(n5264) );
  NAND U9941 ( .A(n6112), .B(e_input[484]), .Z(n9397) );
  XOR U9942 ( .A(n9398), .B(n9399), .Z(n9392) );
  ANDN U9943 ( .A(n9400), .B(n5265), .Z(n9399) );
  XOR U9944 ( .A(n9401), .B(n9402), .Z(n5265) );
  IV U9945 ( .A(n9398), .Z(n9401) );
  XNOR U9946 ( .A(n5266), .B(n9398), .Z(n9400) );
  NAND U9947 ( .A(n9403), .B(e_input[483]), .Z(n5266) );
  NAND U9948 ( .A(n6112), .B(e_input[483]), .Z(n9403) );
  XOR U9949 ( .A(n9404), .B(n9405), .Z(n9398) );
  ANDN U9950 ( .A(n9406), .B(n5267), .Z(n9405) );
  XOR U9951 ( .A(n9407), .B(n9408), .Z(n5267) );
  IV U9952 ( .A(n9404), .Z(n9407) );
  XNOR U9953 ( .A(n5268), .B(n9404), .Z(n9406) );
  NAND U9954 ( .A(n9409), .B(e_input[482]), .Z(n5268) );
  NAND U9955 ( .A(n6112), .B(e_input[482]), .Z(n9409) );
  XOR U9956 ( .A(n9410), .B(n9411), .Z(n9404) );
  ANDN U9957 ( .A(n9412), .B(n5269), .Z(n9411) );
  XOR U9958 ( .A(n9413), .B(n9414), .Z(n5269) );
  IV U9959 ( .A(n9410), .Z(n9413) );
  XNOR U9960 ( .A(n5270), .B(n9410), .Z(n9412) );
  NAND U9961 ( .A(n9415), .B(e_input[481]), .Z(n5270) );
  NAND U9962 ( .A(n6112), .B(e_input[481]), .Z(n9415) );
  XOR U9963 ( .A(n9416), .B(n9417), .Z(n9410) );
  ANDN U9964 ( .A(n9418), .B(n5271), .Z(n9417) );
  XOR U9965 ( .A(n9419), .B(n9420), .Z(n5271) );
  IV U9966 ( .A(n9416), .Z(n9419) );
  XNOR U9967 ( .A(n5272), .B(n9416), .Z(n9418) );
  NAND U9968 ( .A(n9421), .B(e_input[480]), .Z(n5272) );
  NAND U9969 ( .A(n6112), .B(e_input[480]), .Z(n9421) );
  XOR U9970 ( .A(n9422), .B(n9423), .Z(n9416) );
  ANDN U9971 ( .A(n9424), .B(n5275), .Z(n9423) );
  XOR U9972 ( .A(n9425), .B(n9426), .Z(n5275) );
  IV U9973 ( .A(n9422), .Z(n9425) );
  XNOR U9974 ( .A(n5276), .B(n9422), .Z(n9424) );
  NAND U9975 ( .A(n9427), .B(e_input[479]), .Z(n5276) );
  NAND U9976 ( .A(n6112), .B(e_input[479]), .Z(n9427) );
  XOR U9977 ( .A(n9428), .B(n9429), .Z(n9422) );
  ANDN U9978 ( .A(n9430), .B(n5277), .Z(n9429) );
  XOR U9979 ( .A(n9431), .B(n9432), .Z(n5277) );
  IV U9980 ( .A(n9428), .Z(n9431) );
  XNOR U9981 ( .A(n5278), .B(n9428), .Z(n9430) );
  NAND U9982 ( .A(n9433), .B(e_input[478]), .Z(n5278) );
  NAND U9983 ( .A(n6112), .B(e_input[478]), .Z(n9433) );
  XOR U9984 ( .A(n9434), .B(n9435), .Z(n9428) );
  ANDN U9985 ( .A(n9436), .B(n5279), .Z(n9435) );
  XOR U9986 ( .A(n9437), .B(n9438), .Z(n5279) );
  IV U9987 ( .A(n9434), .Z(n9437) );
  XNOR U9988 ( .A(n5280), .B(n9434), .Z(n9436) );
  NAND U9989 ( .A(n9439), .B(e_input[477]), .Z(n5280) );
  NAND U9990 ( .A(n6112), .B(e_input[477]), .Z(n9439) );
  XOR U9991 ( .A(n9440), .B(n9441), .Z(n9434) );
  ANDN U9992 ( .A(n9442), .B(n5281), .Z(n9441) );
  XOR U9993 ( .A(n9443), .B(n9444), .Z(n5281) );
  IV U9994 ( .A(n9440), .Z(n9443) );
  XNOR U9995 ( .A(n5282), .B(n9440), .Z(n9442) );
  NAND U9996 ( .A(n9445), .B(e_input[476]), .Z(n5282) );
  NAND U9997 ( .A(n6112), .B(e_input[476]), .Z(n9445) );
  XOR U9998 ( .A(n9446), .B(n9447), .Z(n9440) );
  ANDN U9999 ( .A(n9448), .B(n5283), .Z(n9447) );
  XOR U10000 ( .A(n9449), .B(n9450), .Z(n5283) );
  IV U10001 ( .A(n9446), .Z(n9449) );
  XNOR U10002 ( .A(n5284), .B(n9446), .Z(n9448) );
  NAND U10003 ( .A(n9451), .B(e_input[475]), .Z(n5284) );
  NAND U10004 ( .A(n6112), .B(e_input[475]), .Z(n9451) );
  XOR U10005 ( .A(n9452), .B(n9453), .Z(n9446) );
  ANDN U10006 ( .A(n9454), .B(n5285), .Z(n9453) );
  XOR U10007 ( .A(n9455), .B(n9456), .Z(n5285) );
  IV U10008 ( .A(n9452), .Z(n9455) );
  XNOR U10009 ( .A(n5286), .B(n9452), .Z(n9454) );
  NAND U10010 ( .A(n9457), .B(e_input[474]), .Z(n5286) );
  NAND U10011 ( .A(n6112), .B(e_input[474]), .Z(n9457) );
  XOR U10012 ( .A(n9458), .B(n9459), .Z(n9452) );
  ANDN U10013 ( .A(n9460), .B(n5287), .Z(n9459) );
  XOR U10014 ( .A(n9461), .B(n9462), .Z(n5287) );
  IV U10015 ( .A(n9458), .Z(n9461) );
  XNOR U10016 ( .A(n5288), .B(n9458), .Z(n9460) );
  NAND U10017 ( .A(n9463), .B(e_input[473]), .Z(n5288) );
  NAND U10018 ( .A(n6112), .B(e_input[473]), .Z(n9463) );
  XOR U10019 ( .A(n9464), .B(n9465), .Z(n9458) );
  ANDN U10020 ( .A(n9466), .B(n5289), .Z(n9465) );
  XOR U10021 ( .A(n9467), .B(n9468), .Z(n5289) );
  IV U10022 ( .A(n9464), .Z(n9467) );
  XNOR U10023 ( .A(n5290), .B(n9464), .Z(n9466) );
  NAND U10024 ( .A(n9469), .B(e_input[472]), .Z(n5290) );
  NAND U10025 ( .A(n6112), .B(e_input[472]), .Z(n9469) );
  XOR U10026 ( .A(n9470), .B(n9471), .Z(n9464) );
  ANDN U10027 ( .A(n9472), .B(n5291), .Z(n9471) );
  XOR U10028 ( .A(n9473), .B(n9474), .Z(n5291) );
  IV U10029 ( .A(n9470), .Z(n9473) );
  XNOR U10030 ( .A(n5292), .B(n9470), .Z(n9472) );
  NAND U10031 ( .A(n9475), .B(e_input[471]), .Z(n5292) );
  NAND U10032 ( .A(n6112), .B(e_input[471]), .Z(n9475) );
  XOR U10033 ( .A(n9476), .B(n9477), .Z(n9470) );
  ANDN U10034 ( .A(n9478), .B(n5293), .Z(n9477) );
  XOR U10035 ( .A(n9479), .B(n9480), .Z(n5293) );
  IV U10036 ( .A(n9476), .Z(n9479) );
  XNOR U10037 ( .A(n5294), .B(n9476), .Z(n9478) );
  NAND U10038 ( .A(n9481), .B(e_input[470]), .Z(n5294) );
  NAND U10039 ( .A(n6112), .B(e_input[470]), .Z(n9481) );
  XOR U10040 ( .A(n9482), .B(n9483), .Z(n9476) );
  ANDN U10041 ( .A(n9484), .B(n5297), .Z(n9483) );
  XOR U10042 ( .A(n9485), .B(n9486), .Z(n5297) );
  IV U10043 ( .A(n9482), .Z(n9485) );
  XNOR U10044 ( .A(n5298), .B(n9482), .Z(n9484) );
  NAND U10045 ( .A(n9487), .B(e_input[469]), .Z(n5298) );
  NAND U10046 ( .A(n6112), .B(e_input[469]), .Z(n9487) );
  XOR U10047 ( .A(n9488), .B(n9489), .Z(n9482) );
  ANDN U10048 ( .A(n9490), .B(n5299), .Z(n9489) );
  XOR U10049 ( .A(n9491), .B(n9492), .Z(n5299) );
  IV U10050 ( .A(n9488), .Z(n9491) );
  XNOR U10051 ( .A(n5300), .B(n9488), .Z(n9490) );
  NAND U10052 ( .A(n9493), .B(e_input[468]), .Z(n5300) );
  NAND U10053 ( .A(n6112), .B(e_input[468]), .Z(n9493) );
  XOR U10054 ( .A(n9494), .B(n9495), .Z(n9488) );
  ANDN U10055 ( .A(n9496), .B(n5301), .Z(n9495) );
  XOR U10056 ( .A(n9497), .B(n9498), .Z(n5301) );
  IV U10057 ( .A(n9494), .Z(n9497) );
  XNOR U10058 ( .A(n5302), .B(n9494), .Z(n9496) );
  NAND U10059 ( .A(n9499), .B(e_input[467]), .Z(n5302) );
  NAND U10060 ( .A(n6112), .B(e_input[467]), .Z(n9499) );
  XOR U10061 ( .A(n9500), .B(n9501), .Z(n9494) );
  ANDN U10062 ( .A(n9502), .B(n5303), .Z(n9501) );
  XOR U10063 ( .A(n9503), .B(n9504), .Z(n5303) );
  IV U10064 ( .A(n9500), .Z(n9503) );
  XNOR U10065 ( .A(n5304), .B(n9500), .Z(n9502) );
  NAND U10066 ( .A(n9505), .B(e_input[466]), .Z(n5304) );
  NAND U10067 ( .A(n6112), .B(e_input[466]), .Z(n9505) );
  XOR U10068 ( .A(n9506), .B(n9507), .Z(n9500) );
  ANDN U10069 ( .A(n9508), .B(n5305), .Z(n9507) );
  XOR U10070 ( .A(n9509), .B(n9510), .Z(n5305) );
  IV U10071 ( .A(n9506), .Z(n9509) );
  XNOR U10072 ( .A(n5306), .B(n9506), .Z(n9508) );
  NAND U10073 ( .A(n9511), .B(e_input[465]), .Z(n5306) );
  NAND U10074 ( .A(n6112), .B(e_input[465]), .Z(n9511) );
  XOR U10075 ( .A(n9512), .B(n9513), .Z(n9506) );
  ANDN U10076 ( .A(n9514), .B(n5307), .Z(n9513) );
  XOR U10077 ( .A(n9515), .B(n9516), .Z(n5307) );
  IV U10078 ( .A(n9512), .Z(n9515) );
  XNOR U10079 ( .A(n5308), .B(n9512), .Z(n9514) );
  NAND U10080 ( .A(n9517), .B(e_input[464]), .Z(n5308) );
  NAND U10081 ( .A(n6112), .B(e_input[464]), .Z(n9517) );
  XOR U10082 ( .A(n9518), .B(n9519), .Z(n9512) );
  ANDN U10083 ( .A(n9520), .B(n5309), .Z(n9519) );
  XOR U10084 ( .A(n9521), .B(n9522), .Z(n5309) );
  IV U10085 ( .A(n9518), .Z(n9521) );
  XNOR U10086 ( .A(n5310), .B(n9518), .Z(n9520) );
  NAND U10087 ( .A(n9523), .B(e_input[463]), .Z(n5310) );
  NAND U10088 ( .A(n6112), .B(e_input[463]), .Z(n9523) );
  XOR U10089 ( .A(n9524), .B(n9525), .Z(n9518) );
  ANDN U10090 ( .A(n9526), .B(n5311), .Z(n9525) );
  XOR U10091 ( .A(n9527), .B(n9528), .Z(n5311) );
  IV U10092 ( .A(n9524), .Z(n9527) );
  XNOR U10093 ( .A(n5312), .B(n9524), .Z(n9526) );
  NAND U10094 ( .A(n9529), .B(e_input[462]), .Z(n5312) );
  NAND U10095 ( .A(n6112), .B(e_input[462]), .Z(n9529) );
  XOR U10096 ( .A(n9530), .B(n9531), .Z(n9524) );
  ANDN U10097 ( .A(n9532), .B(n5313), .Z(n9531) );
  XOR U10098 ( .A(n9533), .B(n9534), .Z(n5313) );
  IV U10099 ( .A(n9530), .Z(n9533) );
  XNOR U10100 ( .A(n5314), .B(n9530), .Z(n9532) );
  NAND U10101 ( .A(n9535), .B(e_input[461]), .Z(n5314) );
  NAND U10102 ( .A(n6112), .B(e_input[461]), .Z(n9535) );
  XOR U10103 ( .A(n9536), .B(n9537), .Z(n9530) );
  ANDN U10104 ( .A(n9538), .B(n5315), .Z(n9537) );
  XOR U10105 ( .A(n9539), .B(n9540), .Z(n5315) );
  IV U10106 ( .A(n9536), .Z(n9539) );
  XNOR U10107 ( .A(n5316), .B(n9536), .Z(n9538) );
  NAND U10108 ( .A(n9541), .B(e_input[460]), .Z(n5316) );
  NAND U10109 ( .A(n6112), .B(e_input[460]), .Z(n9541) );
  XOR U10110 ( .A(n9542), .B(n9543), .Z(n9536) );
  ANDN U10111 ( .A(n9544), .B(n5319), .Z(n9543) );
  XOR U10112 ( .A(n9545), .B(n9546), .Z(n5319) );
  IV U10113 ( .A(n9542), .Z(n9545) );
  XNOR U10114 ( .A(n5320), .B(n9542), .Z(n9544) );
  NAND U10115 ( .A(n9547), .B(e_input[459]), .Z(n5320) );
  NAND U10116 ( .A(n6112), .B(e_input[459]), .Z(n9547) );
  XOR U10117 ( .A(n9548), .B(n9549), .Z(n9542) );
  ANDN U10118 ( .A(n9550), .B(n5321), .Z(n9549) );
  XOR U10119 ( .A(n9551), .B(n9552), .Z(n5321) );
  IV U10120 ( .A(n9548), .Z(n9551) );
  XNOR U10121 ( .A(n5322), .B(n9548), .Z(n9550) );
  NAND U10122 ( .A(n9553), .B(e_input[458]), .Z(n5322) );
  NAND U10123 ( .A(n6112), .B(e_input[458]), .Z(n9553) );
  XOR U10124 ( .A(n9554), .B(n9555), .Z(n9548) );
  ANDN U10125 ( .A(n9556), .B(n5323), .Z(n9555) );
  XOR U10126 ( .A(n9557), .B(n9558), .Z(n5323) );
  IV U10127 ( .A(n9554), .Z(n9557) );
  XNOR U10128 ( .A(n5324), .B(n9554), .Z(n9556) );
  NAND U10129 ( .A(n9559), .B(e_input[457]), .Z(n5324) );
  NAND U10130 ( .A(n6112), .B(e_input[457]), .Z(n9559) );
  XOR U10131 ( .A(n9560), .B(n9561), .Z(n9554) );
  ANDN U10132 ( .A(n9562), .B(n5325), .Z(n9561) );
  XOR U10133 ( .A(n9563), .B(n9564), .Z(n5325) );
  IV U10134 ( .A(n9560), .Z(n9563) );
  XNOR U10135 ( .A(n5326), .B(n9560), .Z(n9562) );
  NAND U10136 ( .A(n9565), .B(e_input[456]), .Z(n5326) );
  NAND U10137 ( .A(n6112), .B(e_input[456]), .Z(n9565) );
  XOR U10138 ( .A(n9566), .B(n9567), .Z(n9560) );
  ANDN U10139 ( .A(n9568), .B(n5327), .Z(n9567) );
  XOR U10140 ( .A(n9569), .B(n9570), .Z(n5327) );
  IV U10141 ( .A(n9566), .Z(n9569) );
  XNOR U10142 ( .A(n5328), .B(n9566), .Z(n9568) );
  NAND U10143 ( .A(n9571), .B(e_input[455]), .Z(n5328) );
  NAND U10144 ( .A(n6112), .B(e_input[455]), .Z(n9571) );
  XOR U10145 ( .A(n9572), .B(n9573), .Z(n9566) );
  ANDN U10146 ( .A(n9574), .B(n5329), .Z(n9573) );
  XOR U10147 ( .A(n9575), .B(n9576), .Z(n5329) );
  IV U10148 ( .A(n9572), .Z(n9575) );
  XNOR U10149 ( .A(n5330), .B(n9572), .Z(n9574) );
  NAND U10150 ( .A(n9577), .B(e_input[454]), .Z(n5330) );
  NAND U10151 ( .A(n6112), .B(e_input[454]), .Z(n9577) );
  XOR U10152 ( .A(n9578), .B(n9579), .Z(n9572) );
  ANDN U10153 ( .A(n9580), .B(n5331), .Z(n9579) );
  XOR U10154 ( .A(n9581), .B(n9582), .Z(n5331) );
  IV U10155 ( .A(n9578), .Z(n9581) );
  XNOR U10156 ( .A(n5332), .B(n9578), .Z(n9580) );
  NAND U10157 ( .A(n9583), .B(e_input[453]), .Z(n5332) );
  NAND U10158 ( .A(n6112), .B(e_input[453]), .Z(n9583) );
  XOR U10159 ( .A(n9584), .B(n9585), .Z(n9578) );
  ANDN U10160 ( .A(n9586), .B(n5333), .Z(n9585) );
  XOR U10161 ( .A(n9587), .B(n9588), .Z(n5333) );
  IV U10162 ( .A(n9584), .Z(n9587) );
  XNOR U10163 ( .A(n5334), .B(n9584), .Z(n9586) );
  NAND U10164 ( .A(n9589), .B(e_input[452]), .Z(n5334) );
  NAND U10165 ( .A(n6112), .B(e_input[452]), .Z(n9589) );
  XOR U10166 ( .A(n9590), .B(n9591), .Z(n9584) );
  ANDN U10167 ( .A(n9592), .B(n5335), .Z(n9591) );
  XOR U10168 ( .A(n9593), .B(n9594), .Z(n5335) );
  IV U10169 ( .A(n9590), .Z(n9593) );
  XNOR U10170 ( .A(n5336), .B(n9590), .Z(n9592) );
  NAND U10171 ( .A(n9595), .B(e_input[451]), .Z(n5336) );
  NAND U10172 ( .A(n6112), .B(e_input[451]), .Z(n9595) );
  XOR U10173 ( .A(n9596), .B(n9597), .Z(n9590) );
  ANDN U10174 ( .A(n9598), .B(n5337), .Z(n9597) );
  XOR U10175 ( .A(n9599), .B(n9600), .Z(n5337) );
  IV U10176 ( .A(n9596), .Z(n9599) );
  XNOR U10177 ( .A(n5338), .B(n9596), .Z(n9598) );
  NAND U10178 ( .A(n9601), .B(e_input[450]), .Z(n5338) );
  NAND U10179 ( .A(n6112), .B(e_input[450]), .Z(n9601) );
  XOR U10180 ( .A(n9602), .B(n9603), .Z(n9596) );
  ANDN U10181 ( .A(n9604), .B(n5341), .Z(n9603) );
  XOR U10182 ( .A(n9605), .B(n9606), .Z(n5341) );
  IV U10183 ( .A(n9602), .Z(n9605) );
  XNOR U10184 ( .A(n5342), .B(n9602), .Z(n9604) );
  NAND U10185 ( .A(n9607), .B(e_input[449]), .Z(n5342) );
  NAND U10186 ( .A(n6112), .B(e_input[449]), .Z(n9607) );
  XOR U10187 ( .A(n9608), .B(n9609), .Z(n9602) );
  ANDN U10188 ( .A(n9610), .B(n5343), .Z(n9609) );
  XOR U10189 ( .A(n9611), .B(n9612), .Z(n5343) );
  IV U10190 ( .A(n9608), .Z(n9611) );
  XNOR U10191 ( .A(n5344), .B(n9608), .Z(n9610) );
  NAND U10192 ( .A(n9613), .B(e_input[448]), .Z(n5344) );
  NAND U10193 ( .A(n6112), .B(e_input[448]), .Z(n9613) );
  XOR U10194 ( .A(n9614), .B(n9615), .Z(n9608) );
  ANDN U10195 ( .A(n9616), .B(n5345), .Z(n9615) );
  XOR U10196 ( .A(n9617), .B(n9618), .Z(n5345) );
  IV U10197 ( .A(n9614), .Z(n9617) );
  XNOR U10198 ( .A(n5346), .B(n9614), .Z(n9616) );
  NAND U10199 ( .A(n9619), .B(e_input[447]), .Z(n5346) );
  NAND U10200 ( .A(n6112), .B(e_input[447]), .Z(n9619) );
  XOR U10201 ( .A(n9620), .B(n9621), .Z(n9614) );
  ANDN U10202 ( .A(n9622), .B(n5347), .Z(n9621) );
  XOR U10203 ( .A(n9623), .B(n9624), .Z(n5347) );
  IV U10204 ( .A(n9620), .Z(n9623) );
  XNOR U10205 ( .A(n5348), .B(n9620), .Z(n9622) );
  NAND U10206 ( .A(n9625), .B(e_input[446]), .Z(n5348) );
  NAND U10207 ( .A(n6112), .B(e_input[446]), .Z(n9625) );
  XOR U10208 ( .A(n9626), .B(n9627), .Z(n9620) );
  ANDN U10209 ( .A(n9628), .B(n5349), .Z(n9627) );
  XOR U10210 ( .A(n9629), .B(n9630), .Z(n5349) );
  IV U10211 ( .A(n9626), .Z(n9629) );
  XNOR U10212 ( .A(n5350), .B(n9626), .Z(n9628) );
  NAND U10213 ( .A(n9631), .B(e_input[445]), .Z(n5350) );
  NAND U10214 ( .A(n6112), .B(e_input[445]), .Z(n9631) );
  XOR U10215 ( .A(n9632), .B(n9633), .Z(n9626) );
  ANDN U10216 ( .A(n9634), .B(n5351), .Z(n9633) );
  XOR U10217 ( .A(n9635), .B(n9636), .Z(n5351) );
  IV U10218 ( .A(n9632), .Z(n9635) );
  XNOR U10219 ( .A(n5352), .B(n9632), .Z(n9634) );
  NAND U10220 ( .A(n9637), .B(e_input[444]), .Z(n5352) );
  NAND U10221 ( .A(n6112), .B(e_input[444]), .Z(n9637) );
  XOR U10222 ( .A(n9638), .B(n9639), .Z(n9632) );
  ANDN U10223 ( .A(n9640), .B(n5353), .Z(n9639) );
  XOR U10224 ( .A(n9641), .B(n9642), .Z(n5353) );
  IV U10225 ( .A(n9638), .Z(n9641) );
  XNOR U10226 ( .A(n5354), .B(n9638), .Z(n9640) );
  NAND U10227 ( .A(n9643), .B(e_input[443]), .Z(n5354) );
  NAND U10228 ( .A(n6112), .B(e_input[443]), .Z(n9643) );
  XOR U10229 ( .A(n9644), .B(n9645), .Z(n9638) );
  ANDN U10230 ( .A(n9646), .B(n5355), .Z(n9645) );
  XOR U10231 ( .A(n9647), .B(n9648), .Z(n5355) );
  IV U10232 ( .A(n9644), .Z(n9647) );
  XNOR U10233 ( .A(n5356), .B(n9644), .Z(n9646) );
  NAND U10234 ( .A(n9649), .B(e_input[442]), .Z(n5356) );
  NAND U10235 ( .A(n6112), .B(e_input[442]), .Z(n9649) );
  XOR U10236 ( .A(n9650), .B(n9651), .Z(n9644) );
  ANDN U10237 ( .A(n9652), .B(n5357), .Z(n9651) );
  XOR U10238 ( .A(n9653), .B(n9654), .Z(n5357) );
  IV U10239 ( .A(n9650), .Z(n9653) );
  XNOR U10240 ( .A(n5358), .B(n9650), .Z(n9652) );
  NAND U10241 ( .A(n9655), .B(e_input[441]), .Z(n5358) );
  NAND U10242 ( .A(n6112), .B(e_input[441]), .Z(n9655) );
  XOR U10243 ( .A(n9656), .B(n9657), .Z(n9650) );
  ANDN U10244 ( .A(n9658), .B(n5359), .Z(n9657) );
  XOR U10245 ( .A(n9659), .B(n9660), .Z(n5359) );
  IV U10246 ( .A(n9656), .Z(n9659) );
  XNOR U10247 ( .A(n5360), .B(n9656), .Z(n9658) );
  NAND U10248 ( .A(n9661), .B(e_input[440]), .Z(n5360) );
  NAND U10249 ( .A(n6112), .B(e_input[440]), .Z(n9661) );
  XOR U10250 ( .A(n9662), .B(n9663), .Z(n9656) );
  ANDN U10251 ( .A(n9664), .B(n5363), .Z(n9663) );
  XOR U10252 ( .A(n9665), .B(n9666), .Z(n5363) );
  IV U10253 ( .A(n9662), .Z(n9665) );
  XNOR U10254 ( .A(n5364), .B(n9662), .Z(n9664) );
  NAND U10255 ( .A(n9667), .B(e_input[439]), .Z(n5364) );
  NAND U10256 ( .A(n6112), .B(e_input[439]), .Z(n9667) );
  XOR U10257 ( .A(n9668), .B(n9669), .Z(n9662) );
  ANDN U10258 ( .A(n9670), .B(n5365), .Z(n9669) );
  XOR U10259 ( .A(n9671), .B(n9672), .Z(n5365) );
  IV U10260 ( .A(n9668), .Z(n9671) );
  XNOR U10261 ( .A(n5366), .B(n9668), .Z(n9670) );
  NAND U10262 ( .A(n9673), .B(e_input[438]), .Z(n5366) );
  NAND U10263 ( .A(n6112), .B(e_input[438]), .Z(n9673) );
  XOR U10264 ( .A(n9674), .B(n9675), .Z(n9668) );
  ANDN U10265 ( .A(n9676), .B(n5367), .Z(n9675) );
  XOR U10266 ( .A(n9677), .B(n9678), .Z(n5367) );
  IV U10267 ( .A(n9674), .Z(n9677) );
  XNOR U10268 ( .A(n5368), .B(n9674), .Z(n9676) );
  NAND U10269 ( .A(n9679), .B(e_input[437]), .Z(n5368) );
  NAND U10270 ( .A(n6112), .B(e_input[437]), .Z(n9679) );
  XOR U10271 ( .A(n9680), .B(n9681), .Z(n9674) );
  ANDN U10272 ( .A(n9682), .B(n5369), .Z(n9681) );
  XOR U10273 ( .A(n9683), .B(n9684), .Z(n5369) );
  IV U10274 ( .A(n9680), .Z(n9683) );
  XNOR U10275 ( .A(n5370), .B(n9680), .Z(n9682) );
  NAND U10276 ( .A(n9685), .B(e_input[436]), .Z(n5370) );
  NAND U10277 ( .A(n6112), .B(e_input[436]), .Z(n9685) );
  XOR U10278 ( .A(n9686), .B(n9687), .Z(n9680) );
  ANDN U10279 ( .A(n9688), .B(n5371), .Z(n9687) );
  XOR U10280 ( .A(n9689), .B(n9690), .Z(n5371) );
  IV U10281 ( .A(n9686), .Z(n9689) );
  XNOR U10282 ( .A(n5372), .B(n9686), .Z(n9688) );
  NAND U10283 ( .A(n9691), .B(e_input[435]), .Z(n5372) );
  NAND U10284 ( .A(n6112), .B(e_input[435]), .Z(n9691) );
  XOR U10285 ( .A(n9692), .B(n9693), .Z(n9686) );
  ANDN U10286 ( .A(n9694), .B(n5373), .Z(n9693) );
  XOR U10287 ( .A(n9695), .B(n9696), .Z(n5373) );
  IV U10288 ( .A(n9692), .Z(n9695) );
  XNOR U10289 ( .A(n5374), .B(n9692), .Z(n9694) );
  NAND U10290 ( .A(n9697), .B(e_input[434]), .Z(n5374) );
  NAND U10291 ( .A(n6112), .B(e_input[434]), .Z(n9697) );
  XOR U10292 ( .A(n9698), .B(n9699), .Z(n9692) );
  ANDN U10293 ( .A(n9700), .B(n5375), .Z(n9699) );
  XOR U10294 ( .A(n9701), .B(n9702), .Z(n5375) );
  IV U10295 ( .A(n9698), .Z(n9701) );
  XNOR U10296 ( .A(n5376), .B(n9698), .Z(n9700) );
  NAND U10297 ( .A(n9703), .B(e_input[433]), .Z(n5376) );
  NAND U10298 ( .A(n6112), .B(e_input[433]), .Z(n9703) );
  XOR U10299 ( .A(n9704), .B(n9705), .Z(n9698) );
  ANDN U10300 ( .A(n9706), .B(n5377), .Z(n9705) );
  XOR U10301 ( .A(n9707), .B(n9708), .Z(n5377) );
  IV U10302 ( .A(n9704), .Z(n9707) );
  XNOR U10303 ( .A(n5378), .B(n9704), .Z(n9706) );
  NAND U10304 ( .A(n9709), .B(e_input[432]), .Z(n5378) );
  NAND U10305 ( .A(n6112), .B(e_input[432]), .Z(n9709) );
  XOR U10306 ( .A(n9710), .B(n9711), .Z(n9704) );
  ANDN U10307 ( .A(n9712), .B(n5379), .Z(n9711) );
  XOR U10308 ( .A(n9713), .B(n9714), .Z(n5379) );
  IV U10309 ( .A(n9710), .Z(n9713) );
  XNOR U10310 ( .A(n5380), .B(n9710), .Z(n9712) );
  NAND U10311 ( .A(n9715), .B(e_input[431]), .Z(n5380) );
  NAND U10312 ( .A(n6112), .B(e_input[431]), .Z(n9715) );
  XOR U10313 ( .A(n9716), .B(n9717), .Z(n9710) );
  ANDN U10314 ( .A(n9718), .B(n5381), .Z(n9717) );
  XOR U10315 ( .A(n9719), .B(n9720), .Z(n5381) );
  IV U10316 ( .A(n9716), .Z(n9719) );
  XNOR U10317 ( .A(n5382), .B(n9716), .Z(n9718) );
  NAND U10318 ( .A(n9721), .B(e_input[430]), .Z(n5382) );
  NAND U10319 ( .A(n6112), .B(e_input[430]), .Z(n9721) );
  XOR U10320 ( .A(n9722), .B(n9723), .Z(n9716) );
  ANDN U10321 ( .A(n9724), .B(n5385), .Z(n9723) );
  XOR U10322 ( .A(n9725), .B(n9726), .Z(n5385) );
  IV U10323 ( .A(n9722), .Z(n9725) );
  XNOR U10324 ( .A(n5386), .B(n9722), .Z(n9724) );
  NAND U10325 ( .A(n9727), .B(e_input[429]), .Z(n5386) );
  NAND U10326 ( .A(n6112), .B(e_input[429]), .Z(n9727) );
  XOR U10327 ( .A(n9728), .B(n9729), .Z(n9722) );
  ANDN U10328 ( .A(n9730), .B(n5387), .Z(n9729) );
  XOR U10329 ( .A(n9731), .B(n9732), .Z(n5387) );
  IV U10330 ( .A(n9728), .Z(n9731) );
  XNOR U10331 ( .A(n5388), .B(n9728), .Z(n9730) );
  NAND U10332 ( .A(n9733), .B(e_input[428]), .Z(n5388) );
  NAND U10333 ( .A(n6112), .B(e_input[428]), .Z(n9733) );
  XOR U10334 ( .A(n9734), .B(n9735), .Z(n9728) );
  ANDN U10335 ( .A(n9736), .B(n5389), .Z(n9735) );
  XOR U10336 ( .A(n9737), .B(n9738), .Z(n5389) );
  IV U10337 ( .A(n9734), .Z(n9737) );
  XNOR U10338 ( .A(n5390), .B(n9734), .Z(n9736) );
  NAND U10339 ( .A(n9739), .B(e_input[427]), .Z(n5390) );
  NAND U10340 ( .A(n6112), .B(e_input[427]), .Z(n9739) );
  XOR U10341 ( .A(n9740), .B(n9741), .Z(n9734) );
  ANDN U10342 ( .A(n9742), .B(n5391), .Z(n9741) );
  XOR U10343 ( .A(n9743), .B(n9744), .Z(n5391) );
  IV U10344 ( .A(n9740), .Z(n9743) );
  XNOR U10345 ( .A(n5392), .B(n9740), .Z(n9742) );
  NAND U10346 ( .A(n9745), .B(e_input[426]), .Z(n5392) );
  NAND U10347 ( .A(n6112), .B(e_input[426]), .Z(n9745) );
  XOR U10348 ( .A(n9746), .B(n9747), .Z(n9740) );
  ANDN U10349 ( .A(n9748), .B(n5393), .Z(n9747) );
  XOR U10350 ( .A(n9749), .B(n9750), .Z(n5393) );
  IV U10351 ( .A(n9746), .Z(n9749) );
  XNOR U10352 ( .A(n5394), .B(n9746), .Z(n9748) );
  NAND U10353 ( .A(n9751), .B(e_input[425]), .Z(n5394) );
  NAND U10354 ( .A(n6112), .B(e_input[425]), .Z(n9751) );
  XOR U10355 ( .A(n9752), .B(n9753), .Z(n9746) );
  ANDN U10356 ( .A(n9754), .B(n5395), .Z(n9753) );
  XOR U10357 ( .A(n9755), .B(n9756), .Z(n5395) );
  IV U10358 ( .A(n9752), .Z(n9755) );
  XNOR U10359 ( .A(n5396), .B(n9752), .Z(n9754) );
  NAND U10360 ( .A(n9757), .B(e_input[424]), .Z(n5396) );
  NAND U10361 ( .A(n6112), .B(e_input[424]), .Z(n9757) );
  XOR U10362 ( .A(n9758), .B(n9759), .Z(n9752) );
  ANDN U10363 ( .A(n9760), .B(n5397), .Z(n9759) );
  XOR U10364 ( .A(n9761), .B(n9762), .Z(n5397) );
  IV U10365 ( .A(n9758), .Z(n9761) );
  XNOR U10366 ( .A(n5398), .B(n9758), .Z(n9760) );
  NAND U10367 ( .A(n9763), .B(e_input[423]), .Z(n5398) );
  NAND U10368 ( .A(n6112), .B(e_input[423]), .Z(n9763) );
  XOR U10369 ( .A(n9764), .B(n9765), .Z(n9758) );
  ANDN U10370 ( .A(n9766), .B(n5399), .Z(n9765) );
  XOR U10371 ( .A(n9767), .B(n9768), .Z(n5399) );
  IV U10372 ( .A(n9764), .Z(n9767) );
  XNOR U10373 ( .A(n5400), .B(n9764), .Z(n9766) );
  NAND U10374 ( .A(n9769), .B(e_input[422]), .Z(n5400) );
  NAND U10375 ( .A(n6112), .B(e_input[422]), .Z(n9769) );
  XOR U10376 ( .A(n9770), .B(n9771), .Z(n9764) );
  ANDN U10377 ( .A(n9772), .B(n5401), .Z(n9771) );
  XOR U10378 ( .A(n9773), .B(n9774), .Z(n5401) );
  IV U10379 ( .A(n9770), .Z(n9773) );
  XNOR U10380 ( .A(n5402), .B(n9770), .Z(n9772) );
  NAND U10381 ( .A(n9775), .B(e_input[421]), .Z(n5402) );
  NAND U10382 ( .A(n6112), .B(e_input[421]), .Z(n9775) );
  XOR U10383 ( .A(n9776), .B(n9777), .Z(n9770) );
  ANDN U10384 ( .A(n9778), .B(n5403), .Z(n9777) );
  XOR U10385 ( .A(n9779), .B(n9780), .Z(n5403) );
  IV U10386 ( .A(n9776), .Z(n9779) );
  XNOR U10387 ( .A(n5404), .B(n9776), .Z(n9778) );
  NAND U10388 ( .A(n9781), .B(e_input[420]), .Z(n5404) );
  NAND U10389 ( .A(n6112), .B(e_input[420]), .Z(n9781) );
  XOR U10390 ( .A(n9782), .B(n9783), .Z(n9776) );
  ANDN U10391 ( .A(n9784), .B(n5407), .Z(n9783) );
  XOR U10392 ( .A(n9785), .B(n9786), .Z(n5407) );
  IV U10393 ( .A(n9782), .Z(n9785) );
  XNOR U10394 ( .A(n5408), .B(n9782), .Z(n9784) );
  NAND U10395 ( .A(n9787), .B(e_input[419]), .Z(n5408) );
  NAND U10396 ( .A(n6112), .B(e_input[419]), .Z(n9787) );
  XOR U10397 ( .A(n9788), .B(n9789), .Z(n9782) );
  ANDN U10398 ( .A(n9790), .B(n5409), .Z(n9789) );
  XOR U10399 ( .A(n9791), .B(n9792), .Z(n5409) );
  IV U10400 ( .A(n9788), .Z(n9791) );
  XNOR U10401 ( .A(n5410), .B(n9788), .Z(n9790) );
  NAND U10402 ( .A(n9793), .B(e_input[418]), .Z(n5410) );
  NAND U10403 ( .A(n6112), .B(e_input[418]), .Z(n9793) );
  XOR U10404 ( .A(n9794), .B(n9795), .Z(n9788) );
  ANDN U10405 ( .A(n9796), .B(n5411), .Z(n9795) );
  XOR U10406 ( .A(n9797), .B(n9798), .Z(n5411) );
  IV U10407 ( .A(n9794), .Z(n9797) );
  XNOR U10408 ( .A(n5412), .B(n9794), .Z(n9796) );
  NAND U10409 ( .A(n9799), .B(e_input[417]), .Z(n5412) );
  NAND U10410 ( .A(n6112), .B(e_input[417]), .Z(n9799) );
  XOR U10411 ( .A(n9800), .B(n9801), .Z(n9794) );
  ANDN U10412 ( .A(n9802), .B(n5413), .Z(n9801) );
  XOR U10413 ( .A(n9803), .B(n9804), .Z(n5413) );
  IV U10414 ( .A(n9800), .Z(n9803) );
  XNOR U10415 ( .A(n5414), .B(n9800), .Z(n9802) );
  NAND U10416 ( .A(n9805), .B(e_input[416]), .Z(n5414) );
  NAND U10417 ( .A(n6112), .B(e_input[416]), .Z(n9805) );
  XOR U10418 ( .A(n9806), .B(n9807), .Z(n9800) );
  ANDN U10419 ( .A(n9808), .B(n5415), .Z(n9807) );
  XOR U10420 ( .A(n9809), .B(n9810), .Z(n5415) );
  IV U10421 ( .A(n9806), .Z(n9809) );
  XNOR U10422 ( .A(n5416), .B(n9806), .Z(n9808) );
  NAND U10423 ( .A(n9811), .B(e_input[415]), .Z(n5416) );
  NAND U10424 ( .A(n6112), .B(e_input[415]), .Z(n9811) );
  XOR U10425 ( .A(n9812), .B(n9813), .Z(n9806) );
  ANDN U10426 ( .A(n9814), .B(n5417), .Z(n9813) );
  XOR U10427 ( .A(n9815), .B(n9816), .Z(n5417) );
  IV U10428 ( .A(n9812), .Z(n9815) );
  XNOR U10429 ( .A(n5418), .B(n9812), .Z(n9814) );
  NAND U10430 ( .A(n9817), .B(e_input[414]), .Z(n5418) );
  NAND U10431 ( .A(n6112), .B(e_input[414]), .Z(n9817) );
  XOR U10432 ( .A(n9818), .B(n9819), .Z(n9812) );
  ANDN U10433 ( .A(n9820), .B(n5419), .Z(n9819) );
  XOR U10434 ( .A(n9821), .B(n9822), .Z(n5419) );
  IV U10435 ( .A(n9818), .Z(n9821) );
  XNOR U10436 ( .A(n5420), .B(n9818), .Z(n9820) );
  NAND U10437 ( .A(n9823), .B(e_input[413]), .Z(n5420) );
  NAND U10438 ( .A(n6112), .B(e_input[413]), .Z(n9823) );
  XOR U10439 ( .A(n9824), .B(n9825), .Z(n9818) );
  ANDN U10440 ( .A(n9826), .B(n5421), .Z(n9825) );
  XOR U10441 ( .A(n9827), .B(n9828), .Z(n5421) );
  IV U10442 ( .A(n9824), .Z(n9827) );
  XNOR U10443 ( .A(n5422), .B(n9824), .Z(n9826) );
  NAND U10444 ( .A(n9829), .B(e_input[412]), .Z(n5422) );
  NAND U10445 ( .A(n6112), .B(e_input[412]), .Z(n9829) );
  XOR U10446 ( .A(n9830), .B(n9831), .Z(n9824) );
  ANDN U10447 ( .A(n9832), .B(n5423), .Z(n9831) );
  XOR U10448 ( .A(n9833), .B(n9834), .Z(n5423) );
  IV U10449 ( .A(n9830), .Z(n9833) );
  XNOR U10450 ( .A(n5424), .B(n9830), .Z(n9832) );
  NAND U10451 ( .A(n9835), .B(e_input[411]), .Z(n5424) );
  NAND U10452 ( .A(n6112), .B(e_input[411]), .Z(n9835) );
  XOR U10453 ( .A(n9836), .B(n9837), .Z(n9830) );
  ANDN U10454 ( .A(n9838), .B(n5425), .Z(n9837) );
  XOR U10455 ( .A(n9839), .B(n9840), .Z(n5425) );
  IV U10456 ( .A(n9836), .Z(n9839) );
  XNOR U10457 ( .A(n5426), .B(n9836), .Z(n9838) );
  NAND U10458 ( .A(n9841), .B(e_input[410]), .Z(n5426) );
  NAND U10459 ( .A(n6112), .B(e_input[410]), .Z(n9841) );
  XOR U10460 ( .A(n9842), .B(n9843), .Z(n9836) );
  ANDN U10461 ( .A(n9844), .B(n5429), .Z(n9843) );
  XOR U10462 ( .A(n9845), .B(n9846), .Z(n5429) );
  IV U10463 ( .A(n9842), .Z(n9845) );
  XNOR U10464 ( .A(n5430), .B(n9842), .Z(n9844) );
  NAND U10465 ( .A(n9847), .B(e_input[409]), .Z(n5430) );
  NAND U10466 ( .A(n6112), .B(e_input[409]), .Z(n9847) );
  XOR U10467 ( .A(n9848), .B(n9849), .Z(n9842) );
  ANDN U10468 ( .A(n9850), .B(n5431), .Z(n9849) );
  XOR U10469 ( .A(n9851), .B(n9852), .Z(n5431) );
  IV U10470 ( .A(n9848), .Z(n9851) );
  XNOR U10471 ( .A(n5432), .B(n9848), .Z(n9850) );
  NAND U10472 ( .A(n9853), .B(e_input[408]), .Z(n5432) );
  NAND U10473 ( .A(n6112), .B(e_input[408]), .Z(n9853) );
  XOR U10474 ( .A(n9854), .B(n9855), .Z(n9848) );
  ANDN U10475 ( .A(n9856), .B(n5433), .Z(n9855) );
  XOR U10476 ( .A(n9857), .B(n9858), .Z(n5433) );
  IV U10477 ( .A(n9854), .Z(n9857) );
  XNOR U10478 ( .A(n5434), .B(n9854), .Z(n9856) );
  NAND U10479 ( .A(n9859), .B(e_input[407]), .Z(n5434) );
  NAND U10480 ( .A(n6112), .B(e_input[407]), .Z(n9859) );
  XOR U10481 ( .A(n9860), .B(n9861), .Z(n9854) );
  ANDN U10482 ( .A(n9862), .B(n5435), .Z(n9861) );
  XOR U10483 ( .A(n9863), .B(n9864), .Z(n5435) );
  IV U10484 ( .A(n9860), .Z(n9863) );
  XNOR U10485 ( .A(n5436), .B(n9860), .Z(n9862) );
  NAND U10486 ( .A(n9865), .B(e_input[406]), .Z(n5436) );
  NAND U10487 ( .A(n6112), .B(e_input[406]), .Z(n9865) );
  XOR U10488 ( .A(n9866), .B(n9867), .Z(n9860) );
  ANDN U10489 ( .A(n9868), .B(n5437), .Z(n9867) );
  XOR U10490 ( .A(n9869), .B(n9870), .Z(n5437) );
  IV U10491 ( .A(n9866), .Z(n9869) );
  XNOR U10492 ( .A(n5438), .B(n9866), .Z(n9868) );
  NAND U10493 ( .A(n9871), .B(e_input[405]), .Z(n5438) );
  NAND U10494 ( .A(n6112), .B(e_input[405]), .Z(n9871) );
  XOR U10495 ( .A(n9872), .B(n9873), .Z(n9866) );
  ANDN U10496 ( .A(n9874), .B(n5439), .Z(n9873) );
  XOR U10497 ( .A(n9875), .B(n9876), .Z(n5439) );
  IV U10498 ( .A(n9872), .Z(n9875) );
  XNOR U10499 ( .A(n5440), .B(n9872), .Z(n9874) );
  NAND U10500 ( .A(n9877), .B(e_input[404]), .Z(n5440) );
  NAND U10501 ( .A(n6112), .B(e_input[404]), .Z(n9877) );
  XOR U10502 ( .A(n9878), .B(n9879), .Z(n9872) );
  ANDN U10503 ( .A(n9880), .B(n5441), .Z(n9879) );
  XOR U10504 ( .A(n9881), .B(n9882), .Z(n5441) );
  IV U10505 ( .A(n9878), .Z(n9881) );
  XNOR U10506 ( .A(n5442), .B(n9878), .Z(n9880) );
  NAND U10507 ( .A(n9883), .B(e_input[403]), .Z(n5442) );
  NAND U10508 ( .A(n6112), .B(e_input[403]), .Z(n9883) );
  XOR U10509 ( .A(n9884), .B(n9885), .Z(n9878) );
  ANDN U10510 ( .A(n9886), .B(n5443), .Z(n9885) );
  XOR U10511 ( .A(n9887), .B(n9888), .Z(n5443) );
  IV U10512 ( .A(n9884), .Z(n9887) );
  XNOR U10513 ( .A(n5444), .B(n9884), .Z(n9886) );
  NAND U10514 ( .A(n9889), .B(e_input[402]), .Z(n5444) );
  NAND U10515 ( .A(n6112), .B(e_input[402]), .Z(n9889) );
  XOR U10516 ( .A(n9890), .B(n9891), .Z(n9884) );
  ANDN U10517 ( .A(n9892), .B(n5445), .Z(n9891) );
  XOR U10518 ( .A(n9893), .B(n9894), .Z(n5445) );
  IV U10519 ( .A(n9890), .Z(n9893) );
  XNOR U10520 ( .A(n5446), .B(n9890), .Z(n9892) );
  NAND U10521 ( .A(n9895), .B(e_input[401]), .Z(n5446) );
  NAND U10522 ( .A(n6112), .B(e_input[401]), .Z(n9895) );
  XOR U10523 ( .A(n9896), .B(n9897), .Z(n9890) );
  ANDN U10524 ( .A(n9898), .B(n5447), .Z(n9897) );
  XOR U10525 ( .A(n9899), .B(n9900), .Z(n5447) );
  IV U10526 ( .A(n9896), .Z(n9899) );
  XNOR U10527 ( .A(n5448), .B(n9896), .Z(n9898) );
  NAND U10528 ( .A(n9901), .B(e_input[400]), .Z(n5448) );
  NAND U10529 ( .A(n6112), .B(e_input[400]), .Z(n9901) );
  XOR U10530 ( .A(n9902), .B(n9903), .Z(n9896) );
  ANDN U10531 ( .A(n9904), .B(n5453), .Z(n9903) );
  XOR U10532 ( .A(n9905), .B(n9906), .Z(n5453) );
  IV U10533 ( .A(n9902), .Z(n9905) );
  XNOR U10534 ( .A(n5454), .B(n9902), .Z(n9904) );
  NAND U10535 ( .A(n9907), .B(e_input[399]), .Z(n5454) );
  NAND U10536 ( .A(n6112), .B(e_input[399]), .Z(n9907) );
  XOR U10537 ( .A(n9908), .B(n9909), .Z(n9902) );
  ANDN U10538 ( .A(n9910), .B(n5455), .Z(n9909) );
  XOR U10539 ( .A(n9911), .B(n9912), .Z(n5455) );
  IV U10540 ( .A(n9908), .Z(n9911) );
  XNOR U10541 ( .A(n5456), .B(n9908), .Z(n9910) );
  NAND U10542 ( .A(n9913), .B(e_input[398]), .Z(n5456) );
  NAND U10543 ( .A(n6112), .B(e_input[398]), .Z(n9913) );
  XOR U10544 ( .A(n9914), .B(n9915), .Z(n9908) );
  ANDN U10545 ( .A(n9916), .B(n5457), .Z(n9915) );
  XOR U10546 ( .A(n9917), .B(n9918), .Z(n5457) );
  IV U10547 ( .A(n9914), .Z(n9917) );
  XNOR U10548 ( .A(n5458), .B(n9914), .Z(n9916) );
  NAND U10549 ( .A(n9919), .B(e_input[397]), .Z(n5458) );
  NAND U10550 ( .A(n6112), .B(e_input[397]), .Z(n9919) );
  XOR U10551 ( .A(n9920), .B(n9921), .Z(n9914) );
  ANDN U10552 ( .A(n9922), .B(n5459), .Z(n9921) );
  XOR U10553 ( .A(n9923), .B(n9924), .Z(n5459) );
  IV U10554 ( .A(n9920), .Z(n9923) );
  XNOR U10555 ( .A(n5460), .B(n9920), .Z(n9922) );
  NAND U10556 ( .A(n9925), .B(e_input[396]), .Z(n5460) );
  NAND U10557 ( .A(n6112), .B(e_input[396]), .Z(n9925) );
  XOR U10558 ( .A(n9926), .B(n9927), .Z(n9920) );
  ANDN U10559 ( .A(n9928), .B(n5461), .Z(n9927) );
  XOR U10560 ( .A(n9929), .B(n9930), .Z(n5461) );
  IV U10561 ( .A(n9926), .Z(n9929) );
  XNOR U10562 ( .A(n5462), .B(n9926), .Z(n9928) );
  NAND U10563 ( .A(n9931), .B(e_input[395]), .Z(n5462) );
  NAND U10564 ( .A(n6112), .B(e_input[395]), .Z(n9931) );
  XOR U10565 ( .A(n9932), .B(n9933), .Z(n9926) );
  ANDN U10566 ( .A(n9934), .B(n5463), .Z(n9933) );
  XOR U10567 ( .A(n9935), .B(n9936), .Z(n5463) );
  IV U10568 ( .A(n9932), .Z(n9935) );
  XNOR U10569 ( .A(n5464), .B(n9932), .Z(n9934) );
  NAND U10570 ( .A(n9937), .B(e_input[394]), .Z(n5464) );
  NAND U10571 ( .A(n6112), .B(e_input[394]), .Z(n9937) );
  XOR U10572 ( .A(n9938), .B(n9939), .Z(n9932) );
  ANDN U10573 ( .A(n9940), .B(n5465), .Z(n9939) );
  XOR U10574 ( .A(n9941), .B(n9942), .Z(n5465) );
  IV U10575 ( .A(n9938), .Z(n9941) );
  XNOR U10576 ( .A(n5466), .B(n9938), .Z(n9940) );
  NAND U10577 ( .A(n9943), .B(e_input[393]), .Z(n5466) );
  NAND U10578 ( .A(n6112), .B(e_input[393]), .Z(n9943) );
  XOR U10579 ( .A(n9944), .B(n9945), .Z(n9938) );
  ANDN U10580 ( .A(n9946), .B(n5467), .Z(n9945) );
  XOR U10581 ( .A(n9947), .B(n9948), .Z(n5467) );
  IV U10582 ( .A(n9944), .Z(n9947) );
  XNOR U10583 ( .A(n5468), .B(n9944), .Z(n9946) );
  NAND U10584 ( .A(n9949), .B(e_input[392]), .Z(n5468) );
  NAND U10585 ( .A(n6112), .B(e_input[392]), .Z(n9949) );
  XOR U10586 ( .A(n9950), .B(n9951), .Z(n9944) );
  ANDN U10587 ( .A(n9952), .B(n5469), .Z(n9951) );
  XOR U10588 ( .A(n9953), .B(n9954), .Z(n5469) );
  IV U10589 ( .A(n9950), .Z(n9953) );
  XNOR U10590 ( .A(n5470), .B(n9950), .Z(n9952) );
  NAND U10591 ( .A(n9955), .B(e_input[391]), .Z(n5470) );
  NAND U10592 ( .A(n6112), .B(e_input[391]), .Z(n9955) );
  XOR U10593 ( .A(n9956), .B(n9957), .Z(n9950) );
  ANDN U10594 ( .A(n9958), .B(n5471), .Z(n9957) );
  XOR U10595 ( .A(n9959), .B(n9960), .Z(n5471) );
  IV U10596 ( .A(n9956), .Z(n9959) );
  XNOR U10597 ( .A(n5472), .B(n9956), .Z(n9958) );
  NAND U10598 ( .A(n9961), .B(e_input[390]), .Z(n5472) );
  NAND U10599 ( .A(n6112), .B(e_input[390]), .Z(n9961) );
  XOR U10600 ( .A(n9962), .B(n9963), .Z(n9956) );
  ANDN U10601 ( .A(n9964), .B(n5475), .Z(n9963) );
  XOR U10602 ( .A(n9965), .B(n9966), .Z(n5475) );
  IV U10603 ( .A(n9962), .Z(n9965) );
  XNOR U10604 ( .A(n5476), .B(n9962), .Z(n9964) );
  NAND U10605 ( .A(n9967), .B(e_input[389]), .Z(n5476) );
  NAND U10606 ( .A(n6112), .B(e_input[389]), .Z(n9967) );
  XOR U10607 ( .A(n9968), .B(n9969), .Z(n9962) );
  ANDN U10608 ( .A(n9970), .B(n5477), .Z(n9969) );
  XOR U10609 ( .A(n9971), .B(n9972), .Z(n5477) );
  IV U10610 ( .A(n9968), .Z(n9971) );
  XNOR U10611 ( .A(n5478), .B(n9968), .Z(n9970) );
  NAND U10612 ( .A(n9973), .B(e_input[388]), .Z(n5478) );
  NAND U10613 ( .A(n6112), .B(e_input[388]), .Z(n9973) );
  XOR U10614 ( .A(n9974), .B(n9975), .Z(n9968) );
  ANDN U10615 ( .A(n9976), .B(n5479), .Z(n9975) );
  XOR U10616 ( .A(n9977), .B(n9978), .Z(n5479) );
  IV U10617 ( .A(n9974), .Z(n9977) );
  XNOR U10618 ( .A(n5480), .B(n9974), .Z(n9976) );
  NAND U10619 ( .A(n9979), .B(e_input[387]), .Z(n5480) );
  NAND U10620 ( .A(n6112), .B(e_input[387]), .Z(n9979) );
  XOR U10621 ( .A(n9980), .B(n9981), .Z(n9974) );
  ANDN U10622 ( .A(n9982), .B(n5481), .Z(n9981) );
  XOR U10623 ( .A(n9983), .B(n9984), .Z(n5481) );
  IV U10624 ( .A(n9980), .Z(n9983) );
  XNOR U10625 ( .A(n5482), .B(n9980), .Z(n9982) );
  NAND U10626 ( .A(n9985), .B(e_input[386]), .Z(n5482) );
  NAND U10627 ( .A(n6112), .B(e_input[386]), .Z(n9985) );
  XOR U10628 ( .A(n9986), .B(n9987), .Z(n9980) );
  ANDN U10629 ( .A(n9988), .B(n5483), .Z(n9987) );
  XOR U10630 ( .A(n9989), .B(n9990), .Z(n5483) );
  IV U10631 ( .A(n9986), .Z(n9989) );
  XNOR U10632 ( .A(n5484), .B(n9986), .Z(n9988) );
  NAND U10633 ( .A(n9991), .B(e_input[385]), .Z(n5484) );
  NAND U10634 ( .A(n6112), .B(e_input[385]), .Z(n9991) );
  XOR U10635 ( .A(n9992), .B(n9993), .Z(n9986) );
  ANDN U10636 ( .A(n9994), .B(n5485), .Z(n9993) );
  XOR U10637 ( .A(n9995), .B(n9996), .Z(n5485) );
  IV U10638 ( .A(n9992), .Z(n9995) );
  XNOR U10639 ( .A(n5486), .B(n9992), .Z(n9994) );
  NAND U10640 ( .A(n9997), .B(e_input[384]), .Z(n5486) );
  NAND U10641 ( .A(n6112), .B(e_input[384]), .Z(n9997) );
  XOR U10642 ( .A(n9998), .B(n9999), .Z(n9992) );
  ANDN U10643 ( .A(n10000), .B(n5487), .Z(n9999) );
  XOR U10644 ( .A(n10001), .B(n10002), .Z(n5487) );
  IV U10645 ( .A(n9998), .Z(n10001) );
  XNOR U10646 ( .A(n5488), .B(n9998), .Z(n10000) );
  NAND U10647 ( .A(n10003), .B(e_input[383]), .Z(n5488) );
  NAND U10648 ( .A(n6112), .B(e_input[383]), .Z(n10003) );
  XOR U10649 ( .A(n10004), .B(n10005), .Z(n9998) );
  ANDN U10650 ( .A(n10006), .B(n5489), .Z(n10005) );
  XOR U10651 ( .A(n10007), .B(n10008), .Z(n5489) );
  IV U10652 ( .A(n10004), .Z(n10007) );
  XNOR U10653 ( .A(n5490), .B(n10004), .Z(n10006) );
  NAND U10654 ( .A(n10009), .B(e_input[382]), .Z(n5490) );
  NAND U10655 ( .A(n6112), .B(e_input[382]), .Z(n10009) );
  XOR U10656 ( .A(n10010), .B(n10011), .Z(n10004) );
  ANDN U10657 ( .A(n10012), .B(n5491), .Z(n10011) );
  XOR U10658 ( .A(n10013), .B(n10014), .Z(n5491) );
  IV U10659 ( .A(n10010), .Z(n10013) );
  XNOR U10660 ( .A(n5492), .B(n10010), .Z(n10012) );
  NAND U10661 ( .A(n10015), .B(e_input[381]), .Z(n5492) );
  NAND U10662 ( .A(n6112), .B(e_input[381]), .Z(n10015) );
  XOR U10663 ( .A(n10016), .B(n10017), .Z(n10010) );
  ANDN U10664 ( .A(n10018), .B(n5493), .Z(n10017) );
  XOR U10665 ( .A(n10019), .B(n10020), .Z(n5493) );
  IV U10666 ( .A(n10016), .Z(n10019) );
  XNOR U10667 ( .A(n5494), .B(n10016), .Z(n10018) );
  NAND U10668 ( .A(n10021), .B(e_input[380]), .Z(n5494) );
  NAND U10669 ( .A(n6112), .B(e_input[380]), .Z(n10021) );
  XOR U10670 ( .A(n10022), .B(n10023), .Z(n10016) );
  ANDN U10671 ( .A(n10024), .B(n5497), .Z(n10023) );
  XOR U10672 ( .A(n10025), .B(n10026), .Z(n5497) );
  IV U10673 ( .A(n10022), .Z(n10025) );
  XNOR U10674 ( .A(n5498), .B(n10022), .Z(n10024) );
  NAND U10675 ( .A(n10027), .B(e_input[379]), .Z(n5498) );
  NAND U10676 ( .A(n6112), .B(e_input[379]), .Z(n10027) );
  XOR U10677 ( .A(n10028), .B(n10029), .Z(n10022) );
  ANDN U10678 ( .A(n10030), .B(n5499), .Z(n10029) );
  XOR U10679 ( .A(n10031), .B(n10032), .Z(n5499) );
  IV U10680 ( .A(n10028), .Z(n10031) );
  XNOR U10681 ( .A(n5500), .B(n10028), .Z(n10030) );
  NAND U10682 ( .A(n10033), .B(e_input[378]), .Z(n5500) );
  NAND U10683 ( .A(n6112), .B(e_input[378]), .Z(n10033) );
  XOR U10684 ( .A(n10034), .B(n10035), .Z(n10028) );
  ANDN U10685 ( .A(n10036), .B(n5501), .Z(n10035) );
  XOR U10686 ( .A(n10037), .B(n10038), .Z(n5501) );
  IV U10687 ( .A(n10034), .Z(n10037) );
  XNOR U10688 ( .A(n5502), .B(n10034), .Z(n10036) );
  NAND U10689 ( .A(n10039), .B(e_input[377]), .Z(n5502) );
  NAND U10690 ( .A(n6112), .B(e_input[377]), .Z(n10039) );
  XOR U10691 ( .A(n10040), .B(n10041), .Z(n10034) );
  ANDN U10692 ( .A(n10042), .B(n5503), .Z(n10041) );
  XOR U10693 ( .A(n10043), .B(n10044), .Z(n5503) );
  IV U10694 ( .A(n10040), .Z(n10043) );
  XNOR U10695 ( .A(n5504), .B(n10040), .Z(n10042) );
  NAND U10696 ( .A(n10045), .B(e_input[376]), .Z(n5504) );
  NAND U10697 ( .A(n6112), .B(e_input[376]), .Z(n10045) );
  XOR U10698 ( .A(n10046), .B(n10047), .Z(n10040) );
  ANDN U10699 ( .A(n10048), .B(n5505), .Z(n10047) );
  XOR U10700 ( .A(n10049), .B(n10050), .Z(n5505) );
  IV U10701 ( .A(n10046), .Z(n10049) );
  XNOR U10702 ( .A(n5506), .B(n10046), .Z(n10048) );
  NAND U10703 ( .A(n10051), .B(e_input[375]), .Z(n5506) );
  NAND U10704 ( .A(n6112), .B(e_input[375]), .Z(n10051) );
  XOR U10705 ( .A(n10052), .B(n10053), .Z(n10046) );
  ANDN U10706 ( .A(n10054), .B(n5507), .Z(n10053) );
  XOR U10707 ( .A(n10055), .B(n10056), .Z(n5507) );
  IV U10708 ( .A(n10052), .Z(n10055) );
  XNOR U10709 ( .A(n5508), .B(n10052), .Z(n10054) );
  NAND U10710 ( .A(n10057), .B(e_input[374]), .Z(n5508) );
  NAND U10711 ( .A(n6112), .B(e_input[374]), .Z(n10057) );
  XOR U10712 ( .A(n10058), .B(n10059), .Z(n10052) );
  ANDN U10713 ( .A(n10060), .B(n5509), .Z(n10059) );
  XOR U10714 ( .A(n10061), .B(n10062), .Z(n5509) );
  IV U10715 ( .A(n10058), .Z(n10061) );
  XNOR U10716 ( .A(n5510), .B(n10058), .Z(n10060) );
  NAND U10717 ( .A(n10063), .B(e_input[373]), .Z(n5510) );
  NAND U10718 ( .A(n6112), .B(e_input[373]), .Z(n10063) );
  XOR U10719 ( .A(n10064), .B(n10065), .Z(n10058) );
  ANDN U10720 ( .A(n10066), .B(n5511), .Z(n10065) );
  XOR U10721 ( .A(n10067), .B(n10068), .Z(n5511) );
  IV U10722 ( .A(n10064), .Z(n10067) );
  XNOR U10723 ( .A(n5512), .B(n10064), .Z(n10066) );
  NAND U10724 ( .A(n10069), .B(e_input[372]), .Z(n5512) );
  NAND U10725 ( .A(n6112), .B(e_input[372]), .Z(n10069) );
  XOR U10726 ( .A(n10070), .B(n10071), .Z(n10064) );
  ANDN U10727 ( .A(n10072), .B(n5513), .Z(n10071) );
  XOR U10728 ( .A(n10073), .B(n10074), .Z(n5513) );
  IV U10729 ( .A(n10070), .Z(n10073) );
  XNOR U10730 ( .A(n5514), .B(n10070), .Z(n10072) );
  NAND U10731 ( .A(n10075), .B(e_input[371]), .Z(n5514) );
  NAND U10732 ( .A(n6112), .B(e_input[371]), .Z(n10075) );
  XOR U10733 ( .A(n10076), .B(n10077), .Z(n10070) );
  ANDN U10734 ( .A(n10078), .B(n5515), .Z(n10077) );
  XOR U10735 ( .A(n10079), .B(n10080), .Z(n5515) );
  IV U10736 ( .A(n10076), .Z(n10079) );
  XNOR U10737 ( .A(n5516), .B(n10076), .Z(n10078) );
  NAND U10738 ( .A(n10081), .B(e_input[370]), .Z(n5516) );
  NAND U10739 ( .A(n6112), .B(e_input[370]), .Z(n10081) );
  XOR U10740 ( .A(n10082), .B(n10083), .Z(n10076) );
  ANDN U10741 ( .A(n10084), .B(n5519), .Z(n10083) );
  XOR U10742 ( .A(n10085), .B(n10086), .Z(n5519) );
  IV U10743 ( .A(n10082), .Z(n10085) );
  XNOR U10744 ( .A(n5520), .B(n10082), .Z(n10084) );
  NAND U10745 ( .A(n10087), .B(e_input[369]), .Z(n5520) );
  NAND U10746 ( .A(n6112), .B(e_input[369]), .Z(n10087) );
  XOR U10747 ( .A(n10088), .B(n10089), .Z(n10082) );
  ANDN U10748 ( .A(n10090), .B(n5521), .Z(n10089) );
  XOR U10749 ( .A(n10091), .B(n10092), .Z(n5521) );
  IV U10750 ( .A(n10088), .Z(n10091) );
  XNOR U10751 ( .A(n5522), .B(n10088), .Z(n10090) );
  NAND U10752 ( .A(n10093), .B(e_input[368]), .Z(n5522) );
  NAND U10753 ( .A(n6112), .B(e_input[368]), .Z(n10093) );
  XOR U10754 ( .A(n10094), .B(n10095), .Z(n10088) );
  ANDN U10755 ( .A(n10096), .B(n5523), .Z(n10095) );
  XOR U10756 ( .A(n10097), .B(n10098), .Z(n5523) );
  IV U10757 ( .A(n10094), .Z(n10097) );
  XNOR U10758 ( .A(n5524), .B(n10094), .Z(n10096) );
  NAND U10759 ( .A(n10099), .B(e_input[367]), .Z(n5524) );
  NAND U10760 ( .A(n6112), .B(e_input[367]), .Z(n10099) );
  XOR U10761 ( .A(n10100), .B(n10101), .Z(n10094) );
  ANDN U10762 ( .A(n10102), .B(n5525), .Z(n10101) );
  XOR U10763 ( .A(n10103), .B(n10104), .Z(n5525) );
  IV U10764 ( .A(n10100), .Z(n10103) );
  XNOR U10765 ( .A(n5526), .B(n10100), .Z(n10102) );
  NAND U10766 ( .A(n10105), .B(e_input[366]), .Z(n5526) );
  NAND U10767 ( .A(n6112), .B(e_input[366]), .Z(n10105) );
  XOR U10768 ( .A(n10106), .B(n10107), .Z(n10100) );
  ANDN U10769 ( .A(n10108), .B(n5527), .Z(n10107) );
  XOR U10770 ( .A(n10109), .B(n10110), .Z(n5527) );
  IV U10771 ( .A(n10106), .Z(n10109) );
  XNOR U10772 ( .A(n5528), .B(n10106), .Z(n10108) );
  NAND U10773 ( .A(n10111), .B(e_input[365]), .Z(n5528) );
  NAND U10774 ( .A(n6112), .B(e_input[365]), .Z(n10111) );
  XOR U10775 ( .A(n10112), .B(n10113), .Z(n10106) );
  ANDN U10776 ( .A(n10114), .B(n5529), .Z(n10113) );
  XOR U10777 ( .A(n10115), .B(n10116), .Z(n5529) );
  IV U10778 ( .A(n10112), .Z(n10115) );
  XNOR U10779 ( .A(n5530), .B(n10112), .Z(n10114) );
  NAND U10780 ( .A(n10117), .B(e_input[364]), .Z(n5530) );
  NAND U10781 ( .A(n6112), .B(e_input[364]), .Z(n10117) );
  XOR U10782 ( .A(n10118), .B(n10119), .Z(n10112) );
  ANDN U10783 ( .A(n10120), .B(n5531), .Z(n10119) );
  XOR U10784 ( .A(n10121), .B(n10122), .Z(n5531) );
  IV U10785 ( .A(n10118), .Z(n10121) );
  XNOR U10786 ( .A(n5532), .B(n10118), .Z(n10120) );
  NAND U10787 ( .A(n10123), .B(e_input[363]), .Z(n5532) );
  NAND U10788 ( .A(n6112), .B(e_input[363]), .Z(n10123) );
  XOR U10789 ( .A(n10124), .B(n10125), .Z(n10118) );
  ANDN U10790 ( .A(n10126), .B(n5533), .Z(n10125) );
  XOR U10791 ( .A(n10127), .B(n10128), .Z(n5533) );
  IV U10792 ( .A(n10124), .Z(n10127) );
  XNOR U10793 ( .A(n5534), .B(n10124), .Z(n10126) );
  NAND U10794 ( .A(n10129), .B(e_input[362]), .Z(n5534) );
  NAND U10795 ( .A(n6112), .B(e_input[362]), .Z(n10129) );
  XOR U10796 ( .A(n10130), .B(n10131), .Z(n10124) );
  ANDN U10797 ( .A(n10132), .B(n5535), .Z(n10131) );
  XOR U10798 ( .A(n10133), .B(n10134), .Z(n5535) );
  IV U10799 ( .A(n10130), .Z(n10133) );
  XNOR U10800 ( .A(n5536), .B(n10130), .Z(n10132) );
  NAND U10801 ( .A(n10135), .B(e_input[361]), .Z(n5536) );
  NAND U10802 ( .A(n6112), .B(e_input[361]), .Z(n10135) );
  XOR U10803 ( .A(n10136), .B(n10137), .Z(n10130) );
  ANDN U10804 ( .A(n10138), .B(n5537), .Z(n10137) );
  XOR U10805 ( .A(n10139), .B(n10140), .Z(n5537) );
  IV U10806 ( .A(n10136), .Z(n10139) );
  XNOR U10807 ( .A(n5538), .B(n10136), .Z(n10138) );
  NAND U10808 ( .A(n10141), .B(e_input[360]), .Z(n5538) );
  NAND U10809 ( .A(n6112), .B(e_input[360]), .Z(n10141) );
  XOR U10810 ( .A(n10142), .B(n10143), .Z(n10136) );
  ANDN U10811 ( .A(n10144), .B(n5541), .Z(n10143) );
  XOR U10812 ( .A(n10145), .B(n10146), .Z(n5541) );
  IV U10813 ( .A(n10142), .Z(n10145) );
  XNOR U10814 ( .A(n5542), .B(n10142), .Z(n10144) );
  NAND U10815 ( .A(n10147), .B(e_input[359]), .Z(n5542) );
  NAND U10816 ( .A(n6112), .B(e_input[359]), .Z(n10147) );
  XOR U10817 ( .A(n10148), .B(n10149), .Z(n10142) );
  ANDN U10818 ( .A(n10150), .B(n5543), .Z(n10149) );
  XOR U10819 ( .A(n10151), .B(n10152), .Z(n5543) );
  IV U10820 ( .A(n10148), .Z(n10151) );
  XNOR U10821 ( .A(n5544), .B(n10148), .Z(n10150) );
  NAND U10822 ( .A(n10153), .B(e_input[358]), .Z(n5544) );
  NAND U10823 ( .A(n6112), .B(e_input[358]), .Z(n10153) );
  XOR U10824 ( .A(n10154), .B(n10155), .Z(n10148) );
  ANDN U10825 ( .A(n10156), .B(n5545), .Z(n10155) );
  XOR U10826 ( .A(n10157), .B(n10158), .Z(n5545) );
  IV U10827 ( .A(n10154), .Z(n10157) );
  XNOR U10828 ( .A(n5546), .B(n10154), .Z(n10156) );
  NAND U10829 ( .A(n10159), .B(e_input[357]), .Z(n5546) );
  NAND U10830 ( .A(n6112), .B(e_input[357]), .Z(n10159) );
  XOR U10831 ( .A(n10160), .B(n10161), .Z(n10154) );
  ANDN U10832 ( .A(n10162), .B(n5547), .Z(n10161) );
  XOR U10833 ( .A(n10163), .B(n10164), .Z(n5547) );
  IV U10834 ( .A(n10160), .Z(n10163) );
  XNOR U10835 ( .A(n5548), .B(n10160), .Z(n10162) );
  NAND U10836 ( .A(n10165), .B(e_input[356]), .Z(n5548) );
  NAND U10837 ( .A(n6112), .B(e_input[356]), .Z(n10165) );
  XOR U10838 ( .A(n10166), .B(n10167), .Z(n10160) );
  ANDN U10839 ( .A(n10168), .B(n5549), .Z(n10167) );
  XOR U10840 ( .A(n10169), .B(n10170), .Z(n5549) );
  IV U10841 ( .A(n10166), .Z(n10169) );
  XNOR U10842 ( .A(n5550), .B(n10166), .Z(n10168) );
  NAND U10843 ( .A(n10171), .B(e_input[355]), .Z(n5550) );
  NAND U10844 ( .A(n6112), .B(e_input[355]), .Z(n10171) );
  XOR U10845 ( .A(n10172), .B(n10173), .Z(n10166) );
  ANDN U10846 ( .A(n10174), .B(n5551), .Z(n10173) );
  XOR U10847 ( .A(n10175), .B(n10176), .Z(n5551) );
  IV U10848 ( .A(n10172), .Z(n10175) );
  XNOR U10849 ( .A(n5552), .B(n10172), .Z(n10174) );
  NAND U10850 ( .A(n10177), .B(e_input[354]), .Z(n5552) );
  NAND U10851 ( .A(n6112), .B(e_input[354]), .Z(n10177) );
  XOR U10852 ( .A(n10178), .B(n10179), .Z(n10172) );
  ANDN U10853 ( .A(n10180), .B(n5553), .Z(n10179) );
  XOR U10854 ( .A(n10181), .B(n10182), .Z(n5553) );
  IV U10855 ( .A(n10178), .Z(n10181) );
  XNOR U10856 ( .A(n5554), .B(n10178), .Z(n10180) );
  NAND U10857 ( .A(n10183), .B(e_input[353]), .Z(n5554) );
  NAND U10858 ( .A(n6112), .B(e_input[353]), .Z(n10183) );
  XOR U10859 ( .A(n10184), .B(n10185), .Z(n10178) );
  ANDN U10860 ( .A(n10186), .B(n5555), .Z(n10185) );
  XOR U10861 ( .A(n10187), .B(n10188), .Z(n5555) );
  IV U10862 ( .A(n10184), .Z(n10187) );
  XNOR U10863 ( .A(n5556), .B(n10184), .Z(n10186) );
  NAND U10864 ( .A(n10189), .B(e_input[352]), .Z(n5556) );
  NAND U10865 ( .A(n6112), .B(e_input[352]), .Z(n10189) );
  XOR U10866 ( .A(n10190), .B(n10191), .Z(n10184) );
  ANDN U10867 ( .A(n10192), .B(n5557), .Z(n10191) );
  XOR U10868 ( .A(n10193), .B(n10194), .Z(n5557) );
  IV U10869 ( .A(n10190), .Z(n10193) );
  XNOR U10870 ( .A(n5558), .B(n10190), .Z(n10192) );
  NAND U10871 ( .A(n10195), .B(e_input[351]), .Z(n5558) );
  NAND U10872 ( .A(n6112), .B(e_input[351]), .Z(n10195) );
  XOR U10873 ( .A(n10196), .B(n10197), .Z(n10190) );
  ANDN U10874 ( .A(n10198), .B(n5559), .Z(n10197) );
  XOR U10875 ( .A(n10199), .B(n10200), .Z(n5559) );
  IV U10876 ( .A(n10196), .Z(n10199) );
  XNOR U10877 ( .A(n5560), .B(n10196), .Z(n10198) );
  NAND U10878 ( .A(n10201), .B(e_input[350]), .Z(n5560) );
  NAND U10879 ( .A(n6112), .B(e_input[350]), .Z(n10201) );
  XOR U10880 ( .A(n10202), .B(n10203), .Z(n10196) );
  ANDN U10881 ( .A(n10204), .B(n5563), .Z(n10203) );
  XOR U10882 ( .A(n10205), .B(n10206), .Z(n5563) );
  IV U10883 ( .A(n10202), .Z(n10205) );
  XNOR U10884 ( .A(n5564), .B(n10202), .Z(n10204) );
  NAND U10885 ( .A(n10207), .B(e_input[349]), .Z(n5564) );
  NAND U10886 ( .A(n6112), .B(e_input[349]), .Z(n10207) );
  XOR U10887 ( .A(n10208), .B(n10209), .Z(n10202) );
  ANDN U10888 ( .A(n10210), .B(n5565), .Z(n10209) );
  XOR U10889 ( .A(n10211), .B(n10212), .Z(n5565) );
  IV U10890 ( .A(n10208), .Z(n10211) );
  XNOR U10891 ( .A(n5566), .B(n10208), .Z(n10210) );
  NAND U10892 ( .A(n10213), .B(e_input[348]), .Z(n5566) );
  NAND U10893 ( .A(n6112), .B(e_input[348]), .Z(n10213) );
  XOR U10894 ( .A(n10214), .B(n10215), .Z(n10208) );
  ANDN U10895 ( .A(n10216), .B(n5567), .Z(n10215) );
  XOR U10896 ( .A(n10217), .B(n10218), .Z(n5567) );
  IV U10897 ( .A(n10214), .Z(n10217) );
  XNOR U10898 ( .A(n5568), .B(n10214), .Z(n10216) );
  NAND U10899 ( .A(n10219), .B(e_input[347]), .Z(n5568) );
  NAND U10900 ( .A(n6112), .B(e_input[347]), .Z(n10219) );
  XOR U10901 ( .A(n10220), .B(n10221), .Z(n10214) );
  ANDN U10902 ( .A(n10222), .B(n5569), .Z(n10221) );
  XOR U10903 ( .A(n10223), .B(n10224), .Z(n5569) );
  IV U10904 ( .A(n10220), .Z(n10223) );
  XNOR U10905 ( .A(n5570), .B(n10220), .Z(n10222) );
  NAND U10906 ( .A(n10225), .B(e_input[346]), .Z(n5570) );
  NAND U10907 ( .A(n6112), .B(e_input[346]), .Z(n10225) );
  XOR U10908 ( .A(n10226), .B(n10227), .Z(n10220) );
  ANDN U10909 ( .A(n10228), .B(n5571), .Z(n10227) );
  XOR U10910 ( .A(n10229), .B(n10230), .Z(n5571) );
  IV U10911 ( .A(n10226), .Z(n10229) );
  XNOR U10912 ( .A(n5572), .B(n10226), .Z(n10228) );
  NAND U10913 ( .A(n10231), .B(e_input[345]), .Z(n5572) );
  NAND U10914 ( .A(n6112), .B(e_input[345]), .Z(n10231) );
  XOR U10915 ( .A(n10232), .B(n10233), .Z(n10226) );
  ANDN U10916 ( .A(n10234), .B(n5573), .Z(n10233) );
  XOR U10917 ( .A(n10235), .B(n10236), .Z(n5573) );
  IV U10918 ( .A(n10232), .Z(n10235) );
  XNOR U10919 ( .A(n5574), .B(n10232), .Z(n10234) );
  NAND U10920 ( .A(n10237), .B(e_input[344]), .Z(n5574) );
  NAND U10921 ( .A(n6112), .B(e_input[344]), .Z(n10237) );
  XOR U10922 ( .A(n10238), .B(n10239), .Z(n10232) );
  ANDN U10923 ( .A(n10240), .B(n5575), .Z(n10239) );
  XOR U10924 ( .A(n10241), .B(n10242), .Z(n5575) );
  IV U10925 ( .A(n10238), .Z(n10241) );
  XNOR U10926 ( .A(n5576), .B(n10238), .Z(n10240) );
  NAND U10927 ( .A(n10243), .B(e_input[343]), .Z(n5576) );
  NAND U10928 ( .A(n6112), .B(e_input[343]), .Z(n10243) );
  XOR U10929 ( .A(n10244), .B(n10245), .Z(n10238) );
  ANDN U10930 ( .A(n10246), .B(n5577), .Z(n10245) );
  XOR U10931 ( .A(n10247), .B(n10248), .Z(n5577) );
  IV U10932 ( .A(n10244), .Z(n10247) );
  XNOR U10933 ( .A(n5578), .B(n10244), .Z(n10246) );
  NAND U10934 ( .A(n10249), .B(e_input[342]), .Z(n5578) );
  NAND U10935 ( .A(n6112), .B(e_input[342]), .Z(n10249) );
  XOR U10936 ( .A(n10250), .B(n10251), .Z(n10244) );
  ANDN U10937 ( .A(n10252), .B(n5579), .Z(n10251) );
  XOR U10938 ( .A(n10253), .B(n10254), .Z(n5579) );
  IV U10939 ( .A(n10250), .Z(n10253) );
  XNOR U10940 ( .A(n5580), .B(n10250), .Z(n10252) );
  NAND U10941 ( .A(n10255), .B(e_input[341]), .Z(n5580) );
  NAND U10942 ( .A(n6112), .B(e_input[341]), .Z(n10255) );
  XOR U10943 ( .A(n10256), .B(n10257), .Z(n10250) );
  ANDN U10944 ( .A(n10258), .B(n5581), .Z(n10257) );
  XOR U10945 ( .A(n10259), .B(n10260), .Z(n5581) );
  IV U10946 ( .A(n10256), .Z(n10259) );
  XNOR U10947 ( .A(n5582), .B(n10256), .Z(n10258) );
  NAND U10948 ( .A(n10261), .B(e_input[340]), .Z(n5582) );
  NAND U10949 ( .A(n6112), .B(e_input[340]), .Z(n10261) );
  XOR U10950 ( .A(n10262), .B(n10263), .Z(n10256) );
  ANDN U10951 ( .A(n10264), .B(n5585), .Z(n10263) );
  XOR U10952 ( .A(n10265), .B(n10266), .Z(n5585) );
  IV U10953 ( .A(n10262), .Z(n10265) );
  XNOR U10954 ( .A(n5586), .B(n10262), .Z(n10264) );
  NAND U10955 ( .A(n10267), .B(e_input[339]), .Z(n5586) );
  NAND U10956 ( .A(n6112), .B(e_input[339]), .Z(n10267) );
  XOR U10957 ( .A(n10268), .B(n10269), .Z(n10262) );
  ANDN U10958 ( .A(n10270), .B(n5587), .Z(n10269) );
  XOR U10959 ( .A(n10271), .B(n10272), .Z(n5587) );
  IV U10960 ( .A(n10268), .Z(n10271) );
  XNOR U10961 ( .A(n5588), .B(n10268), .Z(n10270) );
  NAND U10962 ( .A(n10273), .B(e_input[338]), .Z(n5588) );
  NAND U10963 ( .A(n6112), .B(e_input[338]), .Z(n10273) );
  XOR U10964 ( .A(n10274), .B(n10275), .Z(n10268) );
  ANDN U10965 ( .A(n10276), .B(n5589), .Z(n10275) );
  XOR U10966 ( .A(n10277), .B(n10278), .Z(n5589) );
  IV U10967 ( .A(n10274), .Z(n10277) );
  XNOR U10968 ( .A(n5590), .B(n10274), .Z(n10276) );
  NAND U10969 ( .A(n10279), .B(e_input[337]), .Z(n5590) );
  NAND U10970 ( .A(n6112), .B(e_input[337]), .Z(n10279) );
  XOR U10971 ( .A(n10280), .B(n10281), .Z(n10274) );
  ANDN U10972 ( .A(n10282), .B(n5591), .Z(n10281) );
  XOR U10973 ( .A(n10283), .B(n10284), .Z(n5591) );
  IV U10974 ( .A(n10280), .Z(n10283) );
  XNOR U10975 ( .A(n5592), .B(n10280), .Z(n10282) );
  NAND U10976 ( .A(n10285), .B(e_input[336]), .Z(n5592) );
  NAND U10977 ( .A(n6112), .B(e_input[336]), .Z(n10285) );
  XOR U10978 ( .A(n10286), .B(n10287), .Z(n10280) );
  ANDN U10979 ( .A(n10288), .B(n5593), .Z(n10287) );
  XOR U10980 ( .A(n10289), .B(n10290), .Z(n5593) );
  IV U10981 ( .A(n10286), .Z(n10289) );
  XNOR U10982 ( .A(n5594), .B(n10286), .Z(n10288) );
  NAND U10983 ( .A(n10291), .B(e_input[335]), .Z(n5594) );
  NAND U10984 ( .A(n6112), .B(e_input[335]), .Z(n10291) );
  XOR U10985 ( .A(n10292), .B(n10293), .Z(n10286) );
  ANDN U10986 ( .A(n10294), .B(n5595), .Z(n10293) );
  XOR U10987 ( .A(n10295), .B(n10296), .Z(n5595) );
  IV U10988 ( .A(n10292), .Z(n10295) );
  XNOR U10989 ( .A(n5596), .B(n10292), .Z(n10294) );
  NAND U10990 ( .A(n10297), .B(e_input[334]), .Z(n5596) );
  NAND U10991 ( .A(n6112), .B(e_input[334]), .Z(n10297) );
  XOR U10992 ( .A(n10298), .B(n10299), .Z(n10292) );
  ANDN U10993 ( .A(n10300), .B(n5597), .Z(n10299) );
  XOR U10994 ( .A(n10301), .B(n10302), .Z(n5597) );
  IV U10995 ( .A(n10298), .Z(n10301) );
  XNOR U10996 ( .A(n5598), .B(n10298), .Z(n10300) );
  NAND U10997 ( .A(n10303), .B(e_input[333]), .Z(n5598) );
  NAND U10998 ( .A(n6112), .B(e_input[333]), .Z(n10303) );
  XOR U10999 ( .A(n10304), .B(n10305), .Z(n10298) );
  ANDN U11000 ( .A(n10306), .B(n5599), .Z(n10305) );
  XOR U11001 ( .A(n10307), .B(n10308), .Z(n5599) );
  IV U11002 ( .A(n10304), .Z(n10307) );
  XNOR U11003 ( .A(n5600), .B(n10304), .Z(n10306) );
  NAND U11004 ( .A(n10309), .B(e_input[332]), .Z(n5600) );
  NAND U11005 ( .A(n6112), .B(e_input[332]), .Z(n10309) );
  XOR U11006 ( .A(n10310), .B(n10311), .Z(n10304) );
  ANDN U11007 ( .A(n10312), .B(n5601), .Z(n10311) );
  XOR U11008 ( .A(n10313), .B(n10314), .Z(n5601) );
  IV U11009 ( .A(n10310), .Z(n10313) );
  XNOR U11010 ( .A(n5602), .B(n10310), .Z(n10312) );
  NAND U11011 ( .A(n10315), .B(e_input[331]), .Z(n5602) );
  NAND U11012 ( .A(n6112), .B(e_input[331]), .Z(n10315) );
  XOR U11013 ( .A(n10316), .B(n10317), .Z(n10310) );
  ANDN U11014 ( .A(n10318), .B(n5603), .Z(n10317) );
  XOR U11015 ( .A(n10319), .B(n10320), .Z(n5603) );
  IV U11016 ( .A(n10316), .Z(n10319) );
  XNOR U11017 ( .A(n5604), .B(n10316), .Z(n10318) );
  NAND U11018 ( .A(n10321), .B(e_input[330]), .Z(n5604) );
  NAND U11019 ( .A(n6112), .B(e_input[330]), .Z(n10321) );
  XOR U11020 ( .A(n10322), .B(n10323), .Z(n10316) );
  ANDN U11021 ( .A(n10324), .B(n5607), .Z(n10323) );
  XOR U11022 ( .A(n10325), .B(n10326), .Z(n5607) );
  IV U11023 ( .A(n10322), .Z(n10325) );
  XNOR U11024 ( .A(n5608), .B(n10322), .Z(n10324) );
  NAND U11025 ( .A(n10327), .B(e_input[329]), .Z(n5608) );
  NAND U11026 ( .A(n6112), .B(e_input[329]), .Z(n10327) );
  XOR U11027 ( .A(n10328), .B(n10329), .Z(n10322) );
  ANDN U11028 ( .A(n10330), .B(n5609), .Z(n10329) );
  XOR U11029 ( .A(n10331), .B(n10332), .Z(n5609) );
  IV U11030 ( .A(n10328), .Z(n10331) );
  XNOR U11031 ( .A(n5610), .B(n10328), .Z(n10330) );
  NAND U11032 ( .A(n10333), .B(e_input[328]), .Z(n5610) );
  NAND U11033 ( .A(n6112), .B(e_input[328]), .Z(n10333) );
  XOR U11034 ( .A(n10334), .B(n10335), .Z(n10328) );
  ANDN U11035 ( .A(n10336), .B(n5611), .Z(n10335) );
  XOR U11036 ( .A(n10337), .B(n10338), .Z(n5611) );
  IV U11037 ( .A(n10334), .Z(n10337) );
  XNOR U11038 ( .A(n5612), .B(n10334), .Z(n10336) );
  NAND U11039 ( .A(n10339), .B(e_input[327]), .Z(n5612) );
  NAND U11040 ( .A(n6112), .B(e_input[327]), .Z(n10339) );
  XOR U11041 ( .A(n10340), .B(n10341), .Z(n10334) );
  ANDN U11042 ( .A(n10342), .B(n5613), .Z(n10341) );
  XOR U11043 ( .A(n10343), .B(n10344), .Z(n5613) );
  IV U11044 ( .A(n10340), .Z(n10343) );
  XNOR U11045 ( .A(n5614), .B(n10340), .Z(n10342) );
  NAND U11046 ( .A(n10345), .B(e_input[326]), .Z(n5614) );
  NAND U11047 ( .A(n6112), .B(e_input[326]), .Z(n10345) );
  XOR U11048 ( .A(n10346), .B(n10347), .Z(n10340) );
  ANDN U11049 ( .A(n10348), .B(n5615), .Z(n10347) );
  XOR U11050 ( .A(n10349), .B(n10350), .Z(n5615) );
  IV U11051 ( .A(n10346), .Z(n10349) );
  XNOR U11052 ( .A(n5616), .B(n10346), .Z(n10348) );
  NAND U11053 ( .A(n10351), .B(e_input[325]), .Z(n5616) );
  NAND U11054 ( .A(n6112), .B(e_input[325]), .Z(n10351) );
  XOR U11055 ( .A(n10352), .B(n10353), .Z(n10346) );
  ANDN U11056 ( .A(n10354), .B(n5617), .Z(n10353) );
  XOR U11057 ( .A(n10355), .B(n10356), .Z(n5617) );
  IV U11058 ( .A(n10352), .Z(n10355) );
  XNOR U11059 ( .A(n5618), .B(n10352), .Z(n10354) );
  NAND U11060 ( .A(n10357), .B(e_input[324]), .Z(n5618) );
  NAND U11061 ( .A(n6112), .B(e_input[324]), .Z(n10357) );
  XOR U11062 ( .A(n10358), .B(n10359), .Z(n10352) );
  ANDN U11063 ( .A(n10360), .B(n5619), .Z(n10359) );
  XOR U11064 ( .A(n10361), .B(n10362), .Z(n5619) );
  IV U11065 ( .A(n10358), .Z(n10361) );
  XNOR U11066 ( .A(n5620), .B(n10358), .Z(n10360) );
  NAND U11067 ( .A(n10363), .B(e_input[323]), .Z(n5620) );
  NAND U11068 ( .A(n6112), .B(e_input[323]), .Z(n10363) );
  XOR U11069 ( .A(n10364), .B(n10365), .Z(n10358) );
  ANDN U11070 ( .A(n10366), .B(n5621), .Z(n10365) );
  XOR U11071 ( .A(n10367), .B(n10368), .Z(n5621) );
  IV U11072 ( .A(n10364), .Z(n10367) );
  XNOR U11073 ( .A(n5622), .B(n10364), .Z(n10366) );
  NAND U11074 ( .A(n10369), .B(e_input[322]), .Z(n5622) );
  NAND U11075 ( .A(n6112), .B(e_input[322]), .Z(n10369) );
  XOR U11076 ( .A(n10370), .B(n10371), .Z(n10364) );
  ANDN U11077 ( .A(n10372), .B(n5623), .Z(n10371) );
  XOR U11078 ( .A(n10373), .B(n10374), .Z(n5623) );
  IV U11079 ( .A(n10370), .Z(n10373) );
  XNOR U11080 ( .A(n5624), .B(n10370), .Z(n10372) );
  NAND U11081 ( .A(n10375), .B(e_input[321]), .Z(n5624) );
  NAND U11082 ( .A(n6112), .B(e_input[321]), .Z(n10375) );
  XOR U11083 ( .A(n10376), .B(n10377), .Z(n10370) );
  ANDN U11084 ( .A(n10378), .B(n5625), .Z(n10377) );
  XOR U11085 ( .A(n10379), .B(n10380), .Z(n5625) );
  IV U11086 ( .A(n10376), .Z(n10379) );
  XNOR U11087 ( .A(n5626), .B(n10376), .Z(n10378) );
  NAND U11088 ( .A(n10381), .B(e_input[320]), .Z(n5626) );
  NAND U11089 ( .A(n6112), .B(e_input[320]), .Z(n10381) );
  XOR U11090 ( .A(n10382), .B(n10383), .Z(n10376) );
  ANDN U11091 ( .A(n10384), .B(n5629), .Z(n10383) );
  XOR U11092 ( .A(n10385), .B(n10386), .Z(n5629) );
  IV U11093 ( .A(n10382), .Z(n10385) );
  XNOR U11094 ( .A(n5630), .B(n10382), .Z(n10384) );
  NAND U11095 ( .A(n10387), .B(e_input[319]), .Z(n5630) );
  NAND U11096 ( .A(n6112), .B(e_input[319]), .Z(n10387) );
  XOR U11097 ( .A(n10388), .B(n10389), .Z(n10382) );
  ANDN U11098 ( .A(n10390), .B(n5631), .Z(n10389) );
  XOR U11099 ( .A(n10391), .B(n10392), .Z(n5631) );
  IV U11100 ( .A(n10388), .Z(n10391) );
  XNOR U11101 ( .A(n5632), .B(n10388), .Z(n10390) );
  NAND U11102 ( .A(n10393), .B(e_input[318]), .Z(n5632) );
  NAND U11103 ( .A(n6112), .B(e_input[318]), .Z(n10393) );
  XOR U11104 ( .A(n10394), .B(n10395), .Z(n10388) );
  ANDN U11105 ( .A(n10396), .B(n5633), .Z(n10395) );
  XOR U11106 ( .A(n10397), .B(n10398), .Z(n5633) );
  IV U11107 ( .A(n10394), .Z(n10397) );
  XNOR U11108 ( .A(n5634), .B(n10394), .Z(n10396) );
  NAND U11109 ( .A(n10399), .B(e_input[317]), .Z(n5634) );
  NAND U11110 ( .A(n6112), .B(e_input[317]), .Z(n10399) );
  XOR U11111 ( .A(n10400), .B(n10401), .Z(n10394) );
  ANDN U11112 ( .A(n10402), .B(n5635), .Z(n10401) );
  XOR U11113 ( .A(n10403), .B(n10404), .Z(n5635) );
  IV U11114 ( .A(n10400), .Z(n10403) );
  XNOR U11115 ( .A(n5636), .B(n10400), .Z(n10402) );
  NAND U11116 ( .A(n10405), .B(e_input[316]), .Z(n5636) );
  NAND U11117 ( .A(n6112), .B(e_input[316]), .Z(n10405) );
  XOR U11118 ( .A(n10406), .B(n10407), .Z(n10400) );
  ANDN U11119 ( .A(n10408), .B(n5637), .Z(n10407) );
  XOR U11120 ( .A(n10409), .B(n10410), .Z(n5637) );
  IV U11121 ( .A(n10406), .Z(n10409) );
  XNOR U11122 ( .A(n5638), .B(n10406), .Z(n10408) );
  NAND U11123 ( .A(n10411), .B(e_input[315]), .Z(n5638) );
  NAND U11124 ( .A(n6112), .B(e_input[315]), .Z(n10411) );
  XOR U11125 ( .A(n10412), .B(n10413), .Z(n10406) );
  ANDN U11126 ( .A(n10414), .B(n5639), .Z(n10413) );
  XOR U11127 ( .A(n10415), .B(n10416), .Z(n5639) );
  IV U11128 ( .A(n10412), .Z(n10415) );
  XNOR U11129 ( .A(n5640), .B(n10412), .Z(n10414) );
  NAND U11130 ( .A(n10417), .B(e_input[314]), .Z(n5640) );
  NAND U11131 ( .A(n6112), .B(e_input[314]), .Z(n10417) );
  XOR U11132 ( .A(n10418), .B(n10419), .Z(n10412) );
  ANDN U11133 ( .A(n10420), .B(n5641), .Z(n10419) );
  XOR U11134 ( .A(n10421), .B(n10422), .Z(n5641) );
  IV U11135 ( .A(n10418), .Z(n10421) );
  XNOR U11136 ( .A(n5642), .B(n10418), .Z(n10420) );
  NAND U11137 ( .A(n10423), .B(e_input[313]), .Z(n5642) );
  NAND U11138 ( .A(n6112), .B(e_input[313]), .Z(n10423) );
  XOR U11139 ( .A(n10424), .B(n10425), .Z(n10418) );
  ANDN U11140 ( .A(n10426), .B(n5643), .Z(n10425) );
  XOR U11141 ( .A(n10427), .B(n10428), .Z(n5643) );
  IV U11142 ( .A(n10424), .Z(n10427) );
  XNOR U11143 ( .A(n5644), .B(n10424), .Z(n10426) );
  NAND U11144 ( .A(n10429), .B(e_input[312]), .Z(n5644) );
  NAND U11145 ( .A(n6112), .B(e_input[312]), .Z(n10429) );
  XOR U11146 ( .A(n10430), .B(n10431), .Z(n10424) );
  ANDN U11147 ( .A(n10432), .B(n5645), .Z(n10431) );
  XOR U11148 ( .A(n10433), .B(n10434), .Z(n5645) );
  IV U11149 ( .A(n10430), .Z(n10433) );
  XNOR U11150 ( .A(n5646), .B(n10430), .Z(n10432) );
  NAND U11151 ( .A(n10435), .B(e_input[311]), .Z(n5646) );
  NAND U11152 ( .A(n6112), .B(e_input[311]), .Z(n10435) );
  XOR U11153 ( .A(n10436), .B(n10437), .Z(n10430) );
  ANDN U11154 ( .A(n10438), .B(n5647), .Z(n10437) );
  XOR U11155 ( .A(n10439), .B(n10440), .Z(n5647) );
  IV U11156 ( .A(n10436), .Z(n10439) );
  XNOR U11157 ( .A(n5648), .B(n10436), .Z(n10438) );
  NAND U11158 ( .A(n10441), .B(e_input[310]), .Z(n5648) );
  NAND U11159 ( .A(n6112), .B(e_input[310]), .Z(n10441) );
  XOR U11160 ( .A(n10442), .B(n10443), .Z(n10436) );
  ANDN U11161 ( .A(n10444), .B(n5651), .Z(n10443) );
  XOR U11162 ( .A(n10445), .B(n10446), .Z(n5651) );
  IV U11163 ( .A(n10442), .Z(n10445) );
  XNOR U11164 ( .A(n5652), .B(n10442), .Z(n10444) );
  NAND U11165 ( .A(n10447), .B(e_input[309]), .Z(n5652) );
  NAND U11166 ( .A(n6112), .B(e_input[309]), .Z(n10447) );
  XOR U11167 ( .A(n10448), .B(n10449), .Z(n10442) );
  ANDN U11168 ( .A(n10450), .B(n5653), .Z(n10449) );
  XOR U11169 ( .A(n10451), .B(n10452), .Z(n5653) );
  IV U11170 ( .A(n10448), .Z(n10451) );
  XNOR U11171 ( .A(n5654), .B(n10448), .Z(n10450) );
  NAND U11172 ( .A(n10453), .B(e_input[308]), .Z(n5654) );
  NAND U11173 ( .A(n6112), .B(e_input[308]), .Z(n10453) );
  XOR U11174 ( .A(n10454), .B(n10455), .Z(n10448) );
  ANDN U11175 ( .A(n10456), .B(n5655), .Z(n10455) );
  XOR U11176 ( .A(n10457), .B(n10458), .Z(n5655) );
  IV U11177 ( .A(n10454), .Z(n10457) );
  XNOR U11178 ( .A(n5656), .B(n10454), .Z(n10456) );
  NAND U11179 ( .A(n10459), .B(e_input[307]), .Z(n5656) );
  NAND U11180 ( .A(n6112), .B(e_input[307]), .Z(n10459) );
  XOR U11181 ( .A(n10460), .B(n10461), .Z(n10454) );
  ANDN U11182 ( .A(n10462), .B(n5657), .Z(n10461) );
  XOR U11183 ( .A(n10463), .B(n10464), .Z(n5657) );
  IV U11184 ( .A(n10460), .Z(n10463) );
  XNOR U11185 ( .A(n5658), .B(n10460), .Z(n10462) );
  NAND U11186 ( .A(n10465), .B(e_input[306]), .Z(n5658) );
  NAND U11187 ( .A(n6112), .B(e_input[306]), .Z(n10465) );
  XOR U11188 ( .A(n10466), .B(n10467), .Z(n10460) );
  ANDN U11189 ( .A(n10468), .B(n5659), .Z(n10467) );
  XOR U11190 ( .A(n10469), .B(n10470), .Z(n5659) );
  IV U11191 ( .A(n10466), .Z(n10469) );
  XNOR U11192 ( .A(n5660), .B(n10466), .Z(n10468) );
  NAND U11193 ( .A(n10471), .B(e_input[305]), .Z(n5660) );
  NAND U11194 ( .A(n6112), .B(e_input[305]), .Z(n10471) );
  XOR U11195 ( .A(n10472), .B(n10473), .Z(n10466) );
  ANDN U11196 ( .A(n10474), .B(n5661), .Z(n10473) );
  XOR U11197 ( .A(n10475), .B(n10476), .Z(n5661) );
  IV U11198 ( .A(n10472), .Z(n10475) );
  XNOR U11199 ( .A(n5662), .B(n10472), .Z(n10474) );
  NAND U11200 ( .A(n10477), .B(e_input[304]), .Z(n5662) );
  NAND U11201 ( .A(n6112), .B(e_input[304]), .Z(n10477) );
  XOR U11202 ( .A(n10478), .B(n10479), .Z(n10472) );
  ANDN U11203 ( .A(n10480), .B(n5663), .Z(n10479) );
  XOR U11204 ( .A(n10481), .B(n10482), .Z(n5663) );
  IV U11205 ( .A(n10478), .Z(n10481) );
  XNOR U11206 ( .A(n5664), .B(n10478), .Z(n10480) );
  NAND U11207 ( .A(n10483), .B(e_input[303]), .Z(n5664) );
  NAND U11208 ( .A(n6112), .B(e_input[303]), .Z(n10483) );
  XOR U11209 ( .A(n10484), .B(n10485), .Z(n10478) );
  ANDN U11210 ( .A(n10486), .B(n5665), .Z(n10485) );
  XOR U11211 ( .A(n10487), .B(n10488), .Z(n5665) );
  IV U11212 ( .A(n10484), .Z(n10487) );
  XNOR U11213 ( .A(n5666), .B(n10484), .Z(n10486) );
  NAND U11214 ( .A(n10489), .B(e_input[302]), .Z(n5666) );
  NAND U11215 ( .A(n6112), .B(e_input[302]), .Z(n10489) );
  XOR U11216 ( .A(n10490), .B(n10491), .Z(n10484) );
  ANDN U11217 ( .A(n10492), .B(n5667), .Z(n10491) );
  XOR U11218 ( .A(n10493), .B(n10494), .Z(n5667) );
  IV U11219 ( .A(n10490), .Z(n10493) );
  XNOR U11220 ( .A(n5668), .B(n10490), .Z(n10492) );
  NAND U11221 ( .A(n10495), .B(e_input[301]), .Z(n5668) );
  NAND U11222 ( .A(n6112), .B(e_input[301]), .Z(n10495) );
  XOR U11223 ( .A(n10496), .B(n10497), .Z(n10490) );
  ANDN U11224 ( .A(n10498), .B(n5669), .Z(n10497) );
  XOR U11225 ( .A(n10499), .B(n10500), .Z(n5669) );
  IV U11226 ( .A(n10496), .Z(n10499) );
  XNOR U11227 ( .A(n5670), .B(n10496), .Z(n10498) );
  NAND U11228 ( .A(n10501), .B(e_input[300]), .Z(n5670) );
  NAND U11229 ( .A(n6112), .B(e_input[300]), .Z(n10501) );
  XOR U11230 ( .A(n10502), .B(n10503), .Z(n10496) );
  ANDN U11231 ( .A(n10504), .B(n5675), .Z(n10503) );
  XOR U11232 ( .A(n10505), .B(n10506), .Z(n5675) );
  IV U11233 ( .A(n10502), .Z(n10505) );
  XNOR U11234 ( .A(n5676), .B(n10502), .Z(n10504) );
  NAND U11235 ( .A(n10507), .B(e_input[299]), .Z(n5676) );
  NAND U11236 ( .A(n6112), .B(e_input[299]), .Z(n10507) );
  XOR U11237 ( .A(n10508), .B(n10509), .Z(n10502) );
  ANDN U11238 ( .A(n10510), .B(n5677), .Z(n10509) );
  XOR U11239 ( .A(n10511), .B(n10512), .Z(n5677) );
  IV U11240 ( .A(n10508), .Z(n10511) );
  XNOR U11241 ( .A(n5678), .B(n10508), .Z(n10510) );
  NAND U11242 ( .A(n10513), .B(e_input[298]), .Z(n5678) );
  NAND U11243 ( .A(n6112), .B(e_input[298]), .Z(n10513) );
  XOR U11244 ( .A(n10514), .B(n10515), .Z(n10508) );
  ANDN U11245 ( .A(n10516), .B(n5679), .Z(n10515) );
  XOR U11246 ( .A(n10517), .B(n10518), .Z(n5679) );
  IV U11247 ( .A(n10514), .Z(n10517) );
  XNOR U11248 ( .A(n5680), .B(n10514), .Z(n10516) );
  NAND U11249 ( .A(n10519), .B(e_input[297]), .Z(n5680) );
  NAND U11250 ( .A(n6112), .B(e_input[297]), .Z(n10519) );
  XOR U11251 ( .A(n10520), .B(n10521), .Z(n10514) );
  ANDN U11252 ( .A(n10522), .B(n5681), .Z(n10521) );
  XOR U11253 ( .A(n10523), .B(n10524), .Z(n5681) );
  IV U11254 ( .A(n10520), .Z(n10523) );
  XNOR U11255 ( .A(n5682), .B(n10520), .Z(n10522) );
  NAND U11256 ( .A(n10525), .B(e_input[296]), .Z(n5682) );
  NAND U11257 ( .A(n6112), .B(e_input[296]), .Z(n10525) );
  XOR U11258 ( .A(n10526), .B(n10527), .Z(n10520) );
  ANDN U11259 ( .A(n10528), .B(n5683), .Z(n10527) );
  XOR U11260 ( .A(n10529), .B(n10530), .Z(n5683) );
  IV U11261 ( .A(n10526), .Z(n10529) );
  XNOR U11262 ( .A(n5684), .B(n10526), .Z(n10528) );
  NAND U11263 ( .A(n10531), .B(e_input[295]), .Z(n5684) );
  NAND U11264 ( .A(n6112), .B(e_input[295]), .Z(n10531) );
  XOR U11265 ( .A(n10532), .B(n10533), .Z(n10526) );
  ANDN U11266 ( .A(n10534), .B(n5685), .Z(n10533) );
  XOR U11267 ( .A(n10535), .B(n10536), .Z(n5685) );
  IV U11268 ( .A(n10532), .Z(n10535) );
  XNOR U11269 ( .A(n5686), .B(n10532), .Z(n10534) );
  NAND U11270 ( .A(n10537), .B(e_input[294]), .Z(n5686) );
  NAND U11271 ( .A(n6112), .B(e_input[294]), .Z(n10537) );
  XOR U11272 ( .A(n10538), .B(n10539), .Z(n10532) );
  ANDN U11273 ( .A(n10540), .B(n5687), .Z(n10539) );
  XOR U11274 ( .A(n10541), .B(n10542), .Z(n5687) );
  IV U11275 ( .A(n10538), .Z(n10541) );
  XNOR U11276 ( .A(n5688), .B(n10538), .Z(n10540) );
  NAND U11277 ( .A(n10543), .B(e_input[293]), .Z(n5688) );
  NAND U11278 ( .A(n6112), .B(e_input[293]), .Z(n10543) );
  XOR U11279 ( .A(n10544), .B(n10545), .Z(n10538) );
  ANDN U11280 ( .A(n10546), .B(n5689), .Z(n10545) );
  XOR U11281 ( .A(n10547), .B(n10548), .Z(n5689) );
  IV U11282 ( .A(n10544), .Z(n10547) );
  XNOR U11283 ( .A(n5690), .B(n10544), .Z(n10546) );
  NAND U11284 ( .A(n10549), .B(e_input[292]), .Z(n5690) );
  NAND U11285 ( .A(n6112), .B(e_input[292]), .Z(n10549) );
  XOR U11286 ( .A(n10550), .B(n10551), .Z(n10544) );
  ANDN U11287 ( .A(n10552), .B(n5691), .Z(n10551) );
  XOR U11288 ( .A(n10553), .B(n10554), .Z(n5691) );
  IV U11289 ( .A(n10550), .Z(n10553) );
  XNOR U11290 ( .A(n5692), .B(n10550), .Z(n10552) );
  NAND U11291 ( .A(n10555), .B(e_input[291]), .Z(n5692) );
  NAND U11292 ( .A(n6112), .B(e_input[291]), .Z(n10555) );
  XOR U11293 ( .A(n10556), .B(n10557), .Z(n10550) );
  ANDN U11294 ( .A(n10558), .B(n5693), .Z(n10557) );
  XOR U11295 ( .A(n10559), .B(n10560), .Z(n5693) );
  IV U11296 ( .A(n10556), .Z(n10559) );
  XNOR U11297 ( .A(n5694), .B(n10556), .Z(n10558) );
  NAND U11298 ( .A(n10561), .B(e_input[290]), .Z(n5694) );
  NAND U11299 ( .A(n6112), .B(e_input[290]), .Z(n10561) );
  XOR U11300 ( .A(n10562), .B(n10563), .Z(n10556) );
  ANDN U11301 ( .A(n10564), .B(n5697), .Z(n10563) );
  XOR U11302 ( .A(n10565), .B(n10566), .Z(n5697) );
  IV U11303 ( .A(n10562), .Z(n10565) );
  XNOR U11304 ( .A(n5698), .B(n10562), .Z(n10564) );
  NAND U11305 ( .A(n10567), .B(e_input[289]), .Z(n5698) );
  NAND U11306 ( .A(n6112), .B(e_input[289]), .Z(n10567) );
  XOR U11307 ( .A(n10568), .B(n10569), .Z(n10562) );
  ANDN U11308 ( .A(n10570), .B(n5699), .Z(n10569) );
  XOR U11309 ( .A(n10571), .B(n10572), .Z(n5699) );
  IV U11310 ( .A(n10568), .Z(n10571) );
  XNOR U11311 ( .A(n5700), .B(n10568), .Z(n10570) );
  NAND U11312 ( .A(n10573), .B(e_input[288]), .Z(n5700) );
  NAND U11313 ( .A(n6112), .B(e_input[288]), .Z(n10573) );
  XOR U11314 ( .A(n10574), .B(n10575), .Z(n10568) );
  ANDN U11315 ( .A(n10576), .B(n5701), .Z(n10575) );
  XOR U11316 ( .A(n10577), .B(n10578), .Z(n5701) );
  IV U11317 ( .A(n10574), .Z(n10577) );
  XNOR U11318 ( .A(n5702), .B(n10574), .Z(n10576) );
  NAND U11319 ( .A(n10579), .B(e_input[287]), .Z(n5702) );
  NAND U11320 ( .A(n6112), .B(e_input[287]), .Z(n10579) );
  XOR U11321 ( .A(n10580), .B(n10581), .Z(n10574) );
  ANDN U11322 ( .A(n10582), .B(n5703), .Z(n10581) );
  XOR U11323 ( .A(n10583), .B(n10584), .Z(n5703) );
  IV U11324 ( .A(n10580), .Z(n10583) );
  XNOR U11325 ( .A(n5704), .B(n10580), .Z(n10582) );
  NAND U11326 ( .A(n10585), .B(e_input[286]), .Z(n5704) );
  NAND U11327 ( .A(n6112), .B(e_input[286]), .Z(n10585) );
  XOR U11328 ( .A(n10586), .B(n10587), .Z(n10580) );
  ANDN U11329 ( .A(n10588), .B(n5705), .Z(n10587) );
  XOR U11330 ( .A(n10589), .B(n10590), .Z(n5705) );
  IV U11331 ( .A(n10586), .Z(n10589) );
  XNOR U11332 ( .A(n5706), .B(n10586), .Z(n10588) );
  NAND U11333 ( .A(n10591), .B(e_input[285]), .Z(n5706) );
  NAND U11334 ( .A(n6112), .B(e_input[285]), .Z(n10591) );
  XOR U11335 ( .A(n10592), .B(n10593), .Z(n10586) );
  ANDN U11336 ( .A(n10594), .B(n5707), .Z(n10593) );
  XOR U11337 ( .A(n10595), .B(n10596), .Z(n5707) );
  IV U11338 ( .A(n10592), .Z(n10595) );
  XNOR U11339 ( .A(n5708), .B(n10592), .Z(n10594) );
  NAND U11340 ( .A(n10597), .B(e_input[284]), .Z(n5708) );
  NAND U11341 ( .A(n6112), .B(e_input[284]), .Z(n10597) );
  XOR U11342 ( .A(n10598), .B(n10599), .Z(n10592) );
  ANDN U11343 ( .A(n10600), .B(n5709), .Z(n10599) );
  XOR U11344 ( .A(n10601), .B(n10602), .Z(n5709) );
  IV U11345 ( .A(n10598), .Z(n10601) );
  XNOR U11346 ( .A(n5710), .B(n10598), .Z(n10600) );
  NAND U11347 ( .A(n10603), .B(e_input[283]), .Z(n5710) );
  NAND U11348 ( .A(n6112), .B(e_input[283]), .Z(n10603) );
  XOR U11349 ( .A(n10604), .B(n10605), .Z(n10598) );
  ANDN U11350 ( .A(n10606), .B(n5711), .Z(n10605) );
  XOR U11351 ( .A(n10607), .B(n10608), .Z(n5711) );
  IV U11352 ( .A(n10604), .Z(n10607) );
  XNOR U11353 ( .A(n5712), .B(n10604), .Z(n10606) );
  NAND U11354 ( .A(n10609), .B(e_input[282]), .Z(n5712) );
  NAND U11355 ( .A(n6112), .B(e_input[282]), .Z(n10609) );
  XOR U11356 ( .A(n10610), .B(n10611), .Z(n10604) );
  ANDN U11357 ( .A(n10612), .B(n5713), .Z(n10611) );
  XOR U11358 ( .A(n10613), .B(n10614), .Z(n5713) );
  IV U11359 ( .A(n10610), .Z(n10613) );
  XNOR U11360 ( .A(n5714), .B(n10610), .Z(n10612) );
  NAND U11361 ( .A(n10615), .B(e_input[281]), .Z(n5714) );
  NAND U11362 ( .A(n6112), .B(e_input[281]), .Z(n10615) );
  XOR U11363 ( .A(n10616), .B(n10617), .Z(n10610) );
  ANDN U11364 ( .A(n10618), .B(n5715), .Z(n10617) );
  XOR U11365 ( .A(n10619), .B(n10620), .Z(n5715) );
  IV U11366 ( .A(n10616), .Z(n10619) );
  XNOR U11367 ( .A(n5716), .B(n10616), .Z(n10618) );
  NAND U11368 ( .A(n10621), .B(e_input[280]), .Z(n5716) );
  NAND U11369 ( .A(n6112), .B(e_input[280]), .Z(n10621) );
  XOR U11370 ( .A(n10622), .B(n10623), .Z(n10616) );
  ANDN U11371 ( .A(n10624), .B(n5719), .Z(n10623) );
  XOR U11372 ( .A(n10625), .B(n10626), .Z(n5719) );
  IV U11373 ( .A(n10622), .Z(n10625) );
  XNOR U11374 ( .A(n5720), .B(n10622), .Z(n10624) );
  NAND U11375 ( .A(n10627), .B(e_input[279]), .Z(n5720) );
  NAND U11376 ( .A(n6112), .B(e_input[279]), .Z(n10627) );
  XOR U11377 ( .A(n10628), .B(n10629), .Z(n10622) );
  ANDN U11378 ( .A(n10630), .B(n5721), .Z(n10629) );
  XOR U11379 ( .A(n10631), .B(n10632), .Z(n5721) );
  IV U11380 ( .A(n10628), .Z(n10631) );
  XNOR U11381 ( .A(n5722), .B(n10628), .Z(n10630) );
  NAND U11382 ( .A(n10633), .B(e_input[278]), .Z(n5722) );
  NAND U11383 ( .A(n6112), .B(e_input[278]), .Z(n10633) );
  XOR U11384 ( .A(n10634), .B(n10635), .Z(n10628) );
  ANDN U11385 ( .A(n10636), .B(n5723), .Z(n10635) );
  XOR U11386 ( .A(n10637), .B(n10638), .Z(n5723) );
  IV U11387 ( .A(n10634), .Z(n10637) );
  XNOR U11388 ( .A(n5724), .B(n10634), .Z(n10636) );
  NAND U11389 ( .A(n10639), .B(e_input[277]), .Z(n5724) );
  NAND U11390 ( .A(n6112), .B(e_input[277]), .Z(n10639) );
  XOR U11391 ( .A(n10640), .B(n10641), .Z(n10634) );
  ANDN U11392 ( .A(n10642), .B(n5725), .Z(n10641) );
  XOR U11393 ( .A(n10643), .B(n10644), .Z(n5725) );
  IV U11394 ( .A(n10640), .Z(n10643) );
  XNOR U11395 ( .A(n5726), .B(n10640), .Z(n10642) );
  NAND U11396 ( .A(n10645), .B(e_input[276]), .Z(n5726) );
  NAND U11397 ( .A(n6112), .B(e_input[276]), .Z(n10645) );
  XOR U11398 ( .A(n10646), .B(n10647), .Z(n10640) );
  ANDN U11399 ( .A(n10648), .B(n5727), .Z(n10647) );
  XOR U11400 ( .A(n10649), .B(n10650), .Z(n5727) );
  IV U11401 ( .A(n10646), .Z(n10649) );
  XNOR U11402 ( .A(n5728), .B(n10646), .Z(n10648) );
  NAND U11403 ( .A(n10651), .B(e_input[275]), .Z(n5728) );
  NAND U11404 ( .A(n6112), .B(e_input[275]), .Z(n10651) );
  XOR U11405 ( .A(n10652), .B(n10653), .Z(n10646) );
  ANDN U11406 ( .A(n10654), .B(n5729), .Z(n10653) );
  XOR U11407 ( .A(n10655), .B(n10656), .Z(n5729) );
  IV U11408 ( .A(n10652), .Z(n10655) );
  XNOR U11409 ( .A(n5730), .B(n10652), .Z(n10654) );
  NAND U11410 ( .A(n10657), .B(e_input[274]), .Z(n5730) );
  NAND U11411 ( .A(n6112), .B(e_input[274]), .Z(n10657) );
  XOR U11412 ( .A(n10658), .B(n10659), .Z(n10652) );
  ANDN U11413 ( .A(n10660), .B(n5731), .Z(n10659) );
  XOR U11414 ( .A(n10661), .B(n10662), .Z(n5731) );
  IV U11415 ( .A(n10658), .Z(n10661) );
  XNOR U11416 ( .A(n5732), .B(n10658), .Z(n10660) );
  NAND U11417 ( .A(n10663), .B(e_input[273]), .Z(n5732) );
  NAND U11418 ( .A(n6112), .B(e_input[273]), .Z(n10663) );
  XOR U11419 ( .A(n10664), .B(n10665), .Z(n10658) );
  ANDN U11420 ( .A(n10666), .B(n5733), .Z(n10665) );
  XOR U11421 ( .A(n10667), .B(n10668), .Z(n5733) );
  IV U11422 ( .A(n10664), .Z(n10667) );
  XNOR U11423 ( .A(n5734), .B(n10664), .Z(n10666) );
  NAND U11424 ( .A(n10669), .B(e_input[272]), .Z(n5734) );
  NAND U11425 ( .A(n6112), .B(e_input[272]), .Z(n10669) );
  XOR U11426 ( .A(n10670), .B(n10671), .Z(n10664) );
  ANDN U11427 ( .A(n10672), .B(n5735), .Z(n10671) );
  XOR U11428 ( .A(n10673), .B(n10674), .Z(n5735) );
  IV U11429 ( .A(n10670), .Z(n10673) );
  XNOR U11430 ( .A(n5736), .B(n10670), .Z(n10672) );
  NAND U11431 ( .A(n10675), .B(e_input[271]), .Z(n5736) );
  NAND U11432 ( .A(n6112), .B(e_input[271]), .Z(n10675) );
  XOR U11433 ( .A(n10676), .B(n10677), .Z(n10670) );
  ANDN U11434 ( .A(n10678), .B(n5737), .Z(n10677) );
  XOR U11435 ( .A(n10679), .B(n10680), .Z(n5737) );
  IV U11436 ( .A(n10676), .Z(n10679) );
  XNOR U11437 ( .A(n5738), .B(n10676), .Z(n10678) );
  NAND U11438 ( .A(n10681), .B(e_input[270]), .Z(n5738) );
  NAND U11439 ( .A(n6112), .B(e_input[270]), .Z(n10681) );
  XOR U11440 ( .A(n10682), .B(n10683), .Z(n10676) );
  ANDN U11441 ( .A(n10684), .B(n5741), .Z(n10683) );
  XOR U11442 ( .A(n10685), .B(n10686), .Z(n5741) );
  IV U11443 ( .A(n10682), .Z(n10685) );
  XNOR U11444 ( .A(n5742), .B(n10682), .Z(n10684) );
  NAND U11445 ( .A(n10687), .B(e_input[269]), .Z(n5742) );
  NAND U11446 ( .A(n6112), .B(e_input[269]), .Z(n10687) );
  XOR U11447 ( .A(n10688), .B(n10689), .Z(n10682) );
  ANDN U11448 ( .A(n10690), .B(n5743), .Z(n10689) );
  XOR U11449 ( .A(n10691), .B(n10692), .Z(n5743) );
  IV U11450 ( .A(n10688), .Z(n10691) );
  XNOR U11451 ( .A(n5744), .B(n10688), .Z(n10690) );
  NAND U11452 ( .A(n10693), .B(e_input[268]), .Z(n5744) );
  NAND U11453 ( .A(n6112), .B(e_input[268]), .Z(n10693) );
  XOR U11454 ( .A(n10694), .B(n10695), .Z(n10688) );
  ANDN U11455 ( .A(n10696), .B(n5745), .Z(n10695) );
  XOR U11456 ( .A(n10697), .B(n10698), .Z(n5745) );
  IV U11457 ( .A(n10694), .Z(n10697) );
  XNOR U11458 ( .A(n5746), .B(n10694), .Z(n10696) );
  NAND U11459 ( .A(n10699), .B(e_input[267]), .Z(n5746) );
  NAND U11460 ( .A(n6112), .B(e_input[267]), .Z(n10699) );
  XOR U11461 ( .A(n10700), .B(n10701), .Z(n10694) );
  ANDN U11462 ( .A(n10702), .B(n5747), .Z(n10701) );
  XOR U11463 ( .A(n10703), .B(n10704), .Z(n5747) );
  IV U11464 ( .A(n10700), .Z(n10703) );
  XNOR U11465 ( .A(n5748), .B(n10700), .Z(n10702) );
  NAND U11466 ( .A(n10705), .B(e_input[266]), .Z(n5748) );
  NAND U11467 ( .A(n6112), .B(e_input[266]), .Z(n10705) );
  XOR U11468 ( .A(n10706), .B(n10707), .Z(n10700) );
  ANDN U11469 ( .A(n10708), .B(n5749), .Z(n10707) );
  XOR U11470 ( .A(n10709), .B(n10710), .Z(n5749) );
  IV U11471 ( .A(n10706), .Z(n10709) );
  XNOR U11472 ( .A(n5750), .B(n10706), .Z(n10708) );
  NAND U11473 ( .A(n10711), .B(e_input[265]), .Z(n5750) );
  NAND U11474 ( .A(n6112), .B(e_input[265]), .Z(n10711) );
  XOR U11475 ( .A(n10712), .B(n10713), .Z(n10706) );
  ANDN U11476 ( .A(n10714), .B(n5751), .Z(n10713) );
  XOR U11477 ( .A(n10715), .B(n10716), .Z(n5751) );
  IV U11478 ( .A(n10712), .Z(n10715) );
  XNOR U11479 ( .A(n5752), .B(n10712), .Z(n10714) );
  NAND U11480 ( .A(n10717), .B(e_input[264]), .Z(n5752) );
  NAND U11481 ( .A(n6112), .B(e_input[264]), .Z(n10717) );
  XOR U11482 ( .A(n10718), .B(n10719), .Z(n10712) );
  ANDN U11483 ( .A(n10720), .B(n5753), .Z(n10719) );
  XOR U11484 ( .A(n10721), .B(n10722), .Z(n5753) );
  IV U11485 ( .A(n10718), .Z(n10721) );
  XNOR U11486 ( .A(n5754), .B(n10718), .Z(n10720) );
  NAND U11487 ( .A(n10723), .B(e_input[263]), .Z(n5754) );
  NAND U11488 ( .A(n6112), .B(e_input[263]), .Z(n10723) );
  XOR U11489 ( .A(n10724), .B(n10725), .Z(n10718) );
  ANDN U11490 ( .A(n10726), .B(n5755), .Z(n10725) );
  XOR U11491 ( .A(n10727), .B(n10728), .Z(n5755) );
  IV U11492 ( .A(n10724), .Z(n10727) );
  XNOR U11493 ( .A(n5756), .B(n10724), .Z(n10726) );
  NAND U11494 ( .A(n10729), .B(e_input[262]), .Z(n5756) );
  NAND U11495 ( .A(n6112), .B(e_input[262]), .Z(n10729) );
  XOR U11496 ( .A(n10730), .B(n10731), .Z(n10724) );
  ANDN U11497 ( .A(n10732), .B(n5757), .Z(n10731) );
  XOR U11498 ( .A(n10733), .B(n10734), .Z(n5757) );
  IV U11499 ( .A(n10730), .Z(n10733) );
  XNOR U11500 ( .A(n5758), .B(n10730), .Z(n10732) );
  NAND U11501 ( .A(n10735), .B(e_input[261]), .Z(n5758) );
  NAND U11502 ( .A(n6112), .B(e_input[261]), .Z(n10735) );
  XOR U11503 ( .A(n10736), .B(n10737), .Z(n10730) );
  ANDN U11504 ( .A(n10738), .B(n5759), .Z(n10737) );
  XOR U11505 ( .A(n10739), .B(n10740), .Z(n5759) );
  IV U11506 ( .A(n10736), .Z(n10739) );
  XNOR U11507 ( .A(n5760), .B(n10736), .Z(n10738) );
  NAND U11508 ( .A(n10741), .B(e_input[260]), .Z(n5760) );
  NAND U11509 ( .A(n6112), .B(e_input[260]), .Z(n10741) );
  XOR U11510 ( .A(n10742), .B(n10743), .Z(n10736) );
  ANDN U11511 ( .A(n10744), .B(n5763), .Z(n10743) );
  XOR U11512 ( .A(n10745), .B(n10746), .Z(n5763) );
  IV U11513 ( .A(n10742), .Z(n10745) );
  XNOR U11514 ( .A(n5764), .B(n10742), .Z(n10744) );
  NAND U11515 ( .A(n10747), .B(e_input[259]), .Z(n5764) );
  NAND U11516 ( .A(n6112), .B(e_input[259]), .Z(n10747) );
  XOR U11517 ( .A(n10748), .B(n10749), .Z(n10742) );
  ANDN U11518 ( .A(n10750), .B(n5765), .Z(n10749) );
  XOR U11519 ( .A(n10751), .B(n10752), .Z(n5765) );
  IV U11520 ( .A(n10748), .Z(n10751) );
  XNOR U11521 ( .A(n5766), .B(n10748), .Z(n10750) );
  NAND U11522 ( .A(n10753), .B(e_input[258]), .Z(n5766) );
  NAND U11523 ( .A(n6112), .B(e_input[258]), .Z(n10753) );
  XOR U11524 ( .A(n10754), .B(n10755), .Z(n10748) );
  ANDN U11525 ( .A(n10756), .B(n5767), .Z(n10755) );
  XOR U11526 ( .A(n10757), .B(n10758), .Z(n5767) );
  IV U11527 ( .A(n10754), .Z(n10757) );
  XNOR U11528 ( .A(n5768), .B(n10754), .Z(n10756) );
  NAND U11529 ( .A(n10759), .B(e_input[257]), .Z(n5768) );
  NAND U11530 ( .A(n6112), .B(e_input[257]), .Z(n10759) );
  XOR U11531 ( .A(n10760), .B(n10761), .Z(n10754) );
  ANDN U11532 ( .A(n10762), .B(n5769), .Z(n10761) );
  XOR U11533 ( .A(n10763), .B(n10764), .Z(n5769) );
  IV U11534 ( .A(n10760), .Z(n10763) );
  XNOR U11535 ( .A(n5770), .B(n10760), .Z(n10762) );
  NAND U11536 ( .A(n10765), .B(e_input[256]), .Z(n5770) );
  NAND U11537 ( .A(n6112), .B(e_input[256]), .Z(n10765) );
  XOR U11538 ( .A(n10766), .B(n10767), .Z(n10760) );
  ANDN U11539 ( .A(n10768), .B(n5771), .Z(n10767) );
  XOR U11540 ( .A(n10769), .B(n10770), .Z(n5771) );
  IV U11541 ( .A(n10766), .Z(n10769) );
  XNOR U11542 ( .A(n5772), .B(n10766), .Z(n10768) );
  NAND U11543 ( .A(n10771), .B(e_input[255]), .Z(n5772) );
  NAND U11544 ( .A(n6112), .B(e_input[255]), .Z(n10771) );
  XOR U11545 ( .A(n10772), .B(n10773), .Z(n10766) );
  ANDN U11546 ( .A(n10774), .B(n5773), .Z(n10773) );
  XOR U11547 ( .A(n10775), .B(n10776), .Z(n5773) );
  IV U11548 ( .A(n10772), .Z(n10775) );
  XNOR U11549 ( .A(n5774), .B(n10772), .Z(n10774) );
  NAND U11550 ( .A(n10777), .B(e_input[254]), .Z(n5774) );
  NAND U11551 ( .A(n6112), .B(e_input[254]), .Z(n10777) );
  XOR U11552 ( .A(n10778), .B(n10779), .Z(n10772) );
  ANDN U11553 ( .A(n10780), .B(n5775), .Z(n10779) );
  XOR U11554 ( .A(n10781), .B(n10782), .Z(n5775) );
  IV U11555 ( .A(n10778), .Z(n10781) );
  XNOR U11556 ( .A(n5776), .B(n10778), .Z(n10780) );
  NAND U11557 ( .A(n10783), .B(e_input[253]), .Z(n5776) );
  NAND U11558 ( .A(n6112), .B(e_input[253]), .Z(n10783) );
  XOR U11559 ( .A(n10784), .B(n10785), .Z(n10778) );
  ANDN U11560 ( .A(n10786), .B(n5777), .Z(n10785) );
  XOR U11561 ( .A(n10787), .B(n10788), .Z(n5777) );
  IV U11562 ( .A(n10784), .Z(n10787) );
  XNOR U11563 ( .A(n5778), .B(n10784), .Z(n10786) );
  NAND U11564 ( .A(n10789), .B(e_input[252]), .Z(n5778) );
  NAND U11565 ( .A(n6112), .B(e_input[252]), .Z(n10789) );
  XOR U11566 ( .A(n10790), .B(n10791), .Z(n10784) );
  ANDN U11567 ( .A(n10792), .B(n5779), .Z(n10791) );
  XOR U11568 ( .A(n10793), .B(n10794), .Z(n5779) );
  IV U11569 ( .A(n10790), .Z(n10793) );
  XNOR U11570 ( .A(n5780), .B(n10790), .Z(n10792) );
  NAND U11571 ( .A(n10795), .B(e_input[251]), .Z(n5780) );
  NAND U11572 ( .A(n6112), .B(e_input[251]), .Z(n10795) );
  XOR U11573 ( .A(n10796), .B(n10797), .Z(n10790) );
  ANDN U11574 ( .A(n10798), .B(n5781), .Z(n10797) );
  XOR U11575 ( .A(n10799), .B(n10800), .Z(n5781) );
  IV U11576 ( .A(n10796), .Z(n10799) );
  XNOR U11577 ( .A(n5782), .B(n10796), .Z(n10798) );
  NAND U11578 ( .A(n10801), .B(e_input[250]), .Z(n5782) );
  NAND U11579 ( .A(n6112), .B(e_input[250]), .Z(n10801) );
  XOR U11580 ( .A(n10802), .B(n10803), .Z(n10796) );
  ANDN U11581 ( .A(n10804), .B(n5785), .Z(n10803) );
  XOR U11582 ( .A(n10805), .B(n10806), .Z(n5785) );
  IV U11583 ( .A(n10802), .Z(n10805) );
  XNOR U11584 ( .A(n5786), .B(n10802), .Z(n10804) );
  NAND U11585 ( .A(n10807), .B(e_input[249]), .Z(n5786) );
  NAND U11586 ( .A(n6112), .B(e_input[249]), .Z(n10807) );
  XOR U11587 ( .A(n10808), .B(n10809), .Z(n10802) );
  ANDN U11588 ( .A(n10810), .B(n5787), .Z(n10809) );
  XOR U11589 ( .A(n10811), .B(n10812), .Z(n5787) );
  IV U11590 ( .A(n10808), .Z(n10811) );
  XNOR U11591 ( .A(n5788), .B(n10808), .Z(n10810) );
  NAND U11592 ( .A(n10813), .B(e_input[248]), .Z(n5788) );
  NAND U11593 ( .A(n6112), .B(e_input[248]), .Z(n10813) );
  XOR U11594 ( .A(n10814), .B(n10815), .Z(n10808) );
  ANDN U11595 ( .A(n10816), .B(n5789), .Z(n10815) );
  XOR U11596 ( .A(n10817), .B(n10818), .Z(n5789) );
  IV U11597 ( .A(n10814), .Z(n10817) );
  XNOR U11598 ( .A(n5790), .B(n10814), .Z(n10816) );
  NAND U11599 ( .A(n10819), .B(e_input[247]), .Z(n5790) );
  NAND U11600 ( .A(n6112), .B(e_input[247]), .Z(n10819) );
  XOR U11601 ( .A(n10820), .B(n10821), .Z(n10814) );
  ANDN U11602 ( .A(n10822), .B(n5791), .Z(n10821) );
  XOR U11603 ( .A(n10823), .B(n10824), .Z(n5791) );
  IV U11604 ( .A(n10820), .Z(n10823) );
  XNOR U11605 ( .A(n5792), .B(n10820), .Z(n10822) );
  NAND U11606 ( .A(n10825), .B(e_input[246]), .Z(n5792) );
  NAND U11607 ( .A(n6112), .B(e_input[246]), .Z(n10825) );
  XOR U11608 ( .A(n10826), .B(n10827), .Z(n10820) );
  ANDN U11609 ( .A(n10828), .B(n5793), .Z(n10827) );
  XOR U11610 ( .A(n10829), .B(n10830), .Z(n5793) );
  IV U11611 ( .A(n10826), .Z(n10829) );
  XNOR U11612 ( .A(n5794), .B(n10826), .Z(n10828) );
  NAND U11613 ( .A(n10831), .B(e_input[245]), .Z(n5794) );
  NAND U11614 ( .A(n6112), .B(e_input[245]), .Z(n10831) );
  XOR U11615 ( .A(n10832), .B(n10833), .Z(n10826) );
  ANDN U11616 ( .A(n10834), .B(n5795), .Z(n10833) );
  XOR U11617 ( .A(n10835), .B(n10836), .Z(n5795) );
  IV U11618 ( .A(n10832), .Z(n10835) );
  XNOR U11619 ( .A(n5796), .B(n10832), .Z(n10834) );
  NAND U11620 ( .A(n10837), .B(e_input[244]), .Z(n5796) );
  NAND U11621 ( .A(n6112), .B(e_input[244]), .Z(n10837) );
  XOR U11622 ( .A(n10838), .B(n10839), .Z(n10832) );
  ANDN U11623 ( .A(n10840), .B(n5797), .Z(n10839) );
  XOR U11624 ( .A(n10841), .B(n10842), .Z(n5797) );
  IV U11625 ( .A(n10838), .Z(n10841) );
  XNOR U11626 ( .A(n5798), .B(n10838), .Z(n10840) );
  NAND U11627 ( .A(n10843), .B(e_input[243]), .Z(n5798) );
  NAND U11628 ( .A(n6112), .B(e_input[243]), .Z(n10843) );
  XOR U11629 ( .A(n10844), .B(n10845), .Z(n10838) );
  ANDN U11630 ( .A(n10846), .B(n5799), .Z(n10845) );
  XOR U11631 ( .A(n10847), .B(n10848), .Z(n5799) );
  IV U11632 ( .A(n10844), .Z(n10847) );
  XNOR U11633 ( .A(n5800), .B(n10844), .Z(n10846) );
  NAND U11634 ( .A(n10849), .B(e_input[242]), .Z(n5800) );
  NAND U11635 ( .A(n6112), .B(e_input[242]), .Z(n10849) );
  XOR U11636 ( .A(n10850), .B(n10851), .Z(n10844) );
  ANDN U11637 ( .A(n10852), .B(n5801), .Z(n10851) );
  XOR U11638 ( .A(n10853), .B(n10854), .Z(n5801) );
  IV U11639 ( .A(n10850), .Z(n10853) );
  XNOR U11640 ( .A(n5802), .B(n10850), .Z(n10852) );
  NAND U11641 ( .A(n10855), .B(e_input[241]), .Z(n5802) );
  NAND U11642 ( .A(n6112), .B(e_input[241]), .Z(n10855) );
  XOR U11643 ( .A(n10856), .B(n10857), .Z(n10850) );
  ANDN U11644 ( .A(n10858), .B(n5803), .Z(n10857) );
  XOR U11645 ( .A(n10859), .B(n10860), .Z(n5803) );
  IV U11646 ( .A(n10856), .Z(n10859) );
  XNOR U11647 ( .A(n5804), .B(n10856), .Z(n10858) );
  NAND U11648 ( .A(n10861), .B(e_input[240]), .Z(n5804) );
  NAND U11649 ( .A(n6112), .B(e_input[240]), .Z(n10861) );
  XOR U11650 ( .A(n10862), .B(n10863), .Z(n10856) );
  ANDN U11651 ( .A(n10864), .B(n5807), .Z(n10863) );
  XOR U11652 ( .A(n10865), .B(n10866), .Z(n5807) );
  IV U11653 ( .A(n10862), .Z(n10865) );
  XNOR U11654 ( .A(n5808), .B(n10862), .Z(n10864) );
  NAND U11655 ( .A(n10867), .B(e_input[239]), .Z(n5808) );
  NAND U11656 ( .A(n6112), .B(e_input[239]), .Z(n10867) );
  XOR U11657 ( .A(n10868), .B(n10869), .Z(n10862) );
  ANDN U11658 ( .A(n10870), .B(n5809), .Z(n10869) );
  XOR U11659 ( .A(n10871), .B(n10872), .Z(n5809) );
  IV U11660 ( .A(n10868), .Z(n10871) );
  XNOR U11661 ( .A(n5810), .B(n10868), .Z(n10870) );
  NAND U11662 ( .A(n10873), .B(e_input[238]), .Z(n5810) );
  NAND U11663 ( .A(n6112), .B(e_input[238]), .Z(n10873) );
  XOR U11664 ( .A(n10874), .B(n10875), .Z(n10868) );
  ANDN U11665 ( .A(n10876), .B(n5811), .Z(n10875) );
  XOR U11666 ( .A(n10877), .B(n10878), .Z(n5811) );
  IV U11667 ( .A(n10874), .Z(n10877) );
  XNOR U11668 ( .A(n5812), .B(n10874), .Z(n10876) );
  NAND U11669 ( .A(n10879), .B(e_input[237]), .Z(n5812) );
  NAND U11670 ( .A(n6112), .B(e_input[237]), .Z(n10879) );
  XOR U11671 ( .A(n10880), .B(n10881), .Z(n10874) );
  ANDN U11672 ( .A(n10882), .B(n5813), .Z(n10881) );
  XOR U11673 ( .A(n10883), .B(n10884), .Z(n5813) );
  IV U11674 ( .A(n10880), .Z(n10883) );
  XNOR U11675 ( .A(n5814), .B(n10880), .Z(n10882) );
  NAND U11676 ( .A(n10885), .B(e_input[236]), .Z(n5814) );
  NAND U11677 ( .A(n6112), .B(e_input[236]), .Z(n10885) );
  XOR U11678 ( .A(n10886), .B(n10887), .Z(n10880) );
  ANDN U11679 ( .A(n10888), .B(n5815), .Z(n10887) );
  XOR U11680 ( .A(n10889), .B(n10890), .Z(n5815) );
  IV U11681 ( .A(n10886), .Z(n10889) );
  XNOR U11682 ( .A(n5816), .B(n10886), .Z(n10888) );
  NAND U11683 ( .A(n10891), .B(e_input[235]), .Z(n5816) );
  NAND U11684 ( .A(n6112), .B(e_input[235]), .Z(n10891) );
  XOR U11685 ( .A(n10892), .B(n10893), .Z(n10886) );
  ANDN U11686 ( .A(n10894), .B(n5817), .Z(n10893) );
  XOR U11687 ( .A(n10895), .B(n10896), .Z(n5817) );
  IV U11688 ( .A(n10892), .Z(n10895) );
  XNOR U11689 ( .A(n5818), .B(n10892), .Z(n10894) );
  NAND U11690 ( .A(n10897), .B(e_input[234]), .Z(n5818) );
  NAND U11691 ( .A(n6112), .B(e_input[234]), .Z(n10897) );
  XOR U11692 ( .A(n10898), .B(n10899), .Z(n10892) );
  ANDN U11693 ( .A(n10900), .B(n5819), .Z(n10899) );
  XOR U11694 ( .A(n10901), .B(n10902), .Z(n5819) );
  IV U11695 ( .A(n10898), .Z(n10901) );
  XNOR U11696 ( .A(n5820), .B(n10898), .Z(n10900) );
  NAND U11697 ( .A(n10903), .B(e_input[233]), .Z(n5820) );
  NAND U11698 ( .A(n6112), .B(e_input[233]), .Z(n10903) );
  XOR U11699 ( .A(n10904), .B(n10905), .Z(n10898) );
  ANDN U11700 ( .A(n10906), .B(n5821), .Z(n10905) );
  XOR U11701 ( .A(n10907), .B(n10908), .Z(n5821) );
  IV U11702 ( .A(n10904), .Z(n10907) );
  XNOR U11703 ( .A(n5822), .B(n10904), .Z(n10906) );
  NAND U11704 ( .A(n10909), .B(e_input[232]), .Z(n5822) );
  NAND U11705 ( .A(n6112), .B(e_input[232]), .Z(n10909) );
  XOR U11706 ( .A(n10910), .B(n10911), .Z(n10904) );
  ANDN U11707 ( .A(n10912), .B(n5823), .Z(n10911) );
  XOR U11708 ( .A(n10913), .B(n10914), .Z(n5823) );
  IV U11709 ( .A(n10910), .Z(n10913) );
  XNOR U11710 ( .A(n5824), .B(n10910), .Z(n10912) );
  NAND U11711 ( .A(n10915), .B(e_input[231]), .Z(n5824) );
  NAND U11712 ( .A(n6112), .B(e_input[231]), .Z(n10915) );
  XOR U11713 ( .A(n10916), .B(n10917), .Z(n10910) );
  ANDN U11714 ( .A(n10918), .B(n5825), .Z(n10917) );
  XOR U11715 ( .A(n10919), .B(n10920), .Z(n5825) );
  IV U11716 ( .A(n10916), .Z(n10919) );
  XNOR U11717 ( .A(n5826), .B(n10916), .Z(n10918) );
  NAND U11718 ( .A(n10921), .B(e_input[230]), .Z(n5826) );
  NAND U11719 ( .A(n6112), .B(e_input[230]), .Z(n10921) );
  XOR U11720 ( .A(n10922), .B(n10923), .Z(n10916) );
  ANDN U11721 ( .A(n10924), .B(n5829), .Z(n10923) );
  XOR U11722 ( .A(n10925), .B(n10926), .Z(n5829) );
  IV U11723 ( .A(n10922), .Z(n10925) );
  XNOR U11724 ( .A(n5830), .B(n10922), .Z(n10924) );
  NAND U11725 ( .A(n10927), .B(e_input[229]), .Z(n5830) );
  NAND U11726 ( .A(n6112), .B(e_input[229]), .Z(n10927) );
  XOR U11727 ( .A(n10928), .B(n10929), .Z(n10922) );
  ANDN U11728 ( .A(n10930), .B(n5831), .Z(n10929) );
  XOR U11729 ( .A(n10931), .B(n10932), .Z(n5831) );
  IV U11730 ( .A(n10928), .Z(n10931) );
  XNOR U11731 ( .A(n5832), .B(n10928), .Z(n10930) );
  NAND U11732 ( .A(n10933), .B(e_input[228]), .Z(n5832) );
  NAND U11733 ( .A(n6112), .B(e_input[228]), .Z(n10933) );
  XOR U11734 ( .A(n10934), .B(n10935), .Z(n10928) );
  ANDN U11735 ( .A(n10936), .B(n5833), .Z(n10935) );
  XOR U11736 ( .A(n10937), .B(n10938), .Z(n5833) );
  IV U11737 ( .A(n10934), .Z(n10937) );
  XNOR U11738 ( .A(n5834), .B(n10934), .Z(n10936) );
  NAND U11739 ( .A(n10939), .B(e_input[227]), .Z(n5834) );
  NAND U11740 ( .A(n6112), .B(e_input[227]), .Z(n10939) );
  XOR U11741 ( .A(n10940), .B(n10941), .Z(n10934) );
  ANDN U11742 ( .A(n10942), .B(n5835), .Z(n10941) );
  XOR U11743 ( .A(n10943), .B(n10944), .Z(n5835) );
  IV U11744 ( .A(n10940), .Z(n10943) );
  XNOR U11745 ( .A(n5836), .B(n10940), .Z(n10942) );
  NAND U11746 ( .A(n10945), .B(e_input[226]), .Z(n5836) );
  NAND U11747 ( .A(n6112), .B(e_input[226]), .Z(n10945) );
  XOR U11748 ( .A(n10946), .B(n10947), .Z(n10940) );
  ANDN U11749 ( .A(n10948), .B(n5837), .Z(n10947) );
  XOR U11750 ( .A(n10949), .B(n10950), .Z(n5837) );
  IV U11751 ( .A(n10946), .Z(n10949) );
  XNOR U11752 ( .A(n5838), .B(n10946), .Z(n10948) );
  NAND U11753 ( .A(n10951), .B(e_input[225]), .Z(n5838) );
  NAND U11754 ( .A(n6112), .B(e_input[225]), .Z(n10951) );
  XOR U11755 ( .A(n10952), .B(n10953), .Z(n10946) );
  ANDN U11756 ( .A(n10954), .B(n5839), .Z(n10953) );
  XOR U11757 ( .A(n10955), .B(n10956), .Z(n5839) );
  IV U11758 ( .A(n10952), .Z(n10955) );
  XNOR U11759 ( .A(n5840), .B(n10952), .Z(n10954) );
  NAND U11760 ( .A(n10957), .B(e_input[224]), .Z(n5840) );
  NAND U11761 ( .A(n6112), .B(e_input[224]), .Z(n10957) );
  XOR U11762 ( .A(n10958), .B(n10959), .Z(n10952) );
  ANDN U11763 ( .A(n10960), .B(n5841), .Z(n10959) );
  XOR U11764 ( .A(n10961), .B(n10962), .Z(n5841) );
  IV U11765 ( .A(n10958), .Z(n10961) );
  XNOR U11766 ( .A(n5842), .B(n10958), .Z(n10960) );
  NAND U11767 ( .A(n10963), .B(e_input[223]), .Z(n5842) );
  NAND U11768 ( .A(n6112), .B(e_input[223]), .Z(n10963) );
  XOR U11769 ( .A(n10964), .B(n10965), .Z(n10958) );
  ANDN U11770 ( .A(n10966), .B(n5843), .Z(n10965) );
  XOR U11771 ( .A(n10967), .B(n10968), .Z(n5843) );
  IV U11772 ( .A(n10964), .Z(n10967) );
  XNOR U11773 ( .A(n5844), .B(n10964), .Z(n10966) );
  NAND U11774 ( .A(n10969), .B(e_input[222]), .Z(n5844) );
  NAND U11775 ( .A(n6112), .B(e_input[222]), .Z(n10969) );
  XOR U11776 ( .A(n10970), .B(n10971), .Z(n10964) );
  ANDN U11777 ( .A(n10972), .B(n5845), .Z(n10971) );
  XOR U11778 ( .A(n10973), .B(n10974), .Z(n5845) );
  IV U11779 ( .A(n10970), .Z(n10973) );
  XNOR U11780 ( .A(n5846), .B(n10970), .Z(n10972) );
  NAND U11781 ( .A(n10975), .B(e_input[221]), .Z(n5846) );
  NAND U11782 ( .A(n6112), .B(e_input[221]), .Z(n10975) );
  XOR U11783 ( .A(n10976), .B(n10977), .Z(n10970) );
  ANDN U11784 ( .A(n10978), .B(n5847), .Z(n10977) );
  XOR U11785 ( .A(n10979), .B(n10980), .Z(n5847) );
  IV U11786 ( .A(n10976), .Z(n10979) );
  XNOR U11787 ( .A(n5848), .B(n10976), .Z(n10978) );
  NAND U11788 ( .A(n10981), .B(e_input[220]), .Z(n5848) );
  NAND U11789 ( .A(n6112), .B(e_input[220]), .Z(n10981) );
  XOR U11790 ( .A(n10982), .B(n10983), .Z(n10976) );
  ANDN U11791 ( .A(n10984), .B(n5851), .Z(n10983) );
  XOR U11792 ( .A(n10985), .B(n10986), .Z(n5851) );
  IV U11793 ( .A(n10982), .Z(n10985) );
  XNOR U11794 ( .A(n5852), .B(n10982), .Z(n10984) );
  NAND U11795 ( .A(n10987), .B(e_input[219]), .Z(n5852) );
  NAND U11796 ( .A(n6112), .B(e_input[219]), .Z(n10987) );
  XOR U11797 ( .A(n10988), .B(n10989), .Z(n10982) );
  ANDN U11798 ( .A(n10990), .B(n5853), .Z(n10989) );
  XOR U11799 ( .A(n10991), .B(n10992), .Z(n5853) );
  IV U11800 ( .A(n10988), .Z(n10991) );
  XNOR U11801 ( .A(n5854), .B(n10988), .Z(n10990) );
  NAND U11802 ( .A(n10993), .B(e_input[218]), .Z(n5854) );
  NAND U11803 ( .A(n6112), .B(e_input[218]), .Z(n10993) );
  XOR U11804 ( .A(n10994), .B(n10995), .Z(n10988) );
  ANDN U11805 ( .A(n10996), .B(n5855), .Z(n10995) );
  XOR U11806 ( .A(n10997), .B(n10998), .Z(n5855) );
  IV U11807 ( .A(n10994), .Z(n10997) );
  XNOR U11808 ( .A(n5856), .B(n10994), .Z(n10996) );
  NAND U11809 ( .A(n10999), .B(e_input[217]), .Z(n5856) );
  NAND U11810 ( .A(n6112), .B(e_input[217]), .Z(n10999) );
  XOR U11811 ( .A(n11000), .B(n11001), .Z(n10994) );
  ANDN U11812 ( .A(n11002), .B(n5857), .Z(n11001) );
  XOR U11813 ( .A(n11003), .B(n11004), .Z(n5857) );
  IV U11814 ( .A(n11000), .Z(n11003) );
  XNOR U11815 ( .A(n5858), .B(n11000), .Z(n11002) );
  NAND U11816 ( .A(n11005), .B(e_input[216]), .Z(n5858) );
  NAND U11817 ( .A(n6112), .B(e_input[216]), .Z(n11005) );
  XOR U11818 ( .A(n11006), .B(n11007), .Z(n11000) );
  ANDN U11819 ( .A(n11008), .B(n5859), .Z(n11007) );
  XOR U11820 ( .A(n11009), .B(n11010), .Z(n5859) );
  IV U11821 ( .A(n11006), .Z(n11009) );
  XNOR U11822 ( .A(n5860), .B(n11006), .Z(n11008) );
  NAND U11823 ( .A(n11011), .B(e_input[215]), .Z(n5860) );
  NAND U11824 ( .A(n6112), .B(e_input[215]), .Z(n11011) );
  XOR U11825 ( .A(n11012), .B(n11013), .Z(n11006) );
  ANDN U11826 ( .A(n11014), .B(n5861), .Z(n11013) );
  XOR U11827 ( .A(n11015), .B(n11016), .Z(n5861) );
  IV U11828 ( .A(n11012), .Z(n11015) );
  XNOR U11829 ( .A(n5862), .B(n11012), .Z(n11014) );
  NAND U11830 ( .A(n11017), .B(e_input[214]), .Z(n5862) );
  NAND U11831 ( .A(n6112), .B(e_input[214]), .Z(n11017) );
  XOR U11832 ( .A(n11018), .B(n11019), .Z(n11012) );
  ANDN U11833 ( .A(n11020), .B(n5863), .Z(n11019) );
  XOR U11834 ( .A(n11021), .B(n11022), .Z(n5863) );
  IV U11835 ( .A(n11018), .Z(n11021) );
  XNOR U11836 ( .A(n5864), .B(n11018), .Z(n11020) );
  NAND U11837 ( .A(n11023), .B(e_input[213]), .Z(n5864) );
  NAND U11838 ( .A(n6112), .B(e_input[213]), .Z(n11023) );
  XOR U11839 ( .A(n11024), .B(n11025), .Z(n11018) );
  ANDN U11840 ( .A(n11026), .B(n5865), .Z(n11025) );
  XOR U11841 ( .A(n11027), .B(n11028), .Z(n5865) );
  IV U11842 ( .A(n11024), .Z(n11027) );
  XNOR U11843 ( .A(n5866), .B(n11024), .Z(n11026) );
  NAND U11844 ( .A(n11029), .B(e_input[212]), .Z(n5866) );
  NAND U11845 ( .A(n6112), .B(e_input[212]), .Z(n11029) );
  XOR U11846 ( .A(n11030), .B(n11031), .Z(n11024) );
  ANDN U11847 ( .A(n11032), .B(n5867), .Z(n11031) );
  XOR U11848 ( .A(n11033), .B(n11034), .Z(n5867) );
  IV U11849 ( .A(n11030), .Z(n11033) );
  XNOR U11850 ( .A(n5868), .B(n11030), .Z(n11032) );
  NAND U11851 ( .A(n11035), .B(e_input[211]), .Z(n5868) );
  NAND U11852 ( .A(n6112), .B(e_input[211]), .Z(n11035) );
  XOR U11853 ( .A(n11036), .B(n11037), .Z(n11030) );
  ANDN U11854 ( .A(n11038), .B(n5869), .Z(n11037) );
  XOR U11855 ( .A(n11039), .B(n11040), .Z(n5869) );
  IV U11856 ( .A(n11036), .Z(n11039) );
  XNOR U11857 ( .A(n5870), .B(n11036), .Z(n11038) );
  NAND U11858 ( .A(n11041), .B(e_input[210]), .Z(n5870) );
  NAND U11859 ( .A(n6112), .B(e_input[210]), .Z(n11041) );
  XOR U11860 ( .A(n11042), .B(n11043), .Z(n11036) );
  ANDN U11861 ( .A(n11044), .B(n5873), .Z(n11043) );
  XOR U11862 ( .A(n11045), .B(n11046), .Z(n5873) );
  IV U11863 ( .A(n11042), .Z(n11045) );
  XNOR U11864 ( .A(n5874), .B(n11042), .Z(n11044) );
  NAND U11865 ( .A(n11047), .B(e_input[209]), .Z(n5874) );
  NAND U11866 ( .A(n6112), .B(e_input[209]), .Z(n11047) );
  XOR U11867 ( .A(n11048), .B(n11049), .Z(n11042) );
  ANDN U11868 ( .A(n11050), .B(n5875), .Z(n11049) );
  XOR U11869 ( .A(n11051), .B(n11052), .Z(n5875) );
  IV U11870 ( .A(n11048), .Z(n11051) );
  XNOR U11871 ( .A(n5876), .B(n11048), .Z(n11050) );
  NAND U11872 ( .A(n11053), .B(e_input[208]), .Z(n5876) );
  NAND U11873 ( .A(n6112), .B(e_input[208]), .Z(n11053) );
  XOR U11874 ( .A(n11054), .B(n11055), .Z(n11048) );
  ANDN U11875 ( .A(n11056), .B(n5877), .Z(n11055) );
  XOR U11876 ( .A(n11057), .B(n11058), .Z(n5877) );
  IV U11877 ( .A(n11054), .Z(n11057) );
  XNOR U11878 ( .A(n5878), .B(n11054), .Z(n11056) );
  NAND U11879 ( .A(n11059), .B(e_input[207]), .Z(n5878) );
  NAND U11880 ( .A(n6112), .B(e_input[207]), .Z(n11059) );
  XOR U11881 ( .A(n11060), .B(n11061), .Z(n11054) );
  ANDN U11882 ( .A(n11062), .B(n5879), .Z(n11061) );
  XOR U11883 ( .A(n11063), .B(n11064), .Z(n5879) );
  IV U11884 ( .A(n11060), .Z(n11063) );
  XNOR U11885 ( .A(n5880), .B(n11060), .Z(n11062) );
  NAND U11886 ( .A(n11065), .B(e_input[206]), .Z(n5880) );
  NAND U11887 ( .A(n6112), .B(e_input[206]), .Z(n11065) );
  XOR U11888 ( .A(n11066), .B(n11067), .Z(n11060) );
  ANDN U11889 ( .A(n11068), .B(n5881), .Z(n11067) );
  XOR U11890 ( .A(n11069), .B(n11070), .Z(n5881) );
  IV U11891 ( .A(n11066), .Z(n11069) );
  XNOR U11892 ( .A(n5882), .B(n11066), .Z(n11068) );
  NAND U11893 ( .A(n11071), .B(e_input[205]), .Z(n5882) );
  NAND U11894 ( .A(n6112), .B(e_input[205]), .Z(n11071) );
  XOR U11895 ( .A(n11072), .B(n11073), .Z(n11066) );
  ANDN U11896 ( .A(n11074), .B(n5883), .Z(n11073) );
  XOR U11897 ( .A(n11075), .B(n11076), .Z(n5883) );
  IV U11898 ( .A(n11072), .Z(n11075) );
  XNOR U11899 ( .A(n5884), .B(n11072), .Z(n11074) );
  NAND U11900 ( .A(n11077), .B(e_input[204]), .Z(n5884) );
  NAND U11901 ( .A(n6112), .B(e_input[204]), .Z(n11077) );
  XOR U11902 ( .A(n11078), .B(n11079), .Z(n11072) );
  ANDN U11903 ( .A(n11080), .B(n5885), .Z(n11079) );
  XOR U11904 ( .A(n11081), .B(n11082), .Z(n5885) );
  IV U11905 ( .A(n11078), .Z(n11081) );
  XNOR U11906 ( .A(n5886), .B(n11078), .Z(n11080) );
  NAND U11907 ( .A(n11083), .B(e_input[203]), .Z(n5886) );
  NAND U11908 ( .A(n6112), .B(e_input[203]), .Z(n11083) );
  XOR U11909 ( .A(n11084), .B(n11085), .Z(n11078) );
  ANDN U11910 ( .A(n11086), .B(n5887), .Z(n11085) );
  XOR U11911 ( .A(n11087), .B(n11088), .Z(n5887) );
  IV U11912 ( .A(n11084), .Z(n11087) );
  XNOR U11913 ( .A(n5888), .B(n11084), .Z(n11086) );
  NAND U11914 ( .A(n11089), .B(e_input[202]), .Z(n5888) );
  NAND U11915 ( .A(n6112), .B(e_input[202]), .Z(n11089) );
  XOR U11916 ( .A(n11090), .B(n11091), .Z(n11084) );
  ANDN U11917 ( .A(n11092), .B(n5889), .Z(n11091) );
  XOR U11918 ( .A(n11093), .B(n11094), .Z(n5889) );
  IV U11919 ( .A(n11090), .Z(n11093) );
  XNOR U11920 ( .A(n5890), .B(n11090), .Z(n11092) );
  NAND U11921 ( .A(n11095), .B(e_input[201]), .Z(n5890) );
  NAND U11922 ( .A(n6112), .B(e_input[201]), .Z(n11095) );
  XOR U11923 ( .A(n11096), .B(n11097), .Z(n11090) );
  ANDN U11924 ( .A(n11098), .B(n5891), .Z(n11097) );
  XOR U11925 ( .A(n11099), .B(n11100), .Z(n5891) );
  IV U11926 ( .A(n11096), .Z(n11099) );
  XNOR U11927 ( .A(n5892), .B(n11096), .Z(n11098) );
  NAND U11928 ( .A(n11101), .B(e_input[200]), .Z(n5892) );
  NAND U11929 ( .A(n6112), .B(e_input[200]), .Z(n11101) );
  XOR U11930 ( .A(n11102), .B(n11103), .Z(n11096) );
  ANDN U11931 ( .A(n11104), .B(n5897), .Z(n11103) );
  XOR U11932 ( .A(n11105), .B(n11106), .Z(n5897) );
  IV U11933 ( .A(n11102), .Z(n11105) );
  XNOR U11934 ( .A(n5898), .B(n11102), .Z(n11104) );
  NAND U11935 ( .A(n11107), .B(e_input[199]), .Z(n5898) );
  NAND U11936 ( .A(n6112), .B(e_input[199]), .Z(n11107) );
  XOR U11937 ( .A(n11108), .B(n11109), .Z(n11102) );
  ANDN U11938 ( .A(n11110), .B(n5899), .Z(n11109) );
  XOR U11939 ( .A(n11111), .B(n11112), .Z(n5899) );
  IV U11940 ( .A(n11108), .Z(n11111) );
  XNOR U11941 ( .A(n5900), .B(n11108), .Z(n11110) );
  NAND U11942 ( .A(n11113), .B(e_input[198]), .Z(n5900) );
  NAND U11943 ( .A(n6112), .B(e_input[198]), .Z(n11113) );
  XOR U11944 ( .A(n11114), .B(n11115), .Z(n11108) );
  ANDN U11945 ( .A(n11116), .B(n5901), .Z(n11115) );
  XOR U11946 ( .A(n11117), .B(n11118), .Z(n5901) );
  IV U11947 ( .A(n11114), .Z(n11117) );
  XNOR U11948 ( .A(n5902), .B(n11114), .Z(n11116) );
  NAND U11949 ( .A(n11119), .B(e_input[197]), .Z(n5902) );
  NAND U11950 ( .A(n6112), .B(e_input[197]), .Z(n11119) );
  XOR U11951 ( .A(n11120), .B(n11121), .Z(n11114) );
  ANDN U11952 ( .A(n11122), .B(n5903), .Z(n11121) );
  XOR U11953 ( .A(n11123), .B(n11124), .Z(n5903) );
  IV U11954 ( .A(n11120), .Z(n11123) );
  XNOR U11955 ( .A(n5904), .B(n11120), .Z(n11122) );
  NAND U11956 ( .A(n11125), .B(e_input[196]), .Z(n5904) );
  NAND U11957 ( .A(n6112), .B(e_input[196]), .Z(n11125) );
  XOR U11958 ( .A(n11126), .B(n11127), .Z(n11120) );
  ANDN U11959 ( .A(n11128), .B(n5905), .Z(n11127) );
  XOR U11960 ( .A(n11129), .B(n11130), .Z(n5905) );
  IV U11961 ( .A(n11126), .Z(n11129) );
  XNOR U11962 ( .A(n5906), .B(n11126), .Z(n11128) );
  NAND U11963 ( .A(n11131), .B(e_input[195]), .Z(n5906) );
  NAND U11964 ( .A(n6112), .B(e_input[195]), .Z(n11131) );
  XOR U11965 ( .A(n11132), .B(n11133), .Z(n11126) );
  ANDN U11966 ( .A(n11134), .B(n5907), .Z(n11133) );
  XOR U11967 ( .A(n11135), .B(n11136), .Z(n5907) );
  IV U11968 ( .A(n11132), .Z(n11135) );
  XNOR U11969 ( .A(n5908), .B(n11132), .Z(n11134) );
  NAND U11970 ( .A(n11137), .B(e_input[194]), .Z(n5908) );
  NAND U11971 ( .A(n6112), .B(e_input[194]), .Z(n11137) );
  XOR U11972 ( .A(n11138), .B(n11139), .Z(n11132) );
  ANDN U11973 ( .A(n11140), .B(n5909), .Z(n11139) );
  XOR U11974 ( .A(n11141), .B(n11142), .Z(n5909) );
  IV U11975 ( .A(n11138), .Z(n11141) );
  XNOR U11976 ( .A(n5910), .B(n11138), .Z(n11140) );
  NAND U11977 ( .A(n11143), .B(e_input[193]), .Z(n5910) );
  NAND U11978 ( .A(n6112), .B(e_input[193]), .Z(n11143) );
  XOR U11979 ( .A(n11144), .B(n11145), .Z(n11138) );
  ANDN U11980 ( .A(n11146), .B(n5911), .Z(n11145) );
  XOR U11981 ( .A(n11147), .B(n11148), .Z(n5911) );
  IV U11982 ( .A(n11144), .Z(n11147) );
  XNOR U11983 ( .A(n5912), .B(n11144), .Z(n11146) );
  NAND U11984 ( .A(n11149), .B(e_input[192]), .Z(n5912) );
  NAND U11985 ( .A(n6112), .B(e_input[192]), .Z(n11149) );
  XOR U11986 ( .A(n11150), .B(n11151), .Z(n11144) );
  ANDN U11987 ( .A(n11152), .B(n5913), .Z(n11151) );
  XOR U11988 ( .A(n11153), .B(n11154), .Z(n5913) );
  IV U11989 ( .A(n11150), .Z(n11153) );
  XNOR U11990 ( .A(n5914), .B(n11150), .Z(n11152) );
  NAND U11991 ( .A(n11155), .B(e_input[191]), .Z(n5914) );
  NAND U11992 ( .A(n6112), .B(e_input[191]), .Z(n11155) );
  XOR U11993 ( .A(n11156), .B(n11157), .Z(n11150) );
  ANDN U11994 ( .A(n11158), .B(n5915), .Z(n11157) );
  XOR U11995 ( .A(n11159), .B(n11160), .Z(n5915) );
  IV U11996 ( .A(n11156), .Z(n11159) );
  XNOR U11997 ( .A(n5916), .B(n11156), .Z(n11158) );
  NAND U11998 ( .A(n11161), .B(e_input[190]), .Z(n5916) );
  NAND U11999 ( .A(n6112), .B(e_input[190]), .Z(n11161) );
  XOR U12000 ( .A(n11162), .B(n11163), .Z(n11156) );
  ANDN U12001 ( .A(n11164), .B(n5919), .Z(n11163) );
  XOR U12002 ( .A(n11165), .B(n11166), .Z(n5919) );
  IV U12003 ( .A(n11162), .Z(n11165) );
  XNOR U12004 ( .A(n5920), .B(n11162), .Z(n11164) );
  NAND U12005 ( .A(n11167), .B(e_input[189]), .Z(n5920) );
  NAND U12006 ( .A(n6112), .B(e_input[189]), .Z(n11167) );
  XOR U12007 ( .A(n11168), .B(n11169), .Z(n11162) );
  ANDN U12008 ( .A(n11170), .B(n5921), .Z(n11169) );
  XOR U12009 ( .A(n11171), .B(n11172), .Z(n5921) );
  IV U12010 ( .A(n11168), .Z(n11171) );
  XNOR U12011 ( .A(n5922), .B(n11168), .Z(n11170) );
  NAND U12012 ( .A(n11173), .B(e_input[188]), .Z(n5922) );
  NAND U12013 ( .A(n6112), .B(e_input[188]), .Z(n11173) );
  XOR U12014 ( .A(n11174), .B(n11175), .Z(n11168) );
  ANDN U12015 ( .A(n11176), .B(n5923), .Z(n11175) );
  XOR U12016 ( .A(n11177), .B(n11178), .Z(n5923) );
  IV U12017 ( .A(n11174), .Z(n11177) );
  XNOR U12018 ( .A(n5924), .B(n11174), .Z(n11176) );
  NAND U12019 ( .A(n11179), .B(e_input[187]), .Z(n5924) );
  NAND U12020 ( .A(n6112), .B(e_input[187]), .Z(n11179) );
  XOR U12021 ( .A(n11180), .B(n11181), .Z(n11174) );
  ANDN U12022 ( .A(n11182), .B(n5925), .Z(n11181) );
  XOR U12023 ( .A(n11183), .B(n11184), .Z(n5925) );
  IV U12024 ( .A(n11180), .Z(n11183) );
  XNOR U12025 ( .A(n5926), .B(n11180), .Z(n11182) );
  NAND U12026 ( .A(n11185), .B(e_input[186]), .Z(n5926) );
  NAND U12027 ( .A(n6112), .B(e_input[186]), .Z(n11185) );
  XOR U12028 ( .A(n11186), .B(n11187), .Z(n11180) );
  ANDN U12029 ( .A(n11188), .B(n5927), .Z(n11187) );
  XOR U12030 ( .A(n11189), .B(n11190), .Z(n5927) );
  IV U12031 ( .A(n11186), .Z(n11189) );
  XNOR U12032 ( .A(n5928), .B(n11186), .Z(n11188) );
  NAND U12033 ( .A(n11191), .B(e_input[185]), .Z(n5928) );
  NAND U12034 ( .A(n6112), .B(e_input[185]), .Z(n11191) );
  XOR U12035 ( .A(n11192), .B(n11193), .Z(n11186) );
  ANDN U12036 ( .A(n11194), .B(n5929), .Z(n11193) );
  XOR U12037 ( .A(n11195), .B(n11196), .Z(n5929) );
  IV U12038 ( .A(n11192), .Z(n11195) );
  XNOR U12039 ( .A(n5930), .B(n11192), .Z(n11194) );
  NAND U12040 ( .A(n11197), .B(e_input[184]), .Z(n5930) );
  NAND U12041 ( .A(n6112), .B(e_input[184]), .Z(n11197) );
  XOR U12042 ( .A(n11198), .B(n11199), .Z(n11192) );
  ANDN U12043 ( .A(n11200), .B(n5931), .Z(n11199) );
  XOR U12044 ( .A(n11201), .B(n11202), .Z(n5931) );
  IV U12045 ( .A(n11198), .Z(n11201) );
  XNOR U12046 ( .A(n5932), .B(n11198), .Z(n11200) );
  NAND U12047 ( .A(n11203), .B(e_input[183]), .Z(n5932) );
  NAND U12048 ( .A(n6112), .B(e_input[183]), .Z(n11203) );
  XOR U12049 ( .A(n11204), .B(n11205), .Z(n11198) );
  ANDN U12050 ( .A(n11206), .B(n5933), .Z(n11205) );
  XOR U12051 ( .A(n11207), .B(n11208), .Z(n5933) );
  IV U12052 ( .A(n11204), .Z(n11207) );
  XNOR U12053 ( .A(n5934), .B(n11204), .Z(n11206) );
  NAND U12054 ( .A(n11209), .B(e_input[182]), .Z(n5934) );
  NAND U12055 ( .A(n6112), .B(e_input[182]), .Z(n11209) );
  XOR U12056 ( .A(n11210), .B(n11211), .Z(n11204) );
  ANDN U12057 ( .A(n11212), .B(n5935), .Z(n11211) );
  XOR U12058 ( .A(n11213), .B(n11214), .Z(n5935) );
  IV U12059 ( .A(n11210), .Z(n11213) );
  XNOR U12060 ( .A(n5936), .B(n11210), .Z(n11212) );
  NAND U12061 ( .A(n11215), .B(e_input[181]), .Z(n5936) );
  NAND U12062 ( .A(n6112), .B(e_input[181]), .Z(n11215) );
  XOR U12063 ( .A(n11216), .B(n11217), .Z(n11210) );
  ANDN U12064 ( .A(n11218), .B(n5937), .Z(n11217) );
  XOR U12065 ( .A(n11219), .B(n11220), .Z(n5937) );
  IV U12066 ( .A(n11216), .Z(n11219) );
  XNOR U12067 ( .A(n5938), .B(n11216), .Z(n11218) );
  NAND U12068 ( .A(n11221), .B(e_input[180]), .Z(n5938) );
  NAND U12069 ( .A(n6112), .B(e_input[180]), .Z(n11221) );
  XOR U12070 ( .A(n11222), .B(n11223), .Z(n11216) );
  ANDN U12071 ( .A(n11224), .B(n5941), .Z(n11223) );
  XOR U12072 ( .A(n11225), .B(n11226), .Z(n5941) );
  IV U12073 ( .A(n11222), .Z(n11225) );
  XNOR U12074 ( .A(n5942), .B(n11222), .Z(n11224) );
  NAND U12075 ( .A(n11227), .B(e_input[179]), .Z(n5942) );
  NAND U12076 ( .A(n6112), .B(e_input[179]), .Z(n11227) );
  XOR U12077 ( .A(n11228), .B(n11229), .Z(n11222) );
  ANDN U12078 ( .A(n11230), .B(n5943), .Z(n11229) );
  XOR U12079 ( .A(n11231), .B(n11232), .Z(n5943) );
  IV U12080 ( .A(n11228), .Z(n11231) );
  XNOR U12081 ( .A(n5944), .B(n11228), .Z(n11230) );
  NAND U12082 ( .A(n11233), .B(e_input[178]), .Z(n5944) );
  NAND U12083 ( .A(n6112), .B(e_input[178]), .Z(n11233) );
  XOR U12084 ( .A(n11234), .B(n11235), .Z(n11228) );
  ANDN U12085 ( .A(n11236), .B(n5945), .Z(n11235) );
  XOR U12086 ( .A(n11237), .B(n11238), .Z(n5945) );
  IV U12087 ( .A(n11234), .Z(n11237) );
  XNOR U12088 ( .A(n5946), .B(n11234), .Z(n11236) );
  NAND U12089 ( .A(n11239), .B(e_input[177]), .Z(n5946) );
  NAND U12090 ( .A(n6112), .B(e_input[177]), .Z(n11239) );
  XOR U12091 ( .A(n11240), .B(n11241), .Z(n11234) );
  ANDN U12092 ( .A(n11242), .B(n5947), .Z(n11241) );
  XOR U12093 ( .A(n11243), .B(n11244), .Z(n5947) );
  IV U12094 ( .A(n11240), .Z(n11243) );
  XNOR U12095 ( .A(n5948), .B(n11240), .Z(n11242) );
  NAND U12096 ( .A(n11245), .B(e_input[176]), .Z(n5948) );
  NAND U12097 ( .A(n6112), .B(e_input[176]), .Z(n11245) );
  XOR U12098 ( .A(n11246), .B(n11247), .Z(n11240) );
  ANDN U12099 ( .A(n11248), .B(n5949), .Z(n11247) );
  XOR U12100 ( .A(n11249), .B(n11250), .Z(n5949) );
  IV U12101 ( .A(n11246), .Z(n11249) );
  XNOR U12102 ( .A(n5950), .B(n11246), .Z(n11248) );
  NAND U12103 ( .A(n11251), .B(e_input[175]), .Z(n5950) );
  NAND U12104 ( .A(n6112), .B(e_input[175]), .Z(n11251) );
  XOR U12105 ( .A(n11252), .B(n11253), .Z(n11246) );
  ANDN U12106 ( .A(n11254), .B(n5951), .Z(n11253) );
  XOR U12107 ( .A(n11255), .B(n11256), .Z(n5951) );
  IV U12108 ( .A(n11252), .Z(n11255) );
  XNOR U12109 ( .A(n5952), .B(n11252), .Z(n11254) );
  NAND U12110 ( .A(n11257), .B(e_input[174]), .Z(n5952) );
  NAND U12111 ( .A(n6112), .B(e_input[174]), .Z(n11257) );
  XOR U12112 ( .A(n11258), .B(n11259), .Z(n11252) );
  ANDN U12113 ( .A(n11260), .B(n5953), .Z(n11259) );
  XOR U12114 ( .A(n11261), .B(n11262), .Z(n5953) );
  IV U12115 ( .A(n11258), .Z(n11261) );
  XNOR U12116 ( .A(n5954), .B(n11258), .Z(n11260) );
  NAND U12117 ( .A(n11263), .B(e_input[173]), .Z(n5954) );
  NAND U12118 ( .A(n6112), .B(e_input[173]), .Z(n11263) );
  XOR U12119 ( .A(n11264), .B(n11265), .Z(n11258) );
  ANDN U12120 ( .A(n11266), .B(n5955), .Z(n11265) );
  XOR U12121 ( .A(n11267), .B(n11268), .Z(n5955) );
  IV U12122 ( .A(n11264), .Z(n11267) );
  XNOR U12123 ( .A(n5956), .B(n11264), .Z(n11266) );
  NAND U12124 ( .A(n11269), .B(e_input[172]), .Z(n5956) );
  NAND U12125 ( .A(n6112), .B(e_input[172]), .Z(n11269) );
  XOR U12126 ( .A(n11270), .B(n11271), .Z(n11264) );
  ANDN U12127 ( .A(n11272), .B(n5957), .Z(n11271) );
  XOR U12128 ( .A(n11273), .B(n11274), .Z(n5957) );
  IV U12129 ( .A(n11270), .Z(n11273) );
  XNOR U12130 ( .A(n5958), .B(n11270), .Z(n11272) );
  NAND U12131 ( .A(n11275), .B(e_input[171]), .Z(n5958) );
  NAND U12132 ( .A(n6112), .B(e_input[171]), .Z(n11275) );
  XOR U12133 ( .A(n11276), .B(n11277), .Z(n11270) );
  ANDN U12134 ( .A(n11278), .B(n5959), .Z(n11277) );
  XOR U12135 ( .A(n11279), .B(n11280), .Z(n5959) );
  IV U12136 ( .A(n11276), .Z(n11279) );
  XNOR U12137 ( .A(n5960), .B(n11276), .Z(n11278) );
  NAND U12138 ( .A(n11281), .B(e_input[170]), .Z(n5960) );
  NAND U12139 ( .A(n6112), .B(e_input[170]), .Z(n11281) );
  XOR U12140 ( .A(n11282), .B(n11283), .Z(n11276) );
  ANDN U12141 ( .A(n11284), .B(n5963), .Z(n11283) );
  XOR U12142 ( .A(n11285), .B(n11286), .Z(n5963) );
  IV U12143 ( .A(n11282), .Z(n11285) );
  XNOR U12144 ( .A(n5964), .B(n11282), .Z(n11284) );
  NAND U12145 ( .A(n11287), .B(e_input[169]), .Z(n5964) );
  NAND U12146 ( .A(n6112), .B(e_input[169]), .Z(n11287) );
  XOR U12147 ( .A(n11288), .B(n11289), .Z(n11282) );
  ANDN U12148 ( .A(n11290), .B(n5965), .Z(n11289) );
  XOR U12149 ( .A(n11291), .B(n11292), .Z(n5965) );
  IV U12150 ( .A(n11288), .Z(n11291) );
  XNOR U12151 ( .A(n5966), .B(n11288), .Z(n11290) );
  NAND U12152 ( .A(n11293), .B(e_input[168]), .Z(n5966) );
  NAND U12153 ( .A(n6112), .B(e_input[168]), .Z(n11293) );
  XOR U12154 ( .A(n11294), .B(n11295), .Z(n11288) );
  ANDN U12155 ( .A(n11296), .B(n5967), .Z(n11295) );
  XOR U12156 ( .A(n11297), .B(n11298), .Z(n5967) );
  IV U12157 ( .A(n11294), .Z(n11297) );
  XNOR U12158 ( .A(n5968), .B(n11294), .Z(n11296) );
  NAND U12159 ( .A(n11299), .B(e_input[167]), .Z(n5968) );
  NAND U12160 ( .A(n6112), .B(e_input[167]), .Z(n11299) );
  XOR U12161 ( .A(n11300), .B(n11301), .Z(n11294) );
  ANDN U12162 ( .A(n11302), .B(n5969), .Z(n11301) );
  XOR U12163 ( .A(n11303), .B(n11304), .Z(n5969) );
  IV U12164 ( .A(n11300), .Z(n11303) );
  XNOR U12165 ( .A(n5970), .B(n11300), .Z(n11302) );
  NAND U12166 ( .A(n11305), .B(e_input[166]), .Z(n5970) );
  NAND U12167 ( .A(n6112), .B(e_input[166]), .Z(n11305) );
  XOR U12168 ( .A(n11306), .B(n11307), .Z(n11300) );
  ANDN U12169 ( .A(n11308), .B(n5971), .Z(n11307) );
  XOR U12170 ( .A(n11309), .B(n11310), .Z(n5971) );
  IV U12171 ( .A(n11306), .Z(n11309) );
  XNOR U12172 ( .A(n5972), .B(n11306), .Z(n11308) );
  NAND U12173 ( .A(n11311), .B(e_input[165]), .Z(n5972) );
  NAND U12174 ( .A(n6112), .B(e_input[165]), .Z(n11311) );
  XOR U12175 ( .A(n11312), .B(n11313), .Z(n11306) );
  ANDN U12176 ( .A(n11314), .B(n5973), .Z(n11313) );
  XOR U12177 ( .A(n11315), .B(n11316), .Z(n5973) );
  IV U12178 ( .A(n11312), .Z(n11315) );
  XNOR U12179 ( .A(n5974), .B(n11312), .Z(n11314) );
  NAND U12180 ( .A(n11317), .B(e_input[164]), .Z(n5974) );
  NAND U12181 ( .A(n6112), .B(e_input[164]), .Z(n11317) );
  XOR U12182 ( .A(n11318), .B(n11319), .Z(n11312) );
  ANDN U12183 ( .A(n11320), .B(n5975), .Z(n11319) );
  XOR U12184 ( .A(n11321), .B(n11322), .Z(n5975) );
  IV U12185 ( .A(n11318), .Z(n11321) );
  XNOR U12186 ( .A(n5976), .B(n11318), .Z(n11320) );
  NAND U12187 ( .A(n11323), .B(e_input[163]), .Z(n5976) );
  NAND U12188 ( .A(n6112), .B(e_input[163]), .Z(n11323) );
  XOR U12189 ( .A(n11324), .B(n11325), .Z(n11318) );
  ANDN U12190 ( .A(n11326), .B(n5977), .Z(n11325) );
  XOR U12191 ( .A(n11327), .B(n11328), .Z(n5977) );
  IV U12192 ( .A(n11324), .Z(n11327) );
  XNOR U12193 ( .A(n5978), .B(n11324), .Z(n11326) );
  NAND U12194 ( .A(n11329), .B(e_input[162]), .Z(n5978) );
  NAND U12195 ( .A(n6112), .B(e_input[162]), .Z(n11329) );
  XOR U12196 ( .A(n11330), .B(n11331), .Z(n11324) );
  ANDN U12197 ( .A(n11332), .B(n5979), .Z(n11331) );
  XOR U12198 ( .A(n11333), .B(n11334), .Z(n5979) );
  IV U12199 ( .A(n11330), .Z(n11333) );
  XNOR U12200 ( .A(n5980), .B(n11330), .Z(n11332) );
  NAND U12201 ( .A(n11335), .B(e_input[161]), .Z(n5980) );
  NAND U12202 ( .A(n6112), .B(e_input[161]), .Z(n11335) );
  XOR U12203 ( .A(n11336), .B(n11337), .Z(n11330) );
  ANDN U12204 ( .A(n11338), .B(n5981), .Z(n11337) );
  XOR U12205 ( .A(n11339), .B(n11340), .Z(n5981) );
  IV U12206 ( .A(n11336), .Z(n11339) );
  XNOR U12207 ( .A(n5982), .B(n11336), .Z(n11338) );
  NAND U12208 ( .A(n11341), .B(e_input[160]), .Z(n5982) );
  NAND U12209 ( .A(n6112), .B(e_input[160]), .Z(n11341) );
  XOR U12210 ( .A(n11342), .B(n11343), .Z(n11336) );
  ANDN U12211 ( .A(n11344), .B(n5985), .Z(n11343) );
  XOR U12212 ( .A(n11345), .B(n11346), .Z(n5985) );
  IV U12213 ( .A(n11342), .Z(n11345) );
  XNOR U12214 ( .A(n5986), .B(n11342), .Z(n11344) );
  NAND U12215 ( .A(n11347), .B(e_input[159]), .Z(n5986) );
  NAND U12216 ( .A(n6112), .B(e_input[159]), .Z(n11347) );
  XOR U12217 ( .A(n11348), .B(n11349), .Z(n11342) );
  ANDN U12218 ( .A(n11350), .B(n5987), .Z(n11349) );
  XOR U12219 ( .A(n11351), .B(n11352), .Z(n5987) );
  IV U12220 ( .A(n11348), .Z(n11351) );
  XNOR U12221 ( .A(n5988), .B(n11348), .Z(n11350) );
  NAND U12222 ( .A(n11353), .B(e_input[158]), .Z(n5988) );
  NAND U12223 ( .A(n6112), .B(e_input[158]), .Z(n11353) );
  XOR U12224 ( .A(n11354), .B(n11355), .Z(n11348) );
  ANDN U12225 ( .A(n11356), .B(n5989), .Z(n11355) );
  XOR U12226 ( .A(n11357), .B(n11358), .Z(n5989) );
  IV U12227 ( .A(n11354), .Z(n11357) );
  XNOR U12228 ( .A(n5990), .B(n11354), .Z(n11356) );
  NAND U12229 ( .A(n11359), .B(e_input[157]), .Z(n5990) );
  NAND U12230 ( .A(n6112), .B(e_input[157]), .Z(n11359) );
  XOR U12231 ( .A(n11360), .B(n11361), .Z(n11354) );
  ANDN U12232 ( .A(n11362), .B(n5991), .Z(n11361) );
  XOR U12233 ( .A(n11363), .B(n11364), .Z(n5991) );
  IV U12234 ( .A(n11360), .Z(n11363) );
  XNOR U12235 ( .A(n5992), .B(n11360), .Z(n11362) );
  NAND U12236 ( .A(n11365), .B(e_input[156]), .Z(n5992) );
  NAND U12237 ( .A(n6112), .B(e_input[156]), .Z(n11365) );
  XOR U12238 ( .A(n11366), .B(n11367), .Z(n11360) );
  ANDN U12239 ( .A(n11368), .B(n5993), .Z(n11367) );
  XOR U12240 ( .A(n11369), .B(n11370), .Z(n5993) );
  IV U12241 ( .A(n11366), .Z(n11369) );
  XNOR U12242 ( .A(n5994), .B(n11366), .Z(n11368) );
  NAND U12243 ( .A(n11371), .B(e_input[155]), .Z(n5994) );
  NAND U12244 ( .A(n6112), .B(e_input[155]), .Z(n11371) );
  XOR U12245 ( .A(n11372), .B(n11373), .Z(n11366) );
  ANDN U12246 ( .A(n11374), .B(n5995), .Z(n11373) );
  XOR U12247 ( .A(n11375), .B(n11376), .Z(n5995) );
  IV U12248 ( .A(n11372), .Z(n11375) );
  XNOR U12249 ( .A(n5996), .B(n11372), .Z(n11374) );
  NAND U12250 ( .A(n11377), .B(e_input[154]), .Z(n5996) );
  NAND U12251 ( .A(n6112), .B(e_input[154]), .Z(n11377) );
  XOR U12252 ( .A(n11378), .B(n11379), .Z(n11372) );
  ANDN U12253 ( .A(n11380), .B(n5997), .Z(n11379) );
  XOR U12254 ( .A(n11381), .B(n11382), .Z(n5997) );
  IV U12255 ( .A(n11378), .Z(n11381) );
  XNOR U12256 ( .A(n5998), .B(n11378), .Z(n11380) );
  NAND U12257 ( .A(n11383), .B(e_input[153]), .Z(n5998) );
  NAND U12258 ( .A(n6112), .B(e_input[153]), .Z(n11383) );
  XOR U12259 ( .A(n11384), .B(n11385), .Z(n11378) );
  ANDN U12260 ( .A(n11386), .B(n5999), .Z(n11385) );
  XOR U12261 ( .A(n11387), .B(n11388), .Z(n5999) );
  IV U12262 ( .A(n11384), .Z(n11387) );
  XNOR U12263 ( .A(n6000), .B(n11384), .Z(n11386) );
  NAND U12264 ( .A(n11389), .B(e_input[152]), .Z(n6000) );
  NAND U12265 ( .A(n6112), .B(e_input[152]), .Z(n11389) );
  XOR U12266 ( .A(n11390), .B(n11391), .Z(n11384) );
  ANDN U12267 ( .A(n11392), .B(n6001), .Z(n11391) );
  XOR U12268 ( .A(n11393), .B(n11394), .Z(n6001) );
  IV U12269 ( .A(n11390), .Z(n11393) );
  XNOR U12270 ( .A(n6002), .B(n11390), .Z(n11392) );
  NAND U12271 ( .A(n11395), .B(e_input[151]), .Z(n6002) );
  NAND U12272 ( .A(n6112), .B(e_input[151]), .Z(n11395) );
  XOR U12273 ( .A(n11396), .B(n11397), .Z(n11390) );
  ANDN U12274 ( .A(n11398), .B(n6003), .Z(n11397) );
  XOR U12275 ( .A(n11399), .B(n11400), .Z(n6003) );
  IV U12276 ( .A(n11396), .Z(n11399) );
  XNOR U12277 ( .A(n6004), .B(n11396), .Z(n11398) );
  NAND U12278 ( .A(n11401), .B(e_input[150]), .Z(n6004) );
  NAND U12279 ( .A(n6112), .B(e_input[150]), .Z(n11401) );
  XOR U12280 ( .A(n11402), .B(n11403), .Z(n11396) );
  ANDN U12281 ( .A(n11404), .B(n6007), .Z(n11403) );
  XOR U12282 ( .A(n11405), .B(n11406), .Z(n6007) );
  IV U12283 ( .A(n11402), .Z(n11405) );
  XNOR U12284 ( .A(n6008), .B(n11402), .Z(n11404) );
  NAND U12285 ( .A(n11407), .B(e_input[149]), .Z(n6008) );
  NAND U12286 ( .A(n6112), .B(e_input[149]), .Z(n11407) );
  XOR U12287 ( .A(n11408), .B(n11409), .Z(n11402) );
  ANDN U12288 ( .A(n11410), .B(n6009), .Z(n11409) );
  XOR U12289 ( .A(n11411), .B(n11412), .Z(n6009) );
  IV U12290 ( .A(n11408), .Z(n11411) );
  XNOR U12291 ( .A(n6010), .B(n11408), .Z(n11410) );
  NAND U12292 ( .A(n11413), .B(e_input[148]), .Z(n6010) );
  NAND U12293 ( .A(n6112), .B(e_input[148]), .Z(n11413) );
  XOR U12294 ( .A(n11414), .B(n11415), .Z(n11408) );
  ANDN U12295 ( .A(n11416), .B(n6011), .Z(n11415) );
  XOR U12296 ( .A(n11417), .B(n11418), .Z(n6011) );
  IV U12297 ( .A(n11414), .Z(n11417) );
  XNOR U12298 ( .A(n6012), .B(n11414), .Z(n11416) );
  NAND U12299 ( .A(n11419), .B(e_input[147]), .Z(n6012) );
  NAND U12300 ( .A(n6112), .B(e_input[147]), .Z(n11419) );
  XOR U12301 ( .A(n11420), .B(n11421), .Z(n11414) );
  ANDN U12302 ( .A(n11422), .B(n6013), .Z(n11421) );
  XOR U12303 ( .A(n11423), .B(n11424), .Z(n6013) );
  IV U12304 ( .A(n11420), .Z(n11423) );
  XNOR U12305 ( .A(n6014), .B(n11420), .Z(n11422) );
  NAND U12306 ( .A(n11425), .B(e_input[146]), .Z(n6014) );
  NAND U12307 ( .A(n6112), .B(e_input[146]), .Z(n11425) );
  XOR U12308 ( .A(n11426), .B(n11427), .Z(n11420) );
  ANDN U12309 ( .A(n11428), .B(n6015), .Z(n11427) );
  XOR U12310 ( .A(n11429), .B(n11430), .Z(n6015) );
  IV U12311 ( .A(n11426), .Z(n11429) );
  XNOR U12312 ( .A(n6016), .B(n11426), .Z(n11428) );
  NAND U12313 ( .A(n11431), .B(e_input[145]), .Z(n6016) );
  NAND U12314 ( .A(n6112), .B(e_input[145]), .Z(n11431) );
  XOR U12315 ( .A(n11432), .B(n11433), .Z(n11426) );
  ANDN U12316 ( .A(n11434), .B(n6017), .Z(n11433) );
  XOR U12317 ( .A(n11435), .B(n11436), .Z(n6017) );
  IV U12318 ( .A(n11432), .Z(n11435) );
  XNOR U12319 ( .A(n6018), .B(n11432), .Z(n11434) );
  NAND U12320 ( .A(n11437), .B(e_input[144]), .Z(n6018) );
  NAND U12321 ( .A(n6112), .B(e_input[144]), .Z(n11437) );
  XOR U12322 ( .A(n11438), .B(n11439), .Z(n11432) );
  ANDN U12323 ( .A(n11440), .B(n6019), .Z(n11439) );
  XOR U12324 ( .A(n11441), .B(n11442), .Z(n6019) );
  IV U12325 ( .A(n11438), .Z(n11441) );
  XNOR U12326 ( .A(n6020), .B(n11438), .Z(n11440) );
  NAND U12327 ( .A(n11443), .B(e_input[143]), .Z(n6020) );
  NAND U12328 ( .A(n6112), .B(e_input[143]), .Z(n11443) );
  XOR U12329 ( .A(n11444), .B(n11445), .Z(n11438) );
  ANDN U12330 ( .A(n11446), .B(n6021), .Z(n11445) );
  XOR U12331 ( .A(n11447), .B(n11448), .Z(n6021) );
  IV U12332 ( .A(n11444), .Z(n11447) );
  XNOR U12333 ( .A(n6022), .B(n11444), .Z(n11446) );
  NAND U12334 ( .A(n11449), .B(e_input[142]), .Z(n6022) );
  NAND U12335 ( .A(n6112), .B(e_input[142]), .Z(n11449) );
  XOR U12336 ( .A(n11450), .B(n11451), .Z(n11444) );
  ANDN U12337 ( .A(n11452), .B(n6023), .Z(n11451) );
  XOR U12338 ( .A(n11453), .B(n11454), .Z(n6023) );
  IV U12339 ( .A(n11450), .Z(n11453) );
  XNOR U12340 ( .A(n6024), .B(n11450), .Z(n11452) );
  NAND U12341 ( .A(n11455), .B(e_input[141]), .Z(n6024) );
  NAND U12342 ( .A(n6112), .B(e_input[141]), .Z(n11455) );
  XOR U12343 ( .A(n11456), .B(n11457), .Z(n11450) );
  ANDN U12344 ( .A(n11458), .B(n6025), .Z(n11457) );
  XOR U12345 ( .A(n11459), .B(n11460), .Z(n6025) );
  IV U12346 ( .A(n11456), .Z(n11459) );
  XNOR U12347 ( .A(n6026), .B(n11456), .Z(n11458) );
  NAND U12348 ( .A(n11461), .B(e_input[140]), .Z(n6026) );
  NAND U12349 ( .A(n6112), .B(e_input[140]), .Z(n11461) );
  XOR U12350 ( .A(n11462), .B(n11463), .Z(n11456) );
  ANDN U12351 ( .A(n11464), .B(n6029), .Z(n11463) );
  XOR U12352 ( .A(n11465), .B(n11466), .Z(n6029) );
  IV U12353 ( .A(n11462), .Z(n11465) );
  XNOR U12354 ( .A(n6030), .B(n11462), .Z(n11464) );
  NAND U12355 ( .A(n11467), .B(e_input[139]), .Z(n6030) );
  NAND U12356 ( .A(n6112), .B(e_input[139]), .Z(n11467) );
  XOR U12357 ( .A(n11468), .B(n11469), .Z(n11462) );
  ANDN U12358 ( .A(n11470), .B(n6031), .Z(n11469) );
  XOR U12359 ( .A(n11471), .B(n11472), .Z(n6031) );
  IV U12360 ( .A(n11468), .Z(n11471) );
  XNOR U12361 ( .A(n6032), .B(n11468), .Z(n11470) );
  NAND U12362 ( .A(n11473), .B(e_input[138]), .Z(n6032) );
  NAND U12363 ( .A(n6112), .B(e_input[138]), .Z(n11473) );
  XOR U12364 ( .A(n11474), .B(n11475), .Z(n11468) );
  ANDN U12365 ( .A(n11476), .B(n6033), .Z(n11475) );
  XOR U12366 ( .A(n11477), .B(n11478), .Z(n6033) );
  IV U12367 ( .A(n11474), .Z(n11477) );
  XNOR U12368 ( .A(n6034), .B(n11474), .Z(n11476) );
  NAND U12369 ( .A(n11479), .B(e_input[137]), .Z(n6034) );
  NAND U12370 ( .A(n6112), .B(e_input[137]), .Z(n11479) );
  XOR U12371 ( .A(n11480), .B(n11481), .Z(n11474) );
  ANDN U12372 ( .A(n11482), .B(n6035), .Z(n11481) );
  XOR U12373 ( .A(n11483), .B(n11484), .Z(n6035) );
  IV U12374 ( .A(n11480), .Z(n11483) );
  XNOR U12375 ( .A(n6036), .B(n11480), .Z(n11482) );
  NAND U12376 ( .A(n11485), .B(e_input[136]), .Z(n6036) );
  NAND U12377 ( .A(n6112), .B(e_input[136]), .Z(n11485) );
  XOR U12378 ( .A(n11486), .B(n11487), .Z(n11480) );
  ANDN U12379 ( .A(n11488), .B(n6037), .Z(n11487) );
  XOR U12380 ( .A(n11489), .B(n11490), .Z(n6037) );
  IV U12381 ( .A(n11486), .Z(n11489) );
  XNOR U12382 ( .A(n6038), .B(n11486), .Z(n11488) );
  NAND U12383 ( .A(n11491), .B(e_input[135]), .Z(n6038) );
  NAND U12384 ( .A(n6112), .B(e_input[135]), .Z(n11491) );
  XOR U12385 ( .A(n11492), .B(n11493), .Z(n11486) );
  ANDN U12386 ( .A(n11494), .B(n6039), .Z(n11493) );
  XOR U12387 ( .A(n11495), .B(n11496), .Z(n6039) );
  IV U12388 ( .A(n11492), .Z(n11495) );
  XNOR U12389 ( .A(n6040), .B(n11492), .Z(n11494) );
  NAND U12390 ( .A(n11497), .B(e_input[134]), .Z(n6040) );
  NAND U12391 ( .A(n6112), .B(e_input[134]), .Z(n11497) );
  XOR U12392 ( .A(n11498), .B(n11499), .Z(n11492) );
  ANDN U12393 ( .A(n11500), .B(n6041), .Z(n11499) );
  XOR U12394 ( .A(n11501), .B(n11502), .Z(n6041) );
  IV U12395 ( .A(n11498), .Z(n11501) );
  XNOR U12396 ( .A(n6042), .B(n11498), .Z(n11500) );
  NAND U12397 ( .A(n11503), .B(e_input[133]), .Z(n6042) );
  NAND U12398 ( .A(n6112), .B(e_input[133]), .Z(n11503) );
  XOR U12399 ( .A(n11504), .B(n11505), .Z(n11498) );
  ANDN U12400 ( .A(n11506), .B(n6043), .Z(n11505) );
  XOR U12401 ( .A(n11507), .B(n11508), .Z(n6043) );
  IV U12402 ( .A(n11504), .Z(n11507) );
  XNOR U12403 ( .A(n6044), .B(n11504), .Z(n11506) );
  NAND U12404 ( .A(n11509), .B(e_input[132]), .Z(n6044) );
  NAND U12405 ( .A(n6112), .B(e_input[132]), .Z(n11509) );
  XOR U12406 ( .A(n11510), .B(n11511), .Z(n11504) );
  ANDN U12407 ( .A(n11512), .B(n6045), .Z(n11511) );
  XOR U12408 ( .A(n11513), .B(n11514), .Z(n6045) );
  IV U12409 ( .A(n11510), .Z(n11513) );
  XNOR U12410 ( .A(n6046), .B(n11510), .Z(n11512) );
  NAND U12411 ( .A(n11515), .B(e_input[131]), .Z(n6046) );
  NAND U12412 ( .A(n6112), .B(e_input[131]), .Z(n11515) );
  XOR U12413 ( .A(n11516), .B(n11517), .Z(n11510) );
  ANDN U12414 ( .A(n11518), .B(n6047), .Z(n11517) );
  XOR U12415 ( .A(n11519), .B(n11520), .Z(n6047) );
  IV U12416 ( .A(n11516), .Z(n11519) );
  XNOR U12417 ( .A(n6048), .B(n11516), .Z(n11518) );
  NAND U12418 ( .A(n11521), .B(e_input[130]), .Z(n6048) );
  NAND U12419 ( .A(n6112), .B(e_input[130]), .Z(n11521) );
  XOR U12420 ( .A(n11522), .B(n11523), .Z(n11516) );
  ANDN U12421 ( .A(n11524), .B(n6051), .Z(n11523) );
  XOR U12422 ( .A(n11525), .B(n11526), .Z(n6051) );
  IV U12423 ( .A(n11522), .Z(n11525) );
  XNOR U12424 ( .A(n6052), .B(n11522), .Z(n11524) );
  NAND U12425 ( .A(n11527), .B(e_input[129]), .Z(n6052) );
  NAND U12426 ( .A(n6112), .B(e_input[129]), .Z(n11527) );
  XOR U12427 ( .A(n11528), .B(n11529), .Z(n11522) );
  ANDN U12428 ( .A(n11530), .B(n6053), .Z(n11529) );
  XOR U12429 ( .A(n11531), .B(n11532), .Z(n6053) );
  IV U12430 ( .A(n11528), .Z(n11531) );
  XNOR U12431 ( .A(n6054), .B(n11528), .Z(n11530) );
  NAND U12432 ( .A(n11533), .B(e_input[128]), .Z(n6054) );
  NAND U12433 ( .A(n6112), .B(e_input[128]), .Z(n11533) );
  XOR U12434 ( .A(n11534), .B(n11535), .Z(n11528) );
  ANDN U12435 ( .A(n11536), .B(n6055), .Z(n11535) );
  XOR U12436 ( .A(n11537), .B(n11538), .Z(n6055) );
  IV U12437 ( .A(n11534), .Z(n11537) );
  XNOR U12438 ( .A(n6056), .B(n11534), .Z(n11536) );
  NAND U12439 ( .A(n11539), .B(e_input[127]), .Z(n6056) );
  NAND U12440 ( .A(n6112), .B(e_input[127]), .Z(n11539) );
  XOR U12441 ( .A(n11540), .B(n11541), .Z(n11534) );
  ANDN U12442 ( .A(n11542), .B(n6057), .Z(n11541) );
  XOR U12443 ( .A(n11543), .B(n11544), .Z(n6057) );
  IV U12444 ( .A(n11540), .Z(n11543) );
  XNOR U12445 ( .A(n6058), .B(n11540), .Z(n11542) );
  NAND U12446 ( .A(n11545), .B(e_input[126]), .Z(n6058) );
  NAND U12447 ( .A(n6112), .B(e_input[126]), .Z(n11545) );
  XOR U12448 ( .A(n11546), .B(n11547), .Z(n11540) );
  ANDN U12449 ( .A(n11548), .B(n6059), .Z(n11547) );
  XOR U12450 ( .A(n11549), .B(n11550), .Z(n6059) );
  IV U12451 ( .A(n11546), .Z(n11549) );
  XNOR U12452 ( .A(n6060), .B(n11546), .Z(n11548) );
  NAND U12453 ( .A(n11551), .B(e_input[125]), .Z(n6060) );
  NAND U12454 ( .A(n6112), .B(e_input[125]), .Z(n11551) );
  XOR U12455 ( .A(n11552), .B(n11553), .Z(n11546) );
  ANDN U12456 ( .A(n11554), .B(n6061), .Z(n11553) );
  XOR U12457 ( .A(n11555), .B(n11556), .Z(n6061) );
  IV U12458 ( .A(n11552), .Z(n11555) );
  XNOR U12459 ( .A(n6062), .B(n11552), .Z(n11554) );
  NAND U12460 ( .A(n11557), .B(e_input[124]), .Z(n6062) );
  NAND U12461 ( .A(n6112), .B(e_input[124]), .Z(n11557) );
  XOR U12462 ( .A(n11558), .B(n11559), .Z(n11552) );
  ANDN U12463 ( .A(n11560), .B(n6063), .Z(n11559) );
  XOR U12464 ( .A(n11561), .B(n11562), .Z(n6063) );
  IV U12465 ( .A(n11558), .Z(n11561) );
  XNOR U12466 ( .A(n6064), .B(n11558), .Z(n11560) );
  NAND U12467 ( .A(n11563), .B(e_input[123]), .Z(n6064) );
  NAND U12468 ( .A(n6112), .B(e_input[123]), .Z(n11563) );
  XOR U12469 ( .A(n11564), .B(n11565), .Z(n11558) );
  ANDN U12470 ( .A(n11566), .B(n6065), .Z(n11565) );
  XOR U12471 ( .A(n11567), .B(n11568), .Z(n6065) );
  IV U12472 ( .A(n11564), .Z(n11567) );
  XNOR U12473 ( .A(n6066), .B(n11564), .Z(n11566) );
  NAND U12474 ( .A(n11569), .B(e_input[122]), .Z(n6066) );
  NAND U12475 ( .A(n6112), .B(e_input[122]), .Z(n11569) );
  XOR U12476 ( .A(n11570), .B(n11571), .Z(n11564) );
  ANDN U12477 ( .A(n11572), .B(n6067), .Z(n11571) );
  XOR U12478 ( .A(n11573), .B(n11574), .Z(n6067) );
  IV U12479 ( .A(n11570), .Z(n11573) );
  XNOR U12480 ( .A(n6068), .B(n11570), .Z(n11572) );
  NAND U12481 ( .A(n11575), .B(e_input[121]), .Z(n6068) );
  NAND U12482 ( .A(n6112), .B(e_input[121]), .Z(n11575) );
  XOR U12483 ( .A(n11576), .B(n11577), .Z(n11570) );
  ANDN U12484 ( .A(n11578), .B(n6069), .Z(n11577) );
  XOR U12485 ( .A(n11579), .B(n11580), .Z(n6069) );
  IV U12486 ( .A(n11576), .Z(n11579) );
  XNOR U12487 ( .A(n6070), .B(n11576), .Z(n11578) );
  NAND U12488 ( .A(n11581), .B(e_input[120]), .Z(n6070) );
  NAND U12489 ( .A(n6112), .B(e_input[120]), .Z(n11581) );
  XOR U12490 ( .A(n11582), .B(n11583), .Z(n11576) );
  ANDN U12491 ( .A(n11584), .B(n6073), .Z(n11583) );
  XOR U12492 ( .A(n11585), .B(n11586), .Z(n6073) );
  IV U12493 ( .A(n11582), .Z(n11585) );
  XNOR U12494 ( .A(n6074), .B(n11582), .Z(n11584) );
  NAND U12495 ( .A(n11587), .B(e_input[119]), .Z(n6074) );
  NAND U12496 ( .A(n6112), .B(e_input[119]), .Z(n11587) );
  XOR U12497 ( .A(n11588), .B(n11589), .Z(n11582) );
  ANDN U12498 ( .A(n11590), .B(n6075), .Z(n11589) );
  XOR U12499 ( .A(n11591), .B(n11592), .Z(n6075) );
  IV U12500 ( .A(n11588), .Z(n11591) );
  XNOR U12501 ( .A(n6076), .B(n11588), .Z(n11590) );
  NAND U12502 ( .A(n11593), .B(e_input[118]), .Z(n6076) );
  NAND U12503 ( .A(n6112), .B(e_input[118]), .Z(n11593) );
  XOR U12504 ( .A(n11594), .B(n11595), .Z(n11588) );
  ANDN U12505 ( .A(n11596), .B(n6077), .Z(n11595) );
  XOR U12506 ( .A(n11597), .B(n11598), .Z(n6077) );
  IV U12507 ( .A(n11594), .Z(n11597) );
  XNOR U12508 ( .A(n6078), .B(n11594), .Z(n11596) );
  NAND U12509 ( .A(n11599), .B(e_input[117]), .Z(n6078) );
  NAND U12510 ( .A(n6112), .B(e_input[117]), .Z(n11599) );
  XOR U12511 ( .A(n11600), .B(n11601), .Z(n11594) );
  ANDN U12512 ( .A(n11602), .B(n6079), .Z(n11601) );
  XOR U12513 ( .A(n11603), .B(n11604), .Z(n6079) );
  IV U12514 ( .A(n11600), .Z(n11603) );
  XNOR U12515 ( .A(n6080), .B(n11600), .Z(n11602) );
  NAND U12516 ( .A(n11605), .B(e_input[116]), .Z(n6080) );
  NAND U12517 ( .A(n6112), .B(e_input[116]), .Z(n11605) );
  XOR U12518 ( .A(n11606), .B(n11607), .Z(n11600) );
  ANDN U12519 ( .A(n11608), .B(n6081), .Z(n11607) );
  XOR U12520 ( .A(n11609), .B(n11610), .Z(n6081) );
  IV U12521 ( .A(n11606), .Z(n11609) );
  XNOR U12522 ( .A(n6082), .B(n11606), .Z(n11608) );
  NAND U12523 ( .A(n11611), .B(e_input[115]), .Z(n6082) );
  NAND U12524 ( .A(n6112), .B(e_input[115]), .Z(n11611) );
  XOR U12525 ( .A(n11612), .B(n11613), .Z(n11606) );
  ANDN U12526 ( .A(n11614), .B(n6083), .Z(n11613) );
  XOR U12527 ( .A(n11615), .B(n11616), .Z(n6083) );
  IV U12528 ( .A(n11612), .Z(n11615) );
  XNOR U12529 ( .A(n6084), .B(n11612), .Z(n11614) );
  NAND U12530 ( .A(n11617), .B(e_input[114]), .Z(n6084) );
  NAND U12531 ( .A(n6112), .B(e_input[114]), .Z(n11617) );
  XOR U12532 ( .A(n11618), .B(n11619), .Z(n11612) );
  ANDN U12533 ( .A(n11620), .B(n6085), .Z(n11619) );
  XOR U12534 ( .A(n11621), .B(n11622), .Z(n6085) );
  IV U12535 ( .A(n11618), .Z(n11621) );
  XNOR U12536 ( .A(n6086), .B(n11618), .Z(n11620) );
  NAND U12537 ( .A(n11623), .B(e_input[113]), .Z(n6086) );
  NAND U12538 ( .A(n6112), .B(e_input[113]), .Z(n11623) );
  XOR U12539 ( .A(n11624), .B(n11625), .Z(n11618) );
  ANDN U12540 ( .A(n11626), .B(n6087), .Z(n11625) );
  XOR U12541 ( .A(n11627), .B(n11628), .Z(n6087) );
  IV U12542 ( .A(n11624), .Z(n11627) );
  XNOR U12543 ( .A(n6088), .B(n11624), .Z(n11626) );
  NAND U12544 ( .A(n11629), .B(e_input[112]), .Z(n6088) );
  NAND U12545 ( .A(n6112), .B(e_input[112]), .Z(n11629) );
  XOR U12546 ( .A(n11630), .B(n11631), .Z(n11624) );
  ANDN U12547 ( .A(n11632), .B(n6089), .Z(n11631) );
  XOR U12548 ( .A(n11633), .B(n11634), .Z(n6089) );
  IV U12549 ( .A(n11630), .Z(n11633) );
  XNOR U12550 ( .A(n6090), .B(n11630), .Z(n11632) );
  NAND U12551 ( .A(n11635), .B(e_input[111]), .Z(n6090) );
  NAND U12552 ( .A(n6112), .B(e_input[111]), .Z(n11635) );
  XOR U12553 ( .A(n11636), .B(n11637), .Z(n11630) );
  ANDN U12554 ( .A(n11638), .B(n6091), .Z(n11637) );
  XOR U12555 ( .A(n11639), .B(n11640), .Z(n6091) );
  IV U12556 ( .A(n11636), .Z(n11639) );
  XNOR U12557 ( .A(n6092), .B(n11636), .Z(n11638) );
  NAND U12558 ( .A(n11641), .B(e_input[110]), .Z(n6092) );
  NAND U12559 ( .A(n6112), .B(e_input[110]), .Z(n11641) );
  XOR U12560 ( .A(n11642), .B(n11643), .Z(n11636) );
  ANDN U12561 ( .A(n11644), .B(n6095), .Z(n11643) );
  XOR U12562 ( .A(n11645), .B(n11646), .Z(n6095) );
  IV U12563 ( .A(n11642), .Z(n11645) );
  XNOR U12564 ( .A(n6096), .B(n11642), .Z(n11644) );
  NAND U12565 ( .A(n11647), .B(e_input[109]), .Z(n6096) );
  NAND U12566 ( .A(n6112), .B(e_input[109]), .Z(n11647) );
  XOR U12567 ( .A(n11648), .B(n11649), .Z(n11642) );
  ANDN U12568 ( .A(n11650), .B(n6097), .Z(n11649) );
  XOR U12569 ( .A(n11651), .B(n11652), .Z(n6097) );
  IV U12570 ( .A(n11648), .Z(n11651) );
  XNOR U12571 ( .A(n6098), .B(n11648), .Z(n11650) );
  NAND U12572 ( .A(n11653), .B(e_input[108]), .Z(n6098) );
  NAND U12573 ( .A(n6112), .B(e_input[108]), .Z(n11653) );
  XOR U12574 ( .A(n11654), .B(n11655), .Z(n11648) );
  ANDN U12575 ( .A(n11656), .B(n6099), .Z(n11655) );
  XOR U12576 ( .A(n11657), .B(n11658), .Z(n6099) );
  IV U12577 ( .A(n11654), .Z(n11657) );
  XNOR U12578 ( .A(n6100), .B(n11654), .Z(n11656) );
  NAND U12579 ( .A(n11659), .B(e_input[107]), .Z(n6100) );
  NAND U12580 ( .A(n6112), .B(e_input[107]), .Z(n11659) );
  XOR U12581 ( .A(n11660), .B(n11661), .Z(n11654) );
  ANDN U12582 ( .A(n11662), .B(n6101), .Z(n11661) );
  XOR U12583 ( .A(n11663), .B(n11664), .Z(n6101) );
  IV U12584 ( .A(n11660), .Z(n11663) );
  XNOR U12585 ( .A(n6102), .B(n11660), .Z(n11662) );
  NAND U12586 ( .A(n11665), .B(e_input[106]), .Z(n6102) );
  NAND U12587 ( .A(n6112), .B(e_input[106]), .Z(n11665) );
  XOR U12588 ( .A(n11666), .B(n11667), .Z(n11660) );
  ANDN U12589 ( .A(n11668), .B(n6103), .Z(n11667) );
  XOR U12590 ( .A(n11669), .B(n11670), .Z(n6103) );
  IV U12591 ( .A(n11666), .Z(n11669) );
  XNOR U12592 ( .A(n6104), .B(n11666), .Z(n11668) );
  NAND U12593 ( .A(n11671), .B(e_input[105]), .Z(n6104) );
  NAND U12594 ( .A(n6112), .B(e_input[105]), .Z(n11671) );
  XOR U12595 ( .A(n11672), .B(n11673), .Z(n11666) );
  ANDN U12596 ( .A(n11674), .B(n6105), .Z(n11673) );
  XOR U12597 ( .A(n11675), .B(n11676), .Z(n6105) );
  IV U12598 ( .A(n11672), .Z(n11675) );
  XNOR U12599 ( .A(n6106), .B(n11672), .Z(n11674) );
  NAND U12600 ( .A(n11677), .B(e_input[104]), .Z(n6106) );
  NAND U12601 ( .A(n6112), .B(e_input[104]), .Z(n11677) );
  XOR U12602 ( .A(n11678), .B(n11679), .Z(n11672) );
  ANDN U12603 ( .A(n11680), .B(n6107), .Z(n11679) );
  XOR U12604 ( .A(n11681), .B(n11682), .Z(n6107) );
  IV U12605 ( .A(n11678), .Z(n11681) );
  XNOR U12606 ( .A(n6108), .B(n11678), .Z(n11680) );
  NAND U12607 ( .A(n11683), .B(e_input[103]), .Z(n6108) );
  NAND U12608 ( .A(n6112), .B(e_input[103]), .Z(n11683) );
  XOR U12609 ( .A(n11684), .B(n11685), .Z(n11678) );
  ANDN U12610 ( .A(n11686), .B(n6109), .Z(n11685) );
  XOR U12611 ( .A(n11687), .B(n11688), .Z(n6109) );
  IV U12612 ( .A(n11684), .Z(n11687) );
  XNOR U12613 ( .A(n6110), .B(n11684), .Z(n11686) );
  NAND U12614 ( .A(n11689), .B(e_input[102]), .Z(n6110) );
  NAND U12615 ( .A(n6112), .B(e_input[102]), .Z(n11689) );
  XOR U12616 ( .A(n11690), .B(n11691), .Z(n11684) );
  ANDN U12617 ( .A(n11692), .B(n6143), .Z(n11691) );
  XOR U12618 ( .A(n11693), .B(n11694), .Z(n6143) );
  IV U12619 ( .A(n11690), .Z(n11693) );
  XNOR U12620 ( .A(n6144), .B(n11690), .Z(n11692) );
  NAND U12621 ( .A(n11695), .B(e_input[101]), .Z(n6144) );
  NAND U12622 ( .A(n6112), .B(e_input[101]), .Z(n11695) );
  XOR U12623 ( .A(n11696), .B(n11697), .Z(n11690) );
  ANDN U12624 ( .A(n11698), .B(n6225), .Z(n11697) );
  XOR U12625 ( .A(n11699), .B(n11700), .Z(n6225) );
  IV U12626 ( .A(n11696), .Z(n11699) );
  XNOR U12627 ( .A(n6226), .B(n11696), .Z(n11698) );
  NAND U12628 ( .A(n11701), .B(e_input[100]), .Z(n6226) );
  NAND U12629 ( .A(n6112), .B(e_input[100]), .Z(n11701) );
  XOR U12630 ( .A(n11702), .B(n11703), .Z(n11696) );
  ANDN U12631 ( .A(n11704), .B(n4119), .Z(n11703) );
  XOR U12632 ( .A(n11705), .B(n11706), .Z(n4119) );
  IV U12633 ( .A(n11702), .Z(n11705) );
  XNOR U12634 ( .A(n4120), .B(n11702), .Z(n11704) );
  NAND U12635 ( .A(n11707), .B(e_input[99]), .Z(n4120) );
  NAND U12636 ( .A(n6112), .B(e_input[99]), .Z(n11707) );
  XOR U12637 ( .A(n11708), .B(n11709), .Z(n11702) );
  ANDN U12638 ( .A(n11710), .B(n4141), .Z(n11709) );
  XOR U12639 ( .A(n11711), .B(n11712), .Z(n4141) );
  IV U12640 ( .A(n11708), .Z(n11711) );
  XNOR U12641 ( .A(n4142), .B(n11708), .Z(n11710) );
  NAND U12642 ( .A(n11713), .B(e_input[98]), .Z(n4142) );
  NAND U12643 ( .A(n6112), .B(e_input[98]), .Z(n11713) );
  XOR U12644 ( .A(n11714), .B(n11715), .Z(n11708) );
  ANDN U12645 ( .A(n11716), .B(n4163), .Z(n11715) );
  XOR U12646 ( .A(n11717), .B(n11718), .Z(n4163) );
  IV U12647 ( .A(n11714), .Z(n11717) );
  XNOR U12648 ( .A(n4164), .B(n11714), .Z(n11716) );
  NAND U12649 ( .A(n11719), .B(e_input[97]), .Z(n4164) );
  NAND U12650 ( .A(n6112), .B(e_input[97]), .Z(n11719) );
  XOR U12651 ( .A(n11720), .B(n11721), .Z(n11714) );
  ANDN U12652 ( .A(n11722), .B(n4185), .Z(n11721) );
  XOR U12653 ( .A(n11723), .B(n11724), .Z(n4185) );
  IV U12654 ( .A(n11720), .Z(n11723) );
  XNOR U12655 ( .A(n4186), .B(n11720), .Z(n11722) );
  NAND U12656 ( .A(n11725), .B(e_input[96]), .Z(n4186) );
  NAND U12657 ( .A(n6112), .B(e_input[96]), .Z(n11725) );
  XOR U12658 ( .A(n11726), .B(n11727), .Z(n11720) );
  ANDN U12659 ( .A(n11728), .B(n4207), .Z(n11727) );
  XOR U12660 ( .A(n11729), .B(n11730), .Z(n4207) );
  IV U12661 ( .A(n11726), .Z(n11729) );
  XNOR U12662 ( .A(n4208), .B(n11726), .Z(n11728) );
  NAND U12663 ( .A(n11731), .B(e_input[95]), .Z(n4208) );
  NAND U12664 ( .A(n6112), .B(e_input[95]), .Z(n11731) );
  XOR U12665 ( .A(n11732), .B(n11733), .Z(n11726) );
  ANDN U12666 ( .A(n11734), .B(n4229), .Z(n11733) );
  XOR U12667 ( .A(n11735), .B(n11736), .Z(n4229) );
  IV U12668 ( .A(n11732), .Z(n11735) );
  XNOR U12669 ( .A(n4230), .B(n11732), .Z(n11734) );
  NAND U12670 ( .A(n11737), .B(e_input[94]), .Z(n4230) );
  NAND U12671 ( .A(n6112), .B(e_input[94]), .Z(n11737) );
  XOR U12672 ( .A(n11738), .B(n11739), .Z(n11732) );
  ANDN U12673 ( .A(n11740), .B(n4251), .Z(n11739) );
  XOR U12674 ( .A(n11741), .B(n11742), .Z(n4251) );
  IV U12675 ( .A(n11738), .Z(n11741) );
  XNOR U12676 ( .A(n4252), .B(n11738), .Z(n11740) );
  NAND U12677 ( .A(n11743), .B(e_input[93]), .Z(n4252) );
  NAND U12678 ( .A(n6112), .B(e_input[93]), .Z(n11743) );
  XOR U12679 ( .A(n11744), .B(n11745), .Z(n11738) );
  ANDN U12680 ( .A(n11746), .B(n4273), .Z(n11745) );
  XOR U12681 ( .A(n11747), .B(n11748), .Z(n4273) );
  IV U12682 ( .A(n11744), .Z(n11747) );
  XNOR U12683 ( .A(n4274), .B(n11744), .Z(n11746) );
  NAND U12684 ( .A(n11749), .B(e_input[92]), .Z(n4274) );
  NAND U12685 ( .A(n6112), .B(e_input[92]), .Z(n11749) );
  XOR U12686 ( .A(n11750), .B(n11751), .Z(n11744) );
  ANDN U12687 ( .A(n11752), .B(n4295), .Z(n11751) );
  XOR U12688 ( .A(n11753), .B(n11754), .Z(n4295) );
  IV U12689 ( .A(n11750), .Z(n11753) );
  XNOR U12690 ( .A(n4296), .B(n11750), .Z(n11752) );
  NAND U12691 ( .A(n11755), .B(e_input[91]), .Z(n4296) );
  NAND U12692 ( .A(n6112), .B(e_input[91]), .Z(n11755) );
  XOR U12693 ( .A(n11756), .B(n11757), .Z(n11750) );
  ANDN U12694 ( .A(n11758), .B(n4317), .Z(n11757) );
  XOR U12695 ( .A(n11759), .B(n11760), .Z(n4317) );
  IV U12696 ( .A(n11756), .Z(n11759) );
  XNOR U12697 ( .A(n4318), .B(n11756), .Z(n11758) );
  NAND U12698 ( .A(n11761), .B(e_input[90]), .Z(n4318) );
  NAND U12699 ( .A(n6112), .B(e_input[90]), .Z(n11761) );
  XOR U12700 ( .A(n11762), .B(n11763), .Z(n11756) );
  ANDN U12701 ( .A(n11764), .B(n4341), .Z(n11763) );
  XOR U12702 ( .A(n11765), .B(n11766), .Z(n4341) );
  IV U12703 ( .A(n11762), .Z(n11765) );
  XNOR U12704 ( .A(n4342), .B(n11762), .Z(n11764) );
  NAND U12705 ( .A(n11767), .B(e_input[89]), .Z(n4342) );
  NAND U12706 ( .A(n6112), .B(e_input[89]), .Z(n11767) );
  XOR U12707 ( .A(n11768), .B(n11769), .Z(n11762) );
  ANDN U12708 ( .A(n11770), .B(n4363), .Z(n11769) );
  XOR U12709 ( .A(n11771), .B(n11772), .Z(n4363) );
  IV U12710 ( .A(n11768), .Z(n11771) );
  XNOR U12711 ( .A(n4364), .B(n11768), .Z(n11770) );
  NAND U12712 ( .A(n11773), .B(e_input[88]), .Z(n4364) );
  NAND U12713 ( .A(n6112), .B(e_input[88]), .Z(n11773) );
  XOR U12714 ( .A(n11774), .B(n11775), .Z(n11768) );
  ANDN U12715 ( .A(n11776), .B(n4385), .Z(n11775) );
  XOR U12716 ( .A(n11777), .B(n11778), .Z(n4385) );
  IV U12717 ( .A(n11774), .Z(n11777) );
  XNOR U12718 ( .A(n4386), .B(n11774), .Z(n11776) );
  NAND U12719 ( .A(n11779), .B(e_input[87]), .Z(n4386) );
  NAND U12720 ( .A(n6112), .B(e_input[87]), .Z(n11779) );
  XOR U12721 ( .A(n11780), .B(n11781), .Z(n11774) );
  ANDN U12722 ( .A(n11782), .B(n4407), .Z(n11781) );
  XOR U12723 ( .A(n11783), .B(n11784), .Z(n4407) );
  IV U12724 ( .A(n11780), .Z(n11783) );
  XNOR U12725 ( .A(n4408), .B(n11780), .Z(n11782) );
  NAND U12726 ( .A(n11785), .B(e_input[86]), .Z(n4408) );
  NAND U12727 ( .A(n6112), .B(e_input[86]), .Z(n11785) );
  XOR U12728 ( .A(n11786), .B(n11787), .Z(n11780) );
  ANDN U12729 ( .A(n11788), .B(n4429), .Z(n11787) );
  XOR U12730 ( .A(n11789), .B(n11790), .Z(n4429) );
  IV U12731 ( .A(n11786), .Z(n11789) );
  XNOR U12732 ( .A(n4430), .B(n11786), .Z(n11788) );
  NAND U12733 ( .A(n11791), .B(e_input[85]), .Z(n4430) );
  NAND U12734 ( .A(n6112), .B(e_input[85]), .Z(n11791) );
  XOR U12735 ( .A(n11792), .B(n11793), .Z(n11786) );
  ANDN U12736 ( .A(n11794), .B(n4451), .Z(n11793) );
  XOR U12737 ( .A(n11795), .B(n11796), .Z(n4451) );
  IV U12738 ( .A(n11792), .Z(n11795) );
  XNOR U12739 ( .A(n4452), .B(n11792), .Z(n11794) );
  NAND U12740 ( .A(n11797), .B(e_input[84]), .Z(n4452) );
  NAND U12741 ( .A(n6112), .B(e_input[84]), .Z(n11797) );
  XOR U12742 ( .A(n11798), .B(n11799), .Z(n11792) );
  ANDN U12743 ( .A(n11800), .B(n4473), .Z(n11799) );
  XOR U12744 ( .A(n11801), .B(n11802), .Z(n4473) );
  IV U12745 ( .A(n11798), .Z(n11801) );
  XNOR U12746 ( .A(n4474), .B(n11798), .Z(n11800) );
  NAND U12747 ( .A(n11803), .B(e_input[83]), .Z(n4474) );
  NAND U12748 ( .A(n6112), .B(e_input[83]), .Z(n11803) );
  XOR U12749 ( .A(n11804), .B(n11805), .Z(n11798) );
  ANDN U12750 ( .A(n11806), .B(n4495), .Z(n11805) );
  XOR U12751 ( .A(n11807), .B(n11808), .Z(n4495) );
  IV U12752 ( .A(n11804), .Z(n11807) );
  XNOR U12753 ( .A(n4496), .B(n11804), .Z(n11806) );
  NAND U12754 ( .A(n11809), .B(e_input[82]), .Z(n4496) );
  NAND U12755 ( .A(n6112), .B(e_input[82]), .Z(n11809) );
  XOR U12756 ( .A(n11810), .B(n11811), .Z(n11804) );
  ANDN U12757 ( .A(n11812), .B(n4517), .Z(n11811) );
  XOR U12758 ( .A(n11813), .B(n11814), .Z(n4517) );
  IV U12759 ( .A(n11810), .Z(n11813) );
  XNOR U12760 ( .A(n4518), .B(n11810), .Z(n11812) );
  NAND U12761 ( .A(n11815), .B(e_input[81]), .Z(n4518) );
  NAND U12762 ( .A(n6112), .B(e_input[81]), .Z(n11815) );
  XOR U12763 ( .A(n11816), .B(n11817), .Z(n11810) );
  ANDN U12764 ( .A(n11818), .B(n4539), .Z(n11817) );
  XOR U12765 ( .A(n11819), .B(n11820), .Z(n4539) );
  IV U12766 ( .A(n11816), .Z(n11819) );
  XNOR U12767 ( .A(n4540), .B(n11816), .Z(n11818) );
  NAND U12768 ( .A(n11821), .B(e_input[80]), .Z(n4540) );
  NAND U12769 ( .A(n6112), .B(e_input[80]), .Z(n11821) );
  XOR U12770 ( .A(n11822), .B(n11823), .Z(n11816) );
  ANDN U12771 ( .A(n11824), .B(n4563), .Z(n11823) );
  XOR U12772 ( .A(n11825), .B(n11826), .Z(n4563) );
  IV U12773 ( .A(n11822), .Z(n11825) );
  XNOR U12774 ( .A(n4564), .B(n11822), .Z(n11824) );
  NAND U12775 ( .A(n11827), .B(e_input[79]), .Z(n4564) );
  NAND U12776 ( .A(n6112), .B(e_input[79]), .Z(n11827) );
  XOR U12777 ( .A(n11828), .B(n11829), .Z(n11822) );
  ANDN U12778 ( .A(n11830), .B(n4585), .Z(n11829) );
  XOR U12779 ( .A(n11831), .B(n11832), .Z(n4585) );
  IV U12780 ( .A(n11828), .Z(n11831) );
  XNOR U12781 ( .A(n4586), .B(n11828), .Z(n11830) );
  NAND U12782 ( .A(n11833), .B(e_input[78]), .Z(n4586) );
  NAND U12783 ( .A(n6112), .B(e_input[78]), .Z(n11833) );
  XOR U12784 ( .A(n11834), .B(n11835), .Z(n11828) );
  ANDN U12785 ( .A(n11836), .B(n4607), .Z(n11835) );
  XOR U12786 ( .A(n11837), .B(n11838), .Z(n4607) );
  IV U12787 ( .A(n11834), .Z(n11837) );
  XNOR U12788 ( .A(n4608), .B(n11834), .Z(n11836) );
  NAND U12789 ( .A(n11839), .B(e_input[77]), .Z(n4608) );
  NAND U12790 ( .A(n6112), .B(e_input[77]), .Z(n11839) );
  XOR U12791 ( .A(n11840), .B(n11841), .Z(n11834) );
  ANDN U12792 ( .A(n11842), .B(n4629), .Z(n11841) );
  XOR U12793 ( .A(n11843), .B(n11844), .Z(n4629) );
  IV U12794 ( .A(n11840), .Z(n11843) );
  XNOR U12795 ( .A(n4630), .B(n11840), .Z(n11842) );
  NAND U12796 ( .A(n11845), .B(e_input[76]), .Z(n4630) );
  NAND U12797 ( .A(n6112), .B(e_input[76]), .Z(n11845) );
  XOR U12798 ( .A(n11846), .B(n11847), .Z(n11840) );
  ANDN U12799 ( .A(n11848), .B(n4651), .Z(n11847) );
  XOR U12800 ( .A(n11849), .B(n11850), .Z(n4651) );
  IV U12801 ( .A(n11846), .Z(n11849) );
  XNOR U12802 ( .A(n4652), .B(n11846), .Z(n11848) );
  NAND U12803 ( .A(n11851), .B(e_input[75]), .Z(n4652) );
  NAND U12804 ( .A(n6112), .B(e_input[75]), .Z(n11851) );
  XOR U12805 ( .A(n11852), .B(n11853), .Z(n11846) );
  ANDN U12806 ( .A(n11854), .B(n4673), .Z(n11853) );
  XOR U12807 ( .A(n11855), .B(n11856), .Z(n4673) );
  IV U12808 ( .A(n11852), .Z(n11855) );
  XNOR U12809 ( .A(n4674), .B(n11852), .Z(n11854) );
  NAND U12810 ( .A(n11857), .B(e_input[74]), .Z(n4674) );
  NAND U12811 ( .A(n6112), .B(e_input[74]), .Z(n11857) );
  XOR U12812 ( .A(n11858), .B(n11859), .Z(n11852) );
  ANDN U12813 ( .A(n11860), .B(n4695), .Z(n11859) );
  XOR U12814 ( .A(n11861), .B(n11862), .Z(n4695) );
  IV U12815 ( .A(n11858), .Z(n11861) );
  XNOR U12816 ( .A(n4696), .B(n11858), .Z(n11860) );
  NAND U12817 ( .A(n11863), .B(e_input[73]), .Z(n4696) );
  NAND U12818 ( .A(n6112), .B(e_input[73]), .Z(n11863) );
  XOR U12819 ( .A(n11864), .B(n11865), .Z(n11858) );
  ANDN U12820 ( .A(n11866), .B(n4717), .Z(n11865) );
  XOR U12821 ( .A(n11867), .B(n11868), .Z(n4717) );
  IV U12822 ( .A(n11864), .Z(n11867) );
  XNOR U12823 ( .A(n4718), .B(n11864), .Z(n11866) );
  NAND U12824 ( .A(n11869), .B(e_input[72]), .Z(n4718) );
  NAND U12825 ( .A(n6112), .B(e_input[72]), .Z(n11869) );
  XOR U12826 ( .A(n11870), .B(n11871), .Z(n11864) );
  ANDN U12827 ( .A(n11872), .B(n4739), .Z(n11871) );
  XOR U12828 ( .A(n11873), .B(n11874), .Z(n4739) );
  IV U12829 ( .A(n11870), .Z(n11873) );
  XNOR U12830 ( .A(n4740), .B(n11870), .Z(n11872) );
  NAND U12831 ( .A(n11875), .B(e_input[71]), .Z(n4740) );
  NAND U12832 ( .A(n6112), .B(e_input[71]), .Z(n11875) );
  XOR U12833 ( .A(n11876), .B(n11877), .Z(n11870) );
  ANDN U12834 ( .A(n11878), .B(n4761), .Z(n11877) );
  XOR U12835 ( .A(n11879), .B(n11880), .Z(n4761) );
  IV U12836 ( .A(n11876), .Z(n11879) );
  XNOR U12837 ( .A(n4762), .B(n11876), .Z(n11878) );
  NAND U12838 ( .A(n11881), .B(e_input[70]), .Z(n4762) );
  NAND U12839 ( .A(n6112), .B(e_input[70]), .Z(n11881) );
  XOR U12840 ( .A(n11882), .B(n11883), .Z(n11876) );
  ANDN U12841 ( .A(n11884), .B(n4785), .Z(n11883) );
  XOR U12842 ( .A(n11885), .B(n11886), .Z(n4785) );
  IV U12843 ( .A(n11882), .Z(n11885) );
  XNOR U12844 ( .A(n4786), .B(n11882), .Z(n11884) );
  NAND U12845 ( .A(n11887), .B(e_input[69]), .Z(n4786) );
  NAND U12846 ( .A(n6112), .B(e_input[69]), .Z(n11887) );
  XOR U12847 ( .A(n11888), .B(n11889), .Z(n11882) );
  ANDN U12848 ( .A(n11890), .B(n4807), .Z(n11889) );
  XOR U12849 ( .A(n11891), .B(n11892), .Z(n4807) );
  IV U12850 ( .A(n11888), .Z(n11891) );
  XNOR U12851 ( .A(n4808), .B(n11888), .Z(n11890) );
  NAND U12852 ( .A(n11893), .B(e_input[68]), .Z(n4808) );
  NAND U12853 ( .A(n6112), .B(e_input[68]), .Z(n11893) );
  XOR U12854 ( .A(n11894), .B(n11895), .Z(n11888) );
  ANDN U12855 ( .A(n11896), .B(n4829), .Z(n11895) );
  XOR U12856 ( .A(n11897), .B(n11898), .Z(n4829) );
  IV U12857 ( .A(n11894), .Z(n11897) );
  XNOR U12858 ( .A(n4830), .B(n11894), .Z(n11896) );
  NAND U12859 ( .A(n11899), .B(e_input[67]), .Z(n4830) );
  NAND U12860 ( .A(n6112), .B(e_input[67]), .Z(n11899) );
  XOR U12861 ( .A(n11900), .B(n11901), .Z(n11894) );
  ANDN U12862 ( .A(n11902), .B(n4851), .Z(n11901) );
  XOR U12863 ( .A(n11903), .B(n11904), .Z(n4851) );
  IV U12864 ( .A(n11900), .Z(n11903) );
  XNOR U12865 ( .A(n4852), .B(n11900), .Z(n11902) );
  NAND U12866 ( .A(n11905), .B(e_input[66]), .Z(n4852) );
  NAND U12867 ( .A(n6112), .B(e_input[66]), .Z(n11905) );
  XOR U12868 ( .A(n11906), .B(n11907), .Z(n11900) );
  ANDN U12869 ( .A(n11908), .B(n4873), .Z(n11907) );
  XOR U12870 ( .A(n11909), .B(n11910), .Z(n4873) );
  IV U12871 ( .A(n11906), .Z(n11909) );
  XNOR U12872 ( .A(n4874), .B(n11906), .Z(n11908) );
  NAND U12873 ( .A(n11911), .B(e_input[65]), .Z(n4874) );
  NAND U12874 ( .A(n6112), .B(e_input[65]), .Z(n11911) );
  XOR U12875 ( .A(n11912), .B(n11913), .Z(n11906) );
  ANDN U12876 ( .A(n11914), .B(n4895), .Z(n11913) );
  XOR U12877 ( .A(n11915), .B(n11916), .Z(n4895) );
  IV U12878 ( .A(n11912), .Z(n11915) );
  XNOR U12879 ( .A(n4896), .B(n11912), .Z(n11914) );
  NAND U12880 ( .A(n11917), .B(e_input[64]), .Z(n4896) );
  NAND U12881 ( .A(n6112), .B(e_input[64]), .Z(n11917) );
  XOR U12882 ( .A(n11918), .B(n11919), .Z(n11912) );
  ANDN U12883 ( .A(n11920), .B(n4917), .Z(n11919) );
  XOR U12884 ( .A(n11921), .B(n11922), .Z(n4917) );
  IV U12885 ( .A(n11918), .Z(n11921) );
  XNOR U12886 ( .A(n4918), .B(n11918), .Z(n11920) );
  NAND U12887 ( .A(n11923), .B(e_input[63]), .Z(n4918) );
  NAND U12888 ( .A(n6112), .B(e_input[63]), .Z(n11923) );
  XOR U12889 ( .A(n11924), .B(n11925), .Z(n11918) );
  ANDN U12890 ( .A(n11926), .B(n4939), .Z(n11925) );
  XOR U12891 ( .A(n11927), .B(n11928), .Z(n4939) );
  IV U12892 ( .A(n11924), .Z(n11927) );
  XNOR U12893 ( .A(n4940), .B(n11924), .Z(n11926) );
  NAND U12894 ( .A(n11929), .B(e_input[62]), .Z(n4940) );
  NAND U12895 ( .A(n6112), .B(e_input[62]), .Z(n11929) );
  XOR U12896 ( .A(n11930), .B(n11931), .Z(n11924) );
  ANDN U12897 ( .A(n11932), .B(n4961), .Z(n11931) );
  XOR U12898 ( .A(n11933), .B(n11934), .Z(n4961) );
  IV U12899 ( .A(n11930), .Z(n11933) );
  XNOR U12900 ( .A(n4962), .B(n11930), .Z(n11932) );
  NAND U12901 ( .A(n11935), .B(e_input[61]), .Z(n4962) );
  NAND U12902 ( .A(n6112), .B(e_input[61]), .Z(n11935) );
  XOR U12903 ( .A(n11936), .B(n11937), .Z(n11930) );
  ANDN U12904 ( .A(n11938), .B(n4983), .Z(n11937) );
  XOR U12905 ( .A(n11939), .B(n11940), .Z(n4983) );
  IV U12906 ( .A(n11936), .Z(n11939) );
  XNOR U12907 ( .A(n4984), .B(n11936), .Z(n11938) );
  NAND U12908 ( .A(n11941), .B(e_input[60]), .Z(n4984) );
  NAND U12909 ( .A(n6112), .B(e_input[60]), .Z(n11941) );
  XOR U12910 ( .A(n11942), .B(n11943), .Z(n11936) );
  ANDN U12911 ( .A(n11944), .B(n5007), .Z(n11943) );
  XOR U12912 ( .A(n11945), .B(n11946), .Z(n5007) );
  IV U12913 ( .A(n11942), .Z(n11945) );
  XNOR U12914 ( .A(n5008), .B(n11942), .Z(n11944) );
  NAND U12915 ( .A(n11947), .B(e_input[59]), .Z(n5008) );
  NAND U12916 ( .A(n6112), .B(e_input[59]), .Z(n11947) );
  XOR U12917 ( .A(n11948), .B(n11949), .Z(n11942) );
  ANDN U12918 ( .A(n11950), .B(n5029), .Z(n11949) );
  XOR U12919 ( .A(n11951), .B(n11952), .Z(n5029) );
  IV U12920 ( .A(n11948), .Z(n11951) );
  XNOR U12921 ( .A(n5030), .B(n11948), .Z(n11950) );
  NAND U12922 ( .A(n11953), .B(e_input[58]), .Z(n5030) );
  NAND U12923 ( .A(n6112), .B(e_input[58]), .Z(n11953) );
  XOR U12924 ( .A(n11954), .B(n11955), .Z(n11948) );
  ANDN U12925 ( .A(n11956), .B(n5051), .Z(n11955) );
  XOR U12926 ( .A(n11957), .B(n11958), .Z(n5051) );
  IV U12927 ( .A(n11954), .Z(n11957) );
  XNOR U12928 ( .A(n5052), .B(n11954), .Z(n11956) );
  NAND U12929 ( .A(n11959), .B(e_input[57]), .Z(n5052) );
  NAND U12930 ( .A(n6112), .B(e_input[57]), .Z(n11959) );
  XOR U12931 ( .A(n11960), .B(n11961), .Z(n11954) );
  ANDN U12932 ( .A(n11962), .B(n5073), .Z(n11961) );
  XOR U12933 ( .A(n11963), .B(n11964), .Z(n5073) );
  IV U12934 ( .A(n11960), .Z(n11963) );
  XNOR U12935 ( .A(n5074), .B(n11960), .Z(n11962) );
  NAND U12936 ( .A(n11965), .B(e_input[56]), .Z(n5074) );
  NAND U12937 ( .A(n6112), .B(e_input[56]), .Z(n11965) );
  XOR U12938 ( .A(n11966), .B(n11967), .Z(n11960) );
  ANDN U12939 ( .A(n11968), .B(n5095), .Z(n11967) );
  XOR U12940 ( .A(n11969), .B(n11970), .Z(n5095) );
  IV U12941 ( .A(n11966), .Z(n11969) );
  XNOR U12942 ( .A(n5096), .B(n11966), .Z(n11968) );
  NAND U12943 ( .A(n11971), .B(e_input[55]), .Z(n5096) );
  NAND U12944 ( .A(n6112), .B(e_input[55]), .Z(n11971) );
  XOR U12945 ( .A(n11972), .B(n11973), .Z(n11966) );
  ANDN U12946 ( .A(n11974), .B(n5117), .Z(n11973) );
  XOR U12947 ( .A(n11975), .B(n11976), .Z(n5117) );
  IV U12948 ( .A(n11972), .Z(n11975) );
  XNOR U12949 ( .A(n5118), .B(n11972), .Z(n11974) );
  NAND U12950 ( .A(n11977), .B(e_input[54]), .Z(n5118) );
  NAND U12951 ( .A(n6112), .B(e_input[54]), .Z(n11977) );
  XOR U12952 ( .A(n11978), .B(n11979), .Z(n11972) );
  ANDN U12953 ( .A(n11980), .B(n5139), .Z(n11979) );
  XOR U12954 ( .A(n11981), .B(n11982), .Z(n5139) );
  IV U12955 ( .A(n11978), .Z(n11981) );
  XNOR U12956 ( .A(n5140), .B(n11978), .Z(n11980) );
  NAND U12957 ( .A(n11983), .B(e_input[53]), .Z(n5140) );
  NAND U12958 ( .A(n6112), .B(e_input[53]), .Z(n11983) );
  XOR U12959 ( .A(n11984), .B(n11985), .Z(n11978) );
  ANDN U12960 ( .A(n11986), .B(n5161), .Z(n11985) );
  XOR U12961 ( .A(n11987), .B(n11988), .Z(n5161) );
  IV U12962 ( .A(n11984), .Z(n11987) );
  XNOR U12963 ( .A(n5162), .B(n11984), .Z(n11986) );
  NAND U12964 ( .A(n11989), .B(e_input[52]), .Z(n5162) );
  NAND U12965 ( .A(n6112), .B(e_input[52]), .Z(n11989) );
  XOR U12966 ( .A(n11990), .B(n11991), .Z(n11984) );
  ANDN U12967 ( .A(n11992), .B(n5183), .Z(n11991) );
  XOR U12968 ( .A(n11993), .B(n11994), .Z(n5183) );
  IV U12969 ( .A(n11990), .Z(n11993) );
  XNOR U12970 ( .A(n5184), .B(n11990), .Z(n11992) );
  NAND U12971 ( .A(n11995), .B(e_input[51]), .Z(n5184) );
  NAND U12972 ( .A(n6112), .B(e_input[51]), .Z(n11995) );
  XOR U12973 ( .A(n11996), .B(n11997), .Z(n11990) );
  ANDN U12974 ( .A(n11998), .B(n5205), .Z(n11997) );
  XOR U12975 ( .A(n11999), .B(n12000), .Z(n5205) );
  IV U12976 ( .A(n11996), .Z(n11999) );
  XNOR U12977 ( .A(n5206), .B(n11996), .Z(n11998) );
  NAND U12978 ( .A(n12001), .B(e_input[50]), .Z(n5206) );
  NAND U12979 ( .A(n6112), .B(e_input[50]), .Z(n12001) );
  XOR U12980 ( .A(n12002), .B(n12003), .Z(n11996) );
  ANDN U12981 ( .A(n12004), .B(n5229), .Z(n12003) );
  XOR U12982 ( .A(n12005), .B(n12006), .Z(n5229) );
  IV U12983 ( .A(n12002), .Z(n12005) );
  XNOR U12984 ( .A(n5230), .B(n12002), .Z(n12004) );
  NAND U12985 ( .A(n12007), .B(e_input[49]), .Z(n5230) );
  NAND U12986 ( .A(n6112), .B(e_input[49]), .Z(n12007) );
  XOR U12987 ( .A(n12008), .B(n12009), .Z(n12002) );
  ANDN U12988 ( .A(n12010), .B(n5251), .Z(n12009) );
  XOR U12989 ( .A(n12011), .B(n12012), .Z(n5251) );
  IV U12990 ( .A(n12008), .Z(n12011) );
  XNOR U12991 ( .A(n5252), .B(n12008), .Z(n12010) );
  NAND U12992 ( .A(n12013), .B(e_input[48]), .Z(n5252) );
  NAND U12993 ( .A(n6112), .B(e_input[48]), .Z(n12013) );
  XOR U12994 ( .A(n12014), .B(n12015), .Z(n12008) );
  ANDN U12995 ( .A(n12016), .B(n5273), .Z(n12015) );
  XOR U12996 ( .A(n12017), .B(n12018), .Z(n5273) );
  IV U12997 ( .A(n12014), .Z(n12017) );
  XNOR U12998 ( .A(n5274), .B(n12014), .Z(n12016) );
  NAND U12999 ( .A(n12019), .B(e_input[47]), .Z(n5274) );
  NAND U13000 ( .A(n6112), .B(e_input[47]), .Z(n12019) );
  XOR U13001 ( .A(n12020), .B(n12021), .Z(n12014) );
  ANDN U13002 ( .A(n12022), .B(n5295), .Z(n12021) );
  XOR U13003 ( .A(n12023), .B(n12024), .Z(n5295) );
  IV U13004 ( .A(n12020), .Z(n12023) );
  XNOR U13005 ( .A(n5296), .B(n12020), .Z(n12022) );
  NAND U13006 ( .A(n12025), .B(e_input[46]), .Z(n5296) );
  NAND U13007 ( .A(n6112), .B(e_input[46]), .Z(n12025) );
  XOR U13008 ( .A(n12026), .B(n12027), .Z(n12020) );
  ANDN U13009 ( .A(n12028), .B(n5317), .Z(n12027) );
  XOR U13010 ( .A(n12029), .B(n12030), .Z(n5317) );
  IV U13011 ( .A(n12026), .Z(n12029) );
  XNOR U13012 ( .A(n5318), .B(n12026), .Z(n12028) );
  NAND U13013 ( .A(n12031), .B(e_input[45]), .Z(n5318) );
  NAND U13014 ( .A(n6112), .B(e_input[45]), .Z(n12031) );
  XOR U13015 ( .A(n12032), .B(n12033), .Z(n12026) );
  ANDN U13016 ( .A(n12034), .B(n5339), .Z(n12033) );
  XOR U13017 ( .A(n12035), .B(n12036), .Z(n5339) );
  IV U13018 ( .A(n12032), .Z(n12035) );
  XNOR U13019 ( .A(n5340), .B(n12032), .Z(n12034) );
  NAND U13020 ( .A(n12037), .B(e_input[44]), .Z(n5340) );
  NAND U13021 ( .A(n6112), .B(e_input[44]), .Z(n12037) );
  XOR U13022 ( .A(n12038), .B(n12039), .Z(n12032) );
  ANDN U13023 ( .A(n12040), .B(n5361), .Z(n12039) );
  XOR U13024 ( .A(n12041), .B(n12042), .Z(n5361) );
  IV U13025 ( .A(n12038), .Z(n12041) );
  XNOR U13026 ( .A(n5362), .B(n12038), .Z(n12040) );
  NAND U13027 ( .A(n12043), .B(e_input[43]), .Z(n5362) );
  NAND U13028 ( .A(n6112), .B(e_input[43]), .Z(n12043) );
  XOR U13029 ( .A(n12044), .B(n12045), .Z(n12038) );
  ANDN U13030 ( .A(n12046), .B(n5383), .Z(n12045) );
  XOR U13031 ( .A(n12047), .B(n12048), .Z(n5383) );
  IV U13032 ( .A(n12044), .Z(n12047) );
  XNOR U13033 ( .A(n5384), .B(n12044), .Z(n12046) );
  NAND U13034 ( .A(n12049), .B(e_input[42]), .Z(n5384) );
  NAND U13035 ( .A(n6112), .B(e_input[42]), .Z(n12049) );
  XOR U13036 ( .A(n12050), .B(n12051), .Z(n12044) );
  ANDN U13037 ( .A(n12052), .B(n5405), .Z(n12051) );
  XOR U13038 ( .A(n12053), .B(n12054), .Z(n5405) );
  IV U13039 ( .A(n12050), .Z(n12053) );
  XNOR U13040 ( .A(n5406), .B(n12050), .Z(n12052) );
  NAND U13041 ( .A(n12055), .B(e_input[41]), .Z(n5406) );
  NAND U13042 ( .A(n6112), .B(e_input[41]), .Z(n12055) );
  XOR U13043 ( .A(n12056), .B(n12057), .Z(n12050) );
  ANDN U13044 ( .A(n12058), .B(n5427), .Z(n12057) );
  XOR U13045 ( .A(n12059), .B(n12060), .Z(n5427) );
  IV U13046 ( .A(n12056), .Z(n12059) );
  XNOR U13047 ( .A(n5428), .B(n12056), .Z(n12058) );
  NAND U13048 ( .A(n12061), .B(e_input[40]), .Z(n5428) );
  NAND U13049 ( .A(n6112), .B(e_input[40]), .Z(n12061) );
  XOR U13050 ( .A(n12062), .B(n12063), .Z(n12056) );
  ANDN U13051 ( .A(n12064), .B(n5451), .Z(n12063) );
  XOR U13052 ( .A(n12065), .B(n12066), .Z(n5451) );
  IV U13053 ( .A(n12062), .Z(n12065) );
  XNOR U13054 ( .A(n5452), .B(n12062), .Z(n12064) );
  NAND U13055 ( .A(n12067), .B(e_input[39]), .Z(n5452) );
  NAND U13056 ( .A(n6112), .B(e_input[39]), .Z(n12067) );
  XOR U13057 ( .A(n12068), .B(n12069), .Z(n12062) );
  ANDN U13058 ( .A(n12070), .B(n5473), .Z(n12069) );
  XOR U13059 ( .A(n12071), .B(n12072), .Z(n5473) );
  IV U13060 ( .A(n12068), .Z(n12071) );
  XNOR U13061 ( .A(n5474), .B(n12068), .Z(n12070) );
  NAND U13062 ( .A(n12073), .B(e_input[38]), .Z(n5474) );
  NAND U13063 ( .A(n6112), .B(e_input[38]), .Z(n12073) );
  XOR U13064 ( .A(n12074), .B(n12075), .Z(n12068) );
  ANDN U13065 ( .A(n12076), .B(n5495), .Z(n12075) );
  XOR U13066 ( .A(n12077), .B(n12078), .Z(n5495) );
  IV U13067 ( .A(n12074), .Z(n12077) );
  XNOR U13068 ( .A(n5496), .B(n12074), .Z(n12076) );
  NAND U13069 ( .A(n12079), .B(e_input[37]), .Z(n5496) );
  NAND U13070 ( .A(n6112), .B(e_input[37]), .Z(n12079) );
  XOR U13071 ( .A(n12080), .B(n12081), .Z(n12074) );
  ANDN U13072 ( .A(n12082), .B(n5517), .Z(n12081) );
  XOR U13073 ( .A(n12083), .B(n12084), .Z(n5517) );
  IV U13074 ( .A(n12080), .Z(n12083) );
  XNOR U13075 ( .A(n5518), .B(n12080), .Z(n12082) );
  NAND U13076 ( .A(n12085), .B(e_input[36]), .Z(n5518) );
  NAND U13077 ( .A(n6112), .B(e_input[36]), .Z(n12085) );
  XOR U13078 ( .A(n12086), .B(n12087), .Z(n12080) );
  ANDN U13079 ( .A(n12088), .B(n5539), .Z(n12087) );
  XOR U13080 ( .A(n12089), .B(n12090), .Z(n5539) );
  IV U13081 ( .A(n12086), .Z(n12089) );
  XNOR U13082 ( .A(n5540), .B(n12086), .Z(n12088) );
  NAND U13083 ( .A(n12091), .B(e_input[35]), .Z(n5540) );
  NAND U13084 ( .A(n6112), .B(e_input[35]), .Z(n12091) );
  XOR U13085 ( .A(n12092), .B(n12093), .Z(n12086) );
  ANDN U13086 ( .A(n12094), .B(n5561), .Z(n12093) );
  XOR U13087 ( .A(n12095), .B(n12096), .Z(n5561) );
  IV U13088 ( .A(n12092), .Z(n12095) );
  XNOR U13089 ( .A(n5562), .B(n12092), .Z(n12094) );
  NAND U13090 ( .A(n12097), .B(e_input[34]), .Z(n5562) );
  NAND U13091 ( .A(n6112), .B(e_input[34]), .Z(n12097) );
  XOR U13092 ( .A(n12098), .B(n12099), .Z(n12092) );
  ANDN U13093 ( .A(n12100), .B(n5583), .Z(n12099) );
  XOR U13094 ( .A(n12101), .B(n12102), .Z(n5583) );
  IV U13095 ( .A(n12098), .Z(n12101) );
  XNOR U13096 ( .A(n5584), .B(n12098), .Z(n12100) );
  NAND U13097 ( .A(n12103), .B(e_input[33]), .Z(n5584) );
  NAND U13098 ( .A(n6112), .B(e_input[33]), .Z(n12103) );
  XOR U13099 ( .A(n12104), .B(n12105), .Z(n12098) );
  ANDN U13100 ( .A(n12106), .B(n5605), .Z(n12105) );
  XOR U13101 ( .A(n12107), .B(n12108), .Z(n5605) );
  IV U13102 ( .A(n12104), .Z(n12107) );
  XNOR U13103 ( .A(n5606), .B(n12104), .Z(n12106) );
  NAND U13104 ( .A(n12109), .B(e_input[32]), .Z(n5606) );
  NAND U13105 ( .A(n6112), .B(e_input[32]), .Z(n12109) );
  XOR U13106 ( .A(n12110), .B(n12111), .Z(n12104) );
  ANDN U13107 ( .A(n12112), .B(n5627), .Z(n12111) );
  XOR U13108 ( .A(n12113), .B(n12114), .Z(n5627) );
  IV U13109 ( .A(n12110), .Z(n12113) );
  XNOR U13110 ( .A(n5628), .B(n12110), .Z(n12112) );
  NAND U13111 ( .A(n12115), .B(e_input[31]), .Z(n5628) );
  NAND U13112 ( .A(n6112), .B(e_input[31]), .Z(n12115) );
  XOR U13113 ( .A(n12116), .B(n12117), .Z(n12110) );
  ANDN U13114 ( .A(n12118), .B(n5649), .Z(n12117) );
  XOR U13115 ( .A(n12119), .B(n12120), .Z(n5649) );
  IV U13116 ( .A(n12116), .Z(n12119) );
  XNOR U13117 ( .A(n5650), .B(n12116), .Z(n12118) );
  NAND U13118 ( .A(n12121), .B(e_input[30]), .Z(n5650) );
  NAND U13119 ( .A(n6112), .B(e_input[30]), .Z(n12121) );
  XOR U13120 ( .A(n12122), .B(n12123), .Z(n12116) );
  ANDN U13121 ( .A(n12124), .B(n5673), .Z(n12123) );
  XOR U13122 ( .A(n12125), .B(n12126), .Z(n5673) );
  IV U13123 ( .A(n12122), .Z(n12125) );
  XNOR U13124 ( .A(n5674), .B(n12122), .Z(n12124) );
  NAND U13125 ( .A(n12127), .B(e_input[29]), .Z(n5674) );
  NAND U13126 ( .A(n6112), .B(e_input[29]), .Z(n12127) );
  XOR U13127 ( .A(n12128), .B(n12129), .Z(n12122) );
  ANDN U13128 ( .A(n12130), .B(n5695), .Z(n12129) );
  XOR U13129 ( .A(n12131), .B(n12132), .Z(n5695) );
  IV U13130 ( .A(n12128), .Z(n12131) );
  XNOR U13131 ( .A(n5696), .B(n12128), .Z(n12130) );
  NAND U13132 ( .A(n12133), .B(e_input[28]), .Z(n5696) );
  NAND U13133 ( .A(n6112), .B(e_input[28]), .Z(n12133) );
  XOR U13134 ( .A(n12134), .B(n12135), .Z(n12128) );
  ANDN U13135 ( .A(n12136), .B(n5717), .Z(n12135) );
  XOR U13136 ( .A(n12137), .B(n12138), .Z(n5717) );
  IV U13137 ( .A(n12134), .Z(n12137) );
  XNOR U13138 ( .A(n5718), .B(n12134), .Z(n12136) );
  NAND U13139 ( .A(n12139), .B(e_input[27]), .Z(n5718) );
  NAND U13140 ( .A(n6112), .B(e_input[27]), .Z(n12139) );
  XOR U13141 ( .A(n12140), .B(n12141), .Z(n12134) );
  ANDN U13142 ( .A(n12142), .B(n5739), .Z(n12141) );
  XOR U13143 ( .A(n12143), .B(n12144), .Z(n5739) );
  IV U13144 ( .A(n12140), .Z(n12143) );
  XNOR U13145 ( .A(n5740), .B(n12140), .Z(n12142) );
  NAND U13146 ( .A(n12145), .B(e_input[26]), .Z(n5740) );
  NAND U13147 ( .A(n6112), .B(e_input[26]), .Z(n12145) );
  XOR U13148 ( .A(n12146), .B(n12147), .Z(n12140) );
  ANDN U13149 ( .A(n12148), .B(n5761), .Z(n12147) );
  XOR U13150 ( .A(n12149), .B(n12150), .Z(n5761) );
  IV U13151 ( .A(n12146), .Z(n12149) );
  XNOR U13152 ( .A(n5762), .B(n12146), .Z(n12148) );
  NAND U13153 ( .A(n12151), .B(e_input[25]), .Z(n5762) );
  NAND U13154 ( .A(n6112), .B(e_input[25]), .Z(n12151) );
  XOR U13155 ( .A(n12152), .B(n12153), .Z(n12146) );
  ANDN U13156 ( .A(n12154), .B(n5783), .Z(n12153) );
  XOR U13157 ( .A(n12155), .B(n12156), .Z(n5783) );
  IV U13158 ( .A(n12152), .Z(n12155) );
  XNOR U13159 ( .A(n5784), .B(n12152), .Z(n12154) );
  NAND U13160 ( .A(n12157), .B(e_input[24]), .Z(n5784) );
  NAND U13161 ( .A(n6112), .B(e_input[24]), .Z(n12157) );
  XOR U13162 ( .A(n12158), .B(n12159), .Z(n12152) );
  ANDN U13163 ( .A(n12160), .B(n5805), .Z(n12159) );
  XOR U13164 ( .A(n12161), .B(n12162), .Z(n5805) );
  IV U13165 ( .A(n12158), .Z(n12161) );
  XNOR U13166 ( .A(n5806), .B(n12158), .Z(n12160) );
  NAND U13167 ( .A(n12163), .B(e_input[23]), .Z(n5806) );
  NAND U13168 ( .A(n6112), .B(e_input[23]), .Z(n12163) );
  XOR U13169 ( .A(n12164), .B(n12165), .Z(n12158) );
  ANDN U13170 ( .A(n12166), .B(n5827), .Z(n12165) );
  XOR U13171 ( .A(n12167), .B(n12168), .Z(n5827) );
  IV U13172 ( .A(n12164), .Z(n12167) );
  XNOR U13173 ( .A(n5828), .B(n12164), .Z(n12166) );
  NAND U13174 ( .A(n12169), .B(e_input[22]), .Z(n5828) );
  NAND U13175 ( .A(n6112), .B(e_input[22]), .Z(n12169) );
  XOR U13176 ( .A(n12170), .B(n12171), .Z(n12164) );
  ANDN U13177 ( .A(n12172), .B(n5849), .Z(n12171) );
  XOR U13178 ( .A(n12173), .B(n12174), .Z(n5849) );
  IV U13179 ( .A(n12170), .Z(n12173) );
  XNOR U13180 ( .A(n5850), .B(n12170), .Z(n12172) );
  NAND U13181 ( .A(n12175), .B(e_input[21]), .Z(n5850) );
  NAND U13182 ( .A(n6112), .B(e_input[21]), .Z(n12175) );
  XOR U13183 ( .A(n12176), .B(n12177), .Z(n12170) );
  ANDN U13184 ( .A(n12178), .B(n5871), .Z(n12177) );
  XOR U13185 ( .A(n12179), .B(n12180), .Z(n5871) );
  IV U13186 ( .A(n12176), .Z(n12179) );
  XNOR U13187 ( .A(n5872), .B(n12176), .Z(n12178) );
  NAND U13188 ( .A(n12181), .B(e_input[20]), .Z(n5872) );
  NAND U13189 ( .A(n6112), .B(e_input[20]), .Z(n12181) );
  XOR U13190 ( .A(n12182), .B(n12183), .Z(n12176) );
  ANDN U13191 ( .A(n12184), .B(n5895), .Z(n12183) );
  XOR U13192 ( .A(n12185), .B(n12186), .Z(n5895) );
  IV U13193 ( .A(n12182), .Z(n12185) );
  XNOR U13194 ( .A(n5896), .B(n12182), .Z(n12184) );
  NAND U13195 ( .A(n12187), .B(e_input[19]), .Z(n5896) );
  NAND U13196 ( .A(n6112), .B(e_input[19]), .Z(n12187) );
  XOR U13197 ( .A(n12188), .B(n12189), .Z(n12182) );
  ANDN U13198 ( .A(n12190), .B(n5917), .Z(n12189) );
  XOR U13199 ( .A(n12191), .B(n12192), .Z(n5917) );
  IV U13200 ( .A(n12188), .Z(n12191) );
  XNOR U13201 ( .A(n5918), .B(n12188), .Z(n12190) );
  NAND U13202 ( .A(n12193), .B(e_input[18]), .Z(n5918) );
  NAND U13203 ( .A(n6112), .B(e_input[18]), .Z(n12193) );
  XOR U13204 ( .A(n12194), .B(n12195), .Z(n12188) );
  ANDN U13205 ( .A(n12196), .B(n5939), .Z(n12195) );
  XOR U13206 ( .A(n12197), .B(n12198), .Z(n5939) );
  IV U13207 ( .A(n12194), .Z(n12197) );
  XNOR U13208 ( .A(n5940), .B(n12194), .Z(n12196) );
  NAND U13209 ( .A(n12199), .B(e_input[17]), .Z(n5940) );
  NAND U13210 ( .A(n6112), .B(e_input[17]), .Z(n12199) );
  XOR U13211 ( .A(n12200), .B(n12201), .Z(n12194) );
  ANDN U13212 ( .A(n12202), .B(n5961), .Z(n12201) );
  XOR U13213 ( .A(n12203), .B(n12204), .Z(n5961) );
  IV U13214 ( .A(n12200), .Z(n12203) );
  XNOR U13215 ( .A(n5962), .B(n12200), .Z(n12202) );
  NAND U13216 ( .A(n12205), .B(e_input[16]), .Z(n5962) );
  NAND U13217 ( .A(n6112), .B(e_input[16]), .Z(n12205) );
  XOR U13218 ( .A(n12206), .B(n12207), .Z(n12200) );
  ANDN U13219 ( .A(n12208), .B(n5983), .Z(n12207) );
  XOR U13220 ( .A(n12209), .B(n12210), .Z(n5983) );
  IV U13221 ( .A(n12206), .Z(n12209) );
  XNOR U13222 ( .A(n5984), .B(n12206), .Z(n12208) );
  NAND U13223 ( .A(n12211), .B(e_input[15]), .Z(n5984) );
  NAND U13224 ( .A(n6112), .B(e_input[15]), .Z(n12211) );
  XOR U13225 ( .A(n12212), .B(n12213), .Z(n12206) );
  ANDN U13226 ( .A(n12214), .B(n6005), .Z(n12213) );
  XOR U13227 ( .A(n12215), .B(n12216), .Z(n6005) );
  IV U13228 ( .A(n12212), .Z(n12215) );
  XNOR U13229 ( .A(n6006), .B(n12212), .Z(n12214) );
  NAND U13230 ( .A(n12217), .B(e_input[14]), .Z(n6006) );
  NAND U13231 ( .A(n6112), .B(e_input[14]), .Z(n12217) );
  XOR U13232 ( .A(n12218), .B(n12219), .Z(n12212) );
  ANDN U13233 ( .A(n12220), .B(n6027), .Z(n12219) );
  XOR U13234 ( .A(n12221), .B(n12222), .Z(n6027) );
  IV U13235 ( .A(n12218), .Z(n12221) );
  XNOR U13236 ( .A(n6028), .B(n12218), .Z(n12220) );
  NAND U13237 ( .A(n12223), .B(e_input[13]), .Z(n6028) );
  NAND U13238 ( .A(n6112), .B(e_input[13]), .Z(n12223) );
  XOR U13239 ( .A(n12224), .B(n12225), .Z(n12218) );
  ANDN U13240 ( .A(n12226), .B(n6049), .Z(n12225) );
  XOR U13241 ( .A(n12227), .B(n12228), .Z(n6049) );
  IV U13242 ( .A(n12224), .Z(n12227) );
  XNOR U13243 ( .A(n6050), .B(n12224), .Z(n12226) );
  NAND U13244 ( .A(n12229), .B(e_input[12]), .Z(n6050) );
  NAND U13245 ( .A(n6112), .B(e_input[12]), .Z(n12229) );
  XOR U13246 ( .A(n12230), .B(n12231), .Z(n12224) );
  ANDN U13247 ( .A(n12232), .B(n6071), .Z(n12231) );
  XOR U13248 ( .A(n12233), .B(n12234), .Z(n6071) );
  IV U13249 ( .A(n12230), .Z(n12233) );
  XNOR U13250 ( .A(n6072), .B(n12230), .Z(n12232) );
  NAND U13251 ( .A(n12235), .B(e_input[11]), .Z(n6072) );
  NAND U13252 ( .A(n6112), .B(e_input[11]), .Z(n12235) );
  XOR U13253 ( .A(n12236), .B(n12237), .Z(n12230) );
  ANDN U13254 ( .A(n12238), .B(n6093), .Z(n12237) );
  XOR U13255 ( .A(n12239), .B(n12240), .Z(n6093) );
  IV U13256 ( .A(n12236), .Z(n12239) );
  XNOR U13257 ( .A(n6094), .B(n12236), .Z(n12238) );
  NAND U13258 ( .A(n12241), .B(e_input[10]), .Z(n6094) );
  NAND U13259 ( .A(n6112), .B(e_input[10]), .Z(n12241) );
  XOR U13260 ( .A(n12242), .B(n12243), .Z(n12236) );
  ANDN U13261 ( .A(n12244), .B(n4117), .Z(n12243) );
  XOR U13262 ( .A(n12245), .B(n12246), .Z(n4117) );
  IV U13263 ( .A(n12242), .Z(n12245) );
  XNOR U13264 ( .A(n4118), .B(n12242), .Z(n12244) );
  NAND U13265 ( .A(n12247), .B(e_input[9]), .Z(n4118) );
  NAND U13266 ( .A(n6112), .B(e_input[9]), .Z(n12247) );
  XOR U13267 ( .A(n12248), .B(n12249), .Z(n12242) );
  ANDN U13268 ( .A(n12250), .B(n4339), .Z(n12249) );
  XOR U13269 ( .A(n12251), .B(n12252), .Z(n4339) );
  IV U13270 ( .A(n12248), .Z(n12251) );
  XNOR U13271 ( .A(n4340), .B(n12248), .Z(n12250) );
  NAND U13272 ( .A(n12253), .B(e_input[8]), .Z(n4340) );
  NAND U13273 ( .A(n6112), .B(e_input[8]), .Z(n12253) );
  XOR U13274 ( .A(n12254), .B(n12255), .Z(n12248) );
  ANDN U13275 ( .A(n12256), .B(n4561), .Z(n12255) );
  XOR U13276 ( .A(n12257), .B(n12258), .Z(n4561) );
  IV U13277 ( .A(n12254), .Z(n12257) );
  XNOR U13278 ( .A(n4562), .B(n12254), .Z(n12256) );
  NAND U13279 ( .A(n12259), .B(e_input[7]), .Z(n4562) );
  NAND U13280 ( .A(n6112), .B(e_input[7]), .Z(n12259) );
  XOR U13281 ( .A(n12260), .B(n12261), .Z(n12254) );
  ANDN U13282 ( .A(n12262), .B(n4783), .Z(n12261) );
  XOR U13283 ( .A(n12263), .B(n12264), .Z(n4783) );
  IV U13284 ( .A(n12260), .Z(n12263) );
  XNOR U13285 ( .A(n4784), .B(n12260), .Z(n12262) );
  NAND U13286 ( .A(n12265), .B(e_input[6]), .Z(n4784) );
  NAND U13287 ( .A(n6112), .B(e_input[6]), .Z(n12265) );
  XOR U13288 ( .A(n12266), .B(n12267), .Z(n12260) );
  ANDN U13289 ( .A(n12268), .B(n5005), .Z(n12267) );
  XOR U13290 ( .A(n12269), .B(n12270), .Z(n5005) );
  IV U13291 ( .A(n12266), .Z(n12269) );
  XNOR U13292 ( .A(n5006), .B(n12266), .Z(n12268) );
  NAND U13293 ( .A(n12271), .B(e_input[5]), .Z(n5006) );
  NAND U13294 ( .A(n6112), .B(e_input[5]), .Z(n12271) );
  XOR U13295 ( .A(n12272), .B(n12273), .Z(n12266) );
  ANDN U13296 ( .A(n12274), .B(n5227), .Z(n12273) );
  XOR U13297 ( .A(n12275), .B(n12276), .Z(n5227) );
  IV U13298 ( .A(n12272), .Z(n12275) );
  XNOR U13299 ( .A(n5228), .B(n12272), .Z(n12274) );
  NAND U13300 ( .A(n12277), .B(e_input[4]), .Z(n5228) );
  NAND U13301 ( .A(n6112), .B(e_input[4]), .Z(n12277) );
  XOR U13302 ( .A(n12278), .B(n12279), .Z(n12272) );
  ANDN U13303 ( .A(n12280), .B(n5449), .Z(n12279) );
  XOR U13304 ( .A(n12281), .B(n12282), .Z(n5449) );
  IV U13305 ( .A(n12278), .Z(n12281) );
  XNOR U13306 ( .A(n5450), .B(n12278), .Z(n12280) );
  NAND U13307 ( .A(n12283), .B(e_input[3]), .Z(n5450) );
  NAND U13308 ( .A(n6112), .B(e_input[3]), .Z(n12283) );
  XNOR U13309 ( .A(n12284), .B(n12285), .Z(n12278) );
  ANDN U13310 ( .A(n12286), .B(n5671), .Z(n12285) );
  XOR U13311 ( .A(n12284), .B(n12287), .Z(n5671) );
  XOR U13312 ( .A(n5672), .B(n12284), .Z(n12286) );
  NAND U13313 ( .A(n12288), .B(e_input[2]), .Z(n5672) );
  NAND U13314 ( .A(n6112), .B(e_input[2]), .Z(n12288) );
  XOR U13315 ( .A(n12289), .B(n12290), .Z(n12284) );
  NANDN U13316 ( .B(n5893), .A(n12291), .Z(n12289) );
  XOR U13317 ( .A(n12292), .B(n5894), .Z(n12291) );
  NAND U13318 ( .A(n12293), .B(e_input[1]), .Z(n5894) );
  NAND U13319 ( .A(n6112), .B(e_input[1]), .Z(n12293) );
  XNOR U13320 ( .A(n12294), .B(n12292), .Z(n5893) );
  IV U13321 ( .A(n12290), .Z(n12292) );
  ANDN U13322 ( .A(n12295), .B(n12296), .Z(n12290) );
  XOR U13323 ( .A(n12295), .B(n12296), .Z(mod_mult_o[0]) );
  NAND U13324 ( .A(n12297), .B(e_input[0]), .Z(n12296) );
  NAND U13325 ( .A(n6112), .B(e_input[0]), .Z(n12297) );
  XOR U13326 ( .A(n12298), .B(n12299), .Z(n6112) );
  AND U13327 ( .A(n12300), .B(n12301), .Z(n12299) );
  IV U13328 ( .A(n12298), .Z(n12301) );
  XOR U13329 ( .A(n12302), .B(n12303), .Z(n12300) );
  XOR U13330 ( .A(n12304), .B(n12298), .Z(n12303) );
  XNOR U13331 ( .A(n12305), .B(n12306), .Z(n12302) );
  NOR U13332 ( .A(n12307), .B(n4112), .Z(n12305) );
  XOR U13333 ( .A(n12308), .B(n12309), .Z(n12298) );
  AND U13334 ( .A(n12310), .B(n12311), .Z(n12309) );
  IV U13335 ( .A(n12308), .Z(n12311) );
  XOR U13336 ( .A(n12308), .B(n4112), .Z(n12310) );
  XNOR U13337 ( .A(n12307), .B(n12312), .Z(n4112) );
  IV U13338 ( .A(n12304), .Z(n12307) );
  XOR U13339 ( .A(n12313), .B(n12314), .Z(n12304) );
  AND U13340 ( .A(n12315), .B(n12316), .Z(n12314) );
  XNOR U13341 ( .A(n12317), .B(n12313), .Z(n12316) );
  XOR U13342 ( .A(n12318), .B(n12319), .Z(n12308) );
  AND U13343 ( .A(n12320), .B(n12321), .Z(n12319) );
  XNOR U13344 ( .A(n12318), .B(n6113), .Z(n12321) );
  XNOR U13345 ( .A(n12315), .B(n12317), .Z(n6113) );
  NAND U13346 ( .A(n12322), .B(e_input[1023]), .Z(n12317) );
  NAND U13347 ( .A(n12323), .B(e_input[1023]), .Z(n12322) );
  XNOR U13348 ( .A(n12313), .B(n12324), .Z(n12315) );
  XOR U13349 ( .A(n12325), .B(n12326), .Z(n12313) );
  AND U13350 ( .A(n12327), .B(n12328), .Z(n12326) );
  XNOR U13351 ( .A(n12329), .B(n12325), .Z(n12328) );
  XOR U13352 ( .A(n12330), .B(e_input[1023]), .Z(n12320) );
  IV U13353 ( .A(n12318), .Z(n12330) );
  XOR U13354 ( .A(n12331), .B(n12332), .Z(n12318) );
  AND U13355 ( .A(n12333), .B(n12334), .Z(n12332) );
  XNOR U13356 ( .A(n12331), .B(n6121), .Z(n12334) );
  XNOR U13357 ( .A(n12327), .B(n12329), .Z(n6121) );
  NAND U13358 ( .A(n12335), .B(e_input[1022]), .Z(n12329) );
  NAND U13359 ( .A(n12323), .B(e_input[1022]), .Z(n12335) );
  XNOR U13360 ( .A(n12325), .B(n12336), .Z(n12327) );
  XOR U13361 ( .A(n12337), .B(n12338), .Z(n12325) );
  AND U13362 ( .A(n12339), .B(n12340), .Z(n12338) );
  XNOR U13363 ( .A(n12341), .B(n12337), .Z(n12340) );
  XOR U13364 ( .A(n12342), .B(e_input[1022]), .Z(n12333) );
  IV U13365 ( .A(n12331), .Z(n12342) );
  XOR U13366 ( .A(n12343), .B(n12344), .Z(n12331) );
  AND U13367 ( .A(n12345), .B(n12346), .Z(n12344) );
  XNOR U13368 ( .A(n12343), .B(n6129), .Z(n12346) );
  XNOR U13369 ( .A(n12339), .B(n12341), .Z(n6129) );
  NAND U13370 ( .A(n12347), .B(e_input[1021]), .Z(n12341) );
  NAND U13371 ( .A(n12323), .B(e_input[1021]), .Z(n12347) );
  XNOR U13372 ( .A(n12337), .B(n12348), .Z(n12339) );
  XOR U13373 ( .A(n12349), .B(n12350), .Z(n12337) );
  AND U13374 ( .A(n12351), .B(n12352), .Z(n12350) );
  XNOR U13375 ( .A(n12353), .B(n12349), .Z(n12352) );
  XOR U13376 ( .A(n12354), .B(e_input[1021]), .Z(n12345) );
  IV U13377 ( .A(n12343), .Z(n12354) );
  XOR U13378 ( .A(n12355), .B(n12356), .Z(n12343) );
  AND U13379 ( .A(n12357), .B(n12358), .Z(n12356) );
  XNOR U13380 ( .A(n12355), .B(n6137), .Z(n12358) );
  XNOR U13381 ( .A(n12351), .B(n12353), .Z(n6137) );
  NAND U13382 ( .A(n12359), .B(e_input[1020]), .Z(n12353) );
  NAND U13383 ( .A(n12323), .B(e_input[1020]), .Z(n12359) );
  XNOR U13384 ( .A(n12349), .B(n12360), .Z(n12351) );
  XOR U13385 ( .A(n12361), .B(n12362), .Z(n12349) );
  AND U13386 ( .A(n12363), .B(n12364), .Z(n12362) );
  XNOR U13387 ( .A(n12365), .B(n12361), .Z(n12364) );
  XOR U13388 ( .A(n12366), .B(e_input[1020]), .Z(n12357) );
  IV U13389 ( .A(n12355), .Z(n12366) );
  XOR U13390 ( .A(n12367), .B(n12368), .Z(n12355) );
  AND U13391 ( .A(n12369), .B(n12370), .Z(n12368) );
  XNOR U13392 ( .A(n12367), .B(n6147), .Z(n12370) );
  XNOR U13393 ( .A(n12363), .B(n12365), .Z(n6147) );
  NAND U13394 ( .A(n12371), .B(e_input[1019]), .Z(n12365) );
  NAND U13395 ( .A(n12323), .B(e_input[1019]), .Z(n12371) );
  XNOR U13396 ( .A(n12361), .B(n12372), .Z(n12363) );
  XOR U13397 ( .A(n12373), .B(n12374), .Z(n12361) );
  AND U13398 ( .A(n12375), .B(n12376), .Z(n12374) );
  XNOR U13399 ( .A(n12377), .B(n12373), .Z(n12376) );
  XOR U13400 ( .A(n12378), .B(e_input[1019]), .Z(n12369) );
  IV U13401 ( .A(n12367), .Z(n12378) );
  XOR U13402 ( .A(n12379), .B(n12380), .Z(n12367) );
  AND U13403 ( .A(n12381), .B(n12382), .Z(n12380) );
  XNOR U13404 ( .A(n12379), .B(n6155), .Z(n12382) );
  XNOR U13405 ( .A(n12375), .B(n12377), .Z(n6155) );
  NAND U13406 ( .A(n12383), .B(e_input[1018]), .Z(n12377) );
  NAND U13407 ( .A(n12323), .B(e_input[1018]), .Z(n12383) );
  XNOR U13408 ( .A(n12373), .B(n12384), .Z(n12375) );
  XOR U13409 ( .A(n12385), .B(n12386), .Z(n12373) );
  AND U13410 ( .A(n12387), .B(n12388), .Z(n12386) );
  XNOR U13411 ( .A(n12389), .B(n12385), .Z(n12388) );
  XOR U13412 ( .A(n12390), .B(e_input[1018]), .Z(n12381) );
  IV U13413 ( .A(n12379), .Z(n12390) );
  XOR U13414 ( .A(n12391), .B(n12392), .Z(n12379) );
  AND U13415 ( .A(n12393), .B(n12394), .Z(n12392) );
  XNOR U13416 ( .A(n12391), .B(n6163), .Z(n12394) );
  XNOR U13417 ( .A(n12387), .B(n12389), .Z(n6163) );
  NAND U13418 ( .A(n12395), .B(e_input[1017]), .Z(n12389) );
  NAND U13419 ( .A(n12323), .B(e_input[1017]), .Z(n12395) );
  XNOR U13420 ( .A(n12385), .B(n12396), .Z(n12387) );
  XOR U13421 ( .A(n12397), .B(n12398), .Z(n12385) );
  AND U13422 ( .A(n12399), .B(n12400), .Z(n12398) );
  XNOR U13423 ( .A(n12401), .B(n12397), .Z(n12400) );
  XOR U13424 ( .A(n12402), .B(e_input[1017]), .Z(n12393) );
  IV U13425 ( .A(n12391), .Z(n12402) );
  XOR U13426 ( .A(n12403), .B(n12404), .Z(n12391) );
  AND U13427 ( .A(n12405), .B(n12406), .Z(n12404) );
  XNOR U13428 ( .A(n12403), .B(n6171), .Z(n12406) );
  XNOR U13429 ( .A(n12399), .B(n12401), .Z(n6171) );
  NAND U13430 ( .A(n12407), .B(e_input[1016]), .Z(n12401) );
  NAND U13431 ( .A(n12323), .B(e_input[1016]), .Z(n12407) );
  XNOR U13432 ( .A(n12397), .B(n12408), .Z(n12399) );
  XOR U13433 ( .A(n12409), .B(n12410), .Z(n12397) );
  AND U13434 ( .A(n12411), .B(n12412), .Z(n12410) );
  XNOR U13435 ( .A(n12413), .B(n12409), .Z(n12412) );
  XOR U13436 ( .A(n12414), .B(e_input[1016]), .Z(n12405) );
  IV U13437 ( .A(n12403), .Z(n12414) );
  XOR U13438 ( .A(n12415), .B(n12416), .Z(n12403) );
  AND U13439 ( .A(n12417), .B(n12418), .Z(n12416) );
  XNOR U13440 ( .A(n12415), .B(n6179), .Z(n12418) );
  XNOR U13441 ( .A(n12411), .B(n12413), .Z(n6179) );
  NAND U13442 ( .A(n12419), .B(e_input[1015]), .Z(n12413) );
  NAND U13443 ( .A(n12323), .B(e_input[1015]), .Z(n12419) );
  XNOR U13444 ( .A(n12409), .B(n12420), .Z(n12411) );
  XOR U13445 ( .A(n12421), .B(n12422), .Z(n12409) );
  AND U13446 ( .A(n12423), .B(n12424), .Z(n12422) );
  XNOR U13447 ( .A(n12425), .B(n12421), .Z(n12424) );
  XOR U13448 ( .A(n12426), .B(e_input[1015]), .Z(n12417) );
  IV U13449 ( .A(n12415), .Z(n12426) );
  XOR U13450 ( .A(n12427), .B(n12428), .Z(n12415) );
  AND U13451 ( .A(n12429), .B(n12430), .Z(n12428) );
  XNOR U13452 ( .A(n12427), .B(n6187), .Z(n12430) );
  XNOR U13453 ( .A(n12423), .B(n12425), .Z(n6187) );
  NAND U13454 ( .A(n12431), .B(e_input[1014]), .Z(n12425) );
  NAND U13455 ( .A(n12323), .B(e_input[1014]), .Z(n12431) );
  XNOR U13456 ( .A(n12421), .B(n12432), .Z(n12423) );
  XOR U13457 ( .A(n12433), .B(n12434), .Z(n12421) );
  AND U13458 ( .A(n12435), .B(n12436), .Z(n12434) );
  XNOR U13459 ( .A(n12437), .B(n12433), .Z(n12436) );
  XOR U13460 ( .A(n12438), .B(e_input[1014]), .Z(n12429) );
  IV U13461 ( .A(n12427), .Z(n12438) );
  XOR U13462 ( .A(n12439), .B(n12440), .Z(n12427) );
  AND U13463 ( .A(n12441), .B(n12442), .Z(n12440) );
  XNOR U13464 ( .A(n12439), .B(n6195), .Z(n12442) );
  XNOR U13465 ( .A(n12435), .B(n12437), .Z(n6195) );
  NAND U13466 ( .A(n12443), .B(e_input[1013]), .Z(n12437) );
  NAND U13467 ( .A(n12323), .B(e_input[1013]), .Z(n12443) );
  XNOR U13468 ( .A(n12433), .B(n12444), .Z(n12435) );
  XOR U13469 ( .A(n12445), .B(n12446), .Z(n12433) );
  AND U13470 ( .A(n12447), .B(n12448), .Z(n12446) );
  XNOR U13471 ( .A(n12449), .B(n12445), .Z(n12448) );
  XOR U13472 ( .A(n12450), .B(e_input[1013]), .Z(n12441) );
  IV U13473 ( .A(n12439), .Z(n12450) );
  XOR U13474 ( .A(n12451), .B(n12452), .Z(n12439) );
  AND U13475 ( .A(n12453), .B(n12454), .Z(n12452) );
  XNOR U13476 ( .A(n12451), .B(n6203), .Z(n12454) );
  XNOR U13477 ( .A(n12447), .B(n12449), .Z(n6203) );
  NAND U13478 ( .A(n12455), .B(e_input[1012]), .Z(n12449) );
  NAND U13479 ( .A(n12323), .B(e_input[1012]), .Z(n12455) );
  XNOR U13480 ( .A(n12445), .B(n12456), .Z(n12447) );
  XOR U13481 ( .A(n12457), .B(n12458), .Z(n12445) );
  AND U13482 ( .A(n12459), .B(n12460), .Z(n12458) );
  XNOR U13483 ( .A(n12461), .B(n12457), .Z(n12460) );
  XOR U13484 ( .A(n12462), .B(e_input[1012]), .Z(n12453) );
  IV U13485 ( .A(n12451), .Z(n12462) );
  XOR U13486 ( .A(n12463), .B(n12464), .Z(n12451) );
  AND U13487 ( .A(n12465), .B(n12466), .Z(n12464) );
  XNOR U13488 ( .A(n12463), .B(n6211), .Z(n12466) );
  XNOR U13489 ( .A(n12459), .B(n12461), .Z(n6211) );
  NAND U13490 ( .A(n12467), .B(e_input[1011]), .Z(n12461) );
  NAND U13491 ( .A(n12323), .B(e_input[1011]), .Z(n12467) );
  XNOR U13492 ( .A(n12457), .B(n12468), .Z(n12459) );
  XOR U13493 ( .A(n12469), .B(n12470), .Z(n12457) );
  AND U13494 ( .A(n12471), .B(n12472), .Z(n12470) );
  XNOR U13495 ( .A(n12473), .B(n12469), .Z(n12472) );
  XOR U13496 ( .A(n12474), .B(e_input[1011]), .Z(n12465) );
  IV U13497 ( .A(n12463), .Z(n12474) );
  XOR U13498 ( .A(n12475), .B(n12476), .Z(n12463) );
  AND U13499 ( .A(n12477), .B(n12478), .Z(n12476) );
  XNOR U13500 ( .A(n12475), .B(n6219), .Z(n12478) );
  XNOR U13501 ( .A(n12471), .B(n12473), .Z(n6219) );
  NAND U13502 ( .A(n12479), .B(e_input[1010]), .Z(n12473) );
  NAND U13503 ( .A(n12323), .B(e_input[1010]), .Z(n12479) );
  XNOR U13504 ( .A(n12469), .B(n12480), .Z(n12471) );
  XOR U13505 ( .A(n12481), .B(n12482), .Z(n12469) );
  AND U13506 ( .A(n12483), .B(n12484), .Z(n12482) );
  XNOR U13507 ( .A(n12485), .B(n12481), .Z(n12484) );
  XOR U13508 ( .A(n12486), .B(e_input[1010]), .Z(n12477) );
  IV U13509 ( .A(n12475), .Z(n12486) );
  XOR U13510 ( .A(n12487), .B(n12488), .Z(n12475) );
  AND U13511 ( .A(n12489), .B(n12490), .Z(n12488) );
  XNOR U13512 ( .A(n12487), .B(n6229), .Z(n12490) );
  XNOR U13513 ( .A(n12483), .B(n12485), .Z(n6229) );
  NAND U13514 ( .A(n12491), .B(e_input[1009]), .Z(n12485) );
  NAND U13515 ( .A(n12323), .B(e_input[1009]), .Z(n12491) );
  XNOR U13516 ( .A(n12481), .B(n12492), .Z(n12483) );
  XOR U13517 ( .A(n12493), .B(n12494), .Z(n12481) );
  AND U13518 ( .A(n12495), .B(n12496), .Z(n12494) );
  XNOR U13519 ( .A(n12497), .B(n12493), .Z(n12496) );
  XOR U13520 ( .A(n12498), .B(e_input[1009]), .Z(n12489) );
  IV U13521 ( .A(n12487), .Z(n12498) );
  XOR U13522 ( .A(n12499), .B(n12500), .Z(n12487) );
  AND U13523 ( .A(n12501), .B(n12502), .Z(n12500) );
  XNOR U13524 ( .A(n12499), .B(n6237), .Z(n12502) );
  XNOR U13525 ( .A(n12495), .B(n12497), .Z(n6237) );
  NAND U13526 ( .A(n12503), .B(e_input[1008]), .Z(n12497) );
  NAND U13527 ( .A(n12323), .B(e_input[1008]), .Z(n12503) );
  XNOR U13528 ( .A(n12493), .B(n12504), .Z(n12495) );
  XOR U13529 ( .A(n12505), .B(n12506), .Z(n12493) );
  AND U13530 ( .A(n12507), .B(n12508), .Z(n12506) );
  XNOR U13531 ( .A(n12509), .B(n12505), .Z(n12508) );
  XOR U13532 ( .A(n12510), .B(e_input[1008]), .Z(n12501) );
  IV U13533 ( .A(n12499), .Z(n12510) );
  XOR U13534 ( .A(n12511), .B(n12512), .Z(n12499) );
  AND U13535 ( .A(n12513), .B(n12514), .Z(n12512) );
  XNOR U13536 ( .A(n12511), .B(n6245), .Z(n12514) );
  XNOR U13537 ( .A(n12507), .B(n12509), .Z(n6245) );
  NAND U13538 ( .A(n12515), .B(e_input[1007]), .Z(n12509) );
  NAND U13539 ( .A(n12323), .B(e_input[1007]), .Z(n12515) );
  XNOR U13540 ( .A(n12505), .B(n12516), .Z(n12507) );
  XOR U13541 ( .A(n12517), .B(n12518), .Z(n12505) );
  AND U13542 ( .A(n12519), .B(n12520), .Z(n12518) );
  XNOR U13543 ( .A(n12521), .B(n12517), .Z(n12520) );
  XOR U13544 ( .A(n12522), .B(e_input[1007]), .Z(n12513) );
  IV U13545 ( .A(n12511), .Z(n12522) );
  XOR U13546 ( .A(n12523), .B(n12524), .Z(n12511) );
  AND U13547 ( .A(n12525), .B(n12526), .Z(n12524) );
  XNOR U13548 ( .A(n12523), .B(n6253), .Z(n12526) );
  XNOR U13549 ( .A(n12519), .B(n12521), .Z(n6253) );
  NAND U13550 ( .A(n12527), .B(e_input[1006]), .Z(n12521) );
  NAND U13551 ( .A(n12323), .B(e_input[1006]), .Z(n12527) );
  XNOR U13552 ( .A(n12517), .B(n12528), .Z(n12519) );
  XOR U13553 ( .A(n12529), .B(n12530), .Z(n12517) );
  AND U13554 ( .A(n12531), .B(n12532), .Z(n12530) );
  XNOR U13555 ( .A(n12533), .B(n12529), .Z(n12532) );
  XOR U13556 ( .A(n12534), .B(e_input[1006]), .Z(n12525) );
  IV U13557 ( .A(n12523), .Z(n12534) );
  XOR U13558 ( .A(n12535), .B(n12536), .Z(n12523) );
  AND U13559 ( .A(n12537), .B(n12538), .Z(n12536) );
  XNOR U13560 ( .A(n12535), .B(n6261), .Z(n12538) );
  XNOR U13561 ( .A(n12531), .B(n12533), .Z(n6261) );
  NAND U13562 ( .A(n12539), .B(e_input[1005]), .Z(n12533) );
  NAND U13563 ( .A(n12323), .B(e_input[1005]), .Z(n12539) );
  XNOR U13564 ( .A(n12529), .B(n12540), .Z(n12531) );
  XOR U13565 ( .A(n12541), .B(n12542), .Z(n12529) );
  AND U13566 ( .A(n12543), .B(n12544), .Z(n12542) );
  XNOR U13567 ( .A(n12545), .B(n12541), .Z(n12544) );
  XOR U13568 ( .A(n12546), .B(e_input[1005]), .Z(n12537) );
  IV U13569 ( .A(n12535), .Z(n12546) );
  XOR U13570 ( .A(n12547), .B(n12548), .Z(n12535) );
  AND U13571 ( .A(n12549), .B(n12550), .Z(n12548) );
  XNOR U13572 ( .A(n12547), .B(n6269), .Z(n12550) );
  XNOR U13573 ( .A(n12543), .B(n12545), .Z(n6269) );
  NAND U13574 ( .A(n12551), .B(e_input[1004]), .Z(n12545) );
  NAND U13575 ( .A(n12323), .B(e_input[1004]), .Z(n12551) );
  XNOR U13576 ( .A(n12541), .B(n12552), .Z(n12543) );
  XOR U13577 ( .A(n12553), .B(n12554), .Z(n12541) );
  AND U13578 ( .A(n12555), .B(n12556), .Z(n12554) );
  XNOR U13579 ( .A(n12557), .B(n12553), .Z(n12556) );
  XOR U13580 ( .A(n12558), .B(e_input[1004]), .Z(n12549) );
  IV U13581 ( .A(n12547), .Z(n12558) );
  XOR U13582 ( .A(n12559), .B(n12560), .Z(n12547) );
  AND U13583 ( .A(n12561), .B(n12562), .Z(n12560) );
  XNOR U13584 ( .A(n12559), .B(n6277), .Z(n12562) );
  XNOR U13585 ( .A(n12555), .B(n12557), .Z(n6277) );
  NAND U13586 ( .A(n12563), .B(e_input[1003]), .Z(n12557) );
  NAND U13587 ( .A(n12323), .B(e_input[1003]), .Z(n12563) );
  XNOR U13588 ( .A(n12553), .B(n12564), .Z(n12555) );
  XOR U13589 ( .A(n12565), .B(n12566), .Z(n12553) );
  AND U13590 ( .A(n12567), .B(n12568), .Z(n12566) );
  XNOR U13591 ( .A(n12569), .B(n12565), .Z(n12568) );
  XOR U13592 ( .A(n12570), .B(e_input[1003]), .Z(n12561) );
  IV U13593 ( .A(n12559), .Z(n12570) );
  XOR U13594 ( .A(n12571), .B(n12572), .Z(n12559) );
  AND U13595 ( .A(n12573), .B(n12574), .Z(n12572) );
  XNOR U13596 ( .A(n12571), .B(n6285), .Z(n12574) );
  XNOR U13597 ( .A(n12567), .B(n12569), .Z(n6285) );
  NAND U13598 ( .A(n12575), .B(e_input[1002]), .Z(n12569) );
  NAND U13599 ( .A(n12323), .B(e_input[1002]), .Z(n12575) );
  XNOR U13600 ( .A(n12565), .B(n12576), .Z(n12567) );
  XOR U13601 ( .A(n12577), .B(n12578), .Z(n12565) );
  AND U13602 ( .A(n12579), .B(n12580), .Z(n12578) );
  XNOR U13603 ( .A(n12581), .B(n12577), .Z(n12580) );
  XOR U13604 ( .A(n12582), .B(e_input[1002]), .Z(n12573) );
  IV U13605 ( .A(n12571), .Z(n12582) );
  XOR U13606 ( .A(n12583), .B(n12584), .Z(n12571) );
  AND U13607 ( .A(n12585), .B(n12586), .Z(n12584) );
  XNOR U13608 ( .A(n12583), .B(n6293), .Z(n12586) );
  XNOR U13609 ( .A(n12579), .B(n12581), .Z(n6293) );
  NAND U13610 ( .A(n12587), .B(e_input[1001]), .Z(n12581) );
  NAND U13611 ( .A(n12323), .B(e_input[1001]), .Z(n12587) );
  XNOR U13612 ( .A(n12577), .B(n12588), .Z(n12579) );
  XOR U13613 ( .A(n12589), .B(n12590), .Z(n12577) );
  AND U13614 ( .A(n12591), .B(n12592), .Z(n12590) );
  XNOR U13615 ( .A(n12593), .B(n12589), .Z(n12592) );
  XOR U13616 ( .A(n12594), .B(e_input[1001]), .Z(n12585) );
  IV U13617 ( .A(n12583), .Z(n12594) );
  XOR U13618 ( .A(n12595), .B(n12596), .Z(n12583) );
  AND U13619 ( .A(n12597), .B(n12598), .Z(n12596) );
  XNOR U13620 ( .A(n12595), .B(n6301), .Z(n12598) );
  XNOR U13621 ( .A(n12591), .B(n12593), .Z(n6301) );
  NAND U13622 ( .A(n12599), .B(e_input[1000]), .Z(n12593) );
  NAND U13623 ( .A(n12323), .B(e_input[1000]), .Z(n12599) );
  XNOR U13624 ( .A(n12589), .B(n12600), .Z(n12591) );
  XOR U13625 ( .A(n12601), .B(n12602), .Z(n12589) );
  AND U13626 ( .A(n12603), .B(n12604), .Z(n12602) );
  XNOR U13627 ( .A(n12605), .B(n12601), .Z(n12604) );
  XOR U13628 ( .A(n12606), .B(e_input[1000]), .Z(n12597) );
  IV U13629 ( .A(n12595), .Z(n12606) );
  XOR U13630 ( .A(n12607), .B(n12608), .Z(n12595) );
  AND U13631 ( .A(n12609), .B(n12610), .Z(n12608) );
  XNOR U13632 ( .A(n12607), .B(n6306), .Z(n12610) );
  XNOR U13633 ( .A(n12603), .B(n12605), .Z(n6306) );
  NAND U13634 ( .A(n12611), .B(e_input[999]), .Z(n12605) );
  NAND U13635 ( .A(n12323), .B(e_input[999]), .Z(n12611) );
  XNOR U13636 ( .A(n12601), .B(n12612), .Z(n12603) );
  XOR U13637 ( .A(n12613), .B(n12614), .Z(n12601) );
  AND U13638 ( .A(n12615), .B(n12616), .Z(n12614) );
  XNOR U13639 ( .A(n12617), .B(n12613), .Z(n12616) );
  XOR U13640 ( .A(n12618), .B(e_input[999]), .Z(n12609) );
  IV U13641 ( .A(n12607), .Z(n12618) );
  XOR U13642 ( .A(n12619), .B(n12620), .Z(n12607) );
  AND U13643 ( .A(n12621), .B(n12622), .Z(n12620) );
  XNOR U13644 ( .A(n12619), .B(n6312), .Z(n12622) );
  XNOR U13645 ( .A(n12615), .B(n12617), .Z(n6312) );
  NAND U13646 ( .A(n12623), .B(e_input[998]), .Z(n12617) );
  NAND U13647 ( .A(n12323), .B(e_input[998]), .Z(n12623) );
  XNOR U13648 ( .A(n12613), .B(n12624), .Z(n12615) );
  XOR U13649 ( .A(n12625), .B(n12626), .Z(n12613) );
  AND U13650 ( .A(n12627), .B(n12628), .Z(n12626) );
  XNOR U13651 ( .A(n12629), .B(n12625), .Z(n12628) );
  XOR U13652 ( .A(n12630), .B(e_input[998]), .Z(n12621) );
  IV U13653 ( .A(n12619), .Z(n12630) );
  XOR U13654 ( .A(n12631), .B(n12632), .Z(n12619) );
  AND U13655 ( .A(n12633), .B(n12634), .Z(n12632) );
  XNOR U13656 ( .A(n12631), .B(n6318), .Z(n12634) );
  XNOR U13657 ( .A(n12627), .B(n12629), .Z(n6318) );
  NAND U13658 ( .A(n12635), .B(e_input[997]), .Z(n12629) );
  NAND U13659 ( .A(n12323), .B(e_input[997]), .Z(n12635) );
  XNOR U13660 ( .A(n12625), .B(n12636), .Z(n12627) );
  XOR U13661 ( .A(n12637), .B(n12638), .Z(n12625) );
  AND U13662 ( .A(n12639), .B(n12640), .Z(n12638) );
  XNOR U13663 ( .A(n12641), .B(n12637), .Z(n12640) );
  XOR U13664 ( .A(n12642), .B(e_input[997]), .Z(n12633) );
  IV U13665 ( .A(n12631), .Z(n12642) );
  XOR U13666 ( .A(n12643), .B(n12644), .Z(n12631) );
  AND U13667 ( .A(n12645), .B(n12646), .Z(n12644) );
  XNOR U13668 ( .A(n12643), .B(n6324), .Z(n12646) );
  XNOR U13669 ( .A(n12639), .B(n12641), .Z(n6324) );
  NAND U13670 ( .A(n12647), .B(e_input[996]), .Z(n12641) );
  NAND U13671 ( .A(n12323), .B(e_input[996]), .Z(n12647) );
  XNOR U13672 ( .A(n12637), .B(n12648), .Z(n12639) );
  XOR U13673 ( .A(n12649), .B(n12650), .Z(n12637) );
  AND U13674 ( .A(n12651), .B(n12652), .Z(n12650) );
  XNOR U13675 ( .A(n12653), .B(n12649), .Z(n12652) );
  XOR U13676 ( .A(n12654), .B(e_input[996]), .Z(n12645) );
  IV U13677 ( .A(n12643), .Z(n12654) );
  XOR U13678 ( .A(n12655), .B(n12656), .Z(n12643) );
  AND U13679 ( .A(n12657), .B(n12658), .Z(n12656) );
  XNOR U13680 ( .A(n12655), .B(n6330), .Z(n12658) );
  XNOR U13681 ( .A(n12651), .B(n12653), .Z(n6330) );
  NAND U13682 ( .A(n12659), .B(e_input[995]), .Z(n12653) );
  NAND U13683 ( .A(n12323), .B(e_input[995]), .Z(n12659) );
  XNOR U13684 ( .A(n12649), .B(n12660), .Z(n12651) );
  XOR U13685 ( .A(n12661), .B(n12662), .Z(n12649) );
  AND U13686 ( .A(n12663), .B(n12664), .Z(n12662) );
  XNOR U13687 ( .A(n12665), .B(n12661), .Z(n12664) );
  XOR U13688 ( .A(n12666), .B(e_input[995]), .Z(n12657) );
  IV U13689 ( .A(n12655), .Z(n12666) );
  XOR U13690 ( .A(n12667), .B(n12668), .Z(n12655) );
  AND U13691 ( .A(n12669), .B(n12670), .Z(n12668) );
  XNOR U13692 ( .A(n12667), .B(n6336), .Z(n12670) );
  XNOR U13693 ( .A(n12663), .B(n12665), .Z(n6336) );
  NAND U13694 ( .A(n12671), .B(e_input[994]), .Z(n12665) );
  NAND U13695 ( .A(n12323), .B(e_input[994]), .Z(n12671) );
  XNOR U13696 ( .A(n12661), .B(n12672), .Z(n12663) );
  XOR U13697 ( .A(n12673), .B(n12674), .Z(n12661) );
  AND U13698 ( .A(n12675), .B(n12676), .Z(n12674) );
  XNOR U13699 ( .A(n12677), .B(n12673), .Z(n12676) );
  XOR U13700 ( .A(n12678), .B(e_input[994]), .Z(n12669) );
  IV U13701 ( .A(n12667), .Z(n12678) );
  XOR U13702 ( .A(n12679), .B(n12680), .Z(n12667) );
  AND U13703 ( .A(n12681), .B(n12682), .Z(n12680) );
  XNOR U13704 ( .A(n12679), .B(n6342), .Z(n12682) );
  XNOR U13705 ( .A(n12675), .B(n12677), .Z(n6342) );
  NAND U13706 ( .A(n12683), .B(e_input[993]), .Z(n12677) );
  NAND U13707 ( .A(n12323), .B(e_input[993]), .Z(n12683) );
  XNOR U13708 ( .A(n12673), .B(n12684), .Z(n12675) );
  XOR U13709 ( .A(n12685), .B(n12686), .Z(n12673) );
  AND U13710 ( .A(n12687), .B(n12688), .Z(n12686) );
  XNOR U13711 ( .A(n12689), .B(n12685), .Z(n12688) );
  XOR U13712 ( .A(n12690), .B(e_input[993]), .Z(n12681) );
  IV U13713 ( .A(n12679), .Z(n12690) );
  XOR U13714 ( .A(n12691), .B(n12692), .Z(n12679) );
  AND U13715 ( .A(n12693), .B(n12694), .Z(n12692) );
  XNOR U13716 ( .A(n12691), .B(n6348), .Z(n12694) );
  XNOR U13717 ( .A(n12687), .B(n12689), .Z(n6348) );
  NAND U13718 ( .A(n12695), .B(e_input[992]), .Z(n12689) );
  NAND U13719 ( .A(n12323), .B(e_input[992]), .Z(n12695) );
  XNOR U13720 ( .A(n12685), .B(n12696), .Z(n12687) );
  XOR U13721 ( .A(n12697), .B(n12698), .Z(n12685) );
  AND U13722 ( .A(n12699), .B(n12700), .Z(n12698) );
  XNOR U13723 ( .A(n12701), .B(n12697), .Z(n12700) );
  XOR U13724 ( .A(n12702), .B(e_input[992]), .Z(n12693) );
  IV U13725 ( .A(n12691), .Z(n12702) );
  XOR U13726 ( .A(n12703), .B(n12704), .Z(n12691) );
  AND U13727 ( .A(n12705), .B(n12706), .Z(n12704) );
  XNOR U13728 ( .A(n12703), .B(n6354), .Z(n12706) );
  XNOR U13729 ( .A(n12699), .B(n12701), .Z(n6354) );
  NAND U13730 ( .A(n12707), .B(e_input[991]), .Z(n12701) );
  NAND U13731 ( .A(n12323), .B(e_input[991]), .Z(n12707) );
  XNOR U13732 ( .A(n12697), .B(n12708), .Z(n12699) );
  XOR U13733 ( .A(n12709), .B(n12710), .Z(n12697) );
  AND U13734 ( .A(n12711), .B(n12712), .Z(n12710) );
  XNOR U13735 ( .A(n12713), .B(n12709), .Z(n12712) );
  XOR U13736 ( .A(n12714), .B(e_input[991]), .Z(n12705) );
  IV U13737 ( .A(n12703), .Z(n12714) );
  XOR U13738 ( .A(n12715), .B(n12716), .Z(n12703) );
  AND U13739 ( .A(n12717), .B(n12718), .Z(n12716) );
  XNOR U13740 ( .A(n12715), .B(n6360), .Z(n12718) );
  XNOR U13741 ( .A(n12711), .B(n12713), .Z(n6360) );
  NAND U13742 ( .A(n12719), .B(e_input[990]), .Z(n12713) );
  NAND U13743 ( .A(n12323), .B(e_input[990]), .Z(n12719) );
  XNOR U13744 ( .A(n12709), .B(n12720), .Z(n12711) );
  XOR U13745 ( .A(n12721), .B(n12722), .Z(n12709) );
  AND U13746 ( .A(n12723), .B(n12724), .Z(n12722) );
  XNOR U13747 ( .A(n12725), .B(n12721), .Z(n12724) );
  XOR U13748 ( .A(n12726), .B(e_input[990]), .Z(n12717) );
  IV U13749 ( .A(n12715), .Z(n12726) );
  XOR U13750 ( .A(n12727), .B(n12728), .Z(n12715) );
  AND U13751 ( .A(n12729), .B(n12730), .Z(n12728) );
  XNOR U13752 ( .A(n12727), .B(n6366), .Z(n12730) );
  XNOR U13753 ( .A(n12723), .B(n12725), .Z(n6366) );
  NAND U13754 ( .A(n12731), .B(e_input[989]), .Z(n12725) );
  NAND U13755 ( .A(n12323), .B(e_input[989]), .Z(n12731) );
  XNOR U13756 ( .A(n12721), .B(n12732), .Z(n12723) );
  XOR U13757 ( .A(n12733), .B(n12734), .Z(n12721) );
  AND U13758 ( .A(n12735), .B(n12736), .Z(n12734) );
  XNOR U13759 ( .A(n12737), .B(n12733), .Z(n12736) );
  XOR U13760 ( .A(n12738), .B(e_input[989]), .Z(n12729) );
  IV U13761 ( .A(n12727), .Z(n12738) );
  XOR U13762 ( .A(n12739), .B(n12740), .Z(n12727) );
  AND U13763 ( .A(n12741), .B(n12742), .Z(n12740) );
  XNOR U13764 ( .A(n12739), .B(n6372), .Z(n12742) );
  XNOR U13765 ( .A(n12735), .B(n12737), .Z(n6372) );
  NAND U13766 ( .A(n12743), .B(e_input[988]), .Z(n12737) );
  NAND U13767 ( .A(n12323), .B(e_input[988]), .Z(n12743) );
  XNOR U13768 ( .A(n12733), .B(n12744), .Z(n12735) );
  XOR U13769 ( .A(n12745), .B(n12746), .Z(n12733) );
  AND U13770 ( .A(n12747), .B(n12748), .Z(n12746) );
  XNOR U13771 ( .A(n12749), .B(n12745), .Z(n12748) );
  XOR U13772 ( .A(n12750), .B(e_input[988]), .Z(n12741) );
  IV U13773 ( .A(n12739), .Z(n12750) );
  XOR U13774 ( .A(n12751), .B(n12752), .Z(n12739) );
  AND U13775 ( .A(n12753), .B(n12754), .Z(n12752) );
  XNOR U13776 ( .A(n12751), .B(n6378), .Z(n12754) );
  XNOR U13777 ( .A(n12747), .B(n12749), .Z(n6378) );
  NAND U13778 ( .A(n12755), .B(e_input[987]), .Z(n12749) );
  NAND U13779 ( .A(n12323), .B(e_input[987]), .Z(n12755) );
  XNOR U13780 ( .A(n12745), .B(n12756), .Z(n12747) );
  XOR U13781 ( .A(n12757), .B(n12758), .Z(n12745) );
  AND U13782 ( .A(n12759), .B(n12760), .Z(n12758) );
  XNOR U13783 ( .A(n12761), .B(n12757), .Z(n12760) );
  XOR U13784 ( .A(n12762), .B(e_input[987]), .Z(n12753) );
  IV U13785 ( .A(n12751), .Z(n12762) );
  XOR U13786 ( .A(n12763), .B(n12764), .Z(n12751) );
  AND U13787 ( .A(n12765), .B(n12766), .Z(n12764) );
  XNOR U13788 ( .A(n12763), .B(n6384), .Z(n12766) );
  XNOR U13789 ( .A(n12759), .B(n12761), .Z(n6384) );
  NAND U13790 ( .A(n12767), .B(e_input[986]), .Z(n12761) );
  NAND U13791 ( .A(n12323), .B(e_input[986]), .Z(n12767) );
  XNOR U13792 ( .A(n12757), .B(n12768), .Z(n12759) );
  XOR U13793 ( .A(n12769), .B(n12770), .Z(n12757) );
  AND U13794 ( .A(n12771), .B(n12772), .Z(n12770) );
  XNOR U13795 ( .A(n12773), .B(n12769), .Z(n12772) );
  XOR U13796 ( .A(n12774), .B(e_input[986]), .Z(n12765) );
  IV U13797 ( .A(n12763), .Z(n12774) );
  XOR U13798 ( .A(n12775), .B(n12776), .Z(n12763) );
  AND U13799 ( .A(n12777), .B(n12778), .Z(n12776) );
  XNOR U13800 ( .A(n12775), .B(n6390), .Z(n12778) );
  XNOR U13801 ( .A(n12771), .B(n12773), .Z(n6390) );
  NAND U13802 ( .A(n12779), .B(e_input[985]), .Z(n12773) );
  NAND U13803 ( .A(n12323), .B(e_input[985]), .Z(n12779) );
  XNOR U13804 ( .A(n12769), .B(n12780), .Z(n12771) );
  XOR U13805 ( .A(n12781), .B(n12782), .Z(n12769) );
  AND U13806 ( .A(n12783), .B(n12784), .Z(n12782) );
  XNOR U13807 ( .A(n12785), .B(n12781), .Z(n12784) );
  XOR U13808 ( .A(n12786), .B(e_input[985]), .Z(n12777) );
  IV U13809 ( .A(n12775), .Z(n12786) );
  XOR U13810 ( .A(n12787), .B(n12788), .Z(n12775) );
  AND U13811 ( .A(n12789), .B(n12790), .Z(n12788) );
  XNOR U13812 ( .A(n12787), .B(n6396), .Z(n12790) );
  XNOR U13813 ( .A(n12783), .B(n12785), .Z(n6396) );
  NAND U13814 ( .A(n12791), .B(e_input[984]), .Z(n12785) );
  NAND U13815 ( .A(n12323), .B(e_input[984]), .Z(n12791) );
  XNOR U13816 ( .A(n12781), .B(n12792), .Z(n12783) );
  XOR U13817 ( .A(n12793), .B(n12794), .Z(n12781) );
  AND U13818 ( .A(n12795), .B(n12796), .Z(n12794) );
  XNOR U13819 ( .A(n12797), .B(n12793), .Z(n12796) );
  XOR U13820 ( .A(n12798), .B(e_input[984]), .Z(n12789) );
  IV U13821 ( .A(n12787), .Z(n12798) );
  XOR U13822 ( .A(n12799), .B(n12800), .Z(n12787) );
  AND U13823 ( .A(n12801), .B(n12802), .Z(n12800) );
  XNOR U13824 ( .A(n12799), .B(n6402), .Z(n12802) );
  XNOR U13825 ( .A(n12795), .B(n12797), .Z(n6402) );
  NAND U13826 ( .A(n12803), .B(e_input[983]), .Z(n12797) );
  NAND U13827 ( .A(n12323), .B(e_input[983]), .Z(n12803) );
  XNOR U13828 ( .A(n12793), .B(n12804), .Z(n12795) );
  XOR U13829 ( .A(n12805), .B(n12806), .Z(n12793) );
  AND U13830 ( .A(n12807), .B(n12808), .Z(n12806) );
  XNOR U13831 ( .A(n12809), .B(n12805), .Z(n12808) );
  XOR U13832 ( .A(n12810), .B(e_input[983]), .Z(n12801) );
  IV U13833 ( .A(n12799), .Z(n12810) );
  XOR U13834 ( .A(n12811), .B(n12812), .Z(n12799) );
  AND U13835 ( .A(n12813), .B(n12814), .Z(n12812) );
  XNOR U13836 ( .A(n12811), .B(n6408), .Z(n12814) );
  XNOR U13837 ( .A(n12807), .B(n12809), .Z(n6408) );
  NAND U13838 ( .A(n12815), .B(e_input[982]), .Z(n12809) );
  NAND U13839 ( .A(n12323), .B(e_input[982]), .Z(n12815) );
  XNOR U13840 ( .A(n12805), .B(n12816), .Z(n12807) );
  XOR U13841 ( .A(n12817), .B(n12818), .Z(n12805) );
  AND U13842 ( .A(n12819), .B(n12820), .Z(n12818) );
  XNOR U13843 ( .A(n12821), .B(n12817), .Z(n12820) );
  XOR U13844 ( .A(n12822), .B(e_input[982]), .Z(n12813) );
  IV U13845 ( .A(n12811), .Z(n12822) );
  XOR U13846 ( .A(n12823), .B(n12824), .Z(n12811) );
  AND U13847 ( .A(n12825), .B(n12826), .Z(n12824) );
  XNOR U13848 ( .A(n12823), .B(n6414), .Z(n12826) );
  XNOR U13849 ( .A(n12819), .B(n12821), .Z(n6414) );
  NAND U13850 ( .A(n12827), .B(e_input[981]), .Z(n12821) );
  NAND U13851 ( .A(n12323), .B(e_input[981]), .Z(n12827) );
  XNOR U13852 ( .A(n12817), .B(n12828), .Z(n12819) );
  XOR U13853 ( .A(n12829), .B(n12830), .Z(n12817) );
  AND U13854 ( .A(n12831), .B(n12832), .Z(n12830) );
  XNOR U13855 ( .A(n12833), .B(n12829), .Z(n12832) );
  XOR U13856 ( .A(n12834), .B(e_input[981]), .Z(n12825) );
  IV U13857 ( .A(n12823), .Z(n12834) );
  XOR U13858 ( .A(n12835), .B(n12836), .Z(n12823) );
  AND U13859 ( .A(n12837), .B(n12838), .Z(n12836) );
  XNOR U13860 ( .A(n12835), .B(n6420), .Z(n12838) );
  XNOR U13861 ( .A(n12831), .B(n12833), .Z(n6420) );
  NAND U13862 ( .A(n12839), .B(e_input[980]), .Z(n12833) );
  NAND U13863 ( .A(n12323), .B(e_input[980]), .Z(n12839) );
  XNOR U13864 ( .A(n12829), .B(n12840), .Z(n12831) );
  XOR U13865 ( .A(n12841), .B(n12842), .Z(n12829) );
  AND U13866 ( .A(n12843), .B(n12844), .Z(n12842) );
  XNOR U13867 ( .A(n12845), .B(n12841), .Z(n12844) );
  XOR U13868 ( .A(n12846), .B(e_input[980]), .Z(n12837) );
  IV U13869 ( .A(n12835), .Z(n12846) );
  XOR U13870 ( .A(n12847), .B(n12848), .Z(n12835) );
  AND U13871 ( .A(n12849), .B(n12850), .Z(n12848) );
  XNOR U13872 ( .A(n12847), .B(n6426), .Z(n12850) );
  XNOR U13873 ( .A(n12843), .B(n12845), .Z(n6426) );
  NAND U13874 ( .A(n12851), .B(e_input[979]), .Z(n12845) );
  NAND U13875 ( .A(n12323), .B(e_input[979]), .Z(n12851) );
  XNOR U13876 ( .A(n12841), .B(n12852), .Z(n12843) );
  XOR U13877 ( .A(n12853), .B(n12854), .Z(n12841) );
  AND U13878 ( .A(n12855), .B(n12856), .Z(n12854) );
  XNOR U13879 ( .A(n12857), .B(n12853), .Z(n12856) );
  XOR U13880 ( .A(n12858), .B(e_input[979]), .Z(n12849) );
  IV U13881 ( .A(n12847), .Z(n12858) );
  XOR U13882 ( .A(n12859), .B(n12860), .Z(n12847) );
  AND U13883 ( .A(n12861), .B(n12862), .Z(n12860) );
  XNOR U13884 ( .A(n12859), .B(n6432), .Z(n12862) );
  XNOR U13885 ( .A(n12855), .B(n12857), .Z(n6432) );
  NAND U13886 ( .A(n12863), .B(e_input[978]), .Z(n12857) );
  NAND U13887 ( .A(n12323), .B(e_input[978]), .Z(n12863) );
  XNOR U13888 ( .A(n12853), .B(n12864), .Z(n12855) );
  XOR U13889 ( .A(n12865), .B(n12866), .Z(n12853) );
  AND U13890 ( .A(n12867), .B(n12868), .Z(n12866) );
  XNOR U13891 ( .A(n12869), .B(n12865), .Z(n12868) );
  XOR U13892 ( .A(n12870), .B(e_input[978]), .Z(n12861) );
  IV U13893 ( .A(n12859), .Z(n12870) );
  XOR U13894 ( .A(n12871), .B(n12872), .Z(n12859) );
  AND U13895 ( .A(n12873), .B(n12874), .Z(n12872) );
  XNOR U13896 ( .A(n12871), .B(n6438), .Z(n12874) );
  XNOR U13897 ( .A(n12867), .B(n12869), .Z(n6438) );
  NAND U13898 ( .A(n12875), .B(e_input[977]), .Z(n12869) );
  NAND U13899 ( .A(n12323), .B(e_input[977]), .Z(n12875) );
  XNOR U13900 ( .A(n12865), .B(n12876), .Z(n12867) );
  XOR U13901 ( .A(n12877), .B(n12878), .Z(n12865) );
  AND U13902 ( .A(n12879), .B(n12880), .Z(n12878) );
  XNOR U13903 ( .A(n12881), .B(n12877), .Z(n12880) );
  XOR U13904 ( .A(n12882), .B(e_input[977]), .Z(n12873) );
  IV U13905 ( .A(n12871), .Z(n12882) );
  XOR U13906 ( .A(n12883), .B(n12884), .Z(n12871) );
  AND U13907 ( .A(n12885), .B(n12886), .Z(n12884) );
  XNOR U13908 ( .A(n12883), .B(n6444), .Z(n12886) );
  XNOR U13909 ( .A(n12879), .B(n12881), .Z(n6444) );
  NAND U13910 ( .A(n12887), .B(e_input[976]), .Z(n12881) );
  NAND U13911 ( .A(n12323), .B(e_input[976]), .Z(n12887) );
  XNOR U13912 ( .A(n12877), .B(n12888), .Z(n12879) );
  XOR U13913 ( .A(n12889), .B(n12890), .Z(n12877) );
  AND U13914 ( .A(n12891), .B(n12892), .Z(n12890) );
  XNOR U13915 ( .A(n12893), .B(n12889), .Z(n12892) );
  XOR U13916 ( .A(n12894), .B(e_input[976]), .Z(n12885) );
  IV U13917 ( .A(n12883), .Z(n12894) );
  XOR U13918 ( .A(n12895), .B(n12896), .Z(n12883) );
  AND U13919 ( .A(n12897), .B(n12898), .Z(n12896) );
  XNOR U13920 ( .A(n12895), .B(n6450), .Z(n12898) );
  XNOR U13921 ( .A(n12891), .B(n12893), .Z(n6450) );
  NAND U13922 ( .A(n12899), .B(e_input[975]), .Z(n12893) );
  NAND U13923 ( .A(n12323), .B(e_input[975]), .Z(n12899) );
  XNOR U13924 ( .A(n12889), .B(n12900), .Z(n12891) );
  XOR U13925 ( .A(n12901), .B(n12902), .Z(n12889) );
  AND U13926 ( .A(n12903), .B(n12904), .Z(n12902) );
  XNOR U13927 ( .A(n12905), .B(n12901), .Z(n12904) );
  XOR U13928 ( .A(n12906), .B(e_input[975]), .Z(n12897) );
  IV U13929 ( .A(n12895), .Z(n12906) );
  XOR U13930 ( .A(n12907), .B(n12908), .Z(n12895) );
  AND U13931 ( .A(n12909), .B(n12910), .Z(n12908) );
  XNOR U13932 ( .A(n12907), .B(n6456), .Z(n12910) );
  XNOR U13933 ( .A(n12903), .B(n12905), .Z(n6456) );
  NAND U13934 ( .A(n12911), .B(e_input[974]), .Z(n12905) );
  NAND U13935 ( .A(n12323), .B(e_input[974]), .Z(n12911) );
  XNOR U13936 ( .A(n12901), .B(n12912), .Z(n12903) );
  XOR U13937 ( .A(n12913), .B(n12914), .Z(n12901) );
  AND U13938 ( .A(n12915), .B(n12916), .Z(n12914) );
  XNOR U13939 ( .A(n12917), .B(n12913), .Z(n12916) );
  XOR U13940 ( .A(n12918), .B(e_input[974]), .Z(n12909) );
  IV U13941 ( .A(n12907), .Z(n12918) );
  XOR U13942 ( .A(n12919), .B(n12920), .Z(n12907) );
  AND U13943 ( .A(n12921), .B(n12922), .Z(n12920) );
  XNOR U13944 ( .A(n12919), .B(n6462), .Z(n12922) );
  XNOR U13945 ( .A(n12915), .B(n12917), .Z(n6462) );
  NAND U13946 ( .A(n12923), .B(e_input[973]), .Z(n12917) );
  NAND U13947 ( .A(n12323), .B(e_input[973]), .Z(n12923) );
  XNOR U13948 ( .A(n12913), .B(n12924), .Z(n12915) );
  XOR U13949 ( .A(n12925), .B(n12926), .Z(n12913) );
  AND U13950 ( .A(n12927), .B(n12928), .Z(n12926) );
  XNOR U13951 ( .A(n12929), .B(n12925), .Z(n12928) );
  XOR U13952 ( .A(n12930), .B(e_input[973]), .Z(n12921) );
  IV U13953 ( .A(n12919), .Z(n12930) );
  XOR U13954 ( .A(n12931), .B(n12932), .Z(n12919) );
  AND U13955 ( .A(n12933), .B(n12934), .Z(n12932) );
  XNOR U13956 ( .A(n12931), .B(n6468), .Z(n12934) );
  XNOR U13957 ( .A(n12927), .B(n12929), .Z(n6468) );
  NAND U13958 ( .A(n12935), .B(e_input[972]), .Z(n12929) );
  NAND U13959 ( .A(n12323), .B(e_input[972]), .Z(n12935) );
  XNOR U13960 ( .A(n12925), .B(n12936), .Z(n12927) );
  XOR U13961 ( .A(n12937), .B(n12938), .Z(n12925) );
  AND U13962 ( .A(n12939), .B(n12940), .Z(n12938) );
  XNOR U13963 ( .A(n12941), .B(n12937), .Z(n12940) );
  XOR U13964 ( .A(n12942), .B(e_input[972]), .Z(n12933) );
  IV U13965 ( .A(n12931), .Z(n12942) );
  XOR U13966 ( .A(n12943), .B(n12944), .Z(n12931) );
  AND U13967 ( .A(n12945), .B(n12946), .Z(n12944) );
  XNOR U13968 ( .A(n12943), .B(n6474), .Z(n12946) );
  XNOR U13969 ( .A(n12939), .B(n12941), .Z(n6474) );
  NAND U13970 ( .A(n12947), .B(e_input[971]), .Z(n12941) );
  NAND U13971 ( .A(n12323), .B(e_input[971]), .Z(n12947) );
  XNOR U13972 ( .A(n12937), .B(n12948), .Z(n12939) );
  XOR U13973 ( .A(n12949), .B(n12950), .Z(n12937) );
  AND U13974 ( .A(n12951), .B(n12952), .Z(n12950) );
  XNOR U13975 ( .A(n12953), .B(n12949), .Z(n12952) );
  XOR U13976 ( .A(n12954), .B(e_input[971]), .Z(n12945) );
  IV U13977 ( .A(n12943), .Z(n12954) );
  XOR U13978 ( .A(n12955), .B(n12956), .Z(n12943) );
  AND U13979 ( .A(n12957), .B(n12958), .Z(n12956) );
  XNOR U13980 ( .A(n12955), .B(n6480), .Z(n12958) );
  XNOR U13981 ( .A(n12951), .B(n12953), .Z(n6480) );
  NAND U13982 ( .A(n12959), .B(e_input[970]), .Z(n12953) );
  NAND U13983 ( .A(n12323), .B(e_input[970]), .Z(n12959) );
  XNOR U13984 ( .A(n12949), .B(n12960), .Z(n12951) );
  XOR U13985 ( .A(n12961), .B(n12962), .Z(n12949) );
  AND U13986 ( .A(n12963), .B(n12964), .Z(n12962) );
  XNOR U13987 ( .A(n12965), .B(n12961), .Z(n12964) );
  XOR U13988 ( .A(n12966), .B(e_input[970]), .Z(n12957) );
  IV U13989 ( .A(n12955), .Z(n12966) );
  XOR U13990 ( .A(n12967), .B(n12968), .Z(n12955) );
  AND U13991 ( .A(n12969), .B(n12970), .Z(n12968) );
  XNOR U13992 ( .A(n12967), .B(n6486), .Z(n12970) );
  XNOR U13993 ( .A(n12963), .B(n12965), .Z(n6486) );
  NAND U13994 ( .A(n12971), .B(e_input[969]), .Z(n12965) );
  NAND U13995 ( .A(n12323), .B(e_input[969]), .Z(n12971) );
  XNOR U13996 ( .A(n12961), .B(n12972), .Z(n12963) );
  XOR U13997 ( .A(n12973), .B(n12974), .Z(n12961) );
  AND U13998 ( .A(n12975), .B(n12976), .Z(n12974) );
  XNOR U13999 ( .A(n12977), .B(n12973), .Z(n12976) );
  XOR U14000 ( .A(n12978), .B(e_input[969]), .Z(n12969) );
  IV U14001 ( .A(n12967), .Z(n12978) );
  XOR U14002 ( .A(n12979), .B(n12980), .Z(n12967) );
  AND U14003 ( .A(n12981), .B(n12982), .Z(n12980) );
  XNOR U14004 ( .A(n12979), .B(n6492), .Z(n12982) );
  XNOR U14005 ( .A(n12975), .B(n12977), .Z(n6492) );
  NAND U14006 ( .A(n12983), .B(e_input[968]), .Z(n12977) );
  NAND U14007 ( .A(n12323), .B(e_input[968]), .Z(n12983) );
  XNOR U14008 ( .A(n12973), .B(n12984), .Z(n12975) );
  XOR U14009 ( .A(n12985), .B(n12986), .Z(n12973) );
  AND U14010 ( .A(n12987), .B(n12988), .Z(n12986) );
  XNOR U14011 ( .A(n12989), .B(n12985), .Z(n12988) );
  XOR U14012 ( .A(n12990), .B(e_input[968]), .Z(n12981) );
  IV U14013 ( .A(n12979), .Z(n12990) );
  XOR U14014 ( .A(n12991), .B(n12992), .Z(n12979) );
  AND U14015 ( .A(n12993), .B(n12994), .Z(n12992) );
  XNOR U14016 ( .A(n12991), .B(n6498), .Z(n12994) );
  XNOR U14017 ( .A(n12987), .B(n12989), .Z(n6498) );
  NAND U14018 ( .A(n12995), .B(e_input[967]), .Z(n12989) );
  NAND U14019 ( .A(n12323), .B(e_input[967]), .Z(n12995) );
  XNOR U14020 ( .A(n12985), .B(n12996), .Z(n12987) );
  XOR U14021 ( .A(n12997), .B(n12998), .Z(n12985) );
  AND U14022 ( .A(n12999), .B(n13000), .Z(n12998) );
  XNOR U14023 ( .A(n13001), .B(n12997), .Z(n13000) );
  XOR U14024 ( .A(n13002), .B(e_input[967]), .Z(n12993) );
  IV U14025 ( .A(n12991), .Z(n13002) );
  XOR U14026 ( .A(n13003), .B(n13004), .Z(n12991) );
  AND U14027 ( .A(n13005), .B(n13006), .Z(n13004) );
  XNOR U14028 ( .A(n13003), .B(n6504), .Z(n13006) );
  XNOR U14029 ( .A(n12999), .B(n13001), .Z(n6504) );
  NAND U14030 ( .A(n13007), .B(e_input[966]), .Z(n13001) );
  NAND U14031 ( .A(n12323), .B(e_input[966]), .Z(n13007) );
  XNOR U14032 ( .A(n12997), .B(n13008), .Z(n12999) );
  XOR U14033 ( .A(n13009), .B(n13010), .Z(n12997) );
  AND U14034 ( .A(n13011), .B(n13012), .Z(n13010) );
  XNOR U14035 ( .A(n13013), .B(n13009), .Z(n13012) );
  XOR U14036 ( .A(n13014), .B(e_input[966]), .Z(n13005) );
  IV U14037 ( .A(n13003), .Z(n13014) );
  XOR U14038 ( .A(n13015), .B(n13016), .Z(n13003) );
  AND U14039 ( .A(n13017), .B(n13018), .Z(n13016) );
  XNOR U14040 ( .A(n13015), .B(n6510), .Z(n13018) );
  XNOR U14041 ( .A(n13011), .B(n13013), .Z(n6510) );
  NAND U14042 ( .A(n13019), .B(e_input[965]), .Z(n13013) );
  NAND U14043 ( .A(n12323), .B(e_input[965]), .Z(n13019) );
  XNOR U14044 ( .A(n13009), .B(n13020), .Z(n13011) );
  XOR U14045 ( .A(n13021), .B(n13022), .Z(n13009) );
  AND U14046 ( .A(n13023), .B(n13024), .Z(n13022) );
  XNOR U14047 ( .A(n13025), .B(n13021), .Z(n13024) );
  XOR U14048 ( .A(n13026), .B(e_input[965]), .Z(n13017) );
  IV U14049 ( .A(n13015), .Z(n13026) );
  XOR U14050 ( .A(n13027), .B(n13028), .Z(n13015) );
  AND U14051 ( .A(n13029), .B(n13030), .Z(n13028) );
  XNOR U14052 ( .A(n13027), .B(n6516), .Z(n13030) );
  XNOR U14053 ( .A(n13023), .B(n13025), .Z(n6516) );
  NAND U14054 ( .A(n13031), .B(e_input[964]), .Z(n13025) );
  NAND U14055 ( .A(n12323), .B(e_input[964]), .Z(n13031) );
  XNOR U14056 ( .A(n13021), .B(n13032), .Z(n13023) );
  XOR U14057 ( .A(n13033), .B(n13034), .Z(n13021) );
  AND U14058 ( .A(n13035), .B(n13036), .Z(n13034) );
  XNOR U14059 ( .A(n13037), .B(n13033), .Z(n13036) );
  XOR U14060 ( .A(n13038), .B(e_input[964]), .Z(n13029) );
  IV U14061 ( .A(n13027), .Z(n13038) );
  XOR U14062 ( .A(n13039), .B(n13040), .Z(n13027) );
  AND U14063 ( .A(n13041), .B(n13042), .Z(n13040) );
  XNOR U14064 ( .A(n13039), .B(n6522), .Z(n13042) );
  XNOR U14065 ( .A(n13035), .B(n13037), .Z(n6522) );
  NAND U14066 ( .A(n13043), .B(e_input[963]), .Z(n13037) );
  NAND U14067 ( .A(n12323), .B(e_input[963]), .Z(n13043) );
  XNOR U14068 ( .A(n13033), .B(n13044), .Z(n13035) );
  XOR U14069 ( .A(n13045), .B(n13046), .Z(n13033) );
  AND U14070 ( .A(n13047), .B(n13048), .Z(n13046) );
  XNOR U14071 ( .A(n13049), .B(n13045), .Z(n13048) );
  XOR U14072 ( .A(n13050), .B(e_input[963]), .Z(n13041) );
  IV U14073 ( .A(n13039), .Z(n13050) );
  XOR U14074 ( .A(n13051), .B(n13052), .Z(n13039) );
  AND U14075 ( .A(n13053), .B(n13054), .Z(n13052) );
  XNOR U14076 ( .A(n13051), .B(n6528), .Z(n13054) );
  XNOR U14077 ( .A(n13047), .B(n13049), .Z(n6528) );
  NAND U14078 ( .A(n13055), .B(e_input[962]), .Z(n13049) );
  NAND U14079 ( .A(n12323), .B(e_input[962]), .Z(n13055) );
  XNOR U14080 ( .A(n13045), .B(n13056), .Z(n13047) );
  XOR U14081 ( .A(n13057), .B(n13058), .Z(n13045) );
  AND U14082 ( .A(n13059), .B(n13060), .Z(n13058) );
  XNOR U14083 ( .A(n13061), .B(n13057), .Z(n13060) );
  XOR U14084 ( .A(n13062), .B(e_input[962]), .Z(n13053) );
  IV U14085 ( .A(n13051), .Z(n13062) );
  XOR U14086 ( .A(n13063), .B(n13064), .Z(n13051) );
  AND U14087 ( .A(n13065), .B(n13066), .Z(n13064) );
  XNOR U14088 ( .A(n13063), .B(n6534), .Z(n13066) );
  XNOR U14089 ( .A(n13059), .B(n13061), .Z(n6534) );
  NAND U14090 ( .A(n13067), .B(e_input[961]), .Z(n13061) );
  NAND U14091 ( .A(n12323), .B(e_input[961]), .Z(n13067) );
  XNOR U14092 ( .A(n13057), .B(n13068), .Z(n13059) );
  XOR U14093 ( .A(n13069), .B(n13070), .Z(n13057) );
  AND U14094 ( .A(n13071), .B(n13072), .Z(n13070) );
  XNOR U14095 ( .A(n13073), .B(n13069), .Z(n13072) );
  XOR U14096 ( .A(n13074), .B(e_input[961]), .Z(n13065) );
  IV U14097 ( .A(n13063), .Z(n13074) );
  XOR U14098 ( .A(n13075), .B(n13076), .Z(n13063) );
  AND U14099 ( .A(n13077), .B(n13078), .Z(n13076) );
  XNOR U14100 ( .A(n13075), .B(n6540), .Z(n13078) );
  XNOR U14101 ( .A(n13071), .B(n13073), .Z(n6540) );
  NAND U14102 ( .A(n13079), .B(e_input[960]), .Z(n13073) );
  NAND U14103 ( .A(n12323), .B(e_input[960]), .Z(n13079) );
  XNOR U14104 ( .A(n13069), .B(n13080), .Z(n13071) );
  XOR U14105 ( .A(n13081), .B(n13082), .Z(n13069) );
  AND U14106 ( .A(n13083), .B(n13084), .Z(n13082) );
  XNOR U14107 ( .A(n13085), .B(n13081), .Z(n13084) );
  XOR U14108 ( .A(n13086), .B(e_input[960]), .Z(n13077) );
  IV U14109 ( .A(n13075), .Z(n13086) );
  XOR U14110 ( .A(n13087), .B(n13088), .Z(n13075) );
  AND U14111 ( .A(n13089), .B(n13090), .Z(n13088) );
  XNOR U14112 ( .A(n13087), .B(n6546), .Z(n13090) );
  XNOR U14113 ( .A(n13083), .B(n13085), .Z(n6546) );
  NAND U14114 ( .A(n13091), .B(e_input[959]), .Z(n13085) );
  NAND U14115 ( .A(n12323), .B(e_input[959]), .Z(n13091) );
  XNOR U14116 ( .A(n13081), .B(n13092), .Z(n13083) );
  XOR U14117 ( .A(n13093), .B(n13094), .Z(n13081) );
  AND U14118 ( .A(n13095), .B(n13096), .Z(n13094) );
  XNOR U14119 ( .A(n13097), .B(n13093), .Z(n13096) );
  XOR U14120 ( .A(n13098), .B(e_input[959]), .Z(n13089) );
  IV U14121 ( .A(n13087), .Z(n13098) );
  XOR U14122 ( .A(n13099), .B(n13100), .Z(n13087) );
  AND U14123 ( .A(n13101), .B(n13102), .Z(n13100) );
  XNOR U14124 ( .A(n13099), .B(n6552), .Z(n13102) );
  XNOR U14125 ( .A(n13095), .B(n13097), .Z(n6552) );
  NAND U14126 ( .A(n13103), .B(e_input[958]), .Z(n13097) );
  NAND U14127 ( .A(n12323), .B(e_input[958]), .Z(n13103) );
  XNOR U14128 ( .A(n13093), .B(n13104), .Z(n13095) );
  XOR U14129 ( .A(n13105), .B(n13106), .Z(n13093) );
  AND U14130 ( .A(n13107), .B(n13108), .Z(n13106) );
  XNOR U14131 ( .A(n13109), .B(n13105), .Z(n13108) );
  XOR U14132 ( .A(n13110), .B(e_input[958]), .Z(n13101) );
  IV U14133 ( .A(n13099), .Z(n13110) );
  XOR U14134 ( .A(n13111), .B(n13112), .Z(n13099) );
  AND U14135 ( .A(n13113), .B(n13114), .Z(n13112) );
  XNOR U14136 ( .A(n13111), .B(n6558), .Z(n13114) );
  XNOR U14137 ( .A(n13107), .B(n13109), .Z(n6558) );
  NAND U14138 ( .A(n13115), .B(e_input[957]), .Z(n13109) );
  NAND U14139 ( .A(n12323), .B(e_input[957]), .Z(n13115) );
  XNOR U14140 ( .A(n13105), .B(n13116), .Z(n13107) );
  XOR U14141 ( .A(n13117), .B(n13118), .Z(n13105) );
  AND U14142 ( .A(n13119), .B(n13120), .Z(n13118) );
  XNOR U14143 ( .A(n13121), .B(n13117), .Z(n13120) );
  XOR U14144 ( .A(n13122), .B(e_input[957]), .Z(n13113) );
  IV U14145 ( .A(n13111), .Z(n13122) );
  XOR U14146 ( .A(n13123), .B(n13124), .Z(n13111) );
  AND U14147 ( .A(n13125), .B(n13126), .Z(n13124) );
  XNOR U14148 ( .A(n13123), .B(n6564), .Z(n13126) );
  XNOR U14149 ( .A(n13119), .B(n13121), .Z(n6564) );
  NAND U14150 ( .A(n13127), .B(e_input[956]), .Z(n13121) );
  NAND U14151 ( .A(n12323), .B(e_input[956]), .Z(n13127) );
  XNOR U14152 ( .A(n13117), .B(n13128), .Z(n13119) );
  XOR U14153 ( .A(n13129), .B(n13130), .Z(n13117) );
  AND U14154 ( .A(n13131), .B(n13132), .Z(n13130) );
  XNOR U14155 ( .A(n13133), .B(n13129), .Z(n13132) );
  XOR U14156 ( .A(n13134), .B(e_input[956]), .Z(n13125) );
  IV U14157 ( .A(n13123), .Z(n13134) );
  XOR U14158 ( .A(n13135), .B(n13136), .Z(n13123) );
  AND U14159 ( .A(n13137), .B(n13138), .Z(n13136) );
  XNOR U14160 ( .A(n13135), .B(n6570), .Z(n13138) );
  XNOR U14161 ( .A(n13131), .B(n13133), .Z(n6570) );
  NAND U14162 ( .A(n13139), .B(e_input[955]), .Z(n13133) );
  NAND U14163 ( .A(n12323), .B(e_input[955]), .Z(n13139) );
  XNOR U14164 ( .A(n13129), .B(n13140), .Z(n13131) );
  XOR U14165 ( .A(n13141), .B(n13142), .Z(n13129) );
  AND U14166 ( .A(n13143), .B(n13144), .Z(n13142) );
  XNOR U14167 ( .A(n13145), .B(n13141), .Z(n13144) );
  XOR U14168 ( .A(n13146), .B(e_input[955]), .Z(n13137) );
  IV U14169 ( .A(n13135), .Z(n13146) );
  XOR U14170 ( .A(n13147), .B(n13148), .Z(n13135) );
  AND U14171 ( .A(n13149), .B(n13150), .Z(n13148) );
  XNOR U14172 ( .A(n13147), .B(n6576), .Z(n13150) );
  XNOR U14173 ( .A(n13143), .B(n13145), .Z(n6576) );
  NAND U14174 ( .A(n13151), .B(e_input[954]), .Z(n13145) );
  NAND U14175 ( .A(n12323), .B(e_input[954]), .Z(n13151) );
  XNOR U14176 ( .A(n13141), .B(n13152), .Z(n13143) );
  XOR U14177 ( .A(n13153), .B(n13154), .Z(n13141) );
  AND U14178 ( .A(n13155), .B(n13156), .Z(n13154) );
  XNOR U14179 ( .A(n13157), .B(n13153), .Z(n13156) );
  XOR U14180 ( .A(n13158), .B(e_input[954]), .Z(n13149) );
  IV U14181 ( .A(n13147), .Z(n13158) );
  XOR U14182 ( .A(n13159), .B(n13160), .Z(n13147) );
  AND U14183 ( .A(n13161), .B(n13162), .Z(n13160) );
  XNOR U14184 ( .A(n13159), .B(n6582), .Z(n13162) );
  XNOR U14185 ( .A(n13155), .B(n13157), .Z(n6582) );
  NAND U14186 ( .A(n13163), .B(e_input[953]), .Z(n13157) );
  NAND U14187 ( .A(n12323), .B(e_input[953]), .Z(n13163) );
  XNOR U14188 ( .A(n13153), .B(n13164), .Z(n13155) );
  XOR U14189 ( .A(n13165), .B(n13166), .Z(n13153) );
  AND U14190 ( .A(n13167), .B(n13168), .Z(n13166) );
  XNOR U14191 ( .A(n13169), .B(n13165), .Z(n13168) );
  XOR U14192 ( .A(n13170), .B(e_input[953]), .Z(n13161) );
  IV U14193 ( .A(n13159), .Z(n13170) );
  XOR U14194 ( .A(n13171), .B(n13172), .Z(n13159) );
  AND U14195 ( .A(n13173), .B(n13174), .Z(n13172) );
  XNOR U14196 ( .A(n13171), .B(n6588), .Z(n13174) );
  XNOR U14197 ( .A(n13167), .B(n13169), .Z(n6588) );
  NAND U14198 ( .A(n13175), .B(e_input[952]), .Z(n13169) );
  NAND U14199 ( .A(n12323), .B(e_input[952]), .Z(n13175) );
  XNOR U14200 ( .A(n13165), .B(n13176), .Z(n13167) );
  XOR U14201 ( .A(n13177), .B(n13178), .Z(n13165) );
  AND U14202 ( .A(n13179), .B(n13180), .Z(n13178) );
  XNOR U14203 ( .A(n13181), .B(n13177), .Z(n13180) );
  XOR U14204 ( .A(n13182), .B(e_input[952]), .Z(n13173) );
  IV U14205 ( .A(n13171), .Z(n13182) );
  XOR U14206 ( .A(n13183), .B(n13184), .Z(n13171) );
  AND U14207 ( .A(n13185), .B(n13186), .Z(n13184) );
  XNOR U14208 ( .A(n13183), .B(n6594), .Z(n13186) );
  XNOR U14209 ( .A(n13179), .B(n13181), .Z(n6594) );
  NAND U14210 ( .A(n13187), .B(e_input[951]), .Z(n13181) );
  NAND U14211 ( .A(n12323), .B(e_input[951]), .Z(n13187) );
  XNOR U14212 ( .A(n13177), .B(n13188), .Z(n13179) );
  XOR U14213 ( .A(n13189), .B(n13190), .Z(n13177) );
  AND U14214 ( .A(n13191), .B(n13192), .Z(n13190) );
  XNOR U14215 ( .A(n13193), .B(n13189), .Z(n13192) );
  XOR U14216 ( .A(n13194), .B(e_input[951]), .Z(n13185) );
  IV U14217 ( .A(n13183), .Z(n13194) );
  XOR U14218 ( .A(n13195), .B(n13196), .Z(n13183) );
  AND U14219 ( .A(n13197), .B(n13198), .Z(n13196) );
  XNOR U14220 ( .A(n13195), .B(n6600), .Z(n13198) );
  XNOR U14221 ( .A(n13191), .B(n13193), .Z(n6600) );
  NAND U14222 ( .A(n13199), .B(e_input[950]), .Z(n13193) );
  NAND U14223 ( .A(n12323), .B(e_input[950]), .Z(n13199) );
  XNOR U14224 ( .A(n13189), .B(n13200), .Z(n13191) );
  XOR U14225 ( .A(n13201), .B(n13202), .Z(n13189) );
  AND U14226 ( .A(n13203), .B(n13204), .Z(n13202) );
  XNOR U14227 ( .A(n13205), .B(n13201), .Z(n13204) );
  XOR U14228 ( .A(n13206), .B(e_input[950]), .Z(n13197) );
  IV U14229 ( .A(n13195), .Z(n13206) );
  XOR U14230 ( .A(n13207), .B(n13208), .Z(n13195) );
  AND U14231 ( .A(n13209), .B(n13210), .Z(n13208) );
  XNOR U14232 ( .A(n13207), .B(n6606), .Z(n13210) );
  XNOR U14233 ( .A(n13203), .B(n13205), .Z(n6606) );
  NAND U14234 ( .A(n13211), .B(e_input[949]), .Z(n13205) );
  NAND U14235 ( .A(n12323), .B(e_input[949]), .Z(n13211) );
  XNOR U14236 ( .A(n13201), .B(n13212), .Z(n13203) );
  XOR U14237 ( .A(n13213), .B(n13214), .Z(n13201) );
  AND U14238 ( .A(n13215), .B(n13216), .Z(n13214) );
  XNOR U14239 ( .A(n13217), .B(n13213), .Z(n13216) );
  XOR U14240 ( .A(n13218), .B(e_input[949]), .Z(n13209) );
  IV U14241 ( .A(n13207), .Z(n13218) );
  XOR U14242 ( .A(n13219), .B(n13220), .Z(n13207) );
  AND U14243 ( .A(n13221), .B(n13222), .Z(n13220) );
  XNOR U14244 ( .A(n13219), .B(n6612), .Z(n13222) );
  XNOR U14245 ( .A(n13215), .B(n13217), .Z(n6612) );
  NAND U14246 ( .A(n13223), .B(e_input[948]), .Z(n13217) );
  NAND U14247 ( .A(n12323), .B(e_input[948]), .Z(n13223) );
  XNOR U14248 ( .A(n13213), .B(n13224), .Z(n13215) );
  XOR U14249 ( .A(n13225), .B(n13226), .Z(n13213) );
  AND U14250 ( .A(n13227), .B(n13228), .Z(n13226) );
  XNOR U14251 ( .A(n13229), .B(n13225), .Z(n13228) );
  XOR U14252 ( .A(n13230), .B(e_input[948]), .Z(n13221) );
  IV U14253 ( .A(n13219), .Z(n13230) );
  XOR U14254 ( .A(n13231), .B(n13232), .Z(n13219) );
  AND U14255 ( .A(n13233), .B(n13234), .Z(n13232) );
  XNOR U14256 ( .A(n13231), .B(n6618), .Z(n13234) );
  XNOR U14257 ( .A(n13227), .B(n13229), .Z(n6618) );
  NAND U14258 ( .A(n13235), .B(e_input[947]), .Z(n13229) );
  NAND U14259 ( .A(n12323), .B(e_input[947]), .Z(n13235) );
  XNOR U14260 ( .A(n13225), .B(n13236), .Z(n13227) );
  XOR U14261 ( .A(n13237), .B(n13238), .Z(n13225) );
  AND U14262 ( .A(n13239), .B(n13240), .Z(n13238) );
  XNOR U14263 ( .A(n13241), .B(n13237), .Z(n13240) );
  XOR U14264 ( .A(n13242), .B(e_input[947]), .Z(n13233) );
  IV U14265 ( .A(n13231), .Z(n13242) );
  XOR U14266 ( .A(n13243), .B(n13244), .Z(n13231) );
  AND U14267 ( .A(n13245), .B(n13246), .Z(n13244) );
  XNOR U14268 ( .A(n13243), .B(n6624), .Z(n13246) );
  XNOR U14269 ( .A(n13239), .B(n13241), .Z(n6624) );
  NAND U14270 ( .A(n13247), .B(e_input[946]), .Z(n13241) );
  NAND U14271 ( .A(n12323), .B(e_input[946]), .Z(n13247) );
  XNOR U14272 ( .A(n13237), .B(n13248), .Z(n13239) );
  XOR U14273 ( .A(n13249), .B(n13250), .Z(n13237) );
  AND U14274 ( .A(n13251), .B(n13252), .Z(n13250) );
  XNOR U14275 ( .A(n13253), .B(n13249), .Z(n13252) );
  XOR U14276 ( .A(n13254), .B(e_input[946]), .Z(n13245) );
  IV U14277 ( .A(n13243), .Z(n13254) );
  XOR U14278 ( .A(n13255), .B(n13256), .Z(n13243) );
  AND U14279 ( .A(n13257), .B(n13258), .Z(n13256) );
  XNOR U14280 ( .A(n13255), .B(n6630), .Z(n13258) );
  XNOR U14281 ( .A(n13251), .B(n13253), .Z(n6630) );
  NAND U14282 ( .A(n13259), .B(e_input[945]), .Z(n13253) );
  NAND U14283 ( .A(n12323), .B(e_input[945]), .Z(n13259) );
  XNOR U14284 ( .A(n13249), .B(n13260), .Z(n13251) );
  XOR U14285 ( .A(n13261), .B(n13262), .Z(n13249) );
  AND U14286 ( .A(n13263), .B(n13264), .Z(n13262) );
  XNOR U14287 ( .A(n13265), .B(n13261), .Z(n13264) );
  XOR U14288 ( .A(n13266), .B(e_input[945]), .Z(n13257) );
  IV U14289 ( .A(n13255), .Z(n13266) );
  XOR U14290 ( .A(n13267), .B(n13268), .Z(n13255) );
  AND U14291 ( .A(n13269), .B(n13270), .Z(n13268) );
  XNOR U14292 ( .A(n13267), .B(n6636), .Z(n13270) );
  XNOR U14293 ( .A(n13263), .B(n13265), .Z(n6636) );
  NAND U14294 ( .A(n13271), .B(e_input[944]), .Z(n13265) );
  NAND U14295 ( .A(n12323), .B(e_input[944]), .Z(n13271) );
  XNOR U14296 ( .A(n13261), .B(n13272), .Z(n13263) );
  XOR U14297 ( .A(n13273), .B(n13274), .Z(n13261) );
  AND U14298 ( .A(n13275), .B(n13276), .Z(n13274) );
  XNOR U14299 ( .A(n13277), .B(n13273), .Z(n13276) );
  XOR U14300 ( .A(n13278), .B(e_input[944]), .Z(n13269) );
  IV U14301 ( .A(n13267), .Z(n13278) );
  XOR U14302 ( .A(n13279), .B(n13280), .Z(n13267) );
  AND U14303 ( .A(n13281), .B(n13282), .Z(n13280) );
  XNOR U14304 ( .A(n13279), .B(n6642), .Z(n13282) );
  XNOR U14305 ( .A(n13275), .B(n13277), .Z(n6642) );
  NAND U14306 ( .A(n13283), .B(e_input[943]), .Z(n13277) );
  NAND U14307 ( .A(n12323), .B(e_input[943]), .Z(n13283) );
  XNOR U14308 ( .A(n13273), .B(n13284), .Z(n13275) );
  XOR U14309 ( .A(n13285), .B(n13286), .Z(n13273) );
  AND U14310 ( .A(n13287), .B(n13288), .Z(n13286) );
  XNOR U14311 ( .A(n13289), .B(n13285), .Z(n13288) );
  XOR U14312 ( .A(n13290), .B(e_input[943]), .Z(n13281) );
  IV U14313 ( .A(n13279), .Z(n13290) );
  XOR U14314 ( .A(n13291), .B(n13292), .Z(n13279) );
  AND U14315 ( .A(n13293), .B(n13294), .Z(n13292) );
  XNOR U14316 ( .A(n13291), .B(n6648), .Z(n13294) );
  XNOR U14317 ( .A(n13287), .B(n13289), .Z(n6648) );
  NAND U14318 ( .A(n13295), .B(e_input[942]), .Z(n13289) );
  NAND U14319 ( .A(n12323), .B(e_input[942]), .Z(n13295) );
  XNOR U14320 ( .A(n13285), .B(n13296), .Z(n13287) );
  XOR U14321 ( .A(n13297), .B(n13298), .Z(n13285) );
  AND U14322 ( .A(n13299), .B(n13300), .Z(n13298) );
  XNOR U14323 ( .A(n13301), .B(n13297), .Z(n13300) );
  XOR U14324 ( .A(n13302), .B(e_input[942]), .Z(n13293) );
  IV U14325 ( .A(n13291), .Z(n13302) );
  XOR U14326 ( .A(n13303), .B(n13304), .Z(n13291) );
  AND U14327 ( .A(n13305), .B(n13306), .Z(n13304) );
  XNOR U14328 ( .A(n13303), .B(n6654), .Z(n13306) );
  XNOR U14329 ( .A(n13299), .B(n13301), .Z(n6654) );
  NAND U14330 ( .A(n13307), .B(e_input[941]), .Z(n13301) );
  NAND U14331 ( .A(n12323), .B(e_input[941]), .Z(n13307) );
  XNOR U14332 ( .A(n13297), .B(n13308), .Z(n13299) );
  XOR U14333 ( .A(n13309), .B(n13310), .Z(n13297) );
  AND U14334 ( .A(n13311), .B(n13312), .Z(n13310) );
  XNOR U14335 ( .A(n13313), .B(n13309), .Z(n13312) );
  XOR U14336 ( .A(n13314), .B(e_input[941]), .Z(n13305) );
  IV U14337 ( .A(n13303), .Z(n13314) );
  XOR U14338 ( .A(n13315), .B(n13316), .Z(n13303) );
  AND U14339 ( .A(n13317), .B(n13318), .Z(n13316) );
  XNOR U14340 ( .A(n13315), .B(n6660), .Z(n13318) );
  XNOR U14341 ( .A(n13311), .B(n13313), .Z(n6660) );
  NAND U14342 ( .A(n13319), .B(e_input[940]), .Z(n13313) );
  NAND U14343 ( .A(n12323), .B(e_input[940]), .Z(n13319) );
  XNOR U14344 ( .A(n13309), .B(n13320), .Z(n13311) );
  XOR U14345 ( .A(n13321), .B(n13322), .Z(n13309) );
  AND U14346 ( .A(n13323), .B(n13324), .Z(n13322) );
  XNOR U14347 ( .A(n13325), .B(n13321), .Z(n13324) );
  XOR U14348 ( .A(n13326), .B(e_input[940]), .Z(n13317) );
  IV U14349 ( .A(n13315), .Z(n13326) );
  XOR U14350 ( .A(n13327), .B(n13328), .Z(n13315) );
  AND U14351 ( .A(n13329), .B(n13330), .Z(n13328) );
  XNOR U14352 ( .A(n13327), .B(n6666), .Z(n13330) );
  XNOR U14353 ( .A(n13323), .B(n13325), .Z(n6666) );
  NAND U14354 ( .A(n13331), .B(e_input[939]), .Z(n13325) );
  NAND U14355 ( .A(n12323), .B(e_input[939]), .Z(n13331) );
  XNOR U14356 ( .A(n13321), .B(n13332), .Z(n13323) );
  XOR U14357 ( .A(n13333), .B(n13334), .Z(n13321) );
  AND U14358 ( .A(n13335), .B(n13336), .Z(n13334) );
  XNOR U14359 ( .A(n13337), .B(n13333), .Z(n13336) );
  XOR U14360 ( .A(n13338), .B(e_input[939]), .Z(n13329) );
  IV U14361 ( .A(n13327), .Z(n13338) );
  XOR U14362 ( .A(n13339), .B(n13340), .Z(n13327) );
  AND U14363 ( .A(n13341), .B(n13342), .Z(n13340) );
  XNOR U14364 ( .A(n13339), .B(n6672), .Z(n13342) );
  XNOR U14365 ( .A(n13335), .B(n13337), .Z(n6672) );
  NAND U14366 ( .A(n13343), .B(e_input[938]), .Z(n13337) );
  NAND U14367 ( .A(n12323), .B(e_input[938]), .Z(n13343) );
  XNOR U14368 ( .A(n13333), .B(n13344), .Z(n13335) );
  XOR U14369 ( .A(n13345), .B(n13346), .Z(n13333) );
  AND U14370 ( .A(n13347), .B(n13348), .Z(n13346) );
  XNOR U14371 ( .A(n13349), .B(n13345), .Z(n13348) );
  XOR U14372 ( .A(n13350), .B(e_input[938]), .Z(n13341) );
  IV U14373 ( .A(n13339), .Z(n13350) );
  XOR U14374 ( .A(n13351), .B(n13352), .Z(n13339) );
  AND U14375 ( .A(n13353), .B(n13354), .Z(n13352) );
  XNOR U14376 ( .A(n13351), .B(n6678), .Z(n13354) );
  XNOR U14377 ( .A(n13347), .B(n13349), .Z(n6678) );
  NAND U14378 ( .A(n13355), .B(e_input[937]), .Z(n13349) );
  NAND U14379 ( .A(n12323), .B(e_input[937]), .Z(n13355) );
  XNOR U14380 ( .A(n13345), .B(n13356), .Z(n13347) );
  XOR U14381 ( .A(n13357), .B(n13358), .Z(n13345) );
  AND U14382 ( .A(n13359), .B(n13360), .Z(n13358) );
  XNOR U14383 ( .A(n13361), .B(n13357), .Z(n13360) );
  XOR U14384 ( .A(n13362), .B(e_input[937]), .Z(n13353) );
  IV U14385 ( .A(n13351), .Z(n13362) );
  XOR U14386 ( .A(n13363), .B(n13364), .Z(n13351) );
  AND U14387 ( .A(n13365), .B(n13366), .Z(n13364) );
  XNOR U14388 ( .A(n13363), .B(n6684), .Z(n13366) );
  XNOR U14389 ( .A(n13359), .B(n13361), .Z(n6684) );
  NAND U14390 ( .A(n13367), .B(e_input[936]), .Z(n13361) );
  NAND U14391 ( .A(n12323), .B(e_input[936]), .Z(n13367) );
  XNOR U14392 ( .A(n13357), .B(n13368), .Z(n13359) );
  XOR U14393 ( .A(n13369), .B(n13370), .Z(n13357) );
  AND U14394 ( .A(n13371), .B(n13372), .Z(n13370) );
  XNOR U14395 ( .A(n13373), .B(n13369), .Z(n13372) );
  XOR U14396 ( .A(n13374), .B(e_input[936]), .Z(n13365) );
  IV U14397 ( .A(n13363), .Z(n13374) );
  XOR U14398 ( .A(n13375), .B(n13376), .Z(n13363) );
  AND U14399 ( .A(n13377), .B(n13378), .Z(n13376) );
  XNOR U14400 ( .A(n13375), .B(n6690), .Z(n13378) );
  XNOR U14401 ( .A(n13371), .B(n13373), .Z(n6690) );
  NAND U14402 ( .A(n13379), .B(e_input[935]), .Z(n13373) );
  NAND U14403 ( .A(n12323), .B(e_input[935]), .Z(n13379) );
  XNOR U14404 ( .A(n13369), .B(n13380), .Z(n13371) );
  XOR U14405 ( .A(n13381), .B(n13382), .Z(n13369) );
  AND U14406 ( .A(n13383), .B(n13384), .Z(n13382) );
  XNOR U14407 ( .A(n13385), .B(n13381), .Z(n13384) );
  XOR U14408 ( .A(n13386), .B(e_input[935]), .Z(n13377) );
  IV U14409 ( .A(n13375), .Z(n13386) );
  XOR U14410 ( .A(n13387), .B(n13388), .Z(n13375) );
  AND U14411 ( .A(n13389), .B(n13390), .Z(n13388) );
  XNOR U14412 ( .A(n13387), .B(n6696), .Z(n13390) );
  XNOR U14413 ( .A(n13383), .B(n13385), .Z(n6696) );
  NAND U14414 ( .A(n13391), .B(e_input[934]), .Z(n13385) );
  NAND U14415 ( .A(n12323), .B(e_input[934]), .Z(n13391) );
  XNOR U14416 ( .A(n13381), .B(n13392), .Z(n13383) );
  XOR U14417 ( .A(n13393), .B(n13394), .Z(n13381) );
  AND U14418 ( .A(n13395), .B(n13396), .Z(n13394) );
  XNOR U14419 ( .A(n13397), .B(n13393), .Z(n13396) );
  XOR U14420 ( .A(n13398), .B(e_input[934]), .Z(n13389) );
  IV U14421 ( .A(n13387), .Z(n13398) );
  XOR U14422 ( .A(n13399), .B(n13400), .Z(n13387) );
  AND U14423 ( .A(n13401), .B(n13402), .Z(n13400) );
  XNOR U14424 ( .A(n13399), .B(n6702), .Z(n13402) );
  XNOR U14425 ( .A(n13395), .B(n13397), .Z(n6702) );
  NAND U14426 ( .A(n13403), .B(e_input[933]), .Z(n13397) );
  NAND U14427 ( .A(n12323), .B(e_input[933]), .Z(n13403) );
  XNOR U14428 ( .A(n13393), .B(n13404), .Z(n13395) );
  XOR U14429 ( .A(n13405), .B(n13406), .Z(n13393) );
  AND U14430 ( .A(n13407), .B(n13408), .Z(n13406) );
  XNOR U14431 ( .A(n13409), .B(n13405), .Z(n13408) );
  XOR U14432 ( .A(n13410), .B(e_input[933]), .Z(n13401) );
  IV U14433 ( .A(n13399), .Z(n13410) );
  XOR U14434 ( .A(n13411), .B(n13412), .Z(n13399) );
  AND U14435 ( .A(n13413), .B(n13414), .Z(n13412) );
  XNOR U14436 ( .A(n13411), .B(n6708), .Z(n13414) );
  XNOR U14437 ( .A(n13407), .B(n13409), .Z(n6708) );
  NAND U14438 ( .A(n13415), .B(e_input[932]), .Z(n13409) );
  NAND U14439 ( .A(n12323), .B(e_input[932]), .Z(n13415) );
  XNOR U14440 ( .A(n13405), .B(n13416), .Z(n13407) );
  XOR U14441 ( .A(n13417), .B(n13418), .Z(n13405) );
  AND U14442 ( .A(n13419), .B(n13420), .Z(n13418) );
  XNOR U14443 ( .A(n13421), .B(n13417), .Z(n13420) );
  XOR U14444 ( .A(n13422), .B(e_input[932]), .Z(n13413) );
  IV U14445 ( .A(n13411), .Z(n13422) );
  XOR U14446 ( .A(n13423), .B(n13424), .Z(n13411) );
  AND U14447 ( .A(n13425), .B(n13426), .Z(n13424) );
  XNOR U14448 ( .A(n13423), .B(n6714), .Z(n13426) );
  XNOR U14449 ( .A(n13419), .B(n13421), .Z(n6714) );
  NAND U14450 ( .A(n13427), .B(e_input[931]), .Z(n13421) );
  NAND U14451 ( .A(n12323), .B(e_input[931]), .Z(n13427) );
  XNOR U14452 ( .A(n13417), .B(n13428), .Z(n13419) );
  XOR U14453 ( .A(n13429), .B(n13430), .Z(n13417) );
  AND U14454 ( .A(n13431), .B(n13432), .Z(n13430) );
  XNOR U14455 ( .A(n13433), .B(n13429), .Z(n13432) );
  XOR U14456 ( .A(n13434), .B(e_input[931]), .Z(n13425) );
  IV U14457 ( .A(n13423), .Z(n13434) );
  XOR U14458 ( .A(n13435), .B(n13436), .Z(n13423) );
  AND U14459 ( .A(n13437), .B(n13438), .Z(n13436) );
  XNOR U14460 ( .A(n13435), .B(n6720), .Z(n13438) );
  XNOR U14461 ( .A(n13431), .B(n13433), .Z(n6720) );
  NAND U14462 ( .A(n13439), .B(e_input[930]), .Z(n13433) );
  NAND U14463 ( .A(n12323), .B(e_input[930]), .Z(n13439) );
  XNOR U14464 ( .A(n13429), .B(n13440), .Z(n13431) );
  XOR U14465 ( .A(n13441), .B(n13442), .Z(n13429) );
  AND U14466 ( .A(n13443), .B(n13444), .Z(n13442) );
  XNOR U14467 ( .A(n13445), .B(n13441), .Z(n13444) );
  XOR U14468 ( .A(n13446), .B(e_input[930]), .Z(n13437) );
  IV U14469 ( .A(n13435), .Z(n13446) );
  XOR U14470 ( .A(n13447), .B(n13448), .Z(n13435) );
  AND U14471 ( .A(n13449), .B(n13450), .Z(n13448) );
  XNOR U14472 ( .A(n13447), .B(n6726), .Z(n13450) );
  XNOR U14473 ( .A(n13443), .B(n13445), .Z(n6726) );
  NAND U14474 ( .A(n13451), .B(e_input[929]), .Z(n13445) );
  NAND U14475 ( .A(n12323), .B(e_input[929]), .Z(n13451) );
  XNOR U14476 ( .A(n13441), .B(n13452), .Z(n13443) );
  XOR U14477 ( .A(n13453), .B(n13454), .Z(n13441) );
  AND U14478 ( .A(n13455), .B(n13456), .Z(n13454) );
  XNOR U14479 ( .A(n13457), .B(n13453), .Z(n13456) );
  XOR U14480 ( .A(n13458), .B(e_input[929]), .Z(n13449) );
  IV U14481 ( .A(n13447), .Z(n13458) );
  XOR U14482 ( .A(n13459), .B(n13460), .Z(n13447) );
  AND U14483 ( .A(n13461), .B(n13462), .Z(n13460) );
  XNOR U14484 ( .A(n13459), .B(n6732), .Z(n13462) );
  XNOR U14485 ( .A(n13455), .B(n13457), .Z(n6732) );
  NAND U14486 ( .A(n13463), .B(e_input[928]), .Z(n13457) );
  NAND U14487 ( .A(n12323), .B(e_input[928]), .Z(n13463) );
  XNOR U14488 ( .A(n13453), .B(n13464), .Z(n13455) );
  XOR U14489 ( .A(n13465), .B(n13466), .Z(n13453) );
  AND U14490 ( .A(n13467), .B(n13468), .Z(n13466) );
  XNOR U14491 ( .A(n13469), .B(n13465), .Z(n13468) );
  XOR U14492 ( .A(n13470), .B(e_input[928]), .Z(n13461) );
  IV U14493 ( .A(n13459), .Z(n13470) );
  XOR U14494 ( .A(n13471), .B(n13472), .Z(n13459) );
  AND U14495 ( .A(n13473), .B(n13474), .Z(n13472) );
  XNOR U14496 ( .A(n13471), .B(n6738), .Z(n13474) );
  XNOR U14497 ( .A(n13467), .B(n13469), .Z(n6738) );
  NAND U14498 ( .A(n13475), .B(e_input[927]), .Z(n13469) );
  NAND U14499 ( .A(n12323), .B(e_input[927]), .Z(n13475) );
  XNOR U14500 ( .A(n13465), .B(n13476), .Z(n13467) );
  XOR U14501 ( .A(n13477), .B(n13478), .Z(n13465) );
  AND U14502 ( .A(n13479), .B(n13480), .Z(n13478) );
  XNOR U14503 ( .A(n13481), .B(n13477), .Z(n13480) );
  XOR U14504 ( .A(n13482), .B(e_input[927]), .Z(n13473) );
  IV U14505 ( .A(n13471), .Z(n13482) );
  XOR U14506 ( .A(n13483), .B(n13484), .Z(n13471) );
  AND U14507 ( .A(n13485), .B(n13486), .Z(n13484) );
  XNOR U14508 ( .A(n13483), .B(n6744), .Z(n13486) );
  XNOR U14509 ( .A(n13479), .B(n13481), .Z(n6744) );
  NAND U14510 ( .A(n13487), .B(e_input[926]), .Z(n13481) );
  NAND U14511 ( .A(n12323), .B(e_input[926]), .Z(n13487) );
  XNOR U14512 ( .A(n13477), .B(n13488), .Z(n13479) );
  XOR U14513 ( .A(n13489), .B(n13490), .Z(n13477) );
  AND U14514 ( .A(n13491), .B(n13492), .Z(n13490) );
  XNOR U14515 ( .A(n13493), .B(n13489), .Z(n13492) );
  XOR U14516 ( .A(n13494), .B(e_input[926]), .Z(n13485) );
  IV U14517 ( .A(n13483), .Z(n13494) );
  XOR U14518 ( .A(n13495), .B(n13496), .Z(n13483) );
  AND U14519 ( .A(n13497), .B(n13498), .Z(n13496) );
  XNOR U14520 ( .A(n13495), .B(n6750), .Z(n13498) );
  XNOR U14521 ( .A(n13491), .B(n13493), .Z(n6750) );
  NAND U14522 ( .A(n13499), .B(e_input[925]), .Z(n13493) );
  NAND U14523 ( .A(n12323), .B(e_input[925]), .Z(n13499) );
  XNOR U14524 ( .A(n13489), .B(n13500), .Z(n13491) );
  XOR U14525 ( .A(n13501), .B(n13502), .Z(n13489) );
  AND U14526 ( .A(n13503), .B(n13504), .Z(n13502) );
  XNOR U14527 ( .A(n13505), .B(n13501), .Z(n13504) );
  XOR U14528 ( .A(n13506), .B(e_input[925]), .Z(n13497) );
  IV U14529 ( .A(n13495), .Z(n13506) );
  XOR U14530 ( .A(n13507), .B(n13508), .Z(n13495) );
  AND U14531 ( .A(n13509), .B(n13510), .Z(n13508) );
  XNOR U14532 ( .A(n13507), .B(n6756), .Z(n13510) );
  XNOR U14533 ( .A(n13503), .B(n13505), .Z(n6756) );
  NAND U14534 ( .A(n13511), .B(e_input[924]), .Z(n13505) );
  NAND U14535 ( .A(n12323), .B(e_input[924]), .Z(n13511) );
  XNOR U14536 ( .A(n13501), .B(n13512), .Z(n13503) );
  XOR U14537 ( .A(n13513), .B(n13514), .Z(n13501) );
  AND U14538 ( .A(n13515), .B(n13516), .Z(n13514) );
  XNOR U14539 ( .A(n13517), .B(n13513), .Z(n13516) );
  XOR U14540 ( .A(n13518), .B(e_input[924]), .Z(n13509) );
  IV U14541 ( .A(n13507), .Z(n13518) );
  XOR U14542 ( .A(n13519), .B(n13520), .Z(n13507) );
  AND U14543 ( .A(n13521), .B(n13522), .Z(n13520) );
  XNOR U14544 ( .A(n13519), .B(n6762), .Z(n13522) );
  XNOR U14545 ( .A(n13515), .B(n13517), .Z(n6762) );
  NAND U14546 ( .A(n13523), .B(e_input[923]), .Z(n13517) );
  NAND U14547 ( .A(n12323), .B(e_input[923]), .Z(n13523) );
  XNOR U14548 ( .A(n13513), .B(n13524), .Z(n13515) );
  XOR U14549 ( .A(n13525), .B(n13526), .Z(n13513) );
  AND U14550 ( .A(n13527), .B(n13528), .Z(n13526) );
  XNOR U14551 ( .A(n13529), .B(n13525), .Z(n13528) );
  XOR U14552 ( .A(n13530), .B(e_input[923]), .Z(n13521) );
  IV U14553 ( .A(n13519), .Z(n13530) );
  XOR U14554 ( .A(n13531), .B(n13532), .Z(n13519) );
  AND U14555 ( .A(n13533), .B(n13534), .Z(n13532) );
  XNOR U14556 ( .A(n13531), .B(n6768), .Z(n13534) );
  XNOR U14557 ( .A(n13527), .B(n13529), .Z(n6768) );
  NAND U14558 ( .A(n13535), .B(e_input[922]), .Z(n13529) );
  NAND U14559 ( .A(n12323), .B(e_input[922]), .Z(n13535) );
  XNOR U14560 ( .A(n13525), .B(n13536), .Z(n13527) );
  XOR U14561 ( .A(n13537), .B(n13538), .Z(n13525) );
  AND U14562 ( .A(n13539), .B(n13540), .Z(n13538) );
  XNOR U14563 ( .A(n13541), .B(n13537), .Z(n13540) );
  XOR U14564 ( .A(n13542), .B(e_input[922]), .Z(n13533) );
  IV U14565 ( .A(n13531), .Z(n13542) );
  XOR U14566 ( .A(n13543), .B(n13544), .Z(n13531) );
  AND U14567 ( .A(n13545), .B(n13546), .Z(n13544) );
  XNOR U14568 ( .A(n13543), .B(n6774), .Z(n13546) );
  XNOR U14569 ( .A(n13539), .B(n13541), .Z(n6774) );
  NAND U14570 ( .A(n13547), .B(e_input[921]), .Z(n13541) );
  NAND U14571 ( .A(n12323), .B(e_input[921]), .Z(n13547) );
  XNOR U14572 ( .A(n13537), .B(n13548), .Z(n13539) );
  XOR U14573 ( .A(n13549), .B(n13550), .Z(n13537) );
  AND U14574 ( .A(n13551), .B(n13552), .Z(n13550) );
  XNOR U14575 ( .A(n13553), .B(n13549), .Z(n13552) );
  XOR U14576 ( .A(n13554), .B(e_input[921]), .Z(n13545) );
  IV U14577 ( .A(n13543), .Z(n13554) );
  XOR U14578 ( .A(n13555), .B(n13556), .Z(n13543) );
  AND U14579 ( .A(n13557), .B(n13558), .Z(n13556) );
  XNOR U14580 ( .A(n13555), .B(n6780), .Z(n13558) );
  XNOR U14581 ( .A(n13551), .B(n13553), .Z(n6780) );
  NAND U14582 ( .A(n13559), .B(e_input[920]), .Z(n13553) );
  NAND U14583 ( .A(n12323), .B(e_input[920]), .Z(n13559) );
  XNOR U14584 ( .A(n13549), .B(n13560), .Z(n13551) );
  XOR U14585 ( .A(n13561), .B(n13562), .Z(n13549) );
  AND U14586 ( .A(n13563), .B(n13564), .Z(n13562) );
  XNOR U14587 ( .A(n13565), .B(n13561), .Z(n13564) );
  XOR U14588 ( .A(n13566), .B(e_input[920]), .Z(n13557) );
  IV U14589 ( .A(n13555), .Z(n13566) );
  XOR U14590 ( .A(n13567), .B(n13568), .Z(n13555) );
  AND U14591 ( .A(n13569), .B(n13570), .Z(n13568) );
  XNOR U14592 ( .A(n13567), .B(n6786), .Z(n13570) );
  XNOR U14593 ( .A(n13563), .B(n13565), .Z(n6786) );
  NAND U14594 ( .A(n13571), .B(e_input[919]), .Z(n13565) );
  NAND U14595 ( .A(n12323), .B(e_input[919]), .Z(n13571) );
  XNOR U14596 ( .A(n13561), .B(n13572), .Z(n13563) );
  XOR U14597 ( .A(n13573), .B(n13574), .Z(n13561) );
  AND U14598 ( .A(n13575), .B(n13576), .Z(n13574) );
  XNOR U14599 ( .A(n13577), .B(n13573), .Z(n13576) );
  XOR U14600 ( .A(n13578), .B(e_input[919]), .Z(n13569) );
  IV U14601 ( .A(n13567), .Z(n13578) );
  XOR U14602 ( .A(n13579), .B(n13580), .Z(n13567) );
  AND U14603 ( .A(n13581), .B(n13582), .Z(n13580) );
  XNOR U14604 ( .A(n13579), .B(n6792), .Z(n13582) );
  XNOR U14605 ( .A(n13575), .B(n13577), .Z(n6792) );
  NAND U14606 ( .A(n13583), .B(e_input[918]), .Z(n13577) );
  NAND U14607 ( .A(n12323), .B(e_input[918]), .Z(n13583) );
  XNOR U14608 ( .A(n13573), .B(n13584), .Z(n13575) );
  XOR U14609 ( .A(n13585), .B(n13586), .Z(n13573) );
  AND U14610 ( .A(n13587), .B(n13588), .Z(n13586) );
  XNOR U14611 ( .A(n13589), .B(n13585), .Z(n13588) );
  XOR U14612 ( .A(n13590), .B(e_input[918]), .Z(n13581) );
  IV U14613 ( .A(n13579), .Z(n13590) );
  XOR U14614 ( .A(n13591), .B(n13592), .Z(n13579) );
  AND U14615 ( .A(n13593), .B(n13594), .Z(n13592) );
  XNOR U14616 ( .A(n13591), .B(n6798), .Z(n13594) );
  XNOR U14617 ( .A(n13587), .B(n13589), .Z(n6798) );
  NAND U14618 ( .A(n13595), .B(e_input[917]), .Z(n13589) );
  NAND U14619 ( .A(n12323), .B(e_input[917]), .Z(n13595) );
  XNOR U14620 ( .A(n13585), .B(n13596), .Z(n13587) );
  XOR U14621 ( .A(n13597), .B(n13598), .Z(n13585) );
  AND U14622 ( .A(n13599), .B(n13600), .Z(n13598) );
  XNOR U14623 ( .A(n13601), .B(n13597), .Z(n13600) );
  XOR U14624 ( .A(n13602), .B(e_input[917]), .Z(n13593) );
  IV U14625 ( .A(n13591), .Z(n13602) );
  XOR U14626 ( .A(n13603), .B(n13604), .Z(n13591) );
  AND U14627 ( .A(n13605), .B(n13606), .Z(n13604) );
  XNOR U14628 ( .A(n13603), .B(n6804), .Z(n13606) );
  XNOR U14629 ( .A(n13599), .B(n13601), .Z(n6804) );
  NAND U14630 ( .A(n13607), .B(e_input[916]), .Z(n13601) );
  NAND U14631 ( .A(n12323), .B(e_input[916]), .Z(n13607) );
  XNOR U14632 ( .A(n13597), .B(n13608), .Z(n13599) );
  XOR U14633 ( .A(n13609), .B(n13610), .Z(n13597) );
  AND U14634 ( .A(n13611), .B(n13612), .Z(n13610) );
  XNOR U14635 ( .A(n13613), .B(n13609), .Z(n13612) );
  XOR U14636 ( .A(n13614), .B(e_input[916]), .Z(n13605) );
  IV U14637 ( .A(n13603), .Z(n13614) );
  XOR U14638 ( .A(n13615), .B(n13616), .Z(n13603) );
  AND U14639 ( .A(n13617), .B(n13618), .Z(n13616) );
  XNOR U14640 ( .A(n13615), .B(n6810), .Z(n13618) );
  XNOR U14641 ( .A(n13611), .B(n13613), .Z(n6810) );
  NAND U14642 ( .A(n13619), .B(e_input[915]), .Z(n13613) );
  NAND U14643 ( .A(n12323), .B(e_input[915]), .Z(n13619) );
  XNOR U14644 ( .A(n13609), .B(n13620), .Z(n13611) );
  XOR U14645 ( .A(n13621), .B(n13622), .Z(n13609) );
  AND U14646 ( .A(n13623), .B(n13624), .Z(n13622) );
  XNOR U14647 ( .A(n13625), .B(n13621), .Z(n13624) );
  XOR U14648 ( .A(n13626), .B(e_input[915]), .Z(n13617) );
  IV U14649 ( .A(n13615), .Z(n13626) );
  XOR U14650 ( .A(n13627), .B(n13628), .Z(n13615) );
  AND U14651 ( .A(n13629), .B(n13630), .Z(n13628) );
  XNOR U14652 ( .A(n13627), .B(n6816), .Z(n13630) );
  XNOR U14653 ( .A(n13623), .B(n13625), .Z(n6816) );
  NAND U14654 ( .A(n13631), .B(e_input[914]), .Z(n13625) );
  NAND U14655 ( .A(n12323), .B(e_input[914]), .Z(n13631) );
  XNOR U14656 ( .A(n13621), .B(n13632), .Z(n13623) );
  XOR U14657 ( .A(n13633), .B(n13634), .Z(n13621) );
  AND U14658 ( .A(n13635), .B(n13636), .Z(n13634) );
  XNOR U14659 ( .A(n13637), .B(n13633), .Z(n13636) );
  XOR U14660 ( .A(n13638), .B(e_input[914]), .Z(n13629) );
  IV U14661 ( .A(n13627), .Z(n13638) );
  XOR U14662 ( .A(n13639), .B(n13640), .Z(n13627) );
  AND U14663 ( .A(n13641), .B(n13642), .Z(n13640) );
  XNOR U14664 ( .A(n13639), .B(n6822), .Z(n13642) );
  XNOR U14665 ( .A(n13635), .B(n13637), .Z(n6822) );
  NAND U14666 ( .A(n13643), .B(e_input[913]), .Z(n13637) );
  NAND U14667 ( .A(n12323), .B(e_input[913]), .Z(n13643) );
  XNOR U14668 ( .A(n13633), .B(n13644), .Z(n13635) );
  XOR U14669 ( .A(n13645), .B(n13646), .Z(n13633) );
  AND U14670 ( .A(n13647), .B(n13648), .Z(n13646) );
  XNOR U14671 ( .A(n13649), .B(n13645), .Z(n13648) );
  XOR U14672 ( .A(n13650), .B(e_input[913]), .Z(n13641) );
  IV U14673 ( .A(n13639), .Z(n13650) );
  XOR U14674 ( .A(n13651), .B(n13652), .Z(n13639) );
  AND U14675 ( .A(n13653), .B(n13654), .Z(n13652) );
  XNOR U14676 ( .A(n13651), .B(n6828), .Z(n13654) );
  XNOR U14677 ( .A(n13647), .B(n13649), .Z(n6828) );
  NAND U14678 ( .A(n13655), .B(e_input[912]), .Z(n13649) );
  NAND U14679 ( .A(n12323), .B(e_input[912]), .Z(n13655) );
  XNOR U14680 ( .A(n13645), .B(n13656), .Z(n13647) );
  XOR U14681 ( .A(n13657), .B(n13658), .Z(n13645) );
  AND U14682 ( .A(n13659), .B(n13660), .Z(n13658) );
  XNOR U14683 ( .A(n13661), .B(n13657), .Z(n13660) );
  XOR U14684 ( .A(n13662), .B(e_input[912]), .Z(n13653) );
  IV U14685 ( .A(n13651), .Z(n13662) );
  XOR U14686 ( .A(n13663), .B(n13664), .Z(n13651) );
  AND U14687 ( .A(n13665), .B(n13666), .Z(n13664) );
  XNOR U14688 ( .A(n13663), .B(n6834), .Z(n13666) );
  XNOR U14689 ( .A(n13659), .B(n13661), .Z(n6834) );
  NAND U14690 ( .A(n13667), .B(e_input[911]), .Z(n13661) );
  NAND U14691 ( .A(n12323), .B(e_input[911]), .Z(n13667) );
  XNOR U14692 ( .A(n13657), .B(n13668), .Z(n13659) );
  XOR U14693 ( .A(n13669), .B(n13670), .Z(n13657) );
  AND U14694 ( .A(n13671), .B(n13672), .Z(n13670) );
  XNOR U14695 ( .A(n13673), .B(n13669), .Z(n13672) );
  XOR U14696 ( .A(n13674), .B(e_input[911]), .Z(n13665) );
  IV U14697 ( .A(n13663), .Z(n13674) );
  XOR U14698 ( .A(n13675), .B(n13676), .Z(n13663) );
  AND U14699 ( .A(n13677), .B(n13678), .Z(n13676) );
  XNOR U14700 ( .A(n13675), .B(n6840), .Z(n13678) );
  XNOR U14701 ( .A(n13671), .B(n13673), .Z(n6840) );
  NAND U14702 ( .A(n13679), .B(e_input[910]), .Z(n13673) );
  NAND U14703 ( .A(n12323), .B(e_input[910]), .Z(n13679) );
  XNOR U14704 ( .A(n13669), .B(n13680), .Z(n13671) );
  XOR U14705 ( .A(n13681), .B(n13682), .Z(n13669) );
  AND U14706 ( .A(n13683), .B(n13684), .Z(n13682) );
  XNOR U14707 ( .A(n13685), .B(n13681), .Z(n13684) );
  XOR U14708 ( .A(n13686), .B(e_input[910]), .Z(n13677) );
  IV U14709 ( .A(n13675), .Z(n13686) );
  XOR U14710 ( .A(n13687), .B(n13688), .Z(n13675) );
  AND U14711 ( .A(n13689), .B(n13690), .Z(n13688) );
  XNOR U14712 ( .A(n13687), .B(n6846), .Z(n13690) );
  XNOR U14713 ( .A(n13683), .B(n13685), .Z(n6846) );
  NAND U14714 ( .A(n13691), .B(e_input[909]), .Z(n13685) );
  NAND U14715 ( .A(n12323), .B(e_input[909]), .Z(n13691) );
  XNOR U14716 ( .A(n13681), .B(n13692), .Z(n13683) );
  XOR U14717 ( .A(n13693), .B(n13694), .Z(n13681) );
  AND U14718 ( .A(n13695), .B(n13696), .Z(n13694) );
  XNOR U14719 ( .A(n13697), .B(n13693), .Z(n13696) );
  XOR U14720 ( .A(n13698), .B(e_input[909]), .Z(n13689) );
  IV U14721 ( .A(n13687), .Z(n13698) );
  XOR U14722 ( .A(n13699), .B(n13700), .Z(n13687) );
  AND U14723 ( .A(n13701), .B(n13702), .Z(n13700) );
  XNOR U14724 ( .A(n13699), .B(n6852), .Z(n13702) );
  XNOR U14725 ( .A(n13695), .B(n13697), .Z(n6852) );
  NAND U14726 ( .A(n13703), .B(e_input[908]), .Z(n13697) );
  NAND U14727 ( .A(n12323), .B(e_input[908]), .Z(n13703) );
  XNOR U14728 ( .A(n13693), .B(n13704), .Z(n13695) );
  XOR U14729 ( .A(n13705), .B(n13706), .Z(n13693) );
  AND U14730 ( .A(n13707), .B(n13708), .Z(n13706) );
  XNOR U14731 ( .A(n13709), .B(n13705), .Z(n13708) );
  XOR U14732 ( .A(n13710), .B(e_input[908]), .Z(n13701) );
  IV U14733 ( .A(n13699), .Z(n13710) );
  XOR U14734 ( .A(n13711), .B(n13712), .Z(n13699) );
  AND U14735 ( .A(n13713), .B(n13714), .Z(n13712) );
  XNOR U14736 ( .A(n13711), .B(n6858), .Z(n13714) );
  XNOR U14737 ( .A(n13707), .B(n13709), .Z(n6858) );
  NAND U14738 ( .A(n13715), .B(e_input[907]), .Z(n13709) );
  NAND U14739 ( .A(n12323), .B(e_input[907]), .Z(n13715) );
  XNOR U14740 ( .A(n13705), .B(n13716), .Z(n13707) );
  XOR U14741 ( .A(n13717), .B(n13718), .Z(n13705) );
  AND U14742 ( .A(n13719), .B(n13720), .Z(n13718) );
  XNOR U14743 ( .A(n13721), .B(n13717), .Z(n13720) );
  XOR U14744 ( .A(n13722), .B(e_input[907]), .Z(n13713) );
  IV U14745 ( .A(n13711), .Z(n13722) );
  XOR U14746 ( .A(n13723), .B(n13724), .Z(n13711) );
  AND U14747 ( .A(n13725), .B(n13726), .Z(n13724) );
  XNOR U14748 ( .A(n13723), .B(n6864), .Z(n13726) );
  XNOR U14749 ( .A(n13719), .B(n13721), .Z(n6864) );
  NAND U14750 ( .A(n13727), .B(e_input[906]), .Z(n13721) );
  NAND U14751 ( .A(n12323), .B(e_input[906]), .Z(n13727) );
  XNOR U14752 ( .A(n13717), .B(n13728), .Z(n13719) );
  XOR U14753 ( .A(n13729), .B(n13730), .Z(n13717) );
  AND U14754 ( .A(n13731), .B(n13732), .Z(n13730) );
  XNOR U14755 ( .A(n13733), .B(n13729), .Z(n13732) );
  XOR U14756 ( .A(n13734), .B(e_input[906]), .Z(n13725) );
  IV U14757 ( .A(n13723), .Z(n13734) );
  XOR U14758 ( .A(n13735), .B(n13736), .Z(n13723) );
  AND U14759 ( .A(n13737), .B(n13738), .Z(n13736) );
  XNOR U14760 ( .A(n13735), .B(n6870), .Z(n13738) );
  XNOR U14761 ( .A(n13731), .B(n13733), .Z(n6870) );
  NAND U14762 ( .A(n13739), .B(e_input[905]), .Z(n13733) );
  NAND U14763 ( .A(n12323), .B(e_input[905]), .Z(n13739) );
  XNOR U14764 ( .A(n13729), .B(n13740), .Z(n13731) );
  XOR U14765 ( .A(n13741), .B(n13742), .Z(n13729) );
  AND U14766 ( .A(n13743), .B(n13744), .Z(n13742) );
  XNOR U14767 ( .A(n13745), .B(n13741), .Z(n13744) );
  XOR U14768 ( .A(n13746), .B(e_input[905]), .Z(n13737) );
  IV U14769 ( .A(n13735), .Z(n13746) );
  XOR U14770 ( .A(n13747), .B(n13748), .Z(n13735) );
  AND U14771 ( .A(n13749), .B(n13750), .Z(n13748) );
  XNOR U14772 ( .A(n13747), .B(n6876), .Z(n13750) );
  XNOR U14773 ( .A(n13743), .B(n13745), .Z(n6876) );
  NAND U14774 ( .A(n13751), .B(e_input[904]), .Z(n13745) );
  NAND U14775 ( .A(n12323), .B(e_input[904]), .Z(n13751) );
  XNOR U14776 ( .A(n13741), .B(n13752), .Z(n13743) );
  XOR U14777 ( .A(n13753), .B(n13754), .Z(n13741) );
  AND U14778 ( .A(n13755), .B(n13756), .Z(n13754) );
  XNOR U14779 ( .A(n13757), .B(n13753), .Z(n13756) );
  XOR U14780 ( .A(n13758), .B(e_input[904]), .Z(n13749) );
  IV U14781 ( .A(n13747), .Z(n13758) );
  XOR U14782 ( .A(n13759), .B(n13760), .Z(n13747) );
  AND U14783 ( .A(n13761), .B(n13762), .Z(n13760) );
  XNOR U14784 ( .A(n13759), .B(n6882), .Z(n13762) );
  XNOR U14785 ( .A(n13755), .B(n13757), .Z(n6882) );
  NAND U14786 ( .A(n13763), .B(e_input[903]), .Z(n13757) );
  NAND U14787 ( .A(n12323), .B(e_input[903]), .Z(n13763) );
  XNOR U14788 ( .A(n13753), .B(n13764), .Z(n13755) );
  XOR U14789 ( .A(n13765), .B(n13766), .Z(n13753) );
  AND U14790 ( .A(n13767), .B(n13768), .Z(n13766) );
  XNOR U14791 ( .A(n13769), .B(n13765), .Z(n13768) );
  XOR U14792 ( .A(n13770), .B(e_input[903]), .Z(n13761) );
  IV U14793 ( .A(n13759), .Z(n13770) );
  XOR U14794 ( .A(n13771), .B(n13772), .Z(n13759) );
  AND U14795 ( .A(n13773), .B(n13774), .Z(n13772) );
  XNOR U14796 ( .A(n13771), .B(n6888), .Z(n13774) );
  XNOR U14797 ( .A(n13767), .B(n13769), .Z(n6888) );
  NAND U14798 ( .A(n13775), .B(e_input[902]), .Z(n13769) );
  NAND U14799 ( .A(n12323), .B(e_input[902]), .Z(n13775) );
  XNOR U14800 ( .A(n13765), .B(n13776), .Z(n13767) );
  XOR U14801 ( .A(n13777), .B(n13778), .Z(n13765) );
  AND U14802 ( .A(n13779), .B(n13780), .Z(n13778) );
  XNOR U14803 ( .A(n13781), .B(n13777), .Z(n13780) );
  XOR U14804 ( .A(n13782), .B(e_input[902]), .Z(n13773) );
  IV U14805 ( .A(n13771), .Z(n13782) );
  XOR U14806 ( .A(n13783), .B(n13784), .Z(n13771) );
  AND U14807 ( .A(n13785), .B(n13786), .Z(n13784) );
  XNOR U14808 ( .A(n13783), .B(n6894), .Z(n13786) );
  XNOR U14809 ( .A(n13779), .B(n13781), .Z(n6894) );
  NAND U14810 ( .A(n13787), .B(e_input[901]), .Z(n13781) );
  NAND U14811 ( .A(n12323), .B(e_input[901]), .Z(n13787) );
  XNOR U14812 ( .A(n13777), .B(n13788), .Z(n13779) );
  XOR U14813 ( .A(n13789), .B(n13790), .Z(n13777) );
  AND U14814 ( .A(n13791), .B(n13792), .Z(n13790) );
  XNOR U14815 ( .A(n13793), .B(n13789), .Z(n13792) );
  XOR U14816 ( .A(n13794), .B(e_input[901]), .Z(n13785) );
  IV U14817 ( .A(n13783), .Z(n13794) );
  XOR U14818 ( .A(n13795), .B(n13796), .Z(n13783) );
  AND U14819 ( .A(n13797), .B(n13798), .Z(n13796) );
  XNOR U14820 ( .A(n13795), .B(n6900), .Z(n13798) );
  XNOR U14821 ( .A(n13791), .B(n13793), .Z(n6900) );
  NAND U14822 ( .A(n13799), .B(e_input[900]), .Z(n13793) );
  NAND U14823 ( .A(n12323), .B(e_input[900]), .Z(n13799) );
  XNOR U14824 ( .A(n13789), .B(n13800), .Z(n13791) );
  XOR U14825 ( .A(n13801), .B(n13802), .Z(n13789) );
  AND U14826 ( .A(n13803), .B(n13804), .Z(n13802) );
  XNOR U14827 ( .A(n13805), .B(n13801), .Z(n13804) );
  XOR U14828 ( .A(n13806), .B(e_input[900]), .Z(n13797) );
  IV U14829 ( .A(n13795), .Z(n13806) );
  XOR U14830 ( .A(n13807), .B(n13808), .Z(n13795) );
  AND U14831 ( .A(n13809), .B(n13810), .Z(n13808) );
  XNOR U14832 ( .A(n13807), .B(n6906), .Z(n13810) );
  XNOR U14833 ( .A(n13803), .B(n13805), .Z(n6906) );
  NAND U14834 ( .A(n13811), .B(e_input[899]), .Z(n13805) );
  NAND U14835 ( .A(n12323), .B(e_input[899]), .Z(n13811) );
  XNOR U14836 ( .A(n13801), .B(n13812), .Z(n13803) );
  XOR U14837 ( .A(n13813), .B(n13814), .Z(n13801) );
  AND U14838 ( .A(n13815), .B(n13816), .Z(n13814) );
  XNOR U14839 ( .A(n13817), .B(n13813), .Z(n13816) );
  XOR U14840 ( .A(n13818), .B(e_input[899]), .Z(n13809) );
  IV U14841 ( .A(n13807), .Z(n13818) );
  XOR U14842 ( .A(n13819), .B(n13820), .Z(n13807) );
  AND U14843 ( .A(n13821), .B(n13822), .Z(n13820) );
  XNOR U14844 ( .A(n13819), .B(n6912), .Z(n13822) );
  XNOR U14845 ( .A(n13815), .B(n13817), .Z(n6912) );
  NAND U14846 ( .A(n13823), .B(e_input[898]), .Z(n13817) );
  NAND U14847 ( .A(n12323), .B(e_input[898]), .Z(n13823) );
  XNOR U14848 ( .A(n13813), .B(n13824), .Z(n13815) );
  XOR U14849 ( .A(n13825), .B(n13826), .Z(n13813) );
  AND U14850 ( .A(n13827), .B(n13828), .Z(n13826) );
  XNOR U14851 ( .A(n13829), .B(n13825), .Z(n13828) );
  XOR U14852 ( .A(n13830), .B(e_input[898]), .Z(n13821) );
  IV U14853 ( .A(n13819), .Z(n13830) );
  XOR U14854 ( .A(n13831), .B(n13832), .Z(n13819) );
  AND U14855 ( .A(n13833), .B(n13834), .Z(n13832) );
  XNOR U14856 ( .A(n13831), .B(n6918), .Z(n13834) );
  XNOR U14857 ( .A(n13827), .B(n13829), .Z(n6918) );
  NAND U14858 ( .A(n13835), .B(e_input[897]), .Z(n13829) );
  NAND U14859 ( .A(n12323), .B(e_input[897]), .Z(n13835) );
  XNOR U14860 ( .A(n13825), .B(n13836), .Z(n13827) );
  XOR U14861 ( .A(n13837), .B(n13838), .Z(n13825) );
  AND U14862 ( .A(n13839), .B(n13840), .Z(n13838) );
  XNOR U14863 ( .A(n13841), .B(n13837), .Z(n13840) );
  XOR U14864 ( .A(n13842), .B(e_input[897]), .Z(n13833) );
  IV U14865 ( .A(n13831), .Z(n13842) );
  XOR U14866 ( .A(n13843), .B(n13844), .Z(n13831) );
  AND U14867 ( .A(n13845), .B(n13846), .Z(n13844) );
  XNOR U14868 ( .A(n13843), .B(n6924), .Z(n13846) );
  XNOR U14869 ( .A(n13839), .B(n13841), .Z(n6924) );
  NAND U14870 ( .A(n13847), .B(e_input[896]), .Z(n13841) );
  NAND U14871 ( .A(n12323), .B(e_input[896]), .Z(n13847) );
  XNOR U14872 ( .A(n13837), .B(n13848), .Z(n13839) );
  XOR U14873 ( .A(n13849), .B(n13850), .Z(n13837) );
  AND U14874 ( .A(n13851), .B(n13852), .Z(n13850) );
  XNOR U14875 ( .A(n13853), .B(n13849), .Z(n13852) );
  XOR U14876 ( .A(n13854), .B(e_input[896]), .Z(n13845) );
  IV U14877 ( .A(n13843), .Z(n13854) );
  XOR U14878 ( .A(n13855), .B(n13856), .Z(n13843) );
  AND U14879 ( .A(n13857), .B(n13858), .Z(n13856) );
  XNOR U14880 ( .A(n13855), .B(n6930), .Z(n13858) );
  XNOR U14881 ( .A(n13851), .B(n13853), .Z(n6930) );
  NAND U14882 ( .A(n13859), .B(e_input[895]), .Z(n13853) );
  NAND U14883 ( .A(n12323), .B(e_input[895]), .Z(n13859) );
  XNOR U14884 ( .A(n13849), .B(n13860), .Z(n13851) );
  XOR U14885 ( .A(n13861), .B(n13862), .Z(n13849) );
  AND U14886 ( .A(n13863), .B(n13864), .Z(n13862) );
  XNOR U14887 ( .A(n13865), .B(n13861), .Z(n13864) );
  XOR U14888 ( .A(n13866), .B(e_input[895]), .Z(n13857) );
  IV U14889 ( .A(n13855), .Z(n13866) );
  XOR U14890 ( .A(n13867), .B(n13868), .Z(n13855) );
  AND U14891 ( .A(n13869), .B(n13870), .Z(n13868) );
  XNOR U14892 ( .A(n13867), .B(n6936), .Z(n13870) );
  XNOR U14893 ( .A(n13863), .B(n13865), .Z(n6936) );
  NAND U14894 ( .A(n13871), .B(e_input[894]), .Z(n13865) );
  NAND U14895 ( .A(n12323), .B(e_input[894]), .Z(n13871) );
  XNOR U14896 ( .A(n13861), .B(n13872), .Z(n13863) );
  XOR U14897 ( .A(n13873), .B(n13874), .Z(n13861) );
  AND U14898 ( .A(n13875), .B(n13876), .Z(n13874) );
  XNOR U14899 ( .A(n13877), .B(n13873), .Z(n13876) );
  XOR U14900 ( .A(n13878), .B(e_input[894]), .Z(n13869) );
  IV U14901 ( .A(n13867), .Z(n13878) );
  XOR U14902 ( .A(n13879), .B(n13880), .Z(n13867) );
  AND U14903 ( .A(n13881), .B(n13882), .Z(n13880) );
  XNOR U14904 ( .A(n13879), .B(n6942), .Z(n13882) );
  XNOR U14905 ( .A(n13875), .B(n13877), .Z(n6942) );
  NAND U14906 ( .A(n13883), .B(e_input[893]), .Z(n13877) );
  NAND U14907 ( .A(n12323), .B(e_input[893]), .Z(n13883) );
  XNOR U14908 ( .A(n13873), .B(n13884), .Z(n13875) );
  XOR U14909 ( .A(n13885), .B(n13886), .Z(n13873) );
  AND U14910 ( .A(n13887), .B(n13888), .Z(n13886) );
  XNOR U14911 ( .A(n13889), .B(n13885), .Z(n13888) );
  XOR U14912 ( .A(n13890), .B(e_input[893]), .Z(n13881) );
  IV U14913 ( .A(n13879), .Z(n13890) );
  XOR U14914 ( .A(n13891), .B(n13892), .Z(n13879) );
  AND U14915 ( .A(n13893), .B(n13894), .Z(n13892) );
  XNOR U14916 ( .A(n13891), .B(n6948), .Z(n13894) );
  XNOR U14917 ( .A(n13887), .B(n13889), .Z(n6948) );
  NAND U14918 ( .A(n13895), .B(e_input[892]), .Z(n13889) );
  NAND U14919 ( .A(n12323), .B(e_input[892]), .Z(n13895) );
  XNOR U14920 ( .A(n13885), .B(n13896), .Z(n13887) );
  XOR U14921 ( .A(n13897), .B(n13898), .Z(n13885) );
  AND U14922 ( .A(n13899), .B(n13900), .Z(n13898) );
  XNOR U14923 ( .A(n13901), .B(n13897), .Z(n13900) );
  XOR U14924 ( .A(n13902), .B(e_input[892]), .Z(n13893) );
  IV U14925 ( .A(n13891), .Z(n13902) );
  XOR U14926 ( .A(n13903), .B(n13904), .Z(n13891) );
  AND U14927 ( .A(n13905), .B(n13906), .Z(n13904) );
  XNOR U14928 ( .A(n13903), .B(n6954), .Z(n13906) );
  XNOR U14929 ( .A(n13899), .B(n13901), .Z(n6954) );
  NAND U14930 ( .A(n13907), .B(e_input[891]), .Z(n13901) );
  NAND U14931 ( .A(n12323), .B(e_input[891]), .Z(n13907) );
  XNOR U14932 ( .A(n13897), .B(n13908), .Z(n13899) );
  XOR U14933 ( .A(n13909), .B(n13910), .Z(n13897) );
  AND U14934 ( .A(n13911), .B(n13912), .Z(n13910) );
  XNOR U14935 ( .A(n13913), .B(n13909), .Z(n13912) );
  XOR U14936 ( .A(n13914), .B(e_input[891]), .Z(n13905) );
  IV U14937 ( .A(n13903), .Z(n13914) );
  XOR U14938 ( .A(n13915), .B(n13916), .Z(n13903) );
  AND U14939 ( .A(n13917), .B(n13918), .Z(n13916) );
  XNOR U14940 ( .A(n13915), .B(n6960), .Z(n13918) );
  XNOR U14941 ( .A(n13911), .B(n13913), .Z(n6960) );
  NAND U14942 ( .A(n13919), .B(e_input[890]), .Z(n13913) );
  NAND U14943 ( .A(n12323), .B(e_input[890]), .Z(n13919) );
  XNOR U14944 ( .A(n13909), .B(n13920), .Z(n13911) );
  XOR U14945 ( .A(n13921), .B(n13922), .Z(n13909) );
  AND U14946 ( .A(n13923), .B(n13924), .Z(n13922) );
  XNOR U14947 ( .A(n13925), .B(n13921), .Z(n13924) );
  XOR U14948 ( .A(n13926), .B(e_input[890]), .Z(n13917) );
  IV U14949 ( .A(n13915), .Z(n13926) );
  XOR U14950 ( .A(n13927), .B(n13928), .Z(n13915) );
  AND U14951 ( .A(n13929), .B(n13930), .Z(n13928) );
  XNOR U14952 ( .A(n13927), .B(n6966), .Z(n13930) );
  XNOR U14953 ( .A(n13923), .B(n13925), .Z(n6966) );
  NAND U14954 ( .A(n13931), .B(e_input[889]), .Z(n13925) );
  NAND U14955 ( .A(n12323), .B(e_input[889]), .Z(n13931) );
  XNOR U14956 ( .A(n13921), .B(n13932), .Z(n13923) );
  XOR U14957 ( .A(n13933), .B(n13934), .Z(n13921) );
  AND U14958 ( .A(n13935), .B(n13936), .Z(n13934) );
  XNOR U14959 ( .A(n13937), .B(n13933), .Z(n13936) );
  XOR U14960 ( .A(n13938), .B(e_input[889]), .Z(n13929) );
  IV U14961 ( .A(n13927), .Z(n13938) );
  XOR U14962 ( .A(n13939), .B(n13940), .Z(n13927) );
  AND U14963 ( .A(n13941), .B(n13942), .Z(n13940) );
  XNOR U14964 ( .A(n13939), .B(n6972), .Z(n13942) );
  XNOR U14965 ( .A(n13935), .B(n13937), .Z(n6972) );
  NAND U14966 ( .A(n13943), .B(e_input[888]), .Z(n13937) );
  NAND U14967 ( .A(n12323), .B(e_input[888]), .Z(n13943) );
  XNOR U14968 ( .A(n13933), .B(n13944), .Z(n13935) );
  XOR U14969 ( .A(n13945), .B(n13946), .Z(n13933) );
  AND U14970 ( .A(n13947), .B(n13948), .Z(n13946) );
  XNOR U14971 ( .A(n13949), .B(n13945), .Z(n13948) );
  XOR U14972 ( .A(n13950), .B(e_input[888]), .Z(n13941) );
  IV U14973 ( .A(n13939), .Z(n13950) );
  XOR U14974 ( .A(n13951), .B(n13952), .Z(n13939) );
  AND U14975 ( .A(n13953), .B(n13954), .Z(n13952) );
  XNOR U14976 ( .A(n13951), .B(n6978), .Z(n13954) );
  XNOR U14977 ( .A(n13947), .B(n13949), .Z(n6978) );
  NAND U14978 ( .A(n13955), .B(e_input[887]), .Z(n13949) );
  NAND U14979 ( .A(n12323), .B(e_input[887]), .Z(n13955) );
  XNOR U14980 ( .A(n13945), .B(n13956), .Z(n13947) );
  XOR U14981 ( .A(n13957), .B(n13958), .Z(n13945) );
  AND U14982 ( .A(n13959), .B(n13960), .Z(n13958) );
  XNOR U14983 ( .A(n13961), .B(n13957), .Z(n13960) );
  XOR U14984 ( .A(n13962), .B(e_input[887]), .Z(n13953) );
  IV U14985 ( .A(n13951), .Z(n13962) );
  XOR U14986 ( .A(n13963), .B(n13964), .Z(n13951) );
  AND U14987 ( .A(n13965), .B(n13966), .Z(n13964) );
  XNOR U14988 ( .A(n13963), .B(n6984), .Z(n13966) );
  XNOR U14989 ( .A(n13959), .B(n13961), .Z(n6984) );
  NAND U14990 ( .A(n13967), .B(e_input[886]), .Z(n13961) );
  NAND U14991 ( .A(n12323), .B(e_input[886]), .Z(n13967) );
  XNOR U14992 ( .A(n13957), .B(n13968), .Z(n13959) );
  XOR U14993 ( .A(n13969), .B(n13970), .Z(n13957) );
  AND U14994 ( .A(n13971), .B(n13972), .Z(n13970) );
  XNOR U14995 ( .A(n13973), .B(n13969), .Z(n13972) );
  XOR U14996 ( .A(n13974), .B(e_input[886]), .Z(n13965) );
  IV U14997 ( .A(n13963), .Z(n13974) );
  XOR U14998 ( .A(n13975), .B(n13976), .Z(n13963) );
  AND U14999 ( .A(n13977), .B(n13978), .Z(n13976) );
  XNOR U15000 ( .A(n13975), .B(n6990), .Z(n13978) );
  XNOR U15001 ( .A(n13971), .B(n13973), .Z(n6990) );
  NAND U15002 ( .A(n13979), .B(e_input[885]), .Z(n13973) );
  NAND U15003 ( .A(n12323), .B(e_input[885]), .Z(n13979) );
  XNOR U15004 ( .A(n13969), .B(n13980), .Z(n13971) );
  XOR U15005 ( .A(n13981), .B(n13982), .Z(n13969) );
  AND U15006 ( .A(n13983), .B(n13984), .Z(n13982) );
  XNOR U15007 ( .A(n13985), .B(n13981), .Z(n13984) );
  XOR U15008 ( .A(n13986), .B(e_input[885]), .Z(n13977) );
  IV U15009 ( .A(n13975), .Z(n13986) );
  XOR U15010 ( .A(n13987), .B(n13988), .Z(n13975) );
  AND U15011 ( .A(n13989), .B(n13990), .Z(n13988) );
  XNOR U15012 ( .A(n13987), .B(n6996), .Z(n13990) );
  XNOR U15013 ( .A(n13983), .B(n13985), .Z(n6996) );
  NAND U15014 ( .A(n13991), .B(e_input[884]), .Z(n13985) );
  NAND U15015 ( .A(n12323), .B(e_input[884]), .Z(n13991) );
  XNOR U15016 ( .A(n13981), .B(n13992), .Z(n13983) );
  XOR U15017 ( .A(n13993), .B(n13994), .Z(n13981) );
  AND U15018 ( .A(n13995), .B(n13996), .Z(n13994) );
  XNOR U15019 ( .A(n13997), .B(n13993), .Z(n13996) );
  XOR U15020 ( .A(n13998), .B(e_input[884]), .Z(n13989) );
  IV U15021 ( .A(n13987), .Z(n13998) );
  XOR U15022 ( .A(n13999), .B(n14000), .Z(n13987) );
  AND U15023 ( .A(n14001), .B(n14002), .Z(n14000) );
  XNOR U15024 ( .A(n13999), .B(n7002), .Z(n14002) );
  XNOR U15025 ( .A(n13995), .B(n13997), .Z(n7002) );
  NAND U15026 ( .A(n14003), .B(e_input[883]), .Z(n13997) );
  NAND U15027 ( .A(n12323), .B(e_input[883]), .Z(n14003) );
  XNOR U15028 ( .A(n13993), .B(n14004), .Z(n13995) );
  XOR U15029 ( .A(n14005), .B(n14006), .Z(n13993) );
  AND U15030 ( .A(n14007), .B(n14008), .Z(n14006) );
  XNOR U15031 ( .A(n14009), .B(n14005), .Z(n14008) );
  XOR U15032 ( .A(n14010), .B(e_input[883]), .Z(n14001) );
  IV U15033 ( .A(n13999), .Z(n14010) );
  XOR U15034 ( .A(n14011), .B(n14012), .Z(n13999) );
  AND U15035 ( .A(n14013), .B(n14014), .Z(n14012) );
  XNOR U15036 ( .A(n14011), .B(n7008), .Z(n14014) );
  XNOR U15037 ( .A(n14007), .B(n14009), .Z(n7008) );
  NAND U15038 ( .A(n14015), .B(e_input[882]), .Z(n14009) );
  NAND U15039 ( .A(n12323), .B(e_input[882]), .Z(n14015) );
  XNOR U15040 ( .A(n14005), .B(n14016), .Z(n14007) );
  XOR U15041 ( .A(n14017), .B(n14018), .Z(n14005) );
  AND U15042 ( .A(n14019), .B(n14020), .Z(n14018) );
  XNOR U15043 ( .A(n14021), .B(n14017), .Z(n14020) );
  XOR U15044 ( .A(n14022), .B(e_input[882]), .Z(n14013) );
  IV U15045 ( .A(n14011), .Z(n14022) );
  XOR U15046 ( .A(n14023), .B(n14024), .Z(n14011) );
  AND U15047 ( .A(n14025), .B(n14026), .Z(n14024) );
  XNOR U15048 ( .A(n14023), .B(n7014), .Z(n14026) );
  XNOR U15049 ( .A(n14019), .B(n14021), .Z(n7014) );
  NAND U15050 ( .A(n14027), .B(e_input[881]), .Z(n14021) );
  NAND U15051 ( .A(n12323), .B(e_input[881]), .Z(n14027) );
  XNOR U15052 ( .A(n14017), .B(n14028), .Z(n14019) );
  XOR U15053 ( .A(n14029), .B(n14030), .Z(n14017) );
  AND U15054 ( .A(n14031), .B(n14032), .Z(n14030) );
  XNOR U15055 ( .A(n14033), .B(n14029), .Z(n14032) );
  XOR U15056 ( .A(n14034), .B(e_input[881]), .Z(n14025) );
  IV U15057 ( .A(n14023), .Z(n14034) );
  XOR U15058 ( .A(n14035), .B(n14036), .Z(n14023) );
  AND U15059 ( .A(n14037), .B(n14038), .Z(n14036) );
  XNOR U15060 ( .A(n14035), .B(n7020), .Z(n14038) );
  XNOR U15061 ( .A(n14031), .B(n14033), .Z(n7020) );
  NAND U15062 ( .A(n14039), .B(e_input[880]), .Z(n14033) );
  NAND U15063 ( .A(n12323), .B(e_input[880]), .Z(n14039) );
  XNOR U15064 ( .A(n14029), .B(n14040), .Z(n14031) );
  XOR U15065 ( .A(n14041), .B(n14042), .Z(n14029) );
  AND U15066 ( .A(n14043), .B(n14044), .Z(n14042) );
  XNOR U15067 ( .A(n14045), .B(n14041), .Z(n14044) );
  XOR U15068 ( .A(n14046), .B(e_input[880]), .Z(n14037) );
  IV U15069 ( .A(n14035), .Z(n14046) );
  XOR U15070 ( .A(n14047), .B(n14048), .Z(n14035) );
  AND U15071 ( .A(n14049), .B(n14050), .Z(n14048) );
  XNOR U15072 ( .A(n14047), .B(n7026), .Z(n14050) );
  XNOR U15073 ( .A(n14043), .B(n14045), .Z(n7026) );
  NAND U15074 ( .A(n14051), .B(e_input[879]), .Z(n14045) );
  NAND U15075 ( .A(n12323), .B(e_input[879]), .Z(n14051) );
  XNOR U15076 ( .A(n14041), .B(n14052), .Z(n14043) );
  XOR U15077 ( .A(n14053), .B(n14054), .Z(n14041) );
  AND U15078 ( .A(n14055), .B(n14056), .Z(n14054) );
  XNOR U15079 ( .A(n14057), .B(n14053), .Z(n14056) );
  XOR U15080 ( .A(n14058), .B(e_input[879]), .Z(n14049) );
  IV U15081 ( .A(n14047), .Z(n14058) );
  XOR U15082 ( .A(n14059), .B(n14060), .Z(n14047) );
  AND U15083 ( .A(n14061), .B(n14062), .Z(n14060) );
  XNOR U15084 ( .A(n14059), .B(n7032), .Z(n14062) );
  XNOR U15085 ( .A(n14055), .B(n14057), .Z(n7032) );
  NAND U15086 ( .A(n14063), .B(e_input[878]), .Z(n14057) );
  NAND U15087 ( .A(n12323), .B(e_input[878]), .Z(n14063) );
  XNOR U15088 ( .A(n14053), .B(n14064), .Z(n14055) );
  XOR U15089 ( .A(n14065), .B(n14066), .Z(n14053) );
  AND U15090 ( .A(n14067), .B(n14068), .Z(n14066) );
  XNOR U15091 ( .A(n14069), .B(n14065), .Z(n14068) );
  XOR U15092 ( .A(n14070), .B(e_input[878]), .Z(n14061) );
  IV U15093 ( .A(n14059), .Z(n14070) );
  XOR U15094 ( .A(n14071), .B(n14072), .Z(n14059) );
  AND U15095 ( .A(n14073), .B(n14074), .Z(n14072) );
  XNOR U15096 ( .A(n14071), .B(n7038), .Z(n14074) );
  XNOR U15097 ( .A(n14067), .B(n14069), .Z(n7038) );
  NAND U15098 ( .A(n14075), .B(e_input[877]), .Z(n14069) );
  NAND U15099 ( .A(n12323), .B(e_input[877]), .Z(n14075) );
  XNOR U15100 ( .A(n14065), .B(n14076), .Z(n14067) );
  XOR U15101 ( .A(n14077), .B(n14078), .Z(n14065) );
  AND U15102 ( .A(n14079), .B(n14080), .Z(n14078) );
  XNOR U15103 ( .A(n14081), .B(n14077), .Z(n14080) );
  XOR U15104 ( .A(n14082), .B(e_input[877]), .Z(n14073) );
  IV U15105 ( .A(n14071), .Z(n14082) );
  XOR U15106 ( .A(n14083), .B(n14084), .Z(n14071) );
  AND U15107 ( .A(n14085), .B(n14086), .Z(n14084) );
  XNOR U15108 ( .A(n14083), .B(n7044), .Z(n14086) );
  XNOR U15109 ( .A(n14079), .B(n14081), .Z(n7044) );
  NAND U15110 ( .A(n14087), .B(e_input[876]), .Z(n14081) );
  NAND U15111 ( .A(n12323), .B(e_input[876]), .Z(n14087) );
  XNOR U15112 ( .A(n14077), .B(n14088), .Z(n14079) );
  XOR U15113 ( .A(n14089), .B(n14090), .Z(n14077) );
  AND U15114 ( .A(n14091), .B(n14092), .Z(n14090) );
  XNOR U15115 ( .A(n14093), .B(n14089), .Z(n14092) );
  XOR U15116 ( .A(n14094), .B(e_input[876]), .Z(n14085) );
  IV U15117 ( .A(n14083), .Z(n14094) );
  XOR U15118 ( .A(n14095), .B(n14096), .Z(n14083) );
  AND U15119 ( .A(n14097), .B(n14098), .Z(n14096) );
  XNOR U15120 ( .A(n14095), .B(n7050), .Z(n14098) );
  XNOR U15121 ( .A(n14091), .B(n14093), .Z(n7050) );
  NAND U15122 ( .A(n14099), .B(e_input[875]), .Z(n14093) );
  NAND U15123 ( .A(n12323), .B(e_input[875]), .Z(n14099) );
  XNOR U15124 ( .A(n14089), .B(n14100), .Z(n14091) );
  XOR U15125 ( .A(n14101), .B(n14102), .Z(n14089) );
  AND U15126 ( .A(n14103), .B(n14104), .Z(n14102) );
  XNOR U15127 ( .A(n14105), .B(n14101), .Z(n14104) );
  XOR U15128 ( .A(n14106), .B(e_input[875]), .Z(n14097) );
  IV U15129 ( .A(n14095), .Z(n14106) );
  XOR U15130 ( .A(n14107), .B(n14108), .Z(n14095) );
  AND U15131 ( .A(n14109), .B(n14110), .Z(n14108) );
  XNOR U15132 ( .A(n14107), .B(n7056), .Z(n14110) );
  XNOR U15133 ( .A(n14103), .B(n14105), .Z(n7056) );
  NAND U15134 ( .A(n14111), .B(e_input[874]), .Z(n14105) );
  NAND U15135 ( .A(n12323), .B(e_input[874]), .Z(n14111) );
  XNOR U15136 ( .A(n14101), .B(n14112), .Z(n14103) );
  XOR U15137 ( .A(n14113), .B(n14114), .Z(n14101) );
  AND U15138 ( .A(n14115), .B(n14116), .Z(n14114) );
  XNOR U15139 ( .A(n14117), .B(n14113), .Z(n14116) );
  XOR U15140 ( .A(n14118), .B(e_input[874]), .Z(n14109) );
  IV U15141 ( .A(n14107), .Z(n14118) );
  XOR U15142 ( .A(n14119), .B(n14120), .Z(n14107) );
  AND U15143 ( .A(n14121), .B(n14122), .Z(n14120) );
  XNOR U15144 ( .A(n14119), .B(n7062), .Z(n14122) );
  XNOR U15145 ( .A(n14115), .B(n14117), .Z(n7062) );
  NAND U15146 ( .A(n14123), .B(e_input[873]), .Z(n14117) );
  NAND U15147 ( .A(n12323), .B(e_input[873]), .Z(n14123) );
  XNOR U15148 ( .A(n14113), .B(n14124), .Z(n14115) );
  XOR U15149 ( .A(n14125), .B(n14126), .Z(n14113) );
  AND U15150 ( .A(n14127), .B(n14128), .Z(n14126) );
  XNOR U15151 ( .A(n14129), .B(n14125), .Z(n14128) );
  XOR U15152 ( .A(n14130), .B(e_input[873]), .Z(n14121) );
  IV U15153 ( .A(n14119), .Z(n14130) );
  XOR U15154 ( .A(n14131), .B(n14132), .Z(n14119) );
  AND U15155 ( .A(n14133), .B(n14134), .Z(n14132) );
  XNOR U15156 ( .A(n14131), .B(n7068), .Z(n14134) );
  XNOR U15157 ( .A(n14127), .B(n14129), .Z(n7068) );
  NAND U15158 ( .A(n14135), .B(e_input[872]), .Z(n14129) );
  NAND U15159 ( .A(n12323), .B(e_input[872]), .Z(n14135) );
  XNOR U15160 ( .A(n14125), .B(n14136), .Z(n14127) );
  XOR U15161 ( .A(n14137), .B(n14138), .Z(n14125) );
  AND U15162 ( .A(n14139), .B(n14140), .Z(n14138) );
  XNOR U15163 ( .A(n14141), .B(n14137), .Z(n14140) );
  XOR U15164 ( .A(n14142), .B(e_input[872]), .Z(n14133) );
  IV U15165 ( .A(n14131), .Z(n14142) );
  XOR U15166 ( .A(n14143), .B(n14144), .Z(n14131) );
  AND U15167 ( .A(n14145), .B(n14146), .Z(n14144) );
  XNOR U15168 ( .A(n14143), .B(n7074), .Z(n14146) );
  XNOR U15169 ( .A(n14139), .B(n14141), .Z(n7074) );
  NAND U15170 ( .A(n14147), .B(e_input[871]), .Z(n14141) );
  NAND U15171 ( .A(n12323), .B(e_input[871]), .Z(n14147) );
  XNOR U15172 ( .A(n14137), .B(n14148), .Z(n14139) );
  XOR U15173 ( .A(n14149), .B(n14150), .Z(n14137) );
  AND U15174 ( .A(n14151), .B(n14152), .Z(n14150) );
  XNOR U15175 ( .A(n14153), .B(n14149), .Z(n14152) );
  XOR U15176 ( .A(n14154), .B(e_input[871]), .Z(n14145) );
  IV U15177 ( .A(n14143), .Z(n14154) );
  XOR U15178 ( .A(n14155), .B(n14156), .Z(n14143) );
  AND U15179 ( .A(n14157), .B(n14158), .Z(n14156) );
  XNOR U15180 ( .A(n14155), .B(n7080), .Z(n14158) );
  XNOR U15181 ( .A(n14151), .B(n14153), .Z(n7080) );
  NAND U15182 ( .A(n14159), .B(e_input[870]), .Z(n14153) );
  NAND U15183 ( .A(n12323), .B(e_input[870]), .Z(n14159) );
  XNOR U15184 ( .A(n14149), .B(n14160), .Z(n14151) );
  XOR U15185 ( .A(n14161), .B(n14162), .Z(n14149) );
  AND U15186 ( .A(n14163), .B(n14164), .Z(n14162) );
  XNOR U15187 ( .A(n14165), .B(n14161), .Z(n14164) );
  XOR U15188 ( .A(n14166), .B(e_input[870]), .Z(n14157) );
  IV U15189 ( .A(n14155), .Z(n14166) );
  XOR U15190 ( .A(n14167), .B(n14168), .Z(n14155) );
  AND U15191 ( .A(n14169), .B(n14170), .Z(n14168) );
  XNOR U15192 ( .A(n14167), .B(n7086), .Z(n14170) );
  XNOR U15193 ( .A(n14163), .B(n14165), .Z(n7086) );
  NAND U15194 ( .A(n14171), .B(e_input[869]), .Z(n14165) );
  NAND U15195 ( .A(n12323), .B(e_input[869]), .Z(n14171) );
  XNOR U15196 ( .A(n14161), .B(n14172), .Z(n14163) );
  XOR U15197 ( .A(n14173), .B(n14174), .Z(n14161) );
  AND U15198 ( .A(n14175), .B(n14176), .Z(n14174) );
  XNOR U15199 ( .A(n14177), .B(n14173), .Z(n14176) );
  XOR U15200 ( .A(n14178), .B(e_input[869]), .Z(n14169) );
  IV U15201 ( .A(n14167), .Z(n14178) );
  XOR U15202 ( .A(n14179), .B(n14180), .Z(n14167) );
  AND U15203 ( .A(n14181), .B(n14182), .Z(n14180) );
  XNOR U15204 ( .A(n14179), .B(n7092), .Z(n14182) );
  XNOR U15205 ( .A(n14175), .B(n14177), .Z(n7092) );
  NAND U15206 ( .A(n14183), .B(e_input[868]), .Z(n14177) );
  NAND U15207 ( .A(n12323), .B(e_input[868]), .Z(n14183) );
  XNOR U15208 ( .A(n14173), .B(n14184), .Z(n14175) );
  XOR U15209 ( .A(n14185), .B(n14186), .Z(n14173) );
  AND U15210 ( .A(n14187), .B(n14188), .Z(n14186) );
  XNOR U15211 ( .A(n14189), .B(n14185), .Z(n14188) );
  XOR U15212 ( .A(n14190), .B(e_input[868]), .Z(n14181) );
  IV U15213 ( .A(n14179), .Z(n14190) );
  XOR U15214 ( .A(n14191), .B(n14192), .Z(n14179) );
  AND U15215 ( .A(n14193), .B(n14194), .Z(n14192) );
  XNOR U15216 ( .A(n14191), .B(n7098), .Z(n14194) );
  XNOR U15217 ( .A(n14187), .B(n14189), .Z(n7098) );
  NAND U15218 ( .A(n14195), .B(e_input[867]), .Z(n14189) );
  NAND U15219 ( .A(n12323), .B(e_input[867]), .Z(n14195) );
  XNOR U15220 ( .A(n14185), .B(n14196), .Z(n14187) );
  XOR U15221 ( .A(n14197), .B(n14198), .Z(n14185) );
  AND U15222 ( .A(n14199), .B(n14200), .Z(n14198) );
  XNOR U15223 ( .A(n14201), .B(n14197), .Z(n14200) );
  XOR U15224 ( .A(n14202), .B(e_input[867]), .Z(n14193) );
  IV U15225 ( .A(n14191), .Z(n14202) );
  XOR U15226 ( .A(n14203), .B(n14204), .Z(n14191) );
  AND U15227 ( .A(n14205), .B(n14206), .Z(n14204) );
  XNOR U15228 ( .A(n14203), .B(n7104), .Z(n14206) );
  XNOR U15229 ( .A(n14199), .B(n14201), .Z(n7104) );
  NAND U15230 ( .A(n14207), .B(e_input[866]), .Z(n14201) );
  NAND U15231 ( .A(n12323), .B(e_input[866]), .Z(n14207) );
  XNOR U15232 ( .A(n14197), .B(n14208), .Z(n14199) );
  XOR U15233 ( .A(n14209), .B(n14210), .Z(n14197) );
  AND U15234 ( .A(n14211), .B(n14212), .Z(n14210) );
  XNOR U15235 ( .A(n14213), .B(n14209), .Z(n14212) );
  XOR U15236 ( .A(n14214), .B(e_input[866]), .Z(n14205) );
  IV U15237 ( .A(n14203), .Z(n14214) );
  XOR U15238 ( .A(n14215), .B(n14216), .Z(n14203) );
  AND U15239 ( .A(n14217), .B(n14218), .Z(n14216) );
  XNOR U15240 ( .A(n14215), .B(n7110), .Z(n14218) );
  XNOR U15241 ( .A(n14211), .B(n14213), .Z(n7110) );
  NAND U15242 ( .A(n14219), .B(e_input[865]), .Z(n14213) );
  NAND U15243 ( .A(n12323), .B(e_input[865]), .Z(n14219) );
  XNOR U15244 ( .A(n14209), .B(n14220), .Z(n14211) );
  XOR U15245 ( .A(n14221), .B(n14222), .Z(n14209) );
  AND U15246 ( .A(n14223), .B(n14224), .Z(n14222) );
  XNOR U15247 ( .A(n14225), .B(n14221), .Z(n14224) );
  XOR U15248 ( .A(n14226), .B(e_input[865]), .Z(n14217) );
  IV U15249 ( .A(n14215), .Z(n14226) );
  XOR U15250 ( .A(n14227), .B(n14228), .Z(n14215) );
  AND U15251 ( .A(n14229), .B(n14230), .Z(n14228) );
  XNOR U15252 ( .A(n14227), .B(n7116), .Z(n14230) );
  XNOR U15253 ( .A(n14223), .B(n14225), .Z(n7116) );
  NAND U15254 ( .A(n14231), .B(e_input[864]), .Z(n14225) );
  NAND U15255 ( .A(n12323), .B(e_input[864]), .Z(n14231) );
  XNOR U15256 ( .A(n14221), .B(n14232), .Z(n14223) );
  XOR U15257 ( .A(n14233), .B(n14234), .Z(n14221) );
  AND U15258 ( .A(n14235), .B(n14236), .Z(n14234) );
  XNOR U15259 ( .A(n14237), .B(n14233), .Z(n14236) );
  XOR U15260 ( .A(n14238), .B(e_input[864]), .Z(n14229) );
  IV U15261 ( .A(n14227), .Z(n14238) );
  XOR U15262 ( .A(n14239), .B(n14240), .Z(n14227) );
  AND U15263 ( .A(n14241), .B(n14242), .Z(n14240) );
  XNOR U15264 ( .A(n14239), .B(n7122), .Z(n14242) );
  XNOR U15265 ( .A(n14235), .B(n14237), .Z(n7122) );
  NAND U15266 ( .A(n14243), .B(e_input[863]), .Z(n14237) );
  NAND U15267 ( .A(n12323), .B(e_input[863]), .Z(n14243) );
  XNOR U15268 ( .A(n14233), .B(n14244), .Z(n14235) );
  XOR U15269 ( .A(n14245), .B(n14246), .Z(n14233) );
  AND U15270 ( .A(n14247), .B(n14248), .Z(n14246) );
  XNOR U15271 ( .A(n14249), .B(n14245), .Z(n14248) );
  XOR U15272 ( .A(n14250), .B(e_input[863]), .Z(n14241) );
  IV U15273 ( .A(n14239), .Z(n14250) );
  XOR U15274 ( .A(n14251), .B(n14252), .Z(n14239) );
  AND U15275 ( .A(n14253), .B(n14254), .Z(n14252) );
  XNOR U15276 ( .A(n14251), .B(n7128), .Z(n14254) );
  XNOR U15277 ( .A(n14247), .B(n14249), .Z(n7128) );
  NAND U15278 ( .A(n14255), .B(e_input[862]), .Z(n14249) );
  NAND U15279 ( .A(n12323), .B(e_input[862]), .Z(n14255) );
  XNOR U15280 ( .A(n14245), .B(n14256), .Z(n14247) );
  XOR U15281 ( .A(n14257), .B(n14258), .Z(n14245) );
  AND U15282 ( .A(n14259), .B(n14260), .Z(n14258) );
  XNOR U15283 ( .A(n14261), .B(n14257), .Z(n14260) );
  XOR U15284 ( .A(n14262), .B(e_input[862]), .Z(n14253) );
  IV U15285 ( .A(n14251), .Z(n14262) );
  XOR U15286 ( .A(n14263), .B(n14264), .Z(n14251) );
  AND U15287 ( .A(n14265), .B(n14266), .Z(n14264) );
  XNOR U15288 ( .A(n14263), .B(n7134), .Z(n14266) );
  XNOR U15289 ( .A(n14259), .B(n14261), .Z(n7134) );
  NAND U15290 ( .A(n14267), .B(e_input[861]), .Z(n14261) );
  NAND U15291 ( .A(n12323), .B(e_input[861]), .Z(n14267) );
  XNOR U15292 ( .A(n14257), .B(n14268), .Z(n14259) );
  XOR U15293 ( .A(n14269), .B(n14270), .Z(n14257) );
  AND U15294 ( .A(n14271), .B(n14272), .Z(n14270) );
  XNOR U15295 ( .A(n14273), .B(n14269), .Z(n14272) );
  XOR U15296 ( .A(n14274), .B(e_input[861]), .Z(n14265) );
  IV U15297 ( .A(n14263), .Z(n14274) );
  XOR U15298 ( .A(n14275), .B(n14276), .Z(n14263) );
  AND U15299 ( .A(n14277), .B(n14278), .Z(n14276) );
  XNOR U15300 ( .A(n14275), .B(n7140), .Z(n14278) );
  XNOR U15301 ( .A(n14271), .B(n14273), .Z(n7140) );
  NAND U15302 ( .A(n14279), .B(e_input[860]), .Z(n14273) );
  NAND U15303 ( .A(n12323), .B(e_input[860]), .Z(n14279) );
  XNOR U15304 ( .A(n14269), .B(n14280), .Z(n14271) );
  XOR U15305 ( .A(n14281), .B(n14282), .Z(n14269) );
  AND U15306 ( .A(n14283), .B(n14284), .Z(n14282) );
  XNOR U15307 ( .A(n14285), .B(n14281), .Z(n14284) );
  XOR U15308 ( .A(n14286), .B(e_input[860]), .Z(n14277) );
  IV U15309 ( .A(n14275), .Z(n14286) );
  XOR U15310 ( .A(n14287), .B(n14288), .Z(n14275) );
  AND U15311 ( .A(n14289), .B(n14290), .Z(n14288) );
  XNOR U15312 ( .A(n14287), .B(n7146), .Z(n14290) );
  XNOR U15313 ( .A(n14283), .B(n14285), .Z(n7146) );
  NAND U15314 ( .A(n14291), .B(e_input[859]), .Z(n14285) );
  NAND U15315 ( .A(n12323), .B(e_input[859]), .Z(n14291) );
  XNOR U15316 ( .A(n14281), .B(n14292), .Z(n14283) );
  XOR U15317 ( .A(n14293), .B(n14294), .Z(n14281) );
  AND U15318 ( .A(n14295), .B(n14296), .Z(n14294) );
  XNOR U15319 ( .A(n14297), .B(n14293), .Z(n14296) );
  XOR U15320 ( .A(n14298), .B(e_input[859]), .Z(n14289) );
  IV U15321 ( .A(n14287), .Z(n14298) );
  XOR U15322 ( .A(n14299), .B(n14300), .Z(n14287) );
  AND U15323 ( .A(n14301), .B(n14302), .Z(n14300) );
  XNOR U15324 ( .A(n14299), .B(n7152), .Z(n14302) );
  XNOR U15325 ( .A(n14295), .B(n14297), .Z(n7152) );
  NAND U15326 ( .A(n14303), .B(e_input[858]), .Z(n14297) );
  NAND U15327 ( .A(n12323), .B(e_input[858]), .Z(n14303) );
  XNOR U15328 ( .A(n14293), .B(n14304), .Z(n14295) );
  XOR U15329 ( .A(n14305), .B(n14306), .Z(n14293) );
  AND U15330 ( .A(n14307), .B(n14308), .Z(n14306) );
  XNOR U15331 ( .A(n14309), .B(n14305), .Z(n14308) );
  XOR U15332 ( .A(n14310), .B(e_input[858]), .Z(n14301) );
  IV U15333 ( .A(n14299), .Z(n14310) );
  XOR U15334 ( .A(n14311), .B(n14312), .Z(n14299) );
  AND U15335 ( .A(n14313), .B(n14314), .Z(n14312) );
  XNOR U15336 ( .A(n14311), .B(n7158), .Z(n14314) );
  XNOR U15337 ( .A(n14307), .B(n14309), .Z(n7158) );
  NAND U15338 ( .A(n14315), .B(e_input[857]), .Z(n14309) );
  NAND U15339 ( .A(n12323), .B(e_input[857]), .Z(n14315) );
  XNOR U15340 ( .A(n14305), .B(n14316), .Z(n14307) );
  XOR U15341 ( .A(n14317), .B(n14318), .Z(n14305) );
  AND U15342 ( .A(n14319), .B(n14320), .Z(n14318) );
  XNOR U15343 ( .A(n14321), .B(n14317), .Z(n14320) );
  XOR U15344 ( .A(n14322), .B(e_input[857]), .Z(n14313) );
  IV U15345 ( .A(n14311), .Z(n14322) );
  XOR U15346 ( .A(n14323), .B(n14324), .Z(n14311) );
  AND U15347 ( .A(n14325), .B(n14326), .Z(n14324) );
  XNOR U15348 ( .A(n14323), .B(n7164), .Z(n14326) );
  XNOR U15349 ( .A(n14319), .B(n14321), .Z(n7164) );
  NAND U15350 ( .A(n14327), .B(e_input[856]), .Z(n14321) );
  NAND U15351 ( .A(n12323), .B(e_input[856]), .Z(n14327) );
  XNOR U15352 ( .A(n14317), .B(n14328), .Z(n14319) );
  XOR U15353 ( .A(n14329), .B(n14330), .Z(n14317) );
  AND U15354 ( .A(n14331), .B(n14332), .Z(n14330) );
  XNOR U15355 ( .A(n14333), .B(n14329), .Z(n14332) );
  XOR U15356 ( .A(n14334), .B(e_input[856]), .Z(n14325) );
  IV U15357 ( .A(n14323), .Z(n14334) );
  XOR U15358 ( .A(n14335), .B(n14336), .Z(n14323) );
  AND U15359 ( .A(n14337), .B(n14338), .Z(n14336) );
  XNOR U15360 ( .A(n14335), .B(n7170), .Z(n14338) );
  XNOR U15361 ( .A(n14331), .B(n14333), .Z(n7170) );
  NAND U15362 ( .A(n14339), .B(e_input[855]), .Z(n14333) );
  NAND U15363 ( .A(n12323), .B(e_input[855]), .Z(n14339) );
  XNOR U15364 ( .A(n14329), .B(n14340), .Z(n14331) );
  XOR U15365 ( .A(n14341), .B(n14342), .Z(n14329) );
  AND U15366 ( .A(n14343), .B(n14344), .Z(n14342) );
  XNOR U15367 ( .A(n14345), .B(n14341), .Z(n14344) );
  XOR U15368 ( .A(n14346), .B(e_input[855]), .Z(n14337) );
  IV U15369 ( .A(n14335), .Z(n14346) );
  XOR U15370 ( .A(n14347), .B(n14348), .Z(n14335) );
  AND U15371 ( .A(n14349), .B(n14350), .Z(n14348) );
  XNOR U15372 ( .A(n14347), .B(n7176), .Z(n14350) );
  XNOR U15373 ( .A(n14343), .B(n14345), .Z(n7176) );
  NAND U15374 ( .A(n14351), .B(e_input[854]), .Z(n14345) );
  NAND U15375 ( .A(n12323), .B(e_input[854]), .Z(n14351) );
  XNOR U15376 ( .A(n14341), .B(n14352), .Z(n14343) );
  XOR U15377 ( .A(n14353), .B(n14354), .Z(n14341) );
  AND U15378 ( .A(n14355), .B(n14356), .Z(n14354) );
  XNOR U15379 ( .A(n14357), .B(n14353), .Z(n14356) );
  XOR U15380 ( .A(n14358), .B(e_input[854]), .Z(n14349) );
  IV U15381 ( .A(n14347), .Z(n14358) );
  XOR U15382 ( .A(n14359), .B(n14360), .Z(n14347) );
  AND U15383 ( .A(n14361), .B(n14362), .Z(n14360) );
  XNOR U15384 ( .A(n14359), .B(n7182), .Z(n14362) );
  XNOR U15385 ( .A(n14355), .B(n14357), .Z(n7182) );
  NAND U15386 ( .A(n14363), .B(e_input[853]), .Z(n14357) );
  NAND U15387 ( .A(n12323), .B(e_input[853]), .Z(n14363) );
  XNOR U15388 ( .A(n14353), .B(n14364), .Z(n14355) );
  XOR U15389 ( .A(n14365), .B(n14366), .Z(n14353) );
  AND U15390 ( .A(n14367), .B(n14368), .Z(n14366) );
  XNOR U15391 ( .A(n14369), .B(n14365), .Z(n14368) );
  XOR U15392 ( .A(n14370), .B(e_input[853]), .Z(n14361) );
  IV U15393 ( .A(n14359), .Z(n14370) );
  XOR U15394 ( .A(n14371), .B(n14372), .Z(n14359) );
  AND U15395 ( .A(n14373), .B(n14374), .Z(n14372) );
  XNOR U15396 ( .A(n14371), .B(n7188), .Z(n14374) );
  XNOR U15397 ( .A(n14367), .B(n14369), .Z(n7188) );
  NAND U15398 ( .A(n14375), .B(e_input[852]), .Z(n14369) );
  NAND U15399 ( .A(n12323), .B(e_input[852]), .Z(n14375) );
  XNOR U15400 ( .A(n14365), .B(n14376), .Z(n14367) );
  XOR U15401 ( .A(n14377), .B(n14378), .Z(n14365) );
  AND U15402 ( .A(n14379), .B(n14380), .Z(n14378) );
  XNOR U15403 ( .A(n14381), .B(n14377), .Z(n14380) );
  XOR U15404 ( .A(n14382), .B(e_input[852]), .Z(n14373) );
  IV U15405 ( .A(n14371), .Z(n14382) );
  XOR U15406 ( .A(n14383), .B(n14384), .Z(n14371) );
  AND U15407 ( .A(n14385), .B(n14386), .Z(n14384) );
  XNOR U15408 ( .A(n14383), .B(n7194), .Z(n14386) );
  XNOR U15409 ( .A(n14379), .B(n14381), .Z(n7194) );
  NAND U15410 ( .A(n14387), .B(e_input[851]), .Z(n14381) );
  NAND U15411 ( .A(n12323), .B(e_input[851]), .Z(n14387) );
  XNOR U15412 ( .A(n14377), .B(n14388), .Z(n14379) );
  XOR U15413 ( .A(n14389), .B(n14390), .Z(n14377) );
  AND U15414 ( .A(n14391), .B(n14392), .Z(n14390) );
  XNOR U15415 ( .A(n14393), .B(n14389), .Z(n14392) );
  XOR U15416 ( .A(n14394), .B(e_input[851]), .Z(n14385) );
  IV U15417 ( .A(n14383), .Z(n14394) );
  XOR U15418 ( .A(n14395), .B(n14396), .Z(n14383) );
  AND U15419 ( .A(n14397), .B(n14398), .Z(n14396) );
  XNOR U15420 ( .A(n14395), .B(n7200), .Z(n14398) );
  XNOR U15421 ( .A(n14391), .B(n14393), .Z(n7200) );
  NAND U15422 ( .A(n14399), .B(e_input[850]), .Z(n14393) );
  NAND U15423 ( .A(n12323), .B(e_input[850]), .Z(n14399) );
  XNOR U15424 ( .A(n14389), .B(n14400), .Z(n14391) );
  XOR U15425 ( .A(n14401), .B(n14402), .Z(n14389) );
  AND U15426 ( .A(n14403), .B(n14404), .Z(n14402) );
  XNOR U15427 ( .A(n14405), .B(n14401), .Z(n14404) );
  XOR U15428 ( .A(n14406), .B(e_input[850]), .Z(n14397) );
  IV U15429 ( .A(n14395), .Z(n14406) );
  XOR U15430 ( .A(n14407), .B(n14408), .Z(n14395) );
  AND U15431 ( .A(n14409), .B(n14410), .Z(n14408) );
  XNOR U15432 ( .A(n14407), .B(n7206), .Z(n14410) );
  XNOR U15433 ( .A(n14403), .B(n14405), .Z(n7206) );
  NAND U15434 ( .A(n14411), .B(e_input[849]), .Z(n14405) );
  NAND U15435 ( .A(n12323), .B(e_input[849]), .Z(n14411) );
  XNOR U15436 ( .A(n14401), .B(n14412), .Z(n14403) );
  XOR U15437 ( .A(n14413), .B(n14414), .Z(n14401) );
  AND U15438 ( .A(n14415), .B(n14416), .Z(n14414) );
  XNOR U15439 ( .A(n14417), .B(n14413), .Z(n14416) );
  XOR U15440 ( .A(n14418), .B(e_input[849]), .Z(n14409) );
  IV U15441 ( .A(n14407), .Z(n14418) );
  XOR U15442 ( .A(n14419), .B(n14420), .Z(n14407) );
  AND U15443 ( .A(n14421), .B(n14422), .Z(n14420) );
  XNOR U15444 ( .A(n14419), .B(n7212), .Z(n14422) );
  XNOR U15445 ( .A(n14415), .B(n14417), .Z(n7212) );
  NAND U15446 ( .A(n14423), .B(e_input[848]), .Z(n14417) );
  NAND U15447 ( .A(n12323), .B(e_input[848]), .Z(n14423) );
  XNOR U15448 ( .A(n14413), .B(n14424), .Z(n14415) );
  XOR U15449 ( .A(n14425), .B(n14426), .Z(n14413) );
  AND U15450 ( .A(n14427), .B(n14428), .Z(n14426) );
  XNOR U15451 ( .A(n14429), .B(n14425), .Z(n14428) );
  XOR U15452 ( .A(n14430), .B(e_input[848]), .Z(n14421) );
  IV U15453 ( .A(n14419), .Z(n14430) );
  XOR U15454 ( .A(n14431), .B(n14432), .Z(n14419) );
  AND U15455 ( .A(n14433), .B(n14434), .Z(n14432) );
  XNOR U15456 ( .A(n14431), .B(n7218), .Z(n14434) );
  XNOR U15457 ( .A(n14427), .B(n14429), .Z(n7218) );
  NAND U15458 ( .A(n14435), .B(e_input[847]), .Z(n14429) );
  NAND U15459 ( .A(n12323), .B(e_input[847]), .Z(n14435) );
  XNOR U15460 ( .A(n14425), .B(n14436), .Z(n14427) );
  XOR U15461 ( .A(n14437), .B(n14438), .Z(n14425) );
  AND U15462 ( .A(n14439), .B(n14440), .Z(n14438) );
  XNOR U15463 ( .A(n14441), .B(n14437), .Z(n14440) );
  XOR U15464 ( .A(n14442), .B(e_input[847]), .Z(n14433) );
  IV U15465 ( .A(n14431), .Z(n14442) );
  XOR U15466 ( .A(n14443), .B(n14444), .Z(n14431) );
  AND U15467 ( .A(n14445), .B(n14446), .Z(n14444) );
  XNOR U15468 ( .A(n14443), .B(n7224), .Z(n14446) );
  XNOR U15469 ( .A(n14439), .B(n14441), .Z(n7224) );
  NAND U15470 ( .A(n14447), .B(e_input[846]), .Z(n14441) );
  NAND U15471 ( .A(n12323), .B(e_input[846]), .Z(n14447) );
  XNOR U15472 ( .A(n14437), .B(n14448), .Z(n14439) );
  XOR U15473 ( .A(n14449), .B(n14450), .Z(n14437) );
  AND U15474 ( .A(n14451), .B(n14452), .Z(n14450) );
  XNOR U15475 ( .A(n14453), .B(n14449), .Z(n14452) );
  XOR U15476 ( .A(n14454), .B(e_input[846]), .Z(n14445) );
  IV U15477 ( .A(n14443), .Z(n14454) );
  XOR U15478 ( .A(n14455), .B(n14456), .Z(n14443) );
  AND U15479 ( .A(n14457), .B(n14458), .Z(n14456) );
  XNOR U15480 ( .A(n14455), .B(n7230), .Z(n14458) );
  XNOR U15481 ( .A(n14451), .B(n14453), .Z(n7230) );
  NAND U15482 ( .A(n14459), .B(e_input[845]), .Z(n14453) );
  NAND U15483 ( .A(n12323), .B(e_input[845]), .Z(n14459) );
  XNOR U15484 ( .A(n14449), .B(n14460), .Z(n14451) );
  XOR U15485 ( .A(n14461), .B(n14462), .Z(n14449) );
  AND U15486 ( .A(n14463), .B(n14464), .Z(n14462) );
  XNOR U15487 ( .A(n14465), .B(n14461), .Z(n14464) );
  XOR U15488 ( .A(n14466), .B(e_input[845]), .Z(n14457) );
  IV U15489 ( .A(n14455), .Z(n14466) );
  XOR U15490 ( .A(n14467), .B(n14468), .Z(n14455) );
  AND U15491 ( .A(n14469), .B(n14470), .Z(n14468) );
  XNOR U15492 ( .A(n14467), .B(n7236), .Z(n14470) );
  XNOR U15493 ( .A(n14463), .B(n14465), .Z(n7236) );
  NAND U15494 ( .A(n14471), .B(e_input[844]), .Z(n14465) );
  NAND U15495 ( .A(n12323), .B(e_input[844]), .Z(n14471) );
  XNOR U15496 ( .A(n14461), .B(n14472), .Z(n14463) );
  XOR U15497 ( .A(n14473), .B(n14474), .Z(n14461) );
  AND U15498 ( .A(n14475), .B(n14476), .Z(n14474) );
  XNOR U15499 ( .A(n14477), .B(n14473), .Z(n14476) );
  XOR U15500 ( .A(n14478), .B(e_input[844]), .Z(n14469) );
  IV U15501 ( .A(n14467), .Z(n14478) );
  XOR U15502 ( .A(n14479), .B(n14480), .Z(n14467) );
  AND U15503 ( .A(n14481), .B(n14482), .Z(n14480) );
  XNOR U15504 ( .A(n14479), .B(n7242), .Z(n14482) );
  XNOR U15505 ( .A(n14475), .B(n14477), .Z(n7242) );
  NAND U15506 ( .A(n14483), .B(e_input[843]), .Z(n14477) );
  NAND U15507 ( .A(n12323), .B(e_input[843]), .Z(n14483) );
  XNOR U15508 ( .A(n14473), .B(n14484), .Z(n14475) );
  XOR U15509 ( .A(n14485), .B(n14486), .Z(n14473) );
  AND U15510 ( .A(n14487), .B(n14488), .Z(n14486) );
  XNOR U15511 ( .A(n14489), .B(n14485), .Z(n14488) );
  XOR U15512 ( .A(n14490), .B(e_input[843]), .Z(n14481) );
  IV U15513 ( .A(n14479), .Z(n14490) );
  XOR U15514 ( .A(n14491), .B(n14492), .Z(n14479) );
  AND U15515 ( .A(n14493), .B(n14494), .Z(n14492) );
  XNOR U15516 ( .A(n14491), .B(n7248), .Z(n14494) );
  XNOR U15517 ( .A(n14487), .B(n14489), .Z(n7248) );
  NAND U15518 ( .A(n14495), .B(e_input[842]), .Z(n14489) );
  NAND U15519 ( .A(n12323), .B(e_input[842]), .Z(n14495) );
  XNOR U15520 ( .A(n14485), .B(n14496), .Z(n14487) );
  XOR U15521 ( .A(n14497), .B(n14498), .Z(n14485) );
  AND U15522 ( .A(n14499), .B(n14500), .Z(n14498) );
  XNOR U15523 ( .A(n14501), .B(n14497), .Z(n14500) );
  XOR U15524 ( .A(n14502), .B(e_input[842]), .Z(n14493) );
  IV U15525 ( .A(n14491), .Z(n14502) );
  XOR U15526 ( .A(n14503), .B(n14504), .Z(n14491) );
  AND U15527 ( .A(n14505), .B(n14506), .Z(n14504) );
  XNOR U15528 ( .A(n14503), .B(n7254), .Z(n14506) );
  XNOR U15529 ( .A(n14499), .B(n14501), .Z(n7254) );
  NAND U15530 ( .A(n14507), .B(e_input[841]), .Z(n14501) );
  NAND U15531 ( .A(n12323), .B(e_input[841]), .Z(n14507) );
  XNOR U15532 ( .A(n14497), .B(n14508), .Z(n14499) );
  XOR U15533 ( .A(n14509), .B(n14510), .Z(n14497) );
  AND U15534 ( .A(n14511), .B(n14512), .Z(n14510) );
  XNOR U15535 ( .A(n14513), .B(n14509), .Z(n14512) );
  XOR U15536 ( .A(n14514), .B(e_input[841]), .Z(n14505) );
  IV U15537 ( .A(n14503), .Z(n14514) );
  XOR U15538 ( .A(n14515), .B(n14516), .Z(n14503) );
  AND U15539 ( .A(n14517), .B(n14518), .Z(n14516) );
  XNOR U15540 ( .A(n14515), .B(n7260), .Z(n14518) );
  XNOR U15541 ( .A(n14511), .B(n14513), .Z(n7260) );
  NAND U15542 ( .A(n14519), .B(e_input[840]), .Z(n14513) );
  NAND U15543 ( .A(n12323), .B(e_input[840]), .Z(n14519) );
  XNOR U15544 ( .A(n14509), .B(n14520), .Z(n14511) );
  XOR U15545 ( .A(n14521), .B(n14522), .Z(n14509) );
  AND U15546 ( .A(n14523), .B(n14524), .Z(n14522) );
  XNOR U15547 ( .A(n14525), .B(n14521), .Z(n14524) );
  XOR U15548 ( .A(n14526), .B(e_input[840]), .Z(n14517) );
  IV U15549 ( .A(n14515), .Z(n14526) );
  XOR U15550 ( .A(n14527), .B(n14528), .Z(n14515) );
  AND U15551 ( .A(n14529), .B(n14530), .Z(n14528) );
  XNOR U15552 ( .A(n14527), .B(n7266), .Z(n14530) );
  XNOR U15553 ( .A(n14523), .B(n14525), .Z(n7266) );
  NAND U15554 ( .A(n14531), .B(e_input[839]), .Z(n14525) );
  NAND U15555 ( .A(n12323), .B(e_input[839]), .Z(n14531) );
  XNOR U15556 ( .A(n14521), .B(n14532), .Z(n14523) );
  XOR U15557 ( .A(n14533), .B(n14534), .Z(n14521) );
  AND U15558 ( .A(n14535), .B(n14536), .Z(n14534) );
  XNOR U15559 ( .A(n14537), .B(n14533), .Z(n14536) );
  XOR U15560 ( .A(n14538), .B(e_input[839]), .Z(n14529) );
  IV U15561 ( .A(n14527), .Z(n14538) );
  XOR U15562 ( .A(n14539), .B(n14540), .Z(n14527) );
  AND U15563 ( .A(n14541), .B(n14542), .Z(n14540) );
  XNOR U15564 ( .A(n14539), .B(n7272), .Z(n14542) );
  XNOR U15565 ( .A(n14535), .B(n14537), .Z(n7272) );
  NAND U15566 ( .A(n14543), .B(e_input[838]), .Z(n14537) );
  NAND U15567 ( .A(n12323), .B(e_input[838]), .Z(n14543) );
  XNOR U15568 ( .A(n14533), .B(n14544), .Z(n14535) );
  XOR U15569 ( .A(n14545), .B(n14546), .Z(n14533) );
  AND U15570 ( .A(n14547), .B(n14548), .Z(n14546) );
  XNOR U15571 ( .A(n14549), .B(n14545), .Z(n14548) );
  XOR U15572 ( .A(n14550), .B(e_input[838]), .Z(n14541) );
  IV U15573 ( .A(n14539), .Z(n14550) );
  XOR U15574 ( .A(n14551), .B(n14552), .Z(n14539) );
  AND U15575 ( .A(n14553), .B(n14554), .Z(n14552) );
  XNOR U15576 ( .A(n14551), .B(n7278), .Z(n14554) );
  XNOR U15577 ( .A(n14547), .B(n14549), .Z(n7278) );
  NAND U15578 ( .A(n14555), .B(e_input[837]), .Z(n14549) );
  NAND U15579 ( .A(n12323), .B(e_input[837]), .Z(n14555) );
  XNOR U15580 ( .A(n14545), .B(n14556), .Z(n14547) );
  XOR U15581 ( .A(n14557), .B(n14558), .Z(n14545) );
  AND U15582 ( .A(n14559), .B(n14560), .Z(n14558) );
  XNOR U15583 ( .A(n14561), .B(n14557), .Z(n14560) );
  XOR U15584 ( .A(n14562), .B(e_input[837]), .Z(n14553) );
  IV U15585 ( .A(n14551), .Z(n14562) );
  XOR U15586 ( .A(n14563), .B(n14564), .Z(n14551) );
  AND U15587 ( .A(n14565), .B(n14566), .Z(n14564) );
  XNOR U15588 ( .A(n14563), .B(n7284), .Z(n14566) );
  XNOR U15589 ( .A(n14559), .B(n14561), .Z(n7284) );
  NAND U15590 ( .A(n14567), .B(e_input[836]), .Z(n14561) );
  NAND U15591 ( .A(n12323), .B(e_input[836]), .Z(n14567) );
  XNOR U15592 ( .A(n14557), .B(n14568), .Z(n14559) );
  XOR U15593 ( .A(n14569), .B(n14570), .Z(n14557) );
  AND U15594 ( .A(n14571), .B(n14572), .Z(n14570) );
  XNOR U15595 ( .A(n14573), .B(n14569), .Z(n14572) );
  XOR U15596 ( .A(n14574), .B(e_input[836]), .Z(n14565) );
  IV U15597 ( .A(n14563), .Z(n14574) );
  XOR U15598 ( .A(n14575), .B(n14576), .Z(n14563) );
  AND U15599 ( .A(n14577), .B(n14578), .Z(n14576) );
  XNOR U15600 ( .A(n14575), .B(n7290), .Z(n14578) );
  XNOR U15601 ( .A(n14571), .B(n14573), .Z(n7290) );
  NAND U15602 ( .A(n14579), .B(e_input[835]), .Z(n14573) );
  NAND U15603 ( .A(n12323), .B(e_input[835]), .Z(n14579) );
  XNOR U15604 ( .A(n14569), .B(n14580), .Z(n14571) );
  XOR U15605 ( .A(n14581), .B(n14582), .Z(n14569) );
  AND U15606 ( .A(n14583), .B(n14584), .Z(n14582) );
  XNOR U15607 ( .A(n14585), .B(n14581), .Z(n14584) );
  XOR U15608 ( .A(n14586), .B(e_input[835]), .Z(n14577) );
  IV U15609 ( .A(n14575), .Z(n14586) );
  XOR U15610 ( .A(n14587), .B(n14588), .Z(n14575) );
  AND U15611 ( .A(n14589), .B(n14590), .Z(n14588) );
  XNOR U15612 ( .A(n14587), .B(n7296), .Z(n14590) );
  XNOR U15613 ( .A(n14583), .B(n14585), .Z(n7296) );
  NAND U15614 ( .A(n14591), .B(e_input[834]), .Z(n14585) );
  NAND U15615 ( .A(n12323), .B(e_input[834]), .Z(n14591) );
  XNOR U15616 ( .A(n14581), .B(n14592), .Z(n14583) );
  XOR U15617 ( .A(n14593), .B(n14594), .Z(n14581) );
  AND U15618 ( .A(n14595), .B(n14596), .Z(n14594) );
  XNOR U15619 ( .A(n14597), .B(n14593), .Z(n14596) );
  XOR U15620 ( .A(n14598), .B(e_input[834]), .Z(n14589) );
  IV U15621 ( .A(n14587), .Z(n14598) );
  XOR U15622 ( .A(n14599), .B(n14600), .Z(n14587) );
  AND U15623 ( .A(n14601), .B(n14602), .Z(n14600) );
  XNOR U15624 ( .A(n14599), .B(n7302), .Z(n14602) );
  XNOR U15625 ( .A(n14595), .B(n14597), .Z(n7302) );
  NAND U15626 ( .A(n14603), .B(e_input[833]), .Z(n14597) );
  NAND U15627 ( .A(n12323), .B(e_input[833]), .Z(n14603) );
  XNOR U15628 ( .A(n14593), .B(n14604), .Z(n14595) );
  XOR U15629 ( .A(n14605), .B(n14606), .Z(n14593) );
  AND U15630 ( .A(n14607), .B(n14608), .Z(n14606) );
  XNOR U15631 ( .A(n14609), .B(n14605), .Z(n14608) );
  XOR U15632 ( .A(n14610), .B(e_input[833]), .Z(n14601) );
  IV U15633 ( .A(n14599), .Z(n14610) );
  XOR U15634 ( .A(n14611), .B(n14612), .Z(n14599) );
  AND U15635 ( .A(n14613), .B(n14614), .Z(n14612) );
  XNOR U15636 ( .A(n14611), .B(n7308), .Z(n14614) );
  XNOR U15637 ( .A(n14607), .B(n14609), .Z(n7308) );
  NAND U15638 ( .A(n14615), .B(e_input[832]), .Z(n14609) );
  NAND U15639 ( .A(n12323), .B(e_input[832]), .Z(n14615) );
  XNOR U15640 ( .A(n14605), .B(n14616), .Z(n14607) );
  XOR U15641 ( .A(n14617), .B(n14618), .Z(n14605) );
  AND U15642 ( .A(n14619), .B(n14620), .Z(n14618) );
  XNOR U15643 ( .A(n14621), .B(n14617), .Z(n14620) );
  XOR U15644 ( .A(n14622), .B(e_input[832]), .Z(n14613) );
  IV U15645 ( .A(n14611), .Z(n14622) );
  XOR U15646 ( .A(n14623), .B(n14624), .Z(n14611) );
  AND U15647 ( .A(n14625), .B(n14626), .Z(n14624) );
  XNOR U15648 ( .A(n14623), .B(n7314), .Z(n14626) );
  XNOR U15649 ( .A(n14619), .B(n14621), .Z(n7314) );
  NAND U15650 ( .A(n14627), .B(e_input[831]), .Z(n14621) );
  NAND U15651 ( .A(n12323), .B(e_input[831]), .Z(n14627) );
  XNOR U15652 ( .A(n14617), .B(n14628), .Z(n14619) );
  XOR U15653 ( .A(n14629), .B(n14630), .Z(n14617) );
  AND U15654 ( .A(n14631), .B(n14632), .Z(n14630) );
  XNOR U15655 ( .A(n14633), .B(n14629), .Z(n14632) );
  XOR U15656 ( .A(n14634), .B(e_input[831]), .Z(n14625) );
  IV U15657 ( .A(n14623), .Z(n14634) );
  XOR U15658 ( .A(n14635), .B(n14636), .Z(n14623) );
  AND U15659 ( .A(n14637), .B(n14638), .Z(n14636) );
  XNOR U15660 ( .A(n14635), .B(n7320), .Z(n14638) );
  XNOR U15661 ( .A(n14631), .B(n14633), .Z(n7320) );
  NAND U15662 ( .A(n14639), .B(e_input[830]), .Z(n14633) );
  NAND U15663 ( .A(n12323), .B(e_input[830]), .Z(n14639) );
  XNOR U15664 ( .A(n14629), .B(n14640), .Z(n14631) );
  XOR U15665 ( .A(n14641), .B(n14642), .Z(n14629) );
  AND U15666 ( .A(n14643), .B(n14644), .Z(n14642) );
  XNOR U15667 ( .A(n14645), .B(n14641), .Z(n14644) );
  XOR U15668 ( .A(n14646), .B(e_input[830]), .Z(n14637) );
  IV U15669 ( .A(n14635), .Z(n14646) );
  XOR U15670 ( .A(n14647), .B(n14648), .Z(n14635) );
  AND U15671 ( .A(n14649), .B(n14650), .Z(n14648) );
  XNOR U15672 ( .A(n14647), .B(n7326), .Z(n14650) );
  XNOR U15673 ( .A(n14643), .B(n14645), .Z(n7326) );
  NAND U15674 ( .A(n14651), .B(e_input[829]), .Z(n14645) );
  NAND U15675 ( .A(n12323), .B(e_input[829]), .Z(n14651) );
  XNOR U15676 ( .A(n14641), .B(n14652), .Z(n14643) );
  XOR U15677 ( .A(n14653), .B(n14654), .Z(n14641) );
  AND U15678 ( .A(n14655), .B(n14656), .Z(n14654) );
  XNOR U15679 ( .A(n14657), .B(n14653), .Z(n14656) );
  XOR U15680 ( .A(n14658), .B(e_input[829]), .Z(n14649) );
  IV U15681 ( .A(n14647), .Z(n14658) );
  XOR U15682 ( .A(n14659), .B(n14660), .Z(n14647) );
  AND U15683 ( .A(n14661), .B(n14662), .Z(n14660) );
  XNOR U15684 ( .A(n14659), .B(n7332), .Z(n14662) );
  XNOR U15685 ( .A(n14655), .B(n14657), .Z(n7332) );
  NAND U15686 ( .A(n14663), .B(e_input[828]), .Z(n14657) );
  NAND U15687 ( .A(n12323), .B(e_input[828]), .Z(n14663) );
  XNOR U15688 ( .A(n14653), .B(n14664), .Z(n14655) );
  XOR U15689 ( .A(n14665), .B(n14666), .Z(n14653) );
  AND U15690 ( .A(n14667), .B(n14668), .Z(n14666) );
  XNOR U15691 ( .A(n14669), .B(n14665), .Z(n14668) );
  XOR U15692 ( .A(n14670), .B(e_input[828]), .Z(n14661) );
  IV U15693 ( .A(n14659), .Z(n14670) );
  XOR U15694 ( .A(n14671), .B(n14672), .Z(n14659) );
  AND U15695 ( .A(n14673), .B(n14674), .Z(n14672) );
  XNOR U15696 ( .A(n14671), .B(n7338), .Z(n14674) );
  XNOR U15697 ( .A(n14667), .B(n14669), .Z(n7338) );
  NAND U15698 ( .A(n14675), .B(e_input[827]), .Z(n14669) );
  NAND U15699 ( .A(n12323), .B(e_input[827]), .Z(n14675) );
  XNOR U15700 ( .A(n14665), .B(n14676), .Z(n14667) );
  XOR U15701 ( .A(n14677), .B(n14678), .Z(n14665) );
  AND U15702 ( .A(n14679), .B(n14680), .Z(n14678) );
  XNOR U15703 ( .A(n14681), .B(n14677), .Z(n14680) );
  XOR U15704 ( .A(n14682), .B(e_input[827]), .Z(n14673) );
  IV U15705 ( .A(n14671), .Z(n14682) );
  XOR U15706 ( .A(n14683), .B(n14684), .Z(n14671) );
  AND U15707 ( .A(n14685), .B(n14686), .Z(n14684) );
  XNOR U15708 ( .A(n14683), .B(n7344), .Z(n14686) );
  XNOR U15709 ( .A(n14679), .B(n14681), .Z(n7344) );
  NAND U15710 ( .A(n14687), .B(e_input[826]), .Z(n14681) );
  NAND U15711 ( .A(n12323), .B(e_input[826]), .Z(n14687) );
  XNOR U15712 ( .A(n14677), .B(n14688), .Z(n14679) );
  XOR U15713 ( .A(n14689), .B(n14690), .Z(n14677) );
  AND U15714 ( .A(n14691), .B(n14692), .Z(n14690) );
  XNOR U15715 ( .A(n14693), .B(n14689), .Z(n14692) );
  XOR U15716 ( .A(n14694), .B(e_input[826]), .Z(n14685) );
  IV U15717 ( .A(n14683), .Z(n14694) );
  XOR U15718 ( .A(n14695), .B(n14696), .Z(n14683) );
  AND U15719 ( .A(n14697), .B(n14698), .Z(n14696) );
  XNOR U15720 ( .A(n14695), .B(n7350), .Z(n14698) );
  XNOR U15721 ( .A(n14691), .B(n14693), .Z(n7350) );
  NAND U15722 ( .A(n14699), .B(e_input[825]), .Z(n14693) );
  NAND U15723 ( .A(n12323), .B(e_input[825]), .Z(n14699) );
  XNOR U15724 ( .A(n14689), .B(n14700), .Z(n14691) );
  XOR U15725 ( .A(n14701), .B(n14702), .Z(n14689) );
  AND U15726 ( .A(n14703), .B(n14704), .Z(n14702) );
  XNOR U15727 ( .A(n14705), .B(n14701), .Z(n14704) );
  XOR U15728 ( .A(n14706), .B(e_input[825]), .Z(n14697) );
  IV U15729 ( .A(n14695), .Z(n14706) );
  XOR U15730 ( .A(n14707), .B(n14708), .Z(n14695) );
  AND U15731 ( .A(n14709), .B(n14710), .Z(n14708) );
  XNOR U15732 ( .A(n14707), .B(n7356), .Z(n14710) );
  XNOR U15733 ( .A(n14703), .B(n14705), .Z(n7356) );
  NAND U15734 ( .A(n14711), .B(e_input[824]), .Z(n14705) );
  NAND U15735 ( .A(n12323), .B(e_input[824]), .Z(n14711) );
  XNOR U15736 ( .A(n14701), .B(n14712), .Z(n14703) );
  XOR U15737 ( .A(n14713), .B(n14714), .Z(n14701) );
  AND U15738 ( .A(n14715), .B(n14716), .Z(n14714) );
  XNOR U15739 ( .A(n14717), .B(n14713), .Z(n14716) );
  XOR U15740 ( .A(n14718), .B(e_input[824]), .Z(n14709) );
  IV U15741 ( .A(n14707), .Z(n14718) );
  XOR U15742 ( .A(n14719), .B(n14720), .Z(n14707) );
  AND U15743 ( .A(n14721), .B(n14722), .Z(n14720) );
  XNOR U15744 ( .A(n14719), .B(n7362), .Z(n14722) );
  XNOR U15745 ( .A(n14715), .B(n14717), .Z(n7362) );
  NAND U15746 ( .A(n14723), .B(e_input[823]), .Z(n14717) );
  NAND U15747 ( .A(n12323), .B(e_input[823]), .Z(n14723) );
  XNOR U15748 ( .A(n14713), .B(n14724), .Z(n14715) );
  XOR U15749 ( .A(n14725), .B(n14726), .Z(n14713) );
  AND U15750 ( .A(n14727), .B(n14728), .Z(n14726) );
  XNOR U15751 ( .A(n14729), .B(n14725), .Z(n14728) );
  XOR U15752 ( .A(n14730), .B(e_input[823]), .Z(n14721) );
  IV U15753 ( .A(n14719), .Z(n14730) );
  XOR U15754 ( .A(n14731), .B(n14732), .Z(n14719) );
  AND U15755 ( .A(n14733), .B(n14734), .Z(n14732) );
  XNOR U15756 ( .A(n14731), .B(n7368), .Z(n14734) );
  XNOR U15757 ( .A(n14727), .B(n14729), .Z(n7368) );
  NAND U15758 ( .A(n14735), .B(e_input[822]), .Z(n14729) );
  NAND U15759 ( .A(n12323), .B(e_input[822]), .Z(n14735) );
  XNOR U15760 ( .A(n14725), .B(n14736), .Z(n14727) );
  XOR U15761 ( .A(n14737), .B(n14738), .Z(n14725) );
  AND U15762 ( .A(n14739), .B(n14740), .Z(n14738) );
  XNOR U15763 ( .A(n14741), .B(n14737), .Z(n14740) );
  XOR U15764 ( .A(n14742), .B(e_input[822]), .Z(n14733) );
  IV U15765 ( .A(n14731), .Z(n14742) );
  XOR U15766 ( .A(n14743), .B(n14744), .Z(n14731) );
  AND U15767 ( .A(n14745), .B(n14746), .Z(n14744) );
  XNOR U15768 ( .A(n14743), .B(n7374), .Z(n14746) );
  XNOR U15769 ( .A(n14739), .B(n14741), .Z(n7374) );
  NAND U15770 ( .A(n14747), .B(e_input[821]), .Z(n14741) );
  NAND U15771 ( .A(n12323), .B(e_input[821]), .Z(n14747) );
  XNOR U15772 ( .A(n14737), .B(n14748), .Z(n14739) );
  XOR U15773 ( .A(n14749), .B(n14750), .Z(n14737) );
  AND U15774 ( .A(n14751), .B(n14752), .Z(n14750) );
  XNOR U15775 ( .A(n14753), .B(n14749), .Z(n14752) );
  XOR U15776 ( .A(n14754), .B(e_input[821]), .Z(n14745) );
  IV U15777 ( .A(n14743), .Z(n14754) );
  XOR U15778 ( .A(n14755), .B(n14756), .Z(n14743) );
  AND U15779 ( .A(n14757), .B(n14758), .Z(n14756) );
  XNOR U15780 ( .A(n14755), .B(n7380), .Z(n14758) );
  XNOR U15781 ( .A(n14751), .B(n14753), .Z(n7380) );
  NAND U15782 ( .A(n14759), .B(e_input[820]), .Z(n14753) );
  NAND U15783 ( .A(n12323), .B(e_input[820]), .Z(n14759) );
  XNOR U15784 ( .A(n14749), .B(n14760), .Z(n14751) );
  XOR U15785 ( .A(n14761), .B(n14762), .Z(n14749) );
  AND U15786 ( .A(n14763), .B(n14764), .Z(n14762) );
  XNOR U15787 ( .A(n14765), .B(n14761), .Z(n14764) );
  XOR U15788 ( .A(n14766), .B(e_input[820]), .Z(n14757) );
  IV U15789 ( .A(n14755), .Z(n14766) );
  XOR U15790 ( .A(n14767), .B(n14768), .Z(n14755) );
  AND U15791 ( .A(n14769), .B(n14770), .Z(n14768) );
  XNOR U15792 ( .A(n14767), .B(n7386), .Z(n14770) );
  XNOR U15793 ( .A(n14763), .B(n14765), .Z(n7386) );
  NAND U15794 ( .A(n14771), .B(e_input[819]), .Z(n14765) );
  NAND U15795 ( .A(n12323), .B(e_input[819]), .Z(n14771) );
  XNOR U15796 ( .A(n14761), .B(n14772), .Z(n14763) );
  XOR U15797 ( .A(n14773), .B(n14774), .Z(n14761) );
  AND U15798 ( .A(n14775), .B(n14776), .Z(n14774) );
  XNOR U15799 ( .A(n14777), .B(n14773), .Z(n14776) );
  XOR U15800 ( .A(n14778), .B(e_input[819]), .Z(n14769) );
  IV U15801 ( .A(n14767), .Z(n14778) );
  XOR U15802 ( .A(n14779), .B(n14780), .Z(n14767) );
  AND U15803 ( .A(n14781), .B(n14782), .Z(n14780) );
  XNOR U15804 ( .A(n14779), .B(n7392), .Z(n14782) );
  XNOR U15805 ( .A(n14775), .B(n14777), .Z(n7392) );
  NAND U15806 ( .A(n14783), .B(e_input[818]), .Z(n14777) );
  NAND U15807 ( .A(n12323), .B(e_input[818]), .Z(n14783) );
  XNOR U15808 ( .A(n14773), .B(n14784), .Z(n14775) );
  XOR U15809 ( .A(n14785), .B(n14786), .Z(n14773) );
  AND U15810 ( .A(n14787), .B(n14788), .Z(n14786) );
  XNOR U15811 ( .A(n14789), .B(n14785), .Z(n14788) );
  XOR U15812 ( .A(n14790), .B(e_input[818]), .Z(n14781) );
  IV U15813 ( .A(n14779), .Z(n14790) );
  XOR U15814 ( .A(n14791), .B(n14792), .Z(n14779) );
  AND U15815 ( .A(n14793), .B(n14794), .Z(n14792) );
  XNOR U15816 ( .A(n14791), .B(n7398), .Z(n14794) );
  XNOR U15817 ( .A(n14787), .B(n14789), .Z(n7398) );
  NAND U15818 ( .A(n14795), .B(e_input[817]), .Z(n14789) );
  NAND U15819 ( .A(n12323), .B(e_input[817]), .Z(n14795) );
  XNOR U15820 ( .A(n14785), .B(n14796), .Z(n14787) );
  XOR U15821 ( .A(n14797), .B(n14798), .Z(n14785) );
  AND U15822 ( .A(n14799), .B(n14800), .Z(n14798) );
  XNOR U15823 ( .A(n14801), .B(n14797), .Z(n14800) );
  XOR U15824 ( .A(n14802), .B(e_input[817]), .Z(n14793) );
  IV U15825 ( .A(n14791), .Z(n14802) );
  XOR U15826 ( .A(n14803), .B(n14804), .Z(n14791) );
  AND U15827 ( .A(n14805), .B(n14806), .Z(n14804) );
  XNOR U15828 ( .A(n14803), .B(n7404), .Z(n14806) );
  XNOR U15829 ( .A(n14799), .B(n14801), .Z(n7404) );
  NAND U15830 ( .A(n14807), .B(e_input[816]), .Z(n14801) );
  NAND U15831 ( .A(n12323), .B(e_input[816]), .Z(n14807) );
  XNOR U15832 ( .A(n14797), .B(n14808), .Z(n14799) );
  XOR U15833 ( .A(n14809), .B(n14810), .Z(n14797) );
  AND U15834 ( .A(n14811), .B(n14812), .Z(n14810) );
  XNOR U15835 ( .A(n14813), .B(n14809), .Z(n14812) );
  XOR U15836 ( .A(n14814), .B(e_input[816]), .Z(n14805) );
  IV U15837 ( .A(n14803), .Z(n14814) );
  XOR U15838 ( .A(n14815), .B(n14816), .Z(n14803) );
  AND U15839 ( .A(n14817), .B(n14818), .Z(n14816) );
  XNOR U15840 ( .A(n14815), .B(n7410), .Z(n14818) );
  XNOR U15841 ( .A(n14811), .B(n14813), .Z(n7410) );
  NAND U15842 ( .A(n14819), .B(e_input[815]), .Z(n14813) );
  NAND U15843 ( .A(n12323), .B(e_input[815]), .Z(n14819) );
  XNOR U15844 ( .A(n14809), .B(n14820), .Z(n14811) );
  XOR U15845 ( .A(n14821), .B(n14822), .Z(n14809) );
  AND U15846 ( .A(n14823), .B(n14824), .Z(n14822) );
  XNOR U15847 ( .A(n14825), .B(n14821), .Z(n14824) );
  XOR U15848 ( .A(n14826), .B(e_input[815]), .Z(n14817) );
  IV U15849 ( .A(n14815), .Z(n14826) );
  XOR U15850 ( .A(n14827), .B(n14828), .Z(n14815) );
  AND U15851 ( .A(n14829), .B(n14830), .Z(n14828) );
  XNOR U15852 ( .A(n14827), .B(n7416), .Z(n14830) );
  XNOR U15853 ( .A(n14823), .B(n14825), .Z(n7416) );
  NAND U15854 ( .A(n14831), .B(e_input[814]), .Z(n14825) );
  NAND U15855 ( .A(n12323), .B(e_input[814]), .Z(n14831) );
  XNOR U15856 ( .A(n14821), .B(n14832), .Z(n14823) );
  XOR U15857 ( .A(n14833), .B(n14834), .Z(n14821) );
  AND U15858 ( .A(n14835), .B(n14836), .Z(n14834) );
  XNOR U15859 ( .A(n14837), .B(n14833), .Z(n14836) );
  XOR U15860 ( .A(n14838), .B(e_input[814]), .Z(n14829) );
  IV U15861 ( .A(n14827), .Z(n14838) );
  XOR U15862 ( .A(n14839), .B(n14840), .Z(n14827) );
  AND U15863 ( .A(n14841), .B(n14842), .Z(n14840) );
  XNOR U15864 ( .A(n14839), .B(n7422), .Z(n14842) );
  XNOR U15865 ( .A(n14835), .B(n14837), .Z(n7422) );
  NAND U15866 ( .A(n14843), .B(e_input[813]), .Z(n14837) );
  NAND U15867 ( .A(n12323), .B(e_input[813]), .Z(n14843) );
  XNOR U15868 ( .A(n14833), .B(n14844), .Z(n14835) );
  XOR U15869 ( .A(n14845), .B(n14846), .Z(n14833) );
  AND U15870 ( .A(n14847), .B(n14848), .Z(n14846) );
  XNOR U15871 ( .A(n14849), .B(n14845), .Z(n14848) );
  XOR U15872 ( .A(n14850), .B(e_input[813]), .Z(n14841) );
  IV U15873 ( .A(n14839), .Z(n14850) );
  XOR U15874 ( .A(n14851), .B(n14852), .Z(n14839) );
  AND U15875 ( .A(n14853), .B(n14854), .Z(n14852) );
  XNOR U15876 ( .A(n14851), .B(n7428), .Z(n14854) );
  XNOR U15877 ( .A(n14847), .B(n14849), .Z(n7428) );
  NAND U15878 ( .A(n14855), .B(e_input[812]), .Z(n14849) );
  NAND U15879 ( .A(n12323), .B(e_input[812]), .Z(n14855) );
  XNOR U15880 ( .A(n14845), .B(n14856), .Z(n14847) );
  XOR U15881 ( .A(n14857), .B(n14858), .Z(n14845) );
  AND U15882 ( .A(n14859), .B(n14860), .Z(n14858) );
  XNOR U15883 ( .A(n14861), .B(n14857), .Z(n14860) );
  XOR U15884 ( .A(n14862), .B(e_input[812]), .Z(n14853) );
  IV U15885 ( .A(n14851), .Z(n14862) );
  XOR U15886 ( .A(n14863), .B(n14864), .Z(n14851) );
  AND U15887 ( .A(n14865), .B(n14866), .Z(n14864) );
  XNOR U15888 ( .A(n14863), .B(n7434), .Z(n14866) );
  XNOR U15889 ( .A(n14859), .B(n14861), .Z(n7434) );
  NAND U15890 ( .A(n14867), .B(e_input[811]), .Z(n14861) );
  NAND U15891 ( .A(n12323), .B(e_input[811]), .Z(n14867) );
  XNOR U15892 ( .A(n14857), .B(n14868), .Z(n14859) );
  XOR U15893 ( .A(n14869), .B(n14870), .Z(n14857) );
  AND U15894 ( .A(n14871), .B(n14872), .Z(n14870) );
  XNOR U15895 ( .A(n14873), .B(n14869), .Z(n14872) );
  XOR U15896 ( .A(n14874), .B(e_input[811]), .Z(n14865) );
  IV U15897 ( .A(n14863), .Z(n14874) );
  XOR U15898 ( .A(n14875), .B(n14876), .Z(n14863) );
  AND U15899 ( .A(n14877), .B(n14878), .Z(n14876) );
  XNOR U15900 ( .A(n14875), .B(n7440), .Z(n14878) );
  XNOR U15901 ( .A(n14871), .B(n14873), .Z(n7440) );
  NAND U15902 ( .A(n14879), .B(e_input[810]), .Z(n14873) );
  NAND U15903 ( .A(n12323), .B(e_input[810]), .Z(n14879) );
  XNOR U15904 ( .A(n14869), .B(n14880), .Z(n14871) );
  XOR U15905 ( .A(n14881), .B(n14882), .Z(n14869) );
  AND U15906 ( .A(n14883), .B(n14884), .Z(n14882) );
  XNOR U15907 ( .A(n14885), .B(n14881), .Z(n14884) );
  XOR U15908 ( .A(n14886), .B(e_input[810]), .Z(n14877) );
  IV U15909 ( .A(n14875), .Z(n14886) );
  XOR U15910 ( .A(n14887), .B(n14888), .Z(n14875) );
  AND U15911 ( .A(n14889), .B(n14890), .Z(n14888) );
  XNOR U15912 ( .A(n14887), .B(n7446), .Z(n14890) );
  XNOR U15913 ( .A(n14883), .B(n14885), .Z(n7446) );
  NAND U15914 ( .A(n14891), .B(e_input[809]), .Z(n14885) );
  NAND U15915 ( .A(n12323), .B(e_input[809]), .Z(n14891) );
  XNOR U15916 ( .A(n14881), .B(n14892), .Z(n14883) );
  XOR U15917 ( .A(n14893), .B(n14894), .Z(n14881) );
  AND U15918 ( .A(n14895), .B(n14896), .Z(n14894) );
  XNOR U15919 ( .A(n14897), .B(n14893), .Z(n14896) );
  XOR U15920 ( .A(n14898), .B(e_input[809]), .Z(n14889) );
  IV U15921 ( .A(n14887), .Z(n14898) );
  XOR U15922 ( .A(n14899), .B(n14900), .Z(n14887) );
  AND U15923 ( .A(n14901), .B(n14902), .Z(n14900) );
  XNOR U15924 ( .A(n14899), .B(n7452), .Z(n14902) );
  XNOR U15925 ( .A(n14895), .B(n14897), .Z(n7452) );
  NAND U15926 ( .A(n14903), .B(e_input[808]), .Z(n14897) );
  NAND U15927 ( .A(n12323), .B(e_input[808]), .Z(n14903) );
  XNOR U15928 ( .A(n14893), .B(n14904), .Z(n14895) );
  XOR U15929 ( .A(n14905), .B(n14906), .Z(n14893) );
  AND U15930 ( .A(n14907), .B(n14908), .Z(n14906) );
  XNOR U15931 ( .A(n14909), .B(n14905), .Z(n14908) );
  XOR U15932 ( .A(n14910), .B(e_input[808]), .Z(n14901) );
  IV U15933 ( .A(n14899), .Z(n14910) );
  XOR U15934 ( .A(n14911), .B(n14912), .Z(n14899) );
  AND U15935 ( .A(n14913), .B(n14914), .Z(n14912) );
  XNOR U15936 ( .A(n14911), .B(n7458), .Z(n14914) );
  XNOR U15937 ( .A(n14907), .B(n14909), .Z(n7458) );
  NAND U15938 ( .A(n14915), .B(e_input[807]), .Z(n14909) );
  NAND U15939 ( .A(n12323), .B(e_input[807]), .Z(n14915) );
  XNOR U15940 ( .A(n14905), .B(n14916), .Z(n14907) );
  XOR U15941 ( .A(n14917), .B(n14918), .Z(n14905) );
  AND U15942 ( .A(n14919), .B(n14920), .Z(n14918) );
  XNOR U15943 ( .A(n14921), .B(n14917), .Z(n14920) );
  XOR U15944 ( .A(n14922), .B(e_input[807]), .Z(n14913) );
  IV U15945 ( .A(n14911), .Z(n14922) );
  XOR U15946 ( .A(n14923), .B(n14924), .Z(n14911) );
  AND U15947 ( .A(n14925), .B(n14926), .Z(n14924) );
  XNOR U15948 ( .A(n14923), .B(n7464), .Z(n14926) );
  XNOR U15949 ( .A(n14919), .B(n14921), .Z(n7464) );
  NAND U15950 ( .A(n14927), .B(e_input[806]), .Z(n14921) );
  NAND U15951 ( .A(n12323), .B(e_input[806]), .Z(n14927) );
  XNOR U15952 ( .A(n14917), .B(n14928), .Z(n14919) );
  XOR U15953 ( .A(n14929), .B(n14930), .Z(n14917) );
  AND U15954 ( .A(n14931), .B(n14932), .Z(n14930) );
  XNOR U15955 ( .A(n14933), .B(n14929), .Z(n14932) );
  XOR U15956 ( .A(n14934), .B(e_input[806]), .Z(n14925) );
  IV U15957 ( .A(n14923), .Z(n14934) );
  XOR U15958 ( .A(n14935), .B(n14936), .Z(n14923) );
  AND U15959 ( .A(n14937), .B(n14938), .Z(n14936) );
  XNOR U15960 ( .A(n14935), .B(n7470), .Z(n14938) );
  XNOR U15961 ( .A(n14931), .B(n14933), .Z(n7470) );
  NAND U15962 ( .A(n14939), .B(e_input[805]), .Z(n14933) );
  NAND U15963 ( .A(n12323), .B(e_input[805]), .Z(n14939) );
  XNOR U15964 ( .A(n14929), .B(n14940), .Z(n14931) );
  XOR U15965 ( .A(n14941), .B(n14942), .Z(n14929) );
  AND U15966 ( .A(n14943), .B(n14944), .Z(n14942) );
  XNOR U15967 ( .A(n14945), .B(n14941), .Z(n14944) );
  XOR U15968 ( .A(n14946), .B(e_input[805]), .Z(n14937) );
  IV U15969 ( .A(n14935), .Z(n14946) );
  XOR U15970 ( .A(n14947), .B(n14948), .Z(n14935) );
  AND U15971 ( .A(n14949), .B(n14950), .Z(n14948) );
  XNOR U15972 ( .A(n14947), .B(n7476), .Z(n14950) );
  XNOR U15973 ( .A(n14943), .B(n14945), .Z(n7476) );
  NAND U15974 ( .A(n14951), .B(e_input[804]), .Z(n14945) );
  NAND U15975 ( .A(n12323), .B(e_input[804]), .Z(n14951) );
  XNOR U15976 ( .A(n14941), .B(n14952), .Z(n14943) );
  XOR U15977 ( .A(n14953), .B(n14954), .Z(n14941) );
  AND U15978 ( .A(n14955), .B(n14956), .Z(n14954) );
  XNOR U15979 ( .A(n14957), .B(n14953), .Z(n14956) );
  XOR U15980 ( .A(n14958), .B(e_input[804]), .Z(n14949) );
  IV U15981 ( .A(n14947), .Z(n14958) );
  XOR U15982 ( .A(n14959), .B(n14960), .Z(n14947) );
  AND U15983 ( .A(n14961), .B(n14962), .Z(n14960) );
  XNOR U15984 ( .A(n14959), .B(n7482), .Z(n14962) );
  XNOR U15985 ( .A(n14955), .B(n14957), .Z(n7482) );
  NAND U15986 ( .A(n14963), .B(e_input[803]), .Z(n14957) );
  NAND U15987 ( .A(n12323), .B(e_input[803]), .Z(n14963) );
  XNOR U15988 ( .A(n14953), .B(n14964), .Z(n14955) );
  XOR U15989 ( .A(n14965), .B(n14966), .Z(n14953) );
  AND U15990 ( .A(n14967), .B(n14968), .Z(n14966) );
  XNOR U15991 ( .A(n14969), .B(n14965), .Z(n14968) );
  XOR U15992 ( .A(n14970), .B(e_input[803]), .Z(n14961) );
  IV U15993 ( .A(n14959), .Z(n14970) );
  XOR U15994 ( .A(n14971), .B(n14972), .Z(n14959) );
  AND U15995 ( .A(n14973), .B(n14974), .Z(n14972) );
  XNOR U15996 ( .A(n14971), .B(n7488), .Z(n14974) );
  XNOR U15997 ( .A(n14967), .B(n14969), .Z(n7488) );
  NAND U15998 ( .A(n14975), .B(e_input[802]), .Z(n14969) );
  NAND U15999 ( .A(n12323), .B(e_input[802]), .Z(n14975) );
  XNOR U16000 ( .A(n14965), .B(n14976), .Z(n14967) );
  XOR U16001 ( .A(n14977), .B(n14978), .Z(n14965) );
  AND U16002 ( .A(n14979), .B(n14980), .Z(n14978) );
  XNOR U16003 ( .A(n14981), .B(n14977), .Z(n14980) );
  XOR U16004 ( .A(n14982), .B(e_input[802]), .Z(n14973) );
  IV U16005 ( .A(n14971), .Z(n14982) );
  XOR U16006 ( .A(n14983), .B(n14984), .Z(n14971) );
  AND U16007 ( .A(n14985), .B(n14986), .Z(n14984) );
  XNOR U16008 ( .A(n14983), .B(n7494), .Z(n14986) );
  XNOR U16009 ( .A(n14979), .B(n14981), .Z(n7494) );
  NAND U16010 ( .A(n14987), .B(e_input[801]), .Z(n14981) );
  NAND U16011 ( .A(n12323), .B(e_input[801]), .Z(n14987) );
  XNOR U16012 ( .A(n14977), .B(n14988), .Z(n14979) );
  XOR U16013 ( .A(n14989), .B(n14990), .Z(n14977) );
  AND U16014 ( .A(n14991), .B(n14992), .Z(n14990) );
  XNOR U16015 ( .A(n14993), .B(n14989), .Z(n14992) );
  XOR U16016 ( .A(n14994), .B(e_input[801]), .Z(n14985) );
  IV U16017 ( .A(n14983), .Z(n14994) );
  XOR U16018 ( .A(n14995), .B(n14996), .Z(n14983) );
  AND U16019 ( .A(n14997), .B(n14998), .Z(n14996) );
  XNOR U16020 ( .A(n14995), .B(n7500), .Z(n14998) );
  XNOR U16021 ( .A(n14991), .B(n14993), .Z(n7500) );
  NAND U16022 ( .A(n14999), .B(e_input[800]), .Z(n14993) );
  NAND U16023 ( .A(n12323), .B(e_input[800]), .Z(n14999) );
  XNOR U16024 ( .A(n14989), .B(n15000), .Z(n14991) );
  XOR U16025 ( .A(n15001), .B(n15002), .Z(n14989) );
  AND U16026 ( .A(n15003), .B(n15004), .Z(n15002) );
  XNOR U16027 ( .A(n15005), .B(n15001), .Z(n15004) );
  XOR U16028 ( .A(n15006), .B(e_input[800]), .Z(n14997) );
  IV U16029 ( .A(n14995), .Z(n15006) );
  XOR U16030 ( .A(n15007), .B(n15008), .Z(n14995) );
  AND U16031 ( .A(n15009), .B(n15010), .Z(n15008) );
  XNOR U16032 ( .A(n15007), .B(n7506), .Z(n15010) );
  XNOR U16033 ( .A(n15003), .B(n15005), .Z(n7506) );
  NAND U16034 ( .A(n15011), .B(e_input[799]), .Z(n15005) );
  NAND U16035 ( .A(n12323), .B(e_input[799]), .Z(n15011) );
  XNOR U16036 ( .A(n15001), .B(n15012), .Z(n15003) );
  XOR U16037 ( .A(n15013), .B(n15014), .Z(n15001) );
  AND U16038 ( .A(n15015), .B(n15016), .Z(n15014) );
  XNOR U16039 ( .A(n15017), .B(n15013), .Z(n15016) );
  XOR U16040 ( .A(n15018), .B(e_input[799]), .Z(n15009) );
  IV U16041 ( .A(n15007), .Z(n15018) );
  XOR U16042 ( .A(n15019), .B(n15020), .Z(n15007) );
  AND U16043 ( .A(n15021), .B(n15022), .Z(n15020) );
  XNOR U16044 ( .A(n15019), .B(n7512), .Z(n15022) );
  XNOR U16045 ( .A(n15015), .B(n15017), .Z(n7512) );
  NAND U16046 ( .A(n15023), .B(e_input[798]), .Z(n15017) );
  NAND U16047 ( .A(n12323), .B(e_input[798]), .Z(n15023) );
  XNOR U16048 ( .A(n15013), .B(n15024), .Z(n15015) );
  XOR U16049 ( .A(n15025), .B(n15026), .Z(n15013) );
  AND U16050 ( .A(n15027), .B(n15028), .Z(n15026) );
  XNOR U16051 ( .A(n15029), .B(n15025), .Z(n15028) );
  XOR U16052 ( .A(n15030), .B(e_input[798]), .Z(n15021) );
  IV U16053 ( .A(n15019), .Z(n15030) );
  XOR U16054 ( .A(n15031), .B(n15032), .Z(n15019) );
  AND U16055 ( .A(n15033), .B(n15034), .Z(n15032) );
  XNOR U16056 ( .A(n15031), .B(n7518), .Z(n15034) );
  XNOR U16057 ( .A(n15027), .B(n15029), .Z(n7518) );
  NAND U16058 ( .A(n15035), .B(e_input[797]), .Z(n15029) );
  NAND U16059 ( .A(n12323), .B(e_input[797]), .Z(n15035) );
  XNOR U16060 ( .A(n15025), .B(n15036), .Z(n15027) );
  XOR U16061 ( .A(n15037), .B(n15038), .Z(n15025) );
  AND U16062 ( .A(n15039), .B(n15040), .Z(n15038) );
  XNOR U16063 ( .A(n15041), .B(n15037), .Z(n15040) );
  XOR U16064 ( .A(n15042), .B(e_input[797]), .Z(n15033) );
  IV U16065 ( .A(n15031), .Z(n15042) );
  XOR U16066 ( .A(n15043), .B(n15044), .Z(n15031) );
  AND U16067 ( .A(n15045), .B(n15046), .Z(n15044) );
  XNOR U16068 ( .A(n15043), .B(n7524), .Z(n15046) );
  XNOR U16069 ( .A(n15039), .B(n15041), .Z(n7524) );
  NAND U16070 ( .A(n15047), .B(e_input[796]), .Z(n15041) );
  NAND U16071 ( .A(n12323), .B(e_input[796]), .Z(n15047) );
  XNOR U16072 ( .A(n15037), .B(n15048), .Z(n15039) );
  XOR U16073 ( .A(n15049), .B(n15050), .Z(n15037) );
  AND U16074 ( .A(n15051), .B(n15052), .Z(n15050) );
  XNOR U16075 ( .A(n15053), .B(n15049), .Z(n15052) );
  XOR U16076 ( .A(n15054), .B(e_input[796]), .Z(n15045) );
  IV U16077 ( .A(n15043), .Z(n15054) );
  XOR U16078 ( .A(n15055), .B(n15056), .Z(n15043) );
  AND U16079 ( .A(n15057), .B(n15058), .Z(n15056) );
  XNOR U16080 ( .A(n15055), .B(n7530), .Z(n15058) );
  XNOR U16081 ( .A(n15051), .B(n15053), .Z(n7530) );
  NAND U16082 ( .A(n15059), .B(e_input[795]), .Z(n15053) );
  NAND U16083 ( .A(n12323), .B(e_input[795]), .Z(n15059) );
  XNOR U16084 ( .A(n15049), .B(n15060), .Z(n15051) );
  XOR U16085 ( .A(n15061), .B(n15062), .Z(n15049) );
  AND U16086 ( .A(n15063), .B(n15064), .Z(n15062) );
  XNOR U16087 ( .A(n15065), .B(n15061), .Z(n15064) );
  XOR U16088 ( .A(n15066), .B(e_input[795]), .Z(n15057) );
  IV U16089 ( .A(n15055), .Z(n15066) );
  XOR U16090 ( .A(n15067), .B(n15068), .Z(n15055) );
  AND U16091 ( .A(n15069), .B(n15070), .Z(n15068) );
  XNOR U16092 ( .A(n15067), .B(n7536), .Z(n15070) );
  XNOR U16093 ( .A(n15063), .B(n15065), .Z(n7536) );
  NAND U16094 ( .A(n15071), .B(e_input[794]), .Z(n15065) );
  NAND U16095 ( .A(n12323), .B(e_input[794]), .Z(n15071) );
  XNOR U16096 ( .A(n15061), .B(n15072), .Z(n15063) );
  XOR U16097 ( .A(n15073), .B(n15074), .Z(n15061) );
  AND U16098 ( .A(n15075), .B(n15076), .Z(n15074) );
  XNOR U16099 ( .A(n15077), .B(n15073), .Z(n15076) );
  XOR U16100 ( .A(n15078), .B(e_input[794]), .Z(n15069) );
  IV U16101 ( .A(n15067), .Z(n15078) );
  XOR U16102 ( .A(n15079), .B(n15080), .Z(n15067) );
  AND U16103 ( .A(n15081), .B(n15082), .Z(n15080) );
  XNOR U16104 ( .A(n15079), .B(n7542), .Z(n15082) );
  XNOR U16105 ( .A(n15075), .B(n15077), .Z(n7542) );
  NAND U16106 ( .A(n15083), .B(e_input[793]), .Z(n15077) );
  NAND U16107 ( .A(n12323), .B(e_input[793]), .Z(n15083) );
  XNOR U16108 ( .A(n15073), .B(n15084), .Z(n15075) );
  XOR U16109 ( .A(n15085), .B(n15086), .Z(n15073) );
  AND U16110 ( .A(n15087), .B(n15088), .Z(n15086) );
  XNOR U16111 ( .A(n15089), .B(n15085), .Z(n15088) );
  XOR U16112 ( .A(n15090), .B(e_input[793]), .Z(n15081) );
  IV U16113 ( .A(n15079), .Z(n15090) );
  XOR U16114 ( .A(n15091), .B(n15092), .Z(n15079) );
  AND U16115 ( .A(n15093), .B(n15094), .Z(n15092) );
  XNOR U16116 ( .A(n15091), .B(n7548), .Z(n15094) );
  XNOR U16117 ( .A(n15087), .B(n15089), .Z(n7548) );
  NAND U16118 ( .A(n15095), .B(e_input[792]), .Z(n15089) );
  NAND U16119 ( .A(n12323), .B(e_input[792]), .Z(n15095) );
  XNOR U16120 ( .A(n15085), .B(n15096), .Z(n15087) );
  XOR U16121 ( .A(n15097), .B(n15098), .Z(n15085) );
  AND U16122 ( .A(n15099), .B(n15100), .Z(n15098) );
  XNOR U16123 ( .A(n15101), .B(n15097), .Z(n15100) );
  XOR U16124 ( .A(n15102), .B(e_input[792]), .Z(n15093) );
  IV U16125 ( .A(n15091), .Z(n15102) );
  XOR U16126 ( .A(n15103), .B(n15104), .Z(n15091) );
  AND U16127 ( .A(n15105), .B(n15106), .Z(n15104) );
  XNOR U16128 ( .A(n15103), .B(n7554), .Z(n15106) );
  XNOR U16129 ( .A(n15099), .B(n15101), .Z(n7554) );
  NAND U16130 ( .A(n15107), .B(e_input[791]), .Z(n15101) );
  NAND U16131 ( .A(n12323), .B(e_input[791]), .Z(n15107) );
  XNOR U16132 ( .A(n15097), .B(n15108), .Z(n15099) );
  XOR U16133 ( .A(n15109), .B(n15110), .Z(n15097) );
  AND U16134 ( .A(n15111), .B(n15112), .Z(n15110) );
  XNOR U16135 ( .A(n15113), .B(n15109), .Z(n15112) );
  XOR U16136 ( .A(n15114), .B(e_input[791]), .Z(n15105) );
  IV U16137 ( .A(n15103), .Z(n15114) );
  XOR U16138 ( .A(n15115), .B(n15116), .Z(n15103) );
  AND U16139 ( .A(n15117), .B(n15118), .Z(n15116) );
  XNOR U16140 ( .A(n15115), .B(n7560), .Z(n15118) );
  XNOR U16141 ( .A(n15111), .B(n15113), .Z(n7560) );
  NAND U16142 ( .A(n15119), .B(e_input[790]), .Z(n15113) );
  NAND U16143 ( .A(n12323), .B(e_input[790]), .Z(n15119) );
  XNOR U16144 ( .A(n15109), .B(n15120), .Z(n15111) );
  XOR U16145 ( .A(n15121), .B(n15122), .Z(n15109) );
  AND U16146 ( .A(n15123), .B(n15124), .Z(n15122) );
  XNOR U16147 ( .A(n15125), .B(n15121), .Z(n15124) );
  XOR U16148 ( .A(n15126), .B(e_input[790]), .Z(n15117) );
  IV U16149 ( .A(n15115), .Z(n15126) );
  XOR U16150 ( .A(n15127), .B(n15128), .Z(n15115) );
  AND U16151 ( .A(n15129), .B(n15130), .Z(n15128) );
  XNOR U16152 ( .A(n15127), .B(n7566), .Z(n15130) );
  XNOR U16153 ( .A(n15123), .B(n15125), .Z(n7566) );
  NAND U16154 ( .A(n15131), .B(e_input[789]), .Z(n15125) );
  NAND U16155 ( .A(n12323), .B(e_input[789]), .Z(n15131) );
  XNOR U16156 ( .A(n15121), .B(n15132), .Z(n15123) );
  XOR U16157 ( .A(n15133), .B(n15134), .Z(n15121) );
  AND U16158 ( .A(n15135), .B(n15136), .Z(n15134) );
  XNOR U16159 ( .A(n15137), .B(n15133), .Z(n15136) );
  XOR U16160 ( .A(n15138), .B(e_input[789]), .Z(n15129) );
  IV U16161 ( .A(n15127), .Z(n15138) );
  XOR U16162 ( .A(n15139), .B(n15140), .Z(n15127) );
  AND U16163 ( .A(n15141), .B(n15142), .Z(n15140) );
  XNOR U16164 ( .A(n15139), .B(n7572), .Z(n15142) );
  XNOR U16165 ( .A(n15135), .B(n15137), .Z(n7572) );
  NAND U16166 ( .A(n15143), .B(e_input[788]), .Z(n15137) );
  NAND U16167 ( .A(n12323), .B(e_input[788]), .Z(n15143) );
  XNOR U16168 ( .A(n15133), .B(n15144), .Z(n15135) );
  XOR U16169 ( .A(n15145), .B(n15146), .Z(n15133) );
  AND U16170 ( .A(n15147), .B(n15148), .Z(n15146) );
  XNOR U16171 ( .A(n15149), .B(n15145), .Z(n15148) );
  XOR U16172 ( .A(n15150), .B(e_input[788]), .Z(n15141) );
  IV U16173 ( .A(n15139), .Z(n15150) );
  XOR U16174 ( .A(n15151), .B(n15152), .Z(n15139) );
  AND U16175 ( .A(n15153), .B(n15154), .Z(n15152) );
  XNOR U16176 ( .A(n15151), .B(n7578), .Z(n15154) );
  XNOR U16177 ( .A(n15147), .B(n15149), .Z(n7578) );
  NAND U16178 ( .A(n15155), .B(e_input[787]), .Z(n15149) );
  NAND U16179 ( .A(n12323), .B(e_input[787]), .Z(n15155) );
  XNOR U16180 ( .A(n15145), .B(n15156), .Z(n15147) );
  XOR U16181 ( .A(n15157), .B(n15158), .Z(n15145) );
  AND U16182 ( .A(n15159), .B(n15160), .Z(n15158) );
  XNOR U16183 ( .A(n15161), .B(n15157), .Z(n15160) );
  XOR U16184 ( .A(n15162), .B(e_input[787]), .Z(n15153) );
  IV U16185 ( .A(n15151), .Z(n15162) );
  XOR U16186 ( .A(n15163), .B(n15164), .Z(n15151) );
  AND U16187 ( .A(n15165), .B(n15166), .Z(n15164) );
  XNOR U16188 ( .A(n15163), .B(n7584), .Z(n15166) );
  XNOR U16189 ( .A(n15159), .B(n15161), .Z(n7584) );
  NAND U16190 ( .A(n15167), .B(e_input[786]), .Z(n15161) );
  NAND U16191 ( .A(n12323), .B(e_input[786]), .Z(n15167) );
  XNOR U16192 ( .A(n15157), .B(n15168), .Z(n15159) );
  XOR U16193 ( .A(n15169), .B(n15170), .Z(n15157) );
  AND U16194 ( .A(n15171), .B(n15172), .Z(n15170) );
  XNOR U16195 ( .A(n15173), .B(n15169), .Z(n15172) );
  XOR U16196 ( .A(n15174), .B(e_input[786]), .Z(n15165) );
  IV U16197 ( .A(n15163), .Z(n15174) );
  XOR U16198 ( .A(n15175), .B(n15176), .Z(n15163) );
  AND U16199 ( .A(n15177), .B(n15178), .Z(n15176) );
  XNOR U16200 ( .A(n15175), .B(n7590), .Z(n15178) );
  XNOR U16201 ( .A(n15171), .B(n15173), .Z(n7590) );
  NAND U16202 ( .A(n15179), .B(e_input[785]), .Z(n15173) );
  NAND U16203 ( .A(n12323), .B(e_input[785]), .Z(n15179) );
  XNOR U16204 ( .A(n15169), .B(n15180), .Z(n15171) );
  XOR U16205 ( .A(n15181), .B(n15182), .Z(n15169) );
  AND U16206 ( .A(n15183), .B(n15184), .Z(n15182) );
  XNOR U16207 ( .A(n15185), .B(n15181), .Z(n15184) );
  XOR U16208 ( .A(n15186), .B(e_input[785]), .Z(n15177) );
  IV U16209 ( .A(n15175), .Z(n15186) );
  XOR U16210 ( .A(n15187), .B(n15188), .Z(n15175) );
  AND U16211 ( .A(n15189), .B(n15190), .Z(n15188) );
  XNOR U16212 ( .A(n15187), .B(n7596), .Z(n15190) );
  XNOR U16213 ( .A(n15183), .B(n15185), .Z(n7596) );
  NAND U16214 ( .A(n15191), .B(e_input[784]), .Z(n15185) );
  NAND U16215 ( .A(n12323), .B(e_input[784]), .Z(n15191) );
  XNOR U16216 ( .A(n15181), .B(n15192), .Z(n15183) );
  XOR U16217 ( .A(n15193), .B(n15194), .Z(n15181) );
  AND U16218 ( .A(n15195), .B(n15196), .Z(n15194) );
  XNOR U16219 ( .A(n15197), .B(n15193), .Z(n15196) );
  XOR U16220 ( .A(n15198), .B(e_input[784]), .Z(n15189) );
  IV U16221 ( .A(n15187), .Z(n15198) );
  XOR U16222 ( .A(n15199), .B(n15200), .Z(n15187) );
  AND U16223 ( .A(n15201), .B(n15202), .Z(n15200) );
  XNOR U16224 ( .A(n15199), .B(n7602), .Z(n15202) );
  XNOR U16225 ( .A(n15195), .B(n15197), .Z(n7602) );
  NAND U16226 ( .A(n15203), .B(e_input[783]), .Z(n15197) );
  NAND U16227 ( .A(n12323), .B(e_input[783]), .Z(n15203) );
  XNOR U16228 ( .A(n15193), .B(n15204), .Z(n15195) );
  XOR U16229 ( .A(n15205), .B(n15206), .Z(n15193) );
  AND U16230 ( .A(n15207), .B(n15208), .Z(n15206) );
  XNOR U16231 ( .A(n15209), .B(n15205), .Z(n15208) );
  XOR U16232 ( .A(n15210), .B(e_input[783]), .Z(n15201) );
  IV U16233 ( .A(n15199), .Z(n15210) );
  XOR U16234 ( .A(n15211), .B(n15212), .Z(n15199) );
  AND U16235 ( .A(n15213), .B(n15214), .Z(n15212) );
  XNOR U16236 ( .A(n15211), .B(n7608), .Z(n15214) );
  XNOR U16237 ( .A(n15207), .B(n15209), .Z(n7608) );
  NAND U16238 ( .A(n15215), .B(e_input[782]), .Z(n15209) );
  NAND U16239 ( .A(n12323), .B(e_input[782]), .Z(n15215) );
  XNOR U16240 ( .A(n15205), .B(n15216), .Z(n15207) );
  XOR U16241 ( .A(n15217), .B(n15218), .Z(n15205) );
  AND U16242 ( .A(n15219), .B(n15220), .Z(n15218) );
  XNOR U16243 ( .A(n15221), .B(n15217), .Z(n15220) );
  XOR U16244 ( .A(n15222), .B(e_input[782]), .Z(n15213) );
  IV U16245 ( .A(n15211), .Z(n15222) );
  XOR U16246 ( .A(n15223), .B(n15224), .Z(n15211) );
  AND U16247 ( .A(n15225), .B(n15226), .Z(n15224) );
  XNOR U16248 ( .A(n15223), .B(n7614), .Z(n15226) );
  XNOR U16249 ( .A(n15219), .B(n15221), .Z(n7614) );
  NAND U16250 ( .A(n15227), .B(e_input[781]), .Z(n15221) );
  NAND U16251 ( .A(n12323), .B(e_input[781]), .Z(n15227) );
  XNOR U16252 ( .A(n15217), .B(n15228), .Z(n15219) );
  XOR U16253 ( .A(n15229), .B(n15230), .Z(n15217) );
  AND U16254 ( .A(n15231), .B(n15232), .Z(n15230) );
  XNOR U16255 ( .A(n15233), .B(n15229), .Z(n15232) );
  XOR U16256 ( .A(n15234), .B(e_input[781]), .Z(n15225) );
  IV U16257 ( .A(n15223), .Z(n15234) );
  XOR U16258 ( .A(n15235), .B(n15236), .Z(n15223) );
  AND U16259 ( .A(n15237), .B(n15238), .Z(n15236) );
  XNOR U16260 ( .A(n15235), .B(n7620), .Z(n15238) );
  XNOR U16261 ( .A(n15231), .B(n15233), .Z(n7620) );
  NAND U16262 ( .A(n15239), .B(e_input[780]), .Z(n15233) );
  NAND U16263 ( .A(n12323), .B(e_input[780]), .Z(n15239) );
  XNOR U16264 ( .A(n15229), .B(n15240), .Z(n15231) );
  XOR U16265 ( .A(n15241), .B(n15242), .Z(n15229) );
  AND U16266 ( .A(n15243), .B(n15244), .Z(n15242) );
  XNOR U16267 ( .A(n15245), .B(n15241), .Z(n15244) );
  XOR U16268 ( .A(n15246), .B(e_input[780]), .Z(n15237) );
  IV U16269 ( .A(n15235), .Z(n15246) );
  XOR U16270 ( .A(n15247), .B(n15248), .Z(n15235) );
  AND U16271 ( .A(n15249), .B(n15250), .Z(n15248) );
  XNOR U16272 ( .A(n15247), .B(n7626), .Z(n15250) );
  XNOR U16273 ( .A(n15243), .B(n15245), .Z(n7626) );
  NAND U16274 ( .A(n15251), .B(e_input[779]), .Z(n15245) );
  NAND U16275 ( .A(n12323), .B(e_input[779]), .Z(n15251) );
  XNOR U16276 ( .A(n15241), .B(n15252), .Z(n15243) );
  XOR U16277 ( .A(n15253), .B(n15254), .Z(n15241) );
  AND U16278 ( .A(n15255), .B(n15256), .Z(n15254) );
  XNOR U16279 ( .A(n15257), .B(n15253), .Z(n15256) );
  XOR U16280 ( .A(n15258), .B(e_input[779]), .Z(n15249) );
  IV U16281 ( .A(n15247), .Z(n15258) );
  XOR U16282 ( .A(n15259), .B(n15260), .Z(n15247) );
  AND U16283 ( .A(n15261), .B(n15262), .Z(n15260) );
  XNOR U16284 ( .A(n15259), .B(n7632), .Z(n15262) );
  XNOR U16285 ( .A(n15255), .B(n15257), .Z(n7632) );
  NAND U16286 ( .A(n15263), .B(e_input[778]), .Z(n15257) );
  NAND U16287 ( .A(n12323), .B(e_input[778]), .Z(n15263) );
  XNOR U16288 ( .A(n15253), .B(n15264), .Z(n15255) );
  XOR U16289 ( .A(n15265), .B(n15266), .Z(n15253) );
  AND U16290 ( .A(n15267), .B(n15268), .Z(n15266) );
  XNOR U16291 ( .A(n15269), .B(n15265), .Z(n15268) );
  XOR U16292 ( .A(n15270), .B(e_input[778]), .Z(n15261) );
  IV U16293 ( .A(n15259), .Z(n15270) );
  XOR U16294 ( .A(n15271), .B(n15272), .Z(n15259) );
  AND U16295 ( .A(n15273), .B(n15274), .Z(n15272) );
  XNOR U16296 ( .A(n15271), .B(n7638), .Z(n15274) );
  XNOR U16297 ( .A(n15267), .B(n15269), .Z(n7638) );
  NAND U16298 ( .A(n15275), .B(e_input[777]), .Z(n15269) );
  NAND U16299 ( .A(n12323), .B(e_input[777]), .Z(n15275) );
  XNOR U16300 ( .A(n15265), .B(n15276), .Z(n15267) );
  XOR U16301 ( .A(n15277), .B(n15278), .Z(n15265) );
  AND U16302 ( .A(n15279), .B(n15280), .Z(n15278) );
  XNOR U16303 ( .A(n15281), .B(n15277), .Z(n15280) );
  XOR U16304 ( .A(n15282), .B(e_input[777]), .Z(n15273) );
  IV U16305 ( .A(n15271), .Z(n15282) );
  XOR U16306 ( .A(n15283), .B(n15284), .Z(n15271) );
  AND U16307 ( .A(n15285), .B(n15286), .Z(n15284) );
  XNOR U16308 ( .A(n15283), .B(n7644), .Z(n15286) );
  XNOR U16309 ( .A(n15279), .B(n15281), .Z(n7644) );
  NAND U16310 ( .A(n15287), .B(e_input[776]), .Z(n15281) );
  NAND U16311 ( .A(n12323), .B(e_input[776]), .Z(n15287) );
  XNOR U16312 ( .A(n15277), .B(n15288), .Z(n15279) );
  XOR U16313 ( .A(n15289), .B(n15290), .Z(n15277) );
  AND U16314 ( .A(n15291), .B(n15292), .Z(n15290) );
  XNOR U16315 ( .A(n15293), .B(n15289), .Z(n15292) );
  XOR U16316 ( .A(n15294), .B(e_input[776]), .Z(n15285) );
  IV U16317 ( .A(n15283), .Z(n15294) );
  XOR U16318 ( .A(n15295), .B(n15296), .Z(n15283) );
  AND U16319 ( .A(n15297), .B(n15298), .Z(n15296) );
  XNOR U16320 ( .A(n15295), .B(n7650), .Z(n15298) );
  XNOR U16321 ( .A(n15291), .B(n15293), .Z(n7650) );
  NAND U16322 ( .A(n15299), .B(e_input[775]), .Z(n15293) );
  NAND U16323 ( .A(n12323), .B(e_input[775]), .Z(n15299) );
  XNOR U16324 ( .A(n15289), .B(n15300), .Z(n15291) );
  XOR U16325 ( .A(n15301), .B(n15302), .Z(n15289) );
  AND U16326 ( .A(n15303), .B(n15304), .Z(n15302) );
  XNOR U16327 ( .A(n15305), .B(n15301), .Z(n15304) );
  XOR U16328 ( .A(n15306), .B(e_input[775]), .Z(n15297) );
  IV U16329 ( .A(n15295), .Z(n15306) );
  XOR U16330 ( .A(n15307), .B(n15308), .Z(n15295) );
  AND U16331 ( .A(n15309), .B(n15310), .Z(n15308) );
  XNOR U16332 ( .A(n15307), .B(n7656), .Z(n15310) );
  XNOR U16333 ( .A(n15303), .B(n15305), .Z(n7656) );
  NAND U16334 ( .A(n15311), .B(e_input[774]), .Z(n15305) );
  NAND U16335 ( .A(n12323), .B(e_input[774]), .Z(n15311) );
  XNOR U16336 ( .A(n15301), .B(n15312), .Z(n15303) );
  XOR U16337 ( .A(n15313), .B(n15314), .Z(n15301) );
  AND U16338 ( .A(n15315), .B(n15316), .Z(n15314) );
  XNOR U16339 ( .A(n15317), .B(n15313), .Z(n15316) );
  XOR U16340 ( .A(n15318), .B(e_input[774]), .Z(n15309) );
  IV U16341 ( .A(n15307), .Z(n15318) );
  XOR U16342 ( .A(n15319), .B(n15320), .Z(n15307) );
  AND U16343 ( .A(n15321), .B(n15322), .Z(n15320) );
  XNOR U16344 ( .A(n15319), .B(n7662), .Z(n15322) );
  XNOR U16345 ( .A(n15315), .B(n15317), .Z(n7662) );
  NAND U16346 ( .A(n15323), .B(e_input[773]), .Z(n15317) );
  NAND U16347 ( .A(n12323), .B(e_input[773]), .Z(n15323) );
  XNOR U16348 ( .A(n15313), .B(n15324), .Z(n15315) );
  XOR U16349 ( .A(n15325), .B(n15326), .Z(n15313) );
  AND U16350 ( .A(n15327), .B(n15328), .Z(n15326) );
  XNOR U16351 ( .A(n15329), .B(n15325), .Z(n15328) );
  XOR U16352 ( .A(n15330), .B(e_input[773]), .Z(n15321) );
  IV U16353 ( .A(n15319), .Z(n15330) );
  XOR U16354 ( .A(n15331), .B(n15332), .Z(n15319) );
  AND U16355 ( .A(n15333), .B(n15334), .Z(n15332) );
  XNOR U16356 ( .A(n15331), .B(n7668), .Z(n15334) );
  XNOR U16357 ( .A(n15327), .B(n15329), .Z(n7668) );
  NAND U16358 ( .A(n15335), .B(e_input[772]), .Z(n15329) );
  NAND U16359 ( .A(n12323), .B(e_input[772]), .Z(n15335) );
  XNOR U16360 ( .A(n15325), .B(n15336), .Z(n15327) );
  XOR U16361 ( .A(n15337), .B(n15338), .Z(n15325) );
  AND U16362 ( .A(n15339), .B(n15340), .Z(n15338) );
  XNOR U16363 ( .A(n15341), .B(n15337), .Z(n15340) );
  XOR U16364 ( .A(n15342), .B(e_input[772]), .Z(n15333) );
  IV U16365 ( .A(n15331), .Z(n15342) );
  XOR U16366 ( .A(n15343), .B(n15344), .Z(n15331) );
  AND U16367 ( .A(n15345), .B(n15346), .Z(n15344) );
  XNOR U16368 ( .A(n15343), .B(n7674), .Z(n15346) );
  XNOR U16369 ( .A(n15339), .B(n15341), .Z(n7674) );
  NAND U16370 ( .A(n15347), .B(e_input[771]), .Z(n15341) );
  NAND U16371 ( .A(n12323), .B(e_input[771]), .Z(n15347) );
  XNOR U16372 ( .A(n15337), .B(n15348), .Z(n15339) );
  XOR U16373 ( .A(n15349), .B(n15350), .Z(n15337) );
  AND U16374 ( .A(n15351), .B(n15352), .Z(n15350) );
  XNOR U16375 ( .A(n15353), .B(n15349), .Z(n15352) );
  XOR U16376 ( .A(n15354), .B(e_input[771]), .Z(n15345) );
  IV U16377 ( .A(n15343), .Z(n15354) );
  XOR U16378 ( .A(n15355), .B(n15356), .Z(n15343) );
  AND U16379 ( .A(n15357), .B(n15358), .Z(n15356) );
  XNOR U16380 ( .A(n15355), .B(n7680), .Z(n15358) );
  XNOR U16381 ( .A(n15351), .B(n15353), .Z(n7680) );
  NAND U16382 ( .A(n15359), .B(e_input[770]), .Z(n15353) );
  NAND U16383 ( .A(n12323), .B(e_input[770]), .Z(n15359) );
  XNOR U16384 ( .A(n15349), .B(n15360), .Z(n15351) );
  XOR U16385 ( .A(n15361), .B(n15362), .Z(n15349) );
  AND U16386 ( .A(n15363), .B(n15364), .Z(n15362) );
  XNOR U16387 ( .A(n15365), .B(n15361), .Z(n15364) );
  XOR U16388 ( .A(n15366), .B(e_input[770]), .Z(n15357) );
  IV U16389 ( .A(n15355), .Z(n15366) );
  XOR U16390 ( .A(n15367), .B(n15368), .Z(n15355) );
  AND U16391 ( .A(n15369), .B(n15370), .Z(n15368) );
  XNOR U16392 ( .A(n15367), .B(n7686), .Z(n15370) );
  XNOR U16393 ( .A(n15363), .B(n15365), .Z(n7686) );
  NAND U16394 ( .A(n15371), .B(e_input[769]), .Z(n15365) );
  NAND U16395 ( .A(n12323), .B(e_input[769]), .Z(n15371) );
  XNOR U16396 ( .A(n15361), .B(n15372), .Z(n15363) );
  XOR U16397 ( .A(n15373), .B(n15374), .Z(n15361) );
  AND U16398 ( .A(n15375), .B(n15376), .Z(n15374) );
  XNOR U16399 ( .A(n15377), .B(n15373), .Z(n15376) );
  XOR U16400 ( .A(n15378), .B(e_input[769]), .Z(n15369) );
  IV U16401 ( .A(n15367), .Z(n15378) );
  XOR U16402 ( .A(n15379), .B(n15380), .Z(n15367) );
  AND U16403 ( .A(n15381), .B(n15382), .Z(n15380) );
  XNOR U16404 ( .A(n15379), .B(n7692), .Z(n15382) );
  XNOR U16405 ( .A(n15375), .B(n15377), .Z(n7692) );
  NAND U16406 ( .A(n15383), .B(e_input[768]), .Z(n15377) );
  NAND U16407 ( .A(n12323), .B(e_input[768]), .Z(n15383) );
  XNOR U16408 ( .A(n15373), .B(n15384), .Z(n15375) );
  XOR U16409 ( .A(n15385), .B(n15386), .Z(n15373) );
  AND U16410 ( .A(n15387), .B(n15388), .Z(n15386) );
  XNOR U16411 ( .A(n15389), .B(n15385), .Z(n15388) );
  XOR U16412 ( .A(n15390), .B(e_input[768]), .Z(n15381) );
  IV U16413 ( .A(n15379), .Z(n15390) );
  XOR U16414 ( .A(n15391), .B(n15392), .Z(n15379) );
  AND U16415 ( .A(n15393), .B(n15394), .Z(n15392) );
  XNOR U16416 ( .A(n15391), .B(n7698), .Z(n15394) );
  XNOR U16417 ( .A(n15387), .B(n15389), .Z(n7698) );
  NAND U16418 ( .A(n15395), .B(e_input[767]), .Z(n15389) );
  NAND U16419 ( .A(n12323), .B(e_input[767]), .Z(n15395) );
  XNOR U16420 ( .A(n15385), .B(n15396), .Z(n15387) );
  XOR U16421 ( .A(n15397), .B(n15398), .Z(n15385) );
  AND U16422 ( .A(n15399), .B(n15400), .Z(n15398) );
  XNOR U16423 ( .A(n15401), .B(n15397), .Z(n15400) );
  XOR U16424 ( .A(n15402), .B(e_input[767]), .Z(n15393) );
  IV U16425 ( .A(n15391), .Z(n15402) );
  XOR U16426 ( .A(n15403), .B(n15404), .Z(n15391) );
  AND U16427 ( .A(n15405), .B(n15406), .Z(n15404) );
  XNOR U16428 ( .A(n15403), .B(n7704), .Z(n15406) );
  XNOR U16429 ( .A(n15399), .B(n15401), .Z(n7704) );
  NAND U16430 ( .A(n15407), .B(e_input[766]), .Z(n15401) );
  NAND U16431 ( .A(n12323), .B(e_input[766]), .Z(n15407) );
  XNOR U16432 ( .A(n15397), .B(n15408), .Z(n15399) );
  XOR U16433 ( .A(n15409), .B(n15410), .Z(n15397) );
  AND U16434 ( .A(n15411), .B(n15412), .Z(n15410) );
  XNOR U16435 ( .A(n15413), .B(n15409), .Z(n15412) );
  XOR U16436 ( .A(n15414), .B(e_input[766]), .Z(n15405) );
  IV U16437 ( .A(n15403), .Z(n15414) );
  XOR U16438 ( .A(n15415), .B(n15416), .Z(n15403) );
  AND U16439 ( .A(n15417), .B(n15418), .Z(n15416) );
  XNOR U16440 ( .A(n15415), .B(n7710), .Z(n15418) );
  XNOR U16441 ( .A(n15411), .B(n15413), .Z(n7710) );
  NAND U16442 ( .A(n15419), .B(e_input[765]), .Z(n15413) );
  NAND U16443 ( .A(n12323), .B(e_input[765]), .Z(n15419) );
  XNOR U16444 ( .A(n15409), .B(n15420), .Z(n15411) );
  XOR U16445 ( .A(n15421), .B(n15422), .Z(n15409) );
  AND U16446 ( .A(n15423), .B(n15424), .Z(n15422) );
  XNOR U16447 ( .A(n15425), .B(n15421), .Z(n15424) );
  XOR U16448 ( .A(n15426), .B(e_input[765]), .Z(n15417) );
  IV U16449 ( .A(n15415), .Z(n15426) );
  XOR U16450 ( .A(n15427), .B(n15428), .Z(n15415) );
  AND U16451 ( .A(n15429), .B(n15430), .Z(n15428) );
  XNOR U16452 ( .A(n15427), .B(n7716), .Z(n15430) );
  XNOR U16453 ( .A(n15423), .B(n15425), .Z(n7716) );
  NAND U16454 ( .A(n15431), .B(e_input[764]), .Z(n15425) );
  NAND U16455 ( .A(n12323), .B(e_input[764]), .Z(n15431) );
  XNOR U16456 ( .A(n15421), .B(n15432), .Z(n15423) );
  XOR U16457 ( .A(n15433), .B(n15434), .Z(n15421) );
  AND U16458 ( .A(n15435), .B(n15436), .Z(n15434) );
  XNOR U16459 ( .A(n15437), .B(n15433), .Z(n15436) );
  XOR U16460 ( .A(n15438), .B(e_input[764]), .Z(n15429) );
  IV U16461 ( .A(n15427), .Z(n15438) );
  XOR U16462 ( .A(n15439), .B(n15440), .Z(n15427) );
  AND U16463 ( .A(n15441), .B(n15442), .Z(n15440) );
  XNOR U16464 ( .A(n15439), .B(n7722), .Z(n15442) );
  XNOR U16465 ( .A(n15435), .B(n15437), .Z(n7722) );
  NAND U16466 ( .A(n15443), .B(e_input[763]), .Z(n15437) );
  NAND U16467 ( .A(n12323), .B(e_input[763]), .Z(n15443) );
  XNOR U16468 ( .A(n15433), .B(n15444), .Z(n15435) );
  XOR U16469 ( .A(n15445), .B(n15446), .Z(n15433) );
  AND U16470 ( .A(n15447), .B(n15448), .Z(n15446) );
  XNOR U16471 ( .A(n15449), .B(n15445), .Z(n15448) );
  XOR U16472 ( .A(n15450), .B(e_input[763]), .Z(n15441) );
  IV U16473 ( .A(n15439), .Z(n15450) );
  XOR U16474 ( .A(n15451), .B(n15452), .Z(n15439) );
  AND U16475 ( .A(n15453), .B(n15454), .Z(n15452) );
  XNOR U16476 ( .A(n15451), .B(n7728), .Z(n15454) );
  XNOR U16477 ( .A(n15447), .B(n15449), .Z(n7728) );
  NAND U16478 ( .A(n15455), .B(e_input[762]), .Z(n15449) );
  NAND U16479 ( .A(n12323), .B(e_input[762]), .Z(n15455) );
  XNOR U16480 ( .A(n15445), .B(n15456), .Z(n15447) );
  XOR U16481 ( .A(n15457), .B(n15458), .Z(n15445) );
  AND U16482 ( .A(n15459), .B(n15460), .Z(n15458) );
  XNOR U16483 ( .A(n15461), .B(n15457), .Z(n15460) );
  XOR U16484 ( .A(n15462), .B(e_input[762]), .Z(n15453) );
  IV U16485 ( .A(n15451), .Z(n15462) );
  XOR U16486 ( .A(n15463), .B(n15464), .Z(n15451) );
  AND U16487 ( .A(n15465), .B(n15466), .Z(n15464) );
  XNOR U16488 ( .A(n15463), .B(n7734), .Z(n15466) );
  XNOR U16489 ( .A(n15459), .B(n15461), .Z(n7734) );
  NAND U16490 ( .A(n15467), .B(e_input[761]), .Z(n15461) );
  NAND U16491 ( .A(n12323), .B(e_input[761]), .Z(n15467) );
  XNOR U16492 ( .A(n15457), .B(n15468), .Z(n15459) );
  XOR U16493 ( .A(n15469), .B(n15470), .Z(n15457) );
  AND U16494 ( .A(n15471), .B(n15472), .Z(n15470) );
  XNOR U16495 ( .A(n15473), .B(n15469), .Z(n15472) );
  XOR U16496 ( .A(n15474), .B(e_input[761]), .Z(n15465) );
  IV U16497 ( .A(n15463), .Z(n15474) );
  XOR U16498 ( .A(n15475), .B(n15476), .Z(n15463) );
  AND U16499 ( .A(n15477), .B(n15478), .Z(n15476) );
  XNOR U16500 ( .A(n15475), .B(n7740), .Z(n15478) );
  XNOR U16501 ( .A(n15471), .B(n15473), .Z(n7740) );
  NAND U16502 ( .A(n15479), .B(e_input[760]), .Z(n15473) );
  NAND U16503 ( .A(n12323), .B(e_input[760]), .Z(n15479) );
  XNOR U16504 ( .A(n15469), .B(n15480), .Z(n15471) );
  XOR U16505 ( .A(n15481), .B(n15482), .Z(n15469) );
  AND U16506 ( .A(n15483), .B(n15484), .Z(n15482) );
  XNOR U16507 ( .A(n15485), .B(n15481), .Z(n15484) );
  XOR U16508 ( .A(n15486), .B(e_input[760]), .Z(n15477) );
  IV U16509 ( .A(n15475), .Z(n15486) );
  XOR U16510 ( .A(n15487), .B(n15488), .Z(n15475) );
  AND U16511 ( .A(n15489), .B(n15490), .Z(n15488) );
  XNOR U16512 ( .A(n15487), .B(n7746), .Z(n15490) );
  XNOR U16513 ( .A(n15483), .B(n15485), .Z(n7746) );
  NAND U16514 ( .A(n15491), .B(e_input[759]), .Z(n15485) );
  NAND U16515 ( .A(n12323), .B(e_input[759]), .Z(n15491) );
  XNOR U16516 ( .A(n15481), .B(n15492), .Z(n15483) );
  XOR U16517 ( .A(n15493), .B(n15494), .Z(n15481) );
  AND U16518 ( .A(n15495), .B(n15496), .Z(n15494) );
  XNOR U16519 ( .A(n15497), .B(n15493), .Z(n15496) );
  XOR U16520 ( .A(n15498), .B(e_input[759]), .Z(n15489) );
  IV U16521 ( .A(n15487), .Z(n15498) );
  XOR U16522 ( .A(n15499), .B(n15500), .Z(n15487) );
  AND U16523 ( .A(n15501), .B(n15502), .Z(n15500) );
  XNOR U16524 ( .A(n15499), .B(n7752), .Z(n15502) );
  XNOR U16525 ( .A(n15495), .B(n15497), .Z(n7752) );
  NAND U16526 ( .A(n15503), .B(e_input[758]), .Z(n15497) );
  NAND U16527 ( .A(n12323), .B(e_input[758]), .Z(n15503) );
  XNOR U16528 ( .A(n15493), .B(n15504), .Z(n15495) );
  XOR U16529 ( .A(n15505), .B(n15506), .Z(n15493) );
  AND U16530 ( .A(n15507), .B(n15508), .Z(n15506) );
  XNOR U16531 ( .A(n15509), .B(n15505), .Z(n15508) );
  XOR U16532 ( .A(n15510), .B(e_input[758]), .Z(n15501) );
  IV U16533 ( .A(n15499), .Z(n15510) );
  XOR U16534 ( .A(n15511), .B(n15512), .Z(n15499) );
  AND U16535 ( .A(n15513), .B(n15514), .Z(n15512) );
  XNOR U16536 ( .A(n15511), .B(n7758), .Z(n15514) );
  XNOR U16537 ( .A(n15507), .B(n15509), .Z(n7758) );
  NAND U16538 ( .A(n15515), .B(e_input[757]), .Z(n15509) );
  NAND U16539 ( .A(n12323), .B(e_input[757]), .Z(n15515) );
  XNOR U16540 ( .A(n15505), .B(n15516), .Z(n15507) );
  XOR U16541 ( .A(n15517), .B(n15518), .Z(n15505) );
  AND U16542 ( .A(n15519), .B(n15520), .Z(n15518) );
  XNOR U16543 ( .A(n15521), .B(n15517), .Z(n15520) );
  XOR U16544 ( .A(n15522), .B(e_input[757]), .Z(n15513) );
  IV U16545 ( .A(n15511), .Z(n15522) );
  XOR U16546 ( .A(n15523), .B(n15524), .Z(n15511) );
  AND U16547 ( .A(n15525), .B(n15526), .Z(n15524) );
  XNOR U16548 ( .A(n15523), .B(n7764), .Z(n15526) );
  XNOR U16549 ( .A(n15519), .B(n15521), .Z(n7764) );
  NAND U16550 ( .A(n15527), .B(e_input[756]), .Z(n15521) );
  NAND U16551 ( .A(n12323), .B(e_input[756]), .Z(n15527) );
  XNOR U16552 ( .A(n15517), .B(n15528), .Z(n15519) );
  XOR U16553 ( .A(n15529), .B(n15530), .Z(n15517) );
  AND U16554 ( .A(n15531), .B(n15532), .Z(n15530) );
  XNOR U16555 ( .A(n15533), .B(n15529), .Z(n15532) );
  XOR U16556 ( .A(n15534), .B(e_input[756]), .Z(n15525) );
  IV U16557 ( .A(n15523), .Z(n15534) );
  XOR U16558 ( .A(n15535), .B(n15536), .Z(n15523) );
  AND U16559 ( .A(n15537), .B(n15538), .Z(n15536) );
  XNOR U16560 ( .A(n15535), .B(n7770), .Z(n15538) );
  XNOR U16561 ( .A(n15531), .B(n15533), .Z(n7770) );
  NAND U16562 ( .A(n15539), .B(e_input[755]), .Z(n15533) );
  NAND U16563 ( .A(n12323), .B(e_input[755]), .Z(n15539) );
  XNOR U16564 ( .A(n15529), .B(n15540), .Z(n15531) );
  XOR U16565 ( .A(n15541), .B(n15542), .Z(n15529) );
  AND U16566 ( .A(n15543), .B(n15544), .Z(n15542) );
  XNOR U16567 ( .A(n15545), .B(n15541), .Z(n15544) );
  XOR U16568 ( .A(n15546), .B(e_input[755]), .Z(n15537) );
  IV U16569 ( .A(n15535), .Z(n15546) );
  XOR U16570 ( .A(n15547), .B(n15548), .Z(n15535) );
  AND U16571 ( .A(n15549), .B(n15550), .Z(n15548) );
  XNOR U16572 ( .A(n15547), .B(n7776), .Z(n15550) );
  XNOR U16573 ( .A(n15543), .B(n15545), .Z(n7776) );
  NAND U16574 ( .A(n15551), .B(e_input[754]), .Z(n15545) );
  NAND U16575 ( .A(n12323), .B(e_input[754]), .Z(n15551) );
  XNOR U16576 ( .A(n15541), .B(n15552), .Z(n15543) );
  XOR U16577 ( .A(n15553), .B(n15554), .Z(n15541) );
  AND U16578 ( .A(n15555), .B(n15556), .Z(n15554) );
  XNOR U16579 ( .A(n15557), .B(n15553), .Z(n15556) );
  XOR U16580 ( .A(n15558), .B(e_input[754]), .Z(n15549) );
  IV U16581 ( .A(n15547), .Z(n15558) );
  XOR U16582 ( .A(n15559), .B(n15560), .Z(n15547) );
  AND U16583 ( .A(n15561), .B(n15562), .Z(n15560) );
  XNOR U16584 ( .A(n15559), .B(n7782), .Z(n15562) );
  XNOR U16585 ( .A(n15555), .B(n15557), .Z(n7782) );
  NAND U16586 ( .A(n15563), .B(e_input[753]), .Z(n15557) );
  NAND U16587 ( .A(n12323), .B(e_input[753]), .Z(n15563) );
  XNOR U16588 ( .A(n15553), .B(n15564), .Z(n15555) );
  XOR U16589 ( .A(n15565), .B(n15566), .Z(n15553) );
  AND U16590 ( .A(n15567), .B(n15568), .Z(n15566) );
  XNOR U16591 ( .A(n15569), .B(n15565), .Z(n15568) );
  XOR U16592 ( .A(n15570), .B(e_input[753]), .Z(n15561) );
  IV U16593 ( .A(n15559), .Z(n15570) );
  XOR U16594 ( .A(n15571), .B(n15572), .Z(n15559) );
  AND U16595 ( .A(n15573), .B(n15574), .Z(n15572) );
  XNOR U16596 ( .A(n15571), .B(n7788), .Z(n15574) );
  XNOR U16597 ( .A(n15567), .B(n15569), .Z(n7788) );
  NAND U16598 ( .A(n15575), .B(e_input[752]), .Z(n15569) );
  NAND U16599 ( .A(n12323), .B(e_input[752]), .Z(n15575) );
  XNOR U16600 ( .A(n15565), .B(n15576), .Z(n15567) );
  XOR U16601 ( .A(n15577), .B(n15578), .Z(n15565) );
  AND U16602 ( .A(n15579), .B(n15580), .Z(n15578) );
  XNOR U16603 ( .A(n15581), .B(n15577), .Z(n15580) );
  XOR U16604 ( .A(n15582), .B(e_input[752]), .Z(n15573) );
  IV U16605 ( .A(n15571), .Z(n15582) );
  XOR U16606 ( .A(n15583), .B(n15584), .Z(n15571) );
  AND U16607 ( .A(n15585), .B(n15586), .Z(n15584) );
  XNOR U16608 ( .A(n15583), .B(n7794), .Z(n15586) );
  XNOR U16609 ( .A(n15579), .B(n15581), .Z(n7794) );
  NAND U16610 ( .A(n15587), .B(e_input[751]), .Z(n15581) );
  NAND U16611 ( .A(n12323), .B(e_input[751]), .Z(n15587) );
  XNOR U16612 ( .A(n15577), .B(n15588), .Z(n15579) );
  XOR U16613 ( .A(n15589), .B(n15590), .Z(n15577) );
  AND U16614 ( .A(n15591), .B(n15592), .Z(n15590) );
  XNOR U16615 ( .A(n15593), .B(n15589), .Z(n15592) );
  XOR U16616 ( .A(n15594), .B(e_input[751]), .Z(n15585) );
  IV U16617 ( .A(n15583), .Z(n15594) );
  XOR U16618 ( .A(n15595), .B(n15596), .Z(n15583) );
  AND U16619 ( .A(n15597), .B(n15598), .Z(n15596) );
  XNOR U16620 ( .A(n15595), .B(n7800), .Z(n15598) );
  XNOR U16621 ( .A(n15591), .B(n15593), .Z(n7800) );
  NAND U16622 ( .A(n15599), .B(e_input[750]), .Z(n15593) );
  NAND U16623 ( .A(n12323), .B(e_input[750]), .Z(n15599) );
  XNOR U16624 ( .A(n15589), .B(n15600), .Z(n15591) );
  XOR U16625 ( .A(n15601), .B(n15602), .Z(n15589) );
  AND U16626 ( .A(n15603), .B(n15604), .Z(n15602) );
  XNOR U16627 ( .A(n15605), .B(n15601), .Z(n15604) );
  XOR U16628 ( .A(n15606), .B(e_input[750]), .Z(n15597) );
  IV U16629 ( .A(n15595), .Z(n15606) );
  XOR U16630 ( .A(n15607), .B(n15608), .Z(n15595) );
  AND U16631 ( .A(n15609), .B(n15610), .Z(n15608) );
  XNOR U16632 ( .A(n15607), .B(n7806), .Z(n15610) );
  XNOR U16633 ( .A(n15603), .B(n15605), .Z(n7806) );
  NAND U16634 ( .A(n15611), .B(e_input[749]), .Z(n15605) );
  NAND U16635 ( .A(n12323), .B(e_input[749]), .Z(n15611) );
  XNOR U16636 ( .A(n15601), .B(n15612), .Z(n15603) );
  XOR U16637 ( .A(n15613), .B(n15614), .Z(n15601) );
  AND U16638 ( .A(n15615), .B(n15616), .Z(n15614) );
  XNOR U16639 ( .A(n15617), .B(n15613), .Z(n15616) );
  XOR U16640 ( .A(n15618), .B(e_input[749]), .Z(n15609) );
  IV U16641 ( .A(n15607), .Z(n15618) );
  XOR U16642 ( .A(n15619), .B(n15620), .Z(n15607) );
  AND U16643 ( .A(n15621), .B(n15622), .Z(n15620) );
  XNOR U16644 ( .A(n15619), .B(n7812), .Z(n15622) );
  XNOR U16645 ( .A(n15615), .B(n15617), .Z(n7812) );
  NAND U16646 ( .A(n15623), .B(e_input[748]), .Z(n15617) );
  NAND U16647 ( .A(n12323), .B(e_input[748]), .Z(n15623) );
  XNOR U16648 ( .A(n15613), .B(n15624), .Z(n15615) );
  XOR U16649 ( .A(n15625), .B(n15626), .Z(n15613) );
  AND U16650 ( .A(n15627), .B(n15628), .Z(n15626) );
  XNOR U16651 ( .A(n15629), .B(n15625), .Z(n15628) );
  XOR U16652 ( .A(n15630), .B(e_input[748]), .Z(n15621) );
  IV U16653 ( .A(n15619), .Z(n15630) );
  XOR U16654 ( .A(n15631), .B(n15632), .Z(n15619) );
  AND U16655 ( .A(n15633), .B(n15634), .Z(n15632) );
  XNOR U16656 ( .A(n15631), .B(n7818), .Z(n15634) );
  XNOR U16657 ( .A(n15627), .B(n15629), .Z(n7818) );
  NAND U16658 ( .A(n15635), .B(e_input[747]), .Z(n15629) );
  NAND U16659 ( .A(n12323), .B(e_input[747]), .Z(n15635) );
  XNOR U16660 ( .A(n15625), .B(n15636), .Z(n15627) );
  XOR U16661 ( .A(n15637), .B(n15638), .Z(n15625) );
  AND U16662 ( .A(n15639), .B(n15640), .Z(n15638) );
  XNOR U16663 ( .A(n15641), .B(n15637), .Z(n15640) );
  XOR U16664 ( .A(n15642), .B(e_input[747]), .Z(n15633) );
  IV U16665 ( .A(n15631), .Z(n15642) );
  XOR U16666 ( .A(n15643), .B(n15644), .Z(n15631) );
  AND U16667 ( .A(n15645), .B(n15646), .Z(n15644) );
  XNOR U16668 ( .A(n15643), .B(n7824), .Z(n15646) );
  XNOR U16669 ( .A(n15639), .B(n15641), .Z(n7824) );
  NAND U16670 ( .A(n15647), .B(e_input[746]), .Z(n15641) );
  NAND U16671 ( .A(n12323), .B(e_input[746]), .Z(n15647) );
  XNOR U16672 ( .A(n15637), .B(n15648), .Z(n15639) );
  XOR U16673 ( .A(n15649), .B(n15650), .Z(n15637) );
  AND U16674 ( .A(n15651), .B(n15652), .Z(n15650) );
  XNOR U16675 ( .A(n15653), .B(n15649), .Z(n15652) );
  XOR U16676 ( .A(n15654), .B(e_input[746]), .Z(n15645) );
  IV U16677 ( .A(n15643), .Z(n15654) );
  XOR U16678 ( .A(n15655), .B(n15656), .Z(n15643) );
  AND U16679 ( .A(n15657), .B(n15658), .Z(n15656) );
  XNOR U16680 ( .A(n15655), .B(n7830), .Z(n15658) );
  XNOR U16681 ( .A(n15651), .B(n15653), .Z(n7830) );
  NAND U16682 ( .A(n15659), .B(e_input[745]), .Z(n15653) );
  NAND U16683 ( .A(n12323), .B(e_input[745]), .Z(n15659) );
  XNOR U16684 ( .A(n15649), .B(n15660), .Z(n15651) );
  XOR U16685 ( .A(n15661), .B(n15662), .Z(n15649) );
  AND U16686 ( .A(n15663), .B(n15664), .Z(n15662) );
  XNOR U16687 ( .A(n15665), .B(n15661), .Z(n15664) );
  XOR U16688 ( .A(n15666), .B(e_input[745]), .Z(n15657) );
  IV U16689 ( .A(n15655), .Z(n15666) );
  XOR U16690 ( .A(n15667), .B(n15668), .Z(n15655) );
  AND U16691 ( .A(n15669), .B(n15670), .Z(n15668) );
  XNOR U16692 ( .A(n15667), .B(n7836), .Z(n15670) );
  XNOR U16693 ( .A(n15663), .B(n15665), .Z(n7836) );
  NAND U16694 ( .A(n15671), .B(e_input[744]), .Z(n15665) );
  NAND U16695 ( .A(n12323), .B(e_input[744]), .Z(n15671) );
  XNOR U16696 ( .A(n15661), .B(n15672), .Z(n15663) );
  XOR U16697 ( .A(n15673), .B(n15674), .Z(n15661) );
  AND U16698 ( .A(n15675), .B(n15676), .Z(n15674) );
  XNOR U16699 ( .A(n15677), .B(n15673), .Z(n15676) );
  XOR U16700 ( .A(n15678), .B(e_input[744]), .Z(n15669) );
  IV U16701 ( .A(n15667), .Z(n15678) );
  XOR U16702 ( .A(n15679), .B(n15680), .Z(n15667) );
  AND U16703 ( .A(n15681), .B(n15682), .Z(n15680) );
  XNOR U16704 ( .A(n15679), .B(n7842), .Z(n15682) );
  XNOR U16705 ( .A(n15675), .B(n15677), .Z(n7842) );
  NAND U16706 ( .A(n15683), .B(e_input[743]), .Z(n15677) );
  NAND U16707 ( .A(n12323), .B(e_input[743]), .Z(n15683) );
  XNOR U16708 ( .A(n15673), .B(n15684), .Z(n15675) );
  XOR U16709 ( .A(n15685), .B(n15686), .Z(n15673) );
  AND U16710 ( .A(n15687), .B(n15688), .Z(n15686) );
  XNOR U16711 ( .A(n15689), .B(n15685), .Z(n15688) );
  XOR U16712 ( .A(n15690), .B(e_input[743]), .Z(n15681) );
  IV U16713 ( .A(n15679), .Z(n15690) );
  XOR U16714 ( .A(n15691), .B(n15692), .Z(n15679) );
  AND U16715 ( .A(n15693), .B(n15694), .Z(n15692) );
  XNOR U16716 ( .A(n15691), .B(n7848), .Z(n15694) );
  XNOR U16717 ( .A(n15687), .B(n15689), .Z(n7848) );
  NAND U16718 ( .A(n15695), .B(e_input[742]), .Z(n15689) );
  NAND U16719 ( .A(n12323), .B(e_input[742]), .Z(n15695) );
  XNOR U16720 ( .A(n15685), .B(n15696), .Z(n15687) );
  XOR U16721 ( .A(n15697), .B(n15698), .Z(n15685) );
  AND U16722 ( .A(n15699), .B(n15700), .Z(n15698) );
  XNOR U16723 ( .A(n15701), .B(n15697), .Z(n15700) );
  XOR U16724 ( .A(n15702), .B(e_input[742]), .Z(n15693) );
  IV U16725 ( .A(n15691), .Z(n15702) );
  XOR U16726 ( .A(n15703), .B(n15704), .Z(n15691) );
  AND U16727 ( .A(n15705), .B(n15706), .Z(n15704) );
  XNOR U16728 ( .A(n15703), .B(n7854), .Z(n15706) );
  XNOR U16729 ( .A(n15699), .B(n15701), .Z(n7854) );
  NAND U16730 ( .A(n15707), .B(e_input[741]), .Z(n15701) );
  NAND U16731 ( .A(n12323), .B(e_input[741]), .Z(n15707) );
  XNOR U16732 ( .A(n15697), .B(n15708), .Z(n15699) );
  XOR U16733 ( .A(n15709), .B(n15710), .Z(n15697) );
  AND U16734 ( .A(n15711), .B(n15712), .Z(n15710) );
  XNOR U16735 ( .A(n15713), .B(n15709), .Z(n15712) );
  XOR U16736 ( .A(n15714), .B(e_input[741]), .Z(n15705) );
  IV U16737 ( .A(n15703), .Z(n15714) );
  XOR U16738 ( .A(n15715), .B(n15716), .Z(n15703) );
  AND U16739 ( .A(n15717), .B(n15718), .Z(n15716) );
  XNOR U16740 ( .A(n15715), .B(n7860), .Z(n15718) );
  XNOR U16741 ( .A(n15711), .B(n15713), .Z(n7860) );
  NAND U16742 ( .A(n15719), .B(e_input[740]), .Z(n15713) );
  NAND U16743 ( .A(n12323), .B(e_input[740]), .Z(n15719) );
  XNOR U16744 ( .A(n15709), .B(n15720), .Z(n15711) );
  XOR U16745 ( .A(n15721), .B(n15722), .Z(n15709) );
  AND U16746 ( .A(n15723), .B(n15724), .Z(n15722) );
  XNOR U16747 ( .A(n15725), .B(n15721), .Z(n15724) );
  XOR U16748 ( .A(n15726), .B(e_input[740]), .Z(n15717) );
  IV U16749 ( .A(n15715), .Z(n15726) );
  XOR U16750 ( .A(n15727), .B(n15728), .Z(n15715) );
  AND U16751 ( .A(n15729), .B(n15730), .Z(n15728) );
  XNOR U16752 ( .A(n15727), .B(n7866), .Z(n15730) );
  XNOR U16753 ( .A(n15723), .B(n15725), .Z(n7866) );
  NAND U16754 ( .A(n15731), .B(e_input[739]), .Z(n15725) );
  NAND U16755 ( .A(n12323), .B(e_input[739]), .Z(n15731) );
  XNOR U16756 ( .A(n15721), .B(n15732), .Z(n15723) );
  XOR U16757 ( .A(n15733), .B(n15734), .Z(n15721) );
  AND U16758 ( .A(n15735), .B(n15736), .Z(n15734) );
  XNOR U16759 ( .A(n15737), .B(n15733), .Z(n15736) );
  XOR U16760 ( .A(n15738), .B(e_input[739]), .Z(n15729) );
  IV U16761 ( .A(n15727), .Z(n15738) );
  XOR U16762 ( .A(n15739), .B(n15740), .Z(n15727) );
  AND U16763 ( .A(n15741), .B(n15742), .Z(n15740) );
  XNOR U16764 ( .A(n15739), .B(n7872), .Z(n15742) );
  XNOR U16765 ( .A(n15735), .B(n15737), .Z(n7872) );
  NAND U16766 ( .A(n15743), .B(e_input[738]), .Z(n15737) );
  NAND U16767 ( .A(n12323), .B(e_input[738]), .Z(n15743) );
  XNOR U16768 ( .A(n15733), .B(n15744), .Z(n15735) );
  XOR U16769 ( .A(n15745), .B(n15746), .Z(n15733) );
  AND U16770 ( .A(n15747), .B(n15748), .Z(n15746) );
  XNOR U16771 ( .A(n15749), .B(n15745), .Z(n15748) );
  XOR U16772 ( .A(n15750), .B(e_input[738]), .Z(n15741) );
  IV U16773 ( .A(n15739), .Z(n15750) );
  XOR U16774 ( .A(n15751), .B(n15752), .Z(n15739) );
  AND U16775 ( .A(n15753), .B(n15754), .Z(n15752) );
  XNOR U16776 ( .A(n15751), .B(n7878), .Z(n15754) );
  XNOR U16777 ( .A(n15747), .B(n15749), .Z(n7878) );
  NAND U16778 ( .A(n15755), .B(e_input[737]), .Z(n15749) );
  NAND U16779 ( .A(n12323), .B(e_input[737]), .Z(n15755) );
  XNOR U16780 ( .A(n15745), .B(n15756), .Z(n15747) );
  XOR U16781 ( .A(n15757), .B(n15758), .Z(n15745) );
  AND U16782 ( .A(n15759), .B(n15760), .Z(n15758) );
  XNOR U16783 ( .A(n15761), .B(n15757), .Z(n15760) );
  XOR U16784 ( .A(n15762), .B(e_input[737]), .Z(n15753) );
  IV U16785 ( .A(n15751), .Z(n15762) );
  XOR U16786 ( .A(n15763), .B(n15764), .Z(n15751) );
  AND U16787 ( .A(n15765), .B(n15766), .Z(n15764) );
  XNOR U16788 ( .A(n15763), .B(n7884), .Z(n15766) );
  XNOR U16789 ( .A(n15759), .B(n15761), .Z(n7884) );
  NAND U16790 ( .A(n15767), .B(e_input[736]), .Z(n15761) );
  NAND U16791 ( .A(n12323), .B(e_input[736]), .Z(n15767) );
  XNOR U16792 ( .A(n15757), .B(n15768), .Z(n15759) );
  XOR U16793 ( .A(n15769), .B(n15770), .Z(n15757) );
  AND U16794 ( .A(n15771), .B(n15772), .Z(n15770) );
  XNOR U16795 ( .A(n15773), .B(n15769), .Z(n15772) );
  XOR U16796 ( .A(n15774), .B(e_input[736]), .Z(n15765) );
  IV U16797 ( .A(n15763), .Z(n15774) );
  XOR U16798 ( .A(n15775), .B(n15776), .Z(n15763) );
  AND U16799 ( .A(n15777), .B(n15778), .Z(n15776) );
  XNOR U16800 ( .A(n15775), .B(n7890), .Z(n15778) );
  XNOR U16801 ( .A(n15771), .B(n15773), .Z(n7890) );
  NAND U16802 ( .A(n15779), .B(e_input[735]), .Z(n15773) );
  NAND U16803 ( .A(n12323), .B(e_input[735]), .Z(n15779) );
  XNOR U16804 ( .A(n15769), .B(n15780), .Z(n15771) );
  XOR U16805 ( .A(n15781), .B(n15782), .Z(n15769) );
  AND U16806 ( .A(n15783), .B(n15784), .Z(n15782) );
  XNOR U16807 ( .A(n15785), .B(n15781), .Z(n15784) );
  XOR U16808 ( .A(n15786), .B(e_input[735]), .Z(n15777) );
  IV U16809 ( .A(n15775), .Z(n15786) );
  XOR U16810 ( .A(n15787), .B(n15788), .Z(n15775) );
  AND U16811 ( .A(n15789), .B(n15790), .Z(n15788) );
  XNOR U16812 ( .A(n15787), .B(n7896), .Z(n15790) );
  XNOR U16813 ( .A(n15783), .B(n15785), .Z(n7896) );
  NAND U16814 ( .A(n15791), .B(e_input[734]), .Z(n15785) );
  NAND U16815 ( .A(n12323), .B(e_input[734]), .Z(n15791) );
  XNOR U16816 ( .A(n15781), .B(n15792), .Z(n15783) );
  XOR U16817 ( .A(n15793), .B(n15794), .Z(n15781) );
  AND U16818 ( .A(n15795), .B(n15796), .Z(n15794) );
  XNOR U16819 ( .A(n15797), .B(n15793), .Z(n15796) );
  XOR U16820 ( .A(n15798), .B(e_input[734]), .Z(n15789) );
  IV U16821 ( .A(n15787), .Z(n15798) );
  XOR U16822 ( .A(n15799), .B(n15800), .Z(n15787) );
  AND U16823 ( .A(n15801), .B(n15802), .Z(n15800) );
  XNOR U16824 ( .A(n15799), .B(n7902), .Z(n15802) );
  XNOR U16825 ( .A(n15795), .B(n15797), .Z(n7902) );
  NAND U16826 ( .A(n15803), .B(e_input[733]), .Z(n15797) );
  NAND U16827 ( .A(n12323), .B(e_input[733]), .Z(n15803) );
  XNOR U16828 ( .A(n15793), .B(n15804), .Z(n15795) );
  XOR U16829 ( .A(n15805), .B(n15806), .Z(n15793) );
  AND U16830 ( .A(n15807), .B(n15808), .Z(n15806) );
  XNOR U16831 ( .A(n15809), .B(n15805), .Z(n15808) );
  XOR U16832 ( .A(n15810), .B(e_input[733]), .Z(n15801) );
  IV U16833 ( .A(n15799), .Z(n15810) );
  XOR U16834 ( .A(n15811), .B(n15812), .Z(n15799) );
  AND U16835 ( .A(n15813), .B(n15814), .Z(n15812) );
  XNOR U16836 ( .A(n15811), .B(n7908), .Z(n15814) );
  XNOR U16837 ( .A(n15807), .B(n15809), .Z(n7908) );
  NAND U16838 ( .A(n15815), .B(e_input[732]), .Z(n15809) );
  NAND U16839 ( .A(n12323), .B(e_input[732]), .Z(n15815) );
  XNOR U16840 ( .A(n15805), .B(n15816), .Z(n15807) );
  XOR U16841 ( .A(n15817), .B(n15818), .Z(n15805) );
  AND U16842 ( .A(n15819), .B(n15820), .Z(n15818) );
  XNOR U16843 ( .A(n15821), .B(n15817), .Z(n15820) );
  XOR U16844 ( .A(n15822), .B(e_input[732]), .Z(n15813) );
  IV U16845 ( .A(n15811), .Z(n15822) );
  XOR U16846 ( .A(n15823), .B(n15824), .Z(n15811) );
  AND U16847 ( .A(n15825), .B(n15826), .Z(n15824) );
  XNOR U16848 ( .A(n15823), .B(n7914), .Z(n15826) );
  XNOR U16849 ( .A(n15819), .B(n15821), .Z(n7914) );
  NAND U16850 ( .A(n15827), .B(e_input[731]), .Z(n15821) );
  NAND U16851 ( .A(n12323), .B(e_input[731]), .Z(n15827) );
  XNOR U16852 ( .A(n15817), .B(n15828), .Z(n15819) );
  XOR U16853 ( .A(n15829), .B(n15830), .Z(n15817) );
  AND U16854 ( .A(n15831), .B(n15832), .Z(n15830) );
  XNOR U16855 ( .A(n15833), .B(n15829), .Z(n15832) );
  XOR U16856 ( .A(n15834), .B(e_input[731]), .Z(n15825) );
  IV U16857 ( .A(n15823), .Z(n15834) );
  XOR U16858 ( .A(n15835), .B(n15836), .Z(n15823) );
  AND U16859 ( .A(n15837), .B(n15838), .Z(n15836) );
  XNOR U16860 ( .A(n15835), .B(n7920), .Z(n15838) );
  XNOR U16861 ( .A(n15831), .B(n15833), .Z(n7920) );
  NAND U16862 ( .A(n15839), .B(e_input[730]), .Z(n15833) );
  NAND U16863 ( .A(n12323), .B(e_input[730]), .Z(n15839) );
  XNOR U16864 ( .A(n15829), .B(n15840), .Z(n15831) );
  XOR U16865 ( .A(n15841), .B(n15842), .Z(n15829) );
  AND U16866 ( .A(n15843), .B(n15844), .Z(n15842) );
  XNOR U16867 ( .A(n15845), .B(n15841), .Z(n15844) );
  XOR U16868 ( .A(n15846), .B(e_input[730]), .Z(n15837) );
  IV U16869 ( .A(n15835), .Z(n15846) );
  XOR U16870 ( .A(n15847), .B(n15848), .Z(n15835) );
  AND U16871 ( .A(n15849), .B(n15850), .Z(n15848) );
  XNOR U16872 ( .A(n15847), .B(n7926), .Z(n15850) );
  XNOR U16873 ( .A(n15843), .B(n15845), .Z(n7926) );
  NAND U16874 ( .A(n15851), .B(e_input[729]), .Z(n15845) );
  NAND U16875 ( .A(n12323), .B(e_input[729]), .Z(n15851) );
  XNOR U16876 ( .A(n15841), .B(n15852), .Z(n15843) );
  XOR U16877 ( .A(n15853), .B(n15854), .Z(n15841) );
  AND U16878 ( .A(n15855), .B(n15856), .Z(n15854) );
  XNOR U16879 ( .A(n15857), .B(n15853), .Z(n15856) );
  XOR U16880 ( .A(n15858), .B(e_input[729]), .Z(n15849) );
  IV U16881 ( .A(n15847), .Z(n15858) );
  XOR U16882 ( .A(n15859), .B(n15860), .Z(n15847) );
  AND U16883 ( .A(n15861), .B(n15862), .Z(n15860) );
  XNOR U16884 ( .A(n15859), .B(n7932), .Z(n15862) );
  XNOR U16885 ( .A(n15855), .B(n15857), .Z(n7932) );
  NAND U16886 ( .A(n15863), .B(e_input[728]), .Z(n15857) );
  NAND U16887 ( .A(n12323), .B(e_input[728]), .Z(n15863) );
  XNOR U16888 ( .A(n15853), .B(n15864), .Z(n15855) );
  XOR U16889 ( .A(n15865), .B(n15866), .Z(n15853) );
  AND U16890 ( .A(n15867), .B(n15868), .Z(n15866) );
  XNOR U16891 ( .A(n15869), .B(n15865), .Z(n15868) );
  XOR U16892 ( .A(n15870), .B(e_input[728]), .Z(n15861) );
  IV U16893 ( .A(n15859), .Z(n15870) );
  XOR U16894 ( .A(n15871), .B(n15872), .Z(n15859) );
  AND U16895 ( .A(n15873), .B(n15874), .Z(n15872) );
  XNOR U16896 ( .A(n15871), .B(n7938), .Z(n15874) );
  XNOR U16897 ( .A(n15867), .B(n15869), .Z(n7938) );
  NAND U16898 ( .A(n15875), .B(e_input[727]), .Z(n15869) );
  NAND U16899 ( .A(n12323), .B(e_input[727]), .Z(n15875) );
  XNOR U16900 ( .A(n15865), .B(n15876), .Z(n15867) );
  XOR U16901 ( .A(n15877), .B(n15878), .Z(n15865) );
  AND U16902 ( .A(n15879), .B(n15880), .Z(n15878) );
  XNOR U16903 ( .A(n15881), .B(n15877), .Z(n15880) );
  XOR U16904 ( .A(n15882), .B(e_input[727]), .Z(n15873) );
  IV U16905 ( .A(n15871), .Z(n15882) );
  XOR U16906 ( .A(n15883), .B(n15884), .Z(n15871) );
  AND U16907 ( .A(n15885), .B(n15886), .Z(n15884) );
  XNOR U16908 ( .A(n15883), .B(n7944), .Z(n15886) );
  XNOR U16909 ( .A(n15879), .B(n15881), .Z(n7944) );
  NAND U16910 ( .A(n15887), .B(e_input[726]), .Z(n15881) );
  NAND U16911 ( .A(n12323), .B(e_input[726]), .Z(n15887) );
  XNOR U16912 ( .A(n15877), .B(n15888), .Z(n15879) );
  XOR U16913 ( .A(n15889), .B(n15890), .Z(n15877) );
  AND U16914 ( .A(n15891), .B(n15892), .Z(n15890) );
  XNOR U16915 ( .A(n15893), .B(n15889), .Z(n15892) );
  XOR U16916 ( .A(n15894), .B(e_input[726]), .Z(n15885) );
  IV U16917 ( .A(n15883), .Z(n15894) );
  XOR U16918 ( .A(n15895), .B(n15896), .Z(n15883) );
  AND U16919 ( .A(n15897), .B(n15898), .Z(n15896) );
  XNOR U16920 ( .A(n15895), .B(n7950), .Z(n15898) );
  XNOR U16921 ( .A(n15891), .B(n15893), .Z(n7950) );
  NAND U16922 ( .A(n15899), .B(e_input[725]), .Z(n15893) );
  NAND U16923 ( .A(n12323), .B(e_input[725]), .Z(n15899) );
  XNOR U16924 ( .A(n15889), .B(n15900), .Z(n15891) );
  XOR U16925 ( .A(n15901), .B(n15902), .Z(n15889) );
  AND U16926 ( .A(n15903), .B(n15904), .Z(n15902) );
  XNOR U16927 ( .A(n15905), .B(n15901), .Z(n15904) );
  XOR U16928 ( .A(n15906), .B(e_input[725]), .Z(n15897) );
  IV U16929 ( .A(n15895), .Z(n15906) );
  XOR U16930 ( .A(n15907), .B(n15908), .Z(n15895) );
  AND U16931 ( .A(n15909), .B(n15910), .Z(n15908) );
  XNOR U16932 ( .A(n15907), .B(n7956), .Z(n15910) );
  XNOR U16933 ( .A(n15903), .B(n15905), .Z(n7956) );
  NAND U16934 ( .A(n15911), .B(e_input[724]), .Z(n15905) );
  NAND U16935 ( .A(n12323), .B(e_input[724]), .Z(n15911) );
  XNOR U16936 ( .A(n15901), .B(n15912), .Z(n15903) );
  XOR U16937 ( .A(n15913), .B(n15914), .Z(n15901) );
  AND U16938 ( .A(n15915), .B(n15916), .Z(n15914) );
  XNOR U16939 ( .A(n15917), .B(n15913), .Z(n15916) );
  XOR U16940 ( .A(n15918), .B(e_input[724]), .Z(n15909) );
  IV U16941 ( .A(n15907), .Z(n15918) );
  XOR U16942 ( .A(n15919), .B(n15920), .Z(n15907) );
  AND U16943 ( .A(n15921), .B(n15922), .Z(n15920) );
  XNOR U16944 ( .A(n15919), .B(n7962), .Z(n15922) );
  XNOR U16945 ( .A(n15915), .B(n15917), .Z(n7962) );
  NAND U16946 ( .A(n15923), .B(e_input[723]), .Z(n15917) );
  NAND U16947 ( .A(n12323), .B(e_input[723]), .Z(n15923) );
  XNOR U16948 ( .A(n15913), .B(n15924), .Z(n15915) );
  XOR U16949 ( .A(n15925), .B(n15926), .Z(n15913) );
  AND U16950 ( .A(n15927), .B(n15928), .Z(n15926) );
  XNOR U16951 ( .A(n15929), .B(n15925), .Z(n15928) );
  XOR U16952 ( .A(n15930), .B(e_input[723]), .Z(n15921) );
  IV U16953 ( .A(n15919), .Z(n15930) );
  XOR U16954 ( .A(n15931), .B(n15932), .Z(n15919) );
  AND U16955 ( .A(n15933), .B(n15934), .Z(n15932) );
  XNOR U16956 ( .A(n15931), .B(n7968), .Z(n15934) );
  XNOR U16957 ( .A(n15927), .B(n15929), .Z(n7968) );
  NAND U16958 ( .A(n15935), .B(e_input[722]), .Z(n15929) );
  NAND U16959 ( .A(n12323), .B(e_input[722]), .Z(n15935) );
  XNOR U16960 ( .A(n15925), .B(n15936), .Z(n15927) );
  XOR U16961 ( .A(n15937), .B(n15938), .Z(n15925) );
  AND U16962 ( .A(n15939), .B(n15940), .Z(n15938) );
  XNOR U16963 ( .A(n15941), .B(n15937), .Z(n15940) );
  XOR U16964 ( .A(n15942), .B(e_input[722]), .Z(n15933) );
  IV U16965 ( .A(n15931), .Z(n15942) );
  XOR U16966 ( .A(n15943), .B(n15944), .Z(n15931) );
  AND U16967 ( .A(n15945), .B(n15946), .Z(n15944) );
  XNOR U16968 ( .A(n15943), .B(n7974), .Z(n15946) );
  XNOR U16969 ( .A(n15939), .B(n15941), .Z(n7974) );
  NAND U16970 ( .A(n15947), .B(e_input[721]), .Z(n15941) );
  NAND U16971 ( .A(n12323), .B(e_input[721]), .Z(n15947) );
  XNOR U16972 ( .A(n15937), .B(n15948), .Z(n15939) );
  XOR U16973 ( .A(n15949), .B(n15950), .Z(n15937) );
  AND U16974 ( .A(n15951), .B(n15952), .Z(n15950) );
  XNOR U16975 ( .A(n15953), .B(n15949), .Z(n15952) );
  XOR U16976 ( .A(n15954), .B(e_input[721]), .Z(n15945) );
  IV U16977 ( .A(n15943), .Z(n15954) );
  XOR U16978 ( .A(n15955), .B(n15956), .Z(n15943) );
  AND U16979 ( .A(n15957), .B(n15958), .Z(n15956) );
  XNOR U16980 ( .A(n15955), .B(n7980), .Z(n15958) );
  XNOR U16981 ( .A(n15951), .B(n15953), .Z(n7980) );
  NAND U16982 ( .A(n15959), .B(e_input[720]), .Z(n15953) );
  NAND U16983 ( .A(n12323), .B(e_input[720]), .Z(n15959) );
  XNOR U16984 ( .A(n15949), .B(n15960), .Z(n15951) );
  XOR U16985 ( .A(n15961), .B(n15962), .Z(n15949) );
  AND U16986 ( .A(n15963), .B(n15964), .Z(n15962) );
  XNOR U16987 ( .A(n15965), .B(n15961), .Z(n15964) );
  XOR U16988 ( .A(n15966), .B(e_input[720]), .Z(n15957) );
  IV U16989 ( .A(n15955), .Z(n15966) );
  XOR U16990 ( .A(n15967), .B(n15968), .Z(n15955) );
  AND U16991 ( .A(n15969), .B(n15970), .Z(n15968) );
  XNOR U16992 ( .A(n15967), .B(n7986), .Z(n15970) );
  XNOR U16993 ( .A(n15963), .B(n15965), .Z(n7986) );
  NAND U16994 ( .A(n15971), .B(e_input[719]), .Z(n15965) );
  NAND U16995 ( .A(n12323), .B(e_input[719]), .Z(n15971) );
  XNOR U16996 ( .A(n15961), .B(n15972), .Z(n15963) );
  XOR U16997 ( .A(n15973), .B(n15974), .Z(n15961) );
  AND U16998 ( .A(n15975), .B(n15976), .Z(n15974) );
  XNOR U16999 ( .A(n15977), .B(n15973), .Z(n15976) );
  XOR U17000 ( .A(n15978), .B(e_input[719]), .Z(n15969) );
  IV U17001 ( .A(n15967), .Z(n15978) );
  XOR U17002 ( .A(n15979), .B(n15980), .Z(n15967) );
  AND U17003 ( .A(n15981), .B(n15982), .Z(n15980) );
  XNOR U17004 ( .A(n15979), .B(n7992), .Z(n15982) );
  XNOR U17005 ( .A(n15975), .B(n15977), .Z(n7992) );
  NAND U17006 ( .A(n15983), .B(e_input[718]), .Z(n15977) );
  NAND U17007 ( .A(n12323), .B(e_input[718]), .Z(n15983) );
  XNOR U17008 ( .A(n15973), .B(n15984), .Z(n15975) );
  XOR U17009 ( .A(n15985), .B(n15986), .Z(n15973) );
  AND U17010 ( .A(n15987), .B(n15988), .Z(n15986) );
  XNOR U17011 ( .A(n15989), .B(n15985), .Z(n15988) );
  XOR U17012 ( .A(n15990), .B(e_input[718]), .Z(n15981) );
  IV U17013 ( .A(n15979), .Z(n15990) );
  XOR U17014 ( .A(n15991), .B(n15992), .Z(n15979) );
  AND U17015 ( .A(n15993), .B(n15994), .Z(n15992) );
  XNOR U17016 ( .A(n15991), .B(n7998), .Z(n15994) );
  XNOR U17017 ( .A(n15987), .B(n15989), .Z(n7998) );
  NAND U17018 ( .A(n15995), .B(e_input[717]), .Z(n15989) );
  NAND U17019 ( .A(n12323), .B(e_input[717]), .Z(n15995) );
  XNOR U17020 ( .A(n15985), .B(n15996), .Z(n15987) );
  XOR U17021 ( .A(n15997), .B(n15998), .Z(n15985) );
  AND U17022 ( .A(n15999), .B(n16000), .Z(n15998) );
  XNOR U17023 ( .A(n16001), .B(n15997), .Z(n16000) );
  XOR U17024 ( .A(n16002), .B(e_input[717]), .Z(n15993) );
  IV U17025 ( .A(n15991), .Z(n16002) );
  XOR U17026 ( .A(n16003), .B(n16004), .Z(n15991) );
  AND U17027 ( .A(n16005), .B(n16006), .Z(n16004) );
  XNOR U17028 ( .A(n16003), .B(n8004), .Z(n16006) );
  XNOR U17029 ( .A(n15999), .B(n16001), .Z(n8004) );
  NAND U17030 ( .A(n16007), .B(e_input[716]), .Z(n16001) );
  NAND U17031 ( .A(n12323), .B(e_input[716]), .Z(n16007) );
  XNOR U17032 ( .A(n15997), .B(n16008), .Z(n15999) );
  XOR U17033 ( .A(n16009), .B(n16010), .Z(n15997) );
  AND U17034 ( .A(n16011), .B(n16012), .Z(n16010) );
  XNOR U17035 ( .A(n16013), .B(n16009), .Z(n16012) );
  XOR U17036 ( .A(n16014), .B(e_input[716]), .Z(n16005) );
  IV U17037 ( .A(n16003), .Z(n16014) );
  XOR U17038 ( .A(n16015), .B(n16016), .Z(n16003) );
  AND U17039 ( .A(n16017), .B(n16018), .Z(n16016) );
  XNOR U17040 ( .A(n16015), .B(n8010), .Z(n16018) );
  XNOR U17041 ( .A(n16011), .B(n16013), .Z(n8010) );
  NAND U17042 ( .A(n16019), .B(e_input[715]), .Z(n16013) );
  NAND U17043 ( .A(n12323), .B(e_input[715]), .Z(n16019) );
  XNOR U17044 ( .A(n16009), .B(n16020), .Z(n16011) );
  XOR U17045 ( .A(n16021), .B(n16022), .Z(n16009) );
  AND U17046 ( .A(n16023), .B(n16024), .Z(n16022) );
  XNOR U17047 ( .A(n16025), .B(n16021), .Z(n16024) );
  XOR U17048 ( .A(n16026), .B(e_input[715]), .Z(n16017) );
  IV U17049 ( .A(n16015), .Z(n16026) );
  XOR U17050 ( .A(n16027), .B(n16028), .Z(n16015) );
  AND U17051 ( .A(n16029), .B(n16030), .Z(n16028) );
  XNOR U17052 ( .A(n16027), .B(n8016), .Z(n16030) );
  XNOR U17053 ( .A(n16023), .B(n16025), .Z(n8016) );
  NAND U17054 ( .A(n16031), .B(e_input[714]), .Z(n16025) );
  NAND U17055 ( .A(n12323), .B(e_input[714]), .Z(n16031) );
  XNOR U17056 ( .A(n16021), .B(n16032), .Z(n16023) );
  XOR U17057 ( .A(n16033), .B(n16034), .Z(n16021) );
  AND U17058 ( .A(n16035), .B(n16036), .Z(n16034) );
  XNOR U17059 ( .A(n16037), .B(n16033), .Z(n16036) );
  XOR U17060 ( .A(n16038), .B(e_input[714]), .Z(n16029) );
  IV U17061 ( .A(n16027), .Z(n16038) );
  XOR U17062 ( .A(n16039), .B(n16040), .Z(n16027) );
  AND U17063 ( .A(n16041), .B(n16042), .Z(n16040) );
  XNOR U17064 ( .A(n16039), .B(n8022), .Z(n16042) );
  XNOR U17065 ( .A(n16035), .B(n16037), .Z(n8022) );
  NAND U17066 ( .A(n16043), .B(e_input[713]), .Z(n16037) );
  NAND U17067 ( .A(n12323), .B(e_input[713]), .Z(n16043) );
  XNOR U17068 ( .A(n16033), .B(n16044), .Z(n16035) );
  XOR U17069 ( .A(n16045), .B(n16046), .Z(n16033) );
  AND U17070 ( .A(n16047), .B(n16048), .Z(n16046) );
  XNOR U17071 ( .A(n16049), .B(n16045), .Z(n16048) );
  XOR U17072 ( .A(n16050), .B(e_input[713]), .Z(n16041) );
  IV U17073 ( .A(n16039), .Z(n16050) );
  XOR U17074 ( .A(n16051), .B(n16052), .Z(n16039) );
  AND U17075 ( .A(n16053), .B(n16054), .Z(n16052) );
  XNOR U17076 ( .A(n16051), .B(n8028), .Z(n16054) );
  XNOR U17077 ( .A(n16047), .B(n16049), .Z(n8028) );
  NAND U17078 ( .A(n16055), .B(e_input[712]), .Z(n16049) );
  NAND U17079 ( .A(n12323), .B(e_input[712]), .Z(n16055) );
  XNOR U17080 ( .A(n16045), .B(n16056), .Z(n16047) );
  XOR U17081 ( .A(n16057), .B(n16058), .Z(n16045) );
  AND U17082 ( .A(n16059), .B(n16060), .Z(n16058) );
  XNOR U17083 ( .A(n16061), .B(n16057), .Z(n16060) );
  XOR U17084 ( .A(n16062), .B(e_input[712]), .Z(n16053) );
  IV U17085 ( .A(n16051), .Z(n16062) );
  XOR U17086 ( .A(n16063), .B(n16064), .Z(n16051) );
  AND U17087 ( .A(n16065), .B(n16066), .Z(n16064) );
  XNOR U17088 ( .A(n16063), .B(n8034), .Z(n16066) );
  XNOR U17089 ( .A(n16059), .B(n16061), .Z(n8034) );
  NAND U17090 ( .A(n16067), .B(e_input[711]), .Z(n16061) );
  NAND U17091 ( .A(n12323), .B(e_input[711]), .Z(n16067) );
  XNOR U17092 ( .A(n16057), .B(n16068), .Z(n16059) );
  XOR U17093 ( .A(n16069), .B(n16070), .Z(n16057) );
  AND U17094 ( .A(n16071), .B(n16072), .Z(n16070) );
  XNOR U17095 ( .A(n16073), .B(n16069), .Z(n16072) );
  XOR U17096 ( .A(n16074), .B(e_input[711]), .Z(n16065) );
  IV U17097 ( .A(n16063), .Z(n16074) );
  XOR U17098 ( .A(n16075), .B(n16076), .Z(n16063) );
  AND U17099 ( .A(n16077), .B(n16078), .Z(n16076) );
  XNOR U17100 ( .A(n16075), .B(n8040), .Z(n16078) );
  XNOR U17101 ( .A(n16071), .B(n16073), .Z(n8040) );
  NAND U17102 ( .A(n16079), .B(e_input[710]), .Z(n16073) );
  NAND U17103 ( .A(n12323), .B(e_input[710]), .Z(n16079) );
  XNOR U17104 ( .A(n16069), .B(n16080), .Z(n16071) );
  XOR U17105 ( .A(n16081), .B(n16082), .Z(n16069) );
  AND U17106 ( .A(n16083), .B(n16084), .Z(n16082) );
  XNOR U17107 ( .A(n16085), .B(n16081), .Z(n16084) );
  XOR U17108 ( .A(n16086), .B(e_input[710]), .Z(n16077) );
  IV U17109 ( .A(n16075), .Z(n16086) );
  XOR U17110 ( .A(n16087), .B(n16088), .Z(n16075) );
  AND U17111 ( .A(n16089), .B(n16090), .Z(n16088) );
  XNOR U17112 ( .A(n16087), .B(n8046), .Z(n16090) );
  XNOR U17113 ( .A(n16083), .B(n16085), .Z(n8046) );
  NAND U17114 ( .A(n16091), .B(e_input[709]), .Z(n16085) );
  NAND U17115 ( .A(n12323), .B(e_input[709]), .Z(n16091) );
  XNOR U17116 ( .A(n16081), .B(n16092), .Z(n16083) );
  XOR U17117 ( .A(n16093), .B(n16094), .Z(n16081) );
  AND U17118 ( .A(n16095), .B(n16096), .Z(n16094) );
  XNOR U17119 ( .A(n16097), .B(n16093), .Z(n16096) );
  XOR U17120 ( .A(n16098), .B(e_input[709]), .Z(n16089) );
  IV U17121 ( .A(n16087), .Z(n16098) );
  XOR U17122 ( .A(n16099), .B(n16100), .Z(n16087) );
  AND U17123 ( .A(n16101), .B(n16102), .Z(n16100) );
  XNOR U17124 ( .A(n16099), .B(n8052), .Z(n16102) );
  XNOR U17125 ( .A(n16095), .B(n16097), .Z(n8052) );
  NAND U17126 ( .A(n16103), .B(e_input[708]), .Z(n16097) );
  NAND U17127 ( .A(n12323), .B(e_input[708]), .Z(n16103) );
  XNOR U17128 ( .A(n16093), .B(n16104), .Z(n16095) );
  XOR U17129 ( .A(n16105), .B(n16106), .Z(n16093) );
  AND U17130 ( .A(n16107), .B(n16108), .Z(n16106) );
  XNOR U17131 ( .A(n16109), .B(n16105), .Z(n16108) );
  XOR U17132 ( .A(n16110), .B(e_input[708]), .Z(n16101) );
  IV U17133 ( .A(n16099), .Z(n16110) );
  XOR U17134 ( .A(n16111), .B(n16112), .Z(n16099) );
  AND U17135 ( .A(n16113), .B(n16114), .Z(n16112) );
  XNOR U17136 ( .A(n16111), .B(n8058), .Z(n16114) );
  XNOR U17137 ( .A(n16107), .B(n16109), .Z(n8058) );
  NAND U17138 ( .A(n16115), .B(e_input[707]), .Z(n16109) );
  NAND U17139 ( .A(n12323), .B(e_input[707]), .Z(n16115) );
  XNOR U17140 ( .A(n16105), .B(n16116), .Z(n16107) );
  XOR U17141 ( .A(n16117), .B(n16118), .Z(n16105) );
  AND U17142 ( .A(n16119), .B(n16120), .Z(n16118) );
  XNOR U17143 ( .A(n16121), .B(n16117), .Z(n16120) );
  XOR U17144 ( .A(n16122), .B(e_input[707]), .Z(n16113) );
  IV U17145 ( .A(n16111), .Z(n16122) );
  XOR U17146 ( .A(n16123), .B(n16124), .Z(n16111) );
  AND U17147 ( .A(n16125), .B(n16126), .Z(n16124) );
  XNOR U17148 ( .A(n16123), .B(n8064), .Z(n16126) );
  XNOR U17149 ( .A(n16119), .B(n16121), .Z(n8064) );
  NAND U17150 ( .A(n16127), .B(e_input[706]), .Z(n16121) );
  NAND U17151 ( .A(n12323), .B(e_input[706]), .Z(n16127) );
  XNOR U17152 ( .A(n16117), .B(n16128), .Z(n16119) );
  XOR U17153 ( .A(n16129), .B(n16130), .Z(n16117) );
  AND U17154 ( .A(n16131), .B(n16132), .Z(n16130) );
  XNOR U17155 ( .A(n16133), .B(n16129), .Z(n16132) );
  XOR U17156 ( .A(n16134), .B(e_input[706]), .Z(n16125) );
  IV U17157 ( .A(n16123), .Z(n16134) );
  XOR U17158 ( .A(n16135), .B(n16136), .Z(n16123) );
  AND U17159 ( .A(n16137), .B(n16138), .Z(n16136) );
  XNOR U17160 ( .A(n16135), .B(n8070), .Z(n16138) );
  XNOR U17161 ( .A(n16131), .B(n16133), .Z(n8070) );
  NAND U17162 ( .A(n16139), .B(e_input[705]), .Z(n16133) );
  NAND U17163 ( .A(n12323), .B(e_input[705]), .Z(n16139) );
  XNOR U17164 ( .A(n16129), .B(n16140), .Z(n16131) );
  XOR U17165 ( .A(n16141), .B(n16142), .Z(n16129) );
  AND U17166 ( .A(n16143), .B(n16144), .Z(n16142) );
  XNOR U17167 ( .A(n16145), .B(n16141), .Z(n16144) );
  XOR U17168 ( .A(n16146), .B(e_input[705]), .Z(n16137) );
  IV U17169 ( .A(n16135), .Z(n16146) );
  XOR U17170 ( .A(n16147), .B(n16148), .Z(n16135) );
  AND U17171 ( .A(n16149), .B(n16150), .Z(n16148) );
  XNOR U17172 ( .A(n16147), .B(n8076), .Z(n16150) );
  XNOR U17173 ( .A(n16143), .B(n16145), .Z(n8076) );
  NAND U17174 ( .A(n16151), .B(e_input[704]), .Z(n16145) );
  NAND U17175 ( .A(n12323), .B(e_input[704]), .Z(n16151) );
  XNOR U17176 ( .A(n16141), .B(n16152), .Z(n16143) );
  XOR U17177 ( .A(n16153), .B(n16154), .Z(n16141) );
  AND U17178 ( .A(n16155), .B(n16156), .Z(n16154) );
  XNOR U17179 ( .A(n16157), .B(n16153), .Z(n16156) );
  XOR U17180 ( .A(n16158), .B(e_input[704]), .Z(n16149) );
  IV U17181 ( .A(n16147), .Z(n16158) );
  XOR U17182 ( .A(n16159), .B(n16160), .Z(n16147) );
  AND U17183 ( .A(n16161), .B(n16162), .Z(n16160) );
  XNOR U17184 ( .A(n16159), .B(n8082), .Z(n16162) );
  XNOR U17185 ( .A(n16155), .B(n16157), .Z(n8082) );
  NAND U17186 ( .A(n16163), .B(e_input[703]), .Z(n16157) );
  NAND U17187 ( .A(n12323), .B(e_input[703]), .Z(n16163) );
  XNOR U17188 ( .A(n16153), .B(n16164), .Z(n16155) );
  XOR U17189 ( .A(n16165), .B(n16166), .Z(n16153) );
  AND U17190 ( .A(n16167), .B(n16168), .Z(n16166) );
  XNOR U17191 ( .A(n16169), .B(n16165), .Z(n16168) );
  XOR U17192 ( .A(n16170), .B(e_input[703]), .Z(n16161) );
  IV U17193 ( .A(n16159), .Z(n16170) );
  XOR U17194 ( .A(n16171), .B(n16172), .Z(n16159) );
  AND U17195 ( .A(n16173), .B(n16174), .Z(n16172) );
  XNOR U17196 ( .A(n16171), .B(n8088), .Z(n16174) );
  XNOR U17197 ( .A(n16167), .B(n16169), .Z(n8088) );
  NAND U17198 ( .A(n16175), .B(e_input[702]), .Z(n16169) );
  NAND U17199 ( .A(n12323), .B(e_input[702]), .Z(n16175) );
  XNOR U17200 ( .A(n16165), .B(n16176), .Z(n16167) );
  XOR U17201 ( .A(n16177), .B(n16178), .Z(n16165) );
  AND U17202 ( .A(n16179), .B(n16180), .Z(n16178) );
  XNOR U17203 ( .A(n16181), .B(n16177), .Z(n16180) );
  XOR U17204 ( .A(n16182), .B(e_input[702]), .Z(n16173) );
  IV U17205 ( .A(n16171), .Z(n16182) );
  XOR U17206 ( .A(n16183), .B(n16184), .Z(n16171) );
  AND U17207 ( .A(n16185), .B(n16186), .Z(n16184) );
  XNOR U17208 ( .A(n16183), .B(n8094), .Z(n16186) );
  XNOR U17209 ( .A(n16179), .B(n16181), .Z(n8094) );
  NAND U17210 ( .A(n16187), .B(e_input[701]), .Z(n16181) );
  NAND U17211 ( .A(n12323), .B(e_input[701]), .Z(n16187) );
  XNOR U17212 ( .A(n16177), .B(n16188), .Z(n16179) );
  XOR U17213 ( .A(n16189), .B(n16190), .Z(n16177) );
  AND U17214 ( .A(n16191), .B(n16192), .Z(n16190) );
  XNOR U17215 ( .A(n16193), .B(n16189), .Z(n16192) );
  XOR U17216 ( .A(n16194), .B(e_input[701]), .Z(n16185) );
  IV U17217 ( .A(n16183), .Z(n16194) );
  XOR U17218 ( .A(n16195), .B(n16196), .Z(n16183) );
  AND U17219 ( .A(n16197), .B(n16198), .Z(n16196) );
  XNOR U17220 ( .A(n16195), .B(n8100), .Z(n16198) );
  XNOR U17221 ( .A(n16191), .B(n16193), .Z(n8100) );
  NAND U17222 ( .A(n16199), .B(e_input[700]), .Z(n16193) );
  NAND U17223 ( .A(n12323), .B(e_input[700]), .Z(n16199) );
  XNOR U17224 ( .A(n16189), .B(n16200), .Z(n16191) );
  XOR U17225 ( .A(n16201), .B(n16202), .Z(n16189) );
  AND U17226 ( .A(n16203), .B(n16204), .Z(n16202) );
  XNOR U17227 ( .A(n16205), .B(n16201), .Z(n16204) );
  XOR U17228 ( .A(n16206), .B(e_input[700]), .Z(n16197) );
  IV U17229 ( .A(n16195), .Z(n16206) );
  XOR U17230 ( .A(n16207), .B(n16208), .Z(n16195) );
  AND U17231 ( .A(n16209), .B(n16210), .Z(n16208) );
  XNOR U17232 ( .A(n16207), .B(n8106), .Z(n16210) );
  XNOR U17233 ( .A(n16203), .B(n16205), .Z(n8106) );
  NAND U17234 ( .A(n16211), .B(e_input[699]), .Z(n16205) );
  NAND U17235 ( .A(n12323), .B(e_input[699]), .Z(n16211) );
  XNOR U17236 ( .A(n16201), .B(n16212), .Z(n16203) );
  XOR U17237 ( .A(n16213), .B(n16214), .Z(n16201) );
  AND U17238 ( .A(n16215), .B(n16216), .Z(n16214) );
  XNOR U17239 ( .A(n16217), .B(n16213), .Z(n16216) );
  XOR U17240 ( .A(n16218), .B(e_input[699]), .Z(n16209) );
  IV U17241 ( .A(n16207), .Z(n16218) );
  XOR U17242 ( .A(n16219), .B(n16220), .Z(n16207) );
  AND U17243 ( .A(n16221), .B(n16222), .Z(n16220) );
  XNOR U17244 ( .A(n16219), .B(n8112), .Z(n16222) );
  XNOR U17245 ( .A(n16215), .B(n16217), .Z(n8112) );
  NAND U17246 ( .A(n16223), .B(e_input[698]), .Z(n16217) );
  NAND U17247 ( .A(n12323), .B(e_input[698]), .Z(n16223) );
  XNOR U17248 ( .A(n16213), .B(n16224), .Z(n16215) );
  XOR U17249 ( .A(n16225), .B(n16226), .Z(n16213) );
  AND U17250 ( .A(n16227), .B(n16228), .Z(n16226) );
  XNOR U17251 ( .A(n16229), .B(n16225), .Z(n16228) );
  XOR U17252 ( .A(n16230), .B(e_input[698]), .Z(n16221) );
  IV U17253 ( .A(n16219), .Z(n16230) );
  XOR U17254 ( .A(n16231), .B(n16232), .Z(n16219) );
  AND U17255 ( .A(n16233), .B(n16234), .Z(n16232) );
  XNOR U17256 ( .A(n16231), .B(n8118), .Z(n16234) );
  XNOR U17257 ( .A(n16227), .B(n16229), .Z(n8118) );
  NAND U17258 ( .A(n16235), .B(e_input[697]), .Z(n16229) );
  NAND U17259 ( .A(n12323), .B(e_input[697]), .Z(n16235) );
  XNOR U17260 ( .A(n16225), .B(n16236), .Z(n16227) );
  XOR U17261 ( .A(n16237), .B(n16238), .Z(n16225) );
  AND U17262 ( .A(n16239), .B(n16240), .Z(n16238) );
  XNOR U17263 ( .A(n16241), .B(n16237), .Z(n16240) );
  XOR U17264 ( .A(n16242), .B(e_input[697]), .Z(n16233) );
  IV U17265 ( .A(n16231), .Z(n16242) );
  XOR U17266 ( .A(n16243), .B(n16244), .Z(n16231) );
  AND U17267 ( .A(n16245), .B(n16246), .Z(n16244) );
  XNOR U17268 ( .A(n16243), .B(n8124), .Z(n16246) );
  XNOR U17269 ( .A(n16239), .B(n16241), .Z(n8124) );
  NAND U17270 ( .A(n16247), .B(e_input[696]), .Z(n16241) );
  NAND U17271 ( .A(n12323), .B(e_input[696]), .Z(n16247) );
  XNOR U17272 ( .A(n16237), .B(n16248), .Z(n16239) );
  XOR U17273 ( .A(n16249), .B(n16250), .Z(n16237) );
  AND U17274 ( .A(n16251), .B(n16252), .Z(n16250) );
  XNOR U17275 ( .A(n16253), .B(n16249), .Z(n16252) );
  XOR U17276 ( .A(n16254), .B(e_input[696]), .Z(n16245) );
  IV U17277 ( .A(n16243), .Z(n16254) );
  XOR U17278 ( .A(n16255), .B(n16256), .Z(n16243) );
  AND U17279 ( .A(n16257), .B(n16258), .Z(n16256) );
  XNOR U17280 ( .A(n16255), .B(n8130), .Z(n16258) );
  XNOR U17281 ( .A(n16251), .B(n16253), .Z(n8130) );
  NAND U17282 ( .A(n16259), .B(e_input[695]), .Z(n16253) );
  NAND U17283 ( .A(n12323), .B(e_input[695]), .Z(n16259) );
  XNOR U17284 ( .A(n16249), .B(n16260), .Z(n16251) );
  XOR U17285 ( .A(n16261), .B(n16262), .Z(n16249) );
  AND U17286 ( .A(n16263), .B(n16264), .Z(n16262) );
  XNOR U17287 ( .A(n16265), .B(n16261), .Z(n16264) );
  XOR U17288 ( .A(n16266), .B(e_input[695]), .Z(n16257) );
  IV U17289 ( .A(n16255), .Z(n16266) );
  XOR U17290 ( .A(n16267), .B(n16268), .Z(n16255) );
  AND U17291 ( .A(n16269), .B(n16270), .Z(n16268) );
  XNOR U17292 ( .A(n16267), .B(n8136), .Z(n16270) );
  XNOR U17293 ( .A(n16263), .B(n16265), .Z(n8136) );
  NAND U17294 ( .A(n16271), .B(e_input[694]), .Z(n16265) );
  NAND U17295 ( .A(n12323), .B(e_input[694]), .Z(n16271) );
  XNOR U17296 ( .A(n16261), .B(n16272), .Z(n16263) );
  XOR U17297 ( .A(n16273), .B(n16274), .Z(n16261) );
  AND U17298 ( .A(n16275), .B(n16276), .Z(n16274) );
  XNOR U17299 ( .A(n16277), .B(n16273), .Z(n16276) );
  XOR U17300 ( .A(n16278), .B(e_input[694]), .Z(n16269) );
  IV U17301 ( .A(n16267), .Z(n16278) );
  XOR U17302 ( .A(n16279), .B(n16280), .Z(n16267) );
  AND U17303 ( .A(n16281), .B(n16282), .Z(n16280) );
  XNOR U17304 ( .A(n16279), .B(n8142), .Z(n16282) );
  XNOR U17305 ( .A(n16275), .B(n16277), .Z(n8142) );
  NAND U17306 ( .A(n16283), .B(e_input[693]), .Z(n16277) );
  NAND U17307 ( .A(n12323), .B(e_input[693]), .Z(n16283) );
  XNOR U17308 ( .A(n16273), .B(n16284), .Z(n16275) );
  XOR U17309 ( .A(n16285), .B(n16286), .Z(n16273) );
  AND U17310 ( .A(n16287), .B(n16288), .Z(n16286) );
  XNOR U17311 ( .A(n16289), .B(n16285), .Z(n16288) );
  XOR U17312 ( .A(n16290), .B(e_input[693]), .Z(n16281) );
  IV U17313 ( .A(n16279), .Z(n16290) );
  XOR U17314 ( .A(n16291), .B(n16292), .Z(n16279) );
  AND U17315 ( .A(n16293), .B(n16294), .Z(n16292) );
  XNOR U17316 ( .A(n16291), .B(n8148), .Z(n16294) );
  XNOR U17317 ( .A(n16287), .B(n16289), .Z(n8148) );
  NAND U17318 ( .A(n16295), .B(e_input[692]), .Z(n16289) );
  NAND U17319 ( .A(n12323), .B(e_input[692]), .Z(n16295) );
  XNOR U17320 ( .A(n16285), .B(n16296), .Z(n16287) );
  XOR U17321 ( .A(n16297), .B(n16298), .Z(n16285) );
  AND U17322 ( .A(n16299), .B(n16300), .Z(n16298) );
  XNOR U17323 ( .A(n16301), .B(n16297), .Z(n16300) );
  XOR U17324 ( .A(n16302), .B(e_input[692]), .Z(n16293) );
  IV U17325 ( .A(n16291), .Z(n16302) );
  XOR U17326 ( .A(n16303), .B(n16304), .Z(n16291) );
  AND U17327 ( .A(n16305), .B(n16306), .Z(n16304) );
  XNOR U17328 ( .A(n16303), .B(n8154), .Z(n16306) );
  XNOR U17329 ( .A(n16299), .B(n16301), .Z(n8154) );
  NAND U17330 ( .A(n16307), .B(e_input[691]), .Z(n16301) );
  NAND U17331 ( .A(n12323), .B(e_input[691]), .Z(n16307) );
  XNOR U17332 ( .A(n16297), .B(n16308), .Z(n16299) );
  XOR U17333 ( .A(n16309), .B(n16310), .Z(n16297) );
  AND U17334 ( .A(n16311), .B(n16312), .Z(n16310) );
  XNOR U17335 ( .A(n16313), .B(n16309), .Z(n16312) );
  XOR U17336 ( .A(n16314), .B(e_input[691]), .Z(n16305) );
  IV U17337 ( .A(n16303), .Z(n16314) );
  XOR U17338 ( .A(n16315), .B(n16316), .Z(n16303) );
  AND U17339 ( .A(n16317), .B(n16318), .Z(n16316) );
  XNOR U17340 ( .A(n16315), .B(n8160), .Z(n16318) );
  XNOR U17341 ( .A(n16311), .B(n16313), .Z(n8160) );
  NAND U17342 ( .A(n16319), .B(e_input[690]), .Z(n16313) );
  NAND U17343 ( .A(n12323), .B(e_input[690]), .Z(n16319) );
  XNOR U17344 ( .A(n16309), .B(n16320), .Z(n16311) );
  XOR U17345 ( .A(n16321), .B(n16322), .Z(n16309) );
  AND U17346 ( .A(n16323), .B(n16324), .Z(n16322) );
  XNOR U17347 ( .A(n16325), .B(n16321), .Z(n16324) );
  XOR U17348 ( .A(n16326), .B(e_input[690]), .Z(n16317) );
  IV U17349 ( .A(n16315), .Z(n16326) );
  XOR U17350 ( .A(n16327), .B(n16328), .Z(n16315) );
  AND U17351 ( .A(n16329), .B(n16330), .Z(n16328) );
  XNOR U17352 ( .A(n16327), .B(n8166), .Z(n16330) );
  XNOR U17353 ( .A(n16323), .B(n16325), .Z(n8166) );
  NAND U17354 ( .A(n16331), .B(e_input[689]), .Z(n16325) );
  NAND U17355 ( .A(n12323), .B(e_input[689]), .Z(n16331) );
  XNOR U17356 ( .A(n16321), .B(n16332), .Z(n16323) );
  XOR U17357 ( .A(n16333), .B(n16334), .Z(n16321) );
  AND U17358 ( .A(n16335), .B(n16336), .Z(n16334) );
  XNOR U17359 ( .A(n16337), .B(n16333), .Z(n16336) );
  XOR U17360 ( .A(n16338), .B(e_input[689]), .Z(n16329) );
  IV U17361 ( .A(n16327), .Z(n16338) );
  XOR U17362 ( .A(n16339), .B(n16340), .Z(n16327) );
  AND U17363 ( .A(n16341), .B(n16342), .Z(n16340) );
  XNOR U17364 ( .A(n16339), .B(n8172), .Z(n16342) );
  XNOR U17365 ( .A(n16335), .B(n16337), .Z(n8172) );
  NAND U17366 ( .A(n16343), .B(e_input[688]), .Z(n16337) );
  NAND U17367 ( .A(n12323), .B(e_input[688]), .Z(n16343) );
  XNOR U17368 ( .A(n16333), .B(n16344), .Z(n16335) );
  XOR U17369 ( .A(n16345), .B(n16346), .Z(n16333) );
  AND U17370 ( .A(n16347), .B(n16348), .Z(n16346) );
  XNOR U17371 ( .A(n16349), .B(n16345), .Z(n16348) );
  XOR U17372 ( .A(n16350), .B(e_input[688]), .Z(n16341) );
  IV U17373 ( .A(n16339), .Z(n16350) );
  XOR U17374 ( .A(n16351), .B(n16352), .Z(n16339) );
  AND U17375 ( .A(n16353), .B(n16354), .Z(n16352) );
  XNOR U17376 ( .A(n16351), .B(n8178), .Z(n16354) );
  XNOR U17377 ( .A(n16347), .B(n16349), .Z(n8178) );
  NAND U17378 ( .A(n16355), .B(e_input[687]), .Z(n16349) );
  NAND U17379 ( .A(n12323), .B(e_input[687]), .Z(n16355) );
  XNOR U17380 ( .A(n16345), .B(n16356), .Z(n16347) );
  XOR U17381 ( .A(n16357), .B(n16358), .Z(n16345) );
  AND U17382 ( .A(n16359), .B(n16360), .Z(n16358) );
  XNOR U17383 ( .A(n16361), .B(n16357), .Z(n16360) );
  XOR U17384 ( .A(n16362), .B(e_input[687]), .Z(n16353) );
  IV U17385 ( .A(n16351), .Z(n16362) );
  XOR U17386 ( .A(n16363), .B(n16364), .Z(n16351) );
  AND U17387 ( .A(n16365), .B(n16366), .Z(n16364) );
  XNOR U17388 ( .A(n16363), .B(n8184), .Z(n16366) );
  XNOR U17389 ( .A(n16359), .B(n16361), .Z(n8184) );
  NAND U17390 ( .A(n16367), .B(e_input[686]), .Z(n16361) );
  NAND U17391 ( .A(n12323), .B(e_input[686]), .Z(n16367) );
  XNOR U17392 ( .A(n16357), .B(n16368), .Z(n16359) );
  XOR U17393 ( .A(n16369), .B(n16370), .Z(n16357) );
  AND U17394 ( .A(n16371), .B(n16372), .Z(n16370) );
  XNOR U17395 ( .A(n16373), .B(n16369), .Z(n16372) );
  XOR U17396 ( .A(n16374), .B(e_input[686]), .Z(n16365) );
  IV U17397 ( .A(n16363), .Z(n16374) );
  XOR U17398 ( .A(n16375), .B(n16376), .Z(n16363) );
  AND U17399 ( .A(n16377), .B(n16378), .Z(n16376) );
  XNOR U17400 ( .A(n16375), .B(n8190), .Z(n16378) );
  XNOR U17401 ( .A(n16371), .B(n16373), .Z(n8190) );
  NAND U17402 ( .A(n16379), .B(e_input[685]), .Z(n16373) );
  NAND U17403 ( .A(n12323), .B(e_input[685]), .Z(n16379) );
  XNOR U17404 ( .A(n16369), .B(n16380), .Z(n16371) );
  XOR U17405 ( .A(n16381), .B(n16382), .Z(n16369) );
  AND U17406 ( .A(n16383), .B(n16384), .Z(n16382) );
  XNOR U17407 ( .A(n16385), .B(n16381), .Z(n16384) );
  XOR U17408 ( .A(n16386), .B(e_input[685]), .Z(n16377) );
  IV U17409 ( .A(n16375), .Z(n16386) );
  XOR U17410 ( .A(n16387), .B(n16388), .Z(n16375) );
  AND U17411 ( .A(n16389), .B(n16390), .Z(n16388) );
  XNOR U17412 ( .A(n16387), .B(n8196), .Z(n16390) );
  XNOR U17413 ( .A(n16383), .B(n16385), .Z(n8196) );
  NAND U17414 ( .A(n16391), .B(e_input[684]), .Z(n16385) );
  NAND U17415 ( .A(n12323), .B(e_input[684]), .Z(n16391) );
  XNOR U17416 ( .A(n16381), .B(n16392), .Z(n16383) );
  XOR U17417 ( .A(n16393), .B(n16394), .Z(n16381) );
  AND U17418 ( .A(n16395), .B(n16396), .Z(n16394) );
  XNOR U17419 ( .A(n16397), .B(n16393), .Z(n16396) );
  XOR U17420 ( .A(n16398), .B(e_input[684]), .Z(n16389) );
  IV U17421 ( .A(n16387), .Z(n16398) );
  XOR U17422 ( .A(n16399), .B(n16400), .Z(n16387) );
  AND U17423 ( .A(n16401), .B(n16402), .Z(n16400) );
  XNOR U17424 ( .A(n16399), .B(n8202), .Z(n16402) );
  XNOR U17425 ( .A(n16395), .B(n16397), .Z(n8202) );
  NAND U17426 ( .A(n16403), .B(e_input[683]), .Z(n16397) );
  NAND U17427 ( .A(n12323), .B(e_input[683]), .Z(n16403) );
  XNOR U17428 ( .A(n16393), .B(n16404), .Z(n16395) );
  XOR U17429 ( .A(n16405), .B(n16406), .Z(n16393) );
  AND U17430 ( .A(n16407), .B(n16408), .Z(n16406) );
  XNOR U17431 ( .A(n16409), .B(n16405), .Z(n16408) );
  XOR U17432 ( .A(n16410), .B(e_input[683]), .Z(n16401) );
  IV U17433 ( .A(n16399), .Z(n16410) );
  XOR U17434 ( .A(n16411), .B(n16412), .Z(n16399) );
  AND U17435 ( .A(n16413), .B(n16414), .Z(n16412) );
  XNOR U17436 ( .A(n16411), .B(n8208), .Z(n16414) );
  XNOR U17437 ( .A(n16407), .B(n16409), .Z(n8208) );
  NAND U17438 ( .A(n16415), .B(e_input[682]), .Z(n16409) );
  NAND U17439 ( .A(n12323), .B(e_input[682]), .Z(n16415) );
  XNOR U17440 ( .A(n16405), .B(n16416), .Z(n16407) );
  XOR U17441 ( .A(n16417), .B(n16418), .Z(n16405) );
  AND U17442 ( .A(n16419), .B(n16420), .Z(n16418) );
  XNOR U17443 ( .A(n16421), .B(n16417), .Z(n16420) );
  XOR U17444 ( .A(n16422), .B(e_input[682]), .Z(n16413) );
  IV U17445 ( .A(n16411), .Z(n16422) );
  XOR U17446 ( .A(n16423), .B(n16424), .Z(n16411) );
  AND U17447 ( .A(n16425), .B(n16426), .Z(n16424) );
  XNOR U17448 ( .A(n16423), .B(n8214), .Z(n16426) );
  XNOR U17449 ( .A(n16419), .B(n16421), .Z(n8214) );
  NAND U17450 ( .A(n16427), .B(e_input[681]), .Z(n16421) );
  NAND U17451 ( .A(n12323), .B(e_input[681]), .Z(n16427) );
  XNOR U17452 ( .A(n16417), .B(n16428), .Z(n16419) );
  XOR U17453 ( .A(n16429), .B(n16430), .Z(n16417) );
  AND U17454 ( .A(n16431), .B(n16432), .Z(n16430) );
  XNOR U17455 ( .A(n16433), .B(n16429), .Z(n16432) );
  XOR U17456 ( .A(n16434), .B(e_input[681]), .Z(n16425) );
  IV U17457 ( .A(n16423), .Z(n16434) );
  XOR U17458 ( .A(n16435), .B(n16436), .Z(n16423) );
  AND U17459 ( .A(n16437), .B(n16438), .Z(n16436) );
  XNOR U17460 ( .A(n16435), .B(n8220), .Z(n16438) );
  XNOR U17461 ( .A(n16431), .B(n16433), .Z(n8220) );
  NAND U17462 ( .A(n16439), .B(e_input[680]), .Z(n16433) );
  NAND U17463 ( .A(n12323), .B(e_input[680]), .Z(n16439) );
  XNOR U17464 ( .A(n16429), .B(n16440), .Z(n16431) );
  XOR U17465 ( .A(n16441), .B(n16442), .Z(n16429) );
  AND U17466 ( .A(n16443), .B(n16444), .Z(n16442) );
  XNOR U17467 ( .A(n16445), .B(n16441), .Z(n16444) );
  XOR U17468 ( .A(n16446), .B(e_input[680]), .Z(n16437) );
  IV U17469 ( .A(n16435), .Z(n16446) );
  XOR U17470 ( .A(n16447), .B(n16448), .Z(n16435) );
  AND U17471 ( .A(n16449), .B(n16450), .Z(n16448) );
  XNOR U17472 ( .A(n16447), .B(n8226), .Z(n16450) );
  XNOR U17473 ( .A(n16443), .B(n16445), .Z(n8226) );
  NAND U17474 ( .A(n16451), .B(e_input[679]), .Z(n16445) );
  NAND U17475 ( .A(n12323), .B(e_input[679]), .Z(n16451) );
  XNOR U17476 ( .A(n16441), .B(n16452), .Z(n16443) );
  XOR U17477 ( .A(n16453), .B(n16454), .Z(n16441) );
  AND U17478 ( .A(n16455), .B(n16456), .Z(n16454) );
  XNOR U17479 ( .A(n16457), .B(n16453), .Z(n16456) );
  XOR U17480 ( .A(n16458), .B(e_input[679]), .Z(n16449) );
  IV U17481 ( .A(n16447), .Z(n16458) );
  XOR U17482 ( .A(n16459), .B(n16460), .Z(n16447) );
  AND U17483 ( .A(n16461), .B(n16462), .Z(n16460) );
  XNOR U17484 ( .A(n16459), .B(n8232), .Z(n16462) );
  XNOR U17485 ( .A(n16455), .B(n16457), .Z(n8232) );
  NAND U17486 ( .A(n16463), .B(e_input[678]), .Z(n16457) );
  NAND U17487 ( .A(n12323), .B(e_input[678]), .Z(n16463) );
  XNOR U17488 ( .A(n16453), .B(n16464), .Z(n16455) );
  XOR U17489 ( .A(n16465), .B(n16466), .Z(n16453) );
  AND U17490 ( .A(n16467), .B(n16468), .Z(n16466) );
  XNOR U17491 ( .A(n16469), .B(n16465), .Z(n16468) );
  XOR U17492 ( .A(n16470), .B(e_input[678]), .Z(n16461) );
  IV U17493 ( .A(n16459), .Z(n16470) );
  XOR U17494 ( .A(n16471), .B(n16472), .Z(n16459) );
  AND U17495 ( .A(n16473), .B(n16474), .Z(n16472) );
  XNOR U17496 ( .A(n16471), .B(n8238), .Z(n16474) );
  XNOR U17497 ( .A(n16467), .B(n16469), .Z(n8238) );
  NAND U17498 ( .A(n16475), .B(e_input[677]), .Z(n16469) );
  NAND U17499 ( .A(n12323), .B(e_input[677]), .Z(n16475) );
  XNOR U17500 ( .A(n16465), .B(n16476), .Z(n16467) );
  XOR U17501 ( .A(n16477), .B(n16478), .Z(n16465) );
  AND U17502 ( .A(n16479), .B(n16480), .Z(n16478) );
  XNOR U17503 ( .A(n16481), .B(n16477), .Z(n16480) );
  XOR U17504 ( .A(n16482), .B(e_input[677]), .Z(n16473) );
  IV U17505 ( .A(n16471), .Z(n16482) );
  XOR U17506 ( .A(n16483), .B(n16484), .Z(n16471) );
  AND U17507 ( .A(n16485), .B(n16486), .Z(n16484) );
  XNOR U17508 ( .A(n16483), .B(n8244), .Z(n16486) );
  XNOR U17509 ( .A(n16479), .B(n16481), .Z(n8244) );
  NAND U17510 ( .A(n16487), .B(e_input[676]), .Z(n16481) );
  NAND U17511 ( .A(n12323), .B(e_input[676]), .Z(n16487) );
  XNOR U17512 ( .A(n16477), .B(n16488), .Z(n16479) );
  XOR U17513 ( .A(n16489), .B(n16490), .Z(n16477) );
  AND U17514 ( .A(n16491), .B(n16492), .Z(n16490) );
  XNOR U17515 ( .A(n16493), .B(n16489), .Z(n16492) );
  XOR U17516 ( .A(n16494), .B(e_input[676]), .Z(n16485) );
  IV U17517 ( .A(n16483), .Z(n16494) );
  XOR U17518 ( .A(n16495), .B(n16496), .Z(n16483) );
  AND U17519 ( .A(n16497), .B(n16498), .Z(n16496) );
  XNOR U17520 ( .A(n16495), .B(n8250), .Z(n16498) );
  XNOR U17521 ( .A(n16491), .B(n16493), .Z(n8250) );
  NAND U17522 ( .A(n16499), .B(e_input[675]), .Z(n16493) );
  NAND U17523 ( .A(n12323), .B(e_input[675]), .Z(n16499) );
  XNOR U17524 ( .A(n16489), .B(n16500), .Z(n16491) );
  XOR U17525 ( .A(n16501), .B(n16502), .Z(n16489) );
  AND U17526 ( .A(n16503), .B(n16504), .Z(n16502) );
  XNOR U17527 ( .A(n16505), .B(n16501), .Z(n16504) );
  XOR U17528 ( .A(n16506), .B(e_input[675]), .Z(n16497) );
  IV U17529 ( .A(n16495), .Z(n16506) );
  XOR U17530 ( .A(n16507), .B(n16508), .Z(n16495) );
  AND U17531 ( .A(n16509), .B(n16510), .Z(n16508) );
  XNOR U17532 ( .A(n16507), .B(n8256), .Z(n16510) );
  XNOR U17533 ( .A(n16503), .B(n16505), .Z(n8256) );
  NAND U17534 ( .A(n16511), .B(e_input[674]), .Z(n16505) );
  NAND U17535 ( .A(n12323), .B(e_input[674]), .Z(n16511) );
  XNOR U17536 ( .A(n16501), .B(n16512), .Z(n16503) );
  XOR U17537 ( .A(n16513), .B(n16514), .Z(n16501) );
  AND U17538 ( .A(n16515), .B(n16516), .Z(n16514) );
  XNOR U17539 ( .A(n16517), .B(n16513), .Z(n16516) );
  XOR U17540 ( .A(n16518), .B(e_input[674]), .Z(n16509) );
  IV U17541 ( .A(n16507), .Z(n16518) );
  XOR U17542 ( .A(n16519), .B(n16520), .Z(n16507) );
  AND U17543 ( .A(n16521), .B(n16522), .Z(n16520) );
  XNOR U17544 ( .A(n16519), .B(n8262), .Z(n16522) );
  XNOR U17545 ( .A(n16515), .B(n16517), .Z(n8262) );
  NAND U17546 ( .A(n16523), .B(e_input[673]), .Z(n16517) );
  NAND U17547 ( .A(n12323), .B(e_input[673]), .Z(n16523) );
  XNOR U17548 ( .A(n16513), .B(n16524), .Z(n16515) );
  XOR U17549 ( .A(n16525), .B(n16526), .Z(n16513) );
  AND U17550 ( .A(n16527), .B(n16528), .Z(n16526) );
  XNOR U17551 ( .A(n16529), .B(n16525), .Z(n16528) );
  XOR U17552 ( .A(n16530), .B(e_input[673]), .Z(n16521) );
  IV U17553 ( .A(n16519), .Z(n16530) );
  XOR U17554 ( .A(n16531), .B(n16532), .Z(n16519) );
  AND U17555 ( .A(n16533), .B(n16534), .Z(n16532) );
  XNOR U17556 ( .A(n16531), .B(n8268), .Z(n16534) );
  XNOR U17557 ( .A(n16527), .B(n16529), .Z(n8268) );
  NAND U17558 ( .A(n16535), .B(e_input[672]), .Z(n16529) );
  NAND U17559 ( .A(n12323), .B(e_input[672]), .Z(n16535) );
  XNOR U17560 ( .A(n16525), .B(n16536), .Z(n16527) );
  XOR U17561 ( .A(n16537), .B(n16538), .Z(n16525) );
  AND U17562 ( .A(n16539), .B(n16540), .Z(n16538) );
  XNOR U17563 ( .A(n16541), .B(n16537), .Z(n16540) );
  XOR U17564 ( .A(n16542), .B(e_input[672]), .Z(n16533) );
  IV U17565 ( .A(n16531), .Z(n16542) );
  XOR U17566 ( .A(n16543), .B(n16544), .Z(n16531) );
  AND U17567 ( .A(n16545), .B(n16546), .Z(n16544) );
  XNOR U17568 ( .A(n16543), .B(n8274), .Z(n16546) );
  XNOR U17569 ( .A(n16539), .B(n16541), .Z(n8274) );
  NAND U17570 ( .A(n16547), .B(e_input[671]), .Z(n16541) );
  NAND U17571 ( .A(n12323), .B(e_input[671]), .Z(n16547) );
  XNOR U17572 ( .A(n16537), .B(n16548), .Z(n16539) );
  XOR U17573 ( .A(n16549), .B(n16550), .Z(n16537) );
  AND U17574 ( .A(n16551), .B(n16552), .Z(n16550) );
  XNOR U17575 ( .A(n16553), .B(n16549), .Z(n16552) );
  XOR U17576 ( .A(n16554), .B(e_input[671]), .Z(n16545) );
  IV U17577 ( .A(n16543), .Z(n16554) );
  XOR U17578 ( .A(n16555), .B(n16556), .Z(n16543) );
  AND U17579 ( .A(n16557), .B(n16558), .Z(n16556) );
  XNOR U17580 ( .A(n16555), .B(n8280), .Z(n16558) );
  XNOR U17581 ( .A(n16551), .B(n16553), .Z(n8280) );
  NAND U17582 ( .A(n16559), .B(e_input[670]), .Z(n16553) );
  NAND U17583 ( .A(n12323), .B(e_input[670]), .Z(n16559) );
  XNOR U17584 ( .A(n16549), .B(n16560), .Z(n16551) );
  XOR U17585 ( .A(n16561), .B(n16562), .Z(n16549) );
  AND U17586 ( .A(n16563), .B(n16564), .Z(n16562) );
  XNOR U17587 ( .A(n16565), .B(n16561), .Z(n16564) );
  XOR U17588 ( .A(n16566), .B(e_input[670]), .Z(n16557) );
  IV U17589 ( .A(n16555), .Z(n16566) );
  XOR U17590 ( .A(n16567), .B(n16568), .Z(n16555) );
  AND U17591 ( .A(n16569), .B(n16570), .Z(n16568) );
  XNOR U17592 ( .A(n16567), .B(n8286), .Z(n16570) );
  XNOR U17593 ( .A(n16563), .B(n16565), .Z(n8286) );
  NAND U17594 ( .A(n16571), .B(e_input[669]), .Z(n16565) );
  NAND U17595 ( .A(n12323), .B(e_input[669]), .Z(n16571) );
  XNOR U17596 ( .A(n16561), .B(n16572), .Z(n16563) );
  XOR U17597 ( .A(n16573), .B(n16574), .Z(n16561) );
  AND U17598 ( .A(n16575), .B(n16576), .Z(n16574) );
  XNOR U17599 ( .A(n16577), .B(n16573), .Z(n16576) );
  XOR U17600 ( .A(n16578), .B(e_input[669]), .Z(n16569) );
  IV U17601 ( .A(n16567), .Z(n16578) );
  XOR U17602 ( .A(n16579), .B(n16580), .Z(n16567) );
  AND U17603 ( .A(n16581), .B(n16582), .Z(n16580) );
  XNOR U17604 ( .A(n16579), .B(n8292), .Z(n16582) );
  XNOR U17605 ( .A(n16575), .B(n16577), .Z(n8292) );
  NAND U17606 ( .A(n16583), .B(e_input[668]), .Z(n16577) );
  NAND U17607 ( .A(n12323), .B(e_input[668]), .Z(n16583) );
  XNOR U17608 ( .A(n16573), .B(n16584), .Z(n16575) );
  XOR U17609 ( .A(n16585), .B(n16586), .Z(n16573) );
  AND U17610 ( .A(n16587), .B(n16588), .Z(n16586) );
  XNOR U17611 ( .A(n16589), .B(n16585), .Z(n16588) );
  XOR U17612 ( .A(n16590), .B(e_input[668]), .Z(n16581) );
  IV U17613 ( .A(n16579), .Z(n16590) );
  XOR U17614 ( .A(n16591), .B(n16592), .Z(n16579) );
  AND U17615 ( .A(n16593), .B(n16594), .Z(n16592) );
  XNOR U17616 ( .A(n16591), .B(n8298), .Z(n16594) );
  XNOR U17617 ( .A(n16587), .B(n16589), .Z(n8298) );
  NAND U17618 ( .A(n16595), .B(e_input[667]), .Z(n16589) );
  NAND U17619 ( .A(n12323), .B(e_input[667]), .Z(n16595) );
  XNOR U17620 ( .A(n16585), .B(n16596), .Z(n16587) );
  XOR U17621 ( .A(n16597), .B(n16598), .Z(n16585) );
  AND U17622 ( .A(n16599), .B(n16600), .Z(n16598) );
  XNOR U17623 ( .A(n16601), .B(n16597), .Z(n16600) );
  XOR U17624 ( .A(n16602), .B(e_input[667]), .Z(n16593) );
  IV U17625 ( .A(n16591), .Z(n16602) );
  XOR U17626 ( .A(n16603), .B(n16604), .Z(n16591) );
  AND U17627 ( .A(n16605), .B(n16606), .Z(n16604) );
  XNOR U17628 ( .A(n16603), .B(n8304), .Z(n16606) );
  XNOR U17629 ( .A(n16599), .B(n16601), .Z(n8304) );
  NAND U17630 ( .A(n16607), .B(e_input[666]), .Z(n16601) );
  NAND U17631 ( .A(n12323), .B(e_input[666]), .Z(n16607) );
  XNOR U17632 ( .A(n16597), .B(n16608), .Z(n16599) );
  XOR U17633 ( .A(n16609), .B(n16610), .Z(n16597) );
  AND U17634 ( .A(n16611), .B(n16612), .Z(n16610) );
  XNOR U17635 ( .A(n16613), .B(n16609), .Z(n16612) );
  XOR U17636 ( .A(n16614), .B(e_input[666]), .Z(n16605) );
  IV U17637 ( .A(n16603), .Z(n16614) );
  XOR U17638 ( .A(n16615), .B(n16616), .Z(n16603) );
  AND U17639 ( .A(n16617), .B(n16618), .Z(n16616) );
  XNOR U17640 ( .A(n16615), .B(n8310), .Z(n16618) );
  XNOR U17641 ( .A(n16611), .B(n16613), .Z(n8310) );
  NAND U17642 ( .A(n16619), .B(e_input[665]), .Z(n16613) );
  NAND U17643 ( .A(n12323), .B(e_input[665]), .Z(n16619) );
  XNOR U17644 ( .A(n16609), .B(n16620), .Z(n16611) );
  XOR U17645 ( .A(n16621), .B(n16622), .Z(n16609) );
  AND U17646 ( .A(n16623), .B(n16624), .Z(n16622) );
  XNOR U17647 ( .A(n16625), .B(n16621), .Z(n16624) );
  XOR U17648 ( .A(n16626), .B(e_input[665]), .Z(n16617) );
  IV U17649 ( .A(n16615), .Z(n16626) );
  XOR U17650 ( .A(n16627), .B(n16628), .Z(n16615) );
  AND U17651 ( .A(n16629), .B(n16630), .Z(n16628) );
  XNOR U17652 ( .A(n16627), .B(n8316), .Z(n16630) );
  XNOR U17653 ( .A(n16623), .B(n16625), .Z(n8316) );
  NAND U17654 ( .A(n16631), .B(e_input[664]), .Z(n16625) );
  NAND U17655 ( .A(n12323), .B(e_input[664]), .Z(n16631) );
  XNOR U17656 ( .A(n16621), .B(n16632), .Z(n16623) );
  XOR U17657 ( .A(n16633), .B(n16634), .Z(n16621) );
  AND U17658 ( .A(n16635), .B(n16636), .Z(n16634) );
  XNOR U17659 ( .A(n16637), .B(n16633), .Z(n16636) );
  XOR U17660 ( .A(n16638), .B(e_input[664]), .Z(n16629) );
  IV U17661 ( .A(n16627), .Z(n16638) );
  XOR U17662 ( .A(n16639), .B(n16640), .Z(n16627) );
  AND U17663 ( .A(n16641), .B(n16642), .Z(n16640) );
  XNOR U17664 ( .A(n16639), .B(n8322), .Z(n16642) );
  XNOR U17665 ( .A(n16635), .B(n16637), .Z(n8322) );
  NAND U17666 ( .A(n16643), .B(e_input[663]), .Z(n16637) );
  NAND U17667 ( .A(n12323), .B(e_input[663]), .Z(n16643) );
  XNOR U17668 ( .A(n16633), .B(n16644), .Z(n16635) );
  XOR U17669 ( .A(n16645), .B(n16646), .Z(n16633) );
  AND U17670 ( .A(n16647), .B(n16648), .Z(n16646) );
  XNOR U17671 ( .A(n16649), .B(n16645), .Z(n16648) );
  XOR U17672 ( .A(n16650), .B(e_input[663]), .Z(n16641) );
  IV U17673 ( .A(n16639), .Z(n16650) );
  XOR U17674 ( .A(n16651), .B(n16652), .Z(n16639) );
  AND U17675 ( .A(n16653), .B(n16654), .Z(n16652) );
  XNOR U17676 ( .A(n16651), .B(n8328), .Z(n16654) );
  XNOR U17677 ( .A(n16647), .B(n16649), .Z(n8328) );
  NAND U17678 ( .A(n16655), .B(e_input[662]), .Z(n16649) );
  NAND U17679 ( .A(n12323), .B(e_input[662]), .Z(n16655) );
  XNOR U17680 ( .A(n16645), .B(n16656), .Z(n16647) );
  XOR U17681 ( .A(n16657), .B(n16658), .Z(n16645) );
  AND U17682 ( .A(n16659), .B(n16660), .Z(n16658) );
  XNOR U17683 ( .A(n16661), .B(n16657), .Z(n16660) );
  XOR U17684 ( .A(n16662), .B(e_input[662]), .Z(n16653) );
  IV U17685 ( .A(n16651), .Z(n16662) );
  XOR U17686 ( .A(n16663), .B(n16664), .Z(n16651) );
  AND U17687 ( .A(n16665), .B(n16666), .Z(n16664) );
  XNOR U17688 ( .A(n16663), .B(n8334), .Z(n16666) );
  XNOR U17689 ( .A(n16659), .B(n16661), .Z(n8334) );
  NAND U17690 ( .A(n16667), .B(e_input[661]), .Z(n16661) );
  NAND U17691 ( .A(n12323), .B(e_input[661]), .Z(n16667) );
  XNOR U17692 ( .A(n16657), .B(n16668), .Z(n16659) );
  XOR U17693 ( .A(n16669), .B(n16670), .Z(n16657) );
  AND U17694 ( .A(n16671), .B(n16672), .Z(n16670) );
  XNOR U17695 ( .A(n16673), .B(n16669), .Z(n16672) );
  XOR U17696 ( .A(n16674), .B(e_input[661]), .Z(n16665) );
  IV U17697 ( .A(n16663), .Z(n16674) );
  XOR U17698 ( .A(n16675), .B(n16676), .Z(n16663) );
  AND U17699 ( .A(n16677), .B(n16678), .Z(n16676) );
  XNOR U17700 ( .A(n16675), .B(n8340), .Z(n16678) );
  XNOR U17701 ( .A(n16671), .B(n16673), .Z(n8340) );
  NAND U17702 ( .A(n16679), .B(e_input[660]), .Z(n16673) );
  NAND U17703 ( .A(n12323), .B(e_input[660]), .Z(n16679) );
  XNOR U17704 ( .A(n16669), .B(n16680), .Z(n16671) );
  XOR U17705 ( .A(n16681), .B(n16682), .Z(n16669) );
  AND U17706 ( .A(n16683), .B(n16684), .Z(n16682) );
  XNOR U17707 ( .A(n16685), .B(n16681), .Z(n16684) );
  XOR U17708 ( .A(n16686), .B(e_input[660]), .Z(n16677) );
  IV U17709 ( .A(n16675), .Z(n16686) );
  XOR U17710 ( .A(n16687), .B(n16688), .Z(n16675) );
  AND U17711 ( .A(n16689), .B(n16690), .Z(n16688) );
  XNOR U17712 ( .A(n16687), .B(n8346), .Z(n16690) );
  XNOR U17713 ( .A(n16683), .B(n16685), .Z(n8346) );
  NAND U17714 ( .A(n16691), .B(e_input[659]), .Z(n16685) );
  NAND U17715 ( .A(n12323), .B(e_input[659]), .Z(n16691) );
  XNOR U17716 ( .A(n16681), .B(n16692), .Z(n16683) );
  XOR U17717 ( .A(n16693), .B(n16694), .Z(n16681) );
  AND U17718 ( .A(n16695), .B(n16696), .Z(n16694) );
  XNOR U17719 ( .A(n16697), .B(n16693), .Z(n16696) );
  XOR U17720 ( .A(n16698), .B(e_input[659]), .Z(n16689) );
  IV U17721 ( .A(n16687), .Z(n16698) );
  XOR U17722 ( .A(n16699), .B(n16700), .Z(n16687) );
  AND U17723 ( .A(n16701), .B(n16702), .Z(n16700) );
  XNOR U17724 ( .A(n16699), .B(n8352), .Z(n16702) );
  XNOR U17725 ( .A(n16695), .B(n16697), .Z(n8352) );
  NAND U17726 ( .A(n16703), .B(e_input[658]), .Z(n16697) );
  NAND U17727 ( .A(n12323), .B(e_input[658]), .Z(n16703) );
  XNOR U17728 ( .A(n16693), .B(n16704), .Z(n16695) );
  XOR U17729 ( .A(n16705), .B(n16706), .Z(n16693) );
  AND U17730 ( .A(n16707), .B(n16708), .Z(n16706) );
  XNOR U17731 ( .A(n16709), .B(n16705), .Z(n16708) );
  XOR U17732 ( .A(n16710), .B(e_input[658]), .Z(n16701) );
  IV U17733 ( .A(n16699), .Z(n16710) );
  XOR U17734 ( .A(n16711), .B(n16712), .Z(n16699) );
  AND U17735 ( .A(n16713), .B(n16714), .Z(n16712) );
  XNOR U17736 ( .A(n16711), .B(n8358), .Z(n16714) );
  XNOR U17737 ( .A(n16707), .B(n16709), .Z(n8358) );
  NAND U17738 ( .A(n16715), .B(e_input[657]), .Z(n16709) );
  NAND U17739 ( .A(n12323), .B(e_input[657]), .Z(n16715) );
  XNOR U17740 ( .A(n16705), .B(n16716), .Z(n16707) );
  XOR U17741 ( .A(n16717), .B(n16718), .Z(n16705) );
  AND U17742 ( .A(n16719), .B(n16720), .Z(n16718) );
  XNOR U17743 ( .A(n16721), .B(n16717), .Z(n16720) );
  XOR U17744 ( .A(n16722), .B(e_input[657]), .Z(n16713) );
  IV U17745 ( .A(n16711), .Z(n16722) );
  XOR U17746 ( .A(n16723), .B(n16724), .Z(n16711) );
  AND U17747 ( .A(n16725), .B(n16726), .Z(n16724) );
  XNOR U17748 ( .A(n16723), .B(n8364), .Z(n16726) );
  XNOR U17749 ( .A(n16719), .B(n16721), .Z(n8364) );
  NAND U17750 ( .A(n16727), .B(e_input[656]), .Z(n16721) );
  NAND U17751 ( .A(n12323), .B(e_input[656]), .Z(n16727) );
  XNOR U17752 ( .A(n16717), .B(n16728), .Z(n16719) );
  XOR U17753 ( .A(n16729), .B(n16730), .Z(n16717) );
  AND U17754 ( .A(n16731), .B(n16732), .Z(n16730) );
  XNOR U17755 ( .A(n16733), .B(n16729), .Z(n16732) );
  XOR U17756 ( .A(n16734), .B(e_input[656]), .Z(n16725) );
  IV U17757 ( .A(n16723), .Z(n16734) );
  XOR U17758 ( .A(n16735), .B(n16736), .Z(n16723) );
  AND U17759 ( .A(n16737), .B(n16738), .Z(n16736) );
  XNOR U17760 ( .A(n16735), .B(n8370), .Z(n16738) );
  XNOR U17761 ( .A(n16731), .B(n16733), .Z(n8370) );
  NAND U17762 ( .A(n16739), .B(e_input[655]), .Z(n16733) );
  NAND U17763 ( .A(n12323), .B(e_input[655]), .Z(n16739) );
  XNOR U17764 ( .A(n16729), .B(n16740), .Z(n16731) );
  XOR U17765 ( .A(n16741), .B(n16742), .Z(n16729) );
  AND U17766 ( .A(n16743), .B(n16744), .Z(n16742) );
  XNOR U17767 ( .A(n16745), .B(n16741), .Z(n16744) );
  XOR U17768 ( .A(n16746), .B(e_input[655]), .Z(n16737) );
  IV U17769 ( .A(n16735), .Z(n16746) );
  XOR U17770 ( .A(n16747), .B(n16748), .Z(n16735) );
  AND U17771 ( .A(n16749), .B(n16750), .Z(n16748) );
  XNOR U17772 ( .A(n16747), .B(n8376), .Z(n16750) );
  XNOR U17773 ( .A(n16743), .B(n16745), .Z(n8376) );
  NAND U17774 ( .A(n16751), .B(e_input[654]), .Z(n16745) );
  NAND U17775 ( .A(n12323), .B(e_input[654]), .Z(n16751) );
  XNOR U17776 ( .A(n16741), .B(n16752), .Z(n16743) );
  XOR U17777 ( .A(n16753), .B(n16754), .Z(n16741) );
  AND U17778 ( .A(n16755), .B(n16756), .Z(n16754) );
  XNOR U17779 ( .A(n16757), .B(n16753), .Z(n16756) );
  XOR U17780 ( .A(n16758), .B(e_input[654]), .Z(n16749) );
  IV U17781 ( .A(n16747), .Z(n16758) );
  XOR U17782 ( .A(n16759), .B(n16760), .Z(n16747) );
  AND U17783 ( .A(n16761), .B(n16762), .Z(n16760) );
  XNOR U17784 ( .A(n16759), .B(n8382), .Z(n16762) );
  XNOR U17785 ( .A(n16755), .B(n16757), .Z(n8382) );
  NAND U17786 ( .A(n16763), .B(e_input[653]), .Z(n16757) );
  NAND U17787 ( .A(n12323), .B(e_input[653]), .Z(n16763) );
  XNOR U17788 ( .A(n16753), .B(n16764), .Z(n16755) );
  XOR U17789 ( .A(n16765), .B(n16766), .Z(n16753) );
  AND U17790 ( .A(n16767), .B(n16768), .Z(n16766) );
  XNOR U17791 ( .A(n16769), .B(n16765), .Z(n16768) );
  XOR U17792 ( .A(n16770), .B(e_input[653]), .Z(n16761) );
  IV U17793 ( .A(n16759), .Z(n16770) );
  XOR U17794 ( .A(n16771), .B(n16772), .Z(n16759) );
  AND U17795 ( .A(n16773), .B(n16774), .Z(n16772) );
  XNOR U17796 ( .A(n16771), .B(n8388), .Z(n16774) );
  XNOR U17797 ( .A(n16767), .B(n16769), .Z(n8388) );
  NAND U17798 ( .A(n16775), .B(e_input[652]), .Z(n16769) );
  NAND U17799 ( .A(n12323), .B(e_input[652]), .Z(n16775) );
  XNOR U17800 ( .A(n16765), .B(n16776), .Z(n16767) );
  XOR U17801 ( .A(n16777), .B(n16778), .Z(n16765) );
  AND U17802 ( .A(n16779), .B(n16780), .Z(n16778) );
  XNOR U17803 ( .A(n16781), .B(n16777), .Z(n16780) );
  XOR U17804 ( .A(n16782), .B(e_input[652]), .Z(n16773) );
  IV U17805 ( .A(n16771), .Z(n16782) );
  XOR U17806 ( .A(n16783), .B(n16784), .Z(n16771) );
  AND U17807 ( .A(n16785), .B(n16786), .Z(n16784) );
  XNOR U17808 ( .A(n16783), .B(n8394), .Z(n16786) );
  XNOR U17809 ( .A(n16779), .B(n16781), .Z(n8394) );
  NAND U17810 ( .A(n16787), .B(e_input[651]), .Z(n16781) );
  NAND U17811 ( .A(n12323), .B(e_input[651]), .Z(n16787) );
  XNOR U17812 ( .A(n16777), .B(n16788), .Z(n16779) );
  XOR U17813 ( .A(n16789), .B(n16790), .Z(n16777) );
  AND U17814 ( .A(n16791), .B(n16792), .Z(n16790) );
  XNOR U17815 ( .A(n16793), .B(n16789), .Z(n16792) );
  XOR U17816 ( .A(n16794), .B(e_input[651]), .Z(n16785) );
  IV U17817 ( .A(n16783), .Z(n16794) );
  XOR U17818 ( .A(n16795), .B(n16796), .Z(n16783) );
  AND U17819 ( .A(n16797), .B(n16798), .Z(n16796) );
  XNOR U17820 ( .A(n16795), .B(n8400), .Z(n16798) );
  XNOR U17821 ( .A(n16791), .B(n16793), .Z(n8400) );
  NAND U17822 ( .A(n16799), .B(e_input[650]), .Z(n16793) );
  NAND U17823 ( .A(n12323), .B(e_input[650]), .Z(n16799) );
  XNOR U17824 ( .A(n16789), .B(n16800), .Z(n16791) );
  XOR U17825 ( .A(n16801), .B(n16802), .Z(n16789) );
  AND U17826 ( .A(n16803), .B(n16804), .Z(n16802) );
  XNOR U17827 ( .A(n16805), .B(n16801), .Z(n16804) );
  XOR U17828 ( .A(n16806), .B(e_input[650]), .Z(n16797) );
  IV U17829 ( .A(n16795), .Z(n16806) );
  XOR U17830 ( .A(n16807), .B(n16808), .Z(n16795) );
  AND U17831 ( .A(n16809), .B(n16810), .Z(n16808) );
  XNOR U17832 ( .A(n16807), .B(n8406), .Z(n16810) );
  XNOR U17833 ( .A(n16803), .B(n16805), .Z(n8406) );
  NAND U17834 ( .A(n16811), .B(e_input[649]), .Z(n16805) );
  NAND U17835 ( .A(n12323), .B(e_input[649]), .Z(n16811) );
  XNOR U17836 ( .A(n16801), .B(n16812), .Z(n16803) );
  XOR U17837 ( .A(n16813), .B(n16814), .Z(n16801) );
  AND U17838 ( .A(n16815), .B(n16816), .Z(n16814) );
  XNOR U17839 ( .A(n16817), .B(n16813), .Z(n16816) );
  XOR U17840 ( .A(n16818), .B(e_input[649]), .Z(n16809) );
  IV U17841 ( .A(n16807), .Z(n16818) );
  XOR U17842 ( .A(n16819), .B(n16820), .Z(n16807) );
  AND U17843 ( .A(n16821), .B(n16822), .Z(n16820) );
  XNOR U17844 ( .A(n16819), .B(n8412), .Z(n16822) );
  XNOR U17845 ( .A(n16815), .B(n16817), .Z(n8412) );
  NAND U17846 ( .A(n16823), .B(e_input[648]), .Z(n16817) );
  NAND U17847 ( .A(n12323), .B(e_input[648]), .Z(n16823) );
  XNOR U17848 ( .A(n16813), .B(n16824), .Z(n16815) );
  XOR U17849 ( .A(n16825), .B(n16826), .Z(n16813) );
  AND U17850 ( .A(n16827), .B(n16828), .Z(n16826) );
  XNOR U17851 ( .A(n16829), .B(n16825), .Z(n16828) );
  XOR U17852 ( .A(n16830), .B(e_input[648]), .Z(n16821) );
  IV U17853 ( .A(n16819), .Z(n16830) );
  XOR U17854 ( .A(n16831), .B(n16832), .Z(n16819) );
  AND U17855 ( .A(n16833), .B(n16834), .Z(n16832) );
  XNOR U17856 ( .A(n16831), .B(n8418), .Z(n16834) );
  XNOR U17857 ( .A(n16827), .B(n16829), .Z(n8418) );
  NAND U17858 ( .A(n16835), .B(e_input[647]), .Z(n16829) );
  NAND U17859 ( .A(n12323), .B(e_input[647]), .Z(n16835) );
  XNOR U17860 ( .A(n16825), .B(n16836), .Z(n16827) );
  XOR U17861 ( .A(n16837), .B(n16838), .Z(n16825) );
  AND U17862 ( .A(n16839), .B(n16840), .Z(n16838) );
  XNOR U17863 ( .A(n16841), .B(n16837), .Z(n16840) );
  XOR U17864 ( .A(n16842), .B(e_input[647]), .Z(n16833) );
  IV U17865 ( .A(n16831), .Z(n16842) );
  XOR U17866 ( .A(n16843), .B(n16844), .Z(n16831) );
  AND U17867 ( .A(n16845), .B(n16846), .Z(n16844) );
  XNOR U17868 ( .A(n16843), .B(n8424), .Z(n16846) );
  XNOR U17869 ( .A(n16839), .B(n16841), .Z(n8424) );
  NAND U17870 ( .A(n16847), .B(e_input[646]), .Z(n16841) );
  NAND U17871 ( .A(n12323), .B(e_input[646]), .Z(n16847) );
  XNOR U17872 ( .A(n16837), .B(n16848), .Z(n16839) );
  XOR U17873 ( .A(n16849), .B(n16850), .Z(n16837) );
  AND U17874 ( .A(n16851), .B(n16852), .Z(n16850) );
  XNOR U17875 ( .A(n16853), .B(n16849), .Z(n16852) );
  XOR U17876 ( .A(n16854), .B(e_input[646]), .Z(n16845) );
  IV U17877 ( .A(n16843), .Z(n16854) );
  XOR U17878 ( .A(n16855), .B(n16856), .Z(n16843) );
  AND U17879 ( .A(n16857), .B(n16858), .Z(n16856) );
  XNOR U17880 ( .A(n16855), .B(n8430), .Z(n16858) );
  XNOR U17881 ( .A(n16851), .B(n16853), .Z(n8430) );
  NAND U17882 ( .A(n16859), .B(e_input[645]), .Z(n16853) );
  NAND U17883 ( .A(n12323), .B(e_input[645]), .Z(n16859) );
  XNOR U17884 ( .A(n16849), .B(n16860), .Z(n16851) );
  XOR U17885 ( .A(n16861), .B(n16862), .Z(n16849) );
  AND U17886 ( .A(n16863), .B(n16864), .Z(n16862) );
  XNOR U17887 ( .A(n16865), .B(n16861), .Z(n16864) );
  XOR U17888 ( .A(n16866), .B(e_input[645]), .Z(n16857) );
  IV U17889 ( .A(n16855), .Z(n16866) );
  XOR U17890 ( .A(n16867), .B(n16868), .Z(n16855) );
  AND U17891 ( .A(n16869), .B(n16870), .Z(n16868) );
  XNOR U17892 ( .A(n16867), .B(n8436), .Z(n16870) );
  XNOR U17893 ( .A(n16863), .B(n16865), .Z(n8436) );
  NAND U17894 ( .A(n16871), .B(e_input[644]), .Z(n16865) );
  NAND U17895 ( .A(n12323), .B(e_input[644]), .Z(n16871) );
  XNOR U17896 ( .A(n16861), .B(n16872), .Z(n16863) );
  XOR U17897 ( .A(n16873), .B(n16874), .Z(n16861) );
  AND U17898 ( .A(n16875), .B(n16876), .Z(n16874) );
  XNOR U17899 ( .A(n16877), .B(n16873), .Z(n16876) );
  XOR U17900 ( .A(n16878), .B(e_input[644]), .Z(n16869) );
  IV U17901 ( .A(n16867), .Z(n16878) );
  XOR U17902 ( .A(n16879), .B(n16880), .Z(n16867) );
  AND U17903 ( .A(n16881), .B(n16882), .Z(n16880) );
  XNOR U17904 ( .A(n16879), .B(n8442), .Z(n16882) );
  XNOR U17905 ( .A(n16875), .B(n16877), .Z(n8442) );
  NAND U17906 ( .A(n16883), .B(e_input[643]), .Z(n16877) );
  NAND U17907 ( .A(n12323), .B(e_input[643]), .Z(n16883) );
  XNOR U17908 ( .A(n16873), .B(n16884), .Z(n16875) );
  XOR U17909 ( .A(n16885), .B(n16886), .Z(n16873) );
  AND U17910 ( .A(n16887), .B(n16888), .Z(n16886) );
  XNOR U17911 ( .A(n16889), .B(n16885), .Z(n16888) );
  XOR U17912 ( .A(n16890), .B(e_input[643]), .Z(n16881) );
  IV U17913 ( .A(n16879), .Z(n16890) );
  XOR U17914 ( .A(n16891), .B(n16892), .Z(n16879) );
  AND U17915 ( .A(n16893), .B(n16894), .Z(n16892) );
  XNOR U17916 ( .A(n16891), .B(n8448), .Z(n16894) );
  XNOR U17917 ( .A(n16887), .B(n16889), .Z(n8448) );
  NAND U17918 ( .A(n16895), .B(e_input[642]), .Z(n16889) );
  NAND U17919 ( .A(n12323), .B(e_input[642]), .Z(n16895) );
  XNOR U17920 ( .A(n16885), .B(n16896), .Z(n16887) );
  XOR U17921 ( .A(n16897), .B(n16898), .Z(n16885) );
  AND U17922 ( .A(n16899), .B(n16900), .Z(n16898) );
  XNOR U17923 ( .A(n16901), .B(n16897), .Z(n16900) );
  XOR U17924 ( .A(n16902), .B(e_input[642]), .Z(n16893) );
  IV U17925 ( .A(n16891), .Z(n16902) );
  XOR U17926 ( .A(n16903), .B(n16904), .Z(n16891) );
  AND U17927 ( .A(n16905), .B(n16906), .Z(n16904) );
  XNOR U17928 ( .A(n16903), .B(n8454), .Z(n16906) );
  XNOR U17929 ( .A(n16899), .B(n16901), .Z(n8454) );
  NAND U17930 ( .A(n16907), .B(e_input[641]), .Z(n16901) );
  NAND U17931 ( .A(n12323), .B(e_input[641]), .Z(n16907) );
  XNOR U17932 ( .A(n16897), .B(n16908), .Z(n16899) );
  XOR U17933 ( .A(n16909), .B(n16910), .Z(n16897) );
  AND U17934 ( .A(n16911), .B(n16912), .Z(n16910) );
  XNOR U17935 ( .A(n16913), .B(n16909), .Z(n16912) );
  XOR U17936 ( .A(n16914), .B(e_input[641]), .Z(n16905) );
  IV U17937 ( .A(n16903), .Z(n16914) );
  XOR U17938 ( .A(n16915), .B(n16916), .Z(n16903) );
  AND U17939 ( .A(n16917), .B(n16918), .Z(n16916) );
  XNOR U17940 ( .A(n16915), .B(n8460), .Z(n16918) );
  XNOR U17941 ( .A(n16911), .B(n16913), .Z(n8460) );
  NAND U17942 ( .A(n16919), .B(e_input[640]), .Z(n16913) );
  NAND U17943 ( .A(n12323), .B(e_input[640]), .Z(n16919) );
  XNOR U17944 ( .A(n16909), .B(n16920), .Z(n16911) );
  XOR U17945 ( .A(n16921), .B(n16922), .Z(n16909) );
  AND U17946 ( .A(n16923), .B(n16924), .Z(n16922) );
  XNOR U17947 ( .A(n16925), .B(n16921), .Z(n16924) );
  XOR U17948 ( .A(n16926), .B(e_input[640]), .Z(n16917) );
  IV U17949 ( .A(n16915), .Z(n16926) );
  XOR U17950 ( .A(n16927), .B(n16928), .Z(n16915) );
  AND U17951 ( .A(n16929), .B(n16930), .Z(n16928) );
  XNOR U17952 ( .A(n16927), .B(n8466), .Z(n16930) );
  XNOR U17953 ( .A(n16923), .B(n16925), .Z(n8466) );
  NAND U17954 ( .A(n16931), .B(e_input[639]), .Z(n16925) );
  NAND U17955 ( .A(n12323), .B(e_input[639]), .Z(n16931) );
  XNOR U17956 ( .A(n16921), .B(n16932), .Z(n16923) );
  XOR U17957 ( .A(n16933), .B(n16934), .Z(n16921) );
  AND U17958 ( .A(n16935), .B(n16936), .Z(n16934) );
  XNOR U17959 ( .A(n16937), .B(n16933), .Z(n16936) );
  XOR U17960 ( .A(n16938), .B(e_input[639]), .Z(n16929) );
  IV U17961 ( .A(n16927), .Z(n16938) );
  XOR U17962 ( .A(n16939), .B(n16940), .Z(n16927) );
  AND U17963 ( .A(n16941), .B(n16942), .Z(n16940) );
  XNOR U17964 ( .A(n16939), .B(n8472), .Z(n16942) );
  XNOR U17965 ( .A(n16935), .B(n16937), .Z(n8472) );
  NAND U17966 ( .A(n16943), .B(e_input[638]), .Z(n16937) );
  NAND U17967 ( .A(n12323), .B(e_input[638]), .Z(n16943) );
  XNOR U17968 ( .A(n16933), .B(n16944), .Z(n16935) );
  XOR U17969 ( .A(n16945), .B(n16946), .Z(n16933) );
  AND U17970 ( .A(n16947), .B(n16948), .Z(n16946) );
  XNOR U17971 ( .A(n16949), .B(n16945), .Z(n16948) );
  XOR U17972 ( .A(n16950), .B(e_input[638]), .Z(n16941) );
  IV U17973 ( .A(n16939), .Z(n16950) );
  XOR U17974 ( .A(n16951), .B(n16952), .Z(n16939) );
  AND U17975 ( .A(n16953), .B(n16954), .Z(n16952) );
  XNOR U17976 ( .A(n16951), .B(n8478), .Z(n16954) );
  XNOR U17977 ( .A(n16947), .B(n16949), .Z(n8478) );
  NAND U17978 ( .A(n16955), .B(e_input[637]), .Z(n16949) );
  NAND U17979 ( .A(n12323), .B(e_input[637]), .Z(n16955) );
  XNOR U17980 ( .A(n16945), .B(n16956), .Z(n16947) );
  XOR U17981 ( .A(n16957), .B(n16958), .Z(n16945) );
  AND U17982 ( .A(n16959), .B(n16960), .Z(n16958) );
  XNOR U17983 ( .A(n16961), .B(n16957), .Z(n16960) );
  XOR U17984 ( .A(n16962), .B(e_input[637]), .Z(n16953) );
  IV U17985 ( .A(n16951), .Z(n16962) );
  XOR U17986 ( .A(n16963), .B(n16964), .Z(n16951) );
  AND U17987 ( .A(n16965), .B(n16966), .Z(n16964) );
  XNOR U17988 ( .A(n16963), .B(n8484), .Z(n16966) );
  XNOR U17989 ( .A(n16959), .B(n16961), .Z(n8484) );
  NAND U17990 ( .A(n16967), .B(e_input[636]), .Z(n16961) );
  NAND U17991 ( .A(n12323), .B(e_input[636]), .Z(n16967) );
  XNOR U17992 ( .A(n16957), .B(n16968), .Z(n16959) );
  XOR U17993 ( .A(n16969), .B(n16970), .Z(n16957) );
  AND U17994 ( .A(n16971), .B(n16972), .Z(n16970) );
  XNOR U17995 ( .A(n16973), .B(n16969), .Z(n16972) );
  XOR U17996 ( .A(n16974), .B(e_input[636]), .Z(n16965) );
  IV U17997 ( .A(n16963), .Z(n16974) );
  XOR U17998 ( .A(n16975), .B(n16976), .Z(n16963) );
  AND U17999 ( .A(n16977), .B(n16978), .Z(n16976) );
  XNOR U18000 ( .A(n16975), .B(n8490), .Z(n16978) );
  XNOR U18001 ( .A(n16971), .B(n16973), .Z(n8490) );
  NAND U18002 ( .A(n16979), .B(e_input[635]), .Z(n16973) );
  NAND U18003 ( .A(n12323), .B(e_input[635]), .Z(n16979) );
  XNOR U18004 ( .A(n16969), .B(n16980), .Z(n16971) );
  XOR U18005 ( .A(n16981), .B(n16982), .Z(n16969) );
  AND U18006 ( .A(n16983), .B(n16984), .Z(n16982) );
  XNOR U18007 ( .A(n16985), .B(n16981), .Z(n16984) );
  XOR U18008 ( .A(n16986), .B(e_input[635]), .Z(n16977) );
  IV U18009 ( .A(n16975), .Z(n16986) );
  XOR U18010 ( .A(n16987), .B(n16988), .Z(n16975) );
  AND U18011 ( .A(n16989), .B(n16990), .Z(n16988) );
  XNOR U18012 ( .A(n16987), .B(n8496), .Z(n16990) );
  XNOR U18013 ( .A(n16983), .B(n16985), .Z(n8496) );
  NAND U18014 ( .A(n16991), .B(e_input[634]), .Z(n16985) );
  NAND U18015 ( .A(n12323), .B(e_input[634]), .Z(n16991) );
  XNOR U18016 ( .A(n16981), .B(n16992), .Z(n16983) );
  XOR U18017 ( .A(n16993), .B(n16994), .Z(n16981) );
  AND U18018 ( .A(n16995), .B(n16996), .Z(n16994) );
  XNOR U18019 ( .A(n16997), .B(n16993), .Z(n16996) );
  XOR U18020 ( .A(n16998), .B(e_input[634]), .Z(n16989) );
  IV U18021 ( .A(n16987), .Z(n16998) );
  XOR U18022 ( .A(n16999), .B(n17000), .Z(n16987) );
  AND U18023 ( .A(n17001), .B(n17002), .Z(n17000) );
  XNOR U18024 ( .A(n16999), .B(n8502), .Z(n17002) );
  XNOR U18025 ( .A(n16995), .B(n16997), .Z(n8502) );
  NAND U18026 ( .A(n17003), .B(e_input[633]), .Z(n16997) );
  NAND U18027 ( .A(n12323), .B(e_input[633]), .Z(n17003) );
  XNOR U18028 ( .A(n16993), .B(n17004), .Z(n16995) );
  XOR U18029 ( .A(n17005), .B(n17006), .Z(n16993) );
  AND U18030 ( .A(n17007), .B(n17008), .Z(n17006) );
  XNOR U18031 ( .A(n17009), .B(n17005), .Z(n17008) );
  XOR U18032 ( .A(n17010), .B(e_input[633]), .Z(n17001) );
  IV U18033 ( .A(n16999), .Z(n17010) );
  XOR U18034 ( .A(n17011), .B(n17012), .Z(n16999) );
  AND U18035 ( .A(n17013), .B(n17014), .Z(n17012) );
  XNOR U18036 ( .A(n17011), .B(n8508), .Z(n17014) );
  XNOR U18037 ( .A(n17007), .B(n17009), .Z(n8508) );
  NAND U18038 ( .A(n17015), .B(e_input[632]), .Z(n17009) );
  NAND U18039 ( .A(n12323), .B(e_input[632]), .Z(n17015) );
  XNOR U18040 ( .A(n17005), .B(n17016), .Z(n17007) );
  XOR U18041 ( .A(n17017), .B(n17018), .Z(n17005) );
  AND U18042 ( .A(n17019), .B(n17020), .Z(n17018) );
  XNOR U18043 ( .A(n17021), .B(n17017), .Z(n17020) );
  XOR U18044 ( .A(n17022), .B(e_input[632]), .Z(n17013) );
  IV U18045 ( .A(n17011), .Z(n17022) );
  XOR U18046 ( .A(n17023), .B(n17024), .Z(n17011) );
  AND U18047 ( .A(n17025), .B(n17026), .Z(n17024) );
  XNOR U18048 ( .A(n17023), .B(n8514), .Z(n17026) );
  XNOR U18049 ( .A(n17019), .B(n17021), .Z(n8514) );
  NAND U18050 ( .A(n17027), .B(e_input[631]), .Z(n17021) );
  NAND U18051 ( .A(n12323), .B(e_input[631]), .Z(n17027) );
  XNOR U18052 ( .A(n17017), .B(n17028), .Z(n17019) );
  XOR U18053 ( .A(n17029), .B(n17030), .Z(n17017) );
  AND U18054 ( .A(n17031), .B(n17032), .Z(n17030) );
  XNOR U18055 ( .A(n17033), .B(n17029), .Z(n17032) );
  XOR U18056 ( .A(n17034), .B(e_input[631]), .Z(n17025) );
  IV U18057 ( .A(n17023), .Z(n17034) );
  XOR U18058 ( .A(n17035), .B(n17036), .Z(n17023) );
  AND U18059 ( .A(n17037), .B(n17038), .Z(n17036) );
  XNOR U18060 ( .A(n17035), .B(n8520), .Z(n17038) );
  XNOR U18061 ( .A(n17031), .B(n17033), .Z(n8520) );
  NAND U18062 ( .A(n17039), .B(e_input[630]), .Z(n17033) );
  NAND U18063 ( .A(n12323), .B(e_input[630]), .Z(n17039) );
  XNOR U18064 ( .A(n17029), .B(n17040), .Z(n17031) );
  XOR U18065 ( .A(n17041), .B(n17042), .Z(n17029) );
  AND U18066 ( .A(n17043), .B(n17044), .Z(n17042) );
  XNOR U18067 ( .A(n17045), .B(n17041), .Z(n17044) );
  XOR U18068 ( .A(n17046), .B(e_input[630]), .Z(n17037) );
  IV U18069 ( .A(n17035), .Z(n17046) );
  XOR U18070 ( .A(n17047), .B(n17048), .Z(n17035) );
  AND U18071 ( .A(n17049), .B(n17050), .Z(n17048) );
  XNOR U18072 ( .A(n17047), .B(n8526), .Z(n17050) );
  XNOR U18073 ( .A(n17043), .B(n17045), .Z(n8526) );
  NAND U18074 ( .A(n17051), .B(e_input[629]), .Z(n17045) );
  NAND U18075 ( .A(n12323), .B(e_input[629]), .Z(n17051) );
  XNOR U18076 ( .A(n17041), .B(n17052), .Z(n17043) );
  XOR U18077 ( .A(n17053), .B(n17054), .Z(n17041) );
  AND U18078 ( .A(n17055), .B(n17056), .Z(n17054) );
  XNOR U18079 ( .A(n17057), .B(n17053), .Z(n17056) );
  XOR U18080 ( .A(n17058), .B(e_input[629]), .Z(n17049) );
  IV U18081 ( .A(n17047), .Z(n17058) );
  XOR U18082 ( .A(n17059), .B(n17060), .Z(n17047) );
  AND U18083 ( .A(n17061), .B(n17062), .Z(n17060) );
  XNOR U18084 ( .A(n17059), .B(n8532), .Z(n17062) );
  XNOR U18085 ( .A(n17055), .B(n17057), .Z(n8532) );
  NAND U18086 ( .A(n17063), .B(e_input[628]), .Z(n17057) );
  NAND U18087 ( .A(n12323), .B(e_input[628]), .Z(n17063) );
  XNOR U18088 ( .A(n17053), .B(n17064), .Z(n17055) );
  XOR U18089 ( .A(n17065), .B(n17066), .Z(n17053) );
  AND U18090 ( .A(n17067), .B(n17068), .Z(n17066) );
  XNOR U18091 ( .A(n17069), .B(n17065), .Z(n17068) );
  XOR U18092 ( .A(n17070), .B(e_input[628]), .Z(n17061) );
  IV U18093 ( .A(n17059), .Z(n17070) );
  XOR U18094 ( .A(n17071), .B(n17072), .Z(n17059) );
  AND U18095 ( .A(n17073), .B(n17074), .Z(n17072) );
  XNOR U18096 ( .A(n17071), .B(n8538), .Z(n17074) );
  XNOR U18097 ( .A(n17067), .B(n17069), .Z(n8538) );
  NAND U18098 ( .A(n17075), .B(e_input[627]), .Z(n17069) );
  NAND U18099 ( .A(n12323), .B(e_input[627]), .Z(n17075) );
  XNOR U18100 ( .A(n17065), .B(n17076), .Z(n17067) );
  XOR U18101 ( .A(n17077), .B(n17078), .Z(n17065) );
  AND U18102 ( .A(n17079), .B(n17080), .Z(n17078) );
  XNOR U18103 ( .A(n17081), .B(n17077), .Z(n17080) );
  XOR U18104 ( .A(n17082), .B(e_input[627]), .Z(n17073) );
  IV U18105 ( .A(n17071), .Z(n17082) );
  XOR U18106 ( .A(n17083), .B(n17084), .Z(n17071) );
  AND U18107 ( .A(n17085), .B(n17086), .Z(n17084) );
  XNOR U18108 ( .A(n17083), .B(n8544), .Z(n17086) );
  XNOR U18109 ( .A(n17079), .B(n17081), .Z(n8544) );
  NAND U18110 ( .A(n17087), .B(e_input[626]), .Z(n17081) );
  NAND U18111 ( .A(n12323), .B(e_input[626]), .Z(n17087) );
  XNOR U18112 ( .A(n17077), .B(n17088), .Z(n17079) );
  XOR U18113 ( .A(n17089), .B(n17090), .Z(n17077) );
  AND U18114 ( .A(n17091), .B(n17092), .Z(n17090) );
  XNOR U18115 ( .A(n17093), .B(n17089), .Z(n17092) );
  XOR U18116 ( .A(n17094), .B(e_input[626]), .Z(n17085) );
  IV U18117 ( .A(n17083), .Z(n17094) );
  XOR U18118 ( .A(n17095), .B(n17096), .Z(n17083) );
  AND U18119 ( .A(n17097), .B(n17098), .Z(n17096) );
  XNOR U18120 ( .A(n17095), .B(n8550), .Z(n17098) );
  XNOR U18121 ( .A(n17091), .B(n17093), .Z(n8550) );
  NAND U18122 ( .A(n17099), .B(e_input[625]), .Z(n17093) );
  NAND U18123 ( .A(n12323), .B(e_input[625]), .Z(n17099) );
  XNOR U18124 ( .A(n17089), .B(n17100), .Z(n17091) );
  XOR U18125 ( .A(n17101), .B(n17102), .Z(n17089) );
  AND U18126 ( .A(n17103), .B(n17104), .Z(n17102) );
  XNOR U18127 ( .A(n17105), .B(n17101), .Z(n17104) );
  XOR U18128 ( .A(n17106), .B(e_input[625]), .Z(n17097) );
  IV U18129 ( .A(n17095), .Z(n17106) );
  XOR U18130 ( .A(n17107), .B(n17108), .Z(n17095) );
  AND U18131 ( .A(n17109), .B(n17110), .Z(n17108) );
  XNOR U18132 ( .A(n17107), .B(n8556), .Z(n17110) );
  XNOR U18133 ( .A(n17103), .B(n17105), .Z(n8556) );
  NAND U18134 ( .A(n17111), .B(e_input[624]), .Z(n17105) );
  NAND U18135 ( .A(n12323), .B(e_input[624]), .Z(n17111) );
  XNOR U18136 ( .A(n17101), .B(n17112), .Z(n17103) );
  XOR U18137 ( .A(n17113), .B(n17114), .Z(n17101) );
  AND U18138 ( .A(n17115), .B(n17116), .Z(n17114) );
  XNOR U18139 ( .A(n17117), .B(n17113), .Z(n17116) );
  XOR U18140 ( .A(n17118), .B(e_input[624]), .Z(n17109) );
  IV U18141 ( .A(n17107), .Z(n17118) );
  XOR U18142 ( .A(n17119), .B(n17120), .Z(n17107) );
  AND U18143 ( .A(n17121), .B(n17122), .Z(n17120) );
  XNOR U18144 ( .A(n17119), .B(n8562), .Z(n17122) );
  XNOR U18145 ( .A(n17115), .B(n17117), .Z(n8562) );
  NAND U18146 ( .A(n17123), .B(e_input[623]), .Z(n17117) );
  NAND U18147 ( .A(n12323), .B(e_input[623]), .Z(n17123) );
  XNOR U18148 ( .A(n17113), .B(n17124), .Z(n17115) );
  XOR U18149 ( .A(n17125), .B(n17126), .Z(n17113) );
  AND U18150 ( .A(n17127), .B(n17128), .Z(n17126) );
  XNOR U18151 ( .A(n17129), .B(n17125), .Z(n17128) );
  XOR U18152 ( .A(n17130), .B(e_input[623]), .Z(n17121) );
  IV U18153 ( .A(n17119), .Z(n17130) );
  XOR U18154 ( .A(n17131), .B(n17132), .Z(n17119) );
  AND U18155 ( .A(n17133), .B(n17134), .Z(n17132) );
  XNOR U18156 ( .A(n17131), .B(n8568), .Z(n17134) );
  XNOR U18157 ( .A(n17127), .B(n17129), .Z(n8568) );
  NAND U18158 ( .A(n17135), .B(e_input[622]), .Z(n17129) );
  NAND U18159 ( .A(n12323), .B(e_input[622]), .Z(n17135) );
  XNOR U18160 ( .A(n17125), .B(n17136), .Z(n17127) );
  XOR U18161 ( .A(n17137), .B(n17138), .Z(n17125) );
  AND U18162 ( .A(n17139), .B(n17140), .Z(n17138) );
  XNOR U18163 ( .A(n17141), .B(n17137), .Z(n17140) );
  XOR U18164 ( .A(n17142), .B(e_input[622]), .Z(n17133) );
  IV U18165 ( .A(n17131), .Z(n17142) );
  XOR U18166 ( .A(n17143), .B(n17144), .Z(n17131) );
  AND U18167 ( .A(n17145), .B(n17146), .Z(n17144) );
  XNOR U18168 ( .A(n17143), .B(n8574), .Z(n17146) );
  XNOR U18169 ( .A(n17139), .B(n17141), .Z(n8574) );
  NAND U18170 ( .A(n17147), .B(e_input[621]), .Z(n17141) );
  NAND U18171 ( .A(n12323), .B(e_input[621]), .Z(n17147) );
  XNOR U18172 ( .A(n17137), .B(n17148), .Z(n17139) );
  XOR U18173 ( .A(n17149), .B(n17150), .Z(n17137) );
  AND U18174 ( .A(n17151), .B(n17152), .Z(n17150) );
  XNOR U18175 ( .A(n17153), .B(n17149), .Z(n17152) );
  XOR U18176 ( .A(n17154), .B(e_input[621]), .Z(n17145) );
  IV U18177 ( .A(n17143), .Z(n17154) );
  XOR U18178 ( .A(n17155), .B(n17156), .Z(n17143) );
  AND U18179 ( .A(n17157), .B(n17158), .Z(n17156) );
  XNOR U18180 ( .A(n17155), .B(n8580), .Z(n17158) );
  XNOR U18181 ( .A(n17151), .B(n17153), .Z(n8580) );
  NAND U18182 ( .A(n17159), .B(e_input[620]), .Z(n17153) );
  NAND U18183 ( .A(n12323), .B(e_input[620]), .Z(n17159) );
  XNOR U18184 ( .A(n17149), .B(n17160), .Z(n17151) );
  XOR U18185 ( .A(n17161), .B(n17162), .Z(n17149) );
  AND U18186 ( .A(n17163), .B(n17164), .Z(n17162) );
  XNOR U18187 ( .A(n17165), .B(n17161), .Z(n17164) );
  XOR U18188 ( .A(n17166), .B(e_input[620]), .Z(n17157) );
  IV U18189 ( .A(n17155), .Z(n17166) );
  XOR U18190 ( .A(n17167), .B(n17168), .Z(n17155) );
  AND U18191 ( .A(n17169), .B(n17170), .Z(n17168) );
  XNOR U18192 ( .A(n17167), .B(n8586), .Z(n17170) );
  XNOR U18193 ( .A(n17163), .B(n17165), .Z(n8586) );
  NAND U18194 ( .A(n17171), .B(e_input[619]), .Z(n17165) );
  NAND U18195 ( .A(n12323), .B(e_input[619]), .Z(n17171) );
  XNOR U18196 ( .A(n17161), .B(n17172), .Z(n17163) );
  XOR U18197 ( .A(n17173), .B(n17174), .Z(n17161) );
  AND U18198 ( .A(n17175), .B(n17176), .Z(n17174) );
  XNOR U18199 ( .A(n17177), .B(n17173), .Z(n17176) );
  XOR U18200 ( .A(n17178), .B(e_input[619]), .Z(n17169) );
  IV U18201 ( .A(n17167), .Z(n17178) );
  XOR U18202 ( .A(n17179), .B(n17180), .Z(n17167) );
  AND U18203 ( .A(n17181), .B(n17182), .Z(n17180) );
  XNOR U18204 ( .A(n17179), .B(n8592), .Z(n17182) );
  XNOR U18205 ( .A(n17175), .B(n17177), .Z(n8592) );
  NAND U18206 ( .A(n17183), .B(e_input[618]), .Z(n17177) );
  NAND U18207 ( .A(n12323), .B(e_input[618]), .Z(n17183) );
  XNOR U18208 ( .A(n17173), .B(n17184), .Z(n17175) );
  XOR U18209 ( .A(n17185), .B(n17186), .Z(n17173) );
  AND U18210 ( .A(n17187), .B(n17188), .Z(n17186) );
  XNOR U18211 ( .A(n17189), .B(n17185), .Z(n17188) );
  XOR U18212 ( .A(n17190), .B(e_input[618]), .Z(n17181) );
  IV U18213 ( .A(n17179), .Z(n17190) );
  XOR U18214 ( .A(n17191), .B(n17192), .Z(n17179) );
  AND U18215 ( .A(n17193), .B(n17194), .Z(n17192) );
  XNOR U18216 ( .A(n17191), .B(n8598), .Z(n17194) );
  XNOR U18217 ( .A(n17187), .B(n17189), .Z(n8598) );
  NAND U18218 ( .A(n17195), .B(e_input[617]), .Z(n17189) );
  NAND U18219 ( .A(n12323), .B(e_input[617]), .Z(n17195) );
  XNOR U18220 ( .A(n17185), .B(n17196), .Z(n17187) );
  XOR U18221 ( .A(n17197), .B(n17198), .Z(n17185) );
  AND U18222 ( .A(n17199), .B(n17200), .Z(n17198) );
  XNOR U18223 ( .A(n17201), .B(n17197), .Z(n17200) );
  XOR U18224 ( .A(n17202), .B(e_input[617]), .Z(n17193) );
  IV U18225 ( .A(n17191), .Z(n17202) );
  XOR U18226 ( .A(n17203), .B(n17204), .Z(n17191) );
  AND U18227 ( .A(n17205), .B(n17206), .Z(n17204) );
  XNOR U18228 ( .A(n17203), .B(n8604), .Z(n17206) );
  XNOR U18229 ( .A(n17199), .B(n17201), .Z(n8604) );
  NAND U18230 ( .A(n17207), .B(e_input[616]), .Z(n17201) );
  NAND U18231 ( .A(n12323), .B(e_input[616]), .Z(n17207) );
  XNOR U18232 ( .A(n17197), .B(n17208), .Z(n17199) );
  XOR U18233 ( .A(n17209), .B(n17210), .Z(n17197) );
  AND U18234 ( .A(n17211), .B(n17212), .Z(n17210) );
  XNOR U18235 ( .A(n17213), .B(n17209), .Z(n17212) );
  XOR U18236 ( .A(n17214), .B(e_input[616]), .Z(n17205) );
  IV U18237 ( .A(n17203), .Z(n17214) );
  XOR U18238 ( .A(n17215), .B(n17216), .Z(n17203) );
  AND U18239 ( .A(n17217), .B(n17218), .Z(n17216) );
  XNOR U18240 ( .A(n17215), .B(n8610), .Z(n17218) );
  XNOR U18241 ( .A(n17211), .B(n17213), .Z(n8610) );
  NAND U18242 ( .A(n17219), .B(e_input[615]), .Z(n17213) );
  NAND U18243 ( .A(n12323), .B(e_input[615]), .Z(n17219) );
  XNOR U18244 ( .A(n17209), .B(n17220), .Z(n17211) );
  XOR U18245 ( .A(n17221), .B(n17222), .Z(n17209) );
  AND U18246 ( .A(n17223), .B(n17224), .Z(n17222) );
  XNOR U18247 ( .A(n17225), .B(n17221), .Z(n17224) );
  XOR U18248 ( .A(n17226), .B(e_input[615]), .Z(n17217) );
  IV U18249 ( .A(n17215), .Z(n17226) );
  XOR U18250 ( .A(n17227), .B(n17228), .Z(n17215) );
  AND U18251 ( .A(n17229), .B(n17230), .Z(n17228) );
  XNOR U18252 ( .A(n17227), .B(n8616), .Z(n17230) );
  XNOR U18253 ( .A(n17223), .B(n17225), .Z(n8616) );
  NAND U18254 ( .A(n17231), .B(e_input[614]), .Z(n17225) );
  NAND U18255 ( .A(n12323), .B(e_input[614]), .Z(n17231) );
  XNOR U18256 ( .A(n17221), .B(n17232), .Z(n17223) );
  XOR U18257 ( .A(n17233), .B(n17234), .Z(n17221) );
  AND U18258 ( .A(n17235), .B(n17236), .Z(n17234) );
  XNOR U18259 ( .A(n17237), .B(n17233), .Z(n17236) );
  XOR U18260 ( .A(n17238), .B(e_input[614]), .Z(n17229) );
  IV U18261 ( .A(n17227), .Z(n17238) );
  XOR U18262 ( .A(n17239), .B(n17240), .Z(n17227) );
  AND U18263 ( .A(n17241), .B(n17242), .Z(n17240) );
  XNOR U18264 ( .A(n17239), .B(n8622), .Z(n17242) );
  XNOR U18265 ( .A(n17235), .B(n17237), .Z(n8622) );
  NAND U18266 ( .A(n17243), .B(e_input[613]), .Z(n17237) );
  NAND U18267 ( .A(n12323), .B(e_input[613]), .Z(n17243) );
  XNOR U18268 ( .A(n17233), .B(n17244), .Z(n17235) );
  XOR U18269 ( .A(n17245), .B(n17246), .Z(n17233) );
  AND U18270 ( .A(n17247), .B(n17248), .Z(n17246) );
  XNOR U18271 ( .A(n17249), .B(n17245), .Z(n17248) );
  XOR U18272 ( .A(n17250), .B(e_input[613]), .Z(n17241) );
  IV U18273 ( .A(n17239), .Z(n17250) );
  XOR U18274 ( .A(n17251), .B(n17252), .Z(n17239) );
  AND U18275 ( .A(n17253), .B(n17254), .Z(n17252) );
  XNOR U18276 ( .A(n17251), .B(n8628), .Z(n17254) );
  XNOR U18277 ( .A(n17247), .B(n17249), .Z(n8628) );
  NAND U18278 ( .A(n17255), .B(e_input[612]), .Z(n17249) );
  NAND U18279 ( .A(n12323), .B(e_input[612]), .Z(n17255) );
  XNOR U18280 ( .A(n17245), .B(n17256), .Z(n17247) );
  XOR U18281 ( .A(n17257), .B(n17258), .Z(n17245) );
  AND U18282 ( .A(n17259), .B(n17260), .Z(n17258) );
  XNOR U18283 ( .A(n17261), .B(n17257), .Z(n17260) );
  XOR U18284 ( .A(n17262), .B(e_input[612]), .Z(n17253) );
  IV U18285 ( .A(n17251), .Z(n17262) );
  XOR U18286 ( .A(n17263), .B(n17264), .Z(n17251) );
  AND U18287 ( .A(n17265), .B(n17266), .Z(n17264) );
  XNOR U18288 ( .A(n17263), .B(n8634), .Z(n17266) );
  XNOR U18289 ( .A(n17259), .B(n17261), .Z(n8634) );
  NAND U18290 ( .A(n17267), .B(e_input[611]), .Z(n17261) );
  NAND U18291 ( .A(n12323), .B(e_input[611]), .Z(n17267) );
  XNOR U18292 ( .A(n17257), .B(n17268), .Z(n17259) );
  XOR U18293 ( .A(n17269), .B(n17270), .Z(n17257) );
  AND U18294 ( .A(n17271), .B(n17272), .Z(n17270) );
  XNOR U18295 ( .A(n17273), .B(n17269), .Z(n17272) );
  XOR U18296 ( .A(n17274), .B(e_input[611]), .Z(n17265) );
  IV U18297 ( .A(n17263), .Z(n17274) );
  XOR U18298 ( .A(n17275), .B(n17276), .Z(n17263) );
  AND U18299 ( .A(n17277), .B(n17278), .Z(n17276) );
  XNOR U18300 ( .A(n17275), .B(n8640), .Z(n17278) );
  XNOR U18301 ( .A(n17271), .B(n17273), .Z(n8640) );
  NAND U18302 ( .A(n17279), .B(e_input[610]), .Z(n17273) );
  NAND U18303 ( .A(n12323), .B(e_input[610]), .Z(n17279) );
  XNOR U18304 ( .A(n17269), .B(n17280), .Z(n17271) );
  XOR U18305 ( .A(n17281), .B(n17282), .Z(n17269) );
  AND U18306 ( .A(n17283), .B(n17284), .Z(n17282) );
  XNOR U18307 ( .A(n17285), .B(n17281), .Z(n17284) );
  XOR U18308 ( .A(n17286), .B(e_input[610]), .Z(n17277) );
  IV U18309 ( .A(n17275), .Z(n17286) );
  XOR U18310 ( .A(n17287), .B(n17288), .Z(n17275) );
  AND U18311 ( .A(n17289), .B(n17290), .Z(n17288) );
  XNOR U18312 ( .A(n17287), .B(n8646), .Z(n17290) );
  XNOR U18313 ( .A(n17283), .B(n17285), .Z(n8646) );
  NAND U18314 ( .A(n17291), .B(e_input[609]), .Z(n17285) );
  NAND U18315 ( .A(n12323), .B(e_input[609]), .Z(n17291) );
  XNOR U18316 ( .A(n17281), .B(n17292), .Z(n17283) );
  XOR U18317 ( .A(n17293), .B(n17294), .Z(n17281) );
  AND U18318 ( .A(n17295), .B(n17296), .Z(n17294) );
  XNOR U18319 ( .A(n17297), .B(n17293), .Z(n17296) );
  XOR U18320 ( .A(n17298), .B(e_input[609]), .Z(n17289) );
  IV U18321 ( .A(n17287), .Z(n17298) );
  XOR U18322 ( .A(n17299), .B(n17300), .Z(n17287) );
  AND U18323 ( .A(n17301), .B(n17302), .Z(n17300) );
  XNOR U18324 ( .A(n17299), .B(n8652), .Z(n17302) );
  XNOR U18325 ( .A(n17295), .B(n17297), .Z(n8652) );
  NAND U18326 ( .A(n17303), .B(e_input[608]), .Z(n17297) );
  NAND U18327 ( .A(n12323), .B(e_input[608]), .Z(n17303) );
  XNOR U18328 ( .A(n17293), .B(n17304), .Z(n17295) );
  XOR U18329 ( .A(n17305), .B(n17306), .Z(n17293) );
  AND U18330 ( .A(n17307), .B(n17308), .Z(n17306) );
  XNOR U18331 ( .A(n17309), .B(n17305), .Z(n17308) );
  XOR U18332 ( .A(n17310), .B(e_input[608]), .Z(n17301) );
  IV U18333 ( .A(n17299), .Z(n17310) );
  XOR U18334 ( .A(n17311), .B(n17312), .Z(n17299) );
  AND U18335 ( .A(n17313), .B(n17314), .Z(n17312) );
  XNOR U18336 ( .A(n17311), .B(n8658), .Z(n17314) );
  XNOR U18337 ( .A(n17307), .B(n17309), .Z(n8658) );
  NAND U18338 ( .A(n17315), .B(e_input[607]), .Z(n17309) );
  NAND U18339 ( .A(n12323), .B(e_input[607]), .Z(n17315) );
  XNOR U18340 ( .A(n17305), .B(n17316), .Z(n17307) );
  XOR U18341 ( .A(n17317), .B(n17318), .Z(n17305) );
  AND U18342 ( .A(n17319), .B(n17320), .Z(n17318) );
  XNOR U18343 ( .A(n17321), .B(n17317), .Z(n17320) );
  XOR U18344 ( .A(n17322), .B(e_input[607]), .Z(n17313) );
  IV U18345 ( .A(n17311), .Z(n17322) );
  XOR U18346 ( .A(n17323), .B(n17324), .Z(n17311) );
  AND U18347 ( .A(n17325), .B(n17326), .Z(n17324) );
  XNOR U18348 ( .A(n17323), .B(n8664), .Z(n17326) );
  XNOR U18349 ( .A(n17319), .B(n17321), .Z(n8664) );
  NAND U18350 ( .A(n17327), .B(e_input[606]), .Z(n17321) );
  NAND U18351 ( .A(n12323), .B(e_input[606]), .Z(n17327) );
  XNOR U18352 ( .A(n17317), .B(n17328), .Z(n17319) );
  XOR U18353 ( .A(n17329), .B(n17330), .Z(n17317) );
  AND U18354 ( .A(n17331), .B(n17332), .Z(n17330) );
  XNOR U18355 ( .A(n17333), .B(n17329), .Z(n17332) );
  XOR U18356 ( .A(n17334), .B(e_input[606]), .Z(n17325) );
  IV U18357 ( .A(n17323), .Z(n17334) );
  XOR U18358 ( .A(n17335), .B(n17336), .Z(n17323) );
  AND U18359 ( .A(n17337), .B(n17338), .Z(n17336) );
  XNOR U18360 ( .A(n17335), .B(n8670), .Z(n17338) );
  XNOR U18361 ( .A(n17331), .B(n17333), .Z(n8670) );
  NAND U18362 ( .A(n17339), .B(e_input[605]), .Z(n17333) );
  NAND U18363 ( .A(n12323), .B(e_input[605]), .Z(n17339) );
  XNOR U18364 ( .A(n17329), .B(n17340), .Z(n17331) );
  XOR U18365 ( .A(n17341), .B(n17342), .Z(n17329) );
  AND U18366 ( .A(n17343), .B(n17344), .Z(n17342) );
  XNOR U18367 ( .A(n17345), .B(n17341), .Z(n17344) );
  XOR U18368 ( .A(n17346), .B(e_input[605]), .Z(n17337) );
  IV U18369 ( .A(n17335), .Z(n17346) );
  XOR U18370 ( .A(n17347), .B(n17348), .Z(n17335) );
  AND U18371 ( .A(n17349), .B(n17350), .Z(n17348) );
  XNOR U18372 ( .A(n17347), .B(n8676), .Z(n17350) );
  XNOR U18373 ( .A(n17343), .B(n17345), .Z(n8676) );
  NAND U18374 ( .A(n17351), .B(e_input[604]), .Z(n17345) );
  NAND U18375 ( .A(n12323), .B(e_input[604]), .Z(n17351) );
  XNOR U18376 ( .A(n17341), .B(n17352), .Z(n17343) );
  XOR U18377 ( .A(n17353), .B(n17354), .Z(n17341) );
  AND U18378 ( .A(n17355), .B(n17356), .Z(n17354) );
  XNOR U18379 ( .A(n17357), .B(n17353), .Z(n17356) );
  XOR U18380 ( .A(n17358), .B(e_input[604]), .Z(n17349) );
  IV U18381 ( .A(n17347), .Z(n17358) );
  XOR U18382 ( .A(n17359), .B(n17360), .Z(n17347) );
  AND U18383 ( .A(n17361), .B(n17362), .Z(n17360) );
  XNOR U18384 ( .A(n17359), .B(n8682), .Z(n17362) );
  XNOR U18385 ( .A(n17355), .B(n17357), .Z(n8682) );
  NAND U18386 ( .A(n17363), .B(e_input[603]), .Z(n17357) );
  NAND U18387 ( .A(n12323), .B(e_input[603]), .Z(n17363) );
  XNOR U18388 ( .A(n17353), .B(n17364), .Z(n17355) );
  XOR U18389 ( .A(n17365), .B(n17366), .Z(n17353) );
  AND U18390 ( .A(n17367), .B(n17368), .Z(n17366) );
  XNOR U18391 ( .A(n17369), .B(n17365), .Z(n17368) );
  XOR U18392 ( .A(n17370), .B(e_input[603]), .Z(n17361) );
  IV U18393 ( .A(n17359), .Z(n17370) );
  XOR U18394 ( .A(n17371), .B(n17372), .Z(n17359) );
  AND U18395 ( .A(n17373), .B(n17374), .Z(n17372) );
  XNOR U18396 ( .A(n17371), .B(n8688), .Z(n17374) );
  XNOR U18397 ( .A(n17367), .B(n17369), .Z(n8688) );
  NAND U18398 ( .A(n17375), .B(e_input[602]), .Z(n17369) );
  NAND U18399 ( .A(n12323), .B(e_input[602]), .Z(n17375) );
  XNOR U18400 ( .A(n17365), .B(n17376), .Z(n17367) );
  XOR U18401 ( .A(n17377), .B(n17378), .Z(n17365) );
  AND U18402 ( .A(n17379), .B(n17380), .Z(n17378) );
  XNOR U18403 ( .A(n17381), .B(n17377), .Z(n17380) );
  XOR U18404 ( .A(n17382), .B(e_input[602]), .Z(n17373) );
  IV U18405 ( .A(n17371), .Z(n17382) );
  XOR U18406 ( .A(n17383), .B(n17384), .Z(n17371) );
  AND U18407 ( .A(n17385), .B(n17386), .Z(n17384) );
  XNOR U18408 ( .A(n17383), .B(n8694), .Z(n17386) );
  XNOR U18409 ( .A(n17379), .B(n17381), .Z(n8694) );
  NAND U18410 ( .A(n17387), .B(e_input[601]), .Z(n17381) );
  NAND U18411 ( .A(n12323), .B(e_input[601]), .Z(n17387) );
  XNOR U18412 ( .A(n17377), .B(n17388), .Z(n17379) );
  XOR U18413 ( .A(n17389), .B(n17390), .Z(n17377) );
  AND U18414 ( .A(n17391), .B(n17392), .Z(n17390) );
  XNOR U18415 ( .A(n17393), .B(n17389), .Z(n17392) );
  XOR U18416 ( .A(n17394), .B(e_input[601]), .Z(n17385) );
  IV U18417 ( .A(n17383), .Z(n17394) );
  XOR U18418 ( .A(n17395), .B(n17396), .Z(n17383) );
  AND U18419 ( .A(n17397), .B(n17398), .Z(n17396) );
  XNOR U18420 ( .A(n17395), .B(n8700), .Z(n17398) );
  XNOR U18421 ( .A(n17391), .B(n17393), .Z(n8700) );
  NAND U18422 ( .A(n17399), .B(e_input[600]), .Z(n17393) );
  NAND U18423 ( .A(n12323), .B(e_input[600]), .Z(n17399) );
  XNOR U18424 ( .A(n17389), .B(n17400), .Z(n17391) );
  XOR U18425 ( .A(n17401), .B(n17402), .Z(n17389) );
  AND U18426 ( .A(n17403), .B(n17404), .Z(n17402) );
  XNOR U18427 ( .A(n17405), .B(n17401), .Z(n17404) );
  XOR U18428 ( .A(n17406), .B(e_input[600]), .Z(n17397) );
  IV U18429 ( .A(n17395), .Z(n17406) );
  XOR U18430 ( .A(n17407), .B(n17408), .Z(n17395) );
  AND U18431 ( .A(n17409), .B(n17410), .Z(n17408) );
  XNOR U18432 ( .A(n17407), .B(n8706), .Z(n17410) );
  XNOR U18433 ( .A(n17403), .B(n17405), .Z(n8706) );
  NAND U18434 ( .A(n17411), .B(e_input[599]), .Z(n17405) );
  NAND U18435 ( .A(n12323), .B(e_input[599]), .Z(n17411) );
  XNOR U18436 ( .A(n17401), .B(n17412), .Z(n17403) );
  XOR U18437 ( .A(n17413), .B(n17414), .Z(n17401) );
  AND U18438 ( .A(n17415), .B(n17416), .Z(n17414) );
  XNOR U18439 ( .A(n17417), .B(n17413), .Z(n17416) );
  XOR U18440 ( .A(n17418), .B(e_input[599]), .Z(n17409) );
  IV U18441 ( .A(n17407), .Z(n17418) );
  XOR U18442 ( .A(n17419), .B(n17420), .Z(n17407) );
  AND U18443 ( .A(n17421), .B(n17422), .Z(n17420) );
  XNOR U18444 ( .A(n17419), .B(n8712), .Z(n17422) );
  XNOR U18445 ( .A(n17415), .B(n17417), .Z(n8712) );
  NAND U18446 ( .A(n17423), .B(e_input[598]), .Z(n17417) );
  NAND U18447 ( .A(n12323), .B(e_input[598]), .Z(n17423) );
  XNOR U18448 ( .A(n17413), .B(n17424), .Z(n17415) );
  XOR U18449 ( .A(n17425), .B(n17426), .Z(n17413) );
  AND U18450 ( .A(n17427), .B(n17428), .Z(n17426) );
  XNOR U18451 ( .A(n17429), .B(n17425), .Z(n17428) );
  XOR U18452 ( .A(n17430), .B(e_input[598]), .Z(n17421) );
  IV U18453 ( .A(n17419), .Z(n17430) );
  XOR U18454 ( .A(n17431), .B(n17432), .Z(n17419) );
  AND U18455 ( .A(n17433), .B(n17434), .Z(n17432) );
  XNOR U18456 ( .A(n17431), .B(n8718), .Z(n17434) );
  XNOR U18457 ( .A(n17427), .B(n17429), .Z(n8718) );
  NAND U18458 ( .A(n17435), .B(e_input[597]), .Z(n17429) );
  NAND U18459 ( .A(n12323), .B(e_input[597]), .Z(n17435) );
  XNOR U18460 ( .A(n17425), .B(n17436), .Z(n17427) );
  XOR U18461 ( .A(n17437), .B(n17438), .Z(n17425) );
  AND U18462 ( .A(n17439), .B(n17440), .Z(n17438) );
  XNOR U18463 ( .A(n17441), .B(n17437), .Z(n17440) );
  XOR U18464 ( .A(n17442), .B(e_input[597]), .Z(n17433) );
  IV U18465 ( .A(n17431), .Z(n17442) );
  XOR U18466 ( .A(n17443), .B(n17444), .Z(n17431) );
  AND U18467 ( .A(n17445), .B(n17446), .Z(n17444) );
  XNOR U18468 ( .A(n17443), .B(n8724), .Z(n17446) );
  XNOR U18469 ( .A(n17439), .B(n17441), .Z(n8724) );
  NAND U18470 ( .A(n17447), .B(e_input[596]), .Z(n17441) );
  NAND U18471 ( .A(n12323), .B(e_input[596]), .Z(n17447) );
  XNOR U18472 ( .A(n17437), .B(n17448), .Z(n17439) );
  XOR U18473 ( .A(n17449), .B(n17450), .Z(n17437) );
  AND U18474 ( .A(n17451), .B(n17452), .Z(n17450) );
  XNOR U18475 ( .A(n17453), .B(n17449), .Z(n17452) );
  XOR U18476 ( .A(n17454), .B(e_input[596]), .Z(n17445) );
  IV U18477 ( .A(n17443), .Z(n17454) );
  XOR U18478 ( .A(n17455), .B(n17456), .Z(n17443) );
  AND U18479 ( .A(n17457), .B(n17458), .Z(n17456) );
  XNOR U18480 ( .A(n17455), .B(n8730), .Z(n17458) );
  XNOR U18481 ( .A(n17451), .B(n17453), .Z(n8730) );
  NAND U18482 ( .A(n17459), .B(e_input[595]), .Z(n17453) );
  NAND U18483 ( .A(n12323), .B(e_input[595]), .Z(n17459) );
  XNOR U18484 ( .A(n17449), .B(n17460), .Z(n17451) );
  XOR U18485 ( .A(n17461), .B(n17462), .Z(n17449) );
  AND U18486 ( .A(n17463), .B(n17464), .Z(n17462) );
  XNOR U18487 ( .A(n17465), .B(n17461), .Z(n17464) );
  XOR U18488 ( .A(n17466), .B(e_input[595]), .Z(n17457) );
  IV U18489 ( .A(n17455), .Z(n17466) );
  XOR U18490 ( .A(n17467), .B(n17468), .Z(n17455) );
  AND U18491 ( .A(n17469), .B(n17470), .Z(n17468) );
  XNOR U18492 ( .A(n17467), .B(n8736), .Z(n17470) );
  XNOR U18493 ( .A(n17463), .B(n17465), .Z(n8736) );
  NAND U18494 ( .A(n17471), .B(e_input[594]), .Z(n17465) );
  NAND U18495 ( .A(n12323), .B(e_input[594]), .Z(n17471) );
  XNOR U18496 ( .A(n17461), .B(n17472), .Z(n17463) );
  XOR U18497 ( .A(n17473), .B(n17474), .Z(n17461) );
  AND U18498 ( .A(n17475), .B(n17476), .Z(n17474) );
  XNOR U18499 ( .A(n17477), .B(n17473), .Z(n17476) );
  XOR U18500 ( .A(n17478), .B(e_input[594]), .Z(n17469) );
  IV U18501 ( .A(n17467), .Z(n17478) );
  XOR U18502 ( .A(n17479), .B(n17480), .Z(n17467) );
  AND U18503 ( .A(n17481), .B(n17482), .Z(n17480) );
  XNOR U18504 ( .A(n17479), .B(n8742), .Z(n17482) );
  XNOR U18505 ( .A(n17475), .B(n17477), .Z(n8742) );
  NAND U18506 ( .A(n17483), .B(e_input[593]), .Z(n17477) );
  NAND U18507 ( .A(n12323), .B(e_input[593]), .Z(n17483) );
  XNOR U18508 ( .A(n17473), .B(n17484), .Z(n17475) );
  XOR U18509 ( .A(n17485), .B(n17486), .Z(n17473) );
  AND U18510 ( .A(n17487), .B(n17488), .Z(n17486) );
  XNOR U18511 ( .A(n17489), .B(n17485), .Z(n17488) );
  XOR U18512 ( .A(n17490), .B(e_input[593]), .Z(n17481) );
  IV U18513 ( .A(n17479), .Z(n17490) );
  XOR U18514 ( .A(n17491), .B(n17492), .Z(n17479) );
  AND U18515 ( .A(n17493), .B(n17494), .Z(n17492) );
  XNOR U18516 ( .A(n17491), .B(n8748), .Z(n17494) );
  XNOR U18517 ( .A(n17487), .B(n17489), .Z(n8748) );
  NAND U18518 ( .A(n17495), .B(e_input[592]), .Z(n17489) );
  NAND U18519 ( .A(n12323), .B(e_input[592]), .Z(n17495) );
  XNOR U18520 ( .A(n17485), .B(n17496), .Z(n17487) );
  XOR U18521 ( .A(n17497), .B(n17498), .Z(n17485) );
  AND U18522 ( .A(n17499), .B(n17500), .Z(n17498) );
  XNOR U18523 ( .A(n17501), .B(n17497), .Z(n17500) );
  XOR U18524 ( .A(n17502), .B(e_input[592]), .Z(n17493) );
  IV U18525 ( .A(n17491), .Z(n17502) );
  XOR U18526 ( .A(n17503), .B(n17504), .Z(n17491) );
  AND U18527 ( .A(n17505), .B(n17506), .Z(n17504) );
  XNOR U18528 ( .A(n17503), .B(n8754), .Z(n17506) );
  XNOR U18529 ( .A(n17499), .B(n17501), .Z(n8754) );
  NAND U18530 ( .A(n17507), .B(e_input[591]), .Z(n17501) );
  NAND U18531 ( .A(n12323), .B(e_input[591]), .Z(n17507) );
  XNOR U18532 ( .A(n17497), .B(n17508), .Z(n17499) );
  XOR U18533 ( .A(n17509), .B(n17510), .Z(n17497) );
  AND U18534 ( .A(n17511), .B(n17512), .Z(n17510) );
  XNOR U18535 ( .A(n17513), .B(n17509), .Z(n17512) );
  XOR U18536 ( .A(n17514), .B(e_input[591]), .Z(n17505) );
  IV U18537 ( .A(n17503), .Z(n17514) );
  XOR U18538 ( .A(n17515), .B(n17516), .Z(n17503) );
  AND U18539 ( .A(n17517), .B(n17518), .Z(n17516) );
  XNOR U18540 ( .A(n17515), .B(n8760), .Z(n17518) );
  XNOR U18541 ( .A(n17511), .B(n17513), .Z(n8760) );
  NAND U18542 ( .A(n17519), .B(e_input[590]), .Z(n17513) );
  NAND U18543 ( .A(n12323), .B(e_input[590]), .Z(n17519) );
  XNOR U18544 ( .A(n17509), .B(n17520), .Z(n17511) );
  XOR U18545 ( .A(n17521), .B(n17522), .Z(n17509) );
  AND U18546 ( .A(n17523), .B(n17524), .Z(n17522) );
  XNOR U18547 ( .A(n17525), .B(n17521), .Z(n17524) );
  XOR U18548 ( .A(n17526), .B(e_input[590]), .Z(n17517) );
  IV U18549 ( .A(n17515), .Z(n17526) );
  XOR U18550 ( .A(n17527), .B(n17528), .Z(n17515) );
  AND U18551 ( .A(n17529), .B(n17530), .Z(n17528) );
  XNOR U18552 ( .A(n17527), .B(n8766), .Z(n17530) );
  XNOR U18553 ( .A(n17523), .B(n17525), .Z(n8766) );
  NAND U18554 ( .A(n17531), .B(e_input[589]), .Z(n17525) );
  NAND U18555 ( .A(n12323), .B(e_input[589]), .Z(n17531) );
  XNOR U18556 ( .A(n17521), .B(n17532), .Z(n17523) );
  XOR U18557 ( .A(n17533), .B(n17534), .Z(n17521) );
  AND U18558 ( .A(n17535), .B(n17536), .Z(n17534) );
  XNOR U18559 ( .A(n17537), .B(n17533), .Z(n17536) );
  XOR U18560 ( .A(n17538), .B(e_input[589]), .Z(n17529) );
  IV U18561 ( .A(n17527), .Z(n17538) );
  XOR U18562 ( .A(n17539), .B(n17540), .Z(n17527) );
  AND U18563 ( .A(n17541), .B(n17542), .Z(n17540) );
  XNOR U18564 ( .A(n17539), .B(n8772), .Z(n17542) );
  XNOR U18565 ( .A(n17535), .B(n17537), .Z(n8772) );
  NAND U18566 ( .A(n17543), .B(e_input[588]), .Z(n17537) );
  NAND U18567 ( .A(n12323), .B(e_input[588]), .Z(n17543) );
  XNOR U18568 ( .A(n17533), .B(n17544), .Z(n17535) );
  XOR U18569 ( .A(n17545), .B(n17546), .Z(n17533) );
  AND U18570 ( .A(n17547), .B(n17548), .Z(n17546) );
  XNOR U18571 ( .A(n17549), .B(n17545), .Z(n17548) );
  XOR U18572 ( .A(n17550), .B(e_input[588]), .Z(n17541) );
  IV U18573 ( .A(n17539), .Z(n17550) );
  XOR U18574 ( .A(n17551), .B(n17552), .Z(n17539) );
  AND U18575 ( .A(n17553), .B(n17554), .Z(n17552) );
  XNOR U18576 ( .A(n17551), .B(n8778), .Z(n17554) );
  XNOR U18577 ( .A(n17547), .B(n17549), .Z(n8778) );
  NAND U18578 ( .A(n17555), .B(e_input[587]), .Z(n17549) );
  NAND U18579 ( .A(n12323), .B(e_input[587]), .Z(n17555) );
  XNOR U18580 ( .A(n17545), .B(n17556), .Z(n17547) );
  XOR U18581 ( .A(n17557), .B(n17558), .Z(n17545) );
  AND U18582 ( .A(n17559), .B(n17560), .Z(n17558) );
  XNOR U18583 ( .A(n17561), .B(n17557), .Z(n17560) );
  XOR U18584 ( .A(n17562), .B(e_input[587]), .Z(n17553) );
  IV U18585 ( .A(n17551), .Z(n17562) );
  XOR U18586 ( .A(n17563), .B(n17564), .Z(n17551) );
  AND U18587 ( .A(n17565), .B(n17566), .Z(n17564) );
  XNOR U18588 ( .A(n17563), .B(n8784), .Z(n17566) );
  XNOR U18589 ( .A(n17559), .B(n17561), .Z(n8784) );
  NAND U18590 ( .A(n17567), .B(e_input[586]), .Z(n17561) );
  NAND U18591 ( .A(n12323), .B(e_input[586]), .Z(n17567) );
  XNOR U18592 ( .A(n17557), .B(n17568), .Z(n17559) );
  XOR U18593 ( .A(n17569), .B(n17570), .Z(n17557) );
  AND U18594 ( .A(n17571), .B(n17572), .Z(n17570) );
  XNOR U18595 ( .A(n17573), .B(n17569), .Z(n17572) );
  XOR U18596 ( .A(n17574), .B(e_input[586]), .Z(n17565) );
  IV U18597 ( .A(n17563), .Z(n17574) );
  XOR U18598 ( .A(n17575), .B(n17576), .Z(n17563) );
  AND U18599 ( .A(n17577), .B(n17578), .Z(n17576) );
  XNOR U18600 ( .A(n17575), .B(n8790), .Z(n17578) );
  XNOR U18601 ( .A(n17571), .B(n17573), .Z(n8790) );
  NAND U18602 ( .A(n17579), .B(e_input[585]), .Z(n17573) );
  NAND U18603 ( .A(n12323), .B(e_input[585]), .Z(n17579) );
  XNOR U18604 ( .A(n17569), .B(n17580), .Z(n17571) );
  XOR U18605 ( .A(n17581), .B(n17582), .Z(n17569) );
  AND U18606 ( .A(n17583), .B(n17584), .Z(n17582) );
  XNOR U18607 ( .A(n17585), .B(n17581), .Z(n17584) );
  XOR U18608 ( .A(n17586), .B(e_input[585]), .Z(n17577) );
  IV U18609 ( .A(n17575), .Z(n17586) );
  XOR U18610 ( .A(n17587), .B(n17588), .Z(n17575) );
  AND U18611 ( .A(n17589), .B(n17590), .Z(n17588) );
  XNOR U18612 ( .A(n17587), .B(n8796), .Z(n17590) );
  XNOR U18613 ( .A(n17583), .B(n17585), .Z(n8796) );
  NAND U18614 ( .A(n17591), .B(e_input[584]), .Z(n17585) );
  NAND U18615 ( .A(n12323), .B(e_input[584]), .Z(n17591) );
  XNOR U18616 ( .A(n17581), .B(n17592), .Z(n17583) );
  XOR U18617 ( .A(n17593), .B(n17594), .Z(n17581) );
  AND U18618 ( .A(n17595), .B(n17596), .Z(n17594) );
  XNOR U18619 ( .A(n17597), .B(n17593), .Z(n17596) );
  XOR U18620 ( .A(n17598), .B(e_input[584]), .Z(n17589) );
  IV U18621 ( .A(n17587), .Z(n17598) );
  XOR U18622 ( .A(n17599), .B(n17600), .Z(n17587) );
  AND U18623 ( .A(n17601), .B(n17602), .Z(n17600) );
  XNOR U18624 ( .A(n17599), .B(n8802), .Z(n17602) );
  XNOR U18625 ( .A(n17595), .B(n17597), .Z(n8802) );
  NAND U18626 ( .A(n17603), .B(e_input[583]), .Z(n17597) );
  NAND U18627 ( .A(n12323), .B(e_input[583]), .Z(n17603) );
  XNOR U18628 ( .A(n17593), .B(n17604), .Z(n17595) );
  XOR U18629 ( .A(n17605), .B(n17606), .Z(n17593) );
  AND U18630 ( .A(n17607), .B(n17608), .Z(n17606) );
  XNOR U18631 ( .A(n17609), .B(n17605), .Z(n17608) );
  XOR U18632 ( .A(n17610), .B(e_input[583]), .Z(n17601) );
  IV U18633 ( .A(n17599), .Z(n17610) );
  XOR U18634 ( .A(n17611), .B(n17612), .Z(n17599) );
  AND U18635 ( .A(n17613), .B(n17614), .Z(n17612) );
  XNOR U18636 ( .A(n17611), .B(n8808), .Z(n17614) );
  XNOR U18637 ( .A(n17607), .B(n17609), .Z(n8808) );
  NAND U18638 ( .A(n17615), .B(e_input[582]), .Z(n17609) );
  NAND U18639 ( .A(n12323), .B(e_input[582]), .Z(n17615) );
  XNOR U18640 ( .A(n17605), .B(n17616), .Z(n17607) );
  XOR U18641 ( .A(n17617), .B(n17618), .Z(n17605) );
  AND U18642 ( .A(n17619), .B(n17620), .Z(n17618) );
  XNOR U18643 ( .A(n17621), .B(n17617), .Z(n17620) );
  XOR U18644 ( .A(n17622), .B(e_input[582]), .Z(n17613) );
  IV U18645 ( .A(n17611), .Z(n17622) );
  XOR U18646 ( .A(n17623), .B(n17624), .Z(n17611) );
  AND U18647 ( .A(n17625), .B(n17626), .Z(n17624) );
  XNOR U18648 ( .A(n17623), .B(n8814), .Z(n17626) );
  XNOR U18649 ( .A(n17619), .B(n17621), .Z(n8814) );
  NAND U18650 ( .A(n17627), .B(e_input[581]), .Z(n17621) );
  NAND U18651 ( .A(n12323), .B(e_input[581]), .Z(n17627) );
  XNOR U18652 ( .A(n17617), .B(n17628), .Z(n17619) );
  XOR U18653 ( .A(n17629), .B(n17630), .Z(n17617) );
  AND U18654 ( .A(n17631), .B(n17632), .Z(n17630) );
  XNOR U18655 ( .A(n17633), .B(n17629), .Z(n17632) );
  XOR U18656 ( .A(n17634), .B(e_input[581]), .Z(n17625) );
  IV U18657 ( .A(n17623), .Z(n17634) );
  XOR U18658 ( .A(n17635), .B(n17636), .Z(n17623) );
  AND U18659 ( .A(n17637), .B(n17638), .Z(n17636) );
  XNOR U18660 ( .A(n17635), .B(n8820), .Z(n17638) );
  XNOR U18661 ( .A(n17631), .B(n17633), .Z(n8820) );
  NAND U18662 ( .A(n17639), .B(e_input[580]), .Z(n17633) );
  NAND U18663 ( .A(n12323), .B(e_input[580]), .Z(n17639) );
  XNOR U18664 ( .A(n17629), .B(n17640), .Z(n17631) );
  XOR U18665 ( .A(n17641), .B(n17642), .Z(n17629) );
  AND U18666 ( .A(n17643), .B(n17644), .Z(n17642) );
  XNOR U18667 ( .A(n17645), .B(n17641), .Z(n17644) );
  XOR U18668 ( .A(n17646), .B(e_input[580]), .Z(n17637) );
  IV U18669 ( .A(n17635), .Z(n17646) );
  XOR U18670 ( .A(n17647), .B(n17648), .Z(n17635) );
  AND U18671 ( .A(n17649), .B(n17650), .Z(n17648) );
  XNOR U18672 ( .A(n17647), .B(n8826), .Z(n17650) );
  XNOR U18673 ( .A(n17643), .B(n17645), .Z(n8826) );
  NAND U18674 ( .A(n17651), .B(e_input[579]), .Z(n17645) );
  NAND U18675 ( .A(n12323), .B(e_input[579]), .Z(n17651) );
  XNOR U18676 ( .A(n17641), .B(n17652), .Z(n17643) );
  XOR U18677 ( .A(n17653), .B(n17654), .Z(n17641) );
  AND U18678 ( .A(n17655), .B(n17656), .Z(n17654) );
  XNOR U18679 ( .A(n17657), .B(n17653), .Z(n17656) );
  XOR U18680 ( .A(n17658), .B(e_input[579]), .Z(n17649) );
  IV U18681 ( .A(n17647), .Z(n17658) );
  XOR U18682 ( .A(n17659), .B(n17660), .Z(n17647) );
  AND U18683 ( .A(n17661), .B(n17662), .Z(n17660) );
  XNOR U18684 ( .A(n17659), .B(n8832), .Z(n17662) );
  XNOR U18685 ( .A(n17655), .B(n17657), .Z(n8832) );
  NAND U18686 ( .A(n17663), .B(e_input[578]), .Z(n17657) );
  NAND U18687 ( .A(n12323), .B(e_input[578]), .Z(n17663) );
  XNOR U18688 ( .A(n17653), .B(n17664), .Z(n17655) );
  XOR U18689 ( .A(n17665), .B(n17666), .Z(n17653) );
  AND U18690 ( .A(n17667), .B(n17668), .Z(n17666) );
  XNOR U18691 ( .A(n17669), .B(n17665), .Z(n17668) );
  XOR U18692 ( .A(n17670), .B(e_input[578]), .Z(n17661) );
  IV U18693 ( .A(n17659), .Z(n17670) );
  XOR U18694 ( .A(n17671), .B(n17672), .Z(n17659) );
  AND U18695 ( .A(n17673), .B(n17674), .Z(n17672) );
  XNOR U18696 ( .A(n17671), .B(n8838), .Z(n17674) );
  XNOR U18697 ( .A(n17667), .B(n17669), .Z(n8838) );
  NAND U18698 ( .A(n17675), .B(e_input[577]), .Z(n17669) );
  NAND U18699 ( .A(n12323), .B(e_input[577]), .Z(n17675) );
  XNOR U18700 ( .A(n17665), .B(n17676), .Z(n17667) );
  XOR U18701 ( .A(n17677), .B(n17678), .Z(n17665) );
  AND U18702 ( .A(n17679), .B(n17680), .Z(n17678) );
  XNOR U18703 ( .A(n17681), .B(n17677), .Z(n17680) );
  XOR U18704 ( .A(n17682), .B(e_input[577]), .Z(n17673) );
  IV U18705 ( .A(n17671), .Z(n17682) );
  XOR U18706 ( .A(n17683), .B(n17684), .Z(n17671) );
  AND U18707 ( .A(n17685), .B(n17686), .Z(n17684) );
  XNOR U18708 ( .A(n17683), .B(n8844), .Z(n17686) );
  XNOR U18709 ( .A(n17679), .B(n17681), .Z(n8844) );
  NAND U18710 ( .A(n17687), .B(e_input[576]), .Z(n17681) );
  NAND U18711 ( .A(n12323), .B(e_input[576]), .Z(n17687) );
  XNOR U18712 ( .A(n17677), .B(n17688), .Z(n17679) );
  XOR U18713 ( .A(n17689), .B(n17690), .Z(n17677) );
  AND U18714 ( .A(n17691), .B(n17692), .Z(n17690) );
  XNOR U18715 ( .A(n17693), .B(n17689), .Z(n17692) );
  XOR U18716 ( .A(n17694), .B(e_input[576]), .Z(n17685) );
  IV U18717 ( .A(n17683), .Z(n17694) );
  XOR U18718 ( .A(n17695), .B(n17696), .Z(n17683) );
  AND U18719 ( .A(n17697), .B(n17698), .Z(n17696) );
  XNOR U18720 ( .A(n17695), .B(n8850), .Z(n17698) );
  XNOR U18721 ( .A(n17691), .B(n17693), .Z(n8850) );
  NAND U18722 ( .A(n17699), .B(e_input[575]), .Z(n17693) );
  NAND U18723 ( .A(n12323), .B(e_input[575]), .Z(n17699) );
  XNOR U18724 ( .A(n17689), .B(n17700), .Z(n17691) );
  XOR U18725 ( .A(n17701), .B(n17702), .Z(n17689) );
  AND U18726 ( .A(n17703), .B(n17704), .Z(n17702) );
  XNOR U18727 ( .A(n17705), .B(n17701), .Z(n17704) );
  XOR U18728 ( .A(n17706), .B(e_input[575]), .Z(n17697) );
  IV U18729 ( .A(n17695), .Z(n17706) );
  XOR U18730 ( .A(n17707), .B(n17708), .Z(n17695) );
  AND U18731 ( .A(n17709), .B(n17710), .Z(n17708) );
  XNOR U18732 ( .A(n17707), .B(n8856), .Z(n17710) );
  XNOR U18733 ( .A(n17703), .B(n17705), .Z(n8856) );
  NAND U18734 ( .A(n17711), .B(e_input[574]), .Z(n17705) );
  NAND U18735 ( .A(n12323), .B(e_input[574]), .Z(n17711) );
  XNOR U18736 ( .A(n17701), .B(n17712), .Z(n17703) );
  XOR U18737 ( .A(n17713), .B(n17714), .Z(n17701) );
  AND U18738 ( .A(n17715), .B(n17716), .Z(n17714) );
  XNOR U18739 ( .A(n17717), .B(n17713), .Z(n17716) );
  XOR U18740 ( .A(n17718), .B(e_input[574]), .Z(n17709) );
  IV U18741 ( .A(n17707), .Z(n17718) );
  XOR U18742 ( .A(n17719), .B(n17720), .Z(n17707) );
  AND U18743 ( .A(n17721), .B(n17722), .Z(n17720) );
  XNOR U18744 ( .A(n17719), .B(n8862), .Z(n17722) );
  XNOR U18745 ( .A(n17715), .B(n17717), .Z(n8862) );
  NAND U18746 ( .A(n17723), .B(e_input[573]), .Z(n17717) );
  NAND U18747 ( .A(n12323), .B(e_input[573]), .Z(n17723) );
  XNOR U18748 ( .A(n17713), .B(n17724), .Z(n17715) );
  XOR U18749 ( .A(n17725), .B(n17726), .Z(n17713) );
  AND U18750 ( .A(n17727), .B(n17728), .Z(n17726) );
  XNOR U18751 ( .A(n17729), .B(n17725), .Z(n17728) );
  XOR U18752 ( .A(n17730), .B(e_input[573]), .Z(n17721) );
  IV U18753 ( .A(n17719), .Z(n17730) );
  XOR U18754 ( .A(n17731), .B(n17732), .Z(n17719) );
  AND U18755 ( .A(n17733), .B(n17734), .Z(n17732) );
  XNOR U18756 ( .A(n17731), .B(n8868), .Z(n17734) );
  XNOR U18757 ( .A(n17727), .B(n17729), .Z(n8868) );
  NAND U18758 ( .A(n17735), .B(e_input[572]), .Z(n17729) );
  NAND U18759 ( .A(n12323), .B(e_input[572]), .Z(n17735) );
  XNOR U18760 ( .A(n17725), .B(n17736), .Z(n17727) );
  XOR U18761 ( .A(n17737), .B(n17738), .Z(n17725) );
  AND U18762 ( .A(n17739), .B(n17740), .Z(n17738) );
  XNOR U18763 ( .A(n17741), .B(n17737), .Z(n17740) );
  XOR U18764 ( .A(n17742), .B(e_input[572]), .Z(n17733) );
  IV U18765 ( .A(n17731), .Z(n17742) );
  XOR U18766 ( .A(n17743), .B(n17744), .Z(n17731) );
  AND U18767 ( .A(n17745), .B(n17746), .Z(n17744) );
  XNOR U18768 ( .A(n17743), .B(n8874), .Z(n17746) );
  XNOR U18769 ( .A(n17739), .B(n17741), .Z(n8874) );
  NAND U18770 ( .A(n17747), .B(e_input[571]), .Z(n17741) );
  NAND U18771 ( .A(n12323), .B(e_input[571]), .Z(n17747) );
  XNOR U18772 ( .A(n17737), .B(n17748), .Z(n17739) );
  XOR U18773 ( .A(n17749), .B(n17750), .Z(n17737) );
  AND U18774 ( .A(n17751), .B(n17752), .Z(n17750) );
  XNOR U18775 ( .A(n17753), .B(n17749), .Z(n17752) );
  XOR U18776 ( .A(n17754), .B(e_input[571]), .Z(n17745) );
  IV U18777 ( .A(n17743), .Z(n17754) );
  XOR U18778 ( .A(n17755), .B(n17756), .Z(n17743) );
  AND U18779 ( .A(n17757), .B(n17758), .Z(n17756) );
  XNOR U18780 ( .A(n17755), .B(n8880), .Z(n17758) );
  XNOR U18781 ( .A(n17751), .B(n17753), .Z(n8880) );
  NAND U18782 ( .A(n17759), .B(e_input[570]), .Z(n17753) );
  NAND U18783 ( .A(n12323), .B(e_input[570]), .Z(n17759) );
  XNOR U18784 ( .A(n17749), .B(n17760), .Z(n17751) );
  XOR U18785 ( .A(n17761), .B(n17762), .Z(n17749) );
  AND U18786 ( .A(n17763), .B(n17764), .Z(n17762) );
  XNOR U18787 ( .A(n17765), .B(n17761), .Z(n17764) );
  XOR U18788 ( .A(n17766), .B(e_input[570]), .Z(n17757) );
  IV U18789 ( .A(n17755), .Z(n17766) );
  XOR U18790 ( .A(n17767), .B(n17768), .Z(n17755) );
  AND U18791 ( .A(n17769), .B(n17770), .Z(n17768) );
  XNOR U18792 ( .A(n17767), .B(n8886), .Z(n17770) );
  XNOR U18793 ( .A(n17763), .B(n17765), .Z(n8886) );
  NAND U18794 ( .A(n17771), .B(e_input[569]), .Z(n17765) );
  NAND U18795 ( .A(n12323), .B(e_input[569]), .Z(n17771) );
  XNOR U18796 ( .A(n17761), .B(n17772), .Z(n17763) );
  XOR U18797 ( .A(n17773), .B(n17774), .Z(n17761) );
  AND U18798 ( .A(n17775), .B(n17776), .Z(n17774) );
  XNOR U18799 ( .A(n17777), .B(n17773), .Z(n17776) );
  XOR U18800 ( .A(n17778), .B(e_input[569]), .Z(n17769) );
  IV U18801 ( .A(n17767), .Z(n17778) );
  XOR U18802 ( .A(n17779), .B(n17780), .Z(n17767) );
  AND U18803 ( .A(n17781), .B(n17782), .Z(n17780) );
  XNOR U18804 ( .A(n17779), .B(n8892), .Z(n17782) );
  XNOR U18805 ( .A(n17775), .B(n17777), .Z(n8892) );
  NAND U18806 ( .A(n17783), .B(e_input[568]), .Z(n17777) );
  NAND U18807 ( .A(n12323), .B(e_input[568]), .Z(n17783) );
  XNOR U18808 ( .A(n17773), .B(n17784), .Z(n17775) );
  XOR U18809 ( .A(n17785), .B(n17786), .Z(n17773) );
  AND U18810 ( .A(n17787), .B(n17788), .Z(n17786) );
  XNOR U18811 ( .A(n17789), .B(n17785), .Z(n17788) );
  XOR U18812 ( .A(n17790), .B(e_input[568]), .Z(n17781) );
  IV U18813 ( .A(n17779), .Z(n17790) );
  XOR U18814 ( .A(n17791), .B(n17792), .Z(n17779) );
  AND U18815 ( .A(n17793), .B(n17794), .Z(n17792) );
  XNOR U18816 ( .A(n17791), .B(n8898), .Z(n17794) );
  XNOR U18817 ( .A(n17787), .B(n17789), .Z(n8898) );
  NAND U18818 ( .A(n17795), .B(e_input[567]), .Z(n17789) );
  NAND U18819 ( .A(n12323), .B(e_input[567]), .Z(n17795) );
  XNOR U18820 ( .A(n17785), .B(n17796), .Z(n17787) );
  XOR U18821 ( .A(n17797), .B(n17798), .Z(n17785) );
  AND U18822 ( .A(n17799), .B(n17800), .Z(n17798) );
  XNOR U18823 ( .A(n17801), .B(n17797), .Z(n17800) );
  XOR U18824 ( .A(n17802), .B(e_input[567]), .Z(n17793) );
  IV U18825 ( .A(n17791), .Z(n17802) );
  XOR U18826 ( .A(n17803), .B(n17804), .Z(n17791) );
  AND U18827 ( .A(n17805), .B(n17806), .Z(n17804) );
  XNOR U18828 ( .A(n17803), .B(n8904), .Z(n17806) );
  XNOR U18829 ( .A(n17799), .B(n17801), .Z(n8904) );
  NAND U18830 ( .A(n17807), .B(e_input[566]), .Z(n17801) );
  NAND U18831 ( .A(n12323), .B(e_input[566]), .Z(n17807) );
  XNOR U18832 ( .A(n17797), .B(n17808), .Z(n17799) );
  XOR U18833 ( .A(n17809), .B(n17810), .Z(n17797) );
  AND U18834 ( .A(n17811), .B(n17812), .Z(n17810) );
  XNOR U18835 ( .A(n17813), .B(n17809), .Z(n17812) );
  XOR U18836 ( .A(n17814), .B(e_input[566]), .Z(n17805) );
  IV U18837 ( .A(n17803), .Z(n17814) );
  XOR U18838 ( .A(n17815), .B(n17816), .Z(n17803) );
  AND U18839 ( .A(n17817), .B(n17818), .Z(n17816) );
  XNOR U18840 ( .A(n17815), .B(n8910), .Z(n17818) );
  XNOR U18841 ( .A(n17811), .B(n17813), .Z(n8910) );
  NAND U18842 ( .A(n17819), .B(e_input[565]), .Z(n17813) );
  NAND U18843 ( .A(n12323), .B(e_input[565]), .Z(n17819) );
  XNOR U18844 ( .A(n17809), .B(n17820), .Z(n17811) );
  XOR U18845 ( .A(n17821), .B(n17822), .Z(n17809) );
  AND U18846 ( .A(n17823), .B(n17824), .Z(n17822) );
  XNOR U18847 ( .A(n17825), .B(n17821), .Z(n17824) );
  XOR U18848 ( .A(n17826), .B(e_input[565]), .Z(n17817) );
  IV U18849 ( .A(n17815), .Z(n17826) );
  XOR U18850 ( .A(n17827), .B(n17828), .Z(n17815) );
  AND U18851 ( .A(n17829), .B(n17830), .Z(n17828) );
  XNOR U18852 ( .A(n17827), .B(n8916), .Z(n17830) );
  XNOR U18853 ( .A(n17823), .B(n17825), .Z(n8916) );
  NAND U18854 ( .A(n17831), .B(e_input[564]), .Z(n17825) );
  NAND U18855 ( .A(n12323), .B(e_input[564]), .Z(n17831) );
  XNOR U18856 ( .A(n17821), .B(n17832), .Z(n17823) );
  XOR U18857 ( .A(n17833), .B(n17834), .Z(n17821) );
  AND U18858 ( .A(n17835), .B(n17836), .Z(n17834) );
  XNOR U18859 ( .A(n17837), .B(n17833), .Z(n17836) );
  XOR U18860 ( .A(n17838), .B(e_input[564]), .Z(n17829) );
  IV U18861 ( .A(n17827), .Z(n17838) );
  XOR U18862 ( .A(n17839), .B(n17840), .Z(n17827) );
  AND U18863 ( .A(n17841), .B(n17842), .Z(n17840) );
  XNOR U18864 ( .A(n17839), .B(n8922), .Z(n17842) );
  XNOR U18865 ( .A(n17835), .B(n17837), .Z(n8922) );
  NAND U18866 ( .A(n17843), .B(e_input[563]), .Z(n17837) );
  NAND U18867 ( .A(n12323), .B(e_input[563]), .Z(n17843) );
  XNOR U18868 ( .A(n17833), .B(n17844), .Z(n17835) );
  XOR U18869 ( .A(n17845), .B(n17846), .Z(n17833) );
  AND U18870 ( .A(n17847), .B(n17848), .Z(n17846) );
  XNOR U18871 ( .A(n17849), .B(n17845), .Z(n17848) );
  XOR U18872 ( .A(n17850), .B(e_input[563]), .Z(n17841) );
  IV U18873 ( .A(n17839), .Z(n17850) );
  XOR U18874 ( .A(n17851), .B(n17852), .Z(n17839) );
  AND U18875 ( .A(n17853), .B(n17854), .Z(n17852) );
  XNOR U18876 ( .A(n17851), .B(n8928), .Z(n17854) );
  XNOR U18877 ( .A(n17847), .B(n17849), .Z(n8928) );
  NAND U18878 ( .A(n17855), .B(e_input[562]), .Z(n17849) );
  NAND U18879 ( .A(n12323), .B(e_input[562]), .Z(n17855) );
  XNOR U18880 ( .A(n17845), .B(n17856), .Z(n17847) );
  XOR U18881 ( .A(n17857), .B(n17858), .Z(n17845) );
  AND U18882 ( .A(n17859), .B(n17860), .Z(n17858) );
  XNOR U18883 ( .A(n17861), .B(n17857), .Z(n17860) );
  XOR U18884 ( .A(n17862), .B(e_input[562]), .Z(n17853) );
  IV U18885 ( .A(n17851), .Z(n17862) );
  XOR U18886 ( .A(n17863), .B(n17864), .Z(n17851) );
  AND U18887 ( .A(n17865), .B(n17866), .Z(n17864) );
  XNOR U18888 ( .A(n17863), .B(n8934), .Z(n17866) );
  XNOR U18889 ( .A(n17859), .B(n17861), .Z(n8934) );
  NAND U18890 ( .A(n17867), .B(e_input[561]), .Z(n17861) );
  NAND U18891 ( .A(n12323), .B(e_input[561]), .Z(n17867) );
  XNOR U18892 ( .A(n17857), .B(n17868), .Z(n17859) );
  XOR U18893 ( .A(n17869), .B(n17870), .Z(n17857) );
  AND U18894 ( .A(n17871), .B(n17872), .Z(n17870) );
  XNOR U18895 ( .A(n17873), .B(n17869), .Z(n17872) );
  XOR U18896 ( .A(n17874), .B(e_input[561]), .Z(n17865) );
  IV U18897 ( .A(n17863), .Z(n17874) );
  XOR U18898 ( .A(n17875), .B(n17876), .Z(n17863) );
  AND U18899 ( .A(n17877), .B(n17878), .Z(n17876) );
  XNOR U18900 ( .A(n17875), .B(n8940), .Z(n17878) );
  XNOR U18901 ( .A(n17871), .B(n17873), .Z(n8940) );
  NAND U18902 ( .A(n17879), .B(e_input[560]), .Z(n17873) );
  NAND U18903 ( .A(n12323), .B(e_input[560]), .Z(n17879) );
  XNOR U18904 ( .A(n17869), .B(n17880), .Z(n17871) );
  XOR U18905 ( .A(n17881), .B(n17882), .Z(n17869) );
  AND U18906 ( .A(n17883), .B(n17884), .Z(n17882) );
  XNOR U18907 ( .A(n17885), .B(n17881), .Z(n17884) );
  XOR U18908 ( .A(n17886), .B(e_input[560]), .Z(n17877) );
  IV U18909 ( .A(n17875), .Z(n17886) );
  XOR U18910 ( .A(n17887), .B(n17888), .Z(n17875) );
  AND U18911 ( .A(n17889), .B(n17890), .Z(n17888) );
  XNOR U18912 ( .A(n17887), .B(n8946), .Z(n17890) );
  XNOR U18913 ( .A(n17883), .B(n17885), .Z(n8946) );
  NAND U18914 ( .A(n17891), .B(e_input[559]), .Z(n17885) );
  NAND U18915 ( .A(n12323), .B(e_input[559]), .Z(n17891) );
  XNOR U18916 ( .A(n17881), .B(n17892), .Z(n17883) );
  XOR U18917 ( .A(n17893), .B(n17894), .Z(n17881) );
  AND U18918 ( .A(n17895), .B(n17896), .Z(n17894) );
  XNOR U18919 ( .A(n17897), .B(n17893), .Z(n17896) );
  XOR U18920 ( .A(n17898), .B(e_input[559]), .Z(n17889) );
  IV U18921 ( .A(n17887), .Z(n17898) );
  XOR U18922 ( .A(n17899), .B(n17900), .Z(n17887) );
  AND U18923 ( .A(n17901), .B(n17902), .Z(n17900) );
  XNOR U18924 ( .A(n17899), .B(n8952), .Z(n17902) );
  XNOR U18925 ( .A(n17895), .B(n17897), .Z(n8952) );
  NAND U18926 ( .A(n17903), .B(e_input[558]), .Z(n17897) );
  NAND U18927 ( .A(n12323), .B(e_input[558]), .Z(n17903) );
  XNOR U18928 ( .A(n17893), .B(n17904), .Z(n17895) );
  XOR U18929 ( .A(n17905), .B(n17906), .Z(n17893) );
  AND U18930 ( .A(n17907), .B(n17908), .Z(n17906) );
  XNOR U18931 ( .A(n17909), .B(n17905), .Z(n17908) );
  XOR U18932 ( .A(n17910), .B(e_input[558]), .Z(n17901) );
  IV U18933 ( .A(n17899), .Z(n17910) );
  XOR U18934 ( .A(n17911), .B(n17912), .Z(n17899) );
  AND U18935 ( .A(n17913), .B(n17914), .Z(n17912) );
  XNOR U18936 ( .A(n17911), .B(n8958), .Z(n17914) );
  XNOR U18937 ( .A(n17907), .B(n17909), .Z(n8958) );
  NAND U18938 ( .A(n17915), .B(e_input[557]), .Z(n17909) );
  NAND U18939 ( .A(n12323), .B(e_input[557]), .Z(n17915) );
  XNOR U18940 ( .A(n17905), .B(n17916), .Z(n17907) );
  XOR U18941 ( .A(n17917), .B(n17918), .Z(n17905) );
  AND U18942 ( .A(n17919), .B(n17920), .Z(n17918) );
  XNOR U18943 ( .A(n17921), .B(n17917), .Z(n17920) );
  XOR U18944 ( .A(n17922), .B(e_input[557]), .Z(n17913) );
  IV U18945 ( .A(n17911), .Z(n17922) );
  XOR U18946 ( .A(n17923), .B(n17924), .Z(n17911) );
  AND U18947 ( .A(n17925), .B(n17926), .Z(n17924) );
  XNOR U18948 ( .A(n17923), .B(n8964), .Z(n17926) );
  XNOR U18949 ( .A(n17919), .B(n17921), .Z(n8964) );
  NAND U18950 ( .A(n17927), .B(e_input[556]), .Z(n17921) );
  NAND U18951 ( .A(n12323), .B(e_input[556]), .Z(n17927) );
  XNOR U18952 ( .A(n17917), .B(n17928), .Z(n17919) );
  XOR U18953 ( .A(n17929), .B(n17930), .Z(n17917) );
  AND U18954 ( .A(n17931), .B(n17932), .Z(n17930) );
  XNOR U18955 ( .A(n17933), .B(n17929), .Z(n17932) );
  XOR U18956 ( .A(n17934), .B(e_input[556]), .Z(n17925) );
  IV U18957 ( .A(n17923), .Z(n17934) );
  XOR U18958 ( .A(n17935), .B(n17936), .Z(n17923) );
  AND U18959 ( .A(n17937), .B(n17938), .Z(n17936) );
  XNOR U18960 ( .A(n17935), .B(n8970), .Z(n17938) );
  XNOR U18961 ( .A(n17931), .B(n17933), .Z(n8970) );
  NAND U18962 ( .A(n17939), .B(e_input[555]), .Z(n17933) );
  NAND U18963 ( .A(n12323), .B(e_input[555]), .Z(n17939) );
  XNOR U18964 ( .A(n17929), .B(n17940), .Z(n17931) );
  XOR U18965 ( .A(n17941), .B(n17942), .Z(n17929) );
  AND U18966 ( .A(n17943), .B(n17944), .Z(n17942) );
  XNOR U18967 ( .A(n17945), .B(n17941), .Z(n17944) );
  XOR U18968 ( .A(n17946), .B(e_input[555]), .Z(n17937) );
  IV U18969 ( .A(n17935), .Z(n17946) );
  XOR U18970 ( .A(n17947), .B(n17948), .Z(n17935) );
  AND U18971 ( .A(n17949), .B(n17950), .Z(n17948) );
  XNOR U18972 ( .A(n17947), .B(n8976), .Z(n17950) );
  XNOR U18973 ( .A(n17943), .B(n17945), .Z(n8976) );
  NAND U18974 ( .A(n17951), .B(e_input[554]), .Z(n17945) );
  NAND U18975 ( .A(n12323), .B(e_input[554]), .Z(n17951) );
  XNOR U18976 ( .A(n17941), .B(n17952), .Z(n17943) );
  XOR U18977 ( .A(n17953), .B(n17954), .Z(n17941) );
  AND U18978 ( .A(n17955), .B(n17956), .Z(n17954) );
  XNOR U18979 ( .A(n17957), .B(n17953), .Z(n17956) );
  XOR U18980 ( .A(n17958), .B(e_input[554]), .Z(n17949) );
  IV U18981 ( .A(n17947), .Z(n17958) );
  XOR U18982 ( .A(n17959), .B(n17960), .Z(n17947) );
  AND U18983 ( .A(n17961), .B(n17962), .Z(n17960) );
  XNOR U18984 ( .A(n17959), .B(n8982), .Z(n17962) );
  XNOR U18985 ( .A(n17955), .B(n17957), .Z(n8982) );
  NAND U18986 ( .A(n17963), .B(e_input[553]), .Z(n17957) );
  NAND U18987 ( .A(n12323), .B(e_input[553]), .Z(n17963) );
  XNOR U18988 ( .A(n17953), .B(n17964), .Z(n17955) );
  XOR U18989 ( .A(n17965), .B(n17966), .Z(n17953) );
  AND U18990 ( .A(n17967), .B(n17968), .Z(n17966) );
  XNOR U18991 ( .A(n17969), .B(n17965), .Z(n17968) );
  XOR U18992 ( .A(n17970), .B(e_input[553]), .Z(n17961) );
  IV U18993 ( .A(n17959), .Z(n17970) );
  XOR U18994 ( .A(n17971), .B(n17972), .Z(n17959) );
  AND U18995 ( .A(n17973), .B(n17974), .Z(n17972) );
  XNOR U18996 ( .A(n17971), .B(n8988), .Z(n17974) );
  XNOR U18997 ( .A(n17967), .B(n17969), .Z(n8988) );
  NAND U18998 ( .A(n17975), .B(e_input[552]), .Z(n17969) );
  NAND U18999 ( .A(n12323), .B(e_input[552]), .Z(n17975) );
  XNOR U19000 ( .A(n17965), .B(n17976), .Z(n17967) );
  XOR U19001 ( .A(n17977), .B(n17978), .Z(n17965) );
  AND U19002 ( .A(n17979), .B(n17980), .Z(n17978) );
  XNOR U19003 ( .A(n17981), .B(n17977), .Z(n17980) );
  XOR U19004 ( .A(n17982), .B(e_input[552]), .Z(n17973) );
  IV U19005 ( .A(n17971), .Z(n17982) );
  XOR U19006 ( .A(n17983), .B(n17984), .Z(n17971) );
  AND U19007 ( .A(n17985), .B(n17986), .Z(n17984) );
  XNOR U19008 ( .A(n17983), .B(n8994), .Z(n17986) );
  XNOR U19009 ( .A(n17979), .B(n17981), .Z(n8994) );
  NAND U19010 ( .A(n17987), .B(e_input[551]), .Z(n17981) );
  NAND U19011 ( .A(n12323), .B(e_input[551]), .Z(n17987) );
  XNOR U19012 ( .A(n17977), .B(n17988), .Z(n17979) );
  XOR U19013 ( .A(n17989), .B(n17990), .Z(n17977) );
  AND U19014 ( .A(n17991), .B(n17992), .Z(n17990) );
  XNOR U19015 ( .A(n17993), .B(n17989), .Z(n17992) );
  XOR U19016 ( .A(n17994), .B(e_input[551]), .Z(n17985) );
  IV U19017 ( .A(n17983), .Z(n17994) );
  XOR U19018 ( .A(n17995), .B(n17996), .Z(n17983) );
  AND U19019 ( .A(n17997), .B(n17998), .Z(n17996) );
  XNOR U19020 ( .A(n17995), .B(n9000), .Z(n17998) );
  XNOR U19021 ( .A(n17991), .B(n17993), .Z(n9000) );
  NAND U19022 ( .A(n17999), .B(e_input[550]), .Z(n17993) );
  NAND U19023 ( .A(n12323), .B(e_input[550]), .Z(n17999) );
  XNOR U19024 ( .A(n17989), .B(n18000), .Z(n17991) );
  XOR U19025 ( .A(n18001), .B(n18002), .Z(n17989) );
  AND U19026 ( .A(n18003), .B(n18004), .Z(n18002) );
  XNOR U19027 ( .A(n18005), .B(n18001), .Z(n18004) );
  XOR U19028 ( .A(n18006), .B(e_input[550]), .Z(n17997) );
  IV U19029 ( .A(n17995), .Z(n18006) );
  XOR U19030 ( .A(n18007), .B(n18008), .Z(n17995) );
  AND U19031 ( .A(n18009), .B(n18010), .Z(n18008) );
  XNOR U19032 ( .A(n18007), .B(n9006), .Z(n18010) );
  XNOR U19033 ( .A(n18003), .B(n18005), .Z(n9006) );
  NAND U19034 ( .A(n18011), .B(e_input[549]), .Z(n18005) );
  NAND U19035 ( .A(n12323), .B(e_input[549]), .Z(n18011) );
  XNOR U19036 ( .A(n18001), .B(n18012), .Z(n18003) );
  XOR U19037 ( .A(n18013), .B(n18014), .Z(n18001) );
  AND U19038 ( .A(n18015), .B(n18016), .Z(n18014) );
  XNOR U19039 ( .A(n18017), .B(n18013), .Z(n18016) );
  XOR U19040 ( .A(n18018), .B(e_input[549]), .Z(n18009) );
  IV U19041 ( .A(n18007), .Z(n18018) );
  XOR U19042 ( .A(n18019), .B(n18020), .Z(n18007) );
  AND U19043 ( .A(n18021), .B(n18022), .Z(n18020) );
  XNOR U19044 ( .A(n18019), .B(n9012), .Z(n18022) );
  XNOR U19045 ( .A(n18015), .B(n18017), .Z(n9012) );
  NAND U19046 ( .A(n18023), .B(e_input[548]), .Z(n18017) );
  NAND U19047 ( .A(n12323), .B(e_input[548]), .Z(n18023) );
  XNOR U19048 ( .A(n18013), .B(n18024), .Z(n18015) );
  XOR U19049 ( .A(n18025), .B(n18026), .Z(n18013) );
  AND U19050 ( .A(n18027), .B(n18028), .Z(n18026) );
  XNOR U19051 ( .A(n18029), .B(n18025), .Z(n18028) );
  XOR U19052 ( .A(n18030), .B(e_input[548]), .Z(n18021) );
  IV U19053 ( .A(n18019), .Z(n18030) );
  XOR U19054 ( .A(n18031), .B(n18032), .Z(n18019) );
  AND U19055 ( .A(n18033), .B(n18034), .Z(n18032) );
  XNOR U19056 ( .A(n18031), .B(n9018), .Z(n18034) );
  XNOR U19057 ( .A(n18027), .B(n18029), .Z(n9018) );
  NAND U19058 ( .A(n18035), .B(e_input[547]), .Z(n18029) );
  NAND U19059 ( .A(n12323), .B(e_input[547]), .Z(n18035) );
  XNOR U19060 ( .A(n18025), .B(n18036), .Z(n18027) );
  XOR U19061 ( .A(n18037), .B(n18038), .Z(n18025) );
  AND U19062 ( .A(n18039), .B(n18040), .Z(n18038) );
  XNOR U19063 ( .A(n18041), .B(n18037), .Z(n18040) );
  XOR U19064 ( .A(n18042), .B(e_input[547]), .Z(n18033) );
  IV U19065 ( .A(n18031), .Z(n18042) );
  XOR U19066 ( .A(n18043), .B(n18044), .Z(n18031) );
  AND U19067 ( .A(n18045), .B(n18046), .Z(n18044) );
  XNOR U19068 ( .A(n18043), .B(n9024), .Z(n18046) );
  XNOR U19069 ( .A(n18039), .B(n18041), .Z(n9024) );
  NAND U19070 ( .A(n18047), .B(e_input[546]), .Z(n18041) );
  NAND U19071 ( .A(n12323), .B(e_input[546]), .Z(n18047) );
  XNOR U19072 ( .A(n18037), .B(n18048), .Z(n18039) );
  XOR U19073 ( .A(n18049), .B(n18050), .Z(n18037) );
  AND U19074 ( .A(n18051), .B(n18052), .Z(n18050) );
  XNOR U19075 ( .A(n18053), .B(n18049), .Z(n18052) );
  XOR U19076 ( .A(n18054), .B(e_input[546]), .Z(n18045) );
  IV U19077 ( .A(n18043), .Z(n18054) );
  XOR U19078 ( .A(n18055), .B(n18056), .Z(n18043) );
  AND U19079 ( .A(n18057), .B(n18058), .Z(n18056) );
  XNOR U19080 ( .A(n18055), .B(n9030), .Z(n18058) );
  XNOR U19081 ( .A(n18051), .B(n18053), .Z(n9030) );
  NAND U19082 ( .A(n18059), .B(e_input[545]), .Z(n18053) );
  NAND U19083 ( .A(n12323), .B(e_input[545]), .Z(n18059) );
  XNOR U19084 ( .A(n18049), .B(n18060), .Z(n18051) );
  XOR U19085 ( .A(n18061), .B(n18062), .Z(n18049) );
  AND U19086 ( .A(n18063), .B(n18064), .Z(n18062) );
  XNOR U19087 ( .A(n18065), .B(n18061), .Z(n18064) );
  XOR U19088 ( .A(n18066), .B(e_input[545]), .Z(n18057) );
  IV U19089 ( .A(n18055), .Z(n18066) );
  XOR U19090 ( .A(n18067), .B(n18068), .Z(n18055) );
  AND U19091 ( .A(n18069), .B(n18070), .Z(n18068) );
  XNOR U19092 ( .A(n18067), .B(n9036), .Z(n18070) );
  XNOR U19093 ( .A(n18063), .B(n18065), .Z(n9036) );
  NAND U19094 ( .A(n18071), .B(e_input[544]), .Z(n18065) );
  NAND U19095 ( .A(n12323), .B(e_input[544]), .Z(n18071) );
  XNOR U19096 ( .A(n18061), .B(n18072), .Z(n18063) );
  XOR U19097 ( .A(n18073), .B(n18074), .Z(n18061) );
  AND U19098 ( .A(n18075), .B(n18076), .Z(n18074) );
  XNOR U19099 ( .A(n18077), .B(n18073), .Z(n18076) );
  XOR U19100 ( .A(n18078), .B(e_input[544]), .Z(n18069) );
  IV U19101 ( .A(n18067), .Z(n18078) );
  XOR U19102 ( .A(n18079), .B(n18080), .Z(n18067) );
  AND U19103 ( .A(n18081), .B(n18082), .Z(n18080) );
  XNOR U19104 ( .A(n18079), .B(n9042), .Z(n18082) );
  XNOR U19105 ( .A(n18075), .B(n18077), .Z(n9042) );
  NAND U19106 ( .A(n18083), .B(e_input[543]), .Z(n18077) );
  NAND U19107 ( .A(n12323), .B(e_input[543]), .Z(n18083) );
  XNOR U19108 ( .A(n18073), .B(n18084), .Z(n18075) );
  XOR U19109 ( .A(n18085), .B(n18086), .Z(n18073) );
  AND U19110 ( .A(n18087), .B(n18088), .Z(n18086) );
  XNOR U19111 ( .A(n18089), .B(n18085), .Z(n18088) );
  XOR U19112 ( .A(n18090), .B(e_input[543]), .Z(n18081) );
  IV U19113 ( .A(n18079), .Z(n18090) );
  XOR U19114 ( .A(n18091), .B(n18092), .Z(n18079) );
  AND U19115 ( .A(n18093), .B(n18094), .Z(n18092) );
  XNOR U19116 ( .A(n18091), .B(n9048), .Z(n18094) );
  XNOR U19117 ( .A(n18087), .B(n18089), .Z(n9048) );
  NAND U19118 ( .A(n18095), .B(e_input[542]), .Z(n18089) );
  NAND U19119 ( .A(n12323), .B(e_input[542]), .Z(n18095) );
  XNOR U19120 ( .A(n18085), .B(n18096), .Z(n18087) );
  XOR U19121 ( .A(n18097), .B(n18098), .Z(n18085) );
  AND U19122 ( .A(n18099), .B(n18100), .Z(n18098) );
  XNOR U19123 ( .A(n18101), .B(n18097), .Z(n18100) );
  XOR U19124 ( .A(n18102), .B(e_input[542]), .Z(n18093) );
  IV U19125 ( .A(n18091), .Z(n18102) );
  XOR U19126 ( .A(n18103), .B(n18104), .Z(n18091) );
  AND U19127 ( .A(n18105), .B(n18106), .Z(n18104) );
  XNOR U19128 ( .A(n18103), .B(n9054), .Z(n18106) );
  XNOR U19129 ( .A(n18099), .B(n18101), .Z(n9054) );
  NAND U19130 ( .A(n18107), .B(e_input[541]), .Z(n18101) );
  NAND U19131 ( .A(n12323), .B(e_input[541]), .Z(n18107) );
  XNOR U19132 ( .A(n18097), .B(n18108), .Z(n18099) );
  XOR U19133 ( .A(n18109), .B(n18110), .Z(n18097) );
  AND U19134 ( .A(n18111), .B(n18112), .Z(n18110) );
  XNOR U19135 ( .A(n18113), .B(n18109), .Z(n18112) );
  XOR U19136 ( .A(n18114), .B(e_input[541]), .Z(n18105) );
  IV U19137 ( .A(n18103), .Z(n18114) );
  XOR U19138 ( .A(n18115), .B(n18116), .Z(n18103) );
  AND U19139 ( .A(n18117), .B(n18118), .Z(n18116) );
  XNOR U19140 ( .A(n18115), .B(n9060), .Z(n18118) );
  XNOR U19141 ( .A(n18111), .B(n18113), .Z(n9060) );
  NAND U19142 ( .A(n18119), .B(e_input[540]), .Z(n18113) );
  NAND U19143 ( .A(n12323), .B(e_input[540]), .Z(n18119) );
  XNOR U19144 ( .A(n18109), .B(n18120), .Z(n18111) );
  XOR U19145 ( .A(n18121), .B(n18122), .Z(n18109) );
  AND U19146 ( .A(n18123), .B(n18124), .Z(n18122) );
  XNOR U19147 ( .A(n18125), .B(n18121), .Z(n18124) );
  XOR U19148 ( .A(n18126), .B(e_input[540]), .Z(n18117) );
  IV U19149 ( .A(n18115), .Z(n18126) );
  XOR U19150 ( .A(n18127), .B(n18128), .Z(n18115) );
  AND U19151 ( .A(n18129), .B(n18130), .Z(n18128) );
  XNOR U19152 ( .A(n18127), .B(n9066), .Z(n18130) );
  XNOR U19153 ( .A(n18123), .B(n18125), .Z(n9066) );
  NAND U19154 ( .A(n18131), .B(e_input[539]), .Z(n18125) );
  NAND U19155 ( .A(n12323), .B(e_input[539]), .Z(n18131) );
  XNOR U19156 ( .A(n18121), .B(n18132), .Z(n18123) );
  XOR U19157 ( .A(n18133), .B(n18134), .Z(n18121) );
  AND U19158 ( .A(n18135), .B(n18136), .Z(n18134) );
  XNOR U19159 ( .A(n18137), .B(n18133), .Z(n18136) );
  XOR U19160 ( .A(n18138), .B(e_input[539]), .Z(n18129) );
  IV U19161 ( .A(n18127), .Z(n18138) );
  XOR U19162 ( .A(n18139), .B(n18140), .Z(n18127) );
  AND U19163 ( .A(n18141), .B(n18142), .Z(n18140) );
  XNOR U19164 ( .A(n18139), .B(n9072), .Z(n18142) );
  XNOR U19165 ( .A(n18135), .B(n18137), .Z(n9072) );
  NAND U19166 ( .A(n18143), .B(e_input[538]), .Z(n18137) );
  NAND U19167 ( .A(n12323), .B(e_input[538]), .Z(n18143) );
  XNOR U19168 ( .A(n18133), .B(n18144), .Z(n18135) );
  XOR U19169 ( .A(n18145), .B(n18146), .Z(n18133) );
  AND U19170 ( .A(n18147), .B(n18148), .Z(n18146) );
  XNOR U19171 ( .A(n18149), .B(n18145), .Z(n18148) );
  XOR U19172 ( .A(n18150), .B(e_input[538]), .Z(n18141) );
  IV U19173 ( .A(n18139), .Z(n18150) );
  XOR U19174 ( .A(n18151), .B(n18152), .Z(n18139) );
  AND U19175 ( .A(n18153), .B(n18154), .Z(n18152) );
  XNOR U19176 ( .A(n18151), .B(n9078), .Z(n18154) );
  XNOR U19177 ( .A(n18147), .B(n18149), .Z(n9078) );
  NAND U19178 ( .A(n18155), .B(e_input[537]), .Z(n18149) );
  NAND U19179 ( .A(n12323), .B(e_input[537]), .Z(n18155) );
  XNOR U19180 ( .A(n18145), .B(n18156), .Z(n18147) );
  XOR U19181 ( .A(n18157), .B(n18158), .Z(n18145) );
  AND U19182 ( .A(n18159), .B(n18160), .Z(n18158) );
  XNOR U19183 ( .A(n18161), .B(n18157), .Z(n18160) );
  XOR U19184 ( .A(n18162), .B(e_input[537]), .Z(n18153) );
  IV U19185 ( .A(n18151), .Z(n18162) );
  XOR U19186 ( .A(n18163), .B(n18164), .Z(n18151) );
  AND U19187 ( .A(n18165), .B(n18166), .Z(n18164) );
  XNOR U19188 ( .A(n18163), .B(n9084), .Z(n18166) );
  XNOR U19189 ( .A(n18159), .B(n18161), .Z(n9084) );
  NAND U19190 ( .A(n18167), .B(e_input[536]), .Z(n18161) );
  NAND U19191 ( .A(n12323), .B(e_input[536]), .Z(n18167) );
  XNOR U19192 ( .A(n18157), .B(n18168), .Z(n18159) );
  XOR U19193 ( .A(n18169), .B(n18170), .Z(n18157) );
  AND U19194 ( .A(n18171), .B(n18172), .Z(n18170) );
  XNOR U19195 ( .A(n18173), .B(n18169), .Z(n18172) );
  XOR U19196 ( .A(n18174), .B(e_input[536]), .Z(n18165) );
  IV U19197 ( .A(n18163), .Z(n18174) );
  XOR U19198 ( .A(n18175), .B(n18176), .Z(n18163) );
  AND U19199 ( .A(n18177), .B(n18178), .Z(n18176) );
  XNOR U19200 ( .A(n18175), .B(n9090), .Z(n18178) );
  XNOR U19201 ( .A(n18171), .B(n18173), .Z(n9090) );
  NAND U19202 ( .A(n18179), .B(e_input[535]), .Z(n18173) );
  NAND U19203 ( .A(n12323), .B(e_input[535]), .Z(n18179) );
  XNOR U19204 ( .A(n18169), .B(n18180), .Z(n18171) );
  XOR U19205 ( .A(n18181), .B(n18182), .Z(n18169) );
  AND U19206 ( .A(n18183), .B(n18184), .Z(n18182) );
  XNOR U19207 ( .A(n18185), .B(n18181), .Z(n18184) );
  XOR U19208 ( .A(n18186), .B(e_input[535]), .Z(n18177) );
  IV U19209 ( .A(n18175), .Z(n18186) );
  XOR U19210 ( .A(n18187), .B(n18188), .Z(n18175) );
  AND U19211 ( .A(n18189), .B(n18190), .Z(n18188) );
  XNOR U19212 ( .A(n18187), .B(n9096), .Z(n18190) );
  XNOR U19213 ( .A(n18183), .B(n18185), .Z(n9096) );
  NAND U19214 ( .A(n18191), .B(e_input[534]), .Z(n18185) );
  NAND U19215 ( .A(n12323), .B(e_input[534]), .Z(n18191) );
  XNOR U19216 ( .A(n18181), .B(n18192), .Z(n18183) );
  XOR U19217 ( .A(n18193), .B(n18194), .Z(n18181) );
  AND U19218 ( .A(n18195), .B(n18196), .Z(n18194) );
  XNOR U19219 ( .A(n18197), .B(n18193), .Z(n18196) );
  XOR U19220 ( .A(n18198), .B(e_input[534]), .Z(n18189) );
  IV U19221 ( .A(n18187), .Z(n18198) );
  XOR U19222 ( .A(n18199), .B(n18200), .Z(n18187) );
  AND U19223 ( .A(n18201), .B(n18202), .Z(n18200) );
  XNOR U19224 ( .A(n18199), .B(n9102), .Z(n18202) );
  XNOR U19225 ( .A(n18195), .B(n18197), .Z(n9102) );
  NAND U19226 ( .A(n18203), .B(e_input[533]), .Z(n18197) );
  NAND U19227 ( .A(n12323), .B(e_input[533]), .Z(n18203) );
  XNOR U19228 ( .A(n18193), .B(n18204), .Z(n18195) );
  XOR U19229 ( .A(n18205), .B(n18206), .Z(n18193) );
  AND U19230 ( .A(n18207), .B(n18208), .Z(n18206) );
  XNOR U19231 ( .A(n18209), .B(n18205), .Z(n18208) );
  XOR U19232 ( .A(n18210), .B(e_input[533]), .Z(n18201) );
  IV U19233 ( .A(n18199), .Z(n18210) );
  XOR U19234 ( .A(n18211), .B(n18212), .Z(n18199) );
  AND U19235 ( .A(n18213), .B(n18214), .Z(n18212) );
  XNOR U19236 ( .A(n18211), .B(n9108), .Z(n18214) );
  XNOR U19237 ( .A(n18207), .B(n18209), .Z(n9108) );
  NAND U19238 ( .A(n18215), .B(e_input[532]), .Z(n18209) );
  NAND U19239 ( .A(n12323), .B(e_input[532]), .Z(n18215) );
  XNOR U19240 ( .A(n18205), .B(n18216), .Z(n18207) );
  XOR U19241 ( .A(n18217), .B(n18218), .Z(n18205) );
  AND U19242 ( .A(n18219), .B(n18220), .Z(n18218) );
  XNOR U19243 ( .A(n18221), .B(n18217), .Z(n18220) );
  XOR U19244 ( .A(n18222), .B(e_input[532]), .Z(n18213) );
  IV U19245 ( .A(n18211), .Z(n18222) );
  XOR U19246 ( .A(n18223), .B(n18224), .Z(n18211) );
  AND U19247 ( .A(n18225), .B(n18226), .Z(n18224) );
  XNOR U19248 ( .A(n18223), .B(n9114), .Z(n18226) );
  XNOR U19249 ( .A(n18219), .B(n18221), .Z(n9114) );
  NAND U19250 ( .A(n18227), .B(e_input[531]), .Z(n18221) );
  NAND U19251 ( .A(n12323), .B(e_input[531]), .Z(n18227) );
  XNOR U19252 ( .A(n18217), .B(n18228), .Z(n18219) );
  XOR U19253 ( .A(n18229), .B(n18230), .Z(n18217) );
  AND U19254 ( .A(n18231), .B(n18232), .Z(n18230) );
  XNOR U19255 ( .A(n18233), .B(n18229), .Z(n18232) );
  XOR U19256 ( .A(n18234), .B(e_input[531]), .Z(n18225) );
  IV U19257 ( .A(n18223), .Z(n18234) );
  XOR U19258 ( .A(n18235), .B(n18236), .Z(n18223) );
  AND U19259 ( .A(n18237), .B(n18238), .Z(n18236) );
  XNOR U19260 ( .A(n18235), .B(n9120), .Z(n18238) );
  XNOR U19261 ( .A(n18231), .B(n18233), .Z(n9120) );
  NAND U19262 ( .A(n18239), .B(e_input[530]), .Z(n18233) );
  NAND U19263 ( .A(n12323), .B(e_input[530]), .Z(n18239) );
  XNOR U19264 ( .A(n18229), .B(n18240), .Z(n18231) );
  XOR U19265 ( .A(n18241), .B(n18242), .Z(n18229) );
  AND U19266 ( .A(n18243), .B(n18244), .Z(n18242) );
  XNOR U19267 ( .A(n18245), .B(n18241), .Z(n18244) );
  XOR U19268 ( .A(n18246), .B(e_input[530]), .Z(n18237) );
  IV U19269 ( .A(n18235), .Z(n18246) );
  XOR U19270 ( .A(n18247), .B(n18248), .Z(n18235) );
  AND U19271 ( .A(n18249), .B(n18250), .Z(n18248) );
  XNOR U19272 ( .A(n18247), .B(n9126), .Z(n18250) );
  XNOR U19273 ( .A(n18243), .B(n18245), .Z(n9126) );
  NAND U19274 ( .A(n18251), .B(e_input[529]), .Z(n18245) );
  NAND U19275 ( .A(n12323), .B(e_input[529]), .Z(n18251) );
  XNOR U19276 ( .A(n18241), .B(n18252), .Z(n18243) );
  XOR U19277 ( .A(n18253), .B(n18254), .Z(n18241) );
  AND U19278 ( .A(n18255), .B(n18256), .Z(n18254) );
  XNOR U19279 ( .A(n18257), .B(n18253), .Z(n18256) );
  XOR U19280 ( .A(n18258), .B(e_input[529]), .Z(n18249) );
  IV U19281 ( .A(n18247), .Z(n18258) );
  XOR U19282 ( .A(n18259), .B(n18260), .Z(n18247) );
  AND U19283 ( .A(n18261), .B(n18262), .Z(n18260) );
  XNOR U19284 ( .A(n18259), .B(n9132), .Z(n18262) );
  XNOR U19285 ( .A(n18255), .B(n18257), .Z(n9132) );
  NAND U19286 ( .A(n18263), .B(e_input[528]), .Z(n18257) );
  NAND U19287 ( .A(n12323), .B(e_input[528]), .Z(n18263) );
  XNOR U19288 ( .A(n18253), .B(n18264), .Z(n18255) );
  XOR U19289 ( .A(n18265), .B(n18266), .Z(n18253) );
  AND U19290 ( .A(n18267), .B(n18268), .Z(n18266) );
  XNOR U19291 ( .A(n18269), .B(n18265), .Z(n18268) );
  XOR U19292 ( .A(n18270), .B(e_input[528]), .Z(n18261) );
  IV U19293 ( .A(n18259), .Z(n18270) );
  XOR U19294 ( .A(n18271), .B(n18272), .Z(n18259) );
  AND U19295 ( .A(n18273), .B(n18274), .Z(n18272) );
  XNOR U19296 ( .A(n18271), .B(n9138), .Z(n18274) );
  XNOR U19297 ( .A(n18267), .B(n18269), .Z(n9138) );
  NAND U19298 ( .A(n18275), .B(e_input[527]), .Z(n18269) );
  NAND U19299 ( .A(n12323), .B(e_input[527]), .Z(n18275) );
  XNOR U19300 ( .A(n18265), .B(n18276), .Z(n18267) );
  XOR U19301 ( .A(n18277), .B(n18278), .Z(n18265) );
  AND U19302 ( .A(n18279), .B(n18280), .Z(n18278) );
  XNOR U19303 ( .A(n18281), .B(n18277), .Z(n18280) );
  XOR U19304 ( .A(n18282), .B(e_input[527]), .Z(n18273) );
  IV U19305 ( .A(n18271), .Z(n18282) );
  XOR U19306 ( .A(n18283), .B(n18284), .Z(n18271) );
  AND U19307 ( .A(n18285), .B(n18286), .Z(n18284) );
  XNOR U19308 ( .A(n18283), .B(n9144), .Z(n18286) );
  XNOR U19309 ( .A(n18279), .B(n18281), .Z(n9144) );
  NAND U19310 ( .A(n18287), .B(e_input[526]), .Z(n18281) );
  NAND U19311 ( .A(n12323), .B(e_input[526]), .Z(n18287) );
  XNOR U19312 ( .A(n18277), .B(n18288), .Z(n18279) );
  XOR U19313 ( .A(n18289), .B(n18290), .Z(n18277) );
  AND U19314 ( .A(n18291), .B(n18292), .Z(n18290) );
  XNOR U19315 ( .A(n18293), .B(n18289), .Z(n18292) );
  XOR U19316 ( .A(n18294), .B(e_input[526]), .Z(n18285) );
  IV U19317 ( .A(n18283), .Z(n18294) );
  XOR U19318 ( .A(n18295), .B(n18296), .Z(n18283) );
  AND U19319 ( .A(n18297), .B(n18298), .Z(n18296) );
  XNOR U19320 ( .A(n18295), .B(n9150), .Z(n18298) );
  XNOR U19321 ( .A(n18291), .B(n18293), .Z(n9150) );
  NAND U19322 ( .A(n18299), .B(e_input[525]), .Z(n18293) );
  NAND U19323 ( .A(n12323), .B(e_input[525]), .Z(n18299) );
  XNOR U19324 ( .A(n18289), .B(n18300), .Z(n18291) );
  XOR U19325 ( .A(n18301), .B(n18302), .Z(n18289) );
  AND U19326 ( .A(n18303), .B(n18304), .Z(n18302) );
  XNOR U19327 ( .A(n18305), .B(n18301), .Z(n18304) );
  XOR U19328 ( .A(n18306), .B(e_input[525]), .Z(n18297) );
  IV U19329 ( .A(n18295), .Z(n18306) );
  XOR U19330 ( .A(n18307), .B(n18308), .Z(n18295) );
  AND U19331 ( .A(n18309), .B(n18310), .Z(n18308) );
  XNOR U19332 ( .A(n18307), .B(n9156), .Z(n18310) );
  XNOR U19333 ( .A(n18303), .B(n18305), .Z(n9156) );
  NAND U19334 ( .A(n18311), .B(e_input[524]), .Z(n18305) );
  NAND U19335 ( .A(n12323), .B(e_input[524]), .Z(n18311) );
  XNOR U19336 ( .A(n18301), .B(n18312), .Z(n18303) );
  XOR U19337 ( .A(n18313), .B(n18314), .Z(n18301) );
  AND U19338 ( .A(n18315), .B(n18316), .Z(n18314) );
  XNOR U19339 ( .A(n18317), .B(n18313), .Z(n18316) );
  XOR U19340 ( .A(n18318), .B(e_input[524]), .Z(n18309) );
  IV U19341 ( .A(n18307), .Z(n18318) );
  XOR U19342 ( .A(n18319), .B(n18320), .Z(n18307) );
  AND U19343 ( .A(n18321), .B(n18322), .Z(n18320) );
  XNOR U19344 ( .A(n18319), .B(n9162), .Z(n18322) );
  XNOR U19345 ( .A(n18315), .B(n18317), .Z(n9162) );
  NAND U19346 ( .A(n18323), .B(e_input[523]), .Z(n18317) );
  NAND U19347 ( .A(n12323), .B(e_input[523]), .Z(n18323) );
  XNOR U19348 ( .A(n18313), .B(n18324), .Z(n18315) );
  XOR U19349 ( .A(n18325), .B(n18326), .Z(n18313) );
  AND U19350 ( .A(n18327), .B(n18328), .Z(n18326) );
  XNOR U19351 ( .A(n18329), .B(n18325), .Z(n18328) );
  XOR U19352 ( .A(n18330), .B(e_input[523]), .Z(n18321) );
  IV U19353 ( .A(n18319), .Z(n18330) );
  XOR U19354 ( .A(n18331), .B(n18332), .Z(n18319) );
  AND U19355 ( .A(n18333), .B(n18334), .Z(n18332) );
  XNOR U19356 ( .A(n18331), .B(n9168), .Z(n18334) );
  XNOR U19357 ( .A(n18327), .B(n18329), .Z(n9168) );
  NAND U19358 ( .A(n18335), .B(e_input[522]), .Z(n18329) );
  NAND U19359 ( .A(n12323), .B(e_input[522]), .Z(n18335) );
  XNOR U19360 ( .A(n18325), .B(n18336), .Z(n18327) );
  XOR U19361 ( .A(n18337), .B(n18338), .Z(n18325) );
  AND U19362 ( .A(n18339), .B(n18340), .Z(n18338) );
  XNOR U19363 ( .A(n18341), .B(n18337), .Z(n18340) );
  XOR U19364 ( .A(n18342), .B(e_input[522]), .Z(n18333) );
  IV U19365 ( .A(n18331), .Z(n18342) );
  XOR U19366 ( .A(n18343), .B(n18344), .Z(n18331) );
  AND U19367 ( .A(n18345), .B(n18346), .Z(n18344) );
  XNOR U19368 ( .A(n18343), .B(n9174), .Z(n18346) );
  XNOR U19369 ( .A(n18339), .B(n18341), .Z(n9174) );
  NAND U19370 ( .A(n18347), .B(e_input[521]), .Z(n18341) );
  NAND U19371 ( .A(n12323), .B(e_input[521]), .Z(n18347) );
  XNOR U19372 ( .A(n18337), .B(n18348), .Z(n18339) );
  XOR U19373 ( .A(n18349), .B(n18350), .Z(n18337) );
  AND U19374 ( .A(n18351), .B(n18352), .Z(n18350) );
  XNOR U19375 ( .A(n18353), .B(n18349), .Z(n18352) );
  XOR U19376 ( .A(n18354), .B(e_input[521]), .Z(n18345) );
  IV U19377 ( .A(n18343), .Z(n18354) );
  XOR U19378 ( .A(n18355), .B(n18356), .Z(n18343) );
  AND U19379 ( .A(n18357), .B(n18358), .Z(n18356) );
  XNOR U19380 ( .A(n18355), .B(n9180), .Z(n18358) );
  XNOR U19381 ( .A(n18351), .B(n18353), .Z(n9180) );
  NAND U19382 ( .A(n18359), .B(e_input[520]), .Z(n18353) );
  NAND U19383 ( .A(n12323), .B(e_input[520]), .Z(n18359) );
  XNOR U19384 ( .A(n18349), .B(n18360), .Z(n18351) );
  XOR U19385 ( .A(n18361), .B(n18362), .Z(n18349) );
  AND U19386 ( .A(n18363), .B(n18364), .Z(n18362) );
  XNOR U19387 ( .A(n18365), .B(n18361), .Z(n18364) );
  XOR U19388 ( .A(n18366), .B(e_input[520]), .Z(n18357) );
  IV U19389 ( .A(n18355), .Z(n18366) );
  XOR U19390 ( .A(n18367), .B(n18368), .Z(n18355) );
  AND U19391 ( .A(n18369), .B(n18370), .Z(n18368) );
  XNOR U19392 ( .A(n18367), .B(n9186), .Z(n18370) );
  XNOR U19393 ( .A(n18363), .B(n18365), .Z(n9186) );
  NAND U19394 ( .A(n18371), .B(e_input[519]), .Z(n18365) );
  NAND U19395 ( .A(n12323), .B(e_input[519]), .Z(n18371) );
  XNOR U19396 ( .A(n18361), .B(n18372), .Z(n18363) );
  XOR U19397 ( .A(n18373), .B(n18374), .Z(n18361) );
  AND U19398 ( .A(n18375), .B(n18376), .Z(n18374) );
  XNOR U19399 ( .A(n18377), .B(n18373), .Z(n18376) );
  XOR U19400 ( .A(n18378), .B(e_input[519]), .Z(n18369) );
  IV U19401 ( .A(n18367), .Z(n18378) );
  XOR U19402 ( .A(n18379), .B(n18380), .Z(n18367) );
  AND U19403 ( .A(n18381), .B(n18382), .Z(n18380) );
  XNOR U19404 ( .A(n18379), .B(n9192), .Z(n18382) );
  XNOR U19405 ( .A(n18375), .B(n18377), .Z(n9192) );
  NAND U19406 ( .A(n18383), .B(e_input[518]), .Z(n18377) );
  NAND U19407 ( .A(n12323), .B(e_input[518]), .Z(n18383) );
  XNOR U19408 ( .A(n18373), .B(n18384), .Z(n18375) );
  XOR U19409 ( .A(n18385), .B(n18386), .Z(n18373) );
  AND U19410 ( .A(n18387), .B(n18388), .Z(n18386) );
  XNOR U19411 ( .A(n18389), .B(n18385), .Z(n18388) );
  XOR U19412 ( .A(n18390), .B(e_input[518]), .Z(n18381) );
  IV U19413 ( .A(n18379), .Z(n18390) );
  XOR U19414 ( .A(n18391), .B(n18392), .Z(n18379) );
  AND U19415 ( .A(n18393), .B(n18394), .Z(n18392) );
  XNOR U19416 ( .A(n18391), .B(n9198), .Z(n18394) );
  XNOR U19417 ( .A(n18387), .B(n18389), .Z(n9198) );
  NAND U19418 ( .A(n18395), .B(e_input[517]), .Z(n18389) );
  NAND U19419 ( .A(n12323), .B(e_input[517]), .Z(n18395) );
  XNOR U19420 ( .A(n18385), .B(n18396), .Z(n18387) );
  XOR U19421 ( .A(n18397), .B(n18398), .Z(n18385) );
  AND U19422 ( .A(n18399), .B(n18400), .Z(n18398) );
  XNOR U19423 ( .A(n18401), .B(n18397), .Z(n18400) );
  XOR U19424 ( .A(n18402), .B(e_input[517]), .Z(n18393) );
  IV U19425 ( .A(n18391), .Z(n18402) );
  XOR U19426 ( .A(n18403), .B(n18404), .Z(n18391) );
  AND U19427 ( .A(n18405), .B(n18406), .Z(n18404) );
  XNOR U19428 ( .A(n18403), .B(n9204), .Z(n18406) );
  XNOR U19429 ( .A(n18399), .B(n18401), .Z(n9204) );
  NAND U19430 ( .A(n18407), .B(e_input[516]), .Z(n18401) );
  NAND U19431 ( .A(n12323), .B(e_input[516]), .Z(n18407) );
  XNOR U19432 ( .A(n18397), .B(n18408), .Z(n18399) );
  XOR U19433 ( .A(n18409), .B(n18410), .Z(n18397) );
  AND U19434 ( .A(n18411), .B(n18412), .Z(n18410) );
  XNOR U19435 ( .A(n18413), .B(n18409), .Z(n18412) );
  XOR U19436 ( .A(n18414), .B(e_input[516]), .Z(n18405) );
  IV U19437 ( .A(n18403), .Z(n18414) );
  XOR U19438 ( .A(n18415), .B(n18416), .Z(n18403) );
  AND U19439 ( .A(n18417), .B(n18418), .Z(n18416) );
  XNOR U19440 ( .A(n18415), .B(n9210), .Z(n18418) );
  XNOR U19441 ( .A(n18411), .B(n18413), .Z(n9210) );
  NAND U19442 ( .A(n18419), .B(e_input[515]), .Z(n18413) );
  NAND U19443 ( .A(n12323), .B(e_input[515]), .Z(n18419) );
  XNOR U19444 ( .A(n18409), .B(n18420), .Z(n18411) );
  XOR U19445 ( .A(n18421), .B(n18422), .Z(n18409) );
  AND U19446 ( .A(n18423), .B(n18424), .Z(n18422) );
  XNOR U19447 ( .A(n18425), .B(n18421), .Z(n18424) );
  XOR U19448 ( .A(n18426), .B(e_input[515]), .Z(n18417) );
  IV U19449 ( .A(n18415), .Z(n18426) );
  XOR U19450 ( .A(n18427), .B(n18428), .Z(n18415) );
  AND U19451 ( .A(n18429), .B(n18430), .Z(n18428) );
  XNOR U19452 ( .A(n18427), .B(n9216), .Z(n18430) );
  XNOR U19453 ( .A(n18423), .B(n18425), .Z(n9216) );
  NAND U19454 ( .A(n18431), .B(e_input[514]), .Z(n18425) );
  NAND U19455 ( .A(n12323), .B(e_input[514]), .Z(n18431) );
  XNOR U19456 ( .A(n18421), .B(n18432), .Z(n18423) );
  XOR U19457 ( .A(n18433), .B(n18434), .Z(n18421) );
  AND U19458 ( .A(n18435), .B(n18436), .Z(n18434) );
  XNOR U19459 ( .A(n18437), .B(n18433), .Z(n18436) );
  XOR U19460 ( .A(n18438), .B(e_input[514]), .Z(n18429) );
  IV U19461 ( .A(n18427), .Z(n18438) );
  XOR U19462 ( .A(n18439), .B(n18440), .Z(n18427) );
  AND U19463 ( .A(n18441), .B(n18442), .Z(n18440) );
  XNOR U19464 ( .A(n18439), .B(n9222), .Z(n18442) );
  XNOR U19465 ( .A(n18435), .B(n18437), .Z(n9222) );
  NAND U19466 ( .A(n18443), .B(e_input[513]), .Z(n18437) );
  NAND U19467 ( .A(n12323), .B(e_input[513]), .Z(n18443) );
  XNOR U19468 ( .A(n18433), .B(n18444), .Z(n18435) );
  XOR U19469 ( .A(n18445), .B(n18446), .Z(n18433) );
  AND U19470 ( .A(n18447), .B(n18448), .Z(n18446) );
  XNOR U19471 ( .A(n18449), .B(n18445), .Z(n18448) );
  XOR U19472 ( .A(n18450), .B(e_input[513]), .Z(n18441) );
  IV U19473 ( .A(n18439), .Z(n18450) );
  XOR U19474 ( .A(n18451), .B(n18452), .Z(n18439) );
  AND U19475 ( .A(n18453), .B(n18454), .Z(n18452) );
  XNOR U19476 ( .A(n18451), .B(n9228), .Z(n18454) );
  XNOR U19477 ( .A(n18447), .B(n18449), .Z(n9228) );
  NAND U19478 ( .A(n18455), .B(e_input[512]), .Z(n18449) );
  NAND U19479 ( .A(n12323), .B(e_input[512]), .Z(n18455) );
  XNOR U19480 ( .A(n18445), .B(n18456), .Z(n18447) );
  XOR U19481 ( .A(n18457), .B(n18458), .Z(n18445) );
  AND U19482 ( .A(n18459), .B(n18460), .Z(n18458) );
  XNOR U19483 ( .A(n18461), .B(n18457), .Z(n18460) );
  XOR U19484 ( .A(n18462), .B(e_input[512]), .Z(n18453) );
  IV U19485 ( .A(n18451), .Z(n18462) );
  XOR U19486 ( .A(n18463), .B(n18464), .Z(n18451) );
  AND U19487 ( .A(n18465), .B(n18466), .Z(n18464) );
  XNOR U19488 ( .A(n18463), .B(n9234), .Z(n18466) );
  XNOR U19489 ( .A(n18459), .B(n18461), .Z(n9234) );
  NAND U19490 ( .A(n18467), .B(e_input[511]), .Z(n18461) );
  NAND U19491 ( .A(n12323), .B(e_input[511]), .Z(n18467) );
  XNOR U19492 ( .A(n18457), .B(n18468), .Z(n18459) );
  XOR U19493 ( .A(n18469), .B(n18470), .Z(n18457) );
  AND U19494 ( .A(n18471), .B(n18472), .Z(n18470) );
  XNOR U19495 ( .A(n18473), .B(n18469), .Z(n18472) );
  XOR U19496 ( .A(n18474), .B(e_input[511]), .Z(n18465) );
  IV U19497 ( .A(n18463), .Z(n18474) );
  XOR U19498 ( .A(n18475), .B(n18476), .Z(n18463) );
  AND U19499 ( .A(n18477), .B(n18478), .Z(n18476) );
  XNOR U19500 ( .A(n18475), .B(n9240), .Z(n18478) );
  XNOR U19501 ( .A(n18471), .B(n18473), .Z(n9240) );
  NAND U19502 ( .A(n18479), .B(e_input[510]), .Z(n18473) );
  NAND U19503 ( .A(n12323), .B(e_input[510]), .Z(n18479) );
  XNOR U19504 ( .A(n18469), .B(n18480), .Z(n18471) );
  XOR U19505 ( .A(n18481), .B(n18482), .Z(n18469) );
  AND U19506 ( .A(n18483), .B(n18484), .Z(n18482) );
  XNOR U19507 ( .A(n18485), .B(n18481), .Z(n18484) );
  XOR U19508 ( .A(n18486), .B(e_input[510]), .Z(n18477) );
  IV U19509 ( .A(n18475), .Z(n18486) );
  XOR U19510 ( .A(n18487), .B(n18488), .Z(n18475) );
  AND U19511 ( .A(n18489), .B(n18490), .Z(n18488) );
  XNOR U19512 ( .A(n18487), .B(n9246), .Z(n18490) );
  XNOR U19513 ( .A(n18483), .B(n18485), .Z(n9246) );
  NAND U19514 ( .A(n18491), .B(e_input[509]), .Z(n18485) );
  NAND U19515 ( .A(n12323), .B(e_input[509]), .Z(n18491) );
  XNOR U19516 ( .A(n18481), .B(n18492), .Z(n18483) );
  XOR U19517 ( .A(n18493), .B(n18494), .Z(n18481) );
  AND U19518 ( .A(n18495), .B(n18496), .Z(n18494) );
  XNOR U19519 ( .A(n18497), .B(n18493), .Z(n18496) );
  XOR U19520 ( .A(n18498), .B(e_input[509]), .Z(n18489) );
  IV U19521 ( .A(n18487), .Z(n18498) );
  XOR U19522 ( .A(n18499), .B(n18500), .Z(n18487) );
  AND U19523 ( .A(n18501), .B(n18502), .Z(n18500) );
  XNOR U19524 ( .A(n18499), .B(n9252), .Z(n18502) );
  XNOR U19525 ( .A(n18495), .B(n18497), .Z(n9252) );
  NAND U19526 ( .A(n18503), .B(e_input[508]), .Z(n18497) );
  NAND U19527 ( .A(n12323), .B(e_input[508]), .Z(n18503) );
  XNOR U19528 ( .A(n18493), .B(n18504), .Z(n18495) );
  XOR U19529 ( .A(n18505), .B(n18506), .Z(n18493) );
  AND U19530 ( .A(n18507), .B(n18508), .Z(n18506) );
  XNOR U19531 ( .A(n18509), .B(n18505), .Z(n18508) );
  XOR U19532 ( .A(n18510), .B(e_input[508]), .Z(n18501) );
  IV U19533 ( .A(n18499), .Z(n18510) );
  XOR U19534 ( .A(n18511), .B(n18512), .Z(n18499) );
  AND U19535 ( .A(n18513), .B(n18514), .Z(n18512) );
  XNOR U19536 ( .A(n18511), .B(n9258), .Z(n18514) );
  XNOR U19537 ( .A(n18507), .B(n18509), .Z(n9258) );
  NAND U19538 ( .A(n18515), .B(e_input[507]), .Z(n18509) );
  NAND U19539 ( .A(n12323), .B(e_input[507]), .Z(n18515) );
  XNOR U19540 ( .A(n18505), .B(n18516), .Z(n18507) );
  XOR U19541 ( .A(n18517), .B(n18518), .Z(n18505) );
  AND U19542 ( .A(n18519), .B(n18520), .Z(n18518) );
  XNOR U19543 ( .A(n18521), .B(n18517), .Z(n18520) );
  XOR U19544 ( .A(n18522), .B(e_input[507]), .Z(n18513) );
  IV U19545 ( .A(n18511), .Z(n18522) );
  XOR U19546 ( .A(n18523), .B(n18524), .Z(n18511) );
  AND U19547 ( .A(n18525), .B(n18526), .Z(n18524) );
  XNOR U19548 ( .A(n18523), .B(n9264), .Z(n18526) );
  XNOR U19549 ( .A(n18519), .B(n18521), .Z(n9264) );
  NAND U19550 ( .A(n18527), .B(e_input[506]), .Z(n18521) );
  NAND U19551 ( .A(n12323), .B(e_input[506]), .Z(n18527) );
  XNOR U19552 ( .A(n18517), .B(n18528), .Z(n18519) );
  XOR U19553 ( .A(n18529), .B(n18530), .Z(n18517) );
  AND U19554 ( .A(n18531), .B(n18532), .Z(n18530) );
  XNOR U19555 ( .A(n18533), .B(n18529), .Z(n18532) );
  XOR U19556 ( .A(n18534), .B(e_input[506]), .Z(n18525) );
  IV U19557 ( .A(n18523), .Z(n18534) );
  XOR U19558 ( .A(n18535), .B(n18536), .Z(n18523) );
  AND U19559 ( .A(n18537), .B(n18538), .Z(n18536) );
  XNOR U19560 ( .A(n18535), .B(n9270), .Z(n18538) );
  XNOR U19561 ( .A(n18531), .B(n18533), .Z(n9270) );
  NAND U19562 ( .A(n18539), .B(e_input[505]), .Z(n18533) );
  NAND U19563 ( .A(n12323), .B(e_input[505]), .Z(n18539) );
  XNOR U19564 ( .A(n18529), .B(n18540), .Z(n18531) );
  XOR U19565 ( .A(n18541), .B(n18542), .Z(n18529) );
  AND U19566 ( .A(n18543), .B(n18544), .Z(n18542) );
  XNOR U19567 ( .A(n18545), .B(n18541), .Z(n18544) );
  XOR U19568 ( .A(n18546), .B(e_input[505]), .Z(n18537) );
  IV U19569 ( .A(n18535), .Z(n18546) );
  XOR U19570 ( .A(n18547), .B(n18548), .Z(n18535) );
  AND U19571 ( .A(n18549), .B(n18550), .Z(n18548) );
  XNOR U19572 ( .A(n18547), .B(n9276), .Z(n18550) );
  XNOR U19573 ( .A(n18543), .B(n18545), .Z(n9276) );
  NAND U19574 ( .A(n18551), .B(e_input[504]), .Z(n18545) );
  NAND U19575 ( .A(n12323), .B(e_input[504]), .Z(n18551) );
  XNOR U19576 ( .A(n18541), .B(n18552), .Z(n18543) );
  XOR U19577 ( .A(n18553), .B(n18554), .Z(n18541) );
  AND U19578 ( .A(n18555), .B(n18556), .Z(n18554) );
  XNOR U19579 ( .A(n18557), .B(n18553), .Z(n18556) );
  XOR U19580 ( .A(n18558), .B(e_input[504]), .Z(n18549) );
  IV U19581 ( .A(n18547), .Z(n18558) );
  XOR U19582 ( .A(n18559), .B(n18560), .Z(n18547) );
  AND U19583 ( .A(n18561), .B(n18562), .Z(n18560) );
  XNOR U19584 ( .A(n18559), .B(n9282), .Z(n18562) );
  XNOR U19585 ( .A(n18555), .B(n18557), .Z(n9282) );
  NAND U19586 ( .A(n18563), .B(e_input[503]), .Z(n18557) );
  NAND U19587 ( .A(n12323), .B(e_input[503]), .Z(n18563) );
  XNOR U19588 ( .A(n18553), .B(n18564), .Z(n18555) );
  XOR U19589 ( .A(n18565), .B(n18566), .Z(n18553) );
  AND U19590 ( .A(n18567), .B(n18568), .Z(n18566) );
  XNOR U19591 ( .A(n18569), .B(n18565), .Z(n18568) );
  XOR U19592 ( .A(n18570), .B(e_input[503]), .Z(n18561) );
  IV U19593 ( .A(n18559), .Z(n18570) );
  XOR U19594 ( .A(n18571), .B(n18572), .Z(n18559) );
  AND U19595 ( .A(n18573), .B(n18574), .Z(n18572) );
  XNOR U19596 ( .A(n18571), .B(n9288), .Z(n18574) );
  XNOR U19597 ( .A(n18567), .B(n18569), .Z(n9288) );
  NAND U19598 ( .A(n18575), .B(e_input[502]), .Z(n18569) );
  NAND U19599 ( .A(n12323), .B(e_input[502]), .Z(n18575) );
  XNOR U19600 ( .A(n18565), .B(n18576), .Z(n18567) );
  XOR U19601 ( .A(n18577), .B(n18578), .Z(n18565) );
  AND U19602 ( .A(n18579), .B(n18580), .Z(n18578) );
  XNOR U19603 ( .A(n18581), .B(n18577), .Z(n18580) );
  XOR U19604 ( .A(n18582), .B(e_input[502]), .Z(n18573) );
  IV U19605 ( .A(n18571), .Z(n18582) );
  XOR U19606 ( .A(n18583), .B(n18584), .Z(n18571) );
  AND U19607 ( .A(n18585), .B(n18586), .Z(n18584) );
  XNOR U19608 ( .A(n18583), .B(n9294), .Z(n18586) );
  XNOR U19609 ( .A(n18579), .B(n18581), .Z(n9294) );
  NAND U19610 ( .A(n18587), .B(e_input[501]), .Z(n18581) );
  NAND U19611 ( .A(n12323), .B(e_input[501]), .Z(n18587) );
  XNOR U19612 ( .A(n18577), .B(n18588), .Z(n18579) );
  XOR U19613 ( .A(n18589), .B(n18590), .Z(n18577) );
  AND U19614 ( .A(n18591), .B(n18592), .Z(n18590) );
  XNOR U19615 ( .A(n18593), .B(n18589), .Z(n18592) );
  XOR U19616 ( .A(n18594), .B(e_input[501]), .Z(n18585) );
  IV U19617 ( .A(n18583), .Z(n18594) );
  XOR U19618 ( .A(n18595), .B(n18596), .Z(n18583) );
  AND U19619 ( .A(n18597), .B(n18598), .Z(n18596) );
  XNOR U19620 ( .A(n18595), .B(n9300), .Z(n18598) );
  XNOR U19621 ( .A(n18591), .B(n18593), .Z(n9300) );
  NAND U19622 ( .A(n18599), .B(e_input[500]), .Z(n18593) );
  NAND U19623 ( .A(n12323), .B(e_input[500]), .Z(n18599) );
  XNOR U19624 ( .A(n18589), .B(n18600), .Z(n18591) );
  XOR U19625 ( .A(n18601), .B(n18602), .Z(n18589) );
  AND U19626 ( .A(n18603), .B(n18604), .Z(n18602) );
  XNOR U19627 ( .A(n18605), .B(n18601), .Z(n18604) );
  XOR U19628 ( .A(n18606), .B(e_input[500]), .Z(n18597) );
  IV U19629 ( .A(n18595), .Z(n18606) );
  XOR U19630 ( .A(n18607), .B(n18608), .Z(n18595) );
  AND U19631 ( .A(n18609), .B(n18610), .Z(n18608) );
  XNOR U19632 ( .A(n18607), .B(n9306), .Z(n18610) );
  XNOR U19633 ( .A(n18603), .B(n18605), .Z(n9306) );
  NAND U19634 ( .A(n18611), .B(e_input[499]), .Z(n18605) );
  NAND U19635 ( .A(n12323), .B(e_input[499]), .Z(n18611) );
  XNOR U19636 ( .A(n18601), .B(n18612), .Z(n18603) );
  XOR U19637 ( .A(n18613), .B(n18614), .Z(n18601) );
  AND U19638 ( .A(n18615), .B(n18616), .Z(n18614) );
  XNOR U19639 ( .A(n18617), .B(n18613), .Z(n18616) );
  XOR U19640 ( .A(n18618), .B(e_input[499]), .Z(n18609) );
  IV U19641 ( .A(n18607), .Z(n18618) );
  XOR U19642 ( .A(n18619), .B(n18620), .Z(n18607) );
  AND U19643 ( .A(n18621), .B(n18622), .Z(n18620) );
  XNOR U19644 ( .A(n18619), .B(n9312), .Z(n18622) );
  XNOR U19645 ( .A(n18615), .B(n18617), .Z(n9312) );
  NAND U19646 ( .A(n18623), .B(e_input[498]), .Z(n18617) );
  NAND U19647 ( .A(n12323), .B(e_input[498]), .Z(n18623) );
  XNOR U19648 ( .A(n18613), .B(n18624), .Z(n18615) );
  XOR U19649 ( .A(n18625), .B(n18626), .Z(n18613) );
  AND U19650 ( .A(n18627), .B(n18628), .Z(n18626) );
  XNOR U19651 ( .A(n18629), .B(n18625), .Z(n18628) );
  XOR U19652 ( .A(n18630), .B(e_input[498]), .Z(n18621) );
  IV U19653 ( .A(n18619), .Z(n18630) );
  XOR U19654 ( .A(n18631), .B(n18632), .Z(n18619) );
  AND U19655 ( .A(n18633), .B(n18634), .Z(n18632) );
  XNOR U19656 ( .A(n18631), .B(n9318), .Z(n18634) );
  XNOR U19657 ( .A(n18627), .B(n18629), .Z(n9318) );
  NAND U19658 ( .A(n18635), .B(e_input[497]), .Z(n18629) );
  NAND U19659 ( .A(n12323), .B(e_input[497]), .Z(n18635) );
  XNOR U19660 ( .A(n18625), .B(n18636), .Z(n18627) );
  XOR U19661 ( .A(n18637), .B(n18638), .Z(n18625) );
  AND U19662 ( .A(n18639), .B(n18640), .Z(n18638) );
  XNOR U19663 ( .A(n18641), .B(n18637), .Z(n18640) );
  XOR U19664 ( .A(n18642), .B(e_input[497]), .Z(n18633) );
  IV U19665 ( .A(n18631), .Z(n18642) );
  XOR U19666 ( .A(n18643), .B(n18644), .Z(n18631) );
  AND U19667 ( .A(n18645), .B(n18646), .Z(n18644) );
  XNOR U19668 ( .A(n18643), .B(n9324), .Z(n18646) );
  XNOR U19669 ( .A(n18639), .B(n18641), .Z(n9324) );
  NAND U19670 ( .A(n18647), .B(e_input[496]), .Z(n18641) );
  NAND U19671 ( .A(n12323), .B(e_input[496]), .Z(n18647) );
  XNOR U19672 ( .A(n18637), .B(n18648), .Z(n18639) );
  XOR U19673 ( .A(n18649), .B(n18650), .Z(n18637) );
  AND U19674 ( .A(n18651), .B(n18652), .Z(n18650) );
  XNOR U19675 ( .A(n18653), .B(n18649), .Z(n18652) );
  XOR U19676 ( .A(n18654), .B(e_input[496]), .Z(n18645) );
  IV U19677 ( .A(n18643), .Z(n18654) );
  XOR U19678 ( .A(n18655), .B(n18656), .Z(n18643) );
  AND U19679 ( .A(n18657), .B(n18658), .Z(n18656) );
  XNOR U19680 ( .A(n18655), .B(n9330), .Z(n18658) );
  XNOR U19681 ( .A(n18651), .B(n18653), .Z(n9330) );
  NAND U19682 ( .A(n18659), .B(e_input[495]), .Z(n18653) );
  NAND U19683 ( .A(n12323), .B(e_input[495]), .Z(n18659) );
  XNOR U19684 ( .A(n18649), .B(n18660), .Z(n18651) );
  XOR U19685 ( .A(n18661), .B(n18662), .Z(n18649) );
  AND U19686 ( .A(n18663), .B(n18664), .Z(n18662) );
  XNOR U19687 ( .A(n18665), .B(n18661), .Z(n18664) );
  XOR U19688 ( .A(n18666), .B(e_input[495]), .Z(n18657) );
  IV U19689 ( .A(n18655), .Z(n18666) );
  XOR U19690 ( .A(n18667), .B(n18668), .Z(n18655) );
  AND U19691 ( .A(n18669), .B(n18670), .Z(n18668) );
  XNOR U19692 ( .A(n18667), .B(n9336), .Z(n18670) );
  XNOR U19693 ( .A(n18663), .B(n18665), .Z(n9336) );
  NAND U19694 ( .A(n18671), .B(e_input[494]), .Z(n18665) );
  NAND U19695 ( .A(n12323), .B(e_input[494]), .Z(n18671) );
  XNOR U19696 ( .A(n18661), .B(n18672), .Z(n18663) );
  XOR U19697 ( .A(n18673), .B(n18674), .Z(n18661) );
  AND U19698 ( .A(n18675), .B(n18676), .Z(n18674) );
  XNOR U19699 ( .A(n18677), .B(n18673), .Z(n18676) );
  XOR U19700 ( .A(n18678), .B(e_input[494]), .Z(n18669) );
  IV U19701 ( .A(n18667), .Z(n18678) );
  XOR U19702 ( .A(n18679), .B(n18680), .Z(n18667) );
  AND U19703 ( .A(n18681), .B(n18682), .Z(n18680) );
  XNOR U19704 ( .A(n18679), .B(n9342), .Z(n18682) );
  XNOR U19705 ( .A(n18675), .B(n18677), .Z(n9342) );
  NAND U19706 ( .A(n18683), .B(e_input[493]), .Z(n18677) );
  NAND U19707 ( .A(n12323), .B(e_input[493]), .Z(n18683) );
  XNOR U19708 ( .A(n18673), .B(n18684), .Z(n18675) );
  XOR U19709 ( .A(n18685), .B(n18686), .Z(n18673) );
  AND U19710 ( .A(n18687), .B(n18688), .Z(n18686) );
  XNOR U19711 ( .A(n18689), .B(n18685), .Z(n18688) );
  XOR U19712 ( .A(n18690), .B(e_input[493]), .Z(n18681) );
  IV U19713 ( .A(n18679), .Z(n18690) );
  XOR U19714 ( .A(n18691), .B(n18692), .Z(n18679) );
  AND U19715 ( .A(n18693), .B(n18694), .Z(n18692) );
  XNOR U19716 ( .A(n18691), .B(n9348), .Z(n18694) );
  XNOR U19717 ( .A(n18687), .B(n18689), .Z(n9348) );
  NAND U19718 ( .A(n18695), .B(e_input[492]), .Z(n18689) );
  NAND U19719 ( .A(n12323), .B(e_input[492]), .Z(n18695) );
  XNOR U19720 ( .A(n18685), .B(n18696), .Z(n18687) );
  XOR U19721 ( .A(n18697), .B(n18698), .Z(n18685) );
  AND U19722 ( .A(n18699), .B(n18700), .Z(n18698) );
  XNOR U19723 ( .A(n18701), .B(n18697), .Z(n18700) );
  XOR U19724 ( .A(n18702), .B(e_input[492]), .Z(n18693) );
  IV U19725 ( .A(n18691), .Z(n18702) );
  XOR U19726 ( .A(n18703), .B(n18704), .Z(n18691) );
  AND U19727 ( .A(n18705), .B(n18706), .Z(n18704) );
  XNOR U19728 ( .A(n18703), .B(n9354), .Z(n18706) );
  XNOR U19729 ( .A(n18699), .B(n18701), .Z(n9354) );
  NAND U19730 ( .A(n18707), .B(e_input[491]), .Z(n18701) );
  NAND U19731 ( .A(n12323), .B(e_input[491]), .Z(n18707) );
  XNOR U19732 ( .A(n18697), .B(n18708), .Z(n18699) );
  XOR U19733 ( .A(n18709), .B(n18710), .Z(n18697) );
  AND U19734 ( .A(n18711), .B(n18712), .Z(n18710) );
  XNOR U19735 ( .A(n18713), .B(n18709), .Z(n18712) );
  XOR U19736 ( .A(n18714), .B(e_input[491]), .Z(n18705) );
  IV U19737 ( .A(n18703), .Z(n18714) );
  XOR U19738 ( .A(n18715), .B(n18716), .Z(n18703) );
  AND U19739 ( .A(n18717), .B(n18718), .Z(n18716) );
  XNOR U19740 ( .A(n18715), .B(n9360), .Z(n18718) );
  XNOR U19741 ( .A(n18711), .B(n18713), .Z(n9360) );
  NAND U19742 ( .A(n18719), .B(e_input[490]), .Z(n18713) );
  NAND U19743 ( .A(n12323), .B(e_input[490]), .Z(n18719) );
  XNOR U19744 ( .A(n18709), .B(n18720), .Z(n18711) );
  XOR U19745 ( .A(n18721), .B(n18722), .Z(n18709) );
  AND U19746 ( .A(n18723), .B(n18724), .Z(n18722) );
  XNOR U19747 ( .A(n18725), .B(n18721), .Z(n18724) );
  XOR U19748 ( .A(n18726), .B(e_input[490]), .Z(n18717) );
  IV U19749 ( .A(n18715), .Z(n18726) );
  XOR U19750 ( .A(n18727), .B(n18728), .Z(n18715) );
  AND U19751 ( .A(n18729), .B(n18730), .Z(n18728) );
  XNOR U19752 ( .A(n18727), .B(n9366), .Z(n18730) );
  XNOR U19753 ( .A(n18723), .B(n18725), .Z(n9366) );
  NAND U19754 ( .A(n18731), .B(e_input[489]), .Z(n18725) );
  NAND U19755 ( .A(n12323), .B(e_input[489]), .Z(n18731) );
  XNOR U19756 ( .A(n18721), .B(n18732), .Z(n18723) );
  XOR U19757 ( .A(n18733), .B(n18734), .Z(n18721) );
  AND U19758 ( .A(n18735), .B(n18736), .Z(n18734) );
  XNOR U19759 ( .A(n18737), .B(n18733), .Z(n18736) );
  XOR U19760 ( .A(n18738), .B(e_input[489]), .Z(n18729) );
  IV U19761 ( .A(n18727), .Z(n18738) );
  XOR U19762 ( .A(n18739), .B(n18740), .Z(n18727) );
  AND U19763 ( .A(n18741), .B(n18742), .Z(n18740) );
  XNOR U19764 ( .A(n18739), .B(n9372), .Z(n18742) );
  XNOR U19765 ( .A(n18735), .B(n18737), .Z(n9372) );
  NAND U19766 ( .A(n18743), .B(e_input[488]), .Z(n18737) );
  NAND U19767 ( .A(n12323), .B(e_input[488]), .Z(n18743) );
  XNOR U19768 ( .A(n18733), .B(n18744), .Z(n18735) );
  XOR U19769 ( .A(n18745), .B(n18746), .Z(n18733) );
  AND U19770 ( .A(n18747), .B(n18748), .Z(n18746) );
  XNOR U19771 ( .A(n18749), .B(n18745), .Z(n18748) );
  XOR U19772 ( .A(n18750), .B(e_input[488]), .Z(n18741) );
  IV U19773 ( .A(n18739), .Z(n18750) );
  XOR U19774 ( .A(n18751), .B(n18752), .Z(n18739) );
  AND U19775 ( .A(n18753), .B(n18754), .Z(n18752) );
  XNOR U19776 ( .A(n18751), .B(n9378), .Z(n18754) );
  XNOR U19777 ( .A(n18747), .B(n18749), .Z(n9378) );
  NAND U19778 ( .A(n18755), .B(e_input[487]), .Z(n18749) );
  NAND U19779 ( .A(n12323), .B(e_input[487]), .Z(n18755) );
  XNOR U19780 ( .A(n18745), .B(n18756), .Z(n18747) );
  XOR U19781 ( .A(n18757), .B(n18758), .Z(n18745) );
  AND U19782 ( .A(n18759), .B(n18760), .Z(n18758) );
  XNOR U19783 ( .A(n18761), .B(n18757), .Z(n18760) );
  XOR U19784 ( .A(n18762), .B(e_input[487]), .Z(n18753) );
  IV U19785 ( .A(n18751), .Z(n18762) );
  XOR U19786 ( .A(n18763), .B(n18764), .Z(n18751) );
  AND U19787 ( .A(n18765), .B(n18766), .Z(n18764) );
  XNOR U19788 ( .A(n18763), .B(n9384), .Z(n18766) );
  XNOR U19789 ( .A(n18759), .B(n18761), .Z(n9384) );
  NAND U19790 ( .A(n18767), .B(e_input[486]), .Z(n18761) );
  NAND U19791 ( .A(n12323), .B(e_input[486]), .Z(n18767) );
  XNOR U19792 ( .A(n18757), .B(n18768), .Z(n18759) );
  XOR U19793 ( .A(n18769), .B(n18770), .Z(n18757) );
  AND U19794 ( .A(n18771), .B(n18772), .Z(n18770) );
  XNOR U19795 ( .A(n18773), .B(n18769), .Z(n18772) );
  XOR U19796 ( .A(n18774), .B(e_input[486]), .Z(n18765) );
  IV U19797 ( .A(n18763), .Z(n18774) );
  XOR U19798 ( .A(n18775), .B(n18776), .Z(n18763) );
  AND U19799 ( .A(n18777), .B(n18778), .Z(n18776) );
  XNOR U19800 ( .A(n18775), .B(n9390), .Z(n18778) );
  XNOR U19801 ( .A(n18771), .B(n18773), .Z(n9390) );
  NAND U19802 ( .A(n18779), .B(e_input[485]), .Z(n18773) );
  NAND U19803 ( .A(n12323), .B(e_input[485]), .Z(n18779) );
  XNOR U19804 ( .A(n18769), .B(n18780), .Z(n18771) );
  XOR U19805 ( .A(n18781), .B(n18782), .Z(n18769) );
  AND U19806 ( .A(n18783), .B(n18784), .Z(n18782) );
  XNOR U19807 ( .A(n18785), .B(n18781), .Z(n18784) );
  XOR U19808 ( .A(n18786), .B(e_input[485]), .Z(n18777) );
  IV U19809 ( .A(n18775), .Z(n18786) );
  XOR U19810 ( .A(n18787), .B(n18788), .Z(n18775) );
  AND U19811 ( .A(n18789), .B(n18790), .Z(n18788) );
  XNOR U19812 ( .A(n18787), .B(n9396), .Z(n18790) );
  XNOR U19813 ( .A(n18783), .B(n18785), .Z(n9396) );
  NAND U19814 ( .A(n18791), .B(e_input[484]), .Z(n18785) );
  NAND U19815 ( .A(n12323), .B(e_input[484]), .Z(n18791) );
  XNOR U19816 ( .A(n18781), .B(n18792), .Z(n18783) );
  XOR U19817 ( .A(n18793), .B(n18794), .Z(n18781) );
  AND U19818 ( .A(n18795), .B(n18796), .Z(n18794) );
  XNOR U19819 ( .A(n18797), .B(n18793), .Z(n18796) );
  XOR U19820 ( .A(n18798), .B(e_input[484]), .Z(n18789) );
  IV U19821 ( .A(n18787), .Z(n18798) );
  XOR U19822 ( .A(n18799), .B(n18800), .Z(n18787) );
  AND U19823 ( .A(n18801), .B(n18802), .Z(n18800) );
  XNOR U19824 ( .A(n18799), .B(n9402), .Z(n18802) );
  XNOR U19825 ( .A(n18795), .B(n18797), .Z(n9402) );
  NAND U19826 ( .A(n18803), .B(e_input[483]), .Z(n18797) );
  NAND U19827 ( .A(n12323), .B(e_input[483]), .Z(n18803) );
  XNOR U19828 ( .A(n18793), .B(n18804), .Z(n18795) );
  XOR U19829 ( .A(n18805), .B(n18806), .Z(n18793) );
  AND U19830 ( .A(n18807), .B(n18808), .Z(n18806) );
  XNOR U19831 ( .A(n18809), .B(n18805), .Z(n18808) );
  XOR U19832 ( .A(n18810), .B(e_input[483]), .Z(n18801) );
  IV U19833 ( .A(n18799), .Z(n18810) );
  XOR U19834 ( .A(n18811), .B(n18812), .Z(n18799) );
  AND U19835 ( .A(n18813), .B(n18814), .Z(n18812) );
  XNOR U19836 ( .A(n18811), .B(n9408), .Z(n18814) );
  XNOR U19837 ( .A(n18807), .B(n18809), .Z(n9408) );
  NAND U19838 ( .A(n18815), .B(e_input[482]), .Z(n18809) );
  NAND U19839 ( .A(n12323), .B(e_input[482]), .Z(n18815) );
  XNOR U19840 ( .A(n18805), .B(n18816), .Z(n18807) );
  XOR U19841 ( .A(n18817), .B(n18818), .Z(n18805) );
  AND U19842 ( .A(n18819), .B(n18820), .Z(n18818) );
  XNOR U19843 ( .A(n18821), .B(n18817), .Z(n18820) );
  XOR U19844 ( .A(n18822), .B(e_input[482]), .Z(n18813) );
  IV U19845 ( .A(n18811), .Z(n18822) );
  XOR U19846 ( .A(n18823), .B(n18824), .Z(n18811) );
  AND U19847 ( .A(n18825), .B(n18826), .Z(n18824) );
  XNOR U19848 ( .A(n18823), .B(n9414), .Z(n18826) );
  XNOR U19849 ( .A(n18819), .B(n18821), .Z(n9414) );
  NAND U19850 ( .A(n18827), .B(e_input[481]), .Z(n18821) );
  NAND U19851 ( .A(n12323), .B(e_input[481]), .Z(n18827) );
  XNOR U19852 ( .A(n18817), .B(n18828), .Z(n18819) );
  XOR U19853 ( .A(n18829), .B(n18830), .Z(n18817) );
  AND U19854 ( .A(n18831), .B(n18832), .Z(n18830) );
  XNOR U19855 ( .A(n18833), .B(n18829), .Z(n18832) );
  XOR U19856 ( .A(n18834), .B(e_input[481]), .Z(n18825) );
  IV U19857 ( .A(n18823), .Z(n18834) );
  XOR U19858 ( .A(n18835), .B(n18836), .Z(n18823) );
  AND U19859 ( .A(n18837), .B(n18838), .Z(n18836) );
  XNOR U19860 ( .A(n18835), .B(n9420), .Z(n18838) );
  XNOR U19861 ( .A(n18831), .B(n18833), .Z(n9420) );
  NAND U19862 ( .A(n18839), .B(e_input[480]), .Z(n18833) );
  NAND U19863 ( .A(n12323), .B(e_input[480]), .Z(n18839) );
  XNOR U19864 ( .A(n18829), .B(n18840), .Z(n18831) );
  XOR U19865 ( .A(n18841), .B(n18842), .Z(n18829) );
  AND U19866 ( .A(n18843), .B(n18844), .Z(n18842) );
  XNOR U19867 ( .A(n18845), .B(n18841), .Z(n18844) );
  XOR U19868 ( .A(n18846), .B(e_input[480]), .Z(n18837) );
  IV U19869 ( .A(n18835), .Z(n18846) );
  XOR U19870 ( .A(n18847), .B(n18848), .Z(n18835) );
  AND U19871 ( .A(n18849), .B(n18850), .Z(n18848) );
  XNOR U19872 ( .A(n18847), .B(n9426), .Z(n18850) );
  XNOR U19873 ( .A(n18843), .B(n18845), .Z(n9426) );
  NAND U19874 ( .A(n18851), .B(e_input[479]), .Z(n18845) );
  NAND U19875 ( .A(n12323), .B(e_input[479]), .Z(n18851) );
  XNOR U19876 ( .A(n18841), .B(n18852), .Z(n18843) );
  XOR U19877 ( .A(n18853), .B(n18854), .Z(n18841) );
  AND U19878 ( .A(n18855), .B(n18856), .Z(n18854) );
  XNOR U19879 ( .A(n18857), .B(n18853), .Z(n18856) );
  XOR U19880 ( .A(n18858), .B(e_input[479]), .Z(n18849) );
  IV U19881 ( .A(n18847), .Z(n18858) );
  XOR U19882 ( .A(n18859), .B(n18860), .Z(n18847) );
  AND U19883 ( .A(n18861), .B(n18862), .Z(n18860) );
  XNOR U19884 ( .A(n18859), .B(n9432), .Z(n18862) );
  XNOR U19885 ( .A(n18855), .B(n18857), .Z(n9432) );
  NAND U19886 ( .A(n18863), .B(e_input[478]), .Z(n18857) );
  NAND U19887 ( .A(n12323), .B(e_input[478]), .Z(n18863) );
  XNOR U19888 ( .A(n18853), .B(n18864), .Z(n18855) );
  XOR U19889 ( .A(n18865), .B(n18866), .Z(n18853) );
  AND U19890 ( .A(n18867), .B(n18868), .Z(n18866) );
  XNOR U19891 ( .A(n18869), .B(n18865), .Z(n18868) );
  XOR U19892 ( .A(n18870), .B(e_input[478]), .Z(n18861) );
  IV U19893 ( .A(n18859), .Z(n18870) );
  XOR U19894 ( .A(n18871), .B(n18872), .Z(n18859) );
  AND U19895 ( .A(n18873), .B(n18874), .Z(n18872) );
  XNOR U19896 ( .A(n18871), .B(n9438), .Z(n18874) );
  XNOR U19897 ( .A(n18867), .B(n18869), .Z(n9438) );
  NAND U19898 ( .A(n18875), .B(e_input[477]), .Z(n18869) );
  NAND U19899 ( .A(n12323), .B(e_input[477]), .Z(n18875) );
  XNOR U19900 ( .A(n18865), .B(n18876), .Z(n18867) );
  XOR U19901 ( .A(n18877), .B(n18878), .Z(n18865) );
  AND U19902 ( .A(n18879), .B(n18880), .Z(n18878) );
  XNOR U19903 ( .A(n18881), .B(n18877), .Z(n18880) );
  XOR U19904 ( .A(n18882), .B(e_input[477]), .Z(n18873) );
  IV U19905 ( .A(n18871), .Z(n18882) );
  XOR U19906 ( .A(n18883), .B(n18884), .Z(n18871) );
  AND U19907 ( .A(n18885), .B(n18886), .Z(n18884) );
  XNOR U19908 ( .A(n18883), .B(n9444), .Z(n18886) );
  XNOR U19909 ( .A(n18879), .B(n18881), .Z(n9444) );
  NAND U19910 ( .A(n18887), .B(e_input[476]), .Z(n18881) );
  NAND U19911 ( .A(n12323), .B(e_input[476]), .Z(n18887) );
  XNOR U19912 ( .A(n18877), .B(n18888), .Z(n18879) );
  XOR U19913 ( .A(n18889), .B(n18890), .Z(n18877) );
  AND U19914 ( .A(n18891), .B(n18892), .Z(n18890) );
  XNOR U19915 ( .A(n18893), .B(n18889), .Z(n18892) );
  XOR U19916 ( .A(n18894), .B(e_input[476]), .Z(n18885) );
  IV U19917 ( .A(n18883), .Z(n18894) );
  XOR U19918 ( .A(n18895), .B(n18896), .Z(n18883) );
  AND U19919 ( .A(n18897), .B(n18898), .Z(n18896) );
  XNOR U19920 ( .A(n18895), .B(n9450), .Z(n18898) );
  XNOR U19921 ( .A(n18891), .B(n18893), .Z(n9450) );
  NAND U19922 ( .A(n18899), .B(e_input[475]), .Z(n18893) );
  NAND U19923 ( .A(n12323), .B(e_input[475]), .Z(n18899) );
  XNOR U19924 ( .A(n18889), .B(n18900), .Z(n18891) );
  XOR U19925 ( .A(n18901), .B(n18902), .Z(n18889) );
  AND U19926 ( .A(n18903), .B(n18904), .Z(n18902) );
  XNOR U19927 ( .A(n18905), .B(n18901), .Z(n18904) );
  XOR U19928 ( .A(n18906), .B(e_input[475]), .Z(n18897) );
  IV U19929 ( .A(n18895), .Z(n18906) );
  XOR U19930 ( .A(n18907), .B(n18908), .Z(n18895) );
  AND U19931 ( .A(n18909), .B(n18910), .Z(n18908) );
  XNOR U19932 ( .A(n18907), .B(n9456), .Z(n18910) );
  XNOR U19933 ( .A(n18903), .B(n18905), .Z(n9456) );
  NAND U19934 ( .A(n18911), .B(e_input[474]), .Z(n18905) );
  NAND U19935 ( .A(n12323), .B(e_input[474]), .Z(n18911) );
  XNOR U19936 ( .A(n18901), .B(n18912), .Z(n18903) );
  XOR U19937 ( .A(n18913), .B(n18914), .Z(n18901) );
  AND U19938 ( .A(n18915), .B(n18916), .Z(n18914) );
  XNOR U19939 ( .A(n18917), .B(n18913), .Z(n18916) );
  XOR U19940 ( .A(n18918), .B(e_input[474]), .Z(n18909) );
  IV U19941 ( .A(n18907), .Z(n18918) );
  XOR U19942 ( .A(n18919), .B(n18920), .Z(n18907) );
  AND U19943 ( .A(n18921), .B(n18922), .Z(n18920) );
  XNOR U19944 ( .A(n18919), .B(n9462), .Z(n18922) );
  XNOR U19945 ( .A(n18915), .B(n18917), .Z(n9462) );
  NAND U19946 ( .A(n18923), .B(e_input[473]), .Z(n18917) );
  NAND U19947 ( .A(n12323), .B(e_input[473]), .Z(n18923) );
  XNOR U19948 ( .A(n18913), .B(n18924), .Z(n18915) );
  XOR U19949 ( .A(n18925), .B(n18926), .Z(n18913) );
  AND U19950 ( .A(n18927), .B(n18928), .Z(n18926) );
  XNOR U19951 ( .A(n18929), .B(n18925), .Z(n18928) );
  XOR U19952 ( .A(n18930), .B(e_input[473]), .Z(n18921) );
  IV U19953 ( .A(n18919), .Z(n18930) );
  XOR U19954 ( .A(n18931), .B(n18932), .Z(n18919) );
  AND U19955 ( .A(n18933), .B(n18934), .Z(n18932) );
  XNOR U19956 ( .A(n18931), .B(n9468), .Z(n18934) );
  XNOR U19957 ( .A(n18927), .B(n18929), .Z(n9468) );
  NAND U19958 ( .A(n18935), .B(e_input[472]), .Z(n18929) );
  NAND U19959 ( .A(n12323), .B(e_input[472]), .Z(n18935) );
  XNOR U19960 ( .A(n18925), .B(n18936), .Z(n18927) );
  XOR U19961 ( .A(n18937), .B(n18938), .Z(n18925) );
  AND U19962 ( .A(n18939), .B(n18940), .Z(n18938) );
  XNOR U19963 ( .A(n18941), .B(n18937), .Z(n18940) );
  XOR U19964 ( .A(n18942), .B(e_input[472]), .Z(n18933) );
  IV U19965 ( .A(n18931), .Z(n18942) );
  XOR U19966 ( .A(n18943), .B(n18944), .Z(n18931) );
  AND U19967 ( .A(n18945), .B(n18946), .Z(n18944) );
  XNOR U19968 ( .A(n18943), .B(n9474), .Z(n18946) );
  XNOR U19969 ( .A(n18939), .B(n18941), .Z(n9474) );
  NAND U19970 ( .A(n18947), .B(e_input[471]), .Z(n18941) );
  NAND U19971 ( .A(n12323), .B(e_input[471]), .Z(n18947) );
  XNOR U19972 ( .A(n18937), .B(n18948), .Z(n18939) );
  XOR U19973 ( .A(n18949), .B(n18950), .Z(n18937) );
  AND U19974 ( .A(n18951), .B(n18952), .Z(n18950) );
  XNOR U19975 ( .A(n18953), .B(n18949), .Z(n18952) );
  XOR U19976 ( .A(n18954), .B(e_input[471]), .Z(n18945) );
  IV U19977 ( .A(n18943), .Z(n18954) );
  XOR U19978 ( .A(n18955), .B(n18956), .Z(n18943) );
  AND U19979 ( .A(n18957), .B(n18958), .Z(n18956) );
  XNOR U19980 ( .A(n18955), .B(n9480), .Z(n18958) );
  XNOR U19981 ( .A(n18951), .B(n18953), .Z(n9480) );
  NAND U19982 ( .A(n18959), .B(e_input[470]), .Z(n18953) );
  NAND U19983 ( .A(n12323), .B(e_input[470]), .Z(n18959) );
  XNOR U19984 ( .A(n18949), .B(n18960), .Z(n18951) );
  XOR U19985 ( .A(n18961), .B(n18962), .Z(n18949) );
  AND U19986 ( .A(n18963), .B(n18964), .Z(n18962) );
  XNOR U19987 ( .A(n18965), .B(n18961), .Z(n18964) );
  XOR U19988 ( .A(n18966), .B(e_input[470]), .Z(n18957) );
  IV U19989 ( .A(n18955), .Z(n18966) );
  XOR U19990 ( .A(n18967), .B(n18968), .Z(n18955) );
  AND U19991 ( .A(n18969), .B(n18970), .Z(n18968) );
  XNOR U19992 ( .A(n18967), .B(n9486), .Z(n18970) );
  XNOR U19993 ( .A(n18963), .B(n18965), .Z(n9486) );
  NAND U19994 ( .A(n18971), .B(e_input[469]), .Z(n18965) );
  NAND U19995 ( .A(n12323), .B(e_input[469]), .Z(n18971) );
  XNOR U19996 ( .A(n18961), .B(n18972), .Z(n18963) );
  XOR U19997 ( .A(n18973), .B(n18974), .Z(n18961) );
  AND U19998 ( .A(n18975), .B(n18976), .Z(n18974) );
  XNOR U19999 ( .A(n18977), .B(n18973), .Z(n18976) );
  XOR U20000 ( .A(n18978), .B(e_input[469]), .Z(n18969) );
  IV U20001 ( .A(n18967), .Z(n18978) );
  XOR U20002 ( .A(n18979), .B(n18980), .Z(n18967) );
  AND U20003 ( .A(n18981), .B(n18982), .Z(n18980) );
  XNOR U20004 ( .A(n18979), .B(n9492), .Z(n18982) );
  XNOR U20005 ( .A(n18975), .B(n18977), .Z(n9492) );
  NAND U20006 ( .A(n18983), .B(e_input[468]), .Z(n18977) );
  NAND U20007 ( .A(n12323), .B(e_input[468]), .Z(n18983) );
  XNOR U20008 ( .A(n18973), .B(n18984), .Z(n18975) );
  XOR U20009 ( .A(n18985), .B(n18986), .Z(n18973) );
  AND U20010 ( .A(n18987), .B(n18988), .Z(n18986) );
  XNOR U20011 ( .A(n18989), .B(n18985), .Z(n18988) );
  XOR U20012 ( .A(n18990), .B(e_input[468]), .Z(n18981) );
  IV U20013 ( .A(n18979), .Z(n18990) );
  XOR U20014 ( .A(n18991), .B(n18992), .Z(n18979) );
  AND U20015 ( .A(n18993), .B(n18994), .Z(n18992) );
  XNOR U20016 ( .A(n18991), .B(n9498), .Z(n18994) );
  XNOR U20017 ( .A(n18987), .B(n18989), .Z(n9498) );
  NAND U20018 ( .A(n18995), .B(e_input[467]), .Z(n18989) );
  NAND U20019 ( .A(n12323), .B(e_input[467]), .Z(n18995) );
  XNOR U20020 ( .A(n18985), .B(n18996), .Z(n18987) );
  XOR U20021 ( .A(n18997), .B(n18998), .Z(n18985) );
  AND U20022 ( .A(n18999), .B(n19000), .Z(n18998) );
  XNOR U20023 ( .A(n19001), .B(n18997), .Z(n19000) );
  XOR U20024 ( .A(n19002), .B(e_input[467]), .Z(n18993) );
  IV U20025 ( .A(n18991), .Z(n19002) );
  XOR U20026 ( .A(n19003), .B(n19004), .Z(n18991) );
  AND U20027 ( .A(n19005), .B(n19006), .Z(n19004) );
  XNOR U20028 ( .A(n19003), .B(n9504), .Z(n19006) );
  XNOR U20029 ( .A(n18999), .B(n19001), .Z(n9504) );
  NAND U20030 ( .A(n19007), .B(e_input[466]), .Z(n19001) );
  NAND U20031 ( .A(n12323), .B(e_input[466]), .Z(n19007) );
  XNOR U20032 ( .A(n18997), .B(n19008), .Z(n18999) );
  XOR U20033 ( .A(n19009), .B(n19010), .Z(n18997) );
  AND U20034 ( .A(n19011), .B(n19012), .Z(n19010) );
  XNOR U20035 ( .A(n19013), .B(n19009), .Z(n19012) );
  XOR U20036 ( .A(n19014), .B(e_input[466]), .Z(n19005) );
  IV U20037 ( .A(n19003), .Z(n19014) );
  XOR U20038 ( .A(n19015), .B(n19016), .Z(n19003) );
  AND U20039 ( .A(n19017), .B(n19018), .Z(n19016) );
  XNOR U20040 ( .A(n19015), .B(n9510), .Z(n19018) );
  XNOR U20041 ( .A(n19011), .B(n19013), .Z(n9510) );
  NAND U20042 ( .A(n19019), .B(e_input[465]), .Z(n19013) );
  NAND U20043 ( .A(n12323), .B(e_input[465]), .Z(n19019) );
  XNOR U20044 ( .A(n19009), .B(n19020), .Z(n19011) );
  XOR U20045 ( .A(n19021), .B(n19022), .Z(n19009) );
  AND U20046 ( .A(n19023), .B(n19024), .Z(n19022) );
  XNOR U20047 ( .A(n19025), .B(n19021), .Z(n19024) );
  XOR U20048 ( .A(n19026), .B(e_input[465]), .Z(n19017) );
  IV U20049 ( .A(n19015), .Z(n19026) );
  XOR U20050 ( .A(n19027), .B(n19028), .Z(n19015) );
  AND U20051 ( .A(n19029), .B(n19030), .Z(n19028) );
  XNOR U20052 ( .A(n19027), .B(n9516), .Z(n19030) );
  XNOR U20053 ( .A(n19023), .B(n19025), .Z(n9516) );
  NAND U20054 ( .A(n19031), .B(e_input[464]), .Z(n19025) );
  NAND U20055 ( .A(n12323), .B(e_input[464]), .Z(n19031) );
  XNOR U20056 ( .A(n19021), .B(n19032), .Z(n19023) );
  XOR U20057 ( .A(n19033), .B(n19034), .Z(n19021) );
  AND U20058 ( .A(n19035), .B(n19036), .Z(n19034) );
  XNOR U20059 ( .A(n19037), .B(n19033), .Z(n19036) );
  XOR U20060 ( .A(n19038), .B(e_input[464]), .Z(n19029) );
  IV U20061 ( .A(n19027), .Z(n19038) );
  XOR U20062 ( .A(n19039), .B(n19040), .Z(n19027) );
  AND U20063 ( .A(n19041), .B(n19042), .Z(n19040) );
  XNOR U20064 ( .A(n19039), .B(n9522), .Z(n19042) );
  XNOR U20065 ( .A(n19035), .B(n19037), .Z(n9522) );
  NAND U20066 ( .A(n19043), .B(e_input[463]), .Z(n19037) );
  NAND U20067 ( .A(n12323), .B(e_input[463]), .Z(n19043) );
  XNOR U20068 ( .A(n19033), .B(n19044), .Z(n19035) );
  XOR U20069 ( .A(n19045), .B(n19046), .Z(n19033) );
  AND U20070 ( .A(n19047), .B(n19048), .Z(n19046) );
  XNOR U20071 ( .A(n19049), .B(n19045), .Z(n19048) );
  XOR U20072 ( .A(n19050), .B(e_input[463]), .Z(n19041) );
  IV U20073 ( .A(n19039), .Z(n19050) );
  XOR U20074 ( .A(n19051), .B(n19052), .Z(n19039) );
  AND U20075 ( .A(n19053), .B(n19054), .Z(n19052) );
  XNOR U20076 ( .A(n19051), .B(n9528), .Z(n19054) );
  XNOR U20077 ( .A(n19047), .B(n19049), .Z(n9528) );
  NAND U20078 ( .A(n19055), .B(e_input[462]), .Z(n19049) );
  NAND U20079 ( .A(n12323), .B(e_input[462]), .Z(n19055) );
  XNOR U20080 ( .A(n19045), .B(n19056), .Z(n19047) );
  XOR U20081 ( .A(n19057), .B(n19058), .Z(n19045) );
  AND U20082 ( .A(n19059), .B(n19060), .Z(n19058) );
  XNOR U20083 ( .A(n19061), .B(n19057), .Z(n19060) );
  XOR U20084 ( .A(n19062), .B(e_input[462]), .Z(n19053) );
  IV U20085 ( .A(n19051), .Z(n19062) );
  XOR U20086 ( .A(n19063), .B(n19064), .Z(n19051) );
  AND U20087 ( .A(n19065), .B(n19066), .Z(n19064) );
  XNOR U20088 ( .A(n19063), .B(n9534), .Z(n19066) );
  XNOR U20089 ( .A(n19059), .B(n19061), .Z(n9534) );
  NAND U20090 ( .A(n19067), .B(e_input[461]), .Z(n19061) );
  NAND U20091 ( .A(n12323), .B(e_input[461]), .Z(n19067) );
  XNOR U20092 ( .A(n19057), .B(n19068), .Z(n19059) );
  XOR U20093 ( .A(n19069), .B(n19070), .Z(n19057) );
  AND U20094 ( .A(n19071), .B(n19072), .Z(n19070) );
  XNOR U20095 ( .A(n19073), .B(n19069), .Z(n19072) );
  XOR U20096 ( .A(n19074), .B(e_input[461]), .Z(n19065) );
  IV U20097 ( .A(n19063), .Z(n19074) );
  XOR U20098 ( .A(n19075), .B(n19076), .Z(n19063) );
  AND U20099 ( .A(n19077), .B(n19078), .Z(n19076) );
  XNOR U20100 ( .A(n19075), .B(n9540), .Z(n19078) );
  XNOR U20101 ( .A(n19071), .B(n19073), .Z(n9540) );
  NAND U20102 ( .A(n19079), .B(e_input[460]), .Z(n19073) );
  NAND U20103 ( .A(n12323), .B(e_input[460]), .Z(n19079) );
  XNOR U20104 ( .A(n19069), .B(n19080), .Z(n19071) );
  XOR U20105 ( .A(n19081), .B(n19082), .Z(n19069) );
  AND U20106 ( .A(n19083), .B(n19084), .Z(n19082) );
  XNOR U20107 ( .A(n19085), .B(n19081), .Z(n19084) );
  XOR U20108 ( .A(n19086), .B(e_input[460]), .Z(n19077) );
  IV U20109 ( .A(n19075), .Z(n19086) );
  XOR U20110 ( .A(n19087), .B(n19088), .Z(n19075) );
  AND U20111 ( .A(n19089), .B(n19090), .Z(n19088) );
  XNOR U20112 ( .A(n19087), .B(n9546), .Z(n19090) );
  XNOR U20113 ( .A(n19083), .B(n19085), .Z(n9546) );
  NAND U20114 ( .A(n19091), .B(e_input[459]), .Z(n19085) );
  NAND U20115 ( .A(n12323), .B(e_input[459]), .Z(n19091) );
  XNOR U20116 ( .A(n19081), .B(n19092), .Z(n19083) );
  XOR U20117 ( .A(n19093), .B(n19094), .Z(n19081) );
  AND U20118 ( .A(n19095), .B(n19096), .Z(n19094) );
  XNOR U20119 ( .A(n19097), .B(n19093), .Z(n19096) );
  XOR U20120 ( .A(n19098), .B(e_input[459]), .Z(n19089) );
  IV U20121 ( .A(n19087), .Z(n19098) );
  XOR U20122 ( .A(n19099), .B(n19100), .Z(n19087) );
  AND U20123 ( .A(n19101), .B(n19102), .Z(n19100) );
  XNOR U20124 ( .A(n19099), .B(n9552), .Z(n19102) );
  XNOR U20125 ( .A(n19095), .B(n19097), .Z(n9552) );
  NAND U20126 ( .A(n19103), .B(e_input[458]), .Z(n19097) );
  NAND U20127 ( .A(n12323), .B(e_input[458]), .Z(n19103) );
  XNOR U20128 ( .A(n19093), .B(n19104), .Z(n19095) );
  XOR U20129 ( .A(n19105), .B(n19106), .Z(n19093) );
  AND U20130 ( .A(n19107), .B(n19108), .Z(n19106) );
  XNOR U20131 ( .A(n19109), .B(n19105), .Z(n19108) );
  XOR U20132 ( .A(n19110), .B(e_input[458]), .Z(n19101) );
  IV U20133 ( .A(n19099), .Z(n19110) );
  XOR U20134 ( .A(n19111), .B(n19112), .Z(n19099) );
  AND U20135 ( .A(n19113), .B(n19114), .Z(n19112) );
  XNOR U20136 ( .A(n19111), .B(n9558), .Z(n19114) );
  XNOR U20137 ( .A(n19107), .B(n19109), .Z(n9558) );
  NAND U20138 ( .A(n19115), .B(e_input[457]), .Z(n19109) );
  NAND U20139 ( .A(n12323), .B(e_input[457]), .Z(n19115) );
  XNOR U20140 ( .A(n19105), .B(n19116), .Z(n19107) );
  XOR U20141 ( .A(n19117), .B(n19118), .Z(n19105) );
  AND U20142 ( .A(n19119), .B(n19120), .Z(n19118) );
  XNOR U20143 ( .A(n19121), .B(n19117), .Z(n19120) );
  XOR U20144 ( .A(n19122), .B(e_input[457]), .Z(n19113) );
  IV U20145 ( .A(n19111), .Z(n19122) );
  XOR U20146 ( .A(n19123), .B(n19124), .Z(n19111) );
  AND U20147 ( .A(n19125), .B(n19126), .Z(n19124) );
  XNOR U20148 ( .A(n19123), .B(n9564), .Z(n19126) );
  XNOR U20149 ( .A(n19119), .B(n19121), .Z(n9564) );
  NAND U20150 ( .A(n19127), .B(e_input[456]), .Z(n19121) );
  NAND U20151 ( .A(n12323), .B(e_input[456]), .Z(n19127) );
  XNOR U20152 ( .A(n19117), .B(n19128), .Z(n19119) );
  XOR U20153 ( .A(n19129), .B(n19130), .Z(n19117) );
  AND U20154 ( .A(n19131), .B(n19132), .Z(n19130) );
  XNOR U20155 ( .A(n19133), .B(n19129), .Z(n19132) );
  XOR U20156 ( .A(n19134), .B(e_input[456]), .Z(n19125) );
  IV U20157 ( .A(n19123), .Z(n19134) );
  XOR U20158 ( .A(n19135), .B(n19136), .Z(n19123) );
  AND U20159 ( .A(n19137), .B(n19138), .Z(n19136) );
  XNOR U20160 ( .A(n19135), .B(n9570), .Z(n19138) );
  XNOR U20161 ( .A(n19131), .B(n19133), .Z(n9570) );
  NAND U20162 ( .A(n19139), .B(e_input[455]), .Z(n19133) );
  NAND U20163 ( .A(n12323), .B(e_input[455]), .Z(n19139) );
  XNOR U20164 ( .A(n19129), .B(n19140), .Z(n19131) );
  XOR U20165 ( .A(n19141), .B(n19142), .Z(n19129) );
  AND U20166 ( .A(n19143), .B(n19144), .Z(n19142) );
  XNOR U20167 ( .A(n19145), .B(n19141), .Z(n19144) );
  XOR U20168 ( .A(n19146), .B(e_input[455]), .Z(n19137) );
  IV U20169 ( .A(n19135), .Z(n19146) );
  XOR U20170 ( .A(n19147), .B(n19148), .Z(n19135) );
  AND U20171 ( .A(n19149), .B(n19150), .Z(n19148) );
  XNOR U20172 ( .A(n19147), .B(n9576), .Z(n19150) );
  XNOR U20173 ( .A(n19143), .B(n19145), .Z(n9576) );
  NAND U20174 ( .A(n19151), .B(e_input[454]), .Z(n19145) );
  NAND U20175 ( .A(n12323), .B(e_input[454]), .Z(n19151) );
  XNOR U20176 ( .A(n19141), .B(n19152), .Z(n19143) );
  XOR U20177 ( .A(n19153), .B(n19154), .Z(n19141) );
  AND U20178 ( .A(n19155), .B(n19156), .Z(n19154) );
  XNOR U20179 ( .A(n19157), .B(n19153), .Z(n19156) );
  XOR U20180 ( .A(n19158), .B(e_input[454]), .Z(n19149) );
  IV U20181 ( .A(n19147), .Z(n19158) );
  XOR U20182 ( .A(n19159), .B(n19160), .Z(n19147) );
  AND U20183 ( .A(n19161), .B(n19162), .Z(n19160) );
  XNOR U20184 ( .A(n19159), .B(n9582), .Z(n19162) );
  XNOR U20185 ( .A(n19155), .B(n19157), .Z(n9582) );
  NAND U20186 ( .A(n19163), .B(e_input[453]), .Z(n19157) );
  NAND U20187 ( .A(n12323), .B(e_input[453]), .Z(n19163) );
  XNOR U20188 ( .A(n19153), .B(n19164), .Z(n19155) );
  XOR U20189 ( .A(n19165), .B(n19166), .Z(n19153) );
  AND U20190 ( .A(n19167), .B(n19168), .Z(n19166) );
  XNOR U20191 ( .A(n19169), .B(n19165), .Z(n19168) );
  XOR U20192 ( .A(n19170), .B(e_input[453]), .Z(n19161) );
  IV U20193 ( .A(n19159), .Z(n19170) );
  XOR U20194 ( .A(n19171), .B(n19172), .Z(n19159) );
  AND U20195 ( .A(n19173), .B(n19174), .Z(n19172) );
  XNOR U20196 ( .A(n19171), .B(n9588), .Z(n19174) );
  XNOR U20197 ( .A(n19167), .B(n19169), .Z(n9588) );
  NAND U20198 ( .A(n19175), .B(e_input[452]), .Z(n19169) );
  NAND U20199 ( .A(n12323), .B(e_input[452]), .Z(n19175) );
  XNOR U20200 ( .A(n19165), .B(n19176), .Z(n19167) );
  XOR U20201 ( .A(n19177), .B(n19178), .Z(n19165) );
  AND U20202 ( .A(n19179), .B(n19180), .Z(n19178) );
  XNOR U20203 ( .A(n19181), .B(n19177), .Z(n19180) );
  XOR U20204 ( .A(n19182), .B(e_input[452]), .Z(n19173) );
  IV U20205 ( .A(n19171), .Z(n19182) );
  XOR U20206 ( .A(n19183), .B(n19184), .Z(n19171) );
  AND U20207 ( .A(n19185), .B(n19186), .Z(n19184) );
  XNOR U20208 ( .A(n19183), .B(n9594), .Z(n19186) );
  XNOR U20209 ( .A(n19179), .B(n19181), .Z(n9594) );
  NAND U20210 ( .A(n19187), .B(e_input[451]), .Z(n19181) );
  NAND U20211 ( .A(n12323), .B(e_input[451]), .Z(n19187) );
  XNOR U20212 ( .A(n19177), .B(n19188), .Z(n19179) );
  XOR U20213 ( .A(n19189), .B(n19190), .Z(n19177) );
  AND U20214 ( .A(n19191), .B(n19192), .Z(n19190) );
  XNOR U20215 ( .A(n19193), .B(n19189), .Z(n19192) );
  XOR U20216 ( .A(n19194), .B(e_input[451]), .Z(n19185) );
  IV U20217 ( .A(n19183), .Z(n19194) );
  XOR U20218 ( .A(n19195), .B(n19196), .Z(n19183) );
  AND U20219 ( .A(n19197), .B(n19198), .Z(n19196) );
  XNOR U20220 ( .A(n19195), .B(n9600), .Z(n19198) );
  XNOR U20221 ( .A(n19191), .B(n19193), .Z(n9600) );
  NAND U20222 ( .A(n19199), .B(e_input[450]), .Z(n19193) );
  NAND U20223 ( .A(n12323), .B(e_input[450]), .Z(n19199) );
  XNOR U20224 ( .A(n19189), .B(n19200), .Z(n19191) );
  XOR U20225 ( .A(n19201), .B(n19202), .Z(n19189) );
  AND U20226 ( .A(n19203), .B(n19204), .Z(n19202) );
  XNOR U20227 ( .A(n19205), .B(n19201), .Z(n19204) );
  XOR U20228 ( .A(n19206), .B(e_input[450]), .Z(n19197) );
  IV U20229 ( .A(n19195), .Z(n19206) );
  XOR U20230 ( .A(n19207), .B(n19208), .Z(n19195) );
  AND U20231 ( .A(n19209), .B(n19210), .Z(n19208) );
  XNOR U20232 ( .A(n19207), .B(n9606), .Z(n19210) );
  XNOR U20233 ( .A(n19203), .B(n19205), .Z(n9606) );
  NAND U20234 ( .A(n19211), .B(e_input[449]), .Z(n19205) );
  NAND U20235 ( .A(n12323), .B(e_input[449]), .Z(n19211) );
  XNOR U20236 ( .A(n19201), .B(n19212), .Z(n19203) );
  XOR U20237 ( .A(n19213), .B(n19214), .Z(n19201) );
  AND U20238 ( .A(n19215), .B(n19216), .Z(n19214) );
  XNOR U20239 ( .A(n19217), .B(n19213), .Z(n19216) );
  XOR U20240 ( .A(n19218), .B(e_input[449]), .Z(n19209) );
  IV U20241 ( .A(n19207), .Z(n19218) );
  XOR U20242 ( .A(n19219), .B(n19220), .Z(n19207) );
  AND U20243 ( .A(n19221), .B(n19222), .Z(n19220) );
  XNOR U20244 ( .A(n19219), .B(n9612), .Z(n19222) );
  XNOR U20245 ( .A(n19215), .B(n19217), .Z(n9612) );
  NAND U20246 ( .A(n19223), .B(e_input[448]), .Z(n19217) );
  NAND U20247 ( .A(n12323), .B(e_input[448]), .Z(n19223) );
  XNOR U20248 ( .A(n19213), .B(n19224), .Z(n19215) );
  XOR U20249 ( .A(n19225), .B(n19226), .Z(n19213) );
  AND U20250 ( .A(n19227), .B(n19228), .Z(n19226) );
  XNOR U20251 ( .A(n19229), .B(n19225), .Z(n19228) );
  XOR U20252 ( .A(n19230), .B(e_input[448]), .Z(n19221) );
  IV U20253 ( .A(n19219), .Z(n19230) );
  XOR U20254 ( .A(n19231), .B(n19232), .Z(n19219) );
  AND U20255 ( .A(n19233), .B(n19234), .Z(n19232) );
  XNOR U20256 ( .A(n19231), .B(n9618), .Z(n19234) );
  XNOR U20257 ( .A(n19227), .B(n19229), .Z(n9618) );
  NAND U20258 ( .A(n19235), .B(e_input[447]), .Z(n19229) );
  NAND U20259 ( .A(n12323), .B(e_input[447]), .Z(n19235) );
  XNOR U20260 ( .A(n19225), .B(n19236), .Z(n19227) );
  XOR U20261 ( .A(n19237), .B(n19238), .Z(n19225) );
  AND U20262 ( .A(n19239), .B(n19240), .Z(n19238) );
  XNOR U20263 ( .A(n19241), .B(n19237), .Z(n19240) );
  XOR U20264 ( .A(n19242), .B(e_input[447]), .Z(n19233) );
  IV U20265 ( .A(n19231), .Z(n19242) );
  XOR U20266 ( .A(n19243), .B(n19244), .Z(n19231) );
  AND U20267 ( .A(n19245), .B(n19246), .Z(n19244) );
  XNOR U20268 ( .A(n19243), .B(n9624), .Z(n19246) );
  XNOR U20269 ( .A(n19239), .B(n19241), .Z(n9624) );
  NAND U20270 ( .A(n19247), .B(e_input[446]), .Z(n19241) );
  NAND U20271 ( .A(n12323), .B(e_input[446]), .Z(n19247) );
  XNOR U20272 ( .A(n19237), .B(n19248), .Z(n19239) );
  XOR U20273 ( .A(n19249), .B(n19250), .Z(n19237) );
  AND U20274 ( .A(n19251), .B(n19252), .Z(n19250) );
  XNOR U20275 ( .A(n19253), .B(n19249), .Z(n19252) );
  XOR U20276 ( .A(n19254), .B(e_input[446]), .Z(n19245) );
  IV U20277 ( .A(n19243), .Z(n19254) );
  XOR U20278 ( .A(n19255), .B(n19256), .Z(n19243) );
  AND U20279 ( .A(n19257), .B(n19258), .Z(n19256) );
  XNOR U20280 ( .A(n19255), .B(n9630), .Z(n19258) );
  XNOR U20281 ( .A(n19251), .B(n19253), .Z(n9630) );
  NAND U20282 ( .A(n19259), .B(e_input[445]), .Z(n19253) );
  NAND U20283 ( .A(n12323), .B(e_input[445]), .Z(n19259) );
  XNOR U20284 ( .A(n19249), .B(n19260), .Z(n19251) );
  XOR U20285 ( .A(n19261), .B(n19262), .Z(n19249) );
  AND U20286 ( .A(n19263), .B(n19264), .Z(n19262) );
  XNOR U20287 ( .A(n19265), .B(n19261), .Z(n19264) );
  XOR U20288 ( .A(n19266), .B(e_input[445]), .Z(n19257) );
  IV U20289 ( .A(n19255), .Z(n19266) );
  XOR U20290 ( .A(n19267), .B(n19268), .Z(n19255) );
  AND U20291 ( .A(n19269), .B(n19270), .Z(n19268) );
  XNOR U20292 ( .A(n19267), .B(n9636), .Z(n19270) );
  XNOR U20293 ( .A(n19263), .B(n19265), .Z(n9636) );
  NAND U20294 ( .A(n19271), .B(e_input[444]), .Z(n19265) );
  NAND U20295 ( .A(n12323), .B(e_input[444]), .Z(n19271) );
  XNOR U20296 ( .A(n19261), .B(n19272), .Z(n19263) );
  XOR U20297 ( .A(n19273), .B(n19274), .Z(n19261) );
  AND U20298 ( .A(n19275), .B(n19276), .Z(n19274) );
  XNOR U20299 ( .A(n19277), .B(n19273), .Z(n19276) );
  XOR U20300 ( .A(n19278), .B(e_input[444]), .Z(n19269) );
  IV U20301 ( .A(n19267), .Z(n19278) );
  XOR U20302 ( .A(n19279), .B(n19280), .Z(n19267) );
  AND U20303 ( .A(n19281), .B(n19282), .Z(n19280) );
  XNOR U20304 ( .A(n19279), .B(n9642), .Z(n19282) );
  XNOR U20305 ( .A(n19275), .B(n19277), .Z(n9642) );
  NAND U20306 ( .A(n19283), .B(e_input[443]), .Z(n19277) );
  NAND U20307 ( .A(n12323), .B(e_input[443]), .Z(n19283) );
  XNOR U20308 ( .A(n19273), .B(n19284), .Z(n19275) );
  XOR U20309 ( .A(n19285), .B(n19286), .Z(n19273) );
  AND U20310 ( .A(n19287), .B(n19288), .Z(n19286) );
  XNOR U20311 ( .A(n19289), .B(n19285), .Z(n19288) );
  XOR U20312 ( .A(n19290), .B(e_input[443]), .Z(n19281) );
  IV U20313 ( .A(n19279), .Z(n19290) );
  XOR U20314 ( .A(n19291), .B(n19292), .Z(n19279) );
  AND U20315 ( .A(n19293), .B(n19294), .Z(n19292) );
  XNOR U20316 ( .A(n19291), .B(n9648), .Z(n19294) );
  XNOR U20317 ( .A(n19287), .B(n19289), .Z(n9648) );
  NAND U20318 ( .A(n19295), .B(e_input[442]), .Z(n19289) );
  NAND U20319 ( .A(n12323), .B(e_input[442]), .Z(n19295) );
  XNOR U20320 ( .A(n19285), .B(n19296), .Z(n19287) );
  XOR U20321 ( .A(n19297), .B(n19298), .Z(n19285) );
  AND U20322 ( .A(n19299), .B(n19300), .Z(n19298) );
  XNOR U20323 ( .A(n19301), .B(n19297), .Z(n19300) );
  XOR U20324 ( .A(n19302), .B(e_input[442]), .Z(n19293) );
  IV U20325 ( .A(n19291), .Z(n19302) );
  XOR U20326 ( .A(n19303), .B(n19304), .Z(n19291) );
  AND U20327 ( .A(n19305), .B(n19306), .Z(n19304) );
  XNOR U20328 ( .A(n19303), .B(n9654), .Z(n19306) );
  XNOR U20329 ( .A(n19299), .B(n19301), .Z(n9654) );
  NAND U20330 ( .A(n19307), .B(e_input[441]), .Z(n19301) );
  NAND U20331 ( .A(n12323), .B(e_input[441]), .Z(n19307) );
  XNOR U20332 ( .A(n19297), .B(n19308), .Z(n19299) );
  XOR U20333 ( .A(n19309), .B(n19310), .Z(n19297) );
  AND U20334 ( .A(n19311), .B(n19312), .Z(n19310) );
  XNOR U20335 ( .A(n19313), .B(n19309), .Z(n19312) );
  XOR U20336 ( .A(n19314), .B(e_input[441]), .Z(n19305) );
  IV U20337 ( .A(n19303), .Z(n19314) );
  XOR U20338 ( .A(n19315), .B(n19316), .Z(n19303) );
  AND U20339 ( .A(n19317), .B(n19318), .Z(n19316) );
  XNOR U20340 ( .A(n19315), .B(n9660), .Z(n19318) );
  XNOR U20341 ( .A(n19311), .B(n19313), .Z(n9660) );
  NAND U20342 ( .A(n19319), .B(e_input[440]), .Z(n19313) );
  NAND U20343 ( .A(n12323), .B(e_input[440]), .Z(n19319) );
  XNOR U20344 ( .A(n19309), .B(n19320), .Z(n19311) );
  XOR U20345 ( .A(n19321), .B(n19322), .Z(n19309) );
  AND U20346 ( .A(n19323), .B(n19324), .Z(n19322) );
  XNOR U20347 ( .A(n19325), .B(n19321), .Z(n19324) );
  XOR U20348 ( .A(n19326), .B(e_input[440]), .Z(n19317) );
  IV U20349 ( .A(n19315), .Z(n19326) );
  XOR U20350 ( .A(n19327), .B(n19328), .Z(n19315) );
  AND U20351 ( .A(n19329), .B(n19330), .Z(n19328) );
  XNOR U20352 ( .A(n19327), .B(n9666), .Z(n19330) );
  XNOR U20353 ( .A(n19323), .B(n19325), .Z(n9666) );
  NAND U20354 ( .A(n19331), .B(e_input[439]), .Z(n19325) );
  NAND U20355 ( .A(n12323), .B(e_input[439]), .Z(n19331) );
  XNOR U20356 ( .A(n19321), .B(n19332), .Z(n19323) );
  XOR U20357 ( .A(n19333), .B(n19334), .Z(n19321) );
  AND U20358 ( .A(n19335), .B(n19336), .Z(n19334) );
  XNOR U20359 ( .A(n19337), .B(n19333), .Z(n19336) );
  XOR U20360 ( .A(n19338), .B(e_input[439]), .Z(n19329) );
  IV U20361 ( .A(n19327), .Z(n19338) );
  XOR U20362 ( .A(n19339), .B(n19340), .Z(n19327) );
  AND U20363 ( .A(n19341), .B(n19342), .Z(n19340) );
  XNOR U20364 ( .A(n19339), .B(n9672), .Z(n19342) );
  XNOR U20365 ( .A(n19335), .B(n19337), .Z(n9672) );
  NAND U20366 ( .A(n19343), .B(e_input[438]), .Z(n19337) );
  NAND U20367 ( .A(n12323), .B(e_input[438]), .Z(n19343) );
  XNOR U20368 ( .A(n19333), .B(n19344), .Z(n19335) );
  XOR U20369 ( .A(n19345), .B(n19346), .Z(n19333) );
  AND U20370 ( .A(n19347), .B(n19348), .Z(n19346) );
  XNOR U20371 ( .A(n19349), .B(n19345), .Z(n19348) );
  XOR U20372 ( .A(n19350), .B(e_input[438]), .Z(n19341) );
  IV U20373 ( .A(n19339), .Z(n19350) );
  XOR U20374 ( .A(n19351), .B(n19352), .Z(n19339) );
  AND U20375 ( .A(n19353), .B(n19354), .Z(n19352) );
  XNOR U20376 ( .A(n19351), .B(n9678), .Z(n19354) );
  XNOR U20377 ( .A(n19347), .B(n19349), .Z(n9678) );
  NAND U20378 ( .A(n19355), .B(e_input[437]), .Z(n19349) );
  NAND U20379 ( .A(n12323), .B(e_input[437]), .Z(n19355) );
  XNOR U20380 ( .A(n19345), .B(n19356), .Z(n19347) );
  XOR U20381 ( .A(n19357), .B(n19358), .Z(n19345) );
  AND U20382 ( .A(n19359), .B(n19360), .Z(n19358) );
  XNOR U20383 ( .A(n19361), .B(n19357), .Z(n19360) );
  XOR U20384 ( .A(n19362), .B(e_input[437]), .Z(n19353) );
  IV U20385 ( .A(n19351), .Z(n19362) );
  XOR U20386 ( .A(n19363), .B(n19364), .Z(n19351) );
  AND U20387 ( .A(n19365), .B(n19366), .Z(n19364) );
  XNOR U20388 ( .A(n19363), .B(n9684), .Z(n19366) );
  XNOR U20389 ( .A(n19359), .B(n19361), .Z(n9684) );
  NAND U20390 ( .A(n19367), .B(e_input[436]), .Z(n19361) );
  NAND U20391 ( .A(n12323), .B(e_input[436]), .Z(n19367) );
  XNOR U20392 ( .A(n19357), .B(n19368), .Z(n19359) );
  XOR U20393 ( .A(n19369), .B(n19370), .Z(n19357) );
  AND U20394 ( .A(n19371), .B(n19372), .Z(n19370) );
  XNOR U20395 ( .A(n19373), .B(n19369), .Z(n19372) );
  XOR U20396 ( .A(n19374), .B(e_input[436]), .Z(n19365) );
  IV U20397 ( .A(n19363), .Z(n19374) );
  XOR U20398 ( .A(n19375), .B(n19376), .Z(n19363) );
  AND U20399 ( .A(n19377), .B(n19378), .Z(n19376) );
  XNOR U20400 ( .A(n19375), .B(n9690), .Z(n19378) );
  XNOR U20401 ( .A(n19371), .B(n19373), .Z(n9690) );
  NAND U20402 ( .A(n19379), .B(e_input[435]), .Z(n19373) );
  NAND U20403 ( .A(n12323), .B(e_input[435]), .Z(n19379) );
  XNOR U20404 ( .A(n19369), .B(n19380), .Z(n19371) );
  XOR U20405 ( .A(n19381), .B(n19382), .Z(n19369) );
  AND U20406 ( .A(n19383), .B(n19384), .Z(n19382) );
  XNOR U20407 ( .A(n19385), .B(n19381), .Z(n19384) );
  XOR U20408 ( .A(n19386), .B(e_input[435]), .Z(n19377) );
  IV U20409 ( .A(n19375), .Z(n19386) );
  XOR U20410 ( .A(n19387), .B(n19388), .Z(n19375) );
  AND U20411 ( .A(n19389), .B(n19390), .Z(n19388) );
  XNOR U20412 ( .A(n19387), .B(n9696), .Z(n19390) );
  XNOR U20413 ( .A(n19383), .B(n19385), .Z(n9696) );
  NAND U20414 ( .A(n19391), .B(e_input[434]), .Z(n19385) );
  NAND U20415 ( .A(n12323), .B(e_input[434]), .Z(n19391) );
  XNOR U20416 ( .A(n19381), .B(n19392), .Z(n19383) );
  XOR U20417 ( .A(n19393), .B(n19394), .Z(n19381) );
  AND U20418 ( .A(n19395), .B(n19396), .Z(n19394) );
  XNOR U20419 ( .A(n19397), .B(n19393), .Z(n19396) );
  XOR U20420 ( .A(n19398), .B(e_input[434]), .Z(n19389) );
  IV U20421 ( .A(n19387), .Z(n19398) );
  XOR U20422 ( .A(n19399), .B(n19400), .Z(n19387) );
  AND U20423 ( .A(n19401), .B(n19402), .Z(n19400) );
  XNOR U20424 ( .A(n19399), .B(n9702), .Z(n19402) );
  XNOR U20425 ( .A(n19395), .B(n19397), .Z(n9702) );
  NAND U20426 ( .A(n19403), .B(e_input[433]), .Z(n19397) );
  NAND U20427 ( .A(n12323), .B(e_input[433]), .Z(n19403) );
  XNOR U20428 ( .A(n19393), .B(n19404), .Z(n19395) );
  XOR U20429 ( .A(n19405), .B(n19406), .Z(n19393) );
  AND U20430 ( .A(n19407), .B(n19408), .Z(n19406) );
  XNOR U20431 ( .A(n19409), .B(n19405), .Z(n19408) );
  XOR U20432 ( .A(n19410), .B(e_input[433]), .Z(n19401) );
  IV U20433 ( .A(n19399), .Z(n19410) );
  XOR U20434 ( .A(n19411), .B(n19412), .Z(n19399) );
  AND U20435 ( .A(n19413), .B(n19414), .Z(n19412) );
  XNOR U20436 ( .A(n19411), .B(n9708), .Z(n19414) );
  XNOR U20437 ( .A(n19407), .B(n19409), .Z(n9708) );
  NAND U20438 ( .A(n19415), .B(e_input[432]), .Z(n19409) );
  NAND U20439 ( .A(n12323), .B(e_input[432]), .Z(n19415) );
  XNOR U20440 ( .A(n19405), .B(n19416), .Z(n19407) );
  XOR U20441 ( .A(n19417), .B(n19418), .Z(n19405) );
  AND U20442 ( .A(n19419), .B(n19420), .Z(n19418) );
  XNOR U20443 ( .A(n19421), .B(n19417), .Z(n19420) );
  XOR U20444 ( .A(n19422), .B(e_input[432]), .Z(n19413) );
  IV U20445 ( .A(n19411), .Z(n19422) );
  XOR U20446 ( .A(n19423), .B(n19424), .Z(n19411) );
  AND U20447 ( .A(n19425), .B(n19426), .Z(n19424) );
  XNOR U20448 ( .A(n19423), .B(n9714), .Z(n19426) );
  XNOR U20449 ( .A(n19419), .B(n19421), .Z(n9714) );
  NAND U20450 ( .A(n19427), .B(e_input[431]), .Z(n19421) );
  NAND U20451 ( .A(n12323), .B(e_input[431]), .Z(n19427) );
  XNOR U20452 ( .A(n19417), .B(n19428), .Z(n19419) );
  XOR U20453 ( .A(n19429), .B(n19430), .Z(n19417) );
  AND U20454 ( .A(n19431), .B(n19432), .Z(n19430) );
  XNOR U20455 ( .A(n19433), .B(n19429), .Z(n19432) );
  XOR U20456 ( .A(n19434), .B(e_input[431]), .Z(n19425) );
  IV U20457 ( .A(n19423), .Z(n19434) );
  XOR U20458 ( .A(n19435), .B(n19436), .Z(n19423) );
  AND U20459 ( .A(n19437), .B(n19438), .Z(n19436) );
  XNOR U20460 ( .A(n19435), .B(n9720), .Z(n19438) );
  XNOR U20461 ( .A(n19431), .B(n19433), .Z(n9720) );
  NAND U20462 ( .A(n19439), .B(e_input[430]), .Z(n19433) );
  NAND U20463 ( .A(n12323), .B(e_input[430]), .Z(n19439) );
  XNOR U20464 ( .A(n19429), .B(n19440), .Z(n19431) );
  XOR U20465 ( .A(n19441), .B(n19442), .Z(n19429) );
  AND U20466 ( .A(n19443), .B(n19444), .Z(n19442) );
  XNOR U20467 ( .A(n19445), .B(n19441), .Z(n19444) );
  XOR U20468 ( .A(n19446), .B(e_input[430]), .Z(n19437) );
  IV U20469 ( .A(n19435), .Z(n19446) );
  XOR U20470 ( .A(n19447), .B(n19448), .Z(n19435) );
  AND U20471 ( .A(n19449), .B(n19450), .Z(n19448) );
  XNOR U20472 ( .A(n19447), .B(n9726), .Z(n19450) );
  XNOR U20473 ( .A(n19443), .B(n19445), .Z(n9726) );
  NAND U20474 ( .A(n19451), .B(e_input[429]), .Z(n19445) );
  NAND U20475 ( .A(n12323), .B(e_input[429]), .Z(n19451) );
  XNOR U20476 ( .A(n19441), .B(n19452), .Z(n19443) );
  XOR U20477 ( .A(n19453), .B(n19454), .Z(n19441) );
  AND U20478 ( .A(n19455), .B(n19456), .Z(n19454) );
  XNOR U20479 ( .A(n19457), .B(n19453), .Z(n19456) );
  XOR U20480 ( .A(n19458), .B(e_input[429]), .Z(n19449) );
  IV U20481 ( .A(n19447), .Z(n19458) );
  XOR U20482 ( .A(n19459), .B(n19460), .Z(n19447) );
  AND U20483 ( .A(n19461), .B(n19462), .Z(n19460) );
  XNOR U20484 ( .A(n19459), .B(n9732), .Z(n19462) );
  XNOR U20485 ( .A(n19455), .B(n19457), .Z(n9732) );
  NAND U20486 ( .A(n19463), .B(e_input[428]), .Z(n19457) );
  NAND U20487 ( .A(n12323), .B(e_input[428]), .Z(n19463) );
  XNOR U20488 ( .A(n19453), .B(n19464), .Z(n19455) );
  XOR U20489 ( .A(n19465), .B(n19466), .Z(n19453) );
  AND U20490 ( .A(n19467), .B(n19468), .Z(n19466) );
  XNOR U20491 ( .A(n19469), .B(n19465), .Z(n19468) );
  XOR U20492 ( .A(n19470), .B(e_input[428]), .Z(n19461) );
  IV U20493 ( .A(n19459), .Z(n19470) );
  XOR U20494 ( .A(n19471), .B(n19472), .Z(n19459) );
  AND U20495 ( .A(n19473), .B(n19474), .Z(n19472) );
  XNOR U20496 ( .A(n19471), .B(n9738), .Z(n19474) );
  XNOR U20497 ( .A(n19467), .B(n19469), .Z(n9738) );
  NAND U20498 ( .A(n19475), .B(e_input[427]), .Z(n19469) );
  NAND U20499 ( .A(n12323), .B(e_input[427]), .Z(n19475) );
  XNOR U20500 ( .A(n19465), .B(n19476), .Z(n19467) );
  XOR U20501 ( .A(n19477), .B(n19478), .Z(n19465) );
  AND U20502 ( .A(n19479), .B(n19480), .Z(n19478) );
  XNOR U20503 ( .A(n19481), .B(n19477), .Z(n19480) );
  XOR U20504 ( .A(n19482), .B(e_input[427]), .Z(n19473) );
  IV U20505 ( .A(n19471), .Z(n19482) );
  XOR U20506 ( .A(n19483), .B(n19484), .Z(n19471) );
  AND U20507 ( .A(n19485), .B(n19486), .Z(n19484) );
  XNOR U20508 ( .A(n19483), .B(n9744), .Z(n19486) );
  XNOR U20509 ( .A(n19479), .B(n19481), .Z(n9744) );
  NAND U20510 ( .A(n19487), .B(e_input[426]), .Z(n19481) );
  NAND U20511 ( .A(n12323), .B(e_input[426]), .Z(n19487) );
  XNOR U20512 ( .A(n19477), .B(n19488), .Z(n19479) );
  XOR U20513 ( .A(n19489), .B(n19490), .Z(n19477) );
  AND U20514 ( .A(n19491), .B(n19492), .Z(n19490) );
  XNOR U20515 ( .A(n19493), .B(n19489), .Z(n19492) );
  XOR U20516 ( .A(n19494), .B(e_input[426]), .Z(n19485) );
  IV U20517 ( .A(n19483), .Z(n19494) );
  XOR U20518 ( .A(n19495), .B(n19496), .Z(n19483) );
  AND U20519 ( .A(n19497), .B(n19498), .Z(n19496) );
  XNOR U20520 ( .A(n19495), .B(n9750), .Z(n19498) );
  XNOR U20521 ( .A(n19491), .B(n19493), .Z(n9750) );
  NAND U20522 ( .A(n19499), .B(e_input[425]), .Z(n19493) );
  NAND U20523 ( .A(n12323), .B(e_input[425]), .Z(n19499) );
  XNOR U20524 ( .A(n19489), .B(n19500), .Z(n19491) );
  XOR U20525 ( .A(n19501), .B(n19502), .Z(n19489) );
  AND U20526 ( .A(n19503), .B(n19504), .Z(n19502) );
  XNOR U20527 ( .A(n19505), .B(n19501), .Z(n19504) );
  XOR U20528 ( .A(n19506), .B(e_input[425]), .Z(n19497) );
  IV U20529 ( .A(n19495), .Z(n19506) );
  XOR U20530 ( .A(n19507), .B(n19508), .Z(n19495) );
  AND U20531 ( .A(n19509), .B(n19510), .Z(n19508) );
  XNOR U20532 ( .A(n19507), .B(n9756), .Z(n19510) );
  XNOR U20533 ( .A(n19503), .B(n19505), .Z(n9756) );
  NAND U20534 ( .A(n19511), .B(e_input[424]), .Z(n19505) );
  NAND U20535 ( .A(n12323), .B(e_input[424]), .Z(n19511) );
  XNOR U20536 ( .A(n19501), .B(n19512), .Z(n19503) );
  XOR U20537 ( .A(n19513), .B(n19514), .Z(n19501) );
  AND U20538 ( .A(n19515), .B(n19516), .Z(n19514) );
  XNOR U20539 ( .A(n19517), .B(n19513), .Z(n19516) );
  XOR U20540 ( .A(n19518), .B(e_input[424]), .Z(n19509) );
  IV U20541 ( .A(n19507), .Z(n19518) );
  XOR U20542 ( .A(n19519), .B(n19520), .Z(n19507) );
  AND U20543 ( .A(n19521), .B(n19522), .Z(n19520) );
  XNOR U20544 ( .A(n19519), .B(n9762), .Z(n19522) );
  XNOR U20545 ( .A(n19515), .B(n19517), .Z(n9762) );
  NAND U20546 ( .A(n19523), .B(e_input[423]), .Z(n19517) );
  NAND U20547 ( .A(n12323), .B(e_input[423]), .Z(n19523) );
  XNOR U20548 ( .A(n19513), .B(n19524), .Z(n19515) );
  XOR U20549 ( .A(n19525), .B(n19526), .Z(n19513) );
  AND U20550 ( .A(n19527), .B(n19528), .Z(n19526) );
  XNOR U20551 ( .A(n19529), .B(n19525), .Z(n19528) );
  XOR U20552 ( .A(n19530), .B(e_input[423]), .Z(n19521) );
  IV U20553 ( .A(n19519), .Z(n19530) );
  XOR U20554 ( .A(n19531), .B(n19532), .Z(n19519) );
  AND U20555 ( .A(n19533), .B(n19534), .Z(n19532) );
  XNOR U20556 ( .A(n19531), .B(n9768), .Z(n19534) );
  XNOR U20557 ( .A(n19527), .B(n19529), .Z(n9768) );
  NAND U20558 ( .A(n19535), .B(e_input[422]), .Z(n19529) );
  NAND U20559 ( .A(n12323), .B(e_input[422]), .Z(n19535) );
  XNOR U20560 ( .A(n19525), .B(n19536), .Z(n19527) );
  XOR U20561 ( .A(n19537), .B(n19538), .Z(n19525) );
  AND U20562 ( .A(n19539), .B(n19540), .Z(n19538) );
  XNOR U20563 ( .A(n19541), .B(n19537), .Z(n19540) );
  XOR U20564 ( .A(n19542), .B(e_input[422]), .Z(n19533) );
  IV U20565 ( .A(n19531), .Z(n19542) );
  XOR U20566 ( .A(n19543), .B(n19544), .Z(n19531) );
  AND U20567 ( .A(n19545), .B(n19546), .Z(n19544) );
  XNOR U20568 ( .A(n19543), .B(n9774), .Z(n19546) );
  XNOR U20569 ( .A(n19539), .B(n19541), .Z(n9774) );
  NAND U20570 ( .A(n19547), .B(e_input[421]), .Z(n19541) );
  NAND U20571 ( .A(n12323), .B(e_input[421]), .Z(n19547) );
  XNOR U20572 ( .A(n19537), .B(n19548), .Z(n19539) );
  XOR U20573 ( .A(n19549), .B(n19550), .Z(n19537) );
  AND U20574 ( .A(n19551), .B(n19552), .Z(n19550) );
  XNOR U20575 ( .A(n19553), .B(n19549), .Z(n19552) );
  XOR U20576 ( .A(n19554), .B(e_input[421]), .Z(n19545) );
  IV U20577 ( .A(n19543), .Z(n19554) );
  XOR U20578 ( .A(n19555), .B(n19556), .Z(n19543) );
  AND U20579 ( .A(n19557), .B(n19558), .Z(n19556) );
  XNOR U20580 ( .A(n19555), .B(n9780), .Z(n19558) );
  XNOR U20581 ( .A(n19551), .B(n19553), .Z(n9780) );
  NAND U20582 ( .A(n19559), .B(e_input[420]), .Z(n19553) );
  NAND U20583 ( .A(n12323), .B(e_input[420]), .Z(n19559) );
  XNOR U20584 ( .A(n19549), .B(n19560), .Z(n19551) );
  XOR U20585 ( .A(n19561), .B(n19562), .Z(n19549) );
  AND U20586 ( .A(n19563), .B(n19564), .Z(n19562) );
  XNOR U20587 ( .A(n19565), .B(n19561), .Z(n19564) );
  XOR U20588 ( .A(n19566), .B(e_input[420]), .Z(n19557) );
  IV U20589 ( .A(n19555), .Z(n19566) );
  XOR U20590 ( .A(n19567), .B(n19568), .Z(n19555) );
  AND U20591 ( .A(n19569), .B(n19570), .Z(n19568) );
  XNOR U20592 ( .A(n19567), .B(n9786), .Z(n19570) );
  XNOR U20593 ( .A(n19563), .B(n19565), .Z(n9786) );
  NAND U20594 ( .A(n19571), .B(e_input[419]), .Z(n19565) );
  NAND U20595 ( .A(n12323), .B(e_input[419]), .Z(n19571) );
  XNOR U20596 ( .A(n19561), .B(n19572), .Z(n19563) );
  XOR U20597 ( .A(n19573), .B(n19574), .Z(n19561) );
  AND U20598 ( .A(n19575), .B(n19576), .Z(n19574) );
  XNOR U20599 ( .A(n19577), .B(n19573), .Z(n19576) );
  XOR U20600 ( .A(n19578), .B(e_input[419]), .Z(n19569) );
  IV U20601 ( .A(n19567), .Z(n19578) );
  XOR U20602 ( .A(n19579), .B(n19580), .Z(n19567) );
  AND U20603 ( .A(n19581), .B(n19582), .Z(n19580) );
  XNOR U20604 ( .A(n19579), .B(n9792), .Z(n19582) );
  XNOR U20605 ( .A(n19575), .B(n19577), .Z(n9792) );
  NAND U20606 ( .A(n19583), .B(e_input[418]), .Z(n19577) );
  NAND U20607 ( .A(n12323), .B(e_input[418]), .Z(n19583) );
  XNOR U20608 ( .A(n19573), .B(n19584), .Z(n19575) );
  XOR U20609 ( .A(n19585), .B(n19586), .Z(n19573) );
  AND U20610 ( .A(n19587), .B(n19588), .Z(n19586) );
  XNOR U20611 ( .A(n19589), .B(n19585), .Z(n19588) );
  XOR U20612 ( .A(n19590), .B(e_input[418]), .Z(n19581) );
  IV U20613 ( .A(n19579), .Z(n19590) );
  XOR U20614 ( .A(n19591), .B(n19592), .Z(n19579) );
  AND U20615 ( .A(n19593), .B(n19594), .Z(n19592) );
  XNOR U20616 ( .A(n19591), .B(n9798), .Z(n19594) );
  XNOR U20617 ( .A(n19587), .B(n19589), .Z(n9798) );
  NAND U20618 ( .A(n19595), .B(e_input[417]), .Z(n19589) );
  NAND U20619 ( .A(n12323), .B(e_input[417]), .Z(n19595) );
  XNOR U20620 ( .A(n19585), .B(n19596), .Z(n19587) );
  XOR U20621 ( .A(n19597), .B(n19598), .Z(n19585) );
  AND U20622 ( .A(n19599), .B(n19600), .Z(n19598) );
  XNOR U20623 ( .A(n19601), .B(n19597), .Z(n19600) );
  XOR U20624 ( .A(n19602), .B(e_input[417]), .Z(n19593) );
  IV U20625 ( .A(n19591), .Z(n19602) );
  XOR U20626 ( .A(n19603), .B(n19604), .Z(n19591) );
  AND U20627 ( .A(n19605), .B(n19606), .Z(n19604) );
  XNOR U20628 ( .A(n19603), .B(n9804), .Z(n19606) );
  XNOR U20629 ( .A(n19599), .B(n19601), .Z(n9804) );
  NAND U20630 ( .A(n19607), .B(e_input[416]), .Z(n19601) );
  NAND U20631 ( .A(n12323), .B(e_input[416]), .Z(n19607) );
  XNOR U20632 ( .A(n19597), .B(n19608), .Z(n19599) );
  XOR U20633 ( .A(n19609), .B(n19610), .Z(n19597) );
  AND U20634 ( .A(n19611), .B(n19612), .Z(n19610) );
  XNOR U20635 ( .A(n19613), .B(n19609), .Z(n19612) );
  XOR U20636 ( .A(n19614), .B(e_input[416]), .Z(n19605) );
  IV U20637 ( .A(n19603), .Z(n19614) );
  XOR U20638 ( .A(n19615), .B(n19616), .Z(n19603) );
  AND U20639 ( .A(n19617), .B(n19618), .Z(n19616) );
  XNOR U20640 ( .A(n19615), .B(n9810), .Z(n19618) );
  XNOR U20641 ( .A(n19611), .B(n19613), .Z(n9810) );
  NAND U20642 ( .A(n19619), .B(e_input[415]), .Z(n19613) );
  NAND U20643 ( .A(n12323), .B(e_input[415]), .Z(n19619) );
  XNOR U20644 ( .A(n19609), .B(n19620), .Z(n19611) );
  XOR U20645 ( .A(n19621), .B(n19622), .Z(n19609) );
  AND U20646 ( .A(n19623), .B(n19624), .Z(n19622) );
  XNOR U20647 ( .A(n19625), .B(n19621), .Z(n19624) );
  XOR U20648 ( .A(n19626), .B(e_input[415]), .Z(n19617) );
  IV U20649 ( .A(n19615), .Z(n19626) );
  XOR U20650 ( .A(n19627), .B(n19628), .Z(n19615) );
  AND U20651 ( .A(n19629), .B(n19630), .Z(n19628) );
  XNOR U20652 ( .A(n19627), .B(n9816), .Z(n19630) );
  XNOR U20653 ( .A(n19623), .B(n19625), .Z(n9816) );
  NAND U20654 ( .A(n19631), .B(e_input[414]), .Z(n19625) );
  NAND U20655 ( .A(n12323), .B(e_input[414]), .Z(n19631) );
  XNOR U20656 ( .A(n19621), .B(n19632), .Z(n19623) );
  XOR U20657 ( .A(n19633), .B(n19634), .Z(n19621) );
  AND U20658 ( .A(n19635), .B(n19636), .Z(n19634) );
  XNOR U20659 ( .A(n19637), .B(n19633), .Z(n19636) );
  XOR U20660 ( .A(n19638), .B(e_input[414]), .Z(n19629) );
  IV U20661 ( .A(n19627), .Z(n19638) );
  XOR U20662 ( .A(n19639), .B(n19640), .Z(n19627) );
  AND U20663 ( .A(n19641), .B(n19642), .Z(n19640) );
  XNOR U20664 ( .A(n19639), .B(n9822), .Z(n19642) );
  XNOR U20665 ( .A(n19635), .B(n19637), .Z(n9822) );
  NAND U20666 ( .A(n19643), .B(e_input[413]), .Z(n19637) );
  NAND U20667 ( .A(n12323), .B(e_input[413]), .Z(n19643) );
  XNOR U20668 ( .A(n19633), .B(n19644), .Z(n19635) );
  XOR U20669 ( .A(n19645), .B(n19646), .Z(n19633) );
  AND U20670 ( .A(n19647), .B(n19648), .Z(n19646) );
  XNOR U20671 ( .A(n19649), .B(n19645), .Z(n19648) );
  XOR U20672 ( .A(n19650), .B(e_input[413]), .Z(n19641) );
  IV U20673 ( .A(n19639), .Z(n19650) );
  XOR U20674 ( .A(n19651), .B(n19652), .Z(n19639) );
  AND U20675 ( .A(n19653), .B(n19654), .Z(n19652) );
  XNOR U20676 ( .A(n19651), .B(n9828), .Z(n19654) );
  XNOR U20677 ( .A(n19647), .B(n19649), .Z(n9828) );
  NAND U20678 ( .A(n19655), .B(e_input[412]), .Z(n19649) );
  NAND U20679 ( .A(n12323), .B(e_input[412]), .Z(n19655) );
  XNOR U20680 ( .A(n19645), .B(n19656), .Z(n19647) );
  XOR U20681 ( .A(n19657), .B(n19658), .Z(n19645) );
  AND U20682 ( .A(n19659), .B(n19660), .Z(n19658) );
  XNOR U20683 ( .A(n19661), .B(n19657), .Z(n19660) );
  XOR U20684 ( .A(n19662), .B(e_input[412]), .Z(n19653) );
  IV U20685 ( .A(n19651), .Z(n19662) );
  XOR U20686 ( .A(n19663), .B(n19664), .Z(n19651) );
  AND U20687 ( .A(n19665), .B(n19666), .Z(n19664) );
  XNOR U20688 ( .A(n19663), .B(n9834), .Z(n19666) );
  XNOR U20689 ( .A(n19659), .B(n19661), .Z(n9834) );
  NAND U20690 ( .A(n19667), .B(e_input[411]), .Z(n19661) );
  NAND U20691 ( .A(n12323), .B(e_input[411]), .Z(n19667) );
  XNOR U20692 ( .A(n19657), .B(n19668), .Z(n19659) );
  XOR U20693 ( .A(n19669), .B(n19670), .Z(n19657) );
  AND U20694 ( .A(n19671), .B(n19672), .Z(n19670) );
  XNOR U20695 ( .A(n19673), .B(n19669), .Z(n19672) );
  XOR U20696 ( .A(n19674), .B(e_input[411]), .Z(n19665) );
  IV U20697 ( .A(n19663), .Z(n19674) );
  XOR U20698 ( .A(n19675), .B(n19676), .Z(n19663) );
  AND U20699 ( .A(n19677), .B(n19678), .Z(n19676) );
  XNOR U20700 ( .A(n19675), .B(n9840), .Z(n19678) );
  XNOR U20701 ( .A(n19671), .B(n19673), .Z(n9840) );
  NAND U20702 ( .A(n19679), .B(e_input[410]), .Z(n19673) );
  NAND U20703 ( .A(n12323), .B(e_input[410]), .Z(n19679) );
  XNOR U20704 ( .A(n19669), .B(n19680), .Z(n19671) );
  XOR U20705 ( .A(n19681), .B(n19682), .Z(n19669) );
  AND U20706 ( .A(n19683), .B(n19684), .Z(n19682) );
  XNOR U20707 ( .A(n19685), .B(n19681), .Z(n19684) );
  XOR U20708 ( .A(n19686), .B(e_input[410]), .Z(n19677) );
  IV U20709 ( .A(n19675), .Z(n19686) );
  XOR U20710 ( .A(n19687), .B(n19688), .Z(n19675) );
  AND U20711 ( .A(n19689), .B(n19690), .Z(n19688) );
  XNOR U20712 ( .A(n19687), .B(n9846), .Z(n19690) );
  XNOR U20713 ( .A(n19683), .B(n19685), .Z(n9846) );
  NAND U20714 ( .A(n19691), .B(e_input[409]), .Z(n19685) );
  NAND U20715 ( .A(n12323), .B(e_input[409]), .Z(n19691) );
  XNOR U20716 ( .A(n19681), .B(n19692), .Z(n19683) );
  XOR U20717 ( .A(n19693), .B(n19694), .Z(n19681) );
  AND U20718 ( .A(n19695), .B(n19696), .Z(n19694) );
  XNOR U20719 ( .A(n19697), .B(n19693), .Z(n19696) );
  XOR U20720 ( .A(n19698), .B(e_input[409]), .Z(n19689) );
  IV U20721 ( .A(n19687), .Z(n19698) );
  XOR U20722 ( .A(n19699), .B(n19700), .Z(n19687) );
  AND U20723 ( .A(n19701), .B(n19702), .Z(n19700) );
  XNOR U20724 ( .A(n19699), .B(n9852), .Z(n19702) );
  XNOR U20725 ( .A(n19695), .B(n19697), .Z(n9852) );
  NAND U20726 ( .A(n19703), .B(e_input[408]), .Z(n19697) );
  NAND U20727 ( .A(n12323), .B(e_input[408]), .Z(n19703) );
  XNOR U20728 ( .A(n19693), .B(n19704), .Z(n19695) );
  XOR U20729 ( .A(n19705), .B(n19706), .Z(n19693) );
  AND U20730 ( .A(n19707), .B(n19708), .Z(n19706) );
  XNOR U20731 ( .A(n19709), .B(n19705), .Z(n19708) );
  XOR U20732 ( .A(n19710), .B(e_input[408]), .Z(n19701) );
  IV U20733 ( .A(n19699), .Z(n19710) );
  XOR U20734 ( .A(n19711), .B(n19712), .Z(n19699) );
  AND U20735 ( .A(n19713), .B(n19714), .Z(n19712) );
  XNOR U20736 ( .A(n19711), .B(n9858), .Z(n19714) );
  XNOR U20737 ( .A(n19707), .B(n19709), .Z(n9858) );
  NAND U20738 ( .A(n19715), .B(e_input[407]), .Z(n19709) );
  NAND U20739 ( .A(n12323), .B(e_input[407]), .Z(n19715) );
  XNOR U20740 ( .A(n19705), .B(n19716), .Z(n19707) );
  XOR U20741 ( .A(n19717), .B(n19718), .Z(n19705) );
  AND U20742 ( .A(n19719), .B(n19720), .Z(n19718) );
  XNOR U20743 ( .A(n19721), .B(n19717), .Z(n19720) );
  XOR U20744 ( .A(n19722), .B(e_input[407]), .Z(n19713) );
  IV U20745 ( .A(n19711), .Z(n19722) );
  XOR U20746 ( .A(n19723), .B(n19724), .Z(n19711) );
  AND U20747 ( .A(n19725), .B(n19726), .Z(n19724) );
  XNOR U20748 ( .A(n19723), .B(n9864), .Z(n19726) );
  XNOR U20749 ( .A(n19719), .B(n19721), .Z(n9864) );
  NAND U20750 ( .A(n19727), .B(e_input[406]), .Z(n19721) );
  NAND U20751 ( .A(n12323), .B(e_input[406]), .Z(n19727) );
  XNOR U20752 ( .A(n19717), .B(n19728), .Z(n19719) );
  XOR U20753 ( .A(n19729), .B(n19730), .Z(n19717) );
  AND U20754 ( .A(n19731), .B(n19732), .Z(n19730) );
  XNOR U20755 ( .A(n19733), .B(n19729), .Z(n19732) );
  XOR U20756 ( .A(n19734), .B(e_input[406]), .Z(n19725) );
  IV U20757 ( .A(n19723), .Z(n19734) );
  XOR U20758 ( .A(n19735), .B(n19736), .Z(n19723) );
  AND U20759 ( .A(n19737), .B(n19738), .Z(n19736) );
  XNOR U20760 ( .A(n19735), .B(n9870), .Z(n19738) );
  XNOR U20761 ( .A(n19731), .B(n19733), .Z(n9870) );
  NAND U20762 ( .A(n19739), .B(e_input[405]), .Z(n19733) );
  NAND U20763 ( .A(n12323), .B(e_input[405]), .Z(n19739) );
  XNOR U20764 ( .A(n19729), .B(n19740), .Z(n19731) );
  XOR U20765 ( .A(n19741), .B(n19742), .Z(n19729) );
  AND U20766 ( .A(n19743), .B(n19744), .Z(n19742) );
  XNOR U20767 ( .A(n19745), .B(n19741), .Z(n19744) );
  XOR U20768 ( .A(n19746), .B(e_input[405]), .Z(n19737) );
  IV U20769 ( .A(n19735), .Z(n19746) );
  XOR U20770 ( .A(n19747), .B(n19748), .Z(n19735) );
  AND U20771 ( .A(n19749), .B(n19750), .Z(n19748) );
  XNOR U20772 ( .A(n19747), .B(n9876), .Z(n19750) );
  XNOR U20773 ( .A(n19743), .B(n19745), .Z(n9876) );
  NAND U20774 ( .A(n19751), .B(e_input[404]), .Z(n19745) );
  NAND U20775 ( .A(n12323), .B(e_input[404]), .Z(n19751) );
  XNOR U20776 ( .A(n19741), .B(n19752), .Z(n19743) );
  XOR U20777 ( .A(n19753), .B(n19754), .Z(n19741) );
  AND U20778 ( .A(n19755), .B(n19756), .Z(n19754) );
  XNOR U20779 ( .A(n19757), .B(n19753), .Z(n19756) );
  XOR U20780 ( .A(n19758), .B(e_input[404]), .Z(n19749) );
  IV U20781 ( .A(n19747), .Z(n19758) );
  XOR U20782 ( .A(n19759), .B(n19760), .Z(n19747) );
  AND U20783 ( .A(n19761), .B(n19762), .Z(n19760) );
  XNOR U20784 ( .A(n19759), .B(n9882), .Z(n19762) );
  XNOR U20785 ( .A(n19755), .B(n19757), .Z(n9882) );
  NAND U20786 ( .A(n19763), .B(e_input[403]), .Z(n19757) );
  NAND U20787 ( .A(n12323), .B(e_input[403]), .Z(n19763) );
  XNOR U20788 ( .A(n19753), .B(n19764), .Z(n19755) );
  XOR U20789 ( .A(n19765), .B(n19766), .Z(n19753) );
  AND U20790 ( .A(n19767), .B(n19768), .Z(n19766) );
  XNOR U20791 ( .A(n19769), .B(n19765), .Z(n19768) );
  XOR U20792 ( .A(n19770), .B(e_input[403]), .Z(n19761) );
  IV U20793 ( .A(n19759), .Z(n19770) );
  XOR U20794 ( .A(n19771), .B(n19772), .Z(n19759) );
  AND U20795 ( .A(n19773), .B(n19774), .Z(n19772) );
  XNOR U20796 ( .A(n19771), .B(n9888), .Z(n19774) );
  XNOR U20797 ( .A(n19767), .B(n19769), .Z(n9888) );
  NAND U20798 ( .A(n19775), .B(e_input[402]), .Z(n19769) );
  NAND U20799 ( .A(n12323), .B(e_input[402]), .Z(n19775) );
  XNOR U20800 ( .A(n19765), .B(n19776), .Z(n19767) );
  XOR U20801 ( .A(n19777), .B(n19778), .Z(n19765) );
  AND U20802 ( .A(n19779), .B(n19780), .Z(n19778) );
  XNOR U20803 ( .A(n19781), .B(n19777), .Z(n19780) );
  XOR U20804 ( .A(n19782), .B(e_input[402]), .Z(n19773) );
  IV U20805 ( .A(n19771), .Z(n19782) );
  XOR U20806 ( .A(n19783), .B(n19784), .Z(n19771) );
  AND U20807 ( .A(n19785), .B(n19786), .Z(n19784) );
  XNOR U20808 ( .A(n19783), .B(n9894), .Z(n19786) );
  XNOR U20809 ( .A(n19779), .B(n19781), .Z(n9894) );
  NAND U20810 ( .A(n19787), .B(e_input[401]), .Z(n19781) );
  NAND U20811 ( .A(n12323), .B(e_input[401]), .Z(n19787) );
  XNOR U20812 ( .A(n19777), .B(n19788), .Z(n19779) );
  XOR U20813 ( .A(n19789), .B(n19790), .Z(n19777) );
  AND U20814 ( .A(n19791), .B(n19792), .Z(n19790) );
  XNOR U20815 ( .A(n19793), .B(n19789), .Z(n19792) );
  XOR U20816 ( .A(n19794), .B(e_input[401]), .Z(n19785) );
  IV U20817 ( .A(n19783), .Z(n19794) );
  XOR U20818 ( .A(n19795), .B(n19796), .Z(n19783) );
  AND U20819 ( .A(n19797), .B(n19798), .Z(n19796) );
  XNOR U20820 ( .A(n19795), .B(n9900), .Z(n19798) );
  XNOR U20821 ( .A(n19791), .B(n19793), .Z(n9900) );
  NAND U20822 ( .A(n19799), .B(e_input[400]), .Z(n19793) );
  NAND U20823 ( .A(n12323), .B(e_input[400]), .Z(n19799) );
  XNOR U20824 ( .A(n19789), .B(n19800), .Z(n19791) );
  XOR U20825 ( .A(n19801), .B(n19802), .Z(n19789) );
  AND U20826 ( .A(n19803), .B(n19804), .Z(n19802) );
  XNOR U20827 ( .A(n19805), .B(n19801), .Z(n19804) );
  XOR U20828 ( .A(n19806), .B(e_input[400]), .Z(n19797) );
  IV U20829 ( .A(n19795), .Z(n19806) );
  XOR U20830 ( .A(n19807), .B(n19808), .Z(n19795) );
  AND U20831 ( .A(n19809), .B(n19810), .Z(n19808) );
  XNOR U20832 ( .A(n19807), .B(n9906), .Z(n19810) );
  XNOR U20833 ( .A(n19803), .B(n19805), .Z(n9906) );
  NAND U20834 ( .A(n19811), .B(e_input[399]), .Z(n19805) );
  NAND U20835 ( .A(n12323), .B(e_input[399]), .Z(n19811) );
  XNOR U20836 ( .A(n19801), .B(n19812), .Z(n19803) );
  XOR U20837 ( .A(n19813), .B(n19814), .Z(n19801) );
  AND U20838 ( .A(n19815), .B(n19816), .Z(n19814) );
  XNOR U20839 ( .A(n19817), .B(n19813), .Z(n19816) );
  XOR U20840 ( .A(n19818), .B(e_input[399]), .Z(n19809) );
  IV U20841 ( .A(n19807), .Z(n19818) );
  XOR U20842 ( .A(n19819), .B(n19820), .Z(n19807) );
  AND U20843 ( .A(n19821), .B(n19822), .Z(n19820) );
  XNOR U20844 ( .A(n19819), .B(n9912), .Z(n19822) );
  XNOR U20845 ( .A(n19815), .B(n19817), .Z(n9912) );
  NAND U20846 ( .A(n19823), .B(e_input[398]), .Z(n19817) );
  NAND U20847 ( .A(n12323), .B(e_input[398]), .Z(n19823) );
  XNOR U20848 ( .A(n19813), .B(n19824), .Z(n19815) );
  XOR U20849 ( .A(n19825), .B(n19826), .Z(n19813) );
  AND U20850 ( .A(n19827), .B(n19828), .Z(n19826) );
  XNOR U20851 ( .A(n19829), .B(n19825), .Z(n19828) );
  XOR U20852 ( .A(n19830), .B(e_input[398]), .Z(n19821) );
  IV U20853 ( .A(n19819), .Z(n19830) );
  XOR U20854 ( .A(n19831), .B(n19832), .Z(n19819) );
  AND U20855 ( .A(n19833), .B(n19834), .Z(n19832) );
  XNOR U20856 ( .A(n19831), .B(n9918), .Z(n19834) );
  XNOR U20857 ( .A(n19827), .B(n19829), .Z(n9918) );
  NAND U20858 ( .A(n19835), .B(e_input[397]), .Z(n19829) );
  NAND U20859 ( .A(n12323), .B(e_input[397]), .Z(n19835) );
  XNOR U20860 ( .A(n19825), .B(n19836), .Z(n19827) );
  XOR U20861 ( .A(n19837), .B(n19838), .Z(n19825) );
  AND U20862 ( .A(n19839), .B(n19840), .Z(n19838) );
  XNOR U20863 ( .A(n19841), .B(n19837), .Z(n19840) );
  XOR U20864 ( .A(n19842), .B(e_input[397]), .Z(n19833) );
  IV U20865 ( .A(n19831), .Z(n19842) );
  XOR U20866 ( .A(n19843), .B(n19844), .Z(n19831) );
  AND U20867 ( .A(n19845), .B(n19846), .Z(n19844) );
  XNOR U20868 ( .A(n19843), .B(n9924), .Z(n19846) );
  XNOR U20869 ( .A(n19839), .B(n19841), .Z(n9924) );
  NAND U20870 ( .A(n19847), .B(e_input[396]), .Z(n19841) );
  NAND U20871 ( .A(n12323), .B(e_input[396]), .Z(n19847) );
  XNOR U20872 ( .A(n19837), .B(n19848), .Z(n19839) );
  XOR U20873 ( .A(n19849), .B(n19850), .Z(n19837) );
  AND U20874 ( .A(n19851), .B(n19852), .Z(n19850) );
  XNOR U20875 ( .A(n19853), .B(n19849), .Z(n19852) );
  XOR U20876 ( .A(n19854), .B(e_input[396]), .Z(n19845) );
  IV U20877 ( .A(n19843), .Z(n19854) );
  XOR U20878 ( .A(n19855), .B(n19856), .Z(n19843) );
  AND U20879 ( .A(n19857), .B(n19858), .Z(n19856) );
  XNOR U20880 ( .A(n19855), .B(n9930), .Z(n19858) );
  XNOR U20881 ( .A(n19851), .B(n19853), .Z(n9930) );
  NAND U20882 ( .A(n19859), .B(e_input[395]), .Z(n19853) );
  NAND U20883 ( .A(n12323), .B(e_input[395]), .Z(n19859) );
  XNOR U20884 ( .A(n19849), .B(n19860), .Z(n19851) );
  XOR U20885 ( .A(n19861), .B(n19862), .Z(n19849) );
  AND U20886 ( .A(n19863), .B(n19864), .Z(n19862) );
  XNOR U20887 ( .A(n19865), .B(n19861), .Z(n19864) );
  XOR U20888 ( .A(n19866), .B(e_input[395]), .Z(n19857) );
  IV U20889 ( .A(n19855), .Z(n19866) );
  XOR U20890 ( .A(n19867), .B(n19868), .Z(n19855) );
  AND U20891 ( .A(n19869), .B(n19870), .Z(n19868) );
  XNOR U20892 ( .A(n19867), .B(n9936), .Z(n19870) );
  XNOR U20893 ( .A(n19863), .B(n19865), .Z(n9936) );
  NAND U20894 ( .A(n19871), .B(e_input[394]), .Z(n19865) );
  NAND U20895 ( .A(n12323), .B(e_input[394]), .Z(n19871) );
  XNOR U20896 ( .A(n19861), .B(n19872), .Z(n19863) );
  XOR U20897 ( .A(n19873), .B(n19874), .Z(n19861) );
  AND U20898 ( .A(n19875), .B(n19876), .Z(n19874) );
  XNOR U20899 ( .A(n19877), .B(n19873), .Z(n19876) );
  XOR U20900 ( .A(n19878), .B(e_input[394]), .Z(n19869) );
  IV U20901 ( .A(n19867), .Z(n19878) );
  XOR U20902 ( .A(n19879), .B(n19880), .Z(n19867) );
  AND U20903 ( .A(n19881), .B(n19882), .Z(n19880) );
  XNOR U20904 ( .A(n19879), .B(n9942), .Z(n19882) );
  XNOR U20905 ( .A(n19875), .B(n19877), .Z(n9942) );
  NAND U20906 ( .A(n19883), .B(e_input[393]), .Z(n19877) );
  NAND U20907 ( .A(n12323), .B(e_input[393]), .Z(n19883) );
  XNOR U20908 ( .A(n19873), .B(n19884), .Z(n19875) );
  XOR U20909 ( .A(n19885), .B(n19886), .Z(n19873) );
  AND U20910 ( .A(n19887), .B(n19888), .Z(n19886) );
  XNOR U20911 ( .A(n19889), .B(n19885), .Z(n19888) );
  XOR U20912 ( .A(n19890), .B(e_input[393]), .Z(n19881) );
  IV U20913 ( .A(n19879), .Z(n19890) );
  XOR U20914 ( .A(n19891), .B(n19892), .Z(n19879) );
  AND U20915 ( .A(n19893), .B(n19894), .Z(n19892) );
  XNOR U20916 ( .A(n19891), .B(n9948), .Z(n19894) );
  XNOR U20917 ( .A(n19887), .B(n19889), .Z(n9948) );
  NAND U20918 ( .A(n19895), .B(e_input[392]), .Z(n19889) );
  NAND U20919 ( .A(n12323), .B(e_input[392]), .Z(n19895) );
  XNOR U20920 ( .A(n19885), .B(n19896), .Z(n19887) );
  XOR U20921 ( .A(n19897), .B(n19898), .Z(n19885) );
  AND U20922 ( .A(n19899), .B(n19900), .Z(n19898) );
  XNOR U20923 ( .A(n19901), .B(n19897), .Z(n19900) );
  XOR U20924 ( .A(n19902), .B(e_input[392]), .Z(n19893) );
  IV U20925 ( .A(n19891), .Z(n19902) );
  XOR U20926 ( .A(n19903), .B(n19904), .Z(n19891) );
  AND U20927 ( .A(n19905), .B(n19906), .Z(n19904) );
  XNOR U20928 ( .A(n19903), .B(n9954), .Z(n19906) );
  XNOR U20929 ( .A(n19899), .B(n19901), .Z(n9954) );
  NAND U20930 ( .A(n19907), .B(e_input[391]), .Z(n19901) );
  NAND U20931 ( .A(n12323), .B(e_input[391]), .Z(n19907) );
  XNOR U20932 ( .A(n19897), .B(n19908), .Z(n19899) );
  XOR U20933 ( .A(n19909), .B(n19910), .Z(n19897) );
  AND U20934 ( .A(n19911), .B(n19912), .Z(n19910) );
  XNOR U20935 ( .A(n19913), .B(n19909), .Z(n19912) );
  XOR U20936 ( .A(n19914), .B(e_input[391]), .Z(n19905) );
  IV U20937 ( .A(n19903), .Z(n19914) );
  XOR U20938 ( .A(n19915), .B(n19916), .Z(n19903) );
  AND U20939 ( .A(n19917), .B(n19918), .Z(n19916) );
  XNOR U20940 ( .A(n19915), .B(n9960), .Z(n19918) );
  XNOR U20941 ( .A(n19911), .B(n19913), .Z(n9960) );
  NAND U20942 ( .A(n19919), .B(e_input[390]), .Z(n19913) );
  NAND U20943 ( .A(n12323), .B(e_input[390]), .Z(n19919) );
  XNOR U20944 ( .A(n19909), .B(n19920), .Z(n19911) );
  XOR U20945 ( .A(n19921), .B(n19922), .Z(n19909) );
  AND U20946 ( .A(n19923), .B(n19924), .Z(n19922) );
  XNOR U20947 ( .A(n19925), .B(n19921), .Z(n19924) );
  XOR U20948 ( .A(n19926), .B(e_input[390]), .Z(n19917) );
  IV U20949 ( .A(n19915), .Z(n19926) );
  XOR U20950 ( .A(n19927), .B(n19928), .Z(n19915) );
  AND U20951 ( .A(n19929), .B(n19930), .Z(n19928) );
  XNOR U20952 ( .A(n19927), .B(n9966), .Z(n19930) );
  XNOR U20953 ( .A(n19923), .B(n19925), .Z(n9966) );
  NAND U20954 ( .A(n19931), .B(e_input[389]), .Z(n19925) );
  NAND U20955 ( .A(n12323), .B(e_input[389]), .Z(n19931) );
  XNOR U20956 ( .A(n19921), .B(n19932), .Z(n19923) );
  XOR U20957 ( .A(n19933), .B(n19934), .Z(n19921) );
  AND U20958 ( .A(n19935), .B(n19936), .Z(n19934) );
  XNOR U20959 ( .A(n19937), .B(n19933), .Z(n19936) );
  XOR U20960 ( .A(n19938), .B(e_input[389]), .Z(n19929) );
  IV U20961 ( .A(n19927), .Z(n19938) );
  XOR U20962 ( .A(n19939), .B(n19940), .Z(n19927) );
  AND U20963 ( .A(n19941), .B(n19942), .Z(n19940) );
  XNOR U20964 ( .A(n19939), .B(n9972), .Z(n19942) );
  XNOR U20965 ( .A(n19935), .B(n19937), .Z(n9972) );
  NAND U20966 ( .A(n19943), .B(e_input[388]), .Z(n19937) );
  NAND U20967 ( .A(n12323), .B(e_input[388]), .Z(n19943) );
  XNOR U20968 ( .A(n19933), .B(n19944), .Z(n19935) );
  XOR U20969 ( .A(n19945), .B(n19946), .Z(n19933) );
  AND U20970 ( .A(n19947), .B(n19948), .Z(n19946) );
  XNOR U20971 ( .A(n19949), .B(n19945), .Z(n19948) );
  XOR U20972 ( .A(n19950), .B(e_input[388]), .Z(n19941) );
  IV U20973 ( .A(n19939), .Z(n19950) );
  XOR U20974 ( .A(n19951), .B(n19952), .Z(n19939) );
  AND U20975 ( .A(n19953), .B(n19954), .Z(n19952) );
  XNOR U20976 ( .A(n19951), .B(n9978), .Z(n19954) );
  XNOR U20977 ( .A(n19947), .B(n19949), .Z(n9978) );
  NAND U20978 ( .A(n19955), .B(e_input[387]), .Z(n19949) );
  NAND U20979 ( .A(n12323), .B(e_input[387]), .Z(n19955) );
  XNOR U20980 ( .A(n19945), .B(n19956), .Z(n19947) );
  XOR U20981 ( .A(n19957), .B(n19958), .Z(n19945) );
  AND U20982 ( .A(n19959), .B(n19960), .Z(n19958) );
  XNOR U20983 ( .A(n19961), .B(n19957), .Z(n19960) );
  XOR U20984 ( .A(n19962), .B(e_input[387]), .Z(n19953) );
  IV U20985 ( .A(n19951), .Z(n19962) );
  XOR U20986 ( .A(n19963), .B(n19964), .Z(n19951) );
  AND U20987 ( .A(n19965), .B(n19966), .Z(n19964) );
  XNOR U20988 ( .A(n19963), .B(n9984), .Z(n19966) );
  XNOR U20989 ( .A(n19959), .B(n19961), .Z(n9984) );
  NAND U20990 ( .A(n19967), .B(e_input[386]), .Z(n19961) );
  NAND U20991 ( .A(n12323), .B(e_input[386]), .Z(n19967) );
  XNOR U20992 ( .A(n19957), .B(n19968), .Z(n19959) );
  XOR U20993 ( .A(n19969), .B(n19970), .Z(n19957) );
  AND U20994 ( .A(n19971), .B(n19972), .Z(n19970) );
  XNOR U20995 ( .A(n19973), .B(n19969), .Z(n19972) );
  XOR U20996 ( .A(n19974), .B(e_input[386]), .Z(n19965) );
  IV U20997 ( .A(n19963), .Z(n19974) );
  XOR U20998 ( .A(n19975), .B(n19976), .Z(n19963) );
  AND U20999 ( .A(n19977), .B(n19978), .Z(n19976) );
  XNOR U21000 ( .A(n19975), .B(n9990), .Z(n19978) );
  XNOR U21001 ( .A(n19971), .B(n19973), .Z(n9990) );
  NAND U21002 ( .A(n19979), .B(e_input[385]), .Z(n19973) );
  NAND U21003 ( .A(n12323), .B(e_input[385]), .Z(n19979) );
  XNOR U21004 ( .A(n19969), .B(n19980), .Z(n19971) );
  XOR U21005 ( .A(n19981), .B(n19982), .Z(n19969) );
  AND U21006 ( .A(n19983), .B(n19984), .Z(n19982) );
  XNOR U21007 ( .A(n19985), .B(n19981), .Z(n19984) );
  XOR U21008 ( .A(n19986), .B(e_input[385]), .Z(n19977) );
  IV U21009 ( .A(n19975), .Z(n19986) );
  XOR U21010 ( .A(n19987), .B(n19988), .Z(n19975) );
  AND U21011 ( .A(n19989), .B(n19990), .Z(n19988) );
  XNOR U21012 ( .A(n19987), .B(n9996), .Z(n19990) );
  XNOR U21013 ( .A(n19983), .B(n19985), .Z(n9996) );
  NAND U21014 ( .A(n19991), .B(e_input[384]), .Z(n19985) );
  NAND U21015 ( .A(n12323), .B(e_input[384]), .Z(n19991) );
  XNOR U21016 ( .A(n19981), .B(n19992), .Z(n19983) );
  XOR U21017 ( .A(n19993), .B(n19994), .Z(n19981) );
  AND U21018 ( .A(n19995), .B(n19996), .Z(n19994) );
  XNOR U21019 ( .A(n19997), .B(n19993), .Z(n19996) );
  XOR U21020 ( .A(n19998), .B(e_input[384]), .Z(n19989) );
  IV U21021 ( .A(n19987), .Z(n19998) );
  XOR U21022 ( .A(n19999), .B(n20000), .Z(n19987) );
  AND U21023 ( .A(n20001), .B(n20002), .Z(n20000) );
  XNOR U21024 ( .A(n19999), .B(n10002), .Z(n20002) );
  XNOR U21025 ( .A(n19995), .B(n19997), .Z(n10002) );
  NAND U21026 ( .A(n20003), .B(e_input[383]), .Z(n19997) );
  NAND U21027 ( .A(n12323), .B(e_input[383]), .Z(n20003) );
  XNOR U21028 ( .A(n19993), .B(n20004), .Z(n19995) );
  XOR U21029 ( .A(n20005), .B(n20006), .Z(n19993) );
  AND U21030 ( .A(n20007), .B(n20008), .Z(n20006) );
  XNOR U21031 ( .A(n20009), .B(n20005), .Z(n20008) );
  XOR U21032 ( .A(n20010), .B(e_input[383]), .Z(n20001) );
  IV U21033 ( .A(n19999), .Z(n20010) );
  XOR U21034 ( .A(n20011), .B(n20012), .Z(n19999) );
  AND U21035 ( .A(n20013), .B(n20014), .Z(n20012) );
  XNOR U21036 ( .A(n20011), .B(n10008), .Z(n20014) );
  XNOR U21037 ( .A(n20007), .B(n20009), .Z(n10008) );
  NAND U21038 ( .A(n20015), .B(e_input[382]), .Z(n20009) );
  NAND U21039 ( .A(n12323), .B(e_input[382]), .Z(n20015) );
  XNOR U21040 ( .A(n20005), .B(n20016), .Z(n20007) );
  XOR U21041 ( .A(n20017), .B(n20018), .Z(n20005) );
  AND U21042 ( .A(n20019), .B(n20020), .Z(n20018) );
  XNOR U21043 ( .A(n20021), .B(n20017), .Z(n20020) );
  XOR U21044 ( .A(n20022), .B(e_input[382]), .Z(n20013) );
  IV U21045 ( .A(n20011), .Z(n20022) );
  XOR U21046 ( .A(n20023), .B(n20024), .Z(n20011) );
  AND U21047 ( .A(n20025), .B(n20026), .Z(n20024) );
  XNOR U21048 ( .A(n20023), .B(n10014), .Z(n20026) );
  XNOR U21049 ( .A(n20019), .B(n20021), .Z(n10014) );
  NAND U21050 ( .A(n20027), .B(e_input[381]), .Z(n20021) );
  NAND U21051 ( .A(n12323), .B(e_input[381]), .Z(n20027) );
  XNOR U21052 ( .A(n20017), .B(n20028), .Z(n20019) );
  XOR U21053 ( .A(n20029), .B(n20030), .Z(n20017) );
  AND U21054 ( .A(n20031), .B(n20032), .Z(n20030) );
  XNOR U21055 ( .A(n20033), .B(n20029), .Z(n20032) );
  XOR U21056 ( .A(n20034), .B(e_input[381]), .Z(n20025) );
  IV U21057 ( .A(n20023), .Z(n20034) );
  XOR U21058 ( .A(n20035), .B(n20036), .Z(n20023) );
  AND U21059 ( .A(n20037), .B(n20038), .Z(n20036) );
  XNOR U21060 ( .A(n20035), .B(n10020), .Z(n20038) );
  XNOR U21061 ( .A(n20031), .B(n20033), .Z(n10020) );
  NAND U21062 ( .A(n20039), .B(e_input[380]), .Z(n20033) );
  NAND U21063 ( .A(n12323), .B(e_input[380]), .Z(n20039) );
  XNOR U21064 ( .A(n20029), .B(n20040), .Z(n20031) );
  XOR U21065 ( .A(n20041), .B(n20042), .Z(n20029) );
  AND U21066 ( .A(n20043), .B(n20044), .Z(n20042) );
  XNOR U21067 ( .A(n20045), .B(n20041), .Z(n20044) );
  XOR U21068 ( .A(n20046), .B(e_input[380]), .Z(n20037) );
  IV U21069 ( .A(n20035), .Z(n20046) );
  XOR U21070 ( .A(n20047), .B(n20048), .Z(n20035) );
  AND U21071 ( .A(n20049), .B(n20050), .Z(n20048) );
  XNOR U21072 ( .A(n20047), .B(n10026), .Z(n20050) );
  XNOR U21073 ( .A(n20043), .B(n20045), .Z(n10026) );
  NAND U21074 ( .A(n20051), .B(e_input[379]), .Z(n20045) );
  NAND U21075 ( .A(n12323), .B(e_input[379]), .Z(n20051) );
  XNOR U21076 ( .A(n20041), .B(n20052), .Z(n20043) );
  XOR U21077 ( .A(n20053), .B(n20054), .Z(n20041) );
  AND U21078 ( .A(n20055), .B(n20056), .Z(n20054) );
  XNOR U21079 ( .A(n20057), .B(n20053), .Z(n20056) );
  XOR U21080 ( .A(n20058), .B(e_input[379]), .Z(n20049) );
  IV U21081 ( .A(n20047), .Z(n20058) );
  XOR U21082 ( .A(n20059), .B(n20060), .Z(n20047) );
  AND U21083 ( .A(n20061), .B(n20062), .Z(n20060) );
  XNOR U21084 ( .A(n20059), .B(n10032), .Z(n20062) );
  XNOR U21085 ( .A(n20055), .B(n20057), .Z(n10032) );
  NAND U21086 ( .A(n20063), .B(e_input[378]), .Z(n20057) );
  NAND U21087 ( .A(n12323), .B(e_input[378]), .Z(n20063) );
  XNOR U21088 ( .A(n20053), .B(n20064), .Z(n20055) );
  XOR U21089 ( .A(n20065), .B(n20066), .Z(n20053) );
  AND U21090 ( .A(n20067), .B(n20068), .Z(n20066) );
  XNOR U21091 ( .A(n20069), .B(n20065), .Z(n20068) );
  XOR U21092 ( .A(n20070), .B(e_input[378]), .Z(n20061) );
  IV U21093 ( .A(n20059), .Z(n20070) );
  XOR U21094 ( .A(n20071), .B(n20072), .Z(n20059) );
  AND U21095 ( .A(n20073), .B(n20074), .Z(n20072) );
  XNOR U21096 ( .A(n20071), .B(n10038), .Z(n20074) );
  XNOR U21097 ( .A(n20067), .B(n20069), .Z(n10038) );
  NAND U21098 ( .A(n20075), .B(e_input[377]), .Z(n20069) );
  NAND U21099 ( .A(n12323), .B(e_input[377]), .Z(n20075) );
  XNOR U21100 ( .A(n20065), .B(n20076), .Z(n20067) );
  XOR U21101 ( .A(n20077), .B(n20078), .Z(n20065) );
  AND U21102 ( .A(n20079), .B(n20080), .Z(n20078) );
  XNOR U21103 ( .A(n20081), .B(n20077), .Z(n20080) );
  XOR U21104 ( .A(n20082), .B(e_input[377]), .Z(n20073) );
  IV U21105 ( .A(n20071), .Z(n20082) );
  XOR U21106 ( .A(n20083), .B(n20084), .Z(n20071) );
  AND U21107 ( .A(n20085), .B(n20086), .Z(n20084) );
  XNOR U21108 ( .A(n20083), .B(n10044), .Z(n20086) );
  XNOR U21109 ( .A(n20079), .B(n20081), .Z(n10044) );
  NAND U21110 ( .A(n20087), .B(e_input[376]), .Z(n20081) );
  NAND U21111 ( .A(n12323), .B(e_input[376]), .Z(n20087) );
  XNOR U21112 ( .A(n20077), .B(n20088), .Z(n20079) );
  XOR U21113 ( .A(n20089), .B(n20090), .Z(n20077) );
  AND U21114 ( .A(n20091), .B(n20092), .Z(n20090) );
  XNOR U21115 ( .A(n20093), .B(n20089), .Z(n20092) );
  XOR U21116 ( .A(n20094), .B(e_input[376]), .Z(n20085) );
  IV U21117 ( .A(n20083), .Z(n20094) );
  XOR U21118 ( .A(n20095), .B(n20096), .Z(n20083) );
  AND U21119 ( .A(n20097), .B(n20098), .Z(n20096) );
  XNOR U21120 ( .A(n20095), .B(n10050), .Z(n20098) );
  XNOR U21121 ( .A(n20091), .B(n20093), .Z(n10050) );
  NAND U21122 ( .A(n20099), .B(e_input[375]), .Z(n20093) );
  NAND U21123 ( .A(n12323), .B(e_input[375]), .Z(n20099) );
  XNOR U21124 ( .A(n20089), .B(n20100), .Z(n20091) );
  XOR U21125 ( .A(n20101), .B(n20102), .Z(n20089) );
  AND U21126 ( .A(n20103), .B(n20104), .Z(n20102) );
  XNOR U21127 ( .A(n20105), .B(n20101), .Z(n20104) );
  XOR U21128 ( .A(n20106), .B(e_input[375]), .Z(n20097) );
  IV U21129 ( .A(n20095), .Z(n20106) );
  XOR U21130 ( .A(n20107), .B(n20108), .Z(n20095) );
  AND U21131 ( .A(n20109), .B(n20110), .Z(n20108) );
  XNOR U21132 ( .A(n20107), .B(n10056), .Z(n20110) );
  XNOR U21133 ( .A(n20103), .B(n20105), .Z(n10056) );
  NAND U21134 ( .A(n20111), .B(e_input[374]), .Z(n20105) );
  NAND U21135 ( .A(n12323), .B(e_input[374]), .Z(n20111) );
  XNOR U21136 ( .A(n20101), .B(n20112), .Z(n20103) );
  XOR U21137 ( .A(n20113), .B(n20114), .Z(n20101) );
  AND U21138 ( .A(n20115), .B(n20116), .Z(n20114) );
  XNOR U21139 ( .A(n20117), .B(n20113), .Z(n20116) );
  XOR U21140 ( .A(n20118), .B(e_input[374]), .Z(n20109) );
  IV U21141 ( .A(n20107), .Z(n20118) );
  XOR U21142 ( .A(n20119), .B(n20120), .Z(n20107) );
  AND U21143 ( .A(n20121), .B(n20122), .Z(n20120) );
  XNOR U21144 ( .A(n20119), .B(n10062), .Z(n20122) );
  XNOR U21145 ( .A(n20115), .B(n20117), .Z(n10062) );
  NAND U21146 ( .A(n20123), .B(e_input[373]), .Z(n20117) );
  NAND U21147 ( .A(n12323), .B(e_input[373]), .Z(n20123) );
  XNOR U21148 ( .A(n20113), .B(n20124), .Z(n20115) );
  XOR U21149 ( .A(n20125), .B(n20126), .Z(n20113) );
  AND U21150 ( .A(n20127), .B(n20128), .Z(n20126) );
  XNOR U21151 ( .A(n20129), .B(n20125), .Z(n20128) );
  XOR U21152 ( .A(n20130), .B(e_input[373]), .Z(n20121) );
  IV U21153 ( .A(n20119), .Z(n20130) );
  XOR U21154 ( .A(n20131), .B(n20132), .Z(n20119) );
  AND U21155 ( .A(n20133), .B(n20134), .Z(n20132) );
  XNOR U21156 ( .A(n20131), .B(n10068), .Z(n20134) );
  XNOR U21157 ( .A(n20127), .B(n20129), .Z(n10068) );
  NAND U21158 ( .A(n20135), .B(e_input[372]), .Z(n20129) );
  NAND U21159 ( .A(n12323), .B(e_input[372]), .Z(n20135) );
  XNOR U21160 ( .A(n20125), .B(n20136), .Z(n20127) );
  XOR U21161 ( .A(n20137), .B(n20138), .Z(n20125) );
  AND U21162 ( .A(n20139), .B(n20140), .Z(n20138) );
  XNOR U21163 ( .A(n20141), .B(n20137), .Z(n20140) );
  XOR U21164 ( .A(n20142), .B(e_input[372]), .Z(n20133) );
  IV U21165 ( .A(n20131), .Z(n20142) );
  XOR U21166 ( .A(n20143), .B(n20144), .Z(n20131) );
  AND U21167 ( .A(n20145), .B(n20146), .Z(n20144) );
  XNOR U21168 ( .A(n20143), .B(n10074), .Z(n20146) );
  XNOR U21169 ( .A(n20139), .B(n20141), .Z(n10074) );
  NAND U21170 ( .A(n20147), .B(e_input[371]), .Z(n20141) );
  NAND U21171 ( .A(n12323), .B(e_input[371]), .Z(n20147) );
  XNOR U21172 ( .A(n20137), .B(n20148), .Z(n20139) );
  XOR U21173 ( .A(n20149), .B(n20150), .Z(n20137) );
  AND U21174 ( .A(n20151), .B(n20152), .Z(n20150) );
  XNOR U21175 ( .A(n20153), .B(n20149), .Z(n20152) );
  XOR U21176 ( .A(n20154), .B(e_input[371]), .Z(n20145) );
  IV U21177 ( .A(n20143), .Z(n20154) );
  XOR U21178 ( .A(n20155), .B(n20156), .Z(n20143) );
  AND U21179 ( .A(n20157), .B(n20158), .Z(n20156) );
  XNOR U21180 ( .A(n20155), .B(n10080), .Z(n20158) );
  XNOR U21181 ( .A(n20151), .B(n20153), .Z(n10080) );
  NAND U21182 ( .A(n20159), .B(e_input[370]), .Z(n20153) );
  NAND U21183 ( .A(n12323), .B(e_input[370]), .Z(n20159) );
  XNOR U21184 ( .A(n20149), .B(n20160), .Z(n20151) );
  XOR U21185 ( .A(n20161), .B(n20162), .Z(n20149) );
  AND U21186 ( .A(n20163), .B(n20164), .Z(n20162) );
  XNOR U21187 ( .A(n20165), .B(n20161), .Z(n20164) );
  XOR U21188 ( .A(n20166), .B(e_input[370]), .Z(n20157) );
  IV U21189 ( .A(n20155), .Z(n20166) );
  XOR U21190 ( .A(n20167), .B(n20168), .Z(n20155) );
  AND U21191 ( .A(n20169), .B(n20170), .Z(n20168) );
  XNOR U21192 ( .A(n20167), .B(n10086), .Z(n20170) );
  XNOR U21193 ( .A(n20163), .B(n20165), .Z(n10086) );
  NAND U21194 ( .A(n20171), .B(e_input[369]), .Z(n20165) );
  NAND U21195 ( .A(n12323), .B(e_input[369]), .Z(n20171) );
  XNOR U21196 ( .A(n20161), .B(n20172), .Z(n20163) );
  XOR U21197 ( .A(n20173), .B(n20174), .Z(n20161) );
  AND U21198 ( .A(n20175), .B(n20176), .Z(n20174) );
  XNOR U21199 ( .A(n20177), .B(n20173), .Z(n20176) );
  XOR U21200 ( .A(n20178), .B(e_input[369]), .Z(n20169) );
  IV U21201 ( .A(n20167), .Z(n20178) );
  XOR U21202 ( .A(n20179), .B(n20180), .Z(n20167) );
  AND U21203 ( .A(n20181), .B(n20182), .Z(n20180) );
  XNOR U21204 ( .A(n20179), .B(n10092), .Z(n20182) );
  XNOR U21205 ( .A(n20175), .B(n20177), .Z(n10092) );
  NAND U21206 ( .A(n20183), .B(e_input[368]), .Z(n20177) );
  NAND U21207 ( .A(n12323), .B(e_input[368]), .Z(n20183) );
  XNOR U21208 ( .A(n20173), .B(n20184), .Z(n20175) );
  XOR U21209 ( .A(n20185), .B(n20186), .Z(n20173) );
  AND U21210 ( .A(n20187), .B(n20188), .Z(n20186) );
  XNOR U21211 ( .A(n20189), .B(n20185), .Z(n20188) );
  XOR U21212 ( .A(n20190), .B(e_input[368]), .Z(n20181) );
  IV U21213 ( .A(n20179), .Z(n20190) );
  XOR U21214 ( .A(n20191), .B(n20192), .Z(n20179) );
  AND U21215 ( .A(n20193), .B(n20194), .Z(n20192) );
  XNOR U21216 ( .A(n20191), .B(n10098), .Z(n20194) );
  XNOR U21217 ( .A(n20187), .B(n20189), .Z(n10098) );
  NAND U21218 ( .A(n20195), .B(e_input[367]), .Z(n20189) );
  NAND U21219 ( .A(n12323), .B(e_input[367]), .Z(n20195) );
  XNOR U21220 ( .A(n20185), .B(n20196), .Z(n20187) );
  XOR U21221 ( .A(n20197), .B(n20198), .Z(n20185) );
  AND U21222 ( .A(n20199), .B(n20200), .Z(n20198) );
  XNOR U21223 ( .A(n20201), .B(n20197), .Z(n20200) );
  XOR U21224 ( .A(n20202), .B(e_input[367]), .Z(n20193) );
  IV U21225 ( .A(n20191), .Z(n20202) );
  XOR U21226 ( .A(n20203), .B(n20204), .Z(n20191) );
  AND U21227 ( .A(n20205), .B(n20206), .Z(n20204) );
  XNOR U21228 ( .A(n20203), .B(n10104), .Z(n20206) );
  XNOR U21229 ( .A(n20199), .B(n20201), .Z(n10104) );
  NAND U21230 ( .A(n20207), .B(e_input[366]), .Z(n20201) );
  NAND U21231 ( .A(n12323), .B(e_input[366]), .Z(n20207) );
  XNOR U21232 ( .A(n20197), .B(n20208), .Z(n20199) );
  XOR U21233 ( .A(n20209), .B(n20210), .Z(n20197) );
  AND U21234 ( .A(n20211), .B(n20212), .Z(n20210) );
  XNOR U21235 ( .A(n20213), .B(n20209), .Z(n20212) );
  XOR U21236 ( .A(n20214), .B(e_input[366]), .Z(n20205) );
  IV U21237 ( .A(n20203), .Z(n20214) );
  XOR U21238 ( .A(n20215), .B(n20216), .Z(n20203) );
  AND U21239 ( .A(n20217), .B(n20218), .Z(n20216) );
  XNOR U21240 ( .A(n20215), .B(n10110), .Z(n20218) );
  XNOR U21241 ( .A(n20211), .B(n20213), .Z(n10110) );
  NAND U21242 ( .A(n20219), .B(e_input[365]), .Z(n20213) );
  NAND U21243 ( .A(n12323), .B(e_input[365]), .Z(n20219) );
  XNOR U21244 ( .A(n20209), .B(n20220), .Z(n20211) );
  XOR U21245 ( .A(n20221), .B(n20222), .Z(n20209) );
  AND U21246 ( .A(n20223), .B(n20224), .Z(n20222) );
  XNOR U21247 ( .A(n20225), .B(n20221), .Z(n20224) );
  XOR U21248 ( .A(n20226), .B(e_input[365]), .Z(n20217) );
  IV U21249 ( .A(n20215), .Z(n20226) );
  XOR U21250 ( .A(n20227), .B(n20228), .Z(n20215) );
  AND U21251 ( .A(n20229), .B(n20230), .Z(n20228) );
  XNOR U21252 ( .A(n20227), .B(n10116), .Z(n20230) );
  XNOR U21253 ( .A(n20223), .B(n20225), .Z(n10116) );
  NAND U21254 ( .A(n20231), .B(e_input[364]), .Z(n20225) );
  NAND U21255 ( .A(n12323), .B(e_input[364]), .Z(n20231) );
  XNOR U21256 ( .A(n20221), .B(n20232), .Z(n20223) );
  XOR U21257 ( .A(n20233), .B(n20234), .Z(n20221) );
  AND U21258 ( .A(n20235), .B(n20236), .Z(n20234) );
  XNOR U21259 ( .A(n20237), .B(n20233), .Z(n20236) );
  XOR U21260 ( .A(n20238), .B(e_input[364]), .Z(n20229) );
  IV U21261 ( .A(n20227), .Z(n20238) );
  XOR U21262 ( .A(n20239), .B(n20240), .Z(n20227) );
  AND U21263 ( .A(n20241), .B(n20242), .Z(n20240) );
  XNOR U21264 ( .A(n20239), .B(n10122), .Z(n20242) );
  XNOR U21265 ( .A(n20235), .B(n20237), .Z(n10122) );
  NAND U21266 ( .A(n20243), .B(e_input[363]), .Z(n20237) );
  NAND U21267 ( .A(n12323), .B(e_input[363]), .Z(n20243) );
  XNOR U21268 ( .A(n20233), .B(n20244), .Z(n20235) );
  XOR U21269 ( .A(n20245), .B(n20246), .Z(n20233) );
  AND U21270 ( .A(n20247), .B(n20248), .Z(n20246) );
  XNOR U21271 ( .A(n20249), .B(n20245), .Z(n20248) );
  XOR U21272 ( .A(n20250), .B(e_input[363]), .Z(n20241) );
  IV U21273 ( .A(n20239), .Z(n20250) );
  XOR U21274 ( .A(n20251), .B(n20252), .Z(n20239) );
  AND U21275 ( .A(n20253), .B(n20254), .Z(n20252) );
  XNOR U21276 ( .A(n20251), .B(n10128), .Z(n20254) );
  XNOR U21277 ( .A(n20247), .B(n20249), .Z(n10128) );
  NAND U21278 ( .A(n20255), .B(e_input[362]), .Z(n20249) );
  NAND U21279 ( .A(n12323), .B(e_input[362]), .Z(n20255) );
  XNOR U21280 ( .A(n20245), .B(n20256), .Z(n20247) );
  XOR U21281 ( .A(n20257), .B(n20258), .Z(n20245) );
  AND U21282 ( .A(n20259), .B(n20260), .Z(n20258) );
  XNOR U21283 ( .A(n20261), .B(n20257), .Z(n20260) );
  XOR U21284 ( .A(n20262), .B(e_input[362]), .Z(n20253) );
  IV U21285 ( .A(n20251), .Z(n20262) );
  XOR U21286 ( .A(n20263), .B(n20264), .Z(n20251) );
  AND U21287 ( .A(n20265), .B(n20266), .Z(n20264) );
  XNOR U21288 ( .A(n20263), .B(n10134), .Z(n20266) );
  XNOR U21289 ( .A(n20259), .B(n20261), .Z(n10134) );
  NAND U21290 ( .A(n20267), .B(e_input[361]), .Z(n20261) );
  NAND U21291 ( .A(n12323), .B(e_input[361]), .Z(n20267) );
  XNOR U21292 ( .A(n20257), .B(n20268), .Z(n20259) );
  XOR U21293 ( .A(n20269), .B(n20270), .Z(n20257) );
  AND U21294 ( .A(n20271), .B(n20272), .Z(n20270) );
  XNOR U21295 ( .A(n20273), .B(n20269), .Z(n20272) );
  XOR U21296 ( .A(n20274), .B(e_input[361]), .Z(n20265) );
  IV U21297 ( .A(n20263), .Z(n20274) );
  XOR U21298 ( .A(n20275), .B(n20276), .Z(n20263) );
  AND U21299 ( .A(n20277), .B(n20278), .Z(n20276) );
  XNOR U21300 ( .A(n20275), .B(n10140), .Z(n20278) );
  XNOR U21301 ( .A(n20271), .B(n20273), .Z(n10140) );
  NAND U21302 ( .A(n20279), .B(e_input[360]), .Z(n20273) );
  NAND U21303 ( .A(n12323), .B(e_input[360]), .Z(n20279) );
  XNOR U21304 ( .A(n20269), .B(n20280), .Z(n20271) );
  XOR U21305 ( .A(n20281), .B(n20282), .Z(n20269) );
  AND U21306 ( .A(n20283), .B(n20284), .Z(n20282) );
  XNOR U21307 ( .A(n20285), .B(n20281), .Z(n20284) );
  XOR U21308 ( .A(n20286), .B(e_input[360]), .Z(n20277) );
  IV U21309 ( .A(n20275), .Z(n20286) );
  XOR U21310 ( .A(n20287), .B(n20288), .Z(n20275) );
  AND U21311 ( .A(n20289), .B(n20290), .Z(n20288) );
  XNOR U21312 ( .A(n20287), .B(n10146), .Z(n20290) );
  XNOR U21313 ( .A(n20283), .B(n20285), .Z(n10146) );
  NAND U21314 ( .A(n20291), .B(e_input[359]), .Z(n20285) );
  NAND U21315 ( .A(n12323), .B(e_input[359]), .Z(n20291) );
  XNOR U21316 ( .A(n20281), .B(n20292), .Z(n20283) );
  XOR U21317 ( .A(n20293), .B(n20294), .Z(n20281) );
  AND U21318 ( .A(n20295), .B(n20296), .Z(n20294) );
  XNOR U21319 ( .A(n20297), .B(n20293), .Z(n20296) );
  XOR U21320 ( .A(n20298), .B(e_input[359]), .Z(n20289) );
  IV U21321 ( .A(n20287), .Z(n20298) );
  XOR U21322 ( .A(n20299), .B(n20300), .Z(n20287) );
  AND U21323 ( .A(n20301), .B(n20302), .Z(n20300) );
  XNOR U21324 ( .A(n20299), .B(n10152), .Z(n20302) );
  XNOR U21325 ( .A(n20295), .B(n20297), .Z(n10152) );
  NAND U21326 ( .A(n20303), .B(e_input[358]), .Z(n20297) );
  NAND U21327 ( .A(n12323), .B(e_input[358]), .Z(n20303) );
  XNOR U21328 ( .A(n20293), .B(n20304), .Z(n20295) );
  XOR U21329 ( .A(n20305), .B(n20306), .Z(n20293) );
  AND U21330 ( .A(n20307), .B(n20308), .Z(n20306) );
  XNOR U21331 ( .A(n20309), .B(n20305), .Z(n20308) );
  XOR U21332 ( .A(n20310), .B(e_input[358]), .Z(n20301) );
  IV U21333 ( .A(n20299), .Z(n20310) );
  XOR U21334 ( .A(n20311), .B(n20312), .Z(n20299) );
  AND U21335 ( .A(n20313), .B(n20314), .Z(n20312) );
  XNOR U21336 ( .A(n20311), .B(n10158), .Z(n20314) );
  XNOR U21337 ( .A(n20307), .B(n20309), .Z(n10158) );
  NAND U21338 ( .A(n20315), .B(e_input[357]), .Z(n20309) );
  NAND U21339 ( .A(n12323), .B(e_input[357]), .Z(n20315) );
  XNOR U21340 ( .A(n20305), .B(n20316), .Z(n20307) );
  XOR U21341 ( .A(n20317), .B(n20318), .Z(n20305) );
  AND U21342 ( .A(n20319), .B(n20320), .Z(n20318) );
  XNOR U21343 ( .A(n20321), .B(n20317), .Z(n20320) );
  XOR U21344 ( .A(n20322), .B(e_input[357]), .Z(n20313) );
  IV U21345 ( .A(n20311), .Z(n20322) );
  XOR U21346 ( .A(n20323), .B(n20324), .Z(n20311) );
  AND U21347 ( .A(n20325), .B(n20326), .Z(n20324) );
  XNOR U21348 ( .A(n20323), .B(n10164), .Z(n20326) );
  XNOR U21349 ( .A(n20319), .B(n20321), .Z(n10164) );
  NAND U21350 ( .A(n20327), .B(e_input[356]), .Z(n20321) );
  NAND U21351 ( .A(n12323), .B(e_input[356]), .Z(n20327) );
  XNOR U21352 ( .A(n20317), .B(n20328), .Z(n20319) );
  XOR U21353 ( .A(n20329), .B(n20330), .Z(n20317) );
  AND U21354 ( .A(n20331), .B(n20332), .Z(n20330) );
  XNOR U21355 ( .A(n20333), .B(n20329), .Z(n20332) );
  XOR U21356 ( .A(n20334), .B(e_input[356]), .Z(n20325) );
  IV U21357 ( .A(n20323), .Z(n20334) );
  XOR U21358 ( .A(n20335), .B(n20336), .Z(n20323) );
  AND U21359 ( .A(n20337), .B(n20338), .Z(n20336) );
  XNOR U21360 ( .A(n20335), .B(n10170), .Z(n20338) );
  XNOR U21361 ( .A(n20331), .B(n20333), .Z(n10170) );
  NAND U21362 ( .A(n20339), .B(e_input[355]), .Z(n20333) );
  NAND U21363 ( .A(n12323), .B(e_input[355]), .Z(n20339) );
  XNOR U21364 ( .A(n20329), .B(n20340), .Z(n20331) );
  XOR U21365 ( .A(n20341), .B(n20342), .Z(n20329) );
  AND U21366 ( .A(n20343), .B(n20344), .Z(n20342) );
  XNOR U21367 ( .A(n20345), .B(n20341), .Z(n20344) );
  XOR U21368 ( .A(n20346), .B(e_input[355]), .Z(n20337) );
  IV U21369 ( .A(n20335), .Z(n20346) );
  XOR U21370 ( .A(n20347), .B(n20348), .Z(n20335) );
  AND U21371 ( .A(n20349), .B(n20350), .Z(n20348) );
  XNOR U21372 ( .A(n20347), .B(n10176), .Z(n20350) );
  XNOR U21373 ( .A(n20343), .B(n20345), .Z(n10176) );
  NAND U21374 ( .A(n20351), .B(e_input[354]), .Z(n20345) );
  NAND U21375 ( .A(n12323), .B(e_input[354]), .Z(n20351) );
  XNOR U21376 ( .A(n20341), .B(n20352), .Z(n20343) );
  XOR U21377 ( .A(n20353), .B(n20354), .Z(n20341) );
  AND U21378 ( .A(n20355), .B(n20356), .Z(n20354) );
  XNOR U21379 ( .A(n20357), .B(n20353), .Z(n20356) );
  XOR U21380 ( .A(n20358), .B(e_input[354]), .Z(n20349) );
  IV U21381 ( .A(n20347), .Z(n20358) );
  XOR U21382 ( .A(n20359), .B(n20360), .Z(n20347) );
  AND U21383 ( .A(n20361), .B(n20362), .Z(n20360) );
  XNOR U21384 ( .A(n20359), .B(n10182), .Z(n20362) );
  XNOR U21385 ( .A(n20355), .B(n20357), .Z(n10182) );
  NAND U21386 ( .A(n20363), .B(e_input[353]), .Z(n20357) );
  NAND U21387 ( .A(n12323), .B(e_input[353]), .Z(n20363) );
  XNOR U21388 ( .A(n20353), .B(n20364), .Z(n20355) );
  XOR U21389 ( .A(n20365), .B(n20366), .Z(n20353) );
  AND U21390 ( .A(n20367), .B(n20368), .Z(n20366) );
  XNOR U21391 ( .A(n20369), .B(n20365), .Z(n20368) );
  XOR U21392 ( .A(n20370), .B(e_input[353]), .Z(n20361) );
  IV U21393 ( .A(n20359), .Z(n20370) );
  XOR U21394 ( .A(n20371), .B(n20372), .Z(n20359) );
  AND U21395 ( .A(n20373), .B(n20374), .Z(n20372) );
  XNOR U21396 ( .A(n20371), .B(n10188), .Z(n20374) );
  XNOR U21397 ( .A(n20367), .B(n20369), .Z(n10188) );
  NAND U21398 ( .A(n20375), .B(e_input[352]), .Z(n20369) );
  NAND U21399 ( .A(n12323), .B(e_input[352]), .Z(n20375) );
  XNOR U21400 ( .A(n20365), .B(n20376), .Z(n20367) );
  XOR U21401 ( .A(n20377), .B(n20378), .Z(n20365) );
  AND U21402 ( .A(n20379), .B(n20380), .Z(n20378) );
  XNOR U21403 ( .A(n20381), .B(n20377), .Z(n20380) );
  XOR U21404 ( .A(n20382), .B(e_input[352]), .Z(n20373) );
  IV U21405 ( .A(n20371), .Z(n20382) );
  XOR U21406 ( .A(n20383), .B(n20384), .Z(n20371) );
  AND U21407 ( .A(n20385), .B(n20386), .Z(n20384) );
  XNOR U21408 ( .A(n20383), .B(n10194), .Z(n20386) );
  XNOR U21409 ( .A(n20379), .B(n20381), .Z(n10194) );
  NAND U21410 ( .A(n20387), .B(e_input[351]), .Z(n20381) );
  NAND U21411 ( .A(n12323), .B(e_input[351]), .Z(n20387) );
  XNOR U21412 ( .A(n20377), .B(n20388), .Z(n20379) );
  XOR U21413 ( .A(n20389), .B(n20390), .Z(n20377) );
  AND U21414 ( .A(n20391), .B(n20392), .Z(n20390) );
  XNOR U21415 ( .A(n20393), .B(n20389), .Z(n20392) );
  XOR U21416 ( .A(n20394), .B(e_input[351]), .Z(n20385) );
  IV U21417 ( .A(n20383), .Z(n20394) );
  XOR U21418 ( .A(n20395), .B(n20396), .Z(n20383) );
  AND U21419 ( .A(n20397), .B(n20398), .Z(n20396) );
  XNOR U21420 ( .A(n20395), .B(n10200), .Z(n20398) );
  XNOR U21421 ( .A(n20391), .B(n20393), .Z(n10200) );
  NAND U21422 ( .A(n20399), .B(e_input[350]), .Z(n20393) );
  NAND U21423 ( .A(n12323), .B(e_input[350]), .Z(n20399) );
  XNOR U21424 ( .A(n20389), .B(n20400), .Z(n20391) );
  XOR U21425 ( .A(n20401), .B(n20402), .Z(n20389) );
  AND U21426 ( .A(n20403), .B(n20404), .Z(n20402) );
  XNOR U21427 ( .A(n20405), .B(n20401), .Z(n20404) );
  XOR U21428 ( .A(n20406), .B(e_input[350]), .Z(n20397) );
  IV U21429 ( .A(n20395), .Z(n20406) );
  XOR U21430 ( .A(n20407), .B(n20408), .Z(n20395) );
  AND U21431 ( .A(n20409), .B(n20410), .Z(n20408) );
  XNOR U21432 ( .A(n20407), .B(n10206), .Z(n20410) );
  XNOR U21433 ( .A(n20403), .B(n20405), .Z(n10206) );
  NAND U21434 ( .A(n20411), .B(e_input[349]), .Z(n20405) );
  NAND U21435 ( .A(n12323), .B(e_input[349]), .Z(n20411) );
  XNOR U21436 ( .A(n20401), .B(n20412), .Z(n20403) );
  XOR U21437 ( .A(n20413), .B(n20414), .Z(n20401) );
  AND U21438 ( .A(n20415), .B(n20416), .Z(n20414) );
  XNOR U21439 ( .A(n20417), .B(n20413), .Z(n20416) );
  XOR U21440 ( .A(n20418), .B(e_input[349]), .Z(n20409) );
  IV U21441 ( .A(n20407), .Z(n20418) );
  XOR U21442 ( .A(n20419), .B(n20420), .Z(n20407) );
  AND U21443 ( .A(n20421), .B(n20422), .Z(n20420) );
  XNOR U21444 ( .A(n20419), .B(n10212), .Z(n20422) );
  XNOR U21445 ( .A(n20415), .B(n20417), .Z(n10212) );
  NAND U21446 ( .A(n20423), .B(e_input[348]), .Z(n20417) );
  NAND U21447 ( .A(n12323), .B(e_input[348]), .Z(n20423) );
  XNOR U21448 ( .A(n20413), .B(n20424), .Z(n20415) );
  XOR U21449 ( .A(n20425), .B(n20426), .Z(n20413) );
  AND U21450 ( .A(n20427), .B(n20428), .Z(n20426) );
  XNOR U21451 ( .A(n20429), .B(n20425), .Z(n20428) );
  XOR U21452 ( .A(n20430), .B(e_input[348]), .Z(n20421) );
  IV U21453 ( .A(n20419), .Z(n20430) );
  XOR U21454 ( .A(n20431), .B(n20432), .Z(n20419) );
  AND U21455 ( .A(n20433), .B(n20434), .Z(n20432) );
  XNOR U21456 ( .A(n20431), .B(n10218), .Z(n20434) );
  XNOR U21457 ( .A(n20427), .B(n20429), .Z(n10218) );
  NAND U21458 ( .A(n20435), .B(e_input[347]), .Z(n20429) );
  NAND U21459 ( .A(n12323), .B(e_input[347]), .Z(n20435) );
  XNOR U21460 ( .A(n20425), .B(n20436), .Z(n20427) );
  XOR U21461 ( .A(n20437), .B(n20438), .Z(n20425) );
  AND U21462 ( .A(n20439), .B(n20440), .Z(n20438) );
  XNOR U21463 ( .A(n20441), .B(n20437), .Z(n20440) );
  XOR U21464 ( .A(n20442), .B(e_input[347]), .Z(n20433) );
  IV U21465 ( .A(n20431), .Z(n20442) );
  XOR U21466 ( .A(n20443), .B(n20444), .Z(n20431) );
  AND U21467 ( .A(n20445), .B(n20446), .Z(n20444) );
  XNOR U21468 ( .A(n20443), .B(n10224), .Z(n20446) );
  XNOR U21469 ( .A(n20439), .B(n20441), .Z(n10224) );
  NAND U21470 ( .A(n20447), .B(e_input[346]), .Z(n20441) );
  NAND U21471 ( .A(n12323), .B(e_input[346]), .Z(n20447) );
  XNOR U21472 ( .A(n20437), .B(n20448), .Z(n20439) );
  XOR U21473 ( .A(n20449), .B(n20450), .Z(n20437) );
  AND U21474 ( .A(n20451), .B(n20452), .Z(n20450) );
  XNOR U21475 ( .A(n20453), .B(n20449), .Z(n20452) );
  XOR U21476 ( .A(n20454), .B(e_input[346]), .Z(n20445) );
  IV U21477 ( .A(n20443), .Z(n20454) );
  XOR U21478 ( .A(n20455), .B(n20456), .Z(n20443) );
  AND U21479 ( .A(n20457), .B(n20458), .Z(n20456) );
  XNOR U21480 ( .A(n20455), .B(n10230), .Z(n20458) );
  XNOR U21481 ( .A(n20451), .B(n20453), .Z(n10230) );
  NAND U21482 ( .A(n20459), .B(e_input[345]), .Z(n20453) );
  NAND U21483 ( .A(n12323), .B(e_input[345]), .Z(n20459) );
  XNOR U21484 ( .A(n20449), .B(n20460), .Z(n20451) );
  XOR U21485 ( .A(n20461), .B(n20462), .Z(n20449) );
  AND U21486 ( .A(n20463), .B(n20464), .Z(n20462) );
  XNOR U21487 ( .A(n20465), .B(n20461), .Z(n20464) );
  XOR U21488 ( .A(n20466), .B(e_input[345]), .Z(n20457) );
  IV U21489 ( .A(n20455), .Z(n20466) );
  XOR U21490 ( .A(n20467), .B(n20468), .Z(n20455) );
  AND U21491 ( .A(n20469), .B(n20470), .Z(n20468) );
  XNOR U21492 ( .A(n20467), .B(n10236), .Z(n20470) );
  XNOR U21493 ( .A(n20463), .B(n20465), .Z(n10236) );
  NAND U21494 ( .A(n20471), .B(e_input[344]), .Z(n20465) );
  NAND U21495 ( .A(n12323), .B(e_input[344]), .Z(n20471) );
  XNOR U21496 ( .A(n20461), .B(n20472), .Z(n20463) );
  XOR U21497 ( .A(n20473), .B(n20474), .Z(n20461) );
  AND U21498 ( .A(n20475), .B(n20476), .Z(n20474) );
  XNOR U21499 ( .A(n20477), .B(n20473), .Z(n20476) );
  XOR U21500 ( .A(n20478), .B(e_input[344]), .Z(n20469) );
  IV U21501 ( .A(n20467), .Z(n20478) );
  XOR U21502 ( .A(n20479), .B(n20480), .Z(n20467) );
  AND U21503 ( .A(n20481), .B(n20482), .Z(n20480) );
  XNOR U21504 ( .A(n20479), .B(n10242), .Z(n20482) );
  XNOR U21505 ( .A(n20475), .B(n20477), .Z(n10242) );
  NAND U21506 ( .A(n20483), .B(e_input[343]), .Z(n20477) );
  NAND U21507 ( .A(n12323), .B(e_input[343]), .Z(n20483) );
  XNOR U21508 ( .A(n20473), .B(n20484), .Z(n20475) );
  XOR U21509 ( .A(n20485), .B(n20486), .Z(n20473) );
  AND U21510 ( .A(n20487), .B(n20488), .Z(n20486) );
  XNOR U21511 ( .A(n20489), .B(n20485), .Z(n20488) );
  XOR U21512 ( .A(n20490), .B(e_input[343]), .Z(n20481) );
  IV U21513 ( .A(n20479), .Z(n20490) );
  XOR U21514 ( .A(n20491), .B(n20492), .Z(n20479) );
  AND U21515 ( .A(n20493), .B(n20494), .Z(n20492) );
  XNOR U21516 ( .A(n20491), .B(n10248), .Z(n20494) );
  XNOR U21517 ( .A(n20487), .B(n20489), .Z(n10248) );
  NAND U21518 ( .A(n20495), .B(e_input[342]), .Z(n20489) );
  NAND U21519 ( .A(n12323), .B(e_input[342]), .Z(n20495) );
  XNOR U21520 ( .A(n20485), .B(n20496), .Z(n20487) );
  XOR U21521 ( .A(n20497), .B(n20498), .Z(n20485) );
  AND U21522 ( .A(n20499), .B(n20500), .Z(n20498) );
  XNOR U21523 ( .A(n20501), .B(n20497), .Z(n20500) );
  XOR U21524 ( .A(n20502), .B(e_input[342]), .Z(n20493) );
  IV U21525 ( .A(n20491), .Z(n20502) );
  XOR U21526 ( .A(n20503), .B(n20504), .Z(n20491) );
  AND U21527 ( .A(n20505), .B(n20506), .Z(n20504) );
  XNOR U21528 ( .A(n20503), .B(n10254), .Z(n20506) );
  XNOR U21529 ( .A(n20499), .B(n20501), .Z(n10254) );
  NAND U21530 ( .A(n20507), .B(e_input[341]), .Z(n20501) );
  NAND U21531 ( .A(n12323), .B(e_input[341]), .Z(n20507) );
  XNOR U21532 ( .A(n20497), .B(n20508), .Z(n20499) );
  XOR U21533 ( .A(n20509), .B(n20510), .Z(n20497) );
  AND U21534 ( .A(n20511), .B(n20512), .Z(n20510) );
  XNOR U21535 ( .A(n20513), .B(n20509), .Z(n20512) );
  XOR U21536 ( .A(n20514), .B(e_input[341]), .Z(n20505) );
  IV U21537 ( .A(n20503), .Z(n20514) );
  XOR U21538 ( .A(n20515), .B(n20516), .Z(n20503) );
  AND U21539 ( .A(n20517), .B(n20518), .Z(n20516) );
  XNOR U21540 ( .A(n20515), .B(n10260), .Z(n20518) );
  XNOR U21541 ( .A(n20511), .B(n20513), .Z(n10260) );
  NAND U21542 ( .A(n20519), .B(e_input[340]), .Z(n20513) );
  NAND U21543 ( .A(n12323), .B(e_input[340]), .Z(n20519) );
  XNOR U21544 ( .A(n20509), .B(n20520), .Z(n20511) );
  XOR U21545 ( .A(n20521), .B(n20522), .Z(n20509) );
  AND U21546 ( .A(n20523), .B(n20524), .Z(n20522) );
  XNOR U21547 ( .A(n20525), .B(n20521), .Z(n20524) );
  XOR U21548 ( .A(n20526), .B(e_input[340]), .Z(n20517) );
  IV U21549 ( .A(n20515), .Z(n20526) );
  XOR U21550 ( .A(n20527), .B(n20528), .Z(n20515) );
  AND U21551 ( .A(n20529), .B(n20530), .Z(n20528) );
  XNOR U21552 ( .A(n20527), .B(n10266), .Z(n20530) );
  XNOR U21553 ( .A(n20523), .B(n20525), .Z(n10266) );
  NAND U21554 ( .A(n20531), .B(e_input[339]), .Z(n20525) );
  NAND U21555 ( .A(n12323), .B(e_input[339]), .Z(n20531) );
  XNOR U21556 ( .A(n20521), .B(n20532), .Z(n20523) );
  XOR U21557 ( .A(n20533), .B(n20534), .Z(n20521) );
  AND U21558 ( .A(n20535), .B(n20536), .Z(n20534) );
  XNOR U21559 ( .A(n20537), .B(n20533), .Z(n20536) );
  XOR U21560 ( .A(n20538), .B(e_input[339]), .Z(n20529) );
  IV U21561 ( .A(n20527), .Z(n20538) );
  XOR U21562 ( .A(n20539), .B(n20540), .Z(n20527) );
  AND U21563 ( .A(n20541), .B(n20542), .Z(n20540) );
  XNOR U21564 ( .A(n20539), .B(n10272), .Z(n20542) );
  XNOR U21565 ( .A(n20535), .B(n20537), .Z(n10272) );
  NAND U21566 ( .A(n20543), .B(e_input[338]), .Z(n20537) );
  NAND U21567 ( .A(n12323), .B(e_input[338]), .Z(n20543) );
  XNOR U21568 ( .A(n20533), .B(n20544), .Z(n20535) );
  XOR U21569 ( .A(n20545), .B(n20546), .Z(n20533) );
  AND U21570 ( .A(n20547), .B(n20548), .Z(n20546) );
  XNOR U21571 ( .A(n20549), .B(n20545), .Z(n20548) );
  XOR U21572 ( .A(n20550), .B(e_input[338]), .Z(n20541) );
  IV U21573 ( .A(n20539), .Z(n20550) );
  XOR U21574 ( .A(n20551), .B(n20552), .Z(n20539) );
  AND U21575 ( .A(n20553), .B(n20554), .Z(n20552) );
  XNOR U21576 ( .A(n20551), .B(n10278), .Z(n20554) );
  XNOR U21577 ( .A(n20547), .B(n20549), .Z(n10278) );
  NAND U21578 ( .A(n20555), .B(e_input[337]), .Z(n20549) );
  NAND U21579 ( .A(n12323), .B(e_input[337]), .Z(n20555) );
  XNOR U21580 ( .A(n20545), .B(n20556), .Z(n20547) );
  XOR U21581 ( .A(n20557), .B(n20558), .Z(n20545) );
  AND U21582 ( .A(n20559), .B(n20560), .Z(n20558) );
  XNOR U21583 ( .A(n20561), .B(n20557), .Z(n20560) );
  XOR U21584 ( .A(n20562), .B(e_input[337]), .Z(n20553) );
  IV U21585 ( .A(n20551), .Z(n20562) );
  XOR U21586 ( .A(n20563), .B(n20564), .Z(n20551) );
  AND U21587 ( .A(n20565), .B(n20566), .Z(n20564) );
  XNOR U21588 ( .A(n20563), .B(n10284), .Z(n20566) );
  XNOR U21589 ( .A(n20559), .B(n20561), .Z(n10284) );
  NAND U21590 ( .A(n20567), .B(e_input[336]), .Z(n20561) );
  NAND U21591 ( .A(n12323), .B(e_input[336]), .Z(n20567) );
  XNOR U21592 ( .A(n20557), .B(n20568), .Z(n20559) );
  XOR U21593 ( .A(n20569), .B(n20570), .Z(n20557) );
  AND U21594 ( .A(n20571), .B(n20572), .Z(n20570) );
  XNOR U21595 ( .A(n20573), .B(n20569), .Z(n20572) );
  XOR U21596 ( .A(n20574), .B(e_input[336]), .Z(n20565) );
  IV U21597 ( .A(n20563), .Z(n20574) );
  XOR U21598 ( .A(n20575), .B(n20576), .Z(n20563) );
  AND U21599 ( .A(n20577), .B(n20578), .Z(n20576) );
  XNOR U21600 ( .A(n20575), .B(n10290), .Z(n20578) );
  XNOR U21601 ( .A(n20571), .B(n20573), .Z(n10290) );
  NAND U21602 ( .A(n20579), .B(e_input[335]), .Z(n20573) );
  NAND U21603 ( .A(n12323), .B(e_input[335]), .Z(n20579) );
  XNOR U21604 ( .A(n20569), .B(n20580), .Z(n20571) );
  XOR U21605 ( .A(n20581), .B(n20582), .Z(n20569) );
  AND U21606 ( .A(n20583), .B(n20584), .Z(n20582) );
  XNOR U21607 ( .A(n20585), .B(n20581), .Z(n20584) );
  XOR U21608 ( .A(n20586), .B(e_input[335]), .Z(n20577) );
  IV U21609 ( .A(n20575), .Z(n20586) );
  XOR U21610 ( .A(n20587), .B(n20588), .Z(n20575) );
  AND U21611 ( .A(n20589), .B(n20590), .Z(n20588) );
  XNOR U21612 ( .A(n20587), .B(n10296), .Z(n20590) );
  XNOR U21613 ( .A(n20583), .B(n20585), .Z(n10296) );
  NAND U21614 ( .A(n20591), .B(e_input[334]), .Z(n20585) );
  NAND U21615 ( .A(n12323), .B(e_input[334]), .Z(n20591) );
  XNOR U21616 ( .A(n20581), .B(n20592), .Z(n20583) );
  XOR U21617 ( .A(n20593), .B(n20594), .Z(n20581) );
  AND U21618 ( .A(n20595), .B(n20596), .Z(n20594) );
  XNOR U21619 ( .A(n20597), .B(n20593), .Z(n20596) );
  XOR U21620 ( .A(n20598), .B(e_input[334]), .Z(n20589) );
  IV U21621 ( .A(n20587), .Z(n20598) );
  XOR U21622 ( .A(n20599), .B(n20600), .Z(n20587) );
  AND U21623 ( .A(n20601), .B(n20602), .Z(n20600) );
  XNOR U21624 ( .A(n20599), .B(n10302), .Z(n20602) );
  XNOR U21625 ( .A(n20595), .B(n20597), .Z(n10302) );
  NAND U21626 ( .A(n20603), .B(e_input[333]), .Z(n20597) );
  NAND U21627 ( .A(n12323), .B(e_input[333]), .Z(n20603) );
  XNOR U21628 ( .A(n20593), .B(n20604), .Z(n20595) );
  XOR U21629 ( .A(n20605), .B(n20606), .Z(n20593) );
  AND U21630 ( .A(n20607), .B(n20608), .Z(n20606) );
  XNOR U21631 ( .A(n20609), .B(n20605), .Z(n20608) );
  XOR U21632 ( .A(n20610), .B(e_input[333]), .Z(n20601) );
  IV U21633 ( .A(n20599), .Z(n20610) );
  XOR U21634 ( .A(n20611), .B(n20612), .Z(n20599) );
  AND U21635 ( .A(n20613), .B(n20614), .Z(n20612) );
  XNOR U21636 ( .A(n20611), .B(n10308), .Z(n20614) );
  XNOR U21637 ( .A(n20607), .B(n20609), .Z(n10308) );
  NAND U21638 ( .A(n20615), .B(e_input[332]), .Z(n20609) );
  NAND U21639 ( .A(n12323), .B(e_input[332]), .Z(n20615) );
  XNOR U21640 ( .A(n20605), .B(n20616), .Z(n20607) );
  XOR U21641 ( .A(n20617), .B(n20618), .Z(n20605) );
  AND U21642 ( .A(n20619), .B(n20620), .Z(n20618) );
  XNOR U21643 ( .A(n20621), .B(n20617), .Z(n20620) );
  XOR U21644 ( .A(n20622), .B(e_input[332]), .Z(n20613) );
  IV U21645 ( .A(n20611), .Z(n20622) );
  XOR U21646 ( .A(n20623), .B(n20624), .Z(n20611) );
  AND U21647 ( .A(n20625), .B(n20626), .Z(n20624) );
  XNOR U21648 ( .A(n20623), .B(n10314), .Z(n20626) );
  XNOR U21649 ( .A(n20619), .B(n20621), .Z(n10314) );
  NAND U21650 ( .A(n20627), .B(e_input[331]), .Z(n20621) );
  NAND U21651 ( .A(n12323), .B(e_input[331]), .Z(n20627) );
  XNOR U21652 ( .A(n20617), .B(n20628), .Z(n20619) );
  XOR U21653 ( .A(n20629), .B(n20630), .Z(n20617) );
  AND U21654 ( .A(n20631), .B(n20632), .Z(n20630) );
  XNOR U21655 ( .A(n20633), .B(n20629), .Z(n20632) );
  XOR U21656 ( .A(n20634), .B(e_input[331]), .Z(n20625) );
  IV U21657 ( .A(n20623), .Z(n20634) );
  XOR U21658 ( .A(n20635), .B(n20636), .Z(n20623) );
  AND U21659 ( .A(n20637), .B(n20638), .Z(n20636) );
  XNOR U21660 ( .A(n20635), .B(n10320), .Z(n20638) );
  XNOR U21661 ( .A(n20631), .B(n20633), .Z(n10320) );
  NAND U21662 ( .A(n20639), .B(e_input[330]), .Z(n20633) );
  NAND U21663 ( .A(n12323), .B(e_input[330]), .Z(n20639) );
  XNOR U21664 ( .A(n20629), .B(n20640), .Z(n20631) );
  XOR U21665 ( .A(n20641), .B(n20642), .Z(n20629) );
  AND U21666 ( .A(n20643), .B(n20644), .Z(n20642) );
  XNOR U21667 ( .A(n20645), .B(n20641), .Z(n20644) );
  XOR U21668 ( .A(n20646), .B(e_input[330]), .Z(n20637) );
  IV U21669 ( .A(n20635), .Z(n20646) );
  XOR U21670 ( .A(n20647), .B(n20648), .Z(n20635) );
  AND U21671 ( .A(n20649), .B(n20650), .Z(n20648) );
  XNOR U21672 ( .A(n20647), .B(n10326), .Z(n20650) );
  XNOR U21673 ( .A(n20643), .B(n20645), .Z(n10326) );
  NAND U21674 ( .A(n20651), .B(e_input[329]), .Z(n20645) );
  NAND U21675 ( .A(n12323), .B(e_input[329]), .Z(n20651) );
  XNOR U21676 ( .A(n20641), .B(n20652), .Z(n20643) );
  XOR U21677 ( .A(n20653), .B(n20654), .Z(n20641) );
  AND U21678 ( .A(n20655), .B(n20656), .Z(n20654) );
  XNOR U21679 ( .A(n20657), .B(n20653), .Z(n20656) );
  XOR U21680 ( .A(n20658), .B(e_input[329]), .Z(n20649) );
  IV U21681 ( .A(n20647), .Z(n20658) );
  XOR U21682 ( .A(n20659), .B(n20660), .Z(n20647) );
  AND U21683 ( .A(n20661), .B(n20662), .Z(n20660) );
  XNOR U21684 ( .A(n20659), .B(n10332), .Z(n20662) );
  XNOR U21685 ( .A(n20655), .B(n20657), .Z(n10332) );
  NAND U21686 ( .A(n20663), .B(e_input[328]), .Z(n20657) );
  NAND U21687 ( .A(n12323), .B(e_input[328]), .Z(n20663) );
  XNOR U21688 ( .A(n20653), .B(n20664), .Z(n20655) );
  XOR U21689 ( .A(n20665), .B(n20666), .Z(n20653) );
  AND U21690 ( .A(n20667), .B(n20668), .Z(n20666) );
  XNOR U21691 ( .A(n20669), .B(n20665), .Z(n20668) );
  XOR U21692 ( .A(n20670), .B(e_input[328]), .Z(n20661) );
  IV U21693 ( .A(n20659), .Z(n20670) );
  XOR U21694 ( .A(n20671), .B(n20672), .Z(n20659) );
  AND U21695 ( .A(n20673), .B(n20674), .Z(n20672) );
  XNOR U21696 ( .A(n20671), .B(n10338), .Z(n20674) );
  XNOR U21697 ( .A(n20667), .B(n20669), .Z(n10338) );
  NAND U21698 ( .A(n20675), .B(e_input[327]), .Z(n20669) );
  NAND U21699 ( .A(n12323), .B(e_input[327]), .Z(n20675) );
  XNOR U21700 ( .A(n20665), .B(n20676), .Z(n20667) );
  XOR U21701 ( .A(n20677), .B(n20678), .Z(n20665) );
  AND U21702 ( .A(n20679), .B(n20680), .Z(n20678) );
  XNOR U21703 ( .A(n20681), .B(n20677), .Z(n20680) );
  XOR U21704 ( .A(n20682), .B(e_input[327]), .Z(n20673) );
  IV U21705 ( .A(n20671), .Z(n20682) );
  XOR U21706 ( .A(n20683), .B(n20684), .Z(n20671) );
  AND U21707 ( .A(n20685), .B(n20686), .Z(n20684) );
  XNOR U21708 ( .A(n20683), .B(n10344), .Z(n20686) );
  XNOR U21709 ( .A(n20679), .B(n20681), .Z(n10344) );
  NAND U21710 ( .A(n20687), .B(e_input[326]), .Z(n20681) );
  NAND U21711 ( .A(n12323), .B(e_input[326]), .Z(n20687) );
  XNOR U21712 ( .A(n20677), .B(n20688), .Z(n20679) );
  XOR U21713 ( .A(n20689), .B(n20690), .Z(n20677) );
  AND U21714 ( .A(n20691), .B(n20692), .Z(n20690) );
  XNOR U21715 ( .A(n20693), .B(n20689), .Z(n20692) );
  XOR U21716 ( .A(n20694), .B(e_input[326]), .Z(n20685) );
  IV U21717 ( .A(n20683), .Z(n20694) );
  XOR U21718 ( .A(n20695), .B(n20696), .Z(n20683) );
  AND U21719 ( .A(n20697), .B(n20698), .Z(n20696) );
  XNOR U21720 ( .A(n20695), .B(n10350), .Z(n20698) );
  XNOR U21721 ( .A(n20691), .B(n20693), .Z(n10350) );
  NAND U21722 ( .A(n20699), .B(e_input[325]), .Z(n20693) );
  NAND U21723 ( .A(n12323), .B(e_input[325]), .Z(n20699) );
  XNOR U21724 ( .A(n20689), .B(n20700), .Z(n20691) );
  XOR U21725 ( .A(n20701), .B(n20702), .Z(n20689) );
  AND U21726 ( .A(n20703), .B(n20704), .Z(n20702) );
  XNOR U21727 ( .A(n20705), .B(n20701), .Z(n20704) );
  XOR U21728 ( .A(n20706), .B(e_input[325]), .Z(n20697) );
  IV U21729 ( .A(n20695), .Z(n20706) );
  XOR U21730 ( .A(n20707), .B(n20708), .Z(n20695) );
  AND U21731 ( .A(n20709), .B(n20710), .Z(n20708) );
  XNOR U21732 ( .A(n20707), .B(n10356), .Z(n20710) );
  XNOR U21733 ( .A(n20703), .B(n20705), .Z(n10356) );
  NAND U21734 ( .A(n20711), .B(e_input[324]), .Z(n20705) );
  NAND U21735 ( .A(n12323), .B(e_input[324]), .Z(n20711) );
  XNOR U21736 ( .A(n20701), .B(n20712), .Z(n20703) );
  XOR U21737 ( .A(n20713), .B(n20714), .Z(n20701) );
  AND U21738 ( .A(n20715), .B(n20716), .Z(n20714) );
  XNOR U21739 ( .A(n20717), .B(n20713), .Z(n20716) );
  XOR U21740 ( .A(n20718), .B(e_input[324]), .Z(n20709) );
  IV U21741 ( .A(n20707), .Z(n20718) );
  XOR U21742 ( .A(n20719), .B(n20720), .Z(n20707) );
  AND U21743 ( .A(n20721), .B(n20722), .Z(n20720) );
  XNOR U21744 ( .A(n20719), .B(n10362), .Z(n20722) );
  XNOR U21745 ( .A(n20715), .B(n20717), .Z(n10362) );
  NAND U21746 ( .A(n20723), .B(e_input[323]), .Z(n20717) );
  NAND U21747 ( .A(n12323), .B(e_input[323]), .Z(n20723) );
  XNOR U21748 ( .A(n20713), .B(n20724), .Z(n20715) );
  XOR U21749 ( .A(n20725), .B(n20726), .Z(n20713) );
  AND U21750 ( .A(n20727), .B(n20728), .Z(n20726) );
  XNOR U21751 ( .A(n20729), .B(n20725), .Z(n20728) );
  XOR U21752 ( .A(n20730), .B(e_input[323]), .Z(n20721) );
  IV U21753 ( .A(n20719), .Z(n20730) );
  XOR U21754 ( .A(n20731), .B(n20732), .Z(n20719) );
  AND U21755 ( .A(n20733), .B(n20734), .Z(n20732) );
  XNOR U21756 ( .A(n20731), .B(n10368), .Z(n20734) );
  XNOR U21757 ( .A(n20727), .B(n20729), .Z(n10368) );
  NAND U21758 ( .A(n20735), .B(e_input[322]), .Z(n20729) );
  NAND U21759 ( .A(n12323), .B(e_input[322]), .Z(n20735) );
  XNOR U21760 ( .A(n20725), .B(n20736), .Z(n20727) );
  XOR U21761 ( .A(n20737), .B(n20738), .Z(n20725) );
  AND U21762 ( .A(n20739), .B(n20740), .Z(n20738) );
  XNOR U21763 ( .A(n20741), .B(n20737), .Z(n20740) );
  XOR U21764 ( .A(n20742), .B(e_input[322]), .Z(n20733) );
  IV U21765 ( .A(n20731), .Z(n20742) );
  XOR U21766 ( .A(n20743), .B(n20744), .Z(n20731) );
  AND U21767 ( .A(n20745), .B(n20746), .Z(n20744) );
  XNOR U21768 ( .A(n20743), .B(n10374), .Z(n20746) );
  XNOR U21769 ( .A(n20739), .B(n20741), .Z(n10374) );
  NAND U21770 ( .A(n20747), .B(e_input[321]), .Z(n20741) );
  NAND U21771 ( .A(n12323), .B(e_input[321]), .Z(n20747) );
  XNOR U21772 ( .A(n20737), .B(n20748), .Z(n20739) );
  XOR U21773 ( .A(n20749), .B(n20750), .Z(n20737) );
  AND U21774 ( .A(n20751), .B(n20752), .Z(n20750) );
  XNOR U21775 ( .A(n20753), .B(n20749), .Z(n20752) );
  XOR U21776 ( .A(n20754), .B(e_input[321]), .Z(n20745) );
  IV U21777 ( .A(n20743), .Z(n20754) );
  XOR U21778 ( .A(n20755), .B(n20756), .Z(n20743) );
  AND U21779 ( .A(n20757), .B(n20758), .Z(n20756) );
  XNOR U21780 ( .A(n20755), .B(n10380), .Z(n20758) );
  XNOR U21781 ( .A(n20751), .B(n20753), .Z(n10380) );
  NAND U21782 ( .A(n20759), .B(e_input[320]), .Z(n20753) );
  NAND U21783 ( .A(n12323), .B(e_input[320]), .Z(n20759) );
  XNOR U21784 ( .A(n20749), .B(n20760), .Z(n20751) );
  XOR U21785 ( .A(n20761), .B(n20762), .Z(n20749) );
  AND U21786 ( .A(n20763), .B(n20764), .Z(n20762) );
  XNOR U21787 ( .A(n20765), .B(n20761), .Z(n20764) );
  XOR U21788 ( .A(n20766), .B(e_input[320]), .Z(n20757) );
  IV U21789 ( .A(n20755), .Z(n20766) );
  XOR U21790 ( .A(n20767), .B(n20768), .Z(n20755) );
  AND U21791 ( .A(n20769), .B(n20770), .Z(n20768) );
  XNOR U21792 ( .A(n20767), .B(n10386), .Z(n20770) );
  XNOR U21793 ( .A(n20763), .B(n20765), .Z(n10386) );
  NAND U21794 ( .A(n20771), .B(e_input[319]), .Z(n20765) );
  NAND U21795 ( .A(n12323), .B(e_input[319]), .Z(n20771) );
  XNOR U21796 ( .A(n20761), .B(n20772), .Z(n20763) );
  XOR U21797 ( .A(n20773), .B(n20774), .Z(n20761) );
  AND U21798 ( .A(n20775), .B(n20776), .Z(n20774) );
  XNOR U21799 ( .A(n20777), .B(n20773), .Z(n20776) );
  XOR U21800 ( .A(n20778), .B(e_input[319]), .Z(n20769) );
  IV U21801 ( .A(n20767), .Z(n20778) );
  XOR U21802 ( .A(n20779), .B(n20780), .Z(n20767) );
  AND U21803 ( .A(n20781), .B(n20782), .Z(n20780) );
  XNOR U21804 ( .A(n20779), .B(n10392), .Z(n20782) );
  XNOR U21805 ( .A(n20775), .B(n20777), .Z(n10392) );
  NAND U21806 ( .A(n20783), .B(e_input[318]), .Z(n20777) );
  NAND U21807 ( .A(n12323), .B(e_input[318]), .Z(n20783) );
  XNOR U21808 ( .A(n20773), .B(n20784), .Z(n20775) );
  XOR U21809 ( .A(n20785), .B(n20786), .Z(n20773) );
  AND U21810 ( .A(n20787), .B(n20788), .Z(n20786) );
  XNOR U21811 ( .A(n20789), .B(n20785), .Z(n20788) );
  XOR U21812 ( .A(n20790), .B(e_input[318]), .Z(n20781) );
  IV U21813 ( .A(n20779), .Z(n20790) );
  XOR U21814 ( .A(n20791), .B(n20792), .Z(n20779) );
  AND U21815 ( .A(n20793), .B(n20794), .Z(n20792) );
  XNOR U21816 ( .A(n20791), .B(n10398), .Z(n20794) );
  XNOR U21817 ( .A(n20787), .B(n20789), .Z(n10398) );
  NAND U21818 ( .A(n20795), .B(e_input[317]), .Z(n20789) );
  NAND U21819 ( .A(n12323), .B(e_input[317]), .Z(n20795) );
  XNOR U21820 ( .A(n20785), .B(n20796), .Z(n20787) );
  XOR U21821 ( .A(n20797), .B(n20798), .Z(n20785) );
  AND U21822 ( .A(n20799), .B(n20800), .Z(n20798) );
  XNOR U21823 ( .A(n20801), .B(n20797), .Z(n20800) );
  XOR U21824 ( .A(n20802), .B(e_input[317]), .Z(n20793) );
  IV U21825 ( .A(n20791), .Z(n20802) );
  XOR U21826 ( .A(n20803), .B(n20804), .Z(n20791) );
  AND U21827 ( .A(n20805), .B(n20806), .Z(n20804) );
  XNOR U21828 ( .A(n20803), .B(n10404), .Z(n20806) );
  XNOR U21829 ( .A(n20799), .B(n20801), .Z(n10404) );
  NAND U21830 ( .A(n20807), .B(e_input[316]), .Z(n20801) );
  NAND U21831 ( .A(n12323), .B(e_input[316]), .Z(n20807) );
  XNOR U21832 ( .A(n20797), .B(n20808), .Z(n20799) );
  XOR U21833 ( .A(n20809), .B(n20810), .Z(n20797) );
  AND U21834 ( .A(n20811), .B(n20812), .Z(n20810) );
  XNOR U21835 ( .A(n20813), .B(n20809), .Z(n20812) );
  XOR U21836 ( .A(n20814), .B(e_input[316]), .Z(n20805) );
  IV U21837 ( .A(n20803), .Z(n20814) );
  XOR U21838 ( .A(n20815), .B(n20816), .Z(n20803) );
  AND U21839 ( .A(n20817), .B(n20818), .Z(n20816) );
  XNOR U21840 ( .A(n20815), .B(n10410), .Z(n20818) );
  XNOR U21841 ( .A(n20811), .B(n20813), .Z(n10410) );
  NAND U21842 ( .A(n20819), .B(e_input[315]), .Z(n20813) );
  NAND U21843 ( .A(n12323), .B(e_input[315]), .Z(n20819) );
  XNOR U21844 ( .A(n20809), .B(n20820), .Z(n20811) );
  XOR U21845 ( .A(n20821), .B(n20822), .Z(n20809) );
  AND U21846 ( .A(n20823), .B(n20824), .Z(n20822) );
  XNOR U21847 ( .A(n20825), .B(n20821), .Z(n20824) );
  XOR U21848 ( .A(n20826), .B(e_input[315]), .Z(n20817) );
  IV U21849 ( .A(n20815), .Z(n20826) );
  XOR U21850 ( .A(n20827), .B(n20828), .Z(n20815) );
  AND U21851 ( .A(n20829), .B(n20830), .Z(n20828) );
  XNOR U21852 ( .A(n20827), .B(n10416), .Z(n20830) );
  XNOR U21853 ( .A(n20823), .B(n20825), .Z(n10416) );
  NAND U21854 ( .A(n20831), .B(e_input[314]), .Z(n20825) );
  NAND U21855 ( .A(n12323), .B(e_input[314]), .Z(n20831) );
  XNOR U21856 ( .A(n20821), .B(n20832), .Z(n20823) );
  XOR U21857 ( .A(n20833), .B(n20834), .Z(n20821) );
  AND U21858 ( .A(n20835), .B(n20836), .Z(n20834) );
  XNOR U21859 ( .A(n20837), .B(n20833), .Z(n20836) );
  XOR U21860 ( .A(n20838), .B(e_input[314]), .Z(n20829) );
  IV U21861 ( .A(n20827), .Z(n20838) );
  XOR U21862 ( .A(n20839), .B(n20840), .Z(n20827) );
  AND U21863 ( .A(n20841), .B(n20842), .Z(n20840) );
  XNOR U21864 ( .A(n20839), .B(n10422), .Z(n20842) );
  XNOR U21865 ( .A(n20835), .B(n20837), .Z(n10422) );
  NAND U21866 ( .A(n20843), .B(e_input[313]), .Z(n20837) );
  NAND U21867 ( .A(n12323), .B(e_input[313]), .Z(n20843) );
  XNOR U21868 ( .A(n20833), .B(n20844), .Z(n20835) );
  XOR U21869 ( .A(n20845), .B(n20846), .Z(n20833) );
  AND U21870 ( .A(n20847), .B(n20848), .Z(n20846) );
  XNOR U21871 ( .A(n20849), .B(n20845), .Z(n20848) );
  XOR U21872 ( .A(n20850), .B(e_input[313]), .Z(n20841) );
  IV U21873 ( .A(n20839), .Z(n20850) );
  XOR U21874 ( .A(n20851), .B(n20852), .Z(n20839) );
  AND U21875 ( .A(n20853), .B(n20854), .Z(n20852) );
  XNOR U21876 ( .A(n20851), .B(n10428), .Z(n20854) );
  XNOR U21877 ( .A(n20847), .B(n20849), .Z(n10428) );
  NAND U21878 ( .A(n20855), .B(e_input[312]), .Z(n20849) );
  NAND U21879 ( .A(n12323), .B(e_input[312]), .Z(n20855) );
  XNOR U21880 ( .A(n20845), .B(n20856), .Z(n20847) );
  XOR U21881 ( .A(n20857), .B(n20858), .Z(n20845) );
  AND U21882 ( .A(n20859), .B(n20860), .Z(n20858) );
  XNOR U21883 ( .A(n20861), .B(n20857), .Z(n20860) );
  XOR U21884 ( .A(n20862), .B(e_input[312]), .Z(n20853) );
  IV U21885 ( .A(n20851), .Z(n20862) );
  XOR U21886 ( .A(n20863), .B(n20864), .Z(n20851) );
  AND U21887 ( .A(n20865), .B(n20866), .Z(n20864) );
  XNOR U21888 ( .A(n20863), .B(n10434), .Z(n20866) );
  XNOR U21889 ( .A(n20859), .B(n20861), .Z(n10434) );
  NAND U21890 ( .A(n20867), .B(e_input[311]), .Z(n20861) );
  NAND U21891 ( .A(n12323), .B(e_input[311]), .Z(n20867) );
  XNOR U21892 ( .A(n20857), .B(n20868), .Z(n20859) );
  XOR U21893 ( .A(n20869), .B(n20870), .Z(n20857) );
  AND U21894 ( .A(n20871), .B(n20872), .Z(n20870) );
  XNOR U21895 ( .A(n20873), .B(n20869), .Z(n20872) );
  XOR U21896 ( .A(n20874), .B(e_input[311]), .Z(n20865) );
  IV U21897 ( .A(n20863), .Z(n20874) );
  XOR U21898 ( .A(n20875), .B(n20876), .Z(n20863) );
  AND U21899 ( .A(n20877), .B(n20878), .Z(n20876) );
  XNOR U21900 ( .A(n20875), .B(n10440), .Z(n20878) );
  XNOR U21901 ( .A(n20871), .B(n20873), .Z(n10440) );
  NAND U21902 ( .A(n20879), .B(e_input[310]), .Z(n20873) );
  NAND U21903 ( .A(n12323), .B(e_input[310]), .Z(n20879) );
  XNOR U21904 ( .A(n20869), .B(n20880), .Z(n20871) );
  XOR U21905 ( .A(n20881), .B(n20882), .Z(n20869) );
  AND U21906 ( .A(n20883), .B(n20884), .Z(n20882) );
  XNOR U21907 ( .A(n20885), .B(n20881), .Z(n20884) );
  XOR U21908 ( .A(n20886), .B(e_input[310]), .Z(n20877) );
  IV U21909 ( .A(n20875), .Z(n20886) );
  XOR U21910 ( .A(n20887), .B(n20888), .Z(n20875) );
  AND U21911 ( .A(n20889), .B(n20890), .Z(n20888) );
  XNOR U21912 ( .A(n20887), .B(n10446), .Z(n20890) );
  XNOR U21913 ( .A(n20883), .B(n20885), .Z(n10446) );
  NAND U21914 ( .A(n20891), .B(e_input[309]), .Z(n20885) );
  NAND U21915 ( .A(n12323), .B(e_input[309]), .Z(n20891) );
  XNOR U21916 ( .A(n20881), .B(n20892), .Z(n20883) );
  XOR U21917 ( .A(n20893), .B(n20894), .Z(n20881) );
  AND U21918 ( .A(n20895), .B(n20896), .Z(n20894) );
  XNOR U21919 ( .A(n20897), .B(n20893), .Z(n20896) );
  XOR U21920 ( .A(n20898), .B(e_input[309]), .Z(n20889) );
  IV U21921 ( .A(n20887), .Z(n20898) );
  XOR U21922 ( .A(n20899), .B(n20900), .Z(n20887) );
  AND U21923 ( .A(n20901), .B(n20902), .Z(n20900) );
  XNOR U21924 ( .A(n20899), .B(n10452), .Z(n20902) );
  XNOR U21925 ( .A(n20895), .B(n20897), .Z(n10452) );
  NAND U21926 ( .A(n20903), .B(e_input[308]), .Z(n20897) );
  NAND U21927 ( .A(n12323), .B(e_input[308]), .Z(n20903) );
  XNOR U21928 ( .A(n20893), .B(n20904), .Z(n20895) );
  XOR U21929 ( .A(n20905), .B(n20906), .Z(n20893) );
  AND U21930 ( .A(n20907), .B(n20908), .Z(n20906) );
  XNOR U21931 ( .A(n20909), .B(n20905), .Z(n20908) );
  XOR U21932 ( .A(n20910), .B(e_input[308]), .Z(n20901) );
  IV U21933 ( .A(n20899), .Z(n20910) );
  XOR U21934 ( .A(n20911), .B(n20912), .Z(n20899) );
  AND U21935 ( .A(n20913), .B(n20914), .Z(n20912) );
  XNOR U21936 ( .A(n20911), .B(n10458), .Z(n20914) );
  XNOR U21937 ( .A(n20907), .B(n20909), .Z(n10458) );
  NAND U21938 ( .A(n20915), .B(e_input[307]), .Z(n20909) );
  NAND U21939 ( .A(n12323), .B(e_input[307]), .Z(n20915) );
  XNOR U21940 ( .A(n20905), .B(n20916), .Z(n20907) );
  XOR U21941 ( .A(n20917), .B(n20918), .Z(n20905) );
  AND U21942 ( .A(n20919), .B(n20920), .Z(n20918) );
  XNOR U21943 ( .A(n20921), .B(n20917), .Z(n20920) );
  XOR U21944 ( .A(n20922), .B(e_input[307]), .Z(n20913) );
  IV U21945 ( .A(n20911), .Z(n20922) );
  XOR U21946 ( .A(n20923), .B(n20924), .Z(n20911) );
  AND U21947 ( .A(n20925), .B(n20926), .Z(n20924) );
  XNOR U21948 ( .A(n20923), .B(n10464), .Z(n20926) );
  XNOR U21949 ( .A(n20919), .B(n20921), .Z(n10464) );
  NAND U21950 ( .A(n20927), .B(e_input[306]), .Z(n20921) );
  NAND U21951 ( .A(n12323), .B(e_input[306]), .Z(n20927) );
  XNOR U21952 ( .A(n20917), .B(n20928), .Z(n20919) );
  XOR U21953 ( .A(n20929), .B(n20930), .Z(n20917) );
  AND U21954 ( .A(n20931), .B(n20932), .Z(n20930) );
  XNOR U21955 ( .A(n20933), .B(n20929), .Z(n20932) );
  XOR U21956 ( .A(n20934), .B(e_input[306]), .Z(n20925) );
  IV U21957 ( .A(n20923), .Z(n20934) );
  XOR U21958 ( .A(n20935), .B(n20936), .Z(n20923) );
  AND U21959 ( .A(n20937), .B(n20938), .Z(n20936) );
  XNOR U21960 ( .A(n20935), .B(n10470), .Z(n20938) );
  XNOR U21961 ( .A(n20931), .B(n20933), .Z(n10470) );
  NAND U21962 ( .A(n20939), .B(e_input[305]), .Z(n20933) );
  NAND U21963 ( .A(n12323), .B(e_input[305]), .Z(n20939) );
  XNOR U21964 ( .A(n20929), .B(n20940), .Z(n20931) );
  XOR U21965 ( .A(n20941), .B(n20942), .Z(n20929) );
  AND U21966 ( .A(n20943), .B(n20944), .Z(n20942) );
  XNOR U21967 ( .A(n20945), .B(n20941), .Z(n20944) );
  XOR U21968 ( .A(n20946), .B(e_input[305]), .Z(n20937) );
  IV U21969 ( .A(n20935), .Z(n20946) );
  XOR U21970 ( .A(n20947), .B(n20948), .Z(n20935) );
  AND U21971 ( .A(n20949), .B(n20950), .Z(n20948) );
  XNOR U21972 ( .A(n20947), .B(n10476), .Z(n20950) );
  XNOR U21973 ( .A(n20943), .B(n20945), .Z(n10476) );
  NAND U21974 ( .A(n20951), .B(e_input[304]), .Z(n20945) );
  NAND U21975 ( .A(n12323), .B(e_input[304]), .Z(n20951) );
  XNOR U21976 ( .A(n20941), .B(n20952), .Z(n20943) );
  XOR U21977 ( .A(n20953), .B(n20954), .Z(n20941) );
  AND U21978 ( .A(n20955), .B(n20956), .Z(n20954) );
  XNOR U21979 ( .A(n20957), .B(n20953), .Z(n20956) );
  XOR U21980 ( .A(n20958), .B(e_input[304]), .Z(n20949) );
  IV U21981 ( .A(n20947), .Z(n20958) );
  XOR U21982 ( .A(n20959), .B(n20960), .Z(n20947) );
  AND U21983 ( .A(n20961), .B(n20962), .Z(n20960) );
  XNOR U21984 ( .A(n20959), .B(n10482), .Z(n20962) );
  XNOR U21985 ( .A(n20955), .B(n20957), .Z(n10482) );
  NAND U21986 ( .A(n20963), .B(e_input[303]), .Z(n20957) );
  NAND U21987 ( .A(n12323), .B(e_input[303]), .Z(n20963) );
  XNOR U21988 ( .A(n20953), .B(n20964), .Z(n20955) );
  XOR U21989 ( .A(n20965), .B(n20966), .Z(n20953) );
  AND U21990 ( .A(n20967), .B(n20968), .Z(n20966) );
  XNOR U21991 ( .A(n20969), .B(n20965), .Z(n20968) );
  XOR U21992 ( .A(n20970), .B(e_input[303]), .Z(n20961) );
  IV U21993 ( .A(n20959), .Z(n20970) );
  XOR U21994 ( .A(n20971), .B(n20972), .Z(n20959) );
  AND U21995 ( .A(n20973), .B(n20974), .Z(n20972) );
  XNOR U21996 ( .A(n20971), .B(n10488), .Z(n20974) );
  XNOR U21997 ( .A(n20967), .B(n20969), .Z(n10488) );
  NAND U21998 ( .A(n20975), .B(e_input[302]), .Z(n20969) );
  NAND U21999 ( .A(n12323), .B(e_input[302]), .Z(n20975) );
  XNOR U22000 ( .A(n20965), .B(n20976), .Z(n20967) );
  XOR U22001 ( .A(n20977), .B(n20978), .Z(n20965) );
  AND U22002 ( .A(n20979), .B(n20980), .Z(n20978) );
  XNOR U22003 ( .A(n20981), .B(n20977), .Z(n20980) );
  XOR U22004 ( .A(n20982), .B(e_input[302]), .Z(n20973) );
  IV U22005 ( .A(n20971), .Z(n20982) );
  XOR U22006 ( .A(n20983), .B(n20984), .Z(n20971) );
  AND U22007 ( .A(n20985), .B(n20986), .Z(n20984) );
  XNOR U22008 ( .A(n20983), .B(n10494), .Z(n20986) );
  XNOR U22009 ( .A(n20979), .B(n20981), .Z(n10494) );
  NAND U22010 ( .A(n20987), .B(e_input[301]), .Z(n20981) );
  NAND U22011 ( .A(n12323), .B(e_input[301]), .Z(n20987) );
  XNOR U22012 ( .A(n20977), .B(n20988), .Z(n20979) );
  XOR U22013 ( .A(n20989), .B(n20990), .Z(n20977) );
  AND U22014 ( .A(n20991), .B(n20992), .Z(n20990) );
  XNOR U22015 ( .A(n20993), .B(n20989), .Z(n20992) );
  XOR U22016 ( .A(n20994), .B(e_input[301]), .Z(n20985) );
  IV U22017 ( .A(n20983), .Z(n20994) );
  XOR U22018 ( .A(n20995), .B(n20996), .Z(n20983) );
  AND U22019 ( .A(n20997), .B(n20998), .Z(n20996) );
  XNOR U22020 ( .A(n20995), .B(n10500), .Z(n20998) );
  XNOR U22021 ( .A(n20991), .B(n20993), .Z(n10500) );
  NAND U22022 ( .A(n20999), .B(e_input[300]), .Z(n20993) );
  NAND U22023 ( .A(n12323), .B(e_input[300]), .Z(n20999) );
  XNOR U22024 ( .A(n20989), .B(n21000), .Z(n20991) );
  XOR U22025 ( .A(n21001), .B(n21002), .Z(n20989) );
  AND U22026 ( .A(n21003), .B(n21004), .Z(n21002) );
  XNOR U22027 ( .A(n21005), .B(n21001), .Z(n21004) );
  XOR U22028 ( .A(n21006), .B(e_input[300]), .Z(n20997) );
  IV U22029 ( .A(n20995), .Z(n21006) );
  XOR U22030 ( .A(n21007), .B(n21008), .Z(n20995) );
  AND U22031 ( .A(n21009), .B(n21010), .Z(n21008) );
  XNOR U22032 ( .A(n21007), .B(n10506), .Z(n21010) );
  XNOR U22033 ( .A(n21003), .B(n21005), .Z(n10506) );
  NAND U22034 ( .A(n21011), .B(e_input[299]), .Z(n21005) );
  NAND U22035 ( .A(n12323), .B(e_input[299]), .Z(n21011) );
  XNOR U22036 ( .A(n21001), .B(n21012), .Z(n21003) );
  XOR U22037 ( .A(n21013), .B(n21014), .Z(n21001) );
  AND U22038 ( .A(n21015), .B(n21016), .Z(n21014) );
  XNOR U22039 ( .A(n21017), .B(n21013), .Z(n21016) );
  XOR U22040 ( .A(n21018), .B(e_input[299]), .Z(n21009) );
  IV U22041 ( .A(n21007), .Z(n21018) );
  XOR U22042 ( .A(n21019), .B(n21020), .Z(n21007) );
  AND U22043 ( .A(n21021), .B(n21022), .Z(n21020) );
  XNOR U22044 ( .A(n21019), .B(n10512), .Z(n21022) );
  XNOR U22045 ( .A(n21015), .B(n21017), .Z(n10512) );
  NAND U22046 ( .A(n21023), .B(e_input[298]), .Z(n21017) );
  NAND U22047 ( .A(n12323), .B(e_input[298]), .Z(n21023) );
  XNOR U22048 ( .A(n21013), .B(n21024), .Z(n21015) );
  XOR U22049 ( .A(n21025), .B(n21026), .Z(n21013) );
  AND U22050 ( .A(n21027), .B(n21028), .Z(n21026) );
  XNOR U22051 ( .A(n21029), .B(n21025), .Z(n21028) );
  XOR U22052 ( .A(n21030), .B(e_input[298]), .Z(n21021) );
  IV U22053 ( .A(n21019), .Z(n21030) );
  XOR U22054 ( .A(n21031), .B(n21032), .Z(n21019) );
  AND U22055 ( .A(n21033), .B(n21034), .Z(n21032) );
  XNOR U22056 ( .A(n21031), .B(n10518), .Z(n21034) );
  XNOR U22057 ( .A(n21027), .B(n21029), .Z(n10518) );
  NAND U22058 ( .A(n21035), .B(e_input[297]), .Z(n21029) );
  NAND U22059 ( .A(n12323), .B(e_input[297]), .Z(n21035) );
  XNOR U22060 ( .A(n21025), .B(n21036), .Z(n21027) );
  XOR U22061 ( .A(n21037), .B(n21038), .Z(n21025) );
  AND U22062 ( .A(n21039), .B(n21040), .Z(n21038) );
  XNOR U22063 ( .A(n21041), .B(n21037), .Z(n21040) );
  XOR U22064 ( .A(n21042), .B(e_input[297]), .Z(n21033) );
  IV U22065 ( .A(n21031), .Z(n21042) );
  XOR U22066 ( .A(n21043), .B(n21044), .Z(n21031) );
  AND U22067 ( .A(n21045), .B(n21046), .Z(n21044) );
  XNOR U22068 ( .A(n21043), .B(n10524), .Z(n21046) );
  XNOR U22069 ( .A(n21039), .B(n21041), .Z(n10524) );
  NAND U22070 ( .A(n21047), .B(e_input[296]), .Z(n21041) );
  NAND U22071 ( .A(n12323), .B(e_input[296]), .Z(n21047) );
  XNOR U22072 ( .A(n21037), .B(n21048), .Z(n21039) );
  XOR U22073 ( .A(n21049), .B(n21050), .Z(n21037) );
  AND U22074 ( .A(n21051), .B(n21052), .Z(n21050) );
  XNOR U22075 ( .A(n21053), .B(n21049), .Z(n21052) );
  XOR U22076 ( .A(n21054), .B(e_input[296]), .Z(n21045) );
  IV U22077 ( .A(n21043), .Z(n21054) );
  XOR U22078 ( .A(n21055), .B(n21056), .Z(n21043) );
  AND U22079 ( .A(n21057), .B(n21058), .Z(n21056) );
  XNOR U22080 ( .A(n21055), .B(n10530), .Z(n21058) );
  XNOR U22081 ( .A(n21051), .B(n21053), .Z(n10530) );
  NAND U22082 ( .A(n21059), .B(e_input[295]), .Z(n21053) );
  NAND U22083 ( .A(n12323), .B(e_input[295]), .Z(n21059) );
  XNOR U22084 ( .A(n21049), .B(n21060), .Z(n21051) );
  XOR U22085 ( .A(n21061), .B(n21062), .Z(n21049) );
  AND U22086 ( .A(n21063), .B(n21064), .Z(n21062) );
  XNOR U22087 ( .A(n21065), .B(n21061), .Z(n21064) );
  XOR U22088 ( .A(n21066), .B(e_input[295]), .Z(n21057) );
  IV U22089 ( .A(n21055), .Z(n21066) );
  XOR U22090 ( .A(n21067), .B(n21068), .Z(n21055) );
  AND U22091 ( .A(n21069), .B(n21070), .Z(n21068) );
  XNOR U22092 ( .A(n21067), .B(n10536), .Z(n21070) );
  XNOR U22093 ( .A(n21063), .B(n21065), .Z(n10536) );
  NAND U22094 ( .A(n21071), .B(e_input[294]), .Z(n21065) );
  NAND U22095 ( .A(n12323), .B(e_input[294]), .Z(n21071) );
  XNOR U22096 ( .A(n21061), .B(n21072), .Z(n21063) );
  XOR U22097 ( .A(n21073), .B(n21074), .Z(n21061) );
  AND U22098 ( .A(n21075), .B(n21076), .Z(n21074) );
  XNOR U22099 ( .A(n21077), .B(n21073), .Z(n21076) );
  XOR U22100 ( .A(n21078), .B(e_input[294]), .Z(n21069) );
  IV U22101 ( .A(n21067), .Z(n21078) );
  XOR U22102 ( .A(n21079), .B(n21080), .Z(n21067) );
  AND U22103 ( .A(n21081), .B(n21082), .Z(n21080) );
  XNOR U22104 ( .A(n21079), .B(n10542), .Z(n21082) );
  XNOR U22105 ( .A(n21075), .B(n21077), .Z(n10542) );
  NAND U22106 ( .A(n21083), .B(e_input[293]), .Z(n21077) );
  NAND U22107 ( .A(n12323), .B(e_input[293]), .Z(n21083) );
  XNOR U22108 ( .A(n21073), .B(n21084), .Z(n21075) );
  XOR U22109 ( .A(n21085), .B(n21086), .Z(n21073) );
  AND U22110 ( .A(n21087), .B(n21088), .Z(n21086) );
  XNOR U22111 ( .A(n21089), .B(n21085), .Z(n21088) );
  XOR U22112 ( .A(n21090), .B(e_input[293]), .Z(n21081) );
  IV U22113 ( .A(n21079), .Z(n21090) );
  XOR U22114 ( .A(n21091), .B(n21092), .Z(n21079) );
  AND U22115 ( .A(n21093), .B(n21094), .Z(n21092) );
  XNOR U22116 ( .A(n21091), .B(n10548), .Z(n21094) );
  XNOR U22117 ( .A(n21087), .B(n21089), .Z(n10548) );
  NAND U22118 ( .A(n21095), .B(e_input[292]), .Z(n21089) );
  NAND U22119 ( .A(n12323), .B(e_input[292]), .Z(n21095) );
  XNOR U22120 ( .A(n21085), .B(n21096), .Z(n21087) );
  XOR U22121 ( .A(n21097), .B(n21098), .Z(n21085) );
  AND U22122 ( .A(n21099), .B(n21100), .Z(n21098) );
  XNOR U22123 ( .A(n21101), .B(n21097), .Z(n21100) );
  XOR U22124 ( .A(n21102), .B(e_input[292]), .Z(n21093) );
  IV U22125 ( .A(n21091), .Z(n21102) );
  XOR U22126 ( .A(n21103), .B(n21104), .Z(n21091) );
  AND U22127 ( .A(n21105), .B(n21106), .Z(n21104) );
  XNOR U22128 ( .A(n21103), .B(n10554), .Z(n21106) );
  XNOR U22129 ( .A(n21099), .B(n21101), .Z(n10554) );
  NAND U22130 ( .A(n21107), .B(e_input[291]), .Z(n21101) );
  NAND U22131 ( .A(n12323), .B(e_input[291]), .Z(n21107) );
  XNOR U22132 ( .A(n21097), .B(n21108), .Z(n21099) );
  XOR U22133 ( .A(n21109), .B(n21110), .Z(n21097) );
  AND U22134 ( .A(n21111), .B(n21112), .Z(n21110) );
  XNOR U22135 ( .A(n21113), .B(n21109), .Z(n21112) );
  XOR U22136 ( .A(n21114), .B(e_input[291]), .Z(n21105) );
  IV U22137 ( .A(n21103), .Z(n21114) );
  XOR U22138 ( .A(n21115), .B(n21116), .Z(n21103) );
  AND U22139 ( .A(n21117), .B(n21118), .Z(n21116) );
  XNOR U22140 ( .A(n21115), .B(n10560), .Z(n21118) );
  XNOR U22141 ( .A(n21111), .B(n21113), .Z(n10560) );
  NAND U22142 ( .A(n21119), .B(e_input[290]), .Z(n21113) );
  NAND U22143 ( .A(n12323), .B(e_input[290]), .Z(n21119) );
  XNOR U22144 ( .A(n21109), .B(n21120), .Z(n21111) );
  XOR U22145 ( .A(n21121), .B(n21122), .Z(n21109) );
  AND U22146 ( .A(n21123), .B(n21124), .Z(n21122) );
  XNOR U22147 ( .A(n21125), .B(n21121), .Z(n21124) );
  XOR U22148 ( .A(n21126), .B(e_input[290]), .Z(n21117) );
  IV U22149 ( .A(n21115), .Z(n21126) );
  XOR U22150 ( .A(n21127), .B(n21128), .Z(n21115) );
  AND U22151 ( .A(n21129), .B(n21130), .Z(n21128) );
  XNOR U22152 ( .A(n21127), .B(n10566), .Z(n21130) );
  XNOR U22153 ( .A(n21123), .B(n21125), .Z(n10566) );
  NAND U22154 ( .A(n21131), .B(e_input[289]), .Z(n21125) );
  NAND U22155 ( .A(n12323), .B(e_input[289]), .Z(n21131) );
  XNOR U22156 ( .A(n21121), .B(n21132), .Z(n21123) );
  XOR U22157 ( .A(n21133), .B(n21134), .Z(n21121) );
  AND U22158 ( .A(n21135), .B(n21136), .Z(n21134) );
  XNOR U22159 ( .A(n21137), .B(n21133), .Z(n21136) );
  XOR U22160 ( .A(n21138), .B(e_input[289]), .Z(n21129) );
  IV U22161 ( .A(n21127), .Z(n21138) );
  XOR U22162 ( .A(n21139), .B(n21140), .Z(n21127) );
  AND U22163 ( .A(n21141), .B(n21142), .Z(n21140) );
  XNOR U22164 ( .A(n21139), .B(n10572), .Z(n21142) );
  XNOR U22165 ( .A(n21135), .B(n21137), .Z(n10572) );
  NAND U22166 ( .A(n21143), .B(e_input[288]), .Z(n21137) );
  NAND U22167 ( .A(n12323), .B(e_input[288]), .Z(n21143) );
  XNOR U22168 ( .A(n21133), .B(n21144), .Z(n21135) );
  XOR U22169 ( .A(n21145), .B(n21146), .Z(n21133) );
  AND U22170 ( .A(n21147), .B(n21148), .Z(n21146) );
  XNOR U22171 ( .A(n21149), .B(n21145), .Z(n21148) );
  XOR U22172 ( .A(n21150), .B(e_input[288]), .Z(n21141) );
  IV U22173 ( .A(n21139), .Z(n21150) );
  XOR U22174 ( .A(n21151), .B(n21152), .Z(n21139) );
  AND U22175 ( .A(n21153), .B(n21154), .Z(n21152) );
  XNOR U22176 ( .A(n21151), .B(n10578), .Z(n21154) );
  XNOR U22177 ( .A(n21147), .B(n21149), .Z(n10578) );
  NAND U22178 ( .A(n21155), .B(e_input[287]), .Z(n21149) );
  NAND U22179 ( .A(n12323), .B(e_input[287]), .Z(n21155) );
  XNOR U22180 ( .A(n21145), .B(n21156), .Z(n21147) );
  XOR U22181 ( .A(n21157), .B(n21158), .Z(n21145) );
  AND U22182 ( .A(n21159), .B(n21160), .Z(n21158) );
  XNOR U22183 ( .A(n21161), .B(n21157), .Z(n21160) );
  XOR U22184 ( .A(n21162), .B(e_input[287]), .Z(n21153) );
  IV U22185 ( .A(n21151), .Z(n21162) );
  XOR U22186 ( .A(n21163), .B(n21164), .Z(n21151) );
  AND U22187 ( .A(n21165), .B(n21166), .Z(n21164) );
  XNOR U22188 ( .A(n21163), .B(n10584), .Z(n21166) );
  XNOR U22189 ( .A(n21159), .B(n21161), .Z(n10584) );
  NAND U22190 ( .A(n21167), .B(e_input[286]), .Z(n21161) );
  NAND U22191 ( .A(n12323), .B(e_input[286]), .Z(n21167) );
  XNOR U22192 ( .A(n21157), .B(n21168), .Z(n21159) );
  XOR U22193 ( .A(n21169), .B(n21170), .Z(n21157) );
  AND U22194 ( .A(n21171), .B(n21172), .Z(n21170) );
  XNOR U22195 ( .A(n21173), .B(n21169), .Z(n21172) );
  XOR U22196 ( .A(n21174), .B(e_input[286]), .Z(n21165) );
  IV U22197 ( .A(n21163), .Z(n21174) );
  XOR U22198 ( .A(n21175), .B(n21176), .Z(n21163) );
  AND U22199 ( .A(n21177), .B(n21178), .Z(n21176) );
  XNOR U22200 ( .A(n21175), .B(n10590), .Z(n21178) );
  XNOR U22201 ( .A(n21171), .B(n21173), .Z(n10590) );
  NAND U22202 ( .A(n21179), .B(e_input[285]), .Z(n21173) );
  NAND U22203 ( .A(n12323), .B(e_input[285]), .Z(n21179) );
  XNOR U22204 ( .A(n21169), .B(n21180), .Z(n21171) );
  XOR U22205 ( .A(n21181), .B(n21182), .Z(n21169) );
  AND U22206 ( .A(n21183), .B(n21184), .Z(n21182) );
  XNOR U22207 ( .A(n21185), .B(n21181), .Z(n21184) );
  XOR U22208 ( .A(n21186), .B(e_input[285]), .Z(n21177) );
  IV U22209 ( .A(n21175), .Z(n21186) );
  XOR U22210 ( .A(n21187), .B(n21188), .Z(n21175) );
  AND U22211 ( .A(n21189), .B(n21190), .Z(n21188) );
  XNOR U22212 ( .A(n21187), .B(n10596), .Z(n21190) );
  XNOR U22213 ( .A(n21183), .B(n21185), .Z(n10596) );
  NAND U22214 ( .A(n21191), .B(e_input[284]), .Z(n21185) );
  NAND U22215 ( .A(n12323), .B(e_input[284]), .Z(n21191) );
  XNOR U22216 ( .A(n21181), .B(n21192), .Z(n21183) );
  XOR U22217 ( .A(n21193), .B(n21194), .Z(n21181) );
  AND U22218 ( .A(n21195), .B(n21196), .Z(n21194) );
  XNOR U22219 ( .A(n21197), .B(n21193), .Z(n21196) );
  XOR U22220 ( .A(n21198), .B(e_input[284]), .Z(n21189) );
  IV U22221 ( .A(n21187), .Z(n21198) );
  XOR U22222 ( .A(n21199), .B(n21200), .Z(n21187) );
  AND U22223 ( .A(n21201), .B(n21202), .Z(n21200) );
  XNOR U22224 ( .A(n21199), .B(n10602), .Z(n21202) );
  XNOR U22225 ( .A(n21195), .B(n21197), .Z(n10602) );
  NAND U22226 ( .A(n21203), .B(e_input[283]), .Z(n21197) );
  NAND U22227 ( .A(n12323), .B(e_input[283]), .Z(n21203) );
  XNOR U22228 ( .A(n21193), .B(n21204), .Z(n21195) );
  XOR U22229 ( .A(n21205), .B(n21206), .Z(n21193) );
  AND U22230 ( .A(n21207), .B(n21208), .Z(n21206) );
  XNOR U22231 ( .A(n21209), .B(n21205), .Z(n21208) );
  XOR U22232 ( .A(n21210), .B(e_input[283]), .Z(n21201) );
  IV U22233 ( .A(n21199), .Z(n21210) );
  XOR U22234 ( .A(n21211), .B(n21212), .Z(n21199) );
  AND U22235 ( .A(n21213), .B(n21214), .Z(n21212) );
  XNOR U22236 ( .A(n21211), .B(n10608), .Z(n21214) );
  XNOR U22237 ( .A(n21207), .B(n21209), .Z(n10608) );
  NAND U22238 ( .A(n21215), .B(e_input[282]), .Z(n21209) );
  NAND U22239 ( .A(n12323), .B(e_input[282]), .Z(n21215) );
  XNOR U22240 ( .A(n21205), .B(n21216), .Z(n21207) );
  XOR U22241 ( .A(n21217), .B(n21218), .Z(n21205) );
  AND U22242 ( .A(n21219), .B(n21220), .Z(n21218) );
  XNOR U22243 ( .A(n21221), .B(n21217), .Z(n21220) );
  XOR U22244 ( .A(n21222), .B(e_input[282]), .Z(n21213) );
  IV U22245 ( .A(n21211), .Z(n21222) );
  XOR U22246 ( .A(n21223), .B(n21224), .Z(n21211) );
  AND U22247 ( .A(n21225), .B(n21226), .Z(n21224) );
  XNOR U22248 ( .A(n21223), .B(n10614), .Z(n21226) );
  XNOR U22249 ( .A(n21219), .B(n21221), .Z(n10614) );
  NAND U22250 ( .A(n21227), .B(e_input[281]), .Z(n21221) );
  NAND U22251 ( .A(n12323), .B(e_input[281]), .Z(n21227) );
  XNOR U22252 ( .A(n21217), .B(n21228), .Z(n21219) );
  XOR U22253 ( .A(n21229), .B(n21230), .Z(n21217) );
  AND U22254 ( .A(n21231), .B(n21232), .Z(n21230) );
  XNOR U22255 ( .A(n21233), .B(n21229), .Z(n21232) );
  XOR U22256 ( .A(n21234), .B(e_input[281]), .Z(n21225) );
  IV U22257 ( .A(n21223), .Z(n21234) );
  XOR U22258 ( .A(n21235), .B(n21236), .Z(n21223) );
  AND U22259 ( .A(n21237), .B(n21238), .Z(n21236) );
  XNOR U22260 ( .A(n21235), .B(n10620), .Z(n21238) );
  XNOR U22261 ( .A(n21231), .B(n21233), .Z(n10620) );
  NAND U22262 ( .A(n21239), .B(e_input[280]), .Z(n21233) );
  NAND U22263 ( .A(n12323), .B(e_input[280]), .Z(n21239) );
  XNOR U22264 ( .A(n21229), .B(n21240), .Z(n21231) );
  XOR U22265 ( .A(n21241), .B(n21242), .Z(n21229) );
  AND U22266 ( .A(n21243), .B(n21244), .Z(n21242) );
  XNOR U22267 ( .A(n21245), .B(n21241), .Z(n21244) );
  XOR U22268 ( .A(n21246), .B(e_input[280]), .Z(n21237) );
  IV U22269 ( .A(n21235), .Z(n21246) );
  XOR U22270 ( .A(n21247), .B(n21248), .Z(n21235) );
  AND U22271 ( .A(n21249), .B(n21250), .Z(n21248) );
  XNOR U22272 ( .A(n21247), .B(n10626), .Z(n21250) );
  XNOR U22273 ( .A(n21243), .B(n21245), .Z(n10626) );
  NAND U22274 ( .A(n21251), .B(e_input[279]), .Z(n21245) );
  NAND U22275 ( .A(n12323), .B(e_input[279]), .Z(n21251) );
  XNOR U22276 ( .A(n21241), .B(n21252), .Z(n21243) );
  XOR U22277 ( .A(n21253), .B(n21254), .Z(n21241) );
  AND U22278 ( .A(n21255), .B(n21256), .Z(n21254) );
  XNOR U22279 ( .A(n21257), .B(n21253), .Z(n21256) );
  XOR U22280 ( .A(n21258), .B(e_input[279]), .Z(n21249) );
  IV U22281 ( .A(n21247), .Z(n21258) );
  XOR U22282 ( .A(n21259), .B(n21260), .Z(n21247) );
  AND U22283 ( .A(n21261), .B(n21262), .Z(n21260) );
  XNOR U22284 ( .A(n21259), .B(n10632), .Z(n21262) );
  XNOR U22285 ( .A(n21255), .B(n21257), .Z(n10632) );
  NAND U22286 ( .A(n21263), .B(e_input[278]), .Z(n21257) );
  NAND U22287 ( .A(n12323), .B(e_input[278]), .Z(n21263) );
  XNOR U22288 ( .A(n21253), .B(n21264), .Z(n21255) );
  XOR U22289 ( .A(n21265), .B(n21266), .Z(n21253) );
  AND U22290 ( .A(n21267), .B(n21268), .Z(n21266) );
  XNOR U22291 ( .A(n21269), .B(n21265), .Z(n21268) );
  XOR U22292 ( .A(n21270), .B(e_input[278]), .Z(n21261) );
  IV U22293 ( .A(n21259), .Z(n21270) );
  XOR U22294 ( .A(n21271), .B(n21272), .Z(n21259) );
  AND U22295 ( .A(n21273), .B(n21274), .Z(n21272) );
  XNOR U22296 ( .A(n21271), .B(n10638), .Z(n21274) );
  XNOR U22297 ( .A(n21267), .B(n21269), .Z(n10638) );
  NAND U22298 ( .A(n21275), .B(e_input[277]), .Z(n21269) );
  NAND U22299 ( .A(n12323), .B(e_input[277]), .Z(n21275) );
  XNOR U22300 ( .A(n21265), .B(n21276), .Z(n21267) );
  XOR U22301 ( .A(n21277), .B(n21278), .Z(n21265) );
  AND U22302 ( .A(n21279), .B(n21280), .Z(n21278) );
  XNOR U22303 ( .A(n21281), .B(n21277), .Z(n21280) );
  XOR U22304 ( .A(n21282), .B(e_input[277]), .Z(n21273) );
  IV U22305 ( .A(n21271), .Z(n21282) );
  XOR U22306 ( .A(n21283), .B(n21284), .Z(n21271) );
  AND U22307 ( .A(n21285), .B(n21286), .Z(n21284) );
  XNOR U22308 ( .A(n21283), .B(n10644), .Z(n21286) );
  XNOR U22309 ( .A(n21279), .B(n21281), .Z(n10644) );
  NAND U22310 ( .A(n21287), .B(e_input[276]), .Z(n21281) );
  NAND U22311 ( .A(n12323), .B(e_input[276]), .Z(n21287) );
  XNOR U22312 ( .A(n21277), .B(n21288), .Z(n21279) );
  XOR U22313 ( .A(n21289), .B(n21290), .Z(n21277) );
  AND U22314 ( .A(n21291), .B(n21292), .Z(n21290) );
  XNOR U22315 ( .A(n21293), .B(n21289), .Z(n21292) );
  XOR U22316 ( .A(n21294), .B(e_input[276]), .Z(n21285) );
  IV U22317 ( .A(n21283), .Z(n21294) );
  XOR U22318 ( .A(n21295), .B(n21296), .Z(n21283) );
  AND U22319 ( .A(n21297), .B(n21298), .Z(n21296) );
  XNOR U22320 ( .A(n21295), .B(n10650), .Z(n21298) );
  XNOR U22321 ( .A(n21291), .B(n21293), .Z(n10650) );
  NAND U22322 ( .A(n21299), .B(e_input[275]), .Z(n21293) );
  NAND U22323 ( .A(n12323), .B(e_input[275]), .Z(n21299) );
  XNOR U22324 ( .A(n21289), .B(n21300), .Z(n21291) );
  XOR U22325 ( .A(n21301), .B(n21302), .Z(n21289) );
  AND U22326 ( .A(n21303), .B(n21304), .Z(n21302) );
  XNOR U22327 ( .A(n21305), .B(n21301), .Z(n21304) );
  XOR U22328 ( .A(n21306), .B(e_input[275]), .Z(n21297) );
  IV U22329 ( .A(n21295), .Z(n21306) );
  XOR U22330 ( .A(n21307), .B(n21308), .Z(n21295) );
  AND U22331 ( .A(n21309), .B(n21310), .Z(n21308) );
  XNOR U22332 ( .A(n21307), .B(n10656), .Z(n21310) );
  XNOR U22333 ( .A(n21303), .B(n21305), .Z(n10656) );
  NAND U22334 ( .A(n21311), .B(e_input[274]), .Z(n21305) );
  NAND U22335 ( .A(n12323), .B(e_input[274]), .Z(n21311) );
  XNOR U22336 ( .A(n21301), .B(n21312), .Z(n21303) );
  XOR U22337 ( .A(n21313), .B(n21314), .Z(n21301) );
  AND U22338 ( .A(n21315), .B(n21316), .Z(n21314) );
  XNOR U22339 ( .A(n21317), .B(n21313), .Z(n21316) );
  XOR U22340 ( .A(n21318), .B(e_input[274]), .Z(n21309) );
  IV U22341 ( .A(n21307), .Z(n21318) );
  XOR U22342 ( .A(n21319), .B(n21320), .Z(n21307) );
  AND U22343 ( .A(n21321), .B(n21322), .Z(n21320) );
  XNOR U22344 ( .A(n21319), .B(n10662), .Z(n21322) );
  XNOR U22345 ( .A(n21315), .B(n21317), .Z(n10662) );
  NAND U22346 ( .A(n21323), .B(e_input[273]), .Z(n21317) );
  NAND U22347 ( .A(n12323), .B(e_input[273]), .Z(n21323) );
  XNOR U22348 ( .A(n21313), .B(n21324), .Z(n21315) );
  XOR U22349 ( .A(n21325), .B(n21326), .Z(n21313) );
  AND U22350 ( .A(n21327), .B(n21328), .Z(n21326) );
  XNOR U22351 ( .A(n21329), .B(n21325), .Z(n21328) );
  XOR U22352 ( .A(n21330), .B(e_input[273]), .Z(n21321) );
  IV U22353 ( .A(n21319), .Z(n21330) );
  XOR U22354 ( .A(n21331), .B(n21332), .Z(n21319) );
  AND U22355 ( .A(n21333), .B(n21334), .Z(n21332) );
  XNOR U22356 ( .A(n21331), .B(n10668), .Z(n21334) );
  XNOR U22357 ( .A(n21327), .B(n21329), .Z(n10668) );
  NAND U22358 ( .A(n21335), .B(e_input[272]), .Z(n21329) );
  NAND U22359 ( .A(n12323), .B(e_input[272]), .Z(n21335) );
  XNOR U22360 ( .A(n21325), .B(n21336), .Z(n21327) );
  XOR U22361 ( .A(n21337), .B(n21338), .Z(n21325) );
  AND U22362 ( .A(n21339), .B(n21340), .Z(n21338) );
  XNOR U22363 ( .A(n21341), .B(n21337), .Z(n21340) );
  XOR U22364 ( .A(n21342), .B(e_input[272]), .Z(n21333) );
  IV U22365 ( .A(n21331), .Z(n21342) );
  XOR U22366 ( .A(n21343), .B(n21344), .Z(n21331) );
  AND U22367 ( .A(n21345), .B(n21346), .Z(n21344) );
  XNOR U22368 ( .A(n21343), .B(n10674), .Z(n21346) );
  XNOR U22369 ( .A(n21339), .B(n21341), .Z(n10674) );
  NAND U22370 ( .A(n21347), .B(e_input[271]), .Z(n21341) );
  NAND U22371 ( .A(n12323), .B(e_input[271]), .Z(n21347) );
  XNOR U22372 ( .A(n21337), .B(n21348), .Z(n21339) );
  XOR U22373 ( .A(n21349), .B(n21350), .Z(n21337) );
  AND U22374 ( .A(n21351), .B(n21352), .Z(n21350) );
  XNOR U22375 ( .A(n21353), .B(n21349), .Z(n21352) );
  XOR U22376 ( .A(n21354), .B(e_input[271]), .Z(n21345) );
  IV U22377 ( .A(n21343), .Z(n21354) );
  XOR U22378 ( .A(n21355), .B(n21356), .Z(n21343) );
  AND U22379 ( .A(n21357), .B(n21358), .Z(n21356) );
  XNOR U22380 ( .A(n21355), .B(n10680), .Z(n21358) );
  XNOR U22381 ( .A(n21351), .B(n21353), .Z(n10680) );
  NAND U22382 ( .A(n21359), .B(e_input[270]), .Z(n21353) );
  NAND U22383 ( .A(n12323), .B(e_input[270]), .Z(n21359) );
  XNOR U22384 ( .A(n21349), .B(n21360), .Z(n21351) );
  XOR U22385 ( .A(n21361), .B(n21362), .Z(n21349) );
  AND U22386 ( .A(n21363), .B(n21364), .Z(n21362) );
  XNOR U22387 ( .A(n21365), .B(n21361), .Z(n21364) );
  XOR U22388 ( .A(n21366), .B(e_input[270]), .Z(n21357) );
  IV U22389 ( .A(n21355), .Z(n21366) );
  XOR U22390 ( .A(n21367), .B(n21368), .Z(n21355) );
  AND U22391 ( .A(n21369), .B(n21370), .Z(n21368) );
  XNOR U22392 ( .A(n21367), .B(n10686), .Z(n21370) );
  XNOR U22393 ( .A(n21363), .B(n21365), .Z(n10686) );
  NAND U22394 ( .A(n21371), .B(e_input[269]), .Z(n21365) );
  NAND U22395 ( .A(n12323), .B(e_input[269]), .Z(n21371) );
  XNOR U22396 ( .A(n21361), .B(n21372), .Z(n21363) );
  XOR U22397 ( .A(n21373), .B(n21374), .Z(n21361) );
  AND U22398 ( .A(n21375), .B(n21376), .Z(n21374) );
  XNOR U22399 ( .A(n21377), .B(n21373), .Z(n21376) );
  XOR U22400 ( .A(n21378), .B(e_input[269]), .Z(n21369) );
  IV U22401 ( .A(n21367), .Z(n21378) );
  XOR U22402 ( .A(n21379), .B(n21380), .Z(n21367) );
  AND U22403 ( .A(n21381), .B(n21382), .Z(n21380) );
  XNOR U22404 ( .A(n21379), .B(n10692), .Z(n21382) );
  XNOR U22405 ( .A(n21375), .B(n21377), .Z(n10692) );
  NAND U22406 ( .A(n21383), .B(e_input[268]), .Z(n21377) );
  NAND U22407 ( .A(n12323), .B(e_input[268]), .Z(n21383) );
  XNOR U22408 ( .A(n21373), .B(n21384), .Z(n21375) );
  XOR U22409 ( .A(n21385), .B(n21386), .Z(n21373) );
  AND U22410 ( .A(n21387), .B(n21388), .Z(n21386) );
  XNOR U22411 ( .A(n21389), .B(n21385), .Z(n21388) );
  XOR U22412 ( .A(n21390), .B(e_input[268]), .Z(n21381) );
  IV U22413 ( .A(n21379), .Z(n21390) );
  XOR U22414 ( .A(n21391), .B(n21392), .Z(n21379) );
  AND U22415 ( .A(n21393), .B(n21394), .Z(n21392) );
  XNOR U22416 ( .A(n21391), .B(n10698), .Z(n21394) );
  XNOR U22417 ( .A(n21387), .B(n21389), .Z(n10698) );
  NAND U22418 ( .A(n21395), .B(e_input[267]), .Z(n21389) );
  NAND U22419 ( .A(n12323), .B(e_input[267]), .Z(n21395) );
  XNOR U22420 ( .A(n21385), .B(n21396), .Z(n21387) );
  XOR U22421 ( .A(n21397), .B(n21398), .Z(n21385) );
  AND U22422 ( .A(n21399), .B(n21400), .Z(n21398) );
  XNOR U22423 ( .A(n21401), .B(n21397), .Z(n21400) );
  XOR U22424 ( .A(n21402), .B(e_input[267]), .Z(n21393) );
  IV U22425 ( .A(n21391), .Z(n21402) );
  XOR U22426 ( .A(n21403), .B(n21404), .Z(n21391) );
  AND U22427 ( .A(n21405), .B(n21406), .Z(n21404) );
  XNOR U22428 ( .A(n21403), .B(n10704), .Z(n21406) );
  XNOR U22429 ( .A(n21399), .B(n21401), .Z(n10704) );
  NAND U22430 ( .A(n21407), .B(e_input[266]), .Z(n21401) );
  NAND U22431 ( .A(n12323), .B(e_input[266]), .Z(n21407) );
  XNOR U22432 ( .A(n21397), .B(n21408), .Z(n21399) );
  XOR U22433 ( .A(n21409), .B(n21410), .Z(n21397) );
  AND U22434 ( .A(n21411), .B(n21412), .Z(n21410) );
  XNOR U22435 ( .A(n21413), .B(n21409), .Z(n21412) );
  XOR U22436 ( .A(n21414), .B(e_input[266]), .Z(n21405) );
  IV U22437 ( .A(n21403), .Z(n21414) );
  XOR U22438 ( .A(n21415), .B(n21416), .Z(n21403) );
  AND U22439 ( .A(n21417), .B(n21418), .Z(n21416) );
  XNOR U22440 ( .A(n21415), .B(n10710), .Z(n21418) );
  XNOR U22441 ( .A(n21411), .B(n21413), .Z(n10710) );
  NAND U22442 ( .A(n21419), .B(e_input[265]), .Z(n21413) );
  NAND U22443 ( .A(n12323), .B(e_input[265]), .Z(n21419) );
  XNOR U22444 ( .A(n21409), .B(n21420), .Z(n21411) );
  XOR U22445 ( .A(n21421), .B(n21422), .Z(n21409) );
  AND U22446 ( .A(n21423), .B(n21424), .Z(n21422) );
  XNOR U22447 ( .A(n21425), .B(n21421), .Z(n21424) );
  XOR U22448 ( .A(n21426), .B(e_input[265]), .Z(n21417) );
  IV U22449 ( .A(n21415), .Z(n21426) );
  XOR U22450 ( .A(n21427), .B(n21428), .Z(n21415) );
  AND U22451 ( .A(n21429), .B(n21430), .Z(n21428) );
  XNOR U22452 ( .A(n21427), .B(n10716), .Z(n21430) );
  XNOR U22453 ( .A(n21423), .B(n21425), .Z(n10716) );
  NAND U22454 ( .A(n21431), .B(e_input[264]), .Z(n21425) );
  NAND U22455 ( .A(n12323), .B(e_input[264]), .Z(n21431) );
  XNOR U22456 ( .A(n21421), .B(n21432), .Z(n21423) );
  XOR U22457 ( .A(n21433), .B(n21434), .Z(n21421) );
  AND U22458 ( .A(n21435), .B(n21436), .Z(n21434) );
  XNOR U22459 ( .A(n21437), .B(n21433), .Z(n21436) );
  XOR U22460 ( .A(n21438), .B(e_input[264]), .Z(n21429) );
  IV U22461 ( .A(n21427), .Z(n21438) );
  XOR U22462 ( .A(n21439), .B(n21440), .Z(n21427) );
  AND U22463 ( .A(n21441), .B(n21442), .Z(n21440) );
  XNOR U22464 ( .A(n21439), .B(n10722), .Z(n21442) );
  XNOR U22465 ( .A(n21435), .B(n21437), .Z(n10722) );
  NAND U22466 ( .A(n21443), .B(e_input[263]), .Z(n21437) );
  NAND U22467 ( .A(n12323), .B(e_input[263]), .Z(n21443) );
  XNOR U22468 ( .A(n21433), .B(n21444), .Z(n21435) );
  XOR U22469 ( .A(n21445), .B(n21446), .Z(n21433) );
  AND U22470 ( .A(n21447), .B(n21448), .Z(n21446) );
  XNOR U22471 ( .A(n21449), .B(n21445), .Z(n21448) );
  XOR U22472 ( .A(n21450), .B(e_input[263]), .Z(n21441) );
  IV U22473 ( .A(n21439), .Z(n21450) );
  XOR U22474 ( .A(n21451), .B(n21452), .Z(n21439) );
  AND U22475 ( .A(n21453), .B(n21454), .Z(n21452) );
  XNOR U22476 ( .A(n21451), .B(n10728), .Z(n21454) );
  XNOR U22477 ( .A(n21447), .B(n21449), .Z(n10728) );
  NAND U22478 ( .A(n21455), .B(e_input[262]), .Z(n21449) );
  NAND U22479 ( .A(n12323), .B(e_input[262]), .Z(n21455) );
  XNOR U22480 ( .A(n21445), .B(n21456), .Z(n21447) );
  XOR U22481 ( .A(n21457), .B(n21458), .Z(n21445) );
  AND U22482 ( .A(n21459), .B(n21460), .Z(n21458) );
  XNOR U22483 ( .A(n21461), .B(n21457), .Z(n21460) );
  XOR U22484 ( .A(n21462), .B(e_input[262]), .Z(n21453) );
  IV U22485 ( .A(n21451), .Z(n21462) );
  XOR U22486 ( .A(n21463), .B(n21464), .Z(n21451) );
  AND U22487 ( .A(n21465), .B(n21466), .Z(n21464) );
  XNOR U22488 ( .A(n21463), .B(n10734), .Z(n21466) );
  XNOR U22489 ( .A(n21459), .B(n21461), .Z(n10734) );
  NAND U22490 ( .A(n21467), .B(e_input[261]), .Z(n21461) );
  NAND U22491 ( .A(n12323), .B(e_input[261]), .Z(n21467) );
  XNOR U22492 ( .A(n21457), .B(n21468), .Z(n21459) );
  XOR U22493 ( .A(n21469), .B(n21470), .Z(n21457) );
  AND U22494 ( .A(n21471), .B(n21472), .Z(n21470) );
  XNOR U22495 ( .A(n21473), .B(n21469), .Z(n21472) );
  XOR U22496 ( .A(n21474), .B(e_input[261]), .Z(n21465) );
  IV U22497 ( .A(n21463), .Z(n21474) );
  XOR U22498 ( .A(n21475), .B(n21476), .Z(n21463) );
  AND U22499 ( .A(n21477), .B(n21478), .Z(n21476) );
  XNOR U22500 ( .A(n21475), .B(n10740), .Z(n21478) );
  XNOR U22501 ( .A(n21471), .B(n21473), .Z(n10740) );
  NAND U22502 ( .A(n21479), .B(e_input[260]), .Z(n21473) );
  NAND U22503 ( .A(n12323), .B(e_input[260]), .Z(n21479) );
  XNOR U22504 ( .A(n21469), .B(n21480), .Z(n21471) );
  XOR U22505 ( .A(n21481), .B(n21482), .Z(n21469) );
  AND U22506 ( .A(n21483), .B(n21484), .Z(n21482) );
  XNOR U22507 ( .A(n21485), .B(n21481), .Z(n21484) );
  XOR U22508 ( .A(n21486), .B(e_input[260]), .Z(n21477) );
  IV U22509 ( .A(n21475), .Z(n21486) );
  XOR U22510 ( .A(n21487), .B(n21488), .Z(n21475) );
  AND U22511 ( .A(n21489), .B(n21490), .Z(n21488) );
  XNOR U22512 ( .A(n21487), .B(n10746), .Z(n21490) );
  XNOR U22513 ( .A(n21483), .B(n21485), .Z(n10746) );
  NAND U22514 ( .A(n21491), .B(e_input[259]), .Z(n21485) );
  NAND U22515 ( .A(n12323), .B(e_input[259]), .Z(n21491) );
  XNOR U22516 ( .A(n21481), .B(n21492), .Z(n21483) );
  XOR U22517 ( .A(n21493), .B(n21494), .Z(n21481) );
  AND U22518 ( .A(n21495), .B(n21496), .Z(n21494) );
  XNOR U22519 ( .A(n21497), .B(n21493), .Z(n21496) );
  XOR U22520 ( .A(n21498), .B(e_input[259]), .Z(n21489) );
  IV U22521 ( .A(n21487), .Z(n21498) );
  XOR U22522 ( .A(n21499), .B(n21500), .Z(n21487) );
  AND U22523 ( .A(n21501), .B(n21502), .Z(n21500) );
  XNOR U22524 ( .A(n21499), .B(n10752), .Z(n21502) );
  XNOR U22525 ( .A(n21495), .B(n21497), .Z(n10752) );
  NAND U22526 ( .A(n21503), .B(e_input[258]), .Z(n21497) );
  NAND U22527 ( .A(n12323), .B(e_input[258]), .Z(n21503) );
  XNOR U22528 ( .A(n21493), .B(n21504), .Z(n21495) );
  XOR U22529 ( .A(n21505), .B(n21506), .Z(n21493) );
  AND U22530 ( .A(n21507), .B(n21508), .Z(n21506) );
  XNOR U22531 ( .A(n21509), .B(n21505), .Z(n21508) );
  XOR U22532 ( .A(n21510), .B(e_input[258]), .Z(n21501) );
  IV U22533 ( .A(n21499), .Z(n21510) );
  XOR U22534 ( .A(n21511), .B(n21512), .Z(n21499) );
  AND U22535 ( .A(n21513), .B(n21514), .Z(n21512) );
  XNOR U22536 ( .A(n21511), .B(n10758), .Z(n21514) );
  XNOR U22537 ( .A(n21507), .B(n21509), .Z(n10758) );
  NAND U22538 ( .A(n21515), .B(e_input[257]), .Z(n21509) );
  NAND U22539 ( .A(n12323), .B(e_input[257]), .Z(n21515) );
  XNOR U22540 ( .A(n21505), .B(n21516), .Z(n21507) );
  XOR U22541 ( .A(n21517), .B(n21518), .Z(n21505) );
  AND U22542 ( .A(n21519), .B(n21520), .Z(n21518) );
  XNOR U22543 ( .A(n21521), .B(n21517), .Z(n21520) );
  XOR U22544 ( .A(n21522), .B(e_input[257]), .Z(n21513) );
  IV U22545 ( .A(n21511), .Z(n21522) );
  XOR U22546 ( .A(n21523), .B(n21524), .Z(n21511) );
  AND U22547 ( .A(n21525), .B(n21526), .Z(n21524) );
  XNOR U22548 ( .A(n21523), .B(n10764), .Z(n21526) );
  XNOR U22549 ( .A(n21519), .B(n21521), .Z(n10764) );
  NAND U22550 ( .A(n21527), .B(e_input[256]), .Z(n21521) );
  NAND U22551 ( .A(n12323), .B(e_input[256]), .Z(n21527) );
  XNOR U22552 ( .A(n21517), .B(n21528), .Z(n21519) );
  XOR U22553 ( .A(n21529), .B(n21530), .Z(n21517) );
  AND U22554 ( .A(n21531), .B(n21532), .Z(n21530) );
  XNOR U22555 ( .A(n21533), .B(n21529), .Z(n21532) );
  XOR U22556 ( .A(n21534), .B(e_input[256]), .Z(n21525) );
  IV U22557 ( .A(n21523), .Z(n21534) );
  XOR U22558 ( .A(n21535), .B(n21536), .Z(n21523) );
  AND U22559 ( .A(n21537), .B(n21538), .Z(n21536) );
  XNOR U22560 ( .A(n21535), .B(n10770), .Z(n21538) );
  XNOR U22561 ( .A(n21531), .B(n21533), .Z(n10770) );
  NAND U22562 ( .A(n21539), .B(e_input[255]), .Z(n21533) );
  NAND U22563 ( .A(n12323), .B(e_input[255]), .Z(n21539) );
  XNOR U22564 ( .A(n21529), .B(n21540), .Z(n21531) );
  XOR U22565 ( .A(n21541), .B(n21542), .Z(n21529) );
  AND U22566 ( .A(n21543), .B(n21544), .Z(n21542) );
  XNOR U22567 ( .A(n21545), .B(n21541), .Z(n21544) );
  XOR U22568 ( .A(n21546), .B(e_input[255]), .Z(n21537) );
  IV U22569 ( .A(n21535), .Z(n21546) );
  XOR U22570 ( .A(n21547), .B(n21548), .Z(n21535) );
  AND U22571 ( .A(n21549), .B(n21550), .Z(n21548) );
  XNOR U22572 ( .A(n21547), .B(n10776), .Z(n21550) );
  XNOR U22573 ( .A(n21543), .B(n21545), .Z(n10776) );
  NAND U22574 ( .A(n21551), .B(e_input[254]), .Z(n21545) );
  NAND U22575 ( .A(n12323), .B(e_input[254]), .Z(n21551) );
  XNOR U22576 ( .A(n21541), .B(n21552), .Z(n21543) );
  XOR U22577 ( .A(n21553), .B(n21554), .Z(n21541) );
  AND U22578 ( .A(n21555), .B(n21556), .Z(n21554) );
  XNOR U22579 ( .A(n21557), .B(n21553), .Z(n21556) );
  XOR U22580 ( .A(n21558), .B(e_input[254]), .Z(n21549) );
  IV U22581 ( .A(n21547), .Z(n21558) );
  XOR U22582 ( .A(n21559), .B(n21560), .Z(n21547) );
  AND U22583 ( .A(n21561), .B(n21562), .Z(n21560) );
  XNOR U22584 ( .A(n21559), .B(n10782), .Z(n21562) );
  XNOR U22585 ( .A(n21555), .B(n21557), .Z(n10782) );
  NAND U22586 ( .A(n21563), .B(e_input[253]), .Z(n21557) );
  NAND U22587 ( .A(n12323), .B(e_input[253]), .Z(n21563) );
  XNOR U22588 ( .A(n21553), .B(n21564), .Z(n21555) );
  XOR U22589 ( .A(n21565), .B(n21566), .Z(n21553) );
  AND U22590 ( .A(n21567), .B(n21568), .Z(n21566) );
  XNOR U22591 ( .A(n21569), .B(n21565), .Z(n21568) );
  XOR U22592 ( .A(n21570), .B(e_input[253]), .Z(n21561) );
  IV U22593 ( .A(n21559), .Z(n21570) );
  XOR U22594 ( .A(n21571), .B(n21572), .Z(n21559) );
  AND U22595 ( .A(n21573), .B(n21574), .Z(n21572) );
  XNOR U22596 ( .A(n21571), .B(n10788), .Z(n21574) );
  XNOR U22597 ( .A(n21567), .B(n21569), .Z(n10788) );
  NAND U22598 ( .A(n21575), .B(e_input[252]), .Z(n21569) );
  NAND U22599 ( .A(n12323), .B(e_input[252]), .Z(n21575) );
  XNOR U22600 ( .A(n21565), .B(n21576), .Z(n21567) );
  XOR U22601 ( .A(n21577), .B(n21578), .Z(n21565) );
  AND U22602 ( .A(n21579), .B(n21580), .Z(n21578) );
  XNOR U22603 ( .A(n21581), .B(n21577), .Z(n21580) );
  XOR U22604 ( .A(n21582), .B(e_input[252]), .Z(n21573) );
  IV U22605 ( .A(n21571), .Z(n21582) );
  XOR U22606 ( .A(n21583), .B(n21584), .Z(n21571) );
  AND U22607 ( .A(n21585), .B(n21586), .Z(n21584) );
  XNOR U22608 ( .A(n21583), .B(n10794), .Z(n21586) );
  XNOR U22609 ( .A(n21579), .B(n21581), .Z(n10794) );
  NAND U22610 ( .A(n21587), .B(e_input[251]), .Z(n21581) );
  NAND U22611 ( .A(n12323), .B(e_input[251]), .Z(n21587) );
  XNOR U22612 ( .A(n21577), .B(n21588), .Z(n21579) );
  XOR U22613 ( .A(n21589), .B(n21590), .Z(n21577) );
  AND U22614 ( .A(n21591), .B(n21592), .Z(n21590) );
  XNOR U22615 ( .A(n21593), .B(n21589), .Z(n21592) );
  XOR U22616 ( .A(n21594), .B(e_input[251]), .Z(n21585) );
  IV U22617 ( .A(n21583), .Z(n21594) );
  XOR U22618 ( .A(n21595), .B(n21596), .Z(n21583) );
  AND U22619 ( .A(n21597), .B(n21598), .Z(n21596) );
  XNOR U22620 ( .A(n21595), .B(n10800), .Z(n21598) );
  XNOR U22621 ( .A(n21591), .B(n21593), .Z(n10800) );
  NAND U22622 ( .A(n21599), .B(e_input[250]), .Z(n21593) );
  NAND U22623 ( .A(n12323), .B(e_input[250]), .Z(n21599) );
  XNOR U22624 ( .A(n21589), .B(n21600), .Z(n21591) );
  XOR U22625 ( .A(n21601), .B(n21602), .Z(n21589) );
  AND U22626 ( .A(n21603), .B(n21604), .Z(n21602) );
  XNOR U22627 ( .A(n21605), .B(n21601), .Z(n21604) );
  XOR U22628 ( .A(n21606), .B(e_input[250]), .Z(n21597) );
  IV U22629 ( .A(n21595), .Z(n21606) );
  XOR U22630 ( .A(n21607), .B(n21608), .Z(n21595) );
  AND U22631 ( .A(n21609), .B(n21610), .Z(n21608) );
  XNOR U22632 ( .A(n21607), .B(n10806), .Z(n21610) );
  XNOR U22633 ( .A(n21603), .B(n21605), .Z(n10806) );
  NAND U22634 ( .A(n21611), .B(e_input[249]), .Z(n21605) );
  NAND U22635 ( .A(n12323), .B(e_input[249]), .Z(n21611) );
  XNOR U22636 ( .A(n21601), .B(n21612), .Z(n21603) );
  XOR U22637 ( .A(n21613), .B(n21614), .Z(n21601) );
  AND U22638 ( .A(n21615), .B(n21616), .Z(n21614) );
  XNOR U22639 ( .A(n21617), .B(n21613), .Z(n21616) );
  XOR U22640 ( .A(n21618), .B(e_input[249]), .Z(n21609) );
  IV U22641 ( .A(n21607), .Z(n21618) );
  XOR U22642 ( .A(n21619), .B(n21620), .Z(n21607) );
  AND U22643 ( .A(n21621), .B(n21622), .Z(n21620) );
  XNOR U22644 ( .A(n21619), .B(n10812), .Z(n21622) );
  XNOR U22645 ( .A(n21615), .B(n21617), .Z(n10812) );
  NAND U22646 ( .A(n21623), .B(e_input[248]), .Z(n21617) );
  NAND U22647 ( .A(n12323), .B(e_input[248]), .Z(n21623) );
  XNOR U22648 ( .A(n21613), .B(n21624), .Z(n21615) );
  XOR U22649 ( .A(n21625), .B(n21626), .Z(n21613) );
  AND U22650 ( .A(n21627), .B(n21628), .Z(n21626) );
  XNOR U22651 ( .A(n21629), .B(n21625), .Z(n21628) );
  XOR U22652 ( .A(n21630), .B(e_input[248]), .Z(n21621) );
  IV U22653 ( .A(n21619), .Z(n21630) );
  XOR U22654 ( .A(n21631), .B(n21632), .Z(n21619) );
  AND U22655 ( .A(n21633), .B(n21634), .Z(n21632) );
  XNOR U22656 ( .A(n21631), .B(n10818), .Z(n21634) );
  XNOR U22657 ( .A(n21627), .B(n21629), .Z(n10818) );
  NAND U22658 ( .A(n21635), .B(e_input[247]), .Z(n21629) );
  NAND U22659 ( .A(n12323), .B(e_input[247]), .Z(n21635) );
  XNOR U22660 ( .A(n21625), .B(n21636), .Z(n21627) );
  XOR U22661 ( .A(n21637), .B(n21638), .Z(n21625) );
  AND U22662 ( .A(n21639), .B(n21640), .Z(n21638) );
  XNOR U22663 ( .A(n21641), .B(n21637), .Z(n21640) );
  XOR U22664 ( .A(n21642), .B(e_input[247]), .Z(n21633) );
  IV U22665 ( .A(n21631), .Z(n21642) );
  XOR U22666 ( .A(n21643), .B(n21644), .Z(n21631) );
  AND U22667 ( .A(n21645), .B(n21646), .Z(n21644) );
  XNOR U22668 ( .A(n21643), .B(n10824), .Z(n21646) );
  XNOR U22669 ( .A(n21639), .B(n21641), .Z(n10824) );
  NAND U22670 ( .A(n21647), .B(e_input[246]), .Z(n21641) );
  NAND U22671 ( .A(n12323), .B(e_input[246]), .Z(n21647) );
  XNOR U22672 ( .A(n21637), .B(n21648), .Z(n21639) );
  XOR U22673 ( .A(n21649), .B(n21650), .Z(n21637) );
  AND U22674 ( .A(n21651), .B(n21652), .Z(n21650) );
  XNOR U22675 ( .A(n21653), .B(n21649), .Z(n21652) );
  XOR U22676 ( .A(n21654), .B(e_input[246]), .Z(n21645) );
  IV U22677 ( .A(n21643), .Z(n21654) );
  XOR U22678 ( .A(n21655), .B(n21656), .Z(n21643) );
  AND U22679 ( .A(n21657), .B(n21658), .Z(n21656) );
  XNOR U22680 ( .A(n21655), .B(n10830), .Z(n21658) );
  XNOR U22681 ( .A(n21651), .B(n21653), .Z(n10830) );
  NAND U22682 ( .A(n21659), .B(e_input[245]), .Z(n21653) );
  NAND U22683 ( .A(n12323), .B(e_input[245]), .Z(n21659) );
  XNOR U22684 ( .A(n21649), .B(n21660), .Z(n21651) );
  XOR U22685 ( .A(n21661), .B(n21662), .Z(n21649) );
  AND U22686 ( .A(n21663), .B(n21664), .Z(n21662) );
  XNOR U22687 ( .A(n21665), .B(n21661), .Z(n21664) );
  XOR U22688 ( .A(n21666), .B(e_input[245]), .Z(n21657) );
  IV U22689 ( .A(n21655), .Z(n21666) );
  XOR U22690 ( .A(n21667), .B(n21668), .Z(n21655) );
  AND U22691 ( .A(n21669), .B(n21670), .Z(n21668) );
  XNOR U22692 ( .A(n21667), .B(n10836), .Z(n21670) );
  XNOR U22693 ( .A(n21663), .B(n21665), .Z(n10836) );
  NAND U22694 ( .A(n21671), .B(e_input[244]), .Z(n21665) );
  NAND U22695 ( .A(n12323), .B(e_input[244]), .Z(n21671) );
  XNOR U22696 ( .A(n21661), .B(n21672), .Z(n21663) );
  XOR U22697 ( .A(n21673), .B(n21674), .Z(n21661) );
  AND U22698 ( .A(n21675), .B(n21676), .Z(n21674) );
  XNOR U22699 ( .A(n21677), .B(n21673), .Z(n21676) );
  XOR U22700 ( .A(n21678), .B(e_input[244]), .Z(n21669) );
  IV U22701 ( .A(n21667), .Z(n21678) );
  XOR U22702 ( .A(n21679), .B(n21680), .Z(n21667) );
  AND U22703 ( .A(n21681), .B(n21682), .Z(n21680) );
  XNOR U22704 ( .A(n21679), .B(n10842), .Z(n21682) );
  XNOR U22705 ( .A(n21675), .B(n21677), .Z(n10842) );
  NAND U22706 ( .A(n21683), .B(e_input[243]), .Z(n21677) );
  NAND U22707 ( .A(n12323), .B(e_input[243]), .Z(n21683) );
  XNOR U22708 ( .A(n21673), .B(n21684), .Z(n21675) );
  XOR U22709 ( .A(n21685), .B(n21686), .Z(n21673) );
  AND U22710 ( .A(n21687), .B(n21688), .Z(n21686) );
  XNOR U22711 ( .A(n21689), .B(n21685), .Z(n21688) );
  XOR U22712 ( .A(n21690), .B(e_input[243]), .Z(n21681) );
  IV U22713 ( .A(n21679), .Z(n21690) );
  XOR U22714 ( .A(n21691), .B(n21692), .Z(n21679) );
  AND U22715 ( .A(n21693), .B(n21694), .Z(n21692) );
  XNOR U22716 ( .A(n21691), .B(n10848), .Z(n21694) );
  XNOR U22717 ( .A(n21687), .B(n21689), .Z(n10848) );
  NAND U22718 ( .A(n21695), .B(e_input[242]), .Z(n21689) );
  NAND U22719 ( .A(n12323), .B(e_input[242]), .Z(n21695) );
  XNOR U22720 ( .A(n21685), .B(n21696), .Z(n21687) );
  XOR U22721 ( .A(n21697), .B(n21698), .Z(n21685) );
  AND U22722 ( .A(n21699), .B(n21700), .Z(n21698) );
  XNOR U22723 ( .A(n21701), .B(n21697), .Z(n21700) );
  XOR U22724 ( .A(n21702), .B(e_input[242]), .Z(n21693) );
  IV U22725 ( .A(n21691), .Z(n21702) );
  XOR U22726 ( .A(n21703), .B(n21704), .Z(n21691) );
  AND U22727 ( .A(n21705), .B(n21706), .Z(n21704) );
  XNOR U22728 ( .A(n21703), .B(n10854), .Z(n21706) );
  XNOR U22729 ( .A(n21699), .B(n21701), .Z(n10854) );
  NAND U22730 ( .A(n21707), .B(e_input[241]), .Z(n21701) );
  NAND U22731 ( .A(n12323), .B(e_input[241]), .Z(n21707) );
  XNOR U22732 ( .A(n21697), .B(n21708), .Z(n21699) );
  XOR U22733 ( .A(n21709), .B(n21710), .Z(n21697) );
  AND U22734 ( .A(n21711), .B(n21712), .Z(n21710) );
  XNOR U22735 ( .A(n21713), .B(n21709), .Z(n21712) );
  XOR U22736 ( .A(n21714), .B(e_input[241]), .Z(n21705) );
  IV U22737 ( .A(n21703), .Z(n21714) );
  XOR U22738 ( .A(n21715), .B(n21716), .Z(n21703) );
  AND U22739 ( .A(n21717), .B(n21718), .Z(n21716) );
  XNOR U22740 ( .A(n21715), .B(n10860), .Z(n21718) );
  XNOR U22741 ( .A(n21711), .B(n21713), .Z(n10860) );
  NAND U22742 ( .A(n21719), .B(e_input[240]), .Z(n21713) );
  NAND U22743 ( .A(n12323), .B(e_input[240]), .Z(n21719) );
  XNOR U22744 ( .A(n21709), .B(n21720), .Z(n21711) );
  XOR U22745 ( .A(n21721), .B(n21722), .Z(n21709) );
  AND U22746 ( .A(n21723), .B(n21724), .Z(n21722) );
  XNOR U22747 ( .A(n21725), .B(n21721), .Z(n21724) );
  XOR U22748 ( .A(n21726), .B(e_input[240]), .Z(n21717) );
  IV U22749 ( .A(n21715), .Z(n21726) );
  XOR U22750 ( .A(n21727), .B(n21728), .Z(n21715) );
  AND U22751 ( .A(n21729), .B(n21730), .Z(n21728) );
  XNOR U22752 ( .A(n21727), .B(n10866), .Z(n21730) );
  XNOR U22753 ( .A(n21723), .B(n21725), .Z(n10866) );
  NAND U22754 ( .A(n21731), .B(e_input[239]), .Z(n21725) );
  NAND U22755 ( .A(n12323), .B(e_input[239]), .Z(n21731) );
  XNOR U22756 ( .A(n21721), .B(n21732), .Z(n21723) );
  XOR U22757 ( .A(n21733), .B(n21734), .Z(n21721) );
  AND U22758 ( .A(n21735), .B(n21736), .Z(n21734) );
  XNOR U22759 ( .A(n21737), .B(n21733), .Z(n21736) );
  XOR U22760 ( .A(n21738), .B(e_input[239]), .Z(n21729) );
  IV U22761 ( .A(n21727), .Z(n21738) );
  XOR U22762 ( .A(n21739), .B(n21740), .Z(n21727) );
  AND U22763 ( .A(n21741), .B(n21742), .Z(n21740) );
  XNOR U22764 ( .A(n21739), .B(n10872), .Z(n21742) );
  XNOR U22765 ( .A(n21735), .B(n21737), .Z(n10872) );
  NAND U22766 ( .A(n21743), .B(e_input[238]), .Z(n21737) );
  NAND U22767 ( .A(n12323), .B(e_input[238]), .Z(n21743) );
  XNOR U22768 ( .A(n21733), .B(n21744), .Z(n21735) );
  XOR U22769 ( .A(n21745), .B(n21746), .Z(n21733) );
  AND U22770 ( .A(n21747), .B(n21748), .Z(n21746) );
  XNOR U22771 ( .A(n21749), .B(n21745), .Z(n21748) );
  XOR U22772 ( .A(n21750), .B(e_input[238]), .Z(n21741) );
  IV U22773 ( .A(n21739), .Z(n21750) );
  XOR U22774 ( .A(n21751), .B(n21752), .Z(n21739) );
  AND U22775 ( .A(n21753), .B(n21754), .Z(n21752) );
  XNOR U22776 ( .A(n21751), .B(n10878), .Z(n21754) );
  XNOR U22777 ( .A(n21747), .B(n21749), .Z(n10878) );
  NAND U22778 ( .A(n21755), .B(e_input[237]), .Z(n21749) );
  NAND U22779 ( .A(n12323), .B(e_input[237]), .Z(n21755) );
  XNOR U22780 ( .A(n21745), .B(n21756), .Z(n21747) );
  XOR U22781 ( .A(n21757), .B(n21758), .Z(n21745) );
  AND U22782 ( .A(n21759), .B(n21760), .Z(n21758) );
  XNOR U22783 ( .A(n21761), .B(n21757), .Z(n21760) );
  XOR U22784 ( .A(n21762), .B(e_input[237]), .Z(n21753) );
  IV U22785 ( .A(n21751), .Z(n21762) );
  XOR U22786 ( .A(n21763), .B(n21764), .Z(n21751) );
  AND U22787 ( .A(n21765), .B(n21766), .Z(n21764) );
  XNOR U22788 ( .A(n21763), .B(n10884), .Z(n21766) );
  XNOR U22789 ( .A(n21759), .B(n21761), .Z(n10884) );
  NAND U22790 ( .A(n21767), .B(e_input[236]), .Z(n21761) );
  NAND U22791 ( .A(n12323), .B(e_input[236]), .Z(n21767) );
  XNOR U22792 ( .A(n21757), .B(n21768), .Z(n21759) );
  XOR U22793 ( .A(n21769), .B(n21770), .Z(n21757) );
  AND U22794 ( .A(n21771), .B(n21772), .Z(n21770) );
  XNOR U22795 ( .A(n21773), .B(n21769), .Z(n21772) );
  XOR U22796 ( .A(n21774), .B(e_input[236]), .Z(n21765) );
  IV U22797 ( .A(n21763), .Z(n21774) );
  XOR U22798 ( .A(n21775), .B(n21776), .Z(n21763) );
  AND U22799 ( .A(n21777), .B(n21778), .Z(n21776) );
  XNOR U22800 ( .A(n21775), .B(n10890), .Z(n21778) );
  XNOR U22801 ( .A(n21771), .B(n21773), .Z(n10890) );
  NAND U22802 ( .A(n21779), .B(e_input[235]), .Z(n21773) );
  NAND U22803 ( .A(n12323), .B(e_input[235]), .Z(n21779) );
  XNOR U22804 ( .A(n21769), .B(n21780), .Z(n21771) );
  XOR U22805 ( .A(n21781), .B(n21782), .Z(n21769) );
  AND U22806 ( .A(n21783), .B(n21784), .Z(n21782) );
  XNOR U22807 ( .A(n21785), .B(n21781), .Z(n21784) );
  XOR U22808 ( .A(n21786), .B(e_input[235]), .Z(n21777) );
  IV U22809 ( .A(n21775), .Z(n21786) );
  XOR U22810 ( .A(n21787), .B(n21788), .Z(n21775) );
  AND U22811 ( .A(n21789), .B(n21790), .Z(n21788) );
  XNOR U22812 ( .A(n21787), .B(n10896), .Z(n21790) );
  XNOR U22813 ( .A(n21783), .B(n21785), .Z(n10896) );
  NAND U22814 ( .A(n21791), .B(e_input[234]), .Z(n21785) );
  NAND U22815 ( .A(n12323), .B(e_input[234]), .Z(n21791) );
  XNOR U22816 ( .A(n21781), .B(n21792), .Z(n21783) );
  XOR U22817 ( .A(n21793), .B(n21794), .Z(n21781) );
  AND U22818 ( .A(n21795), .B(n21796), .Z(n21794) );
  XNOR U22819 ( .A(n21797), .B(n21793), .Z(n21796) );
  XOR U22820 ( .A(n21798), .B(e_input[234]), .Z(n21789) );
  IV U22821 ( .A(n21787), .Z(n21798) );
  XOR U22822 ( .A(n21799), .B(n21800), .Z(n21787) );
  AND U22823 ( .A(n21801), .B(n21802), .Z(n21800) );
  XNOR U22824 ( .A(n21799), .B(n10902), .Z(n21802) );
  XNOR U22825 ( .A(n21795), .B(n21797), .Z(n10902) );
  NAND U22826 ( .A(n21803), .B(e_input[233]), .Z(n21797) );
  NAND U22827 ( .A(n12323), .B(e_input[233]), .Z(n21803) );
  XNOR U22828 ( .A(n21793), .B(n21804), .Z(n21795) );
  XOR U22829 ( .A(n21805), .B(n21806), .Z(n21793) );
  AND U22830 ( .A(n21807), .B(n21808), .Z(n21806) );
  XNOR U22831 ( .A(n21809), .B(n21805), .Z(n21808) );
  XOR U22832 ( .A(n21810), .B(e_input[233]), .Z(n21801) );
  IV U22833 ( .A(n21799), .Z(n21810) );
  XOR U22834 ( .A(n21811), .B(n21812), .Z(n21799) );
  AND U22835 ( .A(n21813), .B(n21814), .Z(n21812) );
  XNOR U22836 ( .A(n21811), .B(n10908), .Z(n21814) );
  XNOR U22837 ( .A(n21807), .B(n21809), .Z(n10908) );
  NAND U22838 ( .A(n21815), .B(e_input[232]), .Z(n21809) );
  NAND U22839 ( .A(n12323), .B(e_input[232]), .Z(n21815) );
  XNOR U22840 ( .A(n21805), .B(n21816), .Z(n21807) );
  XOR U22841 ( .A(n21817), .B(n21818), .Z(n21805) );
  AND U22842 ( .A(n21819), .B(n21820), .Z(n21818) );
  XNOR U22843 ( .A(n21821), .B(n21817), .Z(n21820) );
  XOR U22844 ( .A(n21822), .B(e_input[232]), .Z(n21813) );
  IV U22845 ( .A(n21811), .Z(n21822) );
  XOR U22846 ( .A(n21823), .B(n21824), .Z(n21811) );
  AND U22847 ( .A(n21825), .B(n21826), .Z(n21824) );
  XNOR U22848 ( .A(n21823), .B(n10914), .Z(n21826) );
  XNOR U22849 ( .A(n21819), .B(n21821), .Z(n10914) );
  NAND U22850 ( .A(n21827), .B(e_input[231]), .Z(n21821) );
  NAND U22851 ( .A(n12323), .B(e_input[231]), .Z(n21827) );
  XNOR U22852 ( .A(n21817), .B(n21828), .Z(n21819) );
  XOR U22853 ( .A(n21829), .B(n21830), .Z(n21817) );
  AND U22854 ( .A(n21831), .B(n21832), .Z(n21830) );
  XNOR U22855 ( .A(n21833), .B(n21829), .Z(n21832) );
  XOR U22856 ( .A(n21834), .B(e_input[231]), .Z(n21825) );
  IV U22857 ( .A(n21823), .Z(n21834) );
  XOR U22858 ( .A(n21835), .B(n21836), .Z(n21823) );
  AND U22859 ( .A(n21837), .B(n21838), .Z(n21836) );
  XNOR U22860 ( .A(n21835), .B(n10920), .Z(n21838) );
  XNOR U22861 ( .A(n21831), .B(n21833), .Z(n10920) );
  NAND U22862 ( .A(n21839), .B(e_input[230]), .Z(n21833) );
  NAND U22863 ( .A(n12323), .B(e_input[230]), .Z(n21839) );
  XNOR U22864 ( .A(n21829), .B(n21840), .Z(n21831) );
  XOR U22865 ( .A(n21841), .B(n21842), .Z(n21829) );
  AND U22866 ( .A(n21843), .B(n21844), .Z(n21842) );
  XNOR U22867 ( .A(n21845), .B(n21841), .Z(n21844) );
  XOR U22868 ( .A(n21846), .B(e_input[230]), .Z(n21837) );
  IV U22869 ( .A(n21835), .Z(n21846) );
  XOR U22870 ( .A(n21847), .B(n21848), .Z(n21835) );
  AND U22871 ( .A(n21849), .B(n21850), .Z(n21848) );
  XNOR U22872 ( .A(n21847), .B(n10926), .Z(n21850) );
  XNOR U22873 ( .A(n21843), .B(n21845), .Z(n10926) );
  NAND U22874 ( .A(n21851), .B(e_input[229]), .Z(n21845) );
  NAND U22875 ( .A(n12323), .B(e_input[229]), .Z(n21851) );
  XNOR U22876 ( .A(n21841), .B(n21852), .Z(n21843) );
  XOR U22877 ( .A(n21853), .B(n21854), .Z(n21841) );
  AND U22878 ( .A(n21855), .B(n21856), .Z(n21854) );
  XNOR U22879 ( .A(n21857), .B(n21853), .Z(n21856) );
  XOR U22880 ( .A(n21858), .B(e_input[229]), .Z(n21849) );
  IV U22881 ( .A(n21847), .Z(n21858) );
  XOR U22882 ( .A(n21859), .B(n21860), .Z(n21847) );
  AND U22883 ( .A(n21861), .B(n21862), .Z(n21860) );
  XNOR U22884 ( .A(n21859), .B(n10932), .Z(n21862) );
  XNOR U22885 ( .A(n21855), .B(n21857), .Z(n10932) );
  NAND U22886 ( .A(n21863), .B(e_input[228]), .Z(n21857) );
  NAND U22887 ( .A(n12323), .B(e_input[228]), .Z(n21863) );
  XNOR U22888 ( .A(n21853), .B(n21864), .Z(n21855) );
  XOR U22889 ( .A(n21865), .B(n21866), .Z(n21853) );
  AND U22890 ( .A(n21867), .B(n21868), .Z(n21866) );
  XNOR U22891 ( .A(n21869), .B(n21865), .Z(n21868) );
  XOR U22892 ( .A(n21870), .B(e_input[228]), .Z(n21861) );
  IV U22893 ( .A(n21859), .Z(n21870) );
  XOR U22894 ( .A(n21871), .B(n21872), .Z(n21859) );
  AND U22895 ( .A(n21873), .B(n21874), .Z(n21872) );
  XNOR U22896 ( .A(n21871), .B(n10938), .Z(n21874) );
  XNOR U22897 ( .A(n21867), .B(n21869), .Z(n10938) );
  NAND U22898 ( .A(n21875), .B(e_input[227]), .Z(n21869) );
  NAND U22899 ( .A(n12323), .B(e_input[227]), .Z(n21875) );
  XNOR U22900 ( .A(n21865), .B(n21876), .Z(n21867) );
  XOR U22901 ( .A(n21877), .B(n21878), .Z(n21865) );
  AND U22902 ( .A(n21879), .B(n21880), .Z(n21878) );
  XNOR U22903 ( .A(n21881), .B(n21877), .Z(n21880) );
  XOR U22904 ( .A(n21882), .B(e_input[227]), .Z(n21873) );
  IV U22905 ( .A(n21871), .Z(n21882) );
  XOR U22906 ( .A(n21883), .B(n21884), .Z(n21871) );
  AND U22907 ( .A(n21885), .B(n21886), .Z(n21884) );
  XNOR U22908 ( .A(n21883), .B(n10944), .Z(n21886) );
  XNOR U22909 ( .A(n21879), .B(n21881), .Z(n10944) );
  NAND U22910 ( .A(n21887), .B(e_input[226]), .Z(n21881) );
  NAND U22911 ( .A(n12323), .B(e_input[226]), .Z(n21887) );
  XNOR U22912 ( .A(n21877), .B(n21888), .Z(n21879) );
  XOR U22913 ( .A(n21889), .B(n21890), .Z(n21877) );
  AND U22914 ( .A(n21891), .B(n21892), .Z(n21890) );
  XNOR U22915 ( .A(n21893), .B(n21889), .Z(n21892) );
  XOR U22916 ( .A(n21894), .B(e_input[226]), .Z(n21885) );
  IV U22917 ( .A(n21883), .Z(n21894) );
  XOR U22918 ( .A(n21895), .B(n21896), .Z(n21883) );
  AND U22919 ( .A(n21897), .B(n21898), .Z(n21896) );
  XNOR U22920 ( .A(n21895), .B(n10950), .Z(n21898) );
  XNOR U22921 ( .A(n21891), .B(n21893), .Z(n10950) );
  NAND U22922 ( .A(n21899), .B(e_input[225]), .Z(n21893) );
  NAND U22923 ( .A(n12323), .B(e_input[225]), .Z(n21899) );
  XNOR U22924 ( .A(n21889), .B(n21900), .Z(n21891) );
  XOR U22925 ( .A(n21901), .B(n21902), .Z(n21889) );
  AND U22926 ( .A(n21903), .B(n21904), .Z(n21902) );
  XNOR U22927 ( .A(n21905), .B(n21901), .Z(n21904) );
  XOR U22928 ( .A(n21906), .B(e_input[225]), .Z(n21897) );
  IV U22929 ( .A(n21895), .Z(n21906) );
  XOR U22930 ( .A(n21907), .B(n21908), .Z(n21895) );
  AND U22931 ( .A(n21909), .B(n21910), .Z(n21908) );
  XNOR U22932 ( .A(n21907), .B(n10956), .Z(n21910) );
  XNOR U22933 ( .A(n21903), .B(n21905), .Z(n10956) );
  NAND U22934 ( .A(n21911), .B(e_input[224]), .Z(n21905) );
  NAND U22935 ( .A(n12323), .B(e_input[224]), .Z(n21911) );
  XNOR U22936 ( .A(n21901), .B(n21912), .Z(n21903) );
  XOR U22937 ( .A(n21913), .B(n21914), .Z(n21901) );
  AND U22938 ( .A(n21915), .B(n21916), .Z(n21914) );
  XNOR U22939 ( .A(n21917), .B(n21913), .Z(n21916) );
  XOR U22940 ( .A(n21918), .B(e_input[224]), .Z(n21909) );
  IV U22941 ( .A(n21907), .Z(n21918) );
  XOR U22942 ( .A(n21919), .B(n21920), .Z(n21907) );
  AND U22943 ( .A(n21921), .B(n21922), .Z(n21920) );
  XNOR U22944 ( .A(n21919), .B(n10962), .Z(n21922) );
  XNOR U22945 ( .A(n21915), .B(n21917), .Z(n10962) );
  NAND U22946 ( .A(n21923), .B(e_input[223]), .Z(n21917) );
  NAND U22947 ( .A(n12323), .B(e_input[223]), .Z(n21923) );
  XNOR U22948 ( .A(n21913), .B(n21924), .Z(n21915) );
  XOR U22949 ( .A(n21925), .B(n21926), .Z(n21913) );
  AND U22950 ( .A(n21927), .B(n21928), .Z(n21926) );
  XNOR U22951 ( .A(n21929), .B(n21925), .Z(n21928) );
  XOR U22952 ( .A(n21930), .B(e_input[223]), .Z(n21921) );
  IV U22953 ( .A(n21919), .Z(n21930) );
  XOR U22954 ( .A(n21931), .B(n21932), .Z(n21919) );
  AND U22955 ( .A(n21933), .B(n21934), .Z(n21932) );
  XNOR U22956 ( .A(n21931), .B(n10968), .Z(n21934) );
  XNOR U22957 ( .A(n21927), .B(n21929), .Z(n10968) );
  NAND U22958 ( .A(n21935), .B(e_input[222]), .Z(n21929) );
  NAND U22959 ( .A(n12323), .B(e_input[222]), .Z(n21935) );
  XNOR U22960 ( .A(n21925), .B(n21936), .Z(n21927) );
  XOR U22961 ( .A(n21937), .B(n21938), .Z(n21925) );
  AND U22962 ( .A(n21939), .B(n21940), .Z(n21938) );
  XNOR U22963 ( .A(n21941), .B(n21937), .Z(n21940) );
  XOR U22964 ( .A(n21942), .B(e_input[222]), .Z(n21933) );
  IV U22965 ( .A(n21931), .Z(n21942) );
  XOR U22966 ( .A(n21943), .B(n21944), .Z(n21931) );
  AND U22967 ( .A(n21945), .B(n21946), .Z(n21944) );
  XNOR U22968 ( .A(n21943), .B(n10974), .Z(n21946) );
  XNOR U22969 ( .A(n21939), .B(n21941), .Z(n10974) );
  NAND U22970 ( .A(n21947), .B(e_input[221]), .Z(n21941) );
  NAND U22971 ( .A(n12323), .B(e_input[221]), .Z(n21947) );
  XNOR U22972 ( .A(n21937), .B(n21948), .Z(n21939) );
  XOR U22973 ( .A(n21949), .B(n21950), .Z(n21937) );
  AND U22974 ( .A(n21951), .B(n21952), .Z(n21950) );
  XNOR U22975 ( .A(n21953), .B(n21949), .Z(n21952) );
  XOR U22976 ( .A(n21954), .B(e_input[221]), .Z(n21945) );
  IV U22977 ( .A(n21943), .Z(n21954) );
  XOR U22978 ( .A(n21955), .B(n21956), .Z(n21943) );
  AND U22979 ( .A(n21957), .B(n21958), .Z(n21956) );
  XNOR U22980 ( .A(n21955), .B(n10980), .Z(n21958) );
  XNOR U22981 ( .A(n21951), .B(n21953), .Z(n10980) );
  NAND U22982 ( .A(n21959), .B(e_input[220]), .Z(n21953) );
  NAND U22983 ( .A(n12323), .B(e_input[220]), .Z(n21959) );
  XNOR U22984 ( .A(n21949), .B(n21960), .Z(n21951) );
  XOR U22985 ( .A(n21961), .B(n21962), .Z(n21949) );
  AND U22986 ( .A(n21963), .B(n21964), .Z(n21962) );
  XNOR U22987 ( .A(n21965), .B(n21961), .Z(n21964) );
  XOR U22988 ( .A(n21966), .B(e_input[220]), .Z(n21957) );
  IV U22989 ( .A(n21955), .Z(n21966) );
  XOR U22990 ( .A(n21967), .B(n21968), .Z(n21955) );
  AND U22991 ( .A(n21969), .B(n21970), .Z(n21968) );
  XNOR U22992 ( .A(n21967), .B(n10986), .Z(n21970) );
  XNOR U22993 ( .A(n21963), .B(n21965), .Z(n10986) );
  NAND U22994 ( .A(n21971), .B(e_input[219]), .Z(n21965) );
  NAND U22995 ( .A(n12323), .B(e_input[219]), .Z(n21971) );
  XNOR U22996 ( .A(n21961), .B(n21972), .Z(n21963) );
  XOR U22997 ( .A(n21973), .B(n21974), .Z(n21961) );
  AND U22998 ( .A(n21975), .B(n21976), .Z(n21974) );
  XNOR U22999 ( .A(n21977), .B(n21973), .Z(n21976) );
  XOR U23000 ( .A(n21978), .B(e_input[219]), .Z(n21969) );
  IV U23001 ( .A(n21967), .Z(n21978) );
  XOR U23002 ( .A(n21979), .B(n21980), .Z(n21967) );
  AND U23003 ( .A(n21981), .B(n21982), .Z(n21980) );
  XNOR U23004 ( .A(n21979), .B(n10992), .Z(n21982) );
  XNOR U23005 ( .A(n21975), .B(n21977), .Z(n10992) );
  NAND U23006 ( .A(n21983), .B(e_input[218]), .Z(n21977) );
  NAND U23007 ( .A(n12323), .B(e_input[218]), .Z(n21983) );
  XNOR U23008 ( .A(n21973), .B(n21984), .Z(n21975) );
  XOR U23009 ( .A(n21985), .B(n21986), .Z(n21973) );
  AND U23010 ( .A(n21987), .B(n21988), .Z(n21986) );
  XNOR U23011 ( .A(n21989), .B(n21985), .Z(n21988) );
  XOR U23012 ( .A(n21990), .B(e_input[218]), .Z(n21981) );
  IV U23013 ( .A(n21979), .Z(n21990) );
  XOR U23014 ( .A(n21991), .B(n21992), .Z(n21979) );
  AND U23015 ( .A(n21993), .B(n21994), .Z(n21992) );
  XNOR U23016 ( .A(n21991), .B(n10998), .Z(n21994) );
  XNOR U23017 ( .A(n21987), .B(n21989), .Z(n10998) );
  NAND U23018 ( .A(n21995), .B(e_input[217]), .Z(n21989) );
  NAND U23019 ( .A(n12323), .B(e_input[217]), .Z(n21995) );
  XNOR U23020 ( .A(n21985), .B(n21996), .Z(n21987) );
  XOR U23021 ( .A(n21997), .B(n21998), .Z(n21985) );
  AND U23022 ( .A(n21999), .B(n22000), .Z(n21998) );
  XNOR U23023 ( .A(n22001), .B(n21997), .Z(n22000) );
  XOR U23024 ( .A(n22002), .B(e_input[217]), .Z(n21993) );
  IV U23025 ( .A(n21991), .Z(n22002) );
  XOR U23026 ( .A(n22003), .B(n22004), .Z(n21991) );
  AND U23027 ( .A(n22005), .B(n22006), .Z(n22004) );
  XNOR U23028 ( .A(n22003), .B(n11004), .Z(n22006) );
  XNOR U23029 ( .A(n21999), .B(n22001), .Z(n11004) );
  NAND U23030 ( .A(n22007), .B(e_input[216]), .Z(n22001) );
  NAND U23031 ( .A(n12323), .B(e_input[216]), .Z(n22007) );
  XNOR U23032 ( .A(n21997), .B(n22008), .Z(n21999) );
  XOR U23033 ( .A(n22009), .B(n22010), .Z(n21997) );
  AND U23034 ( .A(n22011), .B(n22012), .Z(n22010) );
  XNOR U23035 ( .A(n22013), .B(n22009), .Z(n22012) );
  XOR U23036 ( .A(n22014), .B(e_input[216]), .Z(n22005) );
  IV U23037 ( .A(n22003), .Z(n22014) );
  XOR U23038 ( .A(n22015), .B(n22016), .Z(n22003) );
  AND U23039 ( .A(n22017), .B(n22018), .Z(n22016) );
  XNOR U23040 ( .A(n22015), .B(n11010), .Z(n22018) );
  XNOR U23041 ( .A(n22011), .B(n22013), .Z(n11010) );
  NAND U23042 ( .A(n22019), .B(e_input[215]), .Z(n22013) );
  NAND U23043 ( .A(n12323), .B(e_input[215]), .Z(n22019) );
  XNOR U23044 ( .A(n22009), .B(n22020), .Z(n22011) );
  XOR U23045 ( .A(n22021), .B(n22022), .Z(n22009) );
  AND U23046 ( .A(n22023), .B(n22024), .Z(n22022) );
  XNOR U23047 ( .A(n22025), .B(n22021), .Z(n22024) );
  XOR U23048 ( .A(n22026), .B(e_input[215]), .Z(n22017) );
  IV U23049 ( .A(n22015), .Z(n22026) );
  XOR U23050 ( .A(n22027), .B(n22028), .Z(n22015) );
  AND U23051 ( .A(n22029), .B(n22030), .Z(n22028) );
  XNOR U23052 ( .A(n22027), .B(n11016), .Z(n22030) );
  XNOR U23053 ( .A(n22023), .B(n22025), .Z(n11016) );
  NAND U23054 ( .A(n22031), .B(e_input[214]), .Z(n22025) );
  NAND U23055 ( .A(n12323), .B(e_input[214]), .Z(n22031) );
  XNOR U23056 ( .A(n22021), .B(n22032), .Z(n22023) );
  XOR U23057 ( .A(n22033), .B(n22034), .Z(n22021) );
  AND U23058 ( .A(n22035), .B(n22036), .Z(n22034) );
  XNOR U23059 ( .A(n22037), .B(n22033), .Z(n22036) );
  XOR U23060 ( .A(n22038), .B(e_input[214]), .Z(n22029) );
  IV U23061 ( .A(n22027), .Z(n22038) );
  XOR U23062 ( .A(n22039), .B(n22040), .Z(n22027) );
  AND U23063 ( .A(n22041), .B(n22042), .Z(n22040) );
  XNOR U23064 ( .A(n22039), .B(n11022), .Z(n22042) );
  XNOR U23065 ( .A(n22035), .B(n22037), .Z(n11022) );
  NAND U23066 ( .A(n22043), .B(e_input[213]), .Z(n22037) );
  NAND U23067 ( .A(n12323), .B(e_input[213]), .Z(n22043) );
  XNOR U23068 ( .A(n22033), .B(n22044), .Z(n22035) );
  XOR U23069 ( .A(n22045), .B(n22046), .Z(n22033) );
  AND U23070 ( .A(n22047), .B(n22048), .Z(n22046) );
  XNOR U23071 ( .A(n22049), .B(n22045), .Z(n22048) );
  XOR U23072 ( .A(n22050), .B(e_input[213]), .Z(n22041) );
  IV U23073 ( .A(n22039), .Z(n22050) );
  XOR U23074 ( .A(n22051), .B(n22052), .Z(n22039) );
  AND U23075 ( .A(n22053), .B(n22054), .Z(n22052) );
  XNOR U23076 ( .A(n22051), .B(n11028), .Z(n22054) );
  XNOR U23077 ( .A(n22047), .B(n22049), .Z(n11028) );
  NAND U23078 ( .A(n22055), .B(e_input[212]), .Z(n22049) );
  NAND U23079 ( .A(n12323), .B(e_input[212]), .Z(n22055) );
  XNOR U23080 ( .A(n22045), .B(n22056), .Z(n22047) );
  XOR U23081 ( .A(n22057), .B(n22058), .Z(n22045) );
  AND U23082 ( .A(n22059), .B(n22060), .Z(n22058) );
  XNOR U23083 ( .A(n22061), .B(n22057), .Z(n22060) );
  XOR U23084 ( .A(n22062), .B(e_input[212]), .Z(n22053) );
  IV U23085 ( .A(n22051), .Z(n22062) );
  XOR U23086 ( .A(n22063), .B(n22064), .Z(n22051) );
  AND U23087 ( .A(n22065), .B(n22066), .Z(n22064) );
  XNOR U23088 ( .A(n22063), .B(n11034), .Z(n22066) );
  XNOR U23089 ( .A(n22059), .B(n22061), .Z(n11034) );
  NAND U23090 ( .A(n22067), .B(e_input[211]), .Z(n22061) );
  NAND U23091 ( .A(n12323), .B(e_input[211]), .Z(n22067) );
  XNOR U23092 ( .A(n22057), .B(n22068), .Z(n22059) );
  XOR U23093 ( .A(n22069), .B(n22070), .Z(n22057) );
  AND U23094 ( .A(n22071), .B(n22072), .Z(n22070) );
  XNOR U23095 ( .A(n22073), .B(n22069), .Z(n22072) );
  XOR U23096 ( .A(n22074), .B(e_input[211]), .Z(n22065) );
  IV U23097 ( .A(n22063), .Z(n22074) );
  XOR U23098 ( .A(n22075), .B(n22076), .Z(n22063) );
  AND U23099 ( .A(n22077), .B(n22078), .Z(n22076) );
  XNOR U23100 ( .A(n22075), .B(n11040), .Z(n22078) );
  XNOR U23101 ( .A(n22071), .B(n22073), .Z(n11040) );
  NAND U23102 ( .A(n22079), .B(e_input[210]), .Z(n22073) );
  NAND U23103 ( .A(n12323), .B(e_input[210]), .Z(n22079) );
  XNOR U23104 ( .A(n22069), .B(n22080), .Z(n22071) );
  XOR U23105 ( .A(n22081), .B(n22082), .Z(n22069) );
  AND U23106 ( .A(n22083), .B(n22084), .Z(n22082) );
  XNOR U23107 ( .A(n22085), .B(n22081), .Z(n22084) );
  XOR U23108 ( .A(n22086), .B(e_input[210]), .Z(n22077) );
  IV U23109 ( .A(n22075), .Z(n22086) );
  XOR U23110 ( .A(n22087), .B(n22088), .Z(n22075) );
  AND U23111 ( .A(n22089), .B(n22090), .Z(n22088) );
  XNOR U23112 ( .A(n22087), .B(n11046), .Z(n22090) );
  XNOR U23113 ( .A(n22083), .B(n22085), .Z(n11046) );
  NAND U23114 ( .A(n22091), .B(e_input[209]), .Z(n22085) );
  NAND U23115 ( .A(n12323), .B(e_input[209]), .Z(n22091) );
  XNOR U23116 ( .A(n22081), .B(n22092), .Z(n22083) );
  XOR U23117 ( .A(n22093), .B(n22094), .Z(n22081) );
  AND U23118 ( .A(n22095), .B(n22096), .Z(n22094) );
  XNOR U23119 ( .A(n22097), .B(n22093), .Z(n22096) );
  XOR U23120 ( .A(n22098), .B(e_input[209]), .Z(n22089) );
  IV U23121 ( .A(n22087), .Z(n22098) );
  XOR U23122 ( .A(n22099), .B(n22100), .Z(n22087) );
  AND U23123 ( .A(n22101), .B(n22102), .Z(n22100) );
  XNOR U23124 ( .A(n22099), .B(n11052), .Z(n22102) );
  XNOR U23125 ( .A(n22095), .B(n22097), .Z(n11052) );
  NAND U23126 ( .A(n22103), .B(e_input[208]), .Z(n22097) );
  NAND U23127 ( .A(n12323), .B(e_input[208]), .Z(n22103) );
  XNOR U23128 ( .A(n22093), .B(n22104), .Z(n22095) );
  XOR U23129 ( .A(n22105), .B(n22106), .Z(n22093) );
  AND U23130 ( .A(n22107), .B(n22108), .Z(n22106) );
  XNOR U23131 ( .A(n22109), .B(n22105), .Z(n22108) );
  XOR U23132 ( .A(n22110), .B(e_input[208]), .Z(n22101) );
  IV U23133 ( .A(n22099), .Z(n22110) );
  XOR U23134 ( .A(n22111), .B(n22112), .Z(n22099) );
  AND U23135 ( .A(n22113), .B(n22114), .Z(n22112) );
  XNOR U23136 ( .A(n22111), .B(n11058), .Z(n22114) );
  XNOR U23137 ( .A(n22107), .B(n22109), .Z(n11058) );
  NAND U23138 ( .A(n22115), .B(e_input[207]), .Z(n22109) );
  NAND U23139 ( .A(n12323), .B(e_input[207]), .Z(n22115) );
  XNOR U23140 ( .A(n22105), .B(n22116), .Z(n22107) );
  XOR U23141 ( .A(n22117), .B(n22118), .Z(n22105) );
  AND U23142 ( .A(n22119), .B(n22120), .Z(n22118) );
  XNOR U23143 ( .A(n22121), .B(n22117), .Z(n22120) );
  XOR U23144 ( .A(n22122), .B(e_input[207]), .Z(n22113) );
  IV U23145 ( .A(n22111), .Z(n22122) );
  XOR U23146 ( .A(n22123), .B(n22124), .Z(n22111) );
  AND U23147 ( .A(n22125), .B(n22126), .Z(n22124) );
  XNOR U23148 ( .A(n22123), .B(n11064), .Z(n22126) );
  XNOR U23149 ( .A(n22119), .B(n22121), .Z(n11064) );
  NAND U23150 ( .A(n22127), .B(e_input[206]), .Z(n22121) );
  NAND U23151 ( .A(n12323), .B(e_input[206]), .Z(n22127) );
  XNOR U23152 ( .A(n22117), .B(n22128), .Z(n22119) );
  XOR U23153 ( .A(n22129), .B(n22130), .Z(n22117) );
  AND U23154 ( .A(n22131), .B(n22132), .Z(n22130) );
  XNOR U23155 ( .A(n22133), .B(n22129), .Z(n22132) );
  XOR U23156 ( .A(n22134), .B(e_input[206]), .Z(n22125) );
  IV U23157 ( .A(n22123), .Z(n22134) );
  XOR U23158 ( .A(n22135), .B(n22136), .Z(n22123) );
  AND U23159 ( .A(n22137), .B(n22138), .Z(n22136) );
  XNOR U23160 ( .A(n22135), .B(n11070), .Z(n22138) );
  XNOR U23161 ( .A(n22131), .B(n22133), .Z(n11070) );
  NAND U23162 ( .A(n22139), .B(e_input[205]), .Z(n22133) );
  NAND U23163 ( .A(n12323), .B(e_input[205]), .Z(n22139) );
  XNOR U23164 ( .A(n22129), .B(n22140), .Z(n22131) );
  XOR U23165 ( .A(n22141), .B(n22142), .Z(n22129) );
  AND U23166 ( .A(n22143), .B(n22144), .Z(n22142) );
  XNOR U23167 ( .A(n22145), .B(n22141), .Z(n22144) );
  XOR U23168 ( .A(n22146), .B(e_input[205]), .Z(n22137) );
  IV U23169 ( .A(n22135), .Z(n22146) );
  XOR U23170 ( .A(n22147), .B(n22148), .Z(n22135) );
  AND U23171 ( .A(n22149), .B(n22150), .Z(n22148) );
  XNOR U23172 ( .A(n22147), .B(n11076), .Z(n22150) );
  XNOR U23173 ( .A(n22143), .B(n22145), .Z(n11076) );
  NAND U23174 ( .A(n22151), .B(e_input[204]), .Z(n22145) );
  NAND U23175 ( .A(n12323), .B(e_input[204]), .Z(n22151) );
  XNOR U23176 ( .A(n22141), .B(n22152), .Z(n22143) );
  XOR U23177 ( .A(n22153), .B(n22154), .Z(n22141) );
  AND U23178 ( .A(n22155), .B(n22156), .Z(n22154) );
  XNOR U23179 ( .A(n22157), .B(n22153), .Z(n22156) );
  XOR U23180 ( .A(n22158), .B(e_input[204]), .Z(n22149) );
  IV U23181 ( .A(n22147), .Z(n22158) );
  XOR U23182 ( .A(n22159), .B(n22160), .Z(n22147) );
  AND U23183 ( .A(n22161), .B(n22162), .Z(n22160) );
  XNOR U23184 ( .A(n22159), .B(n11082), .Z(n22162) );
  XNOR U23185 ( .A(n22155), .B(n22157), .Z(n11082) );
  NAND U23186 ( .A(n22163), .B(e_input[203]), .Z(n22157) );
  NAND U23187 ( .A(n12323), .B(e_input[203]), .Z(n22163) );
  XNOR U23188 ( .A(n22153), .B(n22164), .Z(n22155) );
  XOR U23189 ( .A(n22165), .B(n22166), .Z(n22153) );
  AND U23190 ( .A(n22167), .B(n22168), .Z(n22166) );
  XNOR U23191 ( .A(n22169), .B(n22165), .Z(n22168) );
  XOR U23192 ( .A(n22170), .B(e_input[203]), .Z(n22161) );
  IV U23193 ( .A(n22159), .Z(n22170) );
  XOR U23194 ( .A(n22171), .B(n22172), .Z(n22159) );
  AND U23195 ( .A(n22173), .B(n22174), .Z(n22172) );
  XNOR U23196 ( .A(n22171), .B(n11088), .Z(n22174) );
  XNOR U23197 ( .A(n22167), .B(n22169), .Z(n11088) );
  NAND U23198 ( .A(n22175), .B(e_input[202]), .Z(n22169) );
  NAND U23199 ( .A(n12323), .B(e_input[202]), .Z(n22175) );
  XNOR U23200 ( .A(n22165), .B(n22176), .Z(n22167) );
  XOR U23201 ( .A(n22177), .B(n22178), .Z(n22165) );
  AND U23202 ( .A(n22179), .B(n22180), .Z(n22178) );
  XNOR U23203 ( .A(n22181), .B(n22177), .Z(n22180) );
  XOR U23204 ( .A(n22182), .B(e_input[202]), .Z(n22173) );
  IV U23205 ( .A(n22171), .Z(n22182) );
  XOR U23206 ( .A(n22183), .B(n22184), .Z(n22171) );
  AND U23207 ( .A(n22185), .B(n22186), .Z(n22184) );
  XNOR U23208 ( .A(n22183), .B(n11094), .Z(n22186) );
  XNOR U23209 ( .A(n22179), .B(n22181), .Z(n11094) );
  NAND U23210 ( .A(n22187), .B(e_input[201]), .Z(n22181) );
  NAND U23211 ( .A(n12323), .B(e_input[201]), .Z(n22187) );
  XNOR U23212 ( .A(n22177), .B(n22188), .Z(n22179) );
  XOR U23213 ( .A(n22189), .B(n22190), .Z(n22177) );
  AND U23214 ( .A(n22191), .B(n22192), .Z(n22190) );
  XNOR U23215 ( .A(n22193), .B(n22189), .Z(n22192) );
  XOR U23216 ( .A(n22194), .B(e_input[201]), .Z(n22185) );
  IV U23217 ( .A(n22183), .Z(n22194) );
  XOR U23218 ( .A(n22195), .B(n22196), .Z(n22183) );
  AND U23219 ( .A(n22197), .B(n22198), .Z(n22196) );
  XNOR U23220 ( .A(n22195), .B(n11100), .Z(n22198) );
  XNOR U23221 ( .A(n22191), .B(n22193), .Z(n11100) );
  NAND U23222 ( .A(n22199), .B(e_input[200]), .Z(n22193) );
  NAND U23223 ( .A(n12323), .B(e_input[200]), .Z(n22199) );
  XNOR U23224 ( .A(n22189), .B(n22200), .Z(n22191) );
  XOR U23225 ( .A(n22201), .B(n22202), .Z(n22189) );
  AND U23226 ( .A(n22203), .B(n22204), .Z(n22202) );
  XNOR U23227 ( .A(n22205), .B(n22201), .Z(n22204) );
  XOR U23228 ( .A(n22206), .B(e_input[200]), .Z(n22197) );
  IV U23229 ( .A(n22195), .Z(n22206) );
  XOR U23230 ( .A(n22207), .B(n22208), .Z(n22195) );
  AND U23231 ( .A(n22209), .B(n22210), .Z(n22208) );
  XNOR U23232 ( .A(n22207), .B(n11106), .Z(n22210) );
  XNOR U23233 ( .A(n22203), .B(n22205), .Z(n11106) );
  NAND U23234 ( .A(n22211), .B(e_input[199]), .Z(n22205) );
  NAND U23235 ( .A(n12323), .B(e_input[199]), .Z(n22211) );
  XNOR U23236 ( .A(n22201), .B(n22212), .Z(n22203) );
  XOR U23237 ( .A(n22213), .B(n22214), .Z(n22201) );
  AND U23238 ( .A(n22215), .B(n22216), .Z(n22214) );
  XNOR U23239 ( .A(n22217), .B(n22213), .Z(n22216) );
  XOR U23240 ( .A(n22218), .B(e_input[199]), .Z(n22209) );
  IV U23241 ( .A(n22207), .Z(n22218) );
  XOR U23242 ( .A(n22219), .B(n22220), .Z(n22207) );
  AND U23243 ( .A(n22221), .B(n22222), .Z(n22220) );
  XNOR U23244 ( .A(n22219), .B(n11112), .Z(n22222) );
  XNOR U23245 ( .A(n22215), .B(n22217), .Z(n11112) );
  NAND U23246 ( .A(n22223), .B(e_input[198]), .Z(n22217) );
  NAND U23247 ( .A(n12323), .B(e_input[198]), .Z(n22223) );
  XNOR U23248 ( .A(n22213), .B(n22224), .Z(n22215) );
  XOR U23249 ( .A(n22225), .B(n22226), .Z(n22213) );
  AND U23250 ( .A(n22227), .B(n22228), .Z(n22226) );
  XNOR U23251 ( .A(n22229), .B(n22225), .Z(n22228) );
  XOR U23252 ( .A(n22230), .B(e_input[198]), .Z(n22221) );
  IV U23253 ( .A(n22219), .Z(n22230) );
  XOR U23254 ( .A(n22231), .B(n22232), .Z(n22219) );
  AND U23255 ( .A(n22233), .B(n22234), .Z(n22232) );
  XNOR U23256 ( .A(n22231), .B(n11118), .Z(n22234) );
  XNOR U23257 ( .A(n22227), .B(n22229), .Z(n11118) );
  NAND U23258 ( .A(n22235), .B(e_input[197]), .Z(n22229) );
  NAND U23259 ( .A(n12323), .B(e_input[197]), .Z(n22235) );
  XNOR U23260 ( .A(n22225), .B(n22236), .Z(n22227) );
  XOR U23261 ( .A(n22237), .B(n22238), .Z(n22225) );
  AND U23262 ( .A(n22239), .B(n22240), .Z(n22238) );
  XNOR U23263 ( .A(n22241), .B(n22237), .Z(n22240) );
  XOR U23264 ( .A(n22242), .B(e_input[197]), .Z(n22233) );
  IV U23265 ( .A(n22231), .Z(n22242) );
  XOR U23266 ( .A(n22243), .B(n22244), .Z(n22231) );
  AND U23267 ( .A(n22245), .B(n22246), .Z(n22244) );
  XNOR U23268 ( .A(n22243), .B(n11124), .Z(n22246) );
  XNOR U23269 ( .A(n22239), .B(n22241), .Z(n11124) );
  NAND U23270 ( .A(n22247), .B(e_input[196]), .Z(n22241) );
  NAND U23271 ( .A(n12323), .B(e_input[196]), .Z(n22247) );
  XNOR U23272 ( .A(n22237), .B(n22248), .Z(n22239) );
  XOR U23273 ( .A(n22249), .B(n22250), .Z(n22237) );
  AND U23274 ( .A(n22251), .B(n22252), .Z(n22250) );
  XNOR U23275 ( .A(n22253), .B(n22249), .Z(n22252) );
  XOR U23276 ( .A(n22254), .B(e_input[196]), .Z(n22245) );
  IV U23277 ( .A(n22243), .Z(n22254) );
  XOR U23278 ( .A(n22255), .B(n22256), .Z(n22243) );
  AND U23279 ( .A(n22257), .B(n22258), .Z(n22256) );
  XNOR U23280 ( .A(n22255), .B(n11130), .Z(n22258) );
  XNOR U23281 ( .A(n22251), .B(n22253), .Z(n11130) );
  NAND U23282 ( .A(n22259), .B(e_input[195]), .Z(n22253) );
  NAND U23283 ( .A(n12323), .B(e_input[195]), .Z(n22259) );
  XNOR U23284 ( .A(n22249), .B(n22260), .Z(n22251) );
  XOR U23285 ( .A(n22261), .B(n22262), .Z(n22249) );
  AND U23286 ( .A(n22263), .B(n22264), .Z(n22262) );
  XNOR U23287 ( .A(n22265), .B(n22261), .Z(n22264) );
  XOR U23288 ( .A(n22266), .B(e_input[195]), .Z(n22257) );
  IV U23289 ( .A(n22255), .Z(n22266) );
  XOR U23290 ( .A(n22267), .B(n22268), .Z(n22255) );
  AND U23291 ( .A(n22269), .B(n22270), .Z(n22268) );
  XNOR U23292 ( .A(n22267), .B(n11136), .Z(n22270) );
  XNOR U23293 ( .A(n22263), .B(n22265), .Z(n11136) );
  NAND U23294 ( .A(n22271), .B(e_input[194]), .Z(n22265) );
  NAND U23295 ( .A(n12323), .B(e_input[194]), .Z(n22271) );
  XNOR U23296 ( .A(n22261), .B(n22272), .Z(n22263) );
  XOR U23297 ( .A(n22273), .B(n22274), .Z(n22261) );
  AND U23298 ( .A(n22275), .B(n22276), .Z(n22274) );
  XNOR U23299 ( .A(n22277), .B(n22273), .Z(n22276) );
  XOR U23300 ( .A(n22278), .B(e_input[194]), .Z(n22269) );
  IV U23301 ( .A(n22267), .Z(n22278) );
  XOR U23302 ( .A(n22279), .B(n22280), .Z(n22267) );
  AND U23303 ( .A(n22281), .B(n22282), .Z(n22280) );
  XNOR U23304 ( .A(n22279), .B(n11142), .Z(n22282) );
  XNOR U23305 ( .A(n22275), .B(n22277), .Z(n11142) );
  NAND U23306 ( .A(n22283), .B(e_input[193]), .Z(n22277) );
  NAND U23307 ( .A(n12323), .B(e_input[193]), .Z(n22283) );
  XNOR U23308 ( .A(n22273), .B(n22284), .Z(n22275) );
  XOR U23309 ( .A(n22285), .B(n22286), .Z(n22273) );
  AND U23310 ( .A(n22287), .B(n22288), .Z(n22286) );
  XNOR U23311 ( .A(n22289), .B(n22285), .Z(n22288) );
  XOR U23312 ( .A(n22290), .B(e_input[193]), .Z(n22281) );
  IV U23313 ( .A(n22279), .Z(n22290) );
  XOR U23314 ( .A(n22291), .B(n22292), .Z(n22279) );
  AND U23315 ( .A(n22293), .B(n22294), .Z(n22292) );
  XNOR U23316 ( .A(n22291), .B(n11148), .Z(n22294) );
  XNOR U23317 ( .A(n22287), .B(n22289), .Z(n11148) );
  NAND U23318 ( .A(n22295), .B(e_input[192]), .Z(n22289) );
  NAND U23319 ( .A(n12323), .B(e_input[192]), .Z(n22295) );
  XNOR U23320 ( .A(n22285), .B(n22296), .Z(n22287) );
  XOR U23321 ( .A(n22297), .B(n22298), .Z(n22285) );
  AND U23322 ( .A(n22299), .B(n22300), .Z(n22298) );
  XNOR U23323 ( .A(n22301), .B(n22297), .Z(n22300) );
  XOR U23324 ( .A(n22302), .B(e_input[192]), .Z(n22293) );
  IV U23325 ( .A(n22291), .Z(n22302) );
  XOR U23326 ( .A(n22303), .B(n22304), .Z(n22291) );
  AND U23327 ( .A(n22305), .B(n22306), .Z(n22304) );
  XNOR U23328 ( .A(n22303), .B(n11154), .Z(n22306) );
  XNOR U23329 ( .A(n22299), .B(n22301), .Z(n11154) );
  NAND U23330 ( .A(n22307), .B(e_input[191]), .Z(n22301) );
  NAND U23331 ( .A(n12323), .B(e_input[191]), .Z(n22307) );
  XNOR U23332 ( .A(n22297), .B(n22308), .Z(n22299) );
  XOR U23333 ( .A(n22309), .B(n22310), .Z(n22297) );
  AND U23334 ( .A(n22311), .B(n22312), .Z(n22310) );
  XNOR U23335 ( .A(n22313), .B(n22309), .Z(n22312) );
  XOR U23336 ( .A(n22314), .B(e_input[191]), .Z(n22305) );
  IV U23337 ( .A(n22303), .Z(n22314) );
  XOR U23338 ( .A(n22315), .B(n22316), .Z(n22303) );
  AND U23339 ( .A(n22317), .B(n22318), .Z(n22316) );
  XNOR U23340 ( .A(n22315), .B(n11160), .Z(n22318) );
  XNOR U23341 ( .A(n22311), .B(n22313), .Z(n11160) );
  NAND U23342 ( .A(n22319), .B(e_input[190]), .Z(n22313) );
  NAND U23343 ( .A(n12323), .B(e_input[190]), .Z(n22319) );
  XNOR U23344 ( .A(n22309), .B(n22320), .Z(n22311) );
  XOR U23345 ( .A(n22321), .B(n22322), .Z(n22309) );
  AND U23346 ( .A(n22323), .B(n22324), .Z(n22322) );
  XNOR U23347 ( .A(n22325), .B(n22321), .Z(n22324) );
  XOR U23348 ( .A(n22326), .B(e_input[190]), .Z(n22317) );
  IV U23349 ( .A(n22315), .Z(n22326) );
  XOR U23350 ( .A(n22327), .B(n22328), .Z(n22315) );
  AND U23351 ( .A(n22329), .B(n22330), .Z(n22328) );
  XNOR U23352 ( .A(n22327), .B(n11166), .Z(n22330) );
  XNOR U23353 ( .A(n22323), .B(n22325), .Z(n11166) );
  NAND U23354 ( .A(n22331), .B(e_input[189]), .Z(n22325) );
  NAND U23355 ( .A(n12323), .B(e_input[189]), .Z(n22331) );
  XNOR U23356 ( .A(n22321), .B(n22332), .Z(n22323) );
  XOR U23357 ( .A(n22333), .B(n22334), .Z(n22321) );
  AND U23358 ( .A(n22335), .B(n22336), .Z(n22334) );
  XNOR U23359 ( .A(n22337), .B(n22333), .Z(n22336) );
  XOR U23360 ( .A(n22338), .B(e_input[189]), .Z(n22329) );
  IV U23361 ( .A(n22327), .Z(n22338) );
  XOR U23362 ( .A(n22339), .B(n22340), .Z(n22327) );
  AND U23363 ( .A(n22341), .B(n22342), .Z(n22340) );
  XNOR U23364 ( .A(n22339), .B(n11172), .Z(n22342) );
  XNOR U23365 ( .A(n22335), .B(n22337), .Z(n11172) );
  NAND U23366 ( .A(n22343), .B(e_input[188]), .Z(n22337) );
  NAND U23367 ( .A(n12323), .B(e_input[188]), .Z(n22343) );
  XNOR U23368 ( .A(n22333), .B(n22344), .Z(n22335) );
  XOR U23369 ( .A(n22345), .B(n22346), .Z(n22333) );
  AND U23370 ( .A(n22347), .B(n22348), .Z(n22346) );
  XNOR U23371 ( .A(n22349), .B(n22345), .Z(n22348) );
  XOR U23372 ( .A(n22350), .B(e_input[188]), .Z(n22341) );
  IV U23373 ( .A(n22339), .Z(n22350) );
  XOR U23374 ( .A(n22351), .B(n22352), .Z(n22339) );
  AND U23375 ( .A(n22353), .B(n22354), .Z(n22352) );
  XNOR U23376 ( .A(n22351), .B(n11178), .Z(n22354) );
  XNOR U23377 ( .A(n22347), .B(n22349), .Z(n11178) );
  NAND U23378 ( .A(n22355), .B(e_input[187]), .Z(n22349) );
  NAND U23379 ( .A(n12323), .B(e_input[187]), .Z(n22355) );
  XNOR U23380 ( .A(n22345), .B(n22356), .Z(n22347) );
  XOR U23381 ( .A(n22357), .B(n22358), .Z(n22345) );
  AND U23382 ( .A(n22359), .B(n22360), .Z(n22358) );
  XNOR U23383 ( .A(n22361), .B(n22357), .Z(n22360) );
  XOR U23384 ( .A(n22362), .B(e_input[187]), .Z(n22353) );
  IV U23385 ( .A(n22351), .Z(n22362) );
  XOR U23386 ( .A(n22363), .B(n22364), .Z(n22351) );
  AND U23387 ( .A(n22365), .B(n22366), .Z(n22364) );
  XNOR U23388 ( .A(n22363), .B(n11184), .Z(n22366) );
  XNOR U23389 ( .A(n22359), .B(n22361), .Z(n11184) );
  NAND U23390 ( .A(n22367), .B(e_input[186]), .Z(n22361) );
  NAND U23391 ( .A(n12323), .B(e_input[186]), .Z(n22367) );
  XNOR U23392 ( .A(n22357), .B(n22368), .Z(n22359) );
  XOR U23393 ( .A(n22369), .B(n22370), .Z(n22357) );
  AND U23394 ( .A(n22371), .B(n22372), .Z(n22370) );
  XNOR U23395 ( .A(n22373), .B(n22369), .Z(n22372) );
  XOR U23396 ( .A(n22374), .B(e_input[186]), .Z(n22365) );
  IV U23397 ( .A(n22363), .Z(n22374) );
  XOR U23398 ( .A(n22375), .B(n22376), .Z(n22363) );
  AND U23399 ( .A(n22377), .B(n22378), .Z(n22376) );
  XNOR U23400 ( .A(n22375), .B(n11190), .Z(n22378) );
  XNOR U23401 ( .A(n22371), .B(n22373), .Z(n11190) );
  NAND U23402 ( .A(n22379), .B(e_input[185]), .Z(n22373) );
  NAND U23403 ( .A(n12323), .B(e_input[185]), .Z(n22379) );
  XNOR U23404 ( .A(n22369), .B(n22380), .Z(n22371) );
  XOR U23405 ( .A(n22381), .B(n22382), .Z(n22369) );
  AND U23406 ( .A(n22383), .B(n22384), .Z(n22382) );
  XNOR U23407 ( .A(n22385), .B(n22381), .Z(n22384) );
  XOR U23408 ( .A(n22386), .B(e_input[185]), .Z(n22377) );
  IV U23409 ( .A(n22375), .Z(n22386) );
  XOR U23410 ( .A(n22387), .B(n22388), .Z(n22375) );
  AND U23411 ( .A(n22389), .B(n22390), .Z(n22388) );
  XNOR U23412 ( .A(n22387), .B(n11196), .Z(n22390) );
  XNOR U23413 ( .A(n22383), .B(n22385), .Z(n11196) );
  NAND U23414 ( .A(n22391), .B(e_input[184]), .Z(n22385) );
  NAND U23415 ( .A(n12323), .B(e_input[184]), .Z(n22391) );
  XNOR U23416 ( .A(n22381), .B(n22392), .Z(n22383) );
  XOR U23417 ( .A(n22393), .B(n22394), .Z(n22381) );
  AND U23418 ( .A(n22395), .B(n22396), .Z(n22394) );
  XNOR U23419 ( .A(n22397), .B(n22393), .Z(n22396) );
  XOR U23420 ( .A(n22398), .B(e_input[184]), .Z(n22389) );
  IV U23421 ( .A(n22387), .Z(n22398) );
  XOR U23422 ( .A(n22399), .B(n22400), .Z(n22387) );
  AND U23423 ( .A(n22401), .B(n22402), .Z(n22400) );
  XNOR U23424 ( .A(n22399), .B(n11202), .Z(n22402) );
  XNOR U23425 ( .A(n22395), .B(n22397), .Z(n11202) );
  NAND U23426 ( .A(n22403), .B(e_input[183]), .Z(n22397) );
  NAND U23427 ( .A(n12323), .B(e_input[183]), .Z(n22403) );
  XNOR U23428 ( .A(n22393), .B(n22404), .Z(n22395) );
  XOR U23429 ( .A(n22405), .B(n22406), .Z(n22393) );
  AND U23430 ( .A(n22407), .B(n22408), .Z(n22406) );
  XNOR U23431 ( .A(n22409), .B(n22405), .Z(n22408) );
  XOR U23432 ( .A(n22410), .B(e_input[183]), .Z(n22401) );
  IV U23433 ( .A(n22399), .Z(n22410) );
  XOR U23434 ( .A(n22411), .B(n22412), .Z(n22399) );
  AND U23435 ( .A(n22413), .B(n22414), .Z(n22412) );
  XNOR U23436 ( .A(n22411), .B(n11208), .Z(n22414) );
  XNOR U23437 ( .A(n22407), .B(n22409), .Z(n11208) );
  NAND U23438 ( .A(n22415), .B(e_input[182]), .Z(n22409) );
  NAND U23439 ( .A(n12323), .B(e_input[182]), .Z(n22415) );
  XNOR U23440 ( .A(n22405), .B(n22416), .Z(n22407) );
  XOR U23441 ( .A(n22417), .B(n22418), .Z(n22405) );
  AND U23442 ( .A(n22419), .B(n22420), .Z(n22418) );
  XNOR U23443 ( .A(n22421), .B(n22417), .Z(n22420) );
  XOR U23444 ( .A(n22422), .B(e_input[182]), .Z(n22413) );
  IV U23445 ( .A(n22411), .Z(n22422) );
  XOR U23446 ( .A(n22423), .B(n22424), .Z(n22411) );
  AND U23447 ( .A(n22425), .B(n22426), .Z(n22424) );
  XNOR U23448 ( .A(n22423), .B(n11214), .Z(n22426) );
  XNOR U23449 ( .A(n22419), .B(n22421), .Z(n11214) );
  NAND U23450 ( .A(n22427), .B(e_input[181]), .Z(n22421) );
  NAND U23451 ( .A(n12323), .B(e_input[181]), .Z(n22427) );
  XNOR U23452 ( .A(n22417), .B(n22428), .Z(n22419) );
  XOR U23453 ( .A(n22429), .B(n22430), .Z(n22417) );
  AND U23454 ( .A(n22431), .B(n22432), .Z(n22430) );
  XNOR U23455 ( .A(n22433), .B(n22429), .Z(n22432) );
  XOR U23456 ( .A(n22434), .B(e_input[181]), .Z(n22425) );
  IV U23457 ( .A(n22423), .Z(n22434) );
  XOR U23458 ( .A(n22435), .B(n22436), .Z(n22423) );
  AND U23459 ( .A(n22437), .B(n22438), .Z(n22436) );
  XNOR U23460 ( .A(n22435), .B(n11220), .Z(n22438) );
  XNOR U23461 ( .A(n22431), .B(n22433), .Z(n11220) );
  NAND U23462 ( .A(n22439), .B(e_input[180]), .Z(n22433) );
  NAND U23463 ( .A(n12323), .B(e_input[180]), .Z(n22439) );
  XNOR U23464 ( .A(n22429), .B(n22440), .Z(n22431) );
  XOR U23465 ( .A(n22441), .B(n22442), .Z(n22429) );
  AND U23466 ( .A(n22443), .B(n22444), .Z(n22442) );
  XNOR U23467 ( .A(n22445), .B(n22441), .Z(n22444) );
  XOR U23468 ( .A(n22446), .B(e_input[180]), .Z(n22437) );
  IV U23469 ( .A(n22435), .Z(n22446) );
  XOR U23470 ( .A(n22447), .B(n22448), .Z(n22435) );
  AND U23471 ( .A(n22449), .B(n22450), .Z(n22448) );
  XNOR U23472 ( .A(n22447), .B(n11226), .Z(n22450) );
  XNOR U23473 ( .A(n22443), .B(n22445), .Z(n11226) );
  NAND U23474 ( .A(n22451), .B(e_input[179]), .Z(n22445) );
  NAND U23475 ( .A(n12323), .B(e_input[179]), .Z(n22451) );
  XNOR U23476 ( .A(n22441), .B(n22452), .Z(n22443) );
  XOR U23477 ( .A(n22453), .B(n22454), .Z(n22441) );
  AND U23478 ( .A(n22455), .B(n22456), .Z(n22454) );
  XNOR U23479 ( .A(n22457), .B(n22453), .Z(n22456) );
  XOR U23480 ( .A(n22458), .B(e_input[179]), .Z(n22449) );
  IV U23481 ( .A(n22447), .Z(n22458) );
  XOR U23482 ( .A(n22459), .B(n22460), .Z(n22447) );
  AND U23483 ( .A(n22461), .B(n22462), .Z(n22460) );
  XNOR U23484 ( .A(n22459), .B(n11232), .Z(n22462) );
  XNOR U23485 ( .A(n22455), .B(n22457), .Z(n11232) );
  NAND U23486 ( .A(n22463), .B(e_input[178]), .Z(n22457) );
  NAND U23487 ( .A(n12323), .B(e_input[178]), .Z(n22463) );
  XNOR U23488 ( .A(n22453), .B(n22464), .Z(n22455) );
  XOR U23489 ( .A(n22465), .B(n22466), .Z(n22453) );
  AND U23490 ( .A(n22467), .B(n22468), .Z(n22466) );
  XNOR U23491 ( .A(n22469), .B(n22465), .Z(n22468) );
  XOR U23492 ( .A(n22470), .B(e_input[178]), .Z(n22461) );
  IV U23493 ( .A(n22459), .Z(n22470) );
  XOR U23494 ( .A(n22471), .B(n22472), .Z(n22459) );
  AND U23495 ( .A(n22473), .B(n22474), .Z(n22472) );
  XNOR U23496 ( .A(n22471), .B(n11238), .Z(n22474) );
  XNOR U23497 ( .A(n22467), .B(n22469), .Z(n11238) );
  NAND U23498 ( .A(n22475), .B(e_input[177]), .Z(n22469) );
  NAND U23499 ( .A(n12323), .B(e_input[177]), .Z(n22475) );
  XNOR U23500 ( .A(n22465), .B(n22476), .Z(n22467) );
  XOR U23501 ( .A(n22477), .B(n22478), .Z(n22465) );
  AND U23502 ( .A(n22479), .B(n22480), .Z(n22478) );
  XNOR U23503 ( .A(n22481), .B(n22477), .Z(n22480) );
  XOR U23504 ( .A(n22482), .B(e_input[177]), .Z(n22473) );
  IV U23505 ( .A(n22471), .Z(n22482) );
  XOR U23506 ( .A(n22483), .B(n22484), .Z(n22471) );
  AND U23507 ( .A(n22485), .B(n22486), .Z(n22484) );
  XNOR U23508 ( .A(n22483), .B(n11244), .Z(n22486) );
  XNOR U23509 ( .A(n22479), .B(n22481), .Z(n11244) );
  NAND U23510 ( .A(n22487), .B(e_input[176]), .Z(n22481) );
  NAND U23511 ( .A(n12323), .B(e_input[176]), .Z(n22487) );
  XNOR U23512 ( .A(n22477), .B(n22488), .Z(n22479) );
  XOR U23513 ( .A(n22489), .B(n22490), .Z(n22477) );
  AND U23514 ( .A(n22491), .B(n22492), .Z(n22490) );
  XNOR U23515 ( .A(n22493), .B(n22489), .Z(n22492) );
  XOR U23516 ( .A(n22494), .B(e_input[176]), .Z(n22485) );
  IV U23517 ( .A(n22483), .Z(n22494) );
  XOR U23518 ( .A(n22495), .B(n22496), .Z(n22483) );
  AND U23519 ( .A(n22497), .B(n22498), .Z(n22496) );
  XNOR U23520 ( .A(n22495), .B(n11250), .Z(n22498) );
  XNOR U23521 ( .A(n22491), .B(n22493), .Z(n11250) );
  NAND U23522 ( .A(n22499), .B(e_input[175]), .Z(n22493) );
  NAND U23523 ( .A(n12323), .B(e_input[175]), .Z(n22499) );
  XNOR U23524 ( .A(n22489), .B(n22500), .Z(n22491) );
  XOR U23525 ( .A(n22501), .B(n22502), .Z(n22489) );
  AND U23526 ( .A(n22503), .B(n22504), .Z(n22502) );
  XNOR U23527 ( .A(n22505), .B(n22501), .Z(n22504) );
  XOR U23528 ( .A(n22506), .B(e_input[175]), .Z(n22497) );
  IV U23529 ( .A(n22495), .Z(n22506) );
  XOR U23530 ( .A(n22507), .B(n22508), .Z(n22495) );
  AND U23531 ( .A(n22509), .B(n22510), .Z(n22508) );
  XNOR U23532 ( .A(n22507), .B(n11256), .Z(n22510) );
  XNOR U23533 ( .A(n22503), .B(n22505), .Z(n11256) );
  NAND U23534 ( .A(n22511), .B(e_input[174]), .Z(n22505) );
  NAND U23535 ( .A(n12323), .B(e_input[174]), .Z(n22511) );
  XNOR U23536 ( .A(n22501), .B(n22512), .Z(n22503) );
  XOR U23537 ( .A(n22513), .B(n22514), .Z(n22501) );
  AND U23538 ( .A(n22515), .B(n22516), .Z(n22514) );
  XNOR U23539 ( .A(n22517), .B(n22513), .Z(n22516) );
  XOR U23540 ( .A(n22518), .B(e_input[174]), .Z(n22509) );
  IV U23541 ( .A(n22507), .Z(n22518) );
  XOR U23542 ( .A(n22519), .B(n22520), .Z(n22507) );
  AND U23543 ( .A(n22521), .B(n22522), .Z(n22520) );
  XNOR U23544 ( .A(n22519), .B(n11262), .Z(n22522) );
  XNOR U23545 ( .A(n22515), .B(n22517), .Z(n11262) );
  NAND U23546 ( .A(n22523), .B(e_input[173]), .Z(n22517) );
  NAND U23547 ( .A(n12323), .B(e_input[173]), .Z(n22523) );
  XNOR U23548 ( .A(n22513), .B(n22524), .Z(n22515) );
  XOR U23549 ( .A(n22525), .B(n22526), .Z(n22513) );
  AND U23550 ( .A(n22527), .B(n22528), .Z(n22526) );
  XNOR U23551 ( .A(n22529), .B(n22525), .Z(n22528) );
  XOR U23552 ( .A(n22530), .B(e_input[173]), .Z(n22521) );
  IV U23553 ( .A(n22519), .Z(n22530) );
  XOR U23554 ( .A(n22531), .B(n22532), .Z(n22519) );
  AND U23555 ( .A(n22533), .B(n22534), .Z(n22532) );
  XNOR U23556 ( .A(n22531), .B(n11268), .Z(n22534) );
  XNOR U23557 ( .A(n22527), .B(n22529), .Z(n11268) );
  NAND U23558 ( .A(n22535), .B(e_input[172]), .Z(n22529) );
  NAND U23559 ( .A(n12323), .B(e_input[172]), .Z(n22535) );
  XNOR U23560 ( .A(n22525), .B(n22536), .Z(n22527) );
  XOR U23561 ( .A(n22537), .B(n22538), .Z(n22525) );
  AND U23562 ( .A(n22539), .B(n22540), .Z(n22538) );
  XNOR U23563 ( .A(n22541), .B(n22537), .Z(n22540) );
  XOR U23564 ( .A(n22542), .B(e_input[172]), .Z(n22533) );
  IV U23565 ( .A(n22531), .Z(n22542) );
  XOR U23566 ( .A(n22543), .B(n22544), .Z(n22531) );
  AND U23567 ( .A(n22545), .B(n22546), .Z(n22544) );
  XNOR U23568 ( .A(n22543), .B(n11274), .Z(n22546) );
  XNOR U23569 ( .A(n22539), .B(n22541), .Z(n11274) );
  NAND U23570 ( .A(n22547), .B(e_input[171]), .Z(n22541) );
  NAND U23571 ( .A(n12323), .B(e_input[171]), .Z(n22547) );
  XNOR U23572 ( .A(n22537), .B(n22548), .Z(n22539) );
  XOR U23573 ( .A(n22549), .B(n22550), .Z(n22537) );
  AND U23574 ( .A(n22551), .B(n22552), .Z(n22550) );
  XNOR U23575 ( .A(n22553), .B(n22549), .Z(n22552) );
  XOR U23576 ( .A(n22554), .B(e_input[171]), .Z(n22545) );
  IV U23577 ( .A(n22543), .Z(n22554) );
  XOR U23578 ( .A(n22555), .B(n22556), .Z(n22543) );
  AND U23579 ( .A(n22557), .B(n22558), .Z(n22556) );
  XNOR U23580 ( .A(n22555), .B(n11280), .Z(n22558) );
  XNOR U23581 ( .A(n22551), .B(n22553), .Z(n11280) );
  NAND U23582 ( .A(n22559), .B(e_input[170]), .Z(n22553) );
  NAND U23583 ( .A(n12323), .B(e_input[170]), .Z(n22559) );
  XNOR U23584 ( .A(n22549), .B(n22560), .Z(n22551) );
  XOR U23585 ( .A(n22561), .B(n22562), .Z(n22549) );
  AND U23586 ( .A(n22563), .B(n22564), .Z(n22562) );
  XNOR U23587 ( .A(n22565), .B(n22561), .Z(n22564) );
  XOR U23588 ( .A(n22566), .B(e_input[170]), .Z(n22557) );
  IV U23589 ( .A(n22555), .Z(n22566) );
  XOR U23590 ( .A(n22567), .B(n22568), .Z(n22555) );
  AND U23591 ( .A(n22569), .B(n22570), .Z(n22568) );
  XNOR U23592 ( .A(n22567), .B(n11286), .Z(n22570) );
  XNOR U23593 ( .A(n22563), .B(n22565), .Z(n11286) );
  NAND U23594 ( .A(n22571), .B(e_input[169]), .Z(n22565) );
  NAND U23595 ( .A(n12323), .B(e_input[169]), .Z(n22571) );
  XNOR U23596 ( .A(n22561), .B(n22572), .Z(n22563) );
  XOR U23597 ( .A(n22573), .B(n22574), .Z(n22561) );
  AND U23598 ( .A(n22575), .B(n22576), .Z(n22574) );
  XNOR U23599 ( .A(n22577), .B(n22573), .Z(n22576) );
  XOR U23600 ( .A(n22578), .B(e_input[169]), .Z(n22569) );
  IV U23601 ( .A(n22567), .Z(n22578) );
  XOR U23602 ( .A(n22579), .B(n22580), .Z(n22567) );
  AND U23603 ( .A(n22581), .B(n22582), .Z(n22580) );
  XNOR U23604 ( .A(n22579), .B(n11292), .Z(n22582) );
  XNOR U23605 ( .A(n22575), .B(n22577), .Z(n11292) );
  NAND U23606 ( .A(n22583), .B(e_input[168]), .Z(n22577) );
  NAND U23607 ( .A(n12323), .B(e_input[168]), .Z(n22583) );
  XNOR U23608 ( .A(n22573), .B(n22584), .Z(n22575) );
  XOR U23609 ( .A(n22585), .B(n22586), .Z(n22573) );
  AND U23610 ( .A(n22587), .B(n22588), .Z(n22586) );
  XNOR U23611 ( .A(n22589), .B(n22585), .Z(n22588) );
  XOR U23612 ( .A(n22590), .B(e_input[168]), .Z(n22581) );
  IV U23613 ( .A(n22579), .Z(n22590) );
  XOR U23614 ( .A(n22591), .B(n22592), .Z(n22579) );
  AND U23615 ( .A(n22593), .B(n22594), .Z(n22592) );
  XNOR U23616 ( .A(n22591), .B(n11298), .Z(n22594) );
  XNOR U23617 ( .A(n22587), .B(n22589), .Z(n11298) );
  NAND U23618 ( .A(n22595), .B(e_input[167]), .Z(n22589) );
  NAND U23619 ( .A(n12323), .B(e_input[167]), .Z(n22595) );
  XNOR U23620 ( .A(n22585), .B(n22596), .Z(n22587) );
  XOR U23621 ( .A(n22597), .B(n22598), .Z(n22585) );
  AND U23622 ( .A(n22599), .B(n22600), .Z(n22598) );
  XNOR U23623 ( .A(n22601), .B(n22597), .Z(n22600) );
  XOR U23624 ( .A(n22602), .B(e_input[167]), .Z(n22593) );
  IV U23625 ( .A(n22591), .Z(n22602) );
  XOR U23626 ( .A(n22603), .B(n22604), .Z(n22591) );
  AND U23627 ( .A(n22605), .B(n22606), .Z(n22604) );
  XNOR U23628 ( .A(n22603), .B(n11304), .Z(n22606) );
  XNOR U23629 ( .A(n22599), .B(n22601), .Z(n11304) );
  NAND U23630 ( .A(n22607), .B(e_input[166]), .Z(n22601) );
  NAND U23631 ( .A(n12323), .B(e_input[166]), .Z(n22607) );
  XNOR U23632 ( .A(n22597), .B(n22608), .Z(n22599) );
  XOR U23633 ( .A(n22609), .B(n22610), .Z(n22597) );
  AND U23634 ( .A(n22611), .B(n22612), .Z(n22610) );
  XNOR U23635 ( .A(n22613), .B(n22609), .Z(n22612) );
  XOR U23636 ( .A(n22614), .B(e_input[166]), .Z(n22605) );
  IV U23637 ( .A(n22603), .Z(n22614) );
  XOR U23638 ( .A(n22615), .B(n22616), .Z(n22603) );
  AND U23639 ( .A(n22617), .B(n22618), .Z(n22616) );
  XNOR U23640 ( .A(n22615), .B(n11310), .Z(n22618) );
  XNOR U23641 ( .A(n22611), .B(n22613), .Z(n11310) );
  NAND U23642 ( .A(n22619), .B(e_input[165]), .Z(n22613) );
  NAND U23643 ( .A(n12323), .B(e_input[165]), .Z(n22619) );
  XNOR U23644 ( .A(n22609), .B(n22620), .Z(n22611) );
  XOR U23645 ( .A(n22621), .B(n22622), .Z(n22609) );
  AND U23646 ( .A(n22623), .B(n22624), .Z(n22622) );
  XNOR U23647 ( .A(n22625), .B(n22621), .Z(n22624) );
  XOR U23648 ( .A(n22626), .B(e_input[165]), .Z(n22617) );
  IV U23649 ( .A(n22615), .Z(n22626) );
  XOR U23650 ( .A(n22627), .B(n22628), .Z(n22615) );
  AND U23651 ( .A(n22629), .B(n22630), .Z(n22628) );
  XNOR U23652 ( .A(n22627), .B(n11316), .Z(n22630) );
  XNOR U23653 ( .A(n22623), .B(n22625), .Z(n11316) );
  NAND U23654 ( .A(n22631), .B(e_input[164]), .Z(n22625) );
  NAND U23655 ( .A(n12323), .B(e_input[164]), .Z(n22631) );
  XNOR U23656 ( .A(n22621), .B(n22632), .Z(n22623) );
  XOR U23657 ( .A(n22633), .B(n22634), .Z(n22621) );
  AND U23658 ( .A(n22635), .B(n22636), .Z(n22634) );
  XNOR U23659 ( .A(n22637), .B(n22633), .Z(n22636) );
  XOR U23660 ( .A(n22638), .B(e_input[164]), .Z(n22629) );
  IV U23661 ( .A(n22627), .Z(n22638) );
  XOR U23662 ( .A(n22639), .B(n22640), .Z(n22627) );
  AND U23663 ( .A(n22641), .B(n22642), .Z(n22640) );
  XNOR U23664 ( .A(n22639), .B(n11322), .Z(n22642) );
  XNOR U23665 ( .A(n22635), .B(n22637), .Z(n11322) );
  NAND U23666 ( .A(n22643), .B(e_input[163]), .Z(n22637) );
  NAND U23667 ( .A(n12323), .B(e_input[163]), .Z(n22643) );
  XNOR U23668 ( .A(n22633), .B(n22644), .Z(n22635) );
  XOR U23669 ( .A(n22645), .B(n22646), .Z(n22633) );
  AND U23670 ( .A(n22647), .B(n22648), .Z(n22646) );
  XNOR U23671 ( .A(n22649), .B(n22645), .Z(n22648) );
  XOR U23672 ( .A(n22650), .B(e_input[163]), .Z(n22641) );
  IV U23673 ( .A(n22639), .Z(n22650) );
  XOR U23674 ( .A(n22651), .B(n22652), .Z(n22639) );
  AND U23675 ( .A(n22653), .B(n22654), .Z(n22652) );
  XNOR U23676 ( .A(n22651), .B(n11328), .Z(n22654) );
  XNOR U23677 ( .A(n22647), .B(n22649), .Z(n11328) );
  NAND U23678 ( .A(n22655), .B(e_input[162]), .Z(n22649) );
  NAND U23679 ( .A(n12323), .B(e_input[162]), .Z(n22655) );
  XNOR U23680 ( .A(n22645), .B(n22656), .Z(n22647) );
  XOR U23681 ( .A(n22657), .B(n22658), .Z(n22645) );
  AND U23682 ( .A(n22659), .B(n22660), .Z(n22658) );
  XNOR U23683 ( .A(n22661), .B(n22657), .Z(n22660) );
  XOR U23684 ( .A(n22662), .B(e_input[162]), .Z(n22653) );
  IV U23685 ( .A(n22651), .Z(n22662) );
  XOR U23686 ( .A(n22663), .B(n22664), .Z(n22651) );
  AND U23687 ( .A(n22665), .B(n22666), .Z(n22664) );
  XNOR U23688 ( .A(n22663), .B(n11334), .Z(n22666) );
  XNOR U23689 ( .A(n22659), .B(n22661), .Z(n11334) );
  NAND U23690 ( .A(n22667), .B(e_input[161]), .Z(n22661) );
  NAND U23691 ( .A(n12323), .B(e_input[161]), .Z(n22667) );
  XNOR U23692 ( .A(n22657), .B(n22668), .Z(n22659) );
  XOR U23693 ( .A(n22669), .B(n22670), .Z(n22657) );
  AND U23694 ( .A(n22671), .B(n22672), .Z(n22670) );
  XNOR U23695 ( .A(n22673), .B(n22669), .Z(n22672) );
  XOR U23696 ( .A(n22674), .B(e_input[161]), .Z(n22665) );
  IV U23697 ( .A(n22663), .Z(n22674) );
  XOR U23698 ( .A(n22675), .B(n22676), .Z(n22663) );
  AND U23699 ( .A(n22677), .B(n22678), .Z(n22676) );
  XNOR U23700 ( .A(n22675), .B(n11340), .Z(n22678) );
  XNOR U23701 ( .A(n22671), .B(n22673), .Z(n11340) );
  NAND U23702 ( .A(n22679), .B(e_input[160]), .Z(n22673) );
  NAND U23703 ( .A(n12323), .B(e_input[160]), .Z(n22679) );
  XNOR U23704 ( .A(n22669), .B(n22680), .Z(n22671) );
  XOR U23705 ( .A(n22681), .B(n22682), .Z(n22669) );
  AND U23706 ( .A(n22683), .B(n22684), .Z(n22682) );
  XNOR U23707 ( .A(n22685), .B(n22681), .Z(n22684) );
  XOR U23708 ( .A(n22686), .B(e_input[160]), .Z(n22677) );
  IV U23709 ( .A(n22675), .Z(n22686) );
  XOR U23710 ( .A(n22687), .B(n22688), .Z(n22675) );
  AND U23711 ( .A(n22689), .B(n22690), .Z(n22688) );
  XNOR U23712 ( .A(n22687), .B(n11346), .Z(n22690) );
  XNOR U23713 ( .A(n22683), .B(n22685), .Z(n11346) );
  NAND U23714 ( .A(n22691), .B(e_input[159]), .Z(n22685) );
  NAND U23715 ( .A(n12323), .B(e_input[159]), .Z(n22691) );
  XNOR U23716 ( .A(n22681), .B(n22692), .Z(n22683) );
  XOR U23717 ( .A(n22693), .B(n22694), .Z(n22681) );
  AND U23718 ( .A(n22695), .B(n22696), .Z(n22694) );
  XNOR U23719 ( .A(n22697), .B(n22693), .Z(n22696) );
  XOR U23720 ( .A(n22698), .B(e_input[159]), .Z(n22689) );
  IV U23721 ( .A(n22687), .Z(n22698) );
  XOR U23722 ( .A(n22699), .B(n22700), .Z(n22687) );
  AND U23723 ( .A(n22701), .B(n22702), .Z(n22700) );
  XNOR U23724 ( .A(n22699), .B(n11352), .Z(n22702) );
  XNOR U23725 ( .A(n22695), .B(n22697), .Z(n11352) );
  NAND U23726 ( .A(n22703), .B(e_input[158]), .Z(n22697) );
  NAND U23727 ( .A(n12323), .B(e_input[158]), .Z(n22703) );
  XNOR U23728 ( .A(n22693), .B(n22704), .Z(n22695) );
  XOR U23729 ( .A(n22705), .B(n22706), .Z(n22693) );
  AND U23730 ( .A(n22707), .B(n22708), .Z(n22706) );
  XNOR U23731 ( .A(n22709), .B(n22705), .Z(n22708) );
  XOR U23732 ( .A(n22710), .B(e_input[158]), .Z(n22701) );
  IV U23733 ( .A(n22699), .Z(n22710) );
  XOR U23734 ( .A(n22711), .B(n22712), .Z(n22699) );
  AND U23735 ( .A(n22713), .B(n22714), .Z(n22712) );
  XNOR U23736 ( .A(n22711), .B(n11358), .Z(n22714) );
  XNOR U23737 ( .A(n22707), .B(n22709), .Z(n11358) );
  NAND U23738 ( .A(n22715), .B(e_input[157]), .Z(n22709) );
  NAND U23739 ( .A(n12323), .B(e_input[157]), .Z(n22715) );
  XNOR U23740 ( .A(n22705), .B(n22716), .Z(n22707) );
  XOR U23741 ( .A(n22717), .B(n22718), .Z(n22705) );
  AND U23742 ( .A(n22719), .B(n22720), .Z(n22718) );
  XNOR U23743 ( .A(n22721), .B(n22717), .Z(n22720) );
  XOR U23744 ( .A(n22722), .B(e_input[157]), .Z(n22713) );
  IV U23745 ( .A(n22711), .Z(n22722) );
  XOR U23746 ( .A(n22723), .B(n22724), .Z(n22711) );
  AND U23747 ( .A(n22725), .B(n22726), .Z(n22724) );
  XNOR U23748 ( .A(n22723), .B(n11364), .Z(n22726) );
  XNOR U23749 ( .A(n22719), .B(n22721), .Z(n11364) );
  NAND U23750 ( .A(n22727), .B(e_input[156]), .Z(n22721) );
  NAND U23751 ( .A(n12323), .B(e_input[156]), .Z(n22727) );
  XNOR U23752 ( .A(n22717), .B(n22728), .Z(n22719) );
  XOR U23753 ( .A(n22729), .B(n22730), .Z(n22717) );
  AND U23754 ( .A(n22731), .B(n22732), .Z(n22730) );
  XNOR U23755 ( .A(n22733), .B(n22729), .Z(n22732) );
  XOR U23756 ( .A(n22734), .B(e_input[156]), .Z(n22725) );
  IV U23757 ( .A(n22723), .Z(n22734) );
  XOR U23758 ( .A(n22735), .B(n22736), .Z(n22723) );
  AND U23759 ( .A(n22737), .B(n22738), .Z(n22736) );
  XNOR U23760 ( .A(n22735), .B(n11370), .Z(n22738) );
  XNOR U23761 ( .A(n22731), .B(n22733), .Z(n11370) );
  NAND U23762 ( .A(n22739), .B(e_input[155]), .Z(n22733) );
  NAND U23763 ( .A(n12323), .B(e_input[155]), .Z(n22739) );
  XNOR U23764 ( .A(n22729), .B(n22740), .Z(n22731) );
  XOR U23765 ( .A(n22741), .B(n22742), .Z(n22729) );
  AND U23766 ( .A(n22743), .B(n22744), .Z(n22742) );
  XNOR U23767 ( .A(n22745), .B(n22741), .Z(n22744) );
  XOR U23768 ( .A(n22746), .B(e_input[155]), .Z(n22737) );
  IV U23769 ( .A(n22735), .Z(n22746) );
  XOR U23770 ( .A(n22747), .B(n22748), .Z(n22735) );
  AND U23771 ( .A(n22749), .B(n22750), .Z(n22748) );
  XNOR U23772 ( .A(n22747), .B(n11376), .Z(n22750) );
  XNOR U23773 ( .A(n22743), .B(n22745), .Z(n11376) );
  NAND U23774 ( .A(n22751), .B(e_input[154]), .Z(n22745) );
  NAND U23775 ( .A(n12323), .B(e_input[154]), .Z(n22751) );
  XNOR U23776 ( .A(n22741), .B(n22752), .Z(n22743) );
  XOR U23777 ( .A(n22753), .B(n22754), .Z(n22741) );
  AND U23778 ( .A(n22755), .B(n22756), .Z(n22754) );
  XNOR U23779 ( .A(n22757), .B(n22753), .Z(n22756) );
  XOR U23780 ( .A(n22758), .B(e_input[154]), .Z(n22749) );
  IV U23781 ( .A(n22747), .Z(n22758) );
  XOR U23782 ( .A(n22759), .B(n22760), .Z(n22747) );
  AND U23783 ( .A(n22761), .B(n22762), .Z(n22760) );
  XNOR U23784 ( .A(n22759), .B(n11382), .Z(n22762) );
  XNOR U23785 ( .A(n22755), .B(n22757), .Z(n11382) );
  NAND U23786 ( .A(n22763), .B(e_input[153]), .Z(n22757) );
  NAND U23787 ( .A(n12323), .B(e_input[153]), .Z(n22763) );
  XNOR U23788 ( .A(n22753), .B(n22764), .Z(n22755) );
  XOR U23789 ( .A(n22765), .B(n22766), .Z(n22753) );
  AND U23790 ( .A(n22767), .B(n22768), .Z(n22766) );
  XNOR U23791 ( .A(n22769), .B(n22765), .Z(n22768) );
  XOR U23792 ( .A(n22770), .B(e_input[153]), .Z(n22761) );
  IV U23793 ( .A(n22759), .Z(n22770) );
  XOR U23794 ( .A(n22771), .B(n22772), .Z(n22759) );
  AND U23795 ( .A(n22773), .B(n22774), .Z(n22772) );
  XNOR U23796 ( .A(n22771), .B(n11388), .Z(n22774) );
  XNOR U23797 ( .A(n22767), .B(n22769), .Z(n11388) );
  NAND U23798 ( .A(n22775), .B(e_input[152]), .Z(n22769) );
  NAND U23799 ( .A(n12323), .B(e_input[152]), .Z(n22775) );
  XNOR U23800 ( .A(n22765), .B(n22776), .Z(n22767) );
  XOR U23801 ( .A(n22777), .B(n22778), .Z(n22765) );
  AND U23802 ( .A(n22779), .B(n22780), .Z(n22778) );
  XNOR U23803 ( .A(n22781), .B(n22777), .Z(n22780) );
  XOR U23804 ( .A(n22782), .B(e_input[152]), .Z(n22773) );
  IV U23805 ( .A(n22771), .Z(n22782) );
  XOR U23806 ( .A(n22783), .B(n22784), .Z(n22771) );
  AND U23807 ( .A(n22785), .B(n22786), .Z(n22784) );
  XNOR U23808 ( .A(n22783), .B(n11394), .Z(n22786) );
  XNOR U23809 ( .A(n22779), .B(n22781), .Z(n11394) );
  NAND U23810 ( .A(n22787), .B(e_input[151]), .Z(n22781) );
  NAND U23811 ( .A(n12323), .B(e_input[151]), .Z(n22787) );
  XNOR U23812 ( .A(n22777), .B(n22788), .Z(n22779) );
  XOR U23813 ( .A(n22789), .B(n22790), .Z(n22777) );
  AND U23814 ( .A(n22791), .B(n22792), .Z(n22790) );
  XNOR U23815 ( .A(n22793), .B(n22789), .Z(n22792) );
  XOR U23816 ( .A(n22794), .B(e_input[151]), .Z(n22785) );
  IV U23817 ( .A(n22783), .Z(n22794) );
  XOR U23818 ( .A(n22795), .B(n22796), .Z(n22783) );
  AND U23819 ( .A(n22797), .B(n22798), .Z(n22796) );
  XNOR U23820 ( .A(n22795), .B(n11400), .Z(n22798) );
  XNOR U23821 ( .A(n22791), .B(n22793), .Z(n11400) );
  NAND U23822 ( .A(n22799), .B(e_input[150]), .Z(n22793) );
  NAND U23823 ( .A(n12323), .B(e_input[150]), .Z(n22799) );
  XNOR U23824 ( .A(n22789), .B(n22800), .Z(n22791) );
  XOR U23825 ( .A(n22801), .B(n22802), .Z(n22789) );
  AND U23826 ( .A(n22803), .B(n22804), .Z(n22802) );
  XNOR U23827 ( .A(n22805), .B(n22801), .Z(n22804) );
  XOR U23828 ( .A(n22806), .B(e_input[150]), .Z(n22797) );
  IV U23829 ( .A(n22795), .Z(n22806) );
  XOR U23830 ( .A(n22807), .B(n22808), .Z(n22795) );
  AND U23831 ( .A(n22809), .B(n22810), .Z(n22808) );
  XNOR U23832 ( .A(n22807), .B(n11406), .Z(n22810) );
  XNOR U23833 ( .A(n22803), .B(n22805), .Z(n11406) );
  NAND U23834 ( .A(n22811), .B(e_input[149]), .Z(n22805) );
  NAND U23835 ( .A(n12323), .B(e_input[149]), .Z(n22811) );
  XNOR U23836 ( .A(n22801), .B(n22812), .Z(n22803) );
  XOR U23837 ( .A(n22813), .B(n22814), .Z(n22801) );
  AND U23838 ( .A(n22815), .B(n22816), .Z(n22814) );
  XNOR U23839 ( .A(n22817), .B(n22813), .Z(n22816) );
  XOR U23840 ( .A(n22818), .B(e_input[149]), .Z(n22809) );
  IV U23841 ( .A(n22807), .Z(n22818) );
  XOR U23842 ( .A(n22819), .B(n22820), .Z(n22807) );
  AND U23843 ( .A(n22821), .B(n22822), .Z(n22820) );
  XNOR U23844 ( .A(n22819), .B(n11412), .Z(n22822) );
  XNOR U23845 ( .A(n22815), .B(n22817), .Z(n11412) );
  NAND U23846 ( .A(n22823), .B(e_input[148]), .Z(n22817) );
  NAND U23847 ( .A(n12323), .B(e_input[148]), .Z(n22823) );
  XNOR U23848 ( .A(n22813), .B(n22824), .Z(n22815) );
  XOR U23849 ( .A(n22825), .B(n22826), .Z(n22813) );
  AND U23850 ( .A(n22827), .B(n22828), .Z(n22826) );
  XNOR U23851 ( .A(n22829), .B(n22825), .Z(n22828) );
  XOR U23852 ( .A(n22830), .B(e_input[148]), .Z(n22821) );
  IV U23853 ( .A(n22819), .Z(n22830) );
  XOR U23854 ( .A(n22831), .B(n22832), .Z(n22819) );
  AND U23855 ( .A(n22833), .B(n22834), .Z(n22832) );
  XNOR U23856 ( .A(n22831), .B(n11418), .Z(n22834) );
  XNOR U23857 ( .A(n22827), .B(n22829), .Z(n11418) );
  NAND U23858 ( .A(n22835), .B(e_input[147]), .Z(n22829) );
  NAND U23859 ( .A(n12323), .B(e_input[147]), .Z(n22835) );
  XNOR U23860 ( .A(n22825), .B(n22836), .Z(n22827) );
  XOR U23861 ( .A(n22837), .B(n22838), .Z(n22825) );
  AND U23862 ( .A(n22839), .B(n22840), .Z(n22838) );
  XNOR U23863 ( .A(n22841), .B(n22837), .Z(n22840) );
  XOR U23864 ( .A(n22842), .B(e_input[147]), .Z(n22833) );
  IV U23865 ( .A(n22831), .Z(n22842) );
  XOR U23866 ( .A(n22843), .B(n22844), .Z(n22831) );
  AND U23867 ( .A(n22845), .B(n22846), .Z(n22844) );
  XNOR U23868 ( .A(n22843), .B(n11424), .Z(n22846) );
  XNOR U23869 ( .A(n22839), .B(n22841), .Z(n11424) );
  NAND U23870 ( .A(n22847), .B(e_input[146]), .Z(n22841) );
  NAND U23871 ( .A(n12323), .B(e_input[146]), .Z(n22847) );
  XNOR U23872 ( .A(n22837), .B(n22848), .Z(n22839) );
  XOR U23873 ( .A(n22849), .B(n22850), .Z(n22837) );
  AND U23874 ( .A(n22851), .B(n22852), .Z(n22850) );
  XNOR U23875 ( .A(n22853), .B(n22849), .Z(n22852) );
  XOR U23876 ( .A(n22854), .B(e_input[146]), .Z(n22845) );
  IV U23877 ( .A(n22843), .Z(n22854) );
  XOR U23878 ( .A(n22855), .B(n22856), .Z(n22843) );
  AND U23879 ( .A(n22857), .B(n22858), .Z(n22856) );
  XNOR U23880 ( .A(n22855), .B(n11430), .Z(n22858) );
  XNOR U23881 ( .A(n22851), .B(n22853), .Z(n11430) );
  NAND U23882 ( .A(n22859), .B(e_input[145]), .Z(n22853) );
  NAND U23883 ( .A(n12323), .B(e_input[145]), .Z(n22859) );
  XNOR U23884 ( .A(n22849), .B(n22860), .Z(n22851) );
  XOR U23885 ( .A(n22861), .B(n22862), .Z(n22849) );
  AND U23886 ( .A(n22863), .B(n22864), .Z(n22862) );
  XNOR U23887 ( .A(n22865), .B(n22861), .Z(n22864) );
  XOR U23888 ( .A(n22866), .B(e_input[145]), .Z(n22857) );
  IV U23889 ( .A(n22855), .Z(n22866) );
  XOR U23890 ( .A(n22867), .B(n22868), .Z(n22855) );
  AND U23891 ( .A(n22869), .B(n22870), .Z(n22868) );
  XNOR U23892 ( .A(n22867), .B(n11436), .Z(n22870) );
  XNOR U23893 ( .A(n22863), .B(n22865), .Z(n11436) );
  NAND U23894 ( .A(n22871), .B(e_input[144]), .Z(n22865) );
  NAND U23895 ( .A(n12323), .B(e_input[144]), .Z(n22871) );
  XNOR U23896 ( .A(n22861), .B(n22872), .Z(n22863) );
  XOR U23897 ( .A(n22873), .B(n22874), .Z(n22861) );
  AND U23898 ( .A(n22875), .B(n22876), .Z(n22874) );
  XNOR U23899 ( .A(n22877), .B(n22873), .Z(n22876) );
  XOR U23900 ( .A(n22878), .B(e_input[144]), .Z(n22869) );
  IV U23901 ( .A(n22867), .Z(n22878) );
  XOR U23902 ( .A(n22879), .B(n22880), .Z(n22867) );
  AND U23903 ( .A(n22881), .B(n22882), .Z(n22880) );
  XNOR U23904 ( .A(n22879), .B(n11442), .Z(n22882) );
  XNOR U23905 ( .A(n22875), .B(n22877), .Z(n11442) );
  NAND U23906 ( .A(n22883), .B(e_input[143]), .Z(n22877) );
  NAND U23907 ( .A(n12323), .B(e_input[143]), .Z(n22883) );
  XNOR U23908 ( .A(n22873), .B(n22884), .Z(n22875) );
  XOR U23909 ( .A(n22885), .B(n22886), .Z(n22873) );
  AND U23910 ( .A(n22887), .B(n22888), .Z(n22886) );
  XNOR U23911 ( .A(n22889), .B(n22885), .Z(n22888) );
  XOR U23912 ( .A(n22890), .B(e_input[143]), .Z(n22881) );
  IV U23913 ( .A(n22879), .Z(n22890) );
  XOR U23914 ( .A(n22891), .B(n22892), .Z(n22879) );
  AND U23915 ( .A(n22893), .B(n22894), .Z(n22892) );
  XNOR U23916 ( .A(n22891), .B(n11448), .Z(n22894) );
  XNOR U23917 ( .A(n22887), .B(n22889), .Z(n11448) );
  NAND U23918 ( .A(n22895), .B(e_input[142]), .Z(n22889) );
  NAND U23919 ( .A(n12323), .B(e_input[142]), .Z(n22895) );
  XNOR U23920 ( .A(n22885), .B(n22896), .Z(n22887) );
  XOR U23921 ( .A(n22897), .B(n22898), .Z(n22885) );
  AND U23922 ( .A(n22899), .B(n22900), .Z(n22898) );
  XNOR U23923 ( .A(n22901), .B(n22897), .Z(n22900) );
  XOR U23924 ( .A(n22902), .B(e_input[142]), .Z(n22893) );
  IV U23925 ( .A(n22891), .Z(n22902) );
  XOR U23926 ( .A(n22903), .B(n22904), .Z(n22891) );
  AND U23927 ( .A(n22905), .B(n22906), .Z(n22904) );
  XNOR U23928 ( .A(n22903), .B(n11454), .Z(n22906) );
  XNOR U23929 ( .A(n22899), .B(n22901), .Z(n11454) );
  NAND U23930 ( .A(n22907), .B(e_input[141]), .Z(n22901) );
  NAND U23931 ( .A(n12323), .B(e_input[141]), .Z(n22907) );
  XNOR U23932 ( .A(n22897), .B(n22908), .Z(n22899) );
  XOR U23933 ( .A(n22909), .B(n22910), .Z(n22897) );
  AND U23934 ( .A(n22911), .B(n22912), .Z(n22910) );
  XNOR U23935 ( .A(n22913), .B(n22909), .Z(n22912) );
  XOR U23936 ( .A(n22914), .B(e_input[141]), .Z(n22905) );
  IV U23937 ( .A(n22903), .Z(n22914) );
  XOR U23938 ( .A(n22915), .B(n22916), .Z(n22903) );
  AND U23939 ( .A(n22917), .B(n22918), .Z(n22916) );
  XNOR U23940 ( .A(n22915), .B(n11460), .Z(n22918) );
  XNOR U23941 ( .A(n22911), .B(n22913), .Z(n11460) );
  NAND U23942 ( .A(n22919), .B(e_input[140]), .Z(n22913) );
  NAND U23943 ( .A(n12323), .B(e_input[140]), .Z(n22919) );
  XNOR U23944 ( .A(n22909), .B(n22920), .Z(n22911) );
  XOR U23945 ( .A(n22921), .B(n22922), .Z(n22909) );
  AND U23946 ( .A(n22923), .B(n22924), .Z(n22922) );
  XNOR U23947 ( .A(n22925), .B(n22921), .Z(n22924) );
  XOR U23948 ( .A(n22926), .B(e_input[140]), .Z(n22917) );
  IV U23949 ( .A(n22915), .Z(n22926) );
  XOR U23950 ( .A(n22927), .B(n22928), .Z(n22915) );
  AND U23951 ( .A(n22929), .B(n22930), .Z(n22928) );
  XNOR U23952 ( .A(n22927), .B(n11466), .Z(n22930) );
  XNOR U23953 ( .A(n22923), .B(n22925), .Z(n11466) );
  NAND U23954 ( .A(n22931), .B(e_input[139]), .Z(n22925) );
  NAND U23955 ( .A(n12323), .B(e_input[139]), .Z(n22931) );
  XNOR U23956 ( .A(n22921), .B(n22932), .Z(n22923) );
  XOR U23957 ( .A(n22933), .B(n22934), .Z(n22921) );
  AND U23958 ( .A(n22935), .B(n22936), .Z(n22934) );
  XNOR U23959 ( .A(n22937), .B(n22933), .Z(n22936) );
  XOR U23960 ( .A(n22938), .B(e_input[139]), .Z(n22929) );
  IV U23961 ( .A(n22927), .Z(n22938) );
  XOR U23962 ( .A(n22939), .B(n22940), .Z(n22927) );
  AND U23963 ( .A(n22941), .B(n22942), .Z(n22940) );
  XNOR U23964 ( .A(n22939), .B(n11472), .Z(n22942) );
  XNOR U23965 ( .A(n22935), .B(n22937), .Z(n11472) );
  NAND U23966 ( .A(n22943), .B(e_input[138]), .Z(n22937) );
  NAND U23967 ( .A(n12323), .B(e_input[138]), .Z(n22943) );
  XNOR U23968 ( .A(n22933), .B(n22944), .Z(n22935) );
  XOR U23969 ( .A(n22945), .B(n22946), .Z(n22933) );
  AND U23970 ( .A(n22947), .B(n22948), .Z(n22946) );
  XNOR U23971 ( .A(n22949), .B(n22945), .Z(n22948) );
  XOR U23972 ( .A(n22950), .B(e_input[138]), .Z(n22941) );
  IV U23973 ( .A(n22939), .Z(n22950) );
  XOR U23974 ( .A(n22951), .B(n22952), .Z(n22939) );
  AND U23975 ( .A(n22953), .B(n22954), .Z(n22952) );
  XNOR U23976 ( .A(n22951), .B(n11478), .Z(n22954) );
  XNOR U23977 ( .A(n22947), .B(n22949), .Z(n11478) );
  NAND U23978 ( .A(n22955), .B(e_input[137]), .Z(n22949) );
  NAND U23979 ( .A(n12323), .B(e_input[137]), .Z(n22955) );
  XNOR U23980 ( .A(n22945), .B(n22956), .Z(n22947) );
  XOR U23981 ( .A(n22957), .B(n22958), .Z(n22945) );
  AND U23982 ( .A(n22959), .B(n22960), .Z(n22958) );
  XNOR U23983 ( .A(n22961), .B(n22957), .Z(n22960) );
  XOR U23984 ( .A(n22962), .B(e_input[137]), .Z(n22953) );
  IV U23985 ( .A(n22951), .Z(n22962) );
  XOR U23986 ( .A(n22963), .B(n22964), .Z(n22951) );
  AND U23987 ( .A(n22965), .B(n22966), .Z(n22964) );
  XNOR U23988 ( .A(n22963), .B(n11484), .Z(n22966) );
  XNOR U23989 ( .A(n22959), .B(n22961), .Z(n11484) );
  NAND U23990 ( .A(n22967), .B(e_input[136]), .Z(n22961) );
  NAND U23991 ( .A(n12323), .B(e_input[136]), .Z(n22967) );
  XNOR U23992 ( .A(n22957), .B(n22968), .Z(n22959) );
  XOR U23993 ( .A(n22969), .B(n22970), .Z(n22957) );
  AND U23994 ( .A(n22971), .B(n22972), .Z(n22970) );
  XNOR U23995 ( .A(n22973), .B(n22969), .Z(n22972) );
  XOR U23996 ( .A(n22974), .B(e_input[136]), .Z(n22965) );
  IV U23997 ( .A(n22963), .Z(n22974) );
  XOR U23998 ( .A(n22975), .B(n22976), .Z(n22963) );
  AND U23999 ( .A(n22977), .B(n22978), .Z(n22976) );
  XNOR U24000 ( .A(n22975), .B(n11490), .Z(n22978) );
  XNOR U24001 ( .A(n22971), .B(n22973), .Z(n11490) );
  NAND U24002 ( .A(n22979), .B(e_input[135]), .Z(n22973) );
  NAND U24003 ( .A(n12323), .B(e_input[135]), .Z(n22979) );
  XNOR U24004 ( .A(n22969), .B(n22980), .Z(n22971) );
  XOR U24005 ( .A(n22981), .B(n22982), .Z(n22969) );
  AND U24006 ( .A(n22983), .B(n22984), .Z(n22982) );
  XNOR U24007 ( .A(n22985), .B(n22981), .Z(n22984) );
  XOR U24008 ( .A(n22986), .B(e_input[135]), .Z(n22977) );
  IV U24009 ( .A(n22975), .Z(n22986) );
  XOR U24010 ( .A(n22987), .B(n22988), .Z(n22975) );
  AND U24011 ( .A(n22989), .B(n22990), .Z(n22988) );
  XNOR U24012 ( .A(n22987), .B(n11496), .Z(n22990) );
  XNOR U24013 ( .A(n22983), .B(n22985), .Z(n11496) );
  NAND U24014 ( .A(n22991), .B(e_input[134]), .Z(n22985) );
  NAND U24015 ( .A(n12323), .B(e_input[134]), .Z(n22991) );
  XNOR U24016 ( .A(n22981), .B(n22992), .Z(n22983) );
  XOR U24017 ( .A(n22993), .B(n22994), .Z(n22981) );
  AND U24018 ( .A(n22995), .B(n22996), .Z(n22994) );
  XNOR U24019 ( .A(n22997), .B(n22993), .Z(n22996) );
  XOR U24020 ( .A(n22998), .B(e_input[134]), .Z(n22989) );
  IV U24021 ( .A(n22987), .Z(n22998) );
  XOR U24022 ( .A(n22999), .B(n23000), .Z(n22987) );
  AND U24023 ( .A(n23001), .B(n23002), .Z(n23000) );
  XNOR U24024 ( .A(n22999), .B(n11502), .Z(n23002) );
  XNOR U24025 ( .A(n22995), .B(n22997), .Z(n11502) );
  NAND U24026 ( .A(n23003), .B(e_input[133]), .Z(n22997) );
  NAND U24027 ( .A(n12323), .B(e_input[133]), .Z(n23003) );
  XNOR U24028 ( .A(n22993), .B(n23004), .Z(n22995) );
  XOR U24029 ( .A(n23005), .B(n23006), .Z(n22993) );
  AND U24030 ( .A(n23007), .B(n23008), .Z(n23006) );
  XNOR U24031 ( .A(n23009), .B(n23005), .Z(n23008) );
  XOR U24032 ( .A(n23010), .B(e_input[133]), .Z(n23001) );
  IV U24033 ( .A(n22999), .Z(n23010) );
  XOR U24034 ( .A(n23011), .B(n23012), .Z(n22999) );
  AND U24035 ( .A(n23013), .B(n23014), .Z(n23012) );
  XNOR U24036 ( .A(n23011), .B(n11508), .Z(n23014) );
  XNOR U24037 ( .A(n23007), .B(n23009), .Z(n11508) );
  NAND U24038 ( .A(n23015), .B(e_input[132]), .Z(n23009) );
  NAND U24039 ( .A(n12323), .B(e_input[132]), .Z(n23015) );
  XNOR U24040 ( .A(n23005), .B(n23016), .Z(n23007) );
  XOR U24041 ( .A(n23017), .B(n23018), .Z(n23005) );
  AND U24042 ( .A(n23019), .B(n23020), .Z(n23018) );
  XNOR U24043 ( .A(n23021), .B(n23017), .Z(n23020) );
  XOR U24044 ( .A(n23022), .B(e_input[132]), .Z(n23013) );
  IV U24045 ( .A(n23011), .Z(n23022) );
  XOR U24046 ( .A(n23023), .B(n23024), .Z(n23011) );
  AND U24047 ( .A(n23025), .B(n23026), .Z(n23024) );
  XNOR U24048 ( .A(n23023), .B(n11514), .Z(n23026) );
  XNOR U24049 ( .A(n23019), .B(n23021), .Z(n11514) );
  NAND U24050 ( .A(n23027), .B(e_input[131]), .Z(n23021) );
  NAND U24051 ( .A(n12323), .B(e_input[131]), .Z(n23027) );
  XNOR U24052 ( .A(n23017), .B(n23028), .Z(n23019) );
  XOR U24053 ( .A(n23029), .B(n23030), .Z(n23017) );
  AND U24054 ( .A(n23031), .B(n23032), .Z(n23030) );
  XNOR U24055 ( .A(n23033), .B(n23029), .Z(n23032) );
  XOR U24056 ( .A(n23034), .B(e_input[131]), .Z(n23025) );
  IV U24057 ( .A(n23023), .Z(n23034) );
  XOR U24058 ( .A(n23035), .B(n23036), .Z(n23023) );
  AND U24059 ( .A(n23037), .B(n23038), .Z(n23036) );
  XNOR U24060 ( .A(n23035), .B(n11520), .Z(n23038) );
  XNOR U24061 ( .A(n23031), .B(n23033), .Z(n11520) );
  NAND U24062 ( .A(n23039), .B(e_input[130]), .Z(n23033) );
  NAND U24063 ( .A(n12323), .B(e_input[130]), .Z(n23039) );
  XNOR U24064 ( .A(n23029), .B(n23040), .Z(n23031) );
  XOR U24065 ( .A(n23041), .B(n23042), .Z(n23029) );
  AND U24066 ( .A(n23043), .B(n23044), .Z(n23042) );
  XNOR U24067 ( .A(n23045), .B(n23041), .Z(n23044) );
  XOR U24068 ( .A(n23046), .B(e_input[130]), .Z(n23037) );
  IV U24069 ( .A(n23035), .Z(n23046) );
  XOR U24070 ( .A(n23047), .B(n23048), .Z(n23035) );
  AND U24071 ( .A(n23049), .B(n23050), .Z(n23048) );
  XNOR U24072 ( .A(n23047), .B(n11526), .Z(n23050) );
  XNOR U24073 ( .A(n23043), .B(n23045), .Z(n11526) );
  NAND U24074 ( .A(n23051), .B(e_input[129]), .Z(n23045) );
  NAND U24075 ( .A(n12323), .B(e_input[129]), .Z(n23051) );
  XNOR U24076 ( .A(n23041), .B(n23052), .Z(n23043) );
  XOR U24077 ( .A(n23053), .B(n23054), .Z(n23041) );
  AND U24078 ( .A(n23055), .B(n23056), .Z(n23054) );
  XNOR U24079 ( .A(n23057), .B(n23053), .Z(n23056) );
  XOR U24080 ( .A(n23058), .B(e_input[129]), .Z(n23049) );
  IV U24081 ( .A(n23047), .Z(n23058) );
  XOR U24082 ( .A(n23059), .B(n23060), .Z(n23047) );
  AND U24083 ( .A(n23061), .B(n23062), .Z(n23060) );
  XNOR U24084 ( .A(n23059), .B(n11532), .Z(n23062) );
  XNOR U24085 ( .A(n23055), .B(n23057), .Z(n11532) );
  NAND U24086 ( .A(n23063), .B(e_input[128]), .Z(n23057) );
  NAND U24087 ( .A(n12323), .B(e_input[128]), .Z(n23063) );
  XNOR U24088 ( .A(n23053), .B(n23064), .Z(n23055) );
  XOR U24089 ( .A(n23065), .B(n23066), .Z(n23053) );
  AND U24090 ( .A(n23067), .B(n23068), .Z(n23066) );
  XNOR U24091 ( .A(n23069), .B(n23065), .Z(n23068) );
  XOR U24092 ( .A(n23070), .B(e_input[128]), .Z(n23061) );
  IV U24093 ( .A(n23059), .Z(n23070) );
  XOR U24094 ( .A(n23071), .B(n23072), .Z(n23059) );
  AND U24095 ( .A(n23073), .B(n23074), .Z(n23072) );
  XNOR U24096 ( .A(n23071), .B(n11538), .Z(n23074) );
  XNOR U24097 ( .A(n23067), .B(n23069), .Z(n11538) );
  NAND U24098 ( .A(n23075), .B(e_input[127]), .Z(n23069) );
  NAND U24099 ( .A(n12323), .B(e_input[127]), .Z(n23075) );
  XNOR U24100 ( .A(n23065), .B(n23076), .Z(n23067) );
  XOR U24101 ( .A(n23077), .B(n23078), .Z(n23065) );
  AND U24102 ( .A(n23079), .B(n23080), .Z(n23078) );
  XNOR U24103 ( .A(n23081), .B(n23077), .Z(n23080) );
  XOR U24104 ( .A(n23082), .B(e_input[127]), .Z(n23073) );
  IV U24105 ( .A(n23071), .Z(n23082) );
  XOR U24106 ( .A(n23083), .B(n23084), .Z(n23071) );
  AND U24107 ( .A(n23085), .B(n23086), .Z(n23084) );
  XNOR U24108 ( .A(n23083), .B(n11544), .Z(n23086) );
  XNOR U24109 ( .A(n23079), .B(n23081), .Z(n11544) );
  NAND U24110 ( .A(n23087), .B(e_input[126]), .Z(n23081) );
  NAND U24111 ( .A(n12323), .B(e_input[126]), .Z(n23087) );
  XNOR U24112 ( .A(n23077), .B(n23088), .Z(n23079) );
  XOR U24113 ( .A(n23089), .B(n23090), .Z(n23077) );
  AND U24114 ( .A(n23091), .B(n23092), .Z(n23090) );
  XNOR U24115 ( .A(n23093), .B(n23089), .Z(n23092) );
  XOR U24116 ( .A(n23094), .B(e_input[126]), .Z(n23085) );
  IV U24117 ( .A(n23083), .Z(n23094) );
  XOR U24118 ( .A(n23095), .B(n23096), .Z(n23083) );
  AND U24119 ( .A(n23097), .B(n23098), .Z(n23096) );
  XNOR U24120 ( .A(n23095), .B(n11550), .Z(n23098) );
  XNOR U24121 ( .A(n23091), .B(n23093), .Z(n11550) );
  NAND U24122 ( .A(n23099), .B(e_input[125]), .Z(n23093) );
  NAND U24123 ( .A(n12323), .B(e_input[125]), .Z(n23099) );
  XNOR U24124 ( .A(n23089), .B(n23100), .Z(n23091) );
  XOR U24125 ( .A(n23101), .B(n23102), .Z(n23089) );
  AND U24126 ( .A(n23103), .B(n23104), .Z(n23102) );
  XNOR U24127 ( .A(n23105), .B(n23101), .Z(n23104) );
  XOR U24128 ( .A(n23106), .B(e_input[125]), .Z(n23097) );
  IV U24129 ( .A(n23095), .Z(n23106) );
  XOR U24130 ( .A(n23107), .B(n23108), .Z(n23095) );
  AND U24131 ( .A(n23109), .B(n23110), .Z(n23108) );
  XNOR U24132 ( .A(n23107), .B(n11556), .Z(n23110) );
  XNOR U24133 ( .A(n23103), .B(n23105), .Z(n11556) );
  NAND U24134 ( .A(n23111), .B(e_input[124]), .Z(n23105) );
  NAND U24135 ( .A(n12323), .B(e_input[124]), .Z(n23111) );
  XNOR U24136 ( .A(n23101), .B(n23112), .Z(n23103) );
  XOR U24137 ( .A(n23113), .B(n23114), .Z(n23101) );
  AND U24138 ( .A(n23115), .B(n23116), .Z(n23114) );
  XNOR U24139 ( .A(n23117), .B(n23113), .Z(n23116) );
  XOR U24140 ( .A(n23118), .B(e_input[124]), .Z(n23109) );
  IV U24141 ( .A(n23107), .Z(n23118) );
  XOR U24142 ( .A(n23119), .B(n23120), .Z(n23107) );
  AND U24143 ( .A(n23121), .B(n23122), .Z(n23120) );
  XNOR U24144 ( .A(n23119), .B(n11562), .Z(n23122) );
  XNOR U24145 ( .A(n23115), .B(n23117), .Z(n11562) );
  NAND U24146 ( .A(n23123), .B(e_input[123]), .Z(n23117) );
  NAND U24147 ( .A(n12323), .B(e_input[123]), .Z(n23123) );
  XNOR U24148 ( .A(n23113), .B(n23124), .Z(n23115) );
  XOR U24149 ( .A(n23125), .B(n23126), .Z(n23113) );
  AND U24150 ( .A(n23127), .B(n23128), .Z(n23126) );
  XNOR U24151 ( .A(n23129), .B(n23125), .Z(n23128) );
  XOR U24152 ( .A(n23130), .B(e_input[123]), .Z(n23121) );
  IV U24153 ( .A(n23119), .Z(n23130) );
  XOR U24154 ( .A(n23131), .B(n23132), .Z(n23119) );
  AND U24155 ( .A(n23133), .B(n23134), .Z(n23132) );
  XNOR U24156 ( .A(n23131), .B(n11568), .Z(n23134) );
  XNOR U24157 ( .A(n23127), .B(n23129), .Z(n11568) );
  NAND U24158 ( .A(n23135), .B(e_input[122]), .Z(n23129) );
  NAND U24159 ( .A(n12323), .B(e_input[122]), .Z(n23135) );
  XNOR U24160 ( .A(n23125), .B(n23136), .Z(n23127) );
  XOR U24161 ( .A(n23137), .B(n23138), .Z(n23125) );
  AND U24162 ( .A(n23139), .B(n23140), .Z(n23138) );
  XNOR U24163 ( .A(n23141), .B(n23137), .Z(n23140) );
  XOR U24164 ( .A(n23142), .B(e_input[122]), .Z(n23133) );
  IV U24165 ( .A(n23131), .Z(n23142) );
  XOR U24166 ( .A(n23143), .B(n23144), .Z(n23131) );
  AND U24167 ( .A(n23145), .B(n23146), .Z(n23144) );
  XNOR U24168 ( .A(n23143), .B(n11574), .Z(n23146) );
  XNOR U24169 ( .A(n23139), .B(n23141), .Z(n11574) );
  NAND U24170 ( .A(n23147), .B(e_input[121]), .Z(n23141) );
  NAND U24171 ( .A(n12323), .B(e_input[121]), .Z(n23147) );
  XNOR U24172 ( .A(n23137), .B(n23148), .Z(n23139) );
  XOR U24173 ( .A(n23149), .B(n23150), .Z(n23137) );
  AND U24174 ( .A(n23151), .B(n23152), .Z(n23150) );
  XNOR U24175 ( .A(n23153), .B(n23149), .Z(n23152) );
  XOR U24176 ( .A(n23154), .B(e_input[121]), .Z(n23145) );
  IV U24177 ( .A(n23143), .Z(n23154) );
  XOR U24178 ( .A(n23155), .B(n23156), .Z(n23143) );
  AND U24179 ( .A(n23157), .B(n23158), .Z(n23156) );
  XNOR U24180 ( .A(n23155), .B(n11580), .Z(n23158) );
  XNOR U24181 ( .A(n23151), .B(n23153), .Z(n11580) );
  NAND U24182 ( .A(n23159), .B(e_input[120]), .Z(n23153) );
  NAND U24183 ( .A(n12323), .B(e_input[120]), .Z(n23159) );
  XNOR U24184 ( .A(n23149), .B(n23160), .Z(n23151) );
  XOR U24185 ( .A(n23161), .B(n23162), .Z(n23149) );
  AND U24186 ( .A(n23163), .B(n23164), .Z(n23162) );
  XNOR U24187 ( .A(n23165), .B(n23161), .Z(n23164) );
  XOR U24188 ( .A(n23166), .B(e_input[120]), .Z(n23157) );
  IV U24189 ( .A(n23155), .Z(n23166) );
  XOR U24190 ( .A(n23167), .B(n23168), .Z(n23155) );
  AND U24191 ( .A(n23169), .B(n23170), .Z(n23168) );
  XNOR U24192 ( .A(n23167), .B(n11586), .Z(n23170) );
  XNOR U24193 ( .A(n23163), .B(n23165), .Z(n11586) );
  NAND U24194 ( .A(n23171), .B(e_input[119]), .Z(n23165) );
  NAND U24195 ( .A(n12323), .B(e_input[119]), .Z(n23171) );
  XNOR U24196 ( .A(n23161), .B(n23172), .Z(n23163) );
  XOR U24197 ( .A(n23173), .B(n23174), .Z(n23161) );
  AND U24198 ( .A(n23175), .B(n23176), .Z(n23174) );
  XNOR U24199 ( .A(n23177), .B(n23173), .Z(n23176) );
  XOR U24200 ( .A(n23178), .B(e_input[119]), .Z(n23169) );
  IV U24201 ( .A(n23167), .Z(n23178) );
  XOR U24202 ( .A(n23179), .B(n23180), .Z(n23167) );
  AND U24203 ( .A(n23181), .B(n23182), .Z(n23180) );
  XNOR U24204 ( .A(n23179), .B(n11592), .Z(n23182) );
  XNOR U24205 ( .A(n23175), .B(n23177), .Z(n11592) );
  NAND U24206 ( .A(n23183), .B(e_input[118]), .Z(n23177) );
  NAND U24207 ( .A(n12323), .B(e_input[118]), .Z(n23183) );
  XNOR U24208 ( .A(n23173), .B(n23184), .Z(n23175) );
  XOR U24209 ( .A(n23185), .B(n23186), .Z(n23173) );
  AND U24210 ( .A(n23187), .B(n23188), .Z(n23186) );
  XNOR U24211 ( .A(n23189), .B(n23185), .Z(n23188) );
  XOR U24212 ( .A(n23190), .B(e_input[118]), .Z(n23181) );
  IV U24213 ( .A(n23179), .Z(n23190) );
  XOR U24214 ( .A(n23191), .B(n23192), .Z(n23179) );
  AND U24215 ( .A(n23193), .B(n23194), .Z(n23192) );
  XNOR U24216 ( .A(n23191), .B(n11598), .Z(n23194) );
  XNOR U24217 ( .A(n23187), .B(n23189), .Z(n11598) );
  NAND U24218 ( .A(n23195), .B(e_input[117]), .Z(n23189) );
  NAND U24219 ( .A(n12323), .B(e_input[117]), .Z(n23195) );
  XNOR U24220 ( .A(n23185), .B(n23196), .Z(n23187) );
  XOR U24221 ( .A(n23197), .B(n23198), .Z(n23185) );
  AND U24222 ( .A(n23199), .B(n23200), .Z(n23198) );
  XNOR U24223 ( .A(n23201), .B(n23197), .Z(n23200) );
  XOR U24224 ( .A(n23202), .B(e_input[117]), .Z(n23193) );
  IV U24225 ( .A(n23191), .Z(n23202) );
  XOR U24226 ( .A(n23203), .B(n23204), .Z(n23191) );
  AND U24227 ( .A(n23205), .B(n23206), .Z(n23204) );
  XNOR U24228 ( .A(n23203), .B(n11604), .Z(n23206) );
  XNOR U24229 ( .A(n23199), .B(n23201), .Z(n11604) );
  NAND U24230 ( .A(n23207), .B(e_input[116]), .Z(n23201) );
  NAND U24231 ( .A(n12323), .B(e_input[116]), .Z(n23207) );
  XNOR U24232 ( .A(n23197), .B(n23208), .Z(n23199) );
  XOR U24233 ( .A(n23209), .B(n23210), .Z(n23197) );
  AND U24234 ( .A(n23211), .B(n23212), .Z(n23210) );
  XNOR U24235 ( .A(n23213), .B(n23209), .Z(n23212) );
  XOR U24236 ( .A(n23214), .B(e_input[116]), .Z(n23205) );
  IV U24237 ( .A(n23203), .Z(n23214) );
  XOR U24238 ( .A(n23215), .B(n23216), .Z(n23203) );
  AND U24239 ( .A(n23217), .B(n23218), .Z(n23216) );
  XNOR U24240 ( .A(n23215), .B(n11610), .Z(n23218) );
  XNOR U24241 ( .A(n23211), .B(n23213), .Z(n11610) );
  NAND U24242 ( .A(n23219), .B(e_input[115]), .Z(n23213) );
  NAND U24243 ( .A(n12323), .B(e_input[115]), .Z(n23219) );
  XNOR U24244 ( .A(n23209), .B(n23220), .Z(n23211) );
  XOR U24245 ( .A(n23221), .B(n23222), .Z(n23209) );
  AND U24246 ( .A(n23223), .B(n23224), .Z(n23222) );
  XNOR U24247 ( .A(n23225), .B(n23221), .Z(n23224) );
  XOR U24248 ( .A(n23226), .B(e_input[115]), .Z(n23217) );
  IV U24249 ( .A(n23215), .Z(n23226) );
  XOR U24250 ( .A(n23227), .B(n23228), .Z(n23215) );
  AND U24251 ( .A(n23229), .B(n23230), .Z(n23228) );
  XNOR U24252 ( .A(n23227), .B(n11616), .Z(n23230) );
  XNOR U24253 ( .A(n23223), .B(n23225), .Z(n11616) );
  NAND U24254 ( .A(n23231), .B(e_input[114]), .Z(n23225) );
  NAND U24255 ( .A(n12323), .B(e_input[114]), .Z(n23231) );
  XNOR U24256 ( .A(n23221), .B(n23232), .Z(n23223) );
  XOR U24257 ( .A(n23233), .B(n23234), .Z(n23221) );
  AND U24258 ( .A(n23235), .B(n23236), .Z(n23234) );
  XNOR U24259 ( .A(n23237), .B(n23233), .Z(n23236) );
  XOR U24260 ( .A(n23238), .B(e_input[114]), .Z(n23229) );
  IV U24261 ( .A(n23227), .Z(n23238) );
  XOR U24262 ( .A(n23239), .B(n23240), .Z(n23227) );
  AND U24263 ( .A(n23241), .B(n23242), .Z(n23240) );
  XNOR U24264 ( .A(n23239), .B(n11622), .Z(n23242) );
  XNOR U24265 ( .A(n23235), .B(n23237), .Z(n11622) );
  NAND U24266 ( .A(n23243), .B(e_input[113]), .Z(n23237) );
  NAND U24267 ( .A(n12323), .B(e_input[113]), .Z(n23243) );
  XNOR U24268 ( .A(n23233), .B(n23244), .Z(n23235) );
  XOR U24269 ( .A(n23245), .B(n23246), .Z(n23233) );
  AND U24270 ( .A(n23247), .B(n23248), .Z(n23246) );
  XNOR U24271 ( .A(n23249), .B(n23245), .Z(n23248) );
  XOR U24272 ( .A(n23250), .B(e_input[113]), .Z(n23241) );
  IV U24273 ( .A(n23239), .Z(n23250) );
  XOR U24274 ( .A(n23251), .B(n23252), .Z(n23239) );
  AND U24275 ( .A(n23253), .B(n23254), .Z(n23252) );
  XNOR U24276 ( .A(n23251), .B(n11628), .Z(n23254) );
  XNOR U24277 ( .A(n23247), .B(n23249), .Z(n11628) );
  NAND U24278 ( .A(n23255), .B(e_input[112]), .Z(n23249) );
  NAND U24279 ( .A(n12323), .B(e_input[112]), .Z(n23255) );
  XNOR U24280 ( .A(n23245), .B(n23256), .Z(n23247) );
  XOR U24281 ( .A(n23257), .B(n23258), .Z(n23245) );
  AND U24282 ( .A(n23259), .B(n23260), .Z(n23258) );
  XNOR U24283 ( .A(n23261), .B(n23257), .Z(n23260) );
  XOR U24284 ( .A(n23262), .B(e_input[112]), .Z(n23253) );
  IV U24285 ( .A(n23251), .Z(n23262) );
  XOR U24286 ( .A(n23263), .B(n23264), .Z(n23251) );
  AND U24287 ( .A(n23265), .B(n23266), .Z(n23264) );
  XNOR U24288 ( .A(n23263), .B(n11634), .Z(n23266) );
  XNOR U24289 ( .A(n23259), .B(n23261), .Z(n11634) );
  NAND U24290 ( .A(n23267), .B(e_input[111]), .Z(n23261) );
  NAND U24291 ( .A(n12323), .B(e_input[111]), .Z(n23267) );
  XNOR U24292 ( .A(n23257), .B(n23268), .Z(n23259) );
  XOR U24293 ( .A(n23269), .B(n23270), .Z(n23257) );
  AND U24294 ( .A(n23271), .B(n23272), .Z(n23270) );
  XNOR U24295 ( .A(n23273), .B(n23269), .Z(n23272) );
  XOR U24296 ( .A(n23274), .B(e_input[111]), .Z(n23265) );
  IV U24297 ( .A(n23263), .Z(n23274) );
  XOR U24298 ( .A(n23275), .B(n23276), .Z(n23263) );
  AND U24299 ( .A(n23277), .B(n23278), .Z(n23276) );
  XNOR U24300 ( .A(n23275), .B(n11640), .Z(n23278) );
  XNOR U24301 ( .A(n23271), .B(n23273), .Z(n11640) );
  NAND U24302 ( .A(n23279), .B(e_input[110]), .Z(n23273) );
  NAND U24303 ( .A(n12323), .B(e_input[110]), .Z(n23279) );
  XNOR U24304 ( .A(n23269), .B(n23280), .Z(n23271) );
  XOR U24305 ( .A(n23281), .B(n23282), .Z(n23269) );
  AND U24306 ( .A(n23283), .B(n23284), .Z(n23282) );
  XNOR U24307 ( .A(n23285), .B(n23281), .Z(n23284) );
  XOR U24308 ( .A(n23286), .B(e_input[110]), .Z(n23277) );
  IV U24309 ( .A(n23275), .Z(n23286) );
  XOR U24310 ( .A(n23287), .B(n23288), .Z(n23275) );
  AND U24311 ( .A(n23289), .B(n23290), .Z(n23288) );
  XNOR U24312 ( .A(n23287), .B(n11646), .Z(n23290) );
  XNOR U24313 ( .A(n23283), .B(n23285), .Z(n11646) );
  NAND U24314 ( .A(n23291), .B(e_input[109]), .Z(n23285) );
  NAND U24315 ( .A(n12323), .B(e_input[109]), .Z(n23291) );
  XNOR U24316 ( .A(n23281), .B(n23292), .Z(n23283) );
  XOR U24317 ( .A(n23293), .B(n23294), .Z(n23281) );
  AND U24318 ( .A(n23295), .B(n23296), .Z(n23294) );
  XNOR U24319 ( .A(n23297), .B(n23293), .Z(n23296) );
  XOR U24320 ( .A(n23298), .B(e_input[109]), .Z(n23289) );
  IV U24321 ( .A(n23287), .Z(n23298) );
  XOR U24322 ( .A(n23299), .B(n23300), .Z(n23287) );
  AND U24323 ( .A(n23301), .B(n23302), .Z(n23300) );
  XNOR U24324 ( .A(n23299), .B(n11652), .Z(n23302) );
  XNOR U24325 ( .A(n23295), .B(n23297), .Z(n11652) );
  NAND U24326 ( .A(n23303), .B(e_input[108]), .Z(n23297) );
  NAND U24327 ( .A(n12323), .B(e_input[108]), .Z(n23303) );
  XNOR U24328 ( .A(n23293), .B(n23304), .Z(n23295) );
  XOR U24329 ( .A(n23305), .B(n23306), .Z(n23293) );
  AND U24330 ( .A(n23307), .B(n23308), .Z(n23306) );
  XNOR U24331 ( .A(n23309), .B(n23305), .Z(n23308) );
  XOR U24332 ( .A(n23310), .B(e_input[108]), .Z(n23301) );
  IV U24333 ( .A(n23299), .Z(n23310) );
  XOR U24334 ( .A(n23311), .B(n23312), .Z(n23299) );
  AND U24335 ( .A(n23313), .B(n23314), .Z(n23312) );
  XNOR U24336 ( .A(n23311), .B(n11658), .Z(n23314) );
  XNOR U24337 ( .A(n23307), .B(n23309), .Z(n11658) );
  NAND U24338 ( .A(n23315), .B(e_input[107]), .Z(n23309) );
  NAND U24339 ( .A(n12323), .B(e_input[107]), .Z(n23315) );
  XNOR U24340 ( .A(n23305), .B(n23316), .Z(n23307) );
  XOR U24341 ( .A(n23317), .B(n23318), .Z(n23305) );
  AND U24342 ( .A(n23319), .B(n23320), .Z(n23318) );
  XNOR U24343 ( .A(n23321), .B(n23317), .Z(n23320) );
  XOR U24344 ( .A(n23322), .B(e_input[107]), .Z(n23313) );
  IV U24345 ( .A(n23311), .Z(n23322) );
  XOR U24346 ( .A(n23323), .B(n23324), .Z(n23311) );
  AND U24347 ( .A(n23325), .B(n23326), .Z(n23324) );
  XNOR U24348 ( .A(n23323), .B(n11664), .Z(n23326) );
  XNOR U24349 ( .A(n23319), .B(n23321), .Z(n11664) );
  NAND U24350 ( .A(n23327), .B(e_input[106]), .Z(n23321) );
  NAND U24351 ( .A(n12323), .B(e_input[106]), .Z(n23327) );
  XNOR U24352 ( .A(n23317), .B(n23328), .Z(n23319) );
  XOR U24353 ( .A(n23329), .B(n23330), .Z(n23317) );
  AND U24354 ( .A(n23331), .B(n23332), .Z(n23330) );
  XNOR U24355 ( .A(n23333), .B(n23329), .Z(n23332) );
  XOR U24356 ( .A(n23334), .B(e_input[106]), .Z(n23325) );
  IV U24357 ( .A(n23323), .Z(n23334) );
  XOR U24358 ( .A(n23335), .B(n23336), .Z(n23323) );
  AND U24359 ( .A(n23337), .B(n23338), .Z(n23336) );
  XNOR U24360 ( .A(n23335), .B(n11670), .Z(n23338) );
  XNOR U24361 ( .A(n23331), .B(n23333), .Z(n11670) );
  NAND U24362 ( .A(n23339), .B(e_input[105]), .Z(n23333) );
  NAND U24363 ( .A(n12323), .B(e_input[105]), .Z(n23339) );
  XNOR U24364 ( .A(n23329), .B(n23340), .Z(n23331) );
  XOR U24365 ( .A(n23341), .B(n23342), .Z(n23329) );
  AND U24366 ( .A(n23343), .B(n23344), .Z(n23342) );
  XNOR U24367 ( .A(n23345), .B(n23341), .Z(n23344) );
  XOR U24368 ( .A(n23346), .B(e_input[105]), .Z(n23337) );
  IV U24369 ( .A(n23335), .Z(n23346) );
  XOR U24370 ( .A(n23347), .B(n23348), .Z(n23335) );
  AND U24371 ( .A(n23349), .B(n23350), .Z(n23348) );
  XNOR U24372 ( .A(n23347), .B(n11676), .Z(n23350) );
  XNOR U24373 ( .A(n23343), .B(n23345), .Z(n11676) );
  NAND U24374 ( .A(n23351), .B(e_input[104]), .Z(n23345) );
  NAND U24375 ( .A(n12323), .B(e_input[104]), .Z(n23351) );
  XNOR U24376 ( .A(n23341), .B(n23352), .Z(n23343) );
  XOR U24377 ( .A(n23353), .B(n23354), .Z(n23341) );
  AND U24378 ( .A(n23355), .B(n23356), .Z(n23354) );
  XNOR U24379 ( .A(n23357), .B(n23353), .Z(n23356) );
  XOR U24380 ( .A(n23358), .B(e_input[104]), .Z(n23349) );
  IV U24381 ( .A(n23347), .Z(n23358) );
  XOR U24382 ( .A(n23359), .B(n23360), .Z(n23347) );
  AND U24383 ( .A(n23361), .B(n23362), .Z(n23360) );
  XNOR U24384 ( .A(n23359), .B(n11682), .Z(n23362) );
  XNOR U24385 ( .A(n23355), .B(n23357), .Z(n11682) );
  NAND U24386 ( .A(n23363), .B(e_input[103]), .Z(n23357) );
  NAND U24387 ( .A(n12323), .B(e_input[103]), .Z(n23363) );
  XNOR U24388 ( .A(n23353), .B(n23364), .Z(n23355) );
  XOR U24389 ( .A(n23365), .B(n23366), .Z(n23353) );
  AND U24390 ( .A(n23367), .B(n23368), .Z(n23366) );
  XNOR U24391 ( .A(n23369), .B(n23365), .Z(n23368) );
  XOR U24392 ( .A(n23370), .B(e_input[103]), .Z(n23361) );
  IV U24393 ( .A(n23359), .Z(n23370) );
  XOR U24394 ( .A(n23371), .B(n23372), .Z(n23359) );
  AND U24395 ( .A(n23373), .B(n23374), .Z(n23372) );
  XNOR U24396 ( .A(n23371), .B(n11688), .Z(n23374) );
  XNOR U24397 ( .A(n23367), .B(n23369), .Z(n11688) );
  NAND U24398 ( .A(n23375), .B(e_input[102]), .Z(n23369) );
  NAND U24399 ( .A(n12323), .B(e_input[102]), .Z(n23375) );
  XNOR U24400 ( .A(n23365), .B(n23376), .Z(n23367) );
  XOR U24401 ( .A(n23377), .B(n23378), .Z(n23365) );
  AND U24402 ( .A(n23379), .B(n23380), .Z(n23378) );
  XNOR U24403 ( .A(n23381), .B(n23377), .Z(n23380) );
  XOR U24404 ( .A(n23382), .B(e_input[102]), .Z(n23373) );
  IV U24405 ( .A(n23371), .Z(n23382) );
  XOR U24406 ( .A(n23383), .B(n23384), .Z(n23371) );
  AND U24407 ( .A(n23385), .B(n23386), .Z(n23384) );
  XNOR U24408 ( .A(n23383), .B(n11694), .Z(n23386) );
  XNOR U24409 ( .A(n23379), .B(n23381), .Z(n11694) );
  NAND U24410 ( .A(n23387), .B(e_input[101]), .Z(n23381) );
  NAND U24411 ( .A(n12323), .B(e_input[101]), .Z(n23387) );
  XNOR U24412 ( .A(n23377), .B(n23388), .Z(n23379) );
  XOR U24413 ( .A(n23389), .B(n23390), .Z(n23377) );
  AND U24414 ( .A(n23391), .B(n23392), .Z(n23390) );
  XNOR U24415 ( .A(n23393), .B(n23389), .Z(n23392) );
  XOR U24416 ( .A(n23394), .B(e_input[101]), .Z(n23385) );
  IV U24417 ( .A(n23383), .Z(n23394) );
  XOR U24418 ( .A(n23395), .B(n23396), .Z(n23383) );
  AND U24419 ( .A(n23397), .B(n23398), .Z(n23396) );
  XNOR U24420 ( .A(n23395), .B(n11700), .Z(n23398) );
  XNOR U24421 ( .A(n23391), .B(n23393), .Z(n11700) );
  NAND U24422 ( .A(n23399), .B(e_input[100]), .Z(n23393) );
  NAND U24423 ( .A(n12323), .B(e_input[100]), .Z(n23399) );
  XNOR U24424 ( .A(n23389), .B(n23400), .Z(n23391) );
  XOR U24425 ( .A(n23401), .B(n23402), .Z(n23389) );
  AND U24426 ( .A(n23403), .B(n23404), .Z(n23402) );
  XNOR U24427 ( .A(n23405), .B(n23401), .Z(n23404) );
  XOR U24428 ( .A(n23406), .B(e_input[100]), .Z(n23397) );
  IV U24429 ( .A(n23395), .Z(n23406) );
  XOR U24430 ( .A(n23407), .B(n23408), .Z(n23395) );
  AND U24431 ( .A(n23409), .B(n23410), .Z(n23408) );
  XNOR U24432 ( .A(n23407), .B(n11706), .Z(n23410) );
  XNOR U24433 ( .A(n23403), .B(n23405), .Z(n11706) );
  NAND U24434 ( .A(n23411), .B(e_input[99]), .Z(n23405) );
  NAND U24435 ( .A(n12323), .B(e_input[99]), .Z(n23411) );
  XNOR U24436 ( .A(n23401), .B(n23412), .Z(n23403) );
  XOR U24437 ( .A(n23413), .B(n23414), .Z(n23401) );
  AND U24438 ( .A(n23415), .B(n23416), .Z(n23414) );
  XNOR U24439 ( .A(n23417), .B(n23413), .Z(n23416) );
  XOR U24440 ( .A(n23418), .B(e_input[99]), .Z(n23409) );
  IV U24441 ( .A(n23407), .Z(n23418) );
  XOR U24442 ( .A(n23419), .B(n23420), .Z(n23407) );
  AND U24443 ( .A(n23421), .B(n23422), .Z(n23420) );
  XNOR U24444 ( .A(n23419), .B(n11712), .Z(n23422) );
  XNOR U24445 ( .A(n23415), .B(n23417), .Z(n11712) );
  NAND U24446 ( .A(n23423), .B(e_input[98]), .Z(n23417) );
  NAND U24447 ( .A(n12323), .B(e_input[98]), .Z(n23423) );
  XNOR U24448 ( .A(n23413), .B(n23424), .Z(n23415) );
  XOR U24449 ( .A(n23425), .B(n23426), .Z(n23413) );
  AND U24450 ( .A(n23427), .B(n23428), .Z(n23426) );
  XNOR U24451 ( .A(n23429), .B(n23425), .Z(n23428) );
  XOR U24452 ( .A(n23430), .B(e_input[98]), .Z(n23421) );
  IV U24453 ( .A(n23419), .Z(n23430) );
  XOR U24454 ( .A(n23431), .B(n23432), .Z(n23419) );
  AND U24455 ( .A(n23433), .B(n23434), .Z(n23432) );
  XNOR U24456 ( .A(n23431), .B(n11718), .Z(n23434) );
  XNOR U24457 ( .A(n23427), .B(n23429), .Z(n11718) );
  NAND U24458 ( .A(n23435), .B(e_input[97]), .Z(n23429) );
  NAND U24459 ( .A(n12323), .B(e_input[97]), .Z(n23435) );
  XNOR U24460 ( .A(n23425), .B(n23436), .Z(n23427) );
  XOR U24461 ( .A(n23437), .B(n23438), .Z(n23425) );
  AND U24462 ( .A(n23439), .B(n23440), .Z(n23438) );
  XNOR U24463 ( .A(n23441), .B(n23437), .Z(n23440) );
  XOR U24464 ( .A(n23442), .B(e_input[97]), .Z(n23433) );
  IV U24465 ( .A(n23431), .Z(n23442) );
  XOR U24466 ( .A(n23443), .B(n23444), .Z(n23431) );
  AND U24467 ( .A(n23445), .B(n23446), .Z(n23444) );
  XNOR U24468 ( .A(n23443), .B(n11724), .Z(n23446) );
  XNOR U24469 ( .A(n23439), .B(n23441), .Z(n11724) );
  NAND U24470 ( .A(n23447), .B(e_input[96]), .Z(n23441) );
  NAND U24471 ( .A(n12323), .B(e_input[96]), .Z(n23447) );
  XNOR U24472 ( .A(n23437), .B(n23448), .Z(n23439) );
  XOR U24473 ( .A(n23449), .B(n23450), .Z(n23437) );
  AND U24474 ( .A(n23451), .B(n23452), .Z(n23450) );
  XNOR U24475 ( .A(n23453), .B(n23449), .Z(n23452) );
  XOR U24476 ( .A(n23454), .B(e_input[96]), .Z(n23445) );
  IV U24477 ( .A(n23443), .Z(n23454) );
  XOR U24478 ( .A(n23455), .B(n23456), .Z(n23443) );
  AND U24479 ( .A(n23457), .B(n23458), .Z(n23456) );
  XNOR U24480 ( .A(n23455), .B(n11730), .Z(n23458) );
  XNOR U24481 ( .A(n23451), .B(n23453), .Z(n11730) );
  NAND U24482 ( .A(n23459), .B(e_input[95]), .Z(n23453) );
  NAND U24483 ( .A(n12323), .B(e_input[95]), .Z(n23459) );
  XNOR U24484 ( .A(n23449), .B(n23460), .Z(n23451) );
  XOR U24485 ( .A(n23461), .B(n23462), .Z(n23449) );
  AND U24486 ( .A(n23463), .B(n23464), .Z(n23462) );
  XNOR U24487 ( .A(n23465), .B(n23461), .Z(n23464) );
  XOR U24488 ( .A(n23466), .B(e_input[95]), .Z(n23457) );
  IV U24489 ( .A(n23455), .Z(n23466) );
  XOR U24490 ( .A(n23467), .B(n23468), .Z(n23455) );
  AND U24491 ( .A(n23469), .B(n23470), .Z(n23468) );
  XNOR U24492 ( .A(n23467), .B(n11736), .Z(n23470) );
  XNOR U24493 ( .A(n23463), .B(n23465), .Z(n11736) );
  NAND U24494 ( .A(n23471), .B(e_input[94]), .Z(n23465) );
  NAND U24495 ( .A(n12323), .B(e_input[94]), .Z(n23471) );
  XNOR U24496 ( .A(n23461), .B(n23472), .Z(n23463) );
  XOR U24497 ( .A(n23473), .B(n23474), .Z(n23461) );
  AND U24498 ( .A(n23475), .B(n23476), .Z(n23474) );
  XNOR U24499 ( .A(n23477), .B(n23473), .Z(n23476) );
  XOR U24500 ( .A(n23478), .B(e_input[94]), .Z(n23469) );
  IV U24501 ( .A(n23467), .Z(n23478) );
  XOR U24502 ( .A(n23479), .B(n23480), .Z(n23467) );
  AND U24503 ( .A(n23481), .B(n23482), .Z(n23480) );
  XNOR U24504 ( .A(n23479), .B(n11742), .Z(n23482) );
  XNOR U24505 ( .A(n23475), .B(n23477), .Z(n11742) );
  NAND U24506 ( .A(n23483), .B(e_input[93]), .Z(n23477) );
  NAND U24507 ( .A(n12323), .B(e_input[93]), .Z(n23483) );
  XNOR U24508 ( .A(n23473), .B(n23484), .Z(n23475) );
  XOR U24509 ( .A(n23485), .B(n23486), .Z(n23473) );
  AND U24510 ( .A(n23487), .B(n23488), .Z(n23486) );
  XNOR U24511 ( .A(n23489), .B(n23485), .Z(n23488) );
  XOR U24512 ( .A(n23490), .B(e_input[93]), .Z(n23481) );
  IV U24513 ( .A(n23479), .Z(n23490) );
  XOR U24514 ( .A(n23491), .B(n23492), .Z(n23479) );
  AND U24515 ( .A(n23493), .B(n23494), .Z(n23492) );
  XNOR U24516 ( .A(n23491), .B(n11748), .Z(n23494) );
  XNOR U24517 ( .A(n23487), .B(n23489), .Z(n11748) );
  NAND U24518 ( .A(n23495), .B(e_input[92]), .Z(n23489) );
  NAND U24519 ( .A(n12323), .B(e_input[92]), .Z(n23495) );
  XNOR U24520 ( .A(n23485), .B(n23496), .Z(n23487) );
  XOR U24521 ( .A(n23497), .B(n23498), .Z(n23485) );
  AND U24522 ( .A(n23499), .B(n23500), .Z(n23498) );
  XNOR U24523 ( .A(n23501), .B(n23497), .Z(n23500) );
  XOR U24524 ( .A(n23502), .B(e_input[92]), .Z(n23493) );
  IV U24525 ( .A(n23491), .Z(n23502) );
  XOR U24526 ( .A(n23503), .B(n23504), .Z(n23491) );
  AND U24527 ( .A(n23505), .B(n23506), .Z(n23504) );
  XNOR U24528 ( .A(n23503), .B(n11754), .Z(n23506) );
  XNOR U24529 ( .A(n23499), .B(n23501), .Z(n11754) );
  NAND U24530 ( .A(n23507), .B(e_input[91]), .Z(n23501) );
  NAND U24531 ( .A(n12323), .B(e_input[91]), .Z(n23507) );
  XNOR U24532 ( .A(n23497), .B(n23508), .Z(n23499) );
  XOR U24533 ( .A(n23509), .B(n23510), .Z(n23497) );
  AND U24534 ( .A(n23511), .B(n23512), .Z(n23510) );
  XNOR U24535 ( .A(n23513), .B(n23509), .Z(n23512) );
  XOR U24536 ( .A(n23514), .B(e_input[91]), .Z(n23505) );
  IV U24537 ( .A(n23503), .Z(n23514) );
  XOR U24538 ( .A(n23515), .B(n23516), .Z(n23503) );
  AND U24539 ( .A(n23517), .B(n23518), .Z(n23516) );
  XNOR U24540 ( .A(n23515), .B(n11760), .Z(n23518) );
  XNOR U24541 ( .A(n23511), .B(n23513), .Z(n11760) );
  NAND U24542 ( .A(n23519), .B(e_input[90]), .Z(n23513) );
  NAND U24543 ( .A(n12323), .B(e_input[90]), .Z(n23519) );
  XNOR U24544 ( .A(n23509), .B(n23520), .Z(n23511) );
  XOR U24545 ( .A(n23521), .B(n23522), .Z(n23509) );
  AND U24546 ( .A(n23523), .B(n23524), .Z(n23522) );
  XNOR U24547 ( .A(n23525), .B(n23521), .Z(n23524) );
  XOR U24548 ( .A(n23526), .B(e_input[90]), .Z(n23517) );
  IV U24549 ( .A(n23515), .Z(n23526) );
  XOR U24550 ( .A(n23527), .B(n23528), .Z(n23515) );
  AND U24551 ( .A(n23529), .B(n23530), .Z(n23528) );
  XNOR U24552 ( .A(n23527), .B(n11766), .Z(n23530) );
  XNOR U24553 ( .A(n23523), .B(n23525), .Z(n11766) );
  NAND U24554 ( .A(n23531), .B(e_input[89]), .Z(n23525) );
  NAND U24555 ( .A(n12323), .B(e_input[89]), .Z(n23531) );
  XNOR U24556 ( .A(n23521), .B(n23532), .Z(n23523) );
  XOR U24557 ( .A(n23533), .B(n23534), .Z(n23521) );
  AND U24558 ( .A(n23535), .B(n23536), .Z(n23534) );
  XNOR U24559 ( .A(n23537), .B(n23533), .Z(n23536) );
  XOR U24560 ( .A(n23538), .B(e_input[89]), .Z(n23529) );
  IV U24561 ( .A(n23527), .Z(n23538) );
  XOR U24562 ( .A(n23539), .B(n23540), .Z(n23527) );
  AND U24563 ( .A(n23541), .B(n23542), .Z(n23540) );
  XNOR U24564 ( .A(n23539), .B(n11772), .Z(n23542) );
  XNOR U24565 ( .A(n23535), .B(n23537), .Z(n11772) );
  NAND U24566 ( .A(n23543), .B(e_input[88]), .Z(n23537) );
  NAND U24567 ( .A(n12323), .B(e_input[88]), .Z(n23543) );
  XNOR U24568 ( .A(n23533), .B(n23544), .Z(n23535) );
  XOR U24569 ( .A(n23545), .B(n23546), .Z(n23533) );
  AND U24570 ( .A(n23547), .B(n23548), .Z(n23546) );
  XNOR U24571 ( .A(n23549), .B(n23545), .Z(n23548) );
  XOR U24572 ( .A(n23550), .B(e_input[88]), .Z(n23541) );
  IV U24573 ( .A(n23539), .Z(n23550) );
  XOR U24574 ( .A(n23551), .B(n23552), .Z(n23539) );
  AND U24575 ( .A(n23553), .B(n23554), .Z(n23552) );
  XNOR U24576 ( .A(n23551), .B(n11778), .Z(n23554) );
  XNOR U24577 ( .A(n23547), .B(n23549), .Z(n11778) );
  NAND U24578 ( .A(n23555), .B(e_input[87]), .Z(n23549) );
  NAND U24579 ( .A(n12323), .B(e_input[87]), .Z(n23555) );
  XNOR U24580 ( .A(n23545), .B(n23556), .Z(n23547) );
  XOR U24581 ( .A(n23557), .B(n23558), .Z(n23545) );
  AND U24582 ( .A(n23559), .B(n23560), .Z(n23558) );
  XNOR U24583 ( .A(n23561), .B(n23557), .Z(n23560) );
  XOR U24584 ( .A(n23562), .B(e_input[87]), .Z(n23553) );
  IV U24585 ( .A(n23551), .Z(n23562) );
  XOR U24586 ( .A(n23563), .B(n23564), .Z(n23551) );
  AND U24587 ( .A(n23565), .B(n23566), .Z(n23564) );
  XNOR U24588 ( .A(n23563), .B(n11784), .Z(n23566) );
  XNOR U24589 ( .A(n23559), .B(n23561), .Z(n11784) );
  NAND U24590 ( .A(n23567), .B(e_input[86]), .Z(n23561) );
  NAND U24591 ( .A(n12323), .B(e_input[86]), .Z(n23567) );
  XNOR U24592 ( .A(n23557), .B(n23568), .Z(n23559) );
  XOR U24593 ( .A(n23569), .B(n23570), .Z(n23557) );
  AND U24594 ( .A(n23571), .B(n23572), .Z(n23570) );
  XNOR U24595 ( .A(n23573), .B(n23569), .Z(n23572) );
  XOR U24596 ( .A(n23574), .B(e_input[86]), .Z(n23565) );
  IV U24597 ( .A(n23563), .Z(n23574) );
  XOR U24598 ( .A(n23575), .B(n23576), .Z(n23563) );
  AND U24599 ( .A(n23577), .B(n23578), .Z(n23576) );
  XNOR U24600 ( .A(n23575), .B(n11790), .Z(n23578) );
  XNOR U24601 ( .A(n23571), .B(n23573), .Z(n11790) );
  NAND U24602 ( .A(n23579), .B(e_input[85]), .Z(n23573) );
  NAND U24603 ( .A(n12323), .B(e_input[85]), .Z(n23579) );
  XNOR U24604 ( .A(n23569), .B(n23580), .Z(n23571) );
  XOR U24605 ( .A(n23581), .B(n23582), .Z(n23569) );
  AND U24606 ( .A(n23583), .B(n23584), .Z(n23582) );
  XNOR U24607 ( .A(n23585), .B(n23581), .Z(n23584) );
  XOR U24608 ( .A(n23586), .B(e_input[85]), .Z(n23577) );
  IV U24609 ( .A(n23575), .Z(n23586) );
  XOR U24610 ( .A(n23587), .B(n23588), .Z(n23575) );
  AND U24611 ( .A(n23589), .B(n23590), .Z(n23588) );
  XNOR U24612 ( .A(n23587), .B(n11796), .Z(n23590) );
  XNOR U24613 ( .A(n23583), .B(n23585), .Z(n11796) );
  NAND U24614 ( .A(n23591), .B(e_input[84]), .Z(n23585) );
  NAND U24615 ( .A(n12323), .B(e_input[84]), .Z(n23591) );
  XNOR U24616 ( .A(n23581), .B(n23592), .Z(n23583) );
  XOR U24617 ( .A(n23593), .B(n23594), .Z(n23581) );
  AND U24618 ( .A(n23595), .B(n23596), .Z(n23594) );
  XNOR U24619 ( .A(n23597), .B(n23593), .Z(n23596) );
  XOR U24620 ( .A(n23598), .B(e_input[84]), .Z(n23589) );
  IV U24621 ( .A(n23587), .Z(n23598) );
  XOR U24622 ( .A(n23599), .B(n23600), .Z(n23587) );
  AND U24623 ( .A(n23601), .B(n23602), .Z(n23600) );
  XNOR U24624 ( .A(n23599), .B(n11802), .Z(n23602) );
  XNOR U24625 ( .A(n23595), .B(n23597), .Z(n11802) );
  NAND U24626 ( .A(n23603), .B(e_input[83]), .Z(n23597) );
  NAND U24627 ( .A(n12323), .B(e_input[83]), .Z(n23603) );
  XNOR U24628 ( .A(n23593), .B(n23604), .Z(n23595) );
  XOR U24629 ( .A(n23605), .B(n23606), .Z(n23593) );
  AND U24630 ( .A(n23607), .B(n23608), .Z(n23606) );
  XNOR U24631 ( .A(n23609), .B(n23605), .Z(n23608) );
  XOR U24632 ( .A(n23610), .B(e_input[83]), .Z(n23601) );
  IV U24633 ( .A(n23599), .Z(n23610) );
  XOR U24634 ( .A(n23611), .B(n23612), .Z(n23599) );
  AND U24635 ( .A(n23613), .B(n23614), .Z(n23612) );
  XNOR U24636 ( .A(n23611), .B(n11808), .Z(n23614) );
  XNOR U24637 ( .A(n23607), .B(n23609), .Z(n11808) );
  NAND U24638 ( .A(n23615), .B(e_input[82]), .Z(n23609) );
  NAND U24639 ( .A(n12323), .B(e_input[82]), .Z(n23615) );
  XNOR U24640 ( .A(n23605), .B(n23616), .Z(n23607) );
  XOR U24641 ( .A(n23617), .B(n23618), .Z(n23605) );
  AND U24642 ( .A(n23619), .B(n23620), .Z(n23618) );
  XNOR U24643 ( .A(n23621), .B(n23617), .Z(n23620) );
  XOR U24644 ( .A(n23622), .B(e_input[82]), .Z(n23613) );
  IV U24645 ( .A(n23611), .Z(n23622) );
  XOR U24646 ( .A(n23623), .B(n23624), .Z(n23611) );
  AND U24647 ( .A(n23625), .B(n23626), .Z(n23624) );
  XNOR U24648 ( .A(n23623), .B(n11814), .Z(n23626) );
  XNOR U24649 ( .A(n23619), .B(n23621), .Z(n11814) );
  NAND U24650 ( .A(n23627), .B(e_input[81]), .Z(n23621) );
  NAND U24651 ( .A(n12323), .B(e_input[81]), .Z(n23627) );
  XNOR U24652 ( .A(n23617), .B(n23628), .Z(n23619) );
  XOR U24653 ( .A(n23629), .B(n23630), .Z(n23617) );
  AND U24654 ( .A(n23631), .B(n23632), .Z(n23630) );
  XNOR U24655 ( .A(n23633), .B(n23629), .Z(n23632) );
  XOR U24656 ( .A(n23634), .B(e_input[81]), .Z(n23625) );
  IV U24657 ( .A(n23623), .Z(n23634) );
  XOR U24658 ( .A(n23635), .B(n23636), .Z(n23623) );
  AND U24659 ( .A(n23637), .B(n23638), .Z(n23636) );
  XNOR U24660 ( .A(n23635), .B(n11820), .Z(n23638) );
  XNOR U24661 ( .A(n23631), .B(n23633), .Z(n11820) );
  NAND U24662 ( .A(n23639), .B(e_input[80]), .Z(n23633) );
  NAND U24663 ( .A(n12323), .B(e_input[80]), .Z(n23639) );
  XNOR U24664 ( .A(n23629), .B(n23640), .Z(n23631) );
  XOR U24665 ( .A(n23641), .B(n23642), .Z(n23629) );
  AND U24666 ( .A(n23643), .B(n23644), .Z(n23642) );
  XNOR U24667 ( .A(n23645), .B(n23641), .Z(n23644) );
  XOR U24668 ( .A(n23646), .B(e_input[80]), .Z(n23637) );
  IV U24669 ( .A(n23635), .Z(n23646) );
  XOR U24670 ( .A(n23647), .B(n23648), .Z(n23635) );
  AND U24671 ( .A(n23649), .B(n23650), .Z(n23648) );
  XNOR U24672 ( .A(n23647), .B(n11826), .Z(n23650) );
  XNOR U24673 ( .A(n23643), .B(n23645), .Z(n11826) );
  NAND U24674 ( .A(n23651), .B(e_input[79]), .Z(n23645) );
  NAND U24675 ( .A(n12323), .B(e_input[79]), .Z(n23651) );
  XNOR U24676 ( .A(n23641), .B(n23652), .Z(n23643) );
  XOR U24677 ( .A(n23653), .B(n23654), .Z(n23641) );
  AND U24678 ( .A(n23655), .B(n23656), .Z(n23654) );
  XNOR U24679 ( .A(n23657), .B(n23653), .Z(n23656) );
  XOR U24680 ( .A(n23658), .B(e_input[79]), .Z(n23649) );
  IV U24681 ( .A(n23647), .Z(n23658) );
  XOR U24682 ( .A(n23659), .B(n23660), .Z(n23647) );
  AND U24683 ( .A(n23661), .B(n23662), .Z(n23660) );
  XNOR U24684 ( .A(n23659), .B(n11832), .Z(n23662) );
  XNOR U24685 ( .A(n23655), .B(n23657), .Z(n11832) );
  NAND U24686 ( .A(n23663), .B(e_input[78]), .Z(n23657) );
  NAND U24687 ( .A(n12323), .B(e_input[78]), .Z(n23663) );
  XNOR U24688 ( .A(n23653), .B(n23664), .Z(n23655) );
  XOR U24689 ( .A(n23665), .B(n23666), .Z(n23653) );
  AND U24690 ( .A(n23667), .B(n23668), .Z(n23666) );
  XNOR U24691 ( .A(n23669), .B(n23665), .Z(n23668) );
  XOR U24692 ( .A(n23670), .B(e_input[78]), .Z(n23661) );
  IV U24693 ( .A(n23659), .Z(n23670) );
  XOR U24694 ( .A(n23671), .B(n23672), .Z(n23659) );
  AND U24695 ( .A(n23673), .B(n23674), .Z(n23672) );
  XNOR U24696 ( .A(n23671), .B(n11838), .Z(n23674) );
  XNOR U24697 ( .A(n23667), .B(n23669), .Z(n11838) );
  NAND U24698 ( .A(n23675), .B(e_input[77]), .Z(n23669) );
  NAND U24699 ( .A(n12323), .B(e_input[77]), .Z(n23675) );
  XNOR U24700 ( .A(n23665), .B(n23676), .Z(n23667) );
  XOR U24701 ( .A(n23677), .B(n23678), .Z(n23665) );
  AND U24702 ( .A(n23679), .B(n23680), .Z(n23678) );
  XNOR U24703 ( .A(n23681), .B(n23677), .Z(n23680) );
  XOR U24704 ( .A(n23682), .B(e_input[77]), .Z(n23673) );
  IV U24705 ( .A(n23671), .Z(n23682) );
  XOR U24706 ( .A(n23683), .B(n23684), .Z(n23671) );
  AND U24707 ( .A(n23685), .B(n23686), .Z(n23684) );
  XNOR U24708 ( .A(n23683), .B(n11844), .Z(n23686) );
  XNOR U24709 ( .A(n23679), .B(n23681), .Z(n11844) );
  NAND U24710 ( .A(n23687), .B(e_input[76]), .Z(n23681) );
  NAND U24711 ( .A(n12323), .B(e_input[76]), .Z(n23687) );
  XNOR U24712 ( .A(n23677), .B(n23688), .Z(n23679) );
  XOR U24713 ( .A(n23689), .B(n23690), .Z(n23677) );
  AND U24714 ( .A(n23691), .B(n23692), .Z(n23690) );
  XNOR U24715 ( .A(n23693), .B(n23689), .Z(n23692) );
  XOR U24716 ( .A(n23694), .B(e_input[76]), .Z(n23685) );
  IV U24717 ( .A(n23683), .Z(n23694) );
  XOR U24718 ( .A(n23695), .B(n23696), .Z(n23683) );
  AND U24719 ( .A(n23697), .B(n23698), .Z(n23696) );
  XNOR U24720 ( .A(n23695), .B(n11850), .Z(n23698) );
  XNOR U24721 ( .A(n23691), .B(n23693), .Z(n11850) );
  NAND U24722 ( .A(n23699), .B(e_input[75]), .Z(n23693) );
  NAND U24723 ( .A(n12323), .B(e_input[75]), .Z(n23699) );
  XNOR U24724 ( .A(n23689), .B(n23700), .Z(n23691) );
  XOR U24725 ( .A(n23701), .B(n23702), .Z(n23689) );
  AND U24726 ( .A(n23703), .B(n23704), .Z(n23702) );
  XNOR U24727 ( .A(n23705), .B(n23701), .Z(n23704) );
  XOR U24728 ( .A(n23706), .B(e_input[75]), .Z(n23697) );
  IV U24729 ( .A(n23695), .Z(n23706) );
  XOR U24730 ( .A(n23707), .B(n23708), .Z(n23695) );
  AND U24731 ( .A(n23709), .B(n23710), .Z(n23708) );
  XNOR U24732 ( .A(n23707), .B(n11856), .Z(n23710) );
  XNOR U24733 ( .A(n23703), .B(n23705), .Z(n11856) );
  NAND U24734 ( .A(n23711), .B(e_input[74]), .Z(n23705) );
  NAND U24735 ( .A(n12323), .B(e_input[74]), .Z(n23711) );
  XNOR U24736 ( .A(n23701), .B(n23712), .Z(n23703) );
  XOR U24737 ( .A(n23713), .B(n23714), .Z(n23701) );
  AND U24738 ( .A(n23715), .B(n23716), .Z(n23714) );
  XNOR U24739 ( .A(n23717), .B(n23713), .Z(n23716) );
  XOR U24740 ( .A(n23718), .B(e_input[74]), .Z(n23709) );
  IV U24741 ( .A(n23707), .Z(n23718) );
  XOR U24742 ( .A(n23719), .B(n23720), .Z(n23707) );
  AND U24743 ( .A(n23721), .B(n23722), .Z(n23720) );
  XNOR U24744 ( .A(n23719), .B(n11862), .Z(n23722) );
  XNOR U24745 ( .A(n23715), .B(n23717), .Z(n11862) );
  NAND U24746 ( .A(n23723), .B(e_input[73]), .Z(n23717) );
  NAND U24747 ( .A(n12323), .B(e_input[73]), .Z(n23723) );
  XNOR U24748 ( .A(n23713), .B(n23724), .Z(n23715) );
  XOR U24749 ( .A(n23725), .B(n23726), .Z(n23713) );
  AND U24750 ( .A(n23727), .B(n23728), .Z(n23726) );
  XNOR U24751 ( .A(n23729), .B(n23725), .Z(n23728) );
  XOR U24752 ( .A(n23730), .B(e_input[73]), .Z(n23721) );
  IV U24753 ( .A(n23719), .Z(n23730) );
  XOR U24754 ( .A(n23731), .B(n23732), .Z(n23719) );
  AND U24755 ( .A(n23733), .B(n23734), .Z(n23732) );
  XNOR U24756 ( .A(n23731), .B(n11868), .Z(n23734) );
  XNOR U24757 ( .A(n23727), .B(n23729), .Z(n11868) );
  NAND U24758 ( .A(n23735), .B(e_input[72]), .Z(n23729) );
  NAND U24759 ( .A(n12323), .B(e_input[72]), .Z(n23735) );
  XNOR U24760 ( .A(n23725), .B(n23736), .Z(n23727) );
  XOR U24761 ( .A(n23737), .B(n23738), .Z(n23725) );
  AND U24762 ( .A(n23739), .B(n23740), .Z(n23738) );
  XNOR U24763 ( .A(n23741), .B(n23737), .Z(n23740) );
  XOR U24764 ( .A(n23742), .B(e_input[72]), .Z(n23733) );
  IV U24765 ( .A(n23731), .Z(n23742) );
  XOR U24766 ( .A(n23743), .B(n23744), .Z(n23731) );
  AND U24767 ( .A(n23745), .B(n23746), .Z(n23744) );
  XNOR U24768 ( .A(n23743), .B(n11874), .Z(n23746) );
  XNOR U24769 ( .A(n23739), .B(n23741), .Z(n11874) );
  NAND U24770 ( .A(n23747), .B(e_input[71]), .Z(n23741) );
  NAND U24771 ( .A(n12323), .B(e_input[71]), .Z(n23747) );
  XNOR U24772 ( .A(n23737), .B(n23748), .Z(n23739) );
  XOR U24773 ( .A(n23749), .B(n23750), .Z(n23737) );
  AND U24774 ( .A(n23751), .B(n23752), .Z(n23750) );
  XNOR U24775 ( .A(n23753), .B(n23749), .Z(n23752) );
  XOR U24776 ( .A(n23754), .B(e_input[71]), .Z(n23745) );
  IV U24777 ( .A(n23743), .Z(n23754) );
  XOR U24778 ( .A(n23755), .B(n23756), .Z(n23743) );
  AND U24779 ( .A(n23757), .B(n23758), .Z(n23756) );
  XNOR U24780 ( .A(n23755), .B(n11880), .Z(n23758) );
  XNOR U24781 ( .A(n23751), .B(n23753), .Z(n11880) );
  NAND U24782 ( .A(n23759), .B(e_input[70]), .Z(n23753) );
  NAND U24783 ( .A(n12323), .B(e_input[70]), .Z(n23759) );
  XNOR U24784 ( .A(n23749), .B(n23760), .Z(n23751) );
  XOR U24785 ( .A(n23761), .B(n23762), .Z(n23749) );
  AND U24786 ( .A(n23763), .B(n23764), .Z(n23762) );
  XNOR U24787 ( .A(n23765), .B(n23761), .Z(n23764) );
  XOR U24788 ( .A(n23766), .B(e_input[70]), .Z(n23757) );
  IV U24789 ( .A(n23755), .Z(n23766) );
  XOR U24790 ( .A(n23767), .B(n23768), .Z(n23755) );
  AND U24791 ( .A(n23769), .B(n23770), .Z(n23768) );
  XNOR U24792 ( .A(n23767), .B(n11886), .Z(n23770) );
  XNOR U24793 ( .A(n23763), .B(n23765), .Z(n11886) );
  NAND U24794 ( .A(n23771), .B(e_input[69]), .Z(n23765) );
  NAND U24795 ( .A(n12323), .B(e_input[69]), .Z(n23771) );
  XNOR U24796 ( .A(n23761), .B(n23772), .Z(n23763) );
  XOR U24797 ( .A(n23773), .B(n23774), .Z(n23761) );
  AND U24798 ( .A(n23775), .B(n23776), .Z(n23774) );
  XNOR U24799 ( .A(n23777), .B(n23773), .Z(n23776) );
  XOR U24800 ( .A(n23778), .B(e_input[69]), .Z(n23769) );
  IV U24801 ( .A(n23767), .Z(n23778) );
  XOR U24802 ( .A(n23779), .B(n23780), .Z(n23767) );
  AND U24803 ( .A(n23781), .B(n23782), .Z(n23780) );
  XNOR U24804 ( .A(n23779), .B(n11892), .Z(n23782) );
  XNOR U24805 ( .A(n23775), .B(n23777), .Z(n11892) );
  NAND U24806 ( .A(n23783), .B(e_input[68]), .Z(n23777) );
  NAND U24807 ( .A(n12323), .B(e_input[68]), .Z(n23783) );
  XNOR U24808 ( .A(n23773), .B(n23784), .Z(n23775) );
  XOR U24809 ( .A(n23785), .B(n23786), .Z(n23773) );
  AND U24810 ( .A(n23787), .B(n23788), .Z(n23786) );
  XNOR U24811 ( .A(n23789), .B(n23785), .Z(n23788) );
  XOR U24812 ( .A(n23790), .B(e_input[68]), .Z(n23781) );
  IV U24813 ( .A(n23779), .Z(n23790) );
  XOR U24814 ( .A(n23791), .B(n23792), .Z(n23779) );
  AND U24815 ( .A(n23793), .B(n23794), .Z(n23792) );
  XNOR U24816 ( .A(n23791), .B(n11898), .Z(n23794) );
  XNOR U24817 ( .A(n23787), .B(n23789), .Z(n11898) );
  NAND U24818 ( .A(n23795), .B(e_input[67]), .Z(n23789) );
  NAND U24819 ( .A(n12323), .B(e_input[67]), .Z(n23795) );
  XNOR U24820 ( .A(n23785), .B(n23796), .Z(n23787) );
  XOR U24821 ( .A(n23797), .B(n23798), .Z(n23785) );
  AND U24822 ( .A(n23799), .B(n23800), .Z(n23798) );
  XNOR U24823 ( .A(n23801), .B(n23797), .Z(n23800) );
  XOR U24824 ( .A(n23802), .B(e_input[67]), .Z(n23793) );
  IV U24825 ( .A(n23791), .Z(n23802) );
  XOR U24826 ( .A(n23803), .B(n23804), .Z(n23791) );
  AND U24827 ( .A(n23805), .B(n23806), .Z(n23804) );
  XNOR U24828 ( .A(n23803), .B(n11904), .Z(n23806) );
  XNOR U24829 ( .A(n23799), .B(n23801), .Z(n11904) );
  NAND U24830 ( .A(n23807), .B(e_input[66]), .Z(n23801) );
  NAND U24831 ( .A(n12323), .B(e_input[66]), .Z(n23807) );
  XNOR U24832 ( .A(n23797), .B(n23808), .Z(n23799) );
  XOR U24833 ( .A(n23809), .B(n23810), .Z(n23797) );
  AND U24834 ( .A(n23811), .B(n23812), .Z(n23810) );
  XNOR U24835 ( .A(n23813), .B(n23809), .Z(n23812) );
  XOR U24836 ( .A(n23814), .B(e_input[66]), .Z(n23805) );
  IV U24837 ( .A(n23803), .Z(n23814) );
  XOR U24838 ( .A(n23815), .B(n23816), .Z(n23803) );
  AND U24839 ( .A(n23817), .B(n23818), .Z(n23816) );
  XNOR U24840 ( .A(n23815), .B(n11910), .Z(n23818) );
  XNOR U24841 ( .A(n23811), .B(n23813), .Z(n11910) );
  NAND U24842 ( .A(n23819), .B(e_input[65]), .Z(n23813) );
  NAND U24843 ( .A(n12323), .B(e_input[65]), .Z(n23819) );
  XNOR U24844 ( .A(n23809), .B(n23820), .Z(n23811) );
  XOR U24845 ( .A(n23821), .B(n23822), .Z(n23809) );
  AND U24846 ( .A(n23823), .B(n23824), .Z(n23822) );
  XNOR U24847 ( .A(n23825), .B(n23821), .Z(n23824) );
  XOR U24848 ( .A(n23826), .B(e_input[65]), .Z(n23817) );
  IV U24849 ( .A(n23815), .Z(n23826) );
  XOR U24850 ( .A(n23827), .B(n23828), .Z(n23815) );
  AND U24851 ( .A(n23829), .B(n23830), .Z(n23828) );
  XNOR U24852 ( .A(n23827), .B(n11916), .Z(n23830) );
  XNOR U24853 ( .A(n23823), .B(n23825), .Z(n11916) );
  NAND U24854 ( .A(n23831), .B(e_input[64]), .Z(n23825) );
  NAND U24855 ( .A(n12323), .B(e_input[64]), .Z(n23831) );
  XNOR U24856 ( .A(n23821), .B(n23832), .Z(n23823) );
  XOR U24857 ( .A(n23833), .B(n23834), .Z(n23821) );
  AND U24858 ( .A(n23835), .B(n23836), .Z(n23834) );
  XNOR U24859 ( .A(n23837), .B(n23833), .Z(n23836) );
  XOR U24860 ( .A(n23838), .B(e_input[64]), .Z(n23829) );
  IV U24861 ( .A(n23827), .Z(n23838) );
  XOR U24862 ( .A(n23839), .B(n23840), .Z(n23827) );
  AND U24863 ( .A(n23841), .B(n23842), .Z(n23840) );
  XNOR U24864 ( .A(n23839), .B(n11922), .Z(n23842) );
  XNOR U24865 ( .A(n23835), .B(n23837), .Z(n11922) );
  NAND U24866 ( .A(n23843), .B(e_input[63]), .Z(n23837) );
  NAND U24867 ( .A(n12323), .B(e_input[63]), .Z(n23843) );
  XNOR U24868 ( .A(n23833), .B(n23844), .Z(n23835) );
  XOR U24869 ( .A(n23845), .B(n23846), .Z(n23833) );
  AND U24870 ( .A(n23847), .B(n23848), .Z(n23846) );
  XNOR U24871 ( .A(n23849), .B(n23845), .Z(n23848) );
  XOR U24872 ( .A(n23850), .B(e_input[63]), .Z(n23841) );
  IV U24873 ( .A(n23839), .Z(n23850) );
  XOR U24874 ( .A(n23851), .B(n23852), .Z(n23839) );
  AND U24875 ( .A(n23853), .B(n23854), .Z(n23852) );
  XNOR U24876 ( .A(n23851), .B(n11928), .Z(n23854) );
  XNOR U24877 ( .A(n23847), .B(n23849), .Z(n11928) );
  NAND U24878 ( .A(n23855), .B(e_input[62]), .Z(n23849) );
  NAND U24879 ( .A(n12323), .B(e_input[62]), .Z(n23855) );
  XNOR U24880 ( .A(n23845), .B(n23856), .Z(n23847) );
  XOR U24881 ( .A(n23857), .B(n23858), .Z(n23845) );
  AND U24882 ( .A(n23859), .B(n23860), .Z(n23858) );
  XNOR U24883 ( .A(n23861), .B(n23857), .Z(n23860) );
  XOR U24884 ( .A(n23862), .B(e_input[62]), .Z(n23853) );
  IV U24885 ( .A(n23851), .Z(n23862) );
  XOR U24886 ( .A(n23863), .B(n23864), .Z(n23851) );
  AND U24887 ( .A(n23865), .B(n23866), .Z(n23864) );
  XNOR U24888 ( .A(n23863), .B(n11934), .Z(n23866) );
  XNOR U24889 ( .A(n23859), .B(n23861), .Z(n11934) );
  NAND U24890 ( .A(n23867), .B(e_input[61]), .Z(n23861) );
  NAND U24891 ( .A(n12323), .B(e_input[61]), .Z(n23867) );
  XNOR U24892 ( .A(n23857), .B(n23868), .Z(n23859) );
  XOR U24893 ( .A(n23869), .B(n23870), .Z(n23857) );
  AND U24894 ( .A(n23871), .B(n23872), .Z(n23870) );
  XNOR U24895 ( .A(n23873), .B(n23869), .Z(n23872) );
  XOR U24896 ( .A(n23874), .B(e_input[61]), .Z(n23865) );
  IV U24897 ( .A(n23863), .Z(n23874) );
  XOR U24898 ( .A(n23875), .B(n23876), .Z(n23863) );
  AND U24899 ( .A(n23877), .B(n23878), .Z(n23876) );
  XNOR U24900 ( .A(n23875), .B(n11940), .Z(n23878) );
  XNOR U24901 ( .A(n23871), .B(n23873), .Z(n11940) );
  NAND U24902 ( .A(n23879), .B(e_input[60]), .Z(n23873) );
  NAND U24903 ( .A(n12323), .B(e_input[60]), .Z(n23879) );
  XNOR U24904 ( .A(n23869), .B(n23880), .Z(n23871) );
  XOR U24905 ( .A(n23881), .B(n23882), .Z(n23869) );
  AND U24906 ( .A(n23883), .B(n23884), .Z(n23882) );
  XNOR U24907 ( .A(n23885), .B(n23881), .Z(n23884) );
  XOR U24908 ( .A(n23886), .B(e_input[60]), .Z(n23877) );
  IV U24909 ( .A(n23875), .Z(n23886) );
  XOR U24910 ( .A(n23887), .B(n23888), .Z(n23875) );
  AND U24911 ( .A(n23889), .B(n23890), .Z(n23888) );
  XNOR U24912 ( .A(n23887), .B(n11946), .Z(n23890) );
  XNOR U24913 ( .A(n23883), .B(n23885), .Z(n11946) );
  NAND U24914 ( .A(n23891), .B(e_input[59]), .Z(n23885) );
  NAND U24915 ( .A(n12323), .B(e_input[59]), .Z(n23891) );
  XNOR U24916 ( .A(n23881), .B(n23892), .Z(n23883) );
  XOR U24917 ( .A(n23893), .B(n23894), .Z(n23881) );
  AND U24918 ( .A(n23895), .B(n23896), .Z(n23894) );
  XNOR U24919 ( .A(n23897), .B(n23893), .Z(n23896) );
  XOR U24920 ( .A(n23898), .B(e_input[59]), .Z(n23889) );
  IV U24921 ( .A(n23887), .Z(n23898) );
  XOR U24922 ( .A(n23899), .B(n23900), .Z(n23887) );
  AND U24923 ( .A(n23901), .B(n23902), .Z(n23900) );
  XNOR U24924 ( .A(n23899), .B(n11952), .Z(n23902) );
  XNOR U24925 ( .A(n23895), .B(n23897), .Z(n11952) );
  NAND U24926 ( .A(n23903), .B(e_input[58]), .Z(n23897) );
  NAND U24927 ( .A(n12323), .B(e_input[58]), .Z(n23903) );
  XNOR U24928 ( .A(n23893), .B(n23904), .Z(n23895) );
  XOR U24929 ( .A(n23905), .B(n23906), .Z(n23893) );
  AND U24930 ( .A(n23907), .B(n23908), .Z(n23906) );
  XNOR U24931 ( .A(n23909), .B(n23905), .Z(n23908) );
  XOR U24932 ( .A(n23910), .B(e_input[58]), .Z(n23901) );
  IV U24933 ( .A(n23899), .Z(n23910) );
  XOR U24934 ( .A(n23911), .B(n23912), .Z(n23899) );
  AND U24935 ( .A(n23913), .B(n23914), .Z(n23912) );
  XNOR U24936 ( .A(n23911), .B(n11958), .Z(n23914) );
  XNOR U24937 ( .A(n23907), .B(n23909), .Z(n11958) );
  NAND U24938 ( .A(n23915), .B(e_input[57]), .Z(n23909) );
  NAND U24939 ( .A(n12323), .B(e_input[57]), .Z(n23915) );
  XNOR U24940 ( .A(n23905), .B(n23916), .Z(n23907) );
  XOR U24941 ( .A(n23917), .B(n23918), .Z(n23905) );
  AND U24942 ( .A(n23919), .B(n23920), .Z(n23918) );
  XNOR U24943 ( .A(n23921), .B(n23917), .Z(n23920) );
  XOR U24944 ( .A(n23922), .B(e_input[57]), .Z(n23913) );
  IV U24945 ( .A(n23911), .Z(n23922) );
  XOR U24946 ( .A(n23923), .B(n23924), .Z(n23911) );
  AND U24947 ( .A(n23925), .B(n23926), .Z(n23924) );
  XNOR U24948 ( .A(n23923), .B(n11964), .Z(n23926) );
  XNOR U24949 ( .A(n23919), .B(n23921), .Z(n11964) );
  NAND U24950 ( .A(n23927), .B(e_input[56]), .Z(n23921) );
  NAND U24951 ( .A(n12323), .B(e_input[56]), .Z(n23927) );
  XNOR U24952 ( .A(n23917), .B(n23928), .Z(n23919) );
  XOR U24953 ( .A(n23929), .B(n23930), .Z(n23917) );
  AND U24954 ( .A(n23931), .B(n23932), .Z(n23930) );
  XNOR U24955 ( .A(n23933), .B(n23929), .Z(n23932) );
  XOR U24956 ( .A(n23934), .B(e_input[56]), .Z(n23925) );
  IV U24957 ( .A(n23923), .Z(n23934) );
  XOR U24958 ( .A(n23935), .B(n23936), .Z(n23923) );
  AND U24959 ( .A(n23937), .B(n23938), .Z(n23936) );
  XNOR U24960 ( .A(n23935), .B(n11970), .Z(n23938) );
  XNOR U24961 ( .A(n23931), .B(n23933), .Z(n11970) );
  NAND U24962 ( .A(n23939), .B(e_input[55]), .Z(n23933) );
  NAND U24963 ( .A(n12323), .B(e_input[55]), .Z(n23939) );
  XNOR U24964 ( .A(n23929), .B(n23940), .Z(n23931) );
  XOR U24965 ( .A(n23941), .B(n23942), .Z(n23929) );
  AND U24966 ( .A(n23943), .B(n23944), .Z(n23942) );
  XNOR U24967 ( .A(n23945), .B(n23941), .Z(n23944) );
  XOR U24968 ( .A(n23946), .B(e_input[55]), .Z(n23937) );
  IV U24969 ( .A(n23935), .Z(n23946) );
  XOR U24970 ( .A(n23947), .B(n23948), .Z(n23935) );
  AND U24971 ( .A(n23949), .B(n23950), .Z(n23948) );
  XNOR U24972 ( .A(n23947), .B(n11976), .Z(n23950) );
  XNOR U24973 ( .A(n23943), .B(n23945), .Z(n11976) );
  NAND U24974 ( .A(n23951), .B(e_input[54]), .Z(n23945) );
  NAND U24975 ( .A(n12323), .B(e_input[54]), .Z(n23951) );
  XNOR U24976 ( .A(n23941), .B(n23952), .Z(n23943) );
  XOR U24977 ( .A(n23953), .B(n23954), .Z(n23941) );
  AND U24978 ( .A(n23955), .B(n23956), .Z(n23954) );
  XNOR U24979 ( .A(n23957), .B(n23953), .Z(n23956) );
  XOR U24980 ( .A(n23958), .B(e_input[54]), .Z(n23949) );
  IV U24981 ( .A(n23947), .Z(n23958) );
  XOR U24982 ( .A(n23959), .B(n23960), .Z(n23947) );
  AND U24983 ( .A(n23961), .B(n23962), .Z(n23960) );
  XNOR U24984 ( .A(n23959), .B(n11982), .Z(n23962) );
  XNOR U24985 ( .A(n23955), .B(n23957), .Z(n11982) );
  NAND U24986 ( .A(n23963), .B(e_input[53]), .Z(n23957) );
  NAND U24987 ( .A(n12323), .B(e_input[53]), .Z(n23963) );
  XNOR U24988 ( .A(n23953), .B(n23964), .Z(n23955) );
  XOR U24989 ( .A(n23965), .B(n23966), .Z(n23953) );
  AND U24990 ( .A(n23967), .B(n23968), .Z(n23966) );
  XNOR U24991 ( .A(n23969), .B(n23965), .Z(n23968) );
  XOR U24992 ( .A(n23970), .B(e_input[53]), .Z(n23961) );
  IV U24993 ( .A(n23959), .Z(n23970) );
  XOR U24994 ( .A(n23971), .B(n23972), .Z(n23959) );
  AND U24995 ( .A(n23973), .B(n23974), .Z(n23972) );
  XNOR U24996 ( .A(n23971), .B(n11988), .Z(n23974) );
  XNOR U24997 ( .A(n23967), .B(n23969), .Z(n11988) );
  NAND U24998 ( .A(n23975), .B(e_input[52]), .Z(n23969) );
  NAND U24999 ( .A(n12323), .B(e_input[52]), .Z(n23975) );
  XNOR U25000 ( .A(n23965), .B(n23976), .Z(n23967) );
  XOR U25001 ( .A(n23977), .B(n23978), .Z(n23965) );
  AND U25002 ( .A(n23979), .B(n23980), .Z(n23978) );
  XNOR U25003 ( .A(n23981), .B(n23977), .Z(n23980) );
  XOR U25004 ( .A(n23982), .B(e_input[52]), .Z(n23973) );
  IV U25005 ( .A(n23971), .Z(n23982) );
  XOR U25006 ( .A(n23983), .B(n23984), .Z(n23971) );
  AND U25007 ( .A(n23985), .B(n23986), .Z(n23984) );
  XNOR U25008 ( .A(n23983), .B(n11994), .Z(n23986) );
  XNOR U25009 ( .A(n23979), .B(n23981), .Z(n11994) );
  NAND U25010 ( .A(n23987), .B(e_input[51]), .Z(n23981) );
  NAND U25011 ( .A(n12323), .B(e_input[51]), .Z(n23987) );
  XNOR U25012 ( .A(n23977), .B(n23988), .Z(n23979) );
  XOR U25013 ( .A(n23989), .B(n23990), .Z(n23977) );
  AND U25014 ( .A(n23991), .B(n23992), .Z(n23990) );
  XNOR U25015 ( .A(n23993), .B(n23989), .Z(n23992) );
  XOR U25016 ( .A(n23994), .B(e_input[51]), .Z(n23985) );
  IV U25017 ( .A(n23983), .Z(n23994) );
  XOR U25018 ( .A(n23995), .B(n23996), .Z(n23983) );
  AND U25019 ( .A(n23997), .B(n23998), .Z(n23996) );
  XNOR U25020 ( .A(n23995), .B(n12000), .Z(n23998) );
  XNOR U25021 ( .A(n23991), .B(n23993), .Z(n12000) );
  NAND U25022 ( .A(n23999), .B(e_input[50]), .Z(n23993) );
  NAND U25023 ( .A(n12323), .B(e_input[50]), .Z(n23999) );
  XNOR U25024 ( .A(n23989), .B(n24000), .Z(n23991) );
  XOR U25025 ( .A(n24001), .B(n24002), .Z(n23989) );
  AND U25026 ( .A(n24003), .B(n24004), .Z(n24002) );
  XNOR U25027 ( .A(n24005), .B(n24001), .Z(n24004) );
  XOR U25028 ( .A(n24006), .B(e_input[50]), .Z(n23997) );
  IV U25029 ( .A(n23995), .Z(n24006) );
  XOR U25030 ( .A(n24007), .B(n24008), .Z(n23995) );
  AND U25031 ( .A(n24009), .B(n24010), .Z(n24008) );
  XNOR U25032 ( .A(n24007), .B(n12006), .Z(n24010) );
  XNOR U25033 ( .A(n24003), .B(n24005), .Z(n12006) );
  NAND U25034 ( .A(n24011), .B(e_input[49]), .Z(n24005) );
  NAND U25035 ( .A(n12323), .B(e_input[49]), .Z(n24011) );
  XNOR U25036 ( .A(n24001), .B(n24012), .Z(n24003) );
  XOR U25037 ( .A(n24013), .B(n24014), .Z(n24001) );
  AND U25038 ( .A(n24015), .B(n24016), .Z(n24014) );
  XNOR U25039 ( .A(n24017), .B(n24013), .Z(n24016) );
  XOR U25040 ( .A(n24018), .B(e_input[49]), .Z(n24009) );
  IV U25041 ( .A(n24007), .Z(n24018) );
  XOR U25042 ( .A(n24019), .B(n24020), .Z(n24007) );
  AND U25043 ( .A(n24021), .B(n24022), .Z(n24020) );
  XNOR U25044 ( .A(n24019), .B(n12012), .Z(n24022) );
  XNOR U25045 ( .A(n24015), .B(n24017), .Z(n12012) );
  NAND U25046 ( .A(n24023), .B(e_input[48]), .Z(n24017) );
  NAND U25047 ( .A(n12323), .B(e_input[48]), .Z(n24023) );
  XNOR U25048 ( .A(n24013), .B(n24024), .Z(n24015) );
  XOR U25049 ( .A(n24025), .B(n24026), .Z(n24013) );
  AND U25050 ( .A(n24027), .B(n24028), .Z(n24026) );
  XNOR U25051 ( .A(n24029), .B(n24025), .Z(n24028) );
  XOR U25052 ( .A(n24030), .B(e_input[48]), .Z(n24021) );
  IV U25053 ( .A(n24019), .Z(n24030) );
  XOR U25054 ( .A(n24031), .B(n24032), .Z(n24019) );
  AND U25055 ( .A(n24033), .B(n24034), .Z(n24032) );
  XNOR U25056 ( .A(n24031), .B(n12018), .Z(n24034) );
  XNOR U25057 ( .A(n24027), .B(n24029), .Z(n12018) );
  NAND U25058 ( .A(n24035), .B(e_input[47]), .Z(n24029) );
  NAND U25059 ( .A(n12323), .B(e_input[47]), .Z(n24035) );
  XNOR U25060 ( .A(n24025), .B(n24036), .Z(n24027) );
  XOR U25061 ( .A(n24037), .B(n24038), .Z(n24025) );
  AND U25062 ( .A(n24039), .B(n24040), .Z(n24038) );
  XNOR U25063 ( .A(n24041), .B(n24037), .Z(n24040) );
  XOR U25064 ( .A(n24042), .B(e_input[47]), .Z(n24033) );
  IV U25065 ( .A(n24031), .Z(n24042) );
  XOR U25066 ( .A(n24043), .B(n24044), .Z(n24031) );
  AND U25067 ( .A(n24045), .B(n24046), .Z(n24044) );
  XNOR U25068 ( .A(n24043), .B(n12024), .Z(n24046) );
  XNOR U25069 ( .A(n24039), .B(n24041), .Z(n12024) );
  NAND U25070 ( .A(n24047), .B(e_input[46]), .Z(n24041) );
  NAND U25071 ( .A(n12323), .B(e_input[46]), .Z(n24047) );
  XNOR U25072 ( .A(n24037), .B(n24048), .Z(n24039) );
  XOR U25073 ( .A(n24049), .B(n24050), .Z(n24037) );
  AND U25074 ( .A(n24051), .B(n24052), .Z(n24050) );
  XNOR U25075 ( .A(n24053), .B(n24049), .Z(n24052) );
  XOR U25076 ( .A(n24054), .B(e_input[46]), .Z(n24045) );
  IV U25077 ( .A(n24043), .Z(n24054) );
  XOR U25078 ( .A(n24055), .B(n24056), .Z(n24043) );
  AND U25079 ( .A(n24057), .B(n24058), .Z(n24056) );
  XNOR U25080 ( .A(n24055), .B(n12030), .Z(n24058) );
  XNOR U25081 ( .A(n24051), .B(n24053), .Z(n12030) );
  NAND U25082 ( .A(n24059), .B(e_input[45]), .Z(n24053) );
  NAND U25083 ( .A(n12323), .B(e_input[45]), .Z(n24059) );
  XNOR U25084 ( .A(n24049), .B(n24060), .Z(n24051) );
  XOR U25085 ( .A(n24061), .B(n24062), .Z(n24049) );
  AND U25086 ( .A(n24063), .B(n24064), .Z(n24062) );
  XNOR U25087 ( .A(n24065), .B(n24061), .Z(n24064) );
  XOR U25088 ( .A(n24066), .B(e_input[45]), .Z(n24057) );
  IV U25089 ( .A(n24055), .Z(n24066) );
  XOR U25090 ( .A(n24067), .B(n24068), .Z(n24055) );
  AND U25091 ( .A(n24069), .B(n24070), .Z(n24068) );
  XNOR U25092 ( .A(n24067), .B(n12036), .Z(n24070) );
  XNOR U25093 ( .A(n24063), .B(n24065), .Z(n12036) );
  NAND U25094 ( .A(n24071), .B(e_input[44]), .Z(n24065) );
  NAND U25095 ( .A(n12323), .B(e_input[44]), .Z(n24071) );
  XNOR U25096 ( .A(n24061), .B(n24072), .Z(n24063) );
  XOR U25097 ( .A(n24073), .B(n24074), .Z(n24061) );
  AND U25098 ( .A(n24075), .B(n24076), .Z(n24074) );
  XNOR U25099 ( .A(n24077), .B(n24073), .Z(n24076) );
  XOR U25100 ( .A(n24078), .B(e_input[44]), .Z(n24069) );
  IV U25101 ( .A(n24067), .Z(n24078) );
  XOR U25102 ( .A(n24079), .B(n24080), .Z(n24067) );
  AND U25103 ( .A(n24081), .B(n24082), .Z(n24080) );
  XNOR U25104 ( .A(n24079), .B(n12042), .Z(n24082) );
  XNOR U25105 ( .A(n24075), .B(n24077), .Z(n12042) );
  NAND U25106 ( .A(n24083), .B(e_input[43]), .Z(n24077) );
  NAND U25107 ( .A(n12323), .B(e_input[43]), .Z(n24083) );
  XNOR U25108 ( .A(n24073), .B(n24084), .Z(n24075) );
  XOR U25109 ( .A(n24085), .B(n24086), .Z(n24073) );
  AND U25110 ( .A(n24087), .B(n24088), .Z(n24086) );
  XNOR U25111 ( .A(n24089), .B(n24085), .Z(n24088) );
  XOR U25112 ( .A(n24090), .B(e_input[43]), .Z(n24081) );
  IV U25113 ( .A(n24079), .Z(n24090) );
  XOR U25114 ( .A(n24091), .B(n24092), .Z(n24079) );
  AND U25115 ( .A(n24093), .B(n24094), .Z(n24092) );
  XNOR U25116 ( .A(n24091), .B(n12048), .Z(n24094) );
  XNOR U25117 ( .A(n24087), .B(n24089), .Z(n12048) );
  NAND U25118 ( .A(n24095), .B(e_input[42]), .Z(n24089) );
  NAND U25119 ( .A(n12323), .B(e_input[42]), .Z(n24095) );
  XNOR U25120 ( .A(n24085), .B(n24096), .Z(n24087) );
  XOR U25121 ( .A(n24097), .B(n24098), .Z(n24085) );
  AND U25122 ( .A(n24099), .B(n24100), .Z(n24098) );
  XNOR U25123 ( .A(n24101), .B(n24097), .Z(n24100) );
  XOR U25124 ( .A(n24102), .B(e_input[42]), .Z(n24093) );
  IV U25125 ( .A(n24091), .Z(n24102) );
  XOR U25126 ( .A(n24103), .B(n24104), .Z(n24091) );
  AND U25127 ( .A(n24105), .B(n24106), .Z(n24104) );
  XNOR U25128 ( .A(n24103), .B(n12054), .Z(n24106) );
  XNOR U25129 ( .A(n24099), .B(n24101), .Z(n12054) );
  NAND U25130 ( .A(n24107), .B(e_input[41]), .Z(n24101) );
  NAND U25131 ( .A(n12323), .B(e_input[41]), .Z(n24107) );
  XNOR U25132 ( .A(n24097), .B(n24108), .Z(n24099) );
  XOR U25133 ( .A(n24109), .B(n24110), .Z(n24097) );
  AND U25134 ( .A(n24111), .B(n24112), .Z(n24110) );
  XNOR U25135 ( .A(n24113), .B(n24109), .Z(n24112) );
  XOR U25136 ( .A(n24114), .B(e_input[41]), .Z(n24105) );
  IV U25137 ( .A(n24103), .Z(n24114) );
  XOR U25138 ( .A(n24115), .B(n24116), .Z(n24103) );
  AND U25139 ( .A(n24117), .B(n24118), .Z(n24116) );
  XNOR U25140 ( .A(n24115), .B(n12060), .Z(n24118) );
  XNOR U25141 ( .A(n24111), .B(n24113), .Z(n12060) );
  NAND U25142 ( .A(n24119), .B(e_input[40]), .Z(n24113) );
  NAND U25143 ( .A(n12323), .B(e_input[40]), .Z(n24119) );
  XNOR U25144 ( .A(n24109), .B(n24120), .Z(n24111) );
  XOR U25145 ( .A(n24121), .B(n24122), .Z(n24109) );
  AND U25146 ( .A(n24123), .B(n24124), .Z(n24122) );
  XNOR U25147 ( .A(n24125), .B(n24121), .Z(n24124) );
  XOR U25148 ( .A(n24126), .B(e_input[40]), .Z(n24117) );
  IV U25149 ( .A(n24115), .Z(n24126) );
  XOR U25150 ( .A(n24127), .B(n24128), .Z(n24115) );
  AND U25151 ( .A(n24129), .B(n24130), .Z(n24128) );
  XNOR U25152 ( .A(n24127), .B(n12066), .Z(n24130) );
  XNOR U25153 ( .A(n24123), .B(n24125), .Z(n12066) );
  NAND U25154 ( .A(n24131), .B(e_input[39]), .Z(n24125) );
  NAND U25155 ( .A(n12323), .B(e_input[39]), .Z(n24131) );
  XNOR U25156 ( .A(n24121), .B(n24132), .Z(n24123) );
  XOR U25157 ( .A(n24133), .B(n24134), .Z(n24121) );
  AND U25158 ( .A(n24135), .B(n24136), .Z(n24134) );
  XNOR U25159 ( .A(n24137), .B(n24133), .Z(n24136) );
  XOR U25160 ( .A(n24138), .B(e_input[39]), .Z(n24129) );
  IV U25161 ( .A(n24127), .Z(n24138) );
  XOR U25162 ( .A(n24139), .B(n24140), .Z(n24127) );
  AND U25163 ( .A(n24141), .B(n24142), .Z(n24140) );
  XNOR U25164 ( .A(n24139), .B(n12072), .Z(n24142) );
  XNOR U25165 ( .A(n24135), .B(n24137), .Z(n12072) );
  NAND U25166 ( .A(n24143), .B(e_input[38]), .Z(n24137) );
  NAND U25167 ( .A(n12323), .B(e_input[38]), .Z(n24143) );
  XNOR U25168 ( .A(n24133), .B(n24144), .Z(n24135) );
  XOR U25169 ( .A(n24145), .B(n24146), .Z(n24133) );
  AND U25170 ( .A(n24147), .B(n24148), .Z(n24146) );
  XNOR U25171 ( .A(n24149), .B(n24145), .Z(n24148) );
  XOR U25172 ( .A(n24150), .B(e_input[38]), .Z(n24141) );
  IV U25173 ( .A(n24139), .Z(n24150) );
  XOR U25174 ( .A(n24151), .B(n24152), .Z(n24139) );
  AND U25175 ( .A(n24153), .B(n24154), .Z(n24152) );
  XNOR U25176 ( .A(n24151), .B(n12078), .Z(n24154) );
  XNOR U25177 ( .A(n24147), .B(n24149), .Z(n12078) );
  NAND U25178 ( .A(n24155), .B(e_input[37]), .Z(n24149) );
  NAND U25179 ( .A(n12323), .B(e_input[37]), .Z(n24155) );
  XNOR U25180 ( .A(n24145), .B(n24156), .Z(n24147) );
  XOR U25181 ( .A(n24157), .B(n24158), .Z(n24145) );
  AND U25182 ( .A(n24159), .B(n24160), .Z(n24158) );
  XNOR U25183 ( .A(n24161), .B(n24157), .Z(n24160) );
  XOR U25184 ( .A(n24162), .B(e_input[37]), .Z(n24153) );
  IV U25185 ( .A(n24151), .Z(n24162) );
  XOR U25186 ( .A(n24163), .B(n24164), .Z(n24151) );
  AND U25187 ( .A(n24165), .B(n24166), .Z(n24164) );
  XNOR U25188 ( .A(n24163), .B(n12084), .Z(n24166) );
  XNOR U25189 ( .A(n24159), .B(n24161), .Z(n12084) );
  NAND U25190 ( .A(n24167), .B(e_input[36]), .Z(n24161) );
  NAND U25191 ( .A(n12323), .B(e_input[36]), .Z(n24167) );
  XNOR U25192 ( .A(n24157), .B(n24168), .Z(n24159) );
  XOR U25193 ( .A(n24169), .B(n24170), .Z(n24157) );
  AND U25194 ( .A(n24171), .B(n24172), .Z(n24170) );
  XNOR U25195 ( .A(n24173), .B(n24169), .Z(n24172) );
  XOR U25196 ( .A(n24174), .B(e_input[36]), .Z(n24165) );
  IV U25197 ( .A(n24163), .Z(n24174) );
  XOR U25198 ( .A(n24175), .B(n24176), .Z(n24163) );
  AND U25199 ( .A(n24177), .B(n24178), .Z(n24176) );
  XNOR U25200 ( .A(n24175), .B(n12090), .Z(n24178) );
  XNOR U25201 ( .A(n24171), .B(n24173), .Z(n12090) );
  NAND U25202 ( .A(n24179), .B(e_input[35]), .Z(n24173) );
  NAND U25203 ( .A(n12323), .B(e_input[35]), .Z(n24179) );
  XNOR U25204 ( .A(n24169), .B(n24180), .Z(n24171) );
  XOR U25205 ( .A(n24181), .B(n24182), .Z(n24169) );
  AND U25206 ( .A(n24183), .B(n24184), .Z(n24182) );
  XNOR U25207 ( .A(n24185), .B(n24181), .Z(n24184) );
  XOR U25208 ( .A(n24186), .B(e_input[35]), .Z(n24177) );
  IV U25209 ( .A(n24175), .Z(n24186) );
  XOR U25210 ( .A(n24187), .B(n24188), .Z(n24175) );
  AND U25211 ( .A(n24189), .B(n24190), .Z(n24188) );
  XNOR U25212 ( .A(n24187), .B(n12096), .Z(n24190) );
  XNOR U25213 ( .A(n24183), .B(n24185), .Z(n12096) );
  NAND U25214 ( .A(n24191), .B(e_input[34]), .Z(n24185) );
  NAND U25215 ( .A(n12323), .B(e_input[34]), .Z(n24191) );
  XNOR U25216 ( .A(n24181), .B(n24192), .Z(n24183) );
  XOR U25217 ( .A(n24193), .B(n24194), .Z(n24181) );
  AND U25218 ( .A(n24195), .B(n24196), .Z(n24194) );
  XNOR U25219 ( .A(n24197), .B(n24193), .Z(n24196) );
  XOR U25220 ( .A(n24198), .B(e_input[34]), .Z(n24189) );
  IV U25221 ( .A(n24187), .Z(n24198) );
  XOR U25222 ( .A(n24199), .B(n24200), .Z(n24187) );
  AND U25223 ( .A(n24201), .B(n24202), .Z(n24200) );
  XNOR U25224 ( .A(n24199), .B(n12102), .Z(n24202) );
  XNOR U25225 ( .A(n24195), .B(n24197), .Z(n12102) );
  NAND U25226 ( .A(n24203), .B(e_input[33]), .Z(n24197) );
  NAND U25227 ( .A(n12323), .B(e_input[33]), .Z(n24203) );
  XNOR U25228 ( .A(n24193), .B(n24204), .Z(n24195) );
  XOR U25229 ( .A(n24205), .B(n24206), .Z(n24193) );
  AND U25230 ( .A(n24207), .B(n24208), .Z(n24206) );
  XNOR U25231 ( .A(n24209), .B(n24205), .Z(n24208) );
  XOR U25232 ( .A(n24210), .B(e_input[33]), .Z(n24201) );
  IV U25233 ( .A(n24199), .Z(n24210) );
  XOR U25234 ( .A(n24211), .B(n24212), .Z(n24199) );
  AND U25235 ( .A(n24213), .B(n24214), .Z(n24212) );
  XNOR U25236 ( .A(n24211), .B(n12108), .Z(n24214) );
  XNOR U25237 ( .A(n24207), .B(n24209), .Z(n12108) );
  NAND U25238 ( .A(n24215), .B(e_input[32]), .Z(n24209) );
  NAND U25239 ( .A(n12323), .B(e_input[32]), .Z(n24215) );
  XNOR U25240 ( .A(n24205), .B(n24216), .Z(n24207) );
  XOR U25241 ( .A(n24217), .B(n24218), .Z(n24205) );
  AND U25242 ( .A(n24219), .B(n24220), .Z(n24218) );
  XNOR U25243 ( .A(n24221), .B(n24217), .Z(n24220) );
  XOR U25244 ( .A(n24222), .B(e_input[32]), .Z(n24213) );
  IV U25245 ( .A(n24211), .Z(n24222) );
  XOR U25246 ( .A(n24223), .B(n24224), .Z(n24211) );
  AND U25247 ( .A(n24225), .B(n24226), .Z(n24224) );
  XNOR U25248 ( .A(n24223), .B(n12114), .Z(n24226) );
  XNOR U25249 ( .A(n24219), .B(n24221), .Z(n12114) );
  NAND U25250 ( .A(n24227), .B(e_input[31]), .Z(n24221) );
  NAND U25251 ( .A(n12323), .B(e_input[31]), .Z(n24227) );
  XNOR U25252 ( .A(n24217), .B(n24228), .Z(n24219) );
  XOR U25253 ( .A(n24229), .B(n24230), .Z(n24217) );
  AND U25254 ( .A(n24231), .B(n24232), .Z(n24230) );
  XNOR U25255 ( .A(n24233), .B(n24229), .Z(n24232) );
  XOR U25256 ( .A(n24234), .B(e_input[31]), .Z(n24225) );
  IV U25257 ( .A(n24223), .Z(n24234) );
  XOR U25258 ( .A(n24235), .B(n24236), .Z(n24223) );
  AND U25259 ( .A(n24237), .B(n24238), .Z(n24236) );
  XNOR U25260 ( .A(n24235), .B(n12120), .Z(n24238) );
  XNOR U25261 ( .A(n24231), .B(n24233), .Z(n12120) );
  NAND U25262 ( .A(n24239), .B(e_input[30]), .Z(n24233) );
  NAND U25263 ( .A(n12323), .B(e_input[30]), .Z(n24239) );
  XNOR U25264 ( .A(n24229), .B(n24240), .Z(n24231) );
  XOR U25265 ( .A(n24241), .B(n24242), .Z(n24229) );
  AND U25266 ( .A(n24243), .B(n24244), .Z(n24242) );
  XNOR U25267 ( .A(n24245), .B(n24241), .Z(n24244) );
  XOR U25268 ( .A(n24246), .B(e_input[30]), .Z(n24237) );
  IV U25269 ( .A(n24235), .Z(n24246) );
  XOR U25270 ( .A(n24247), .B(n24248), .Z(n24235) );
  AND U25271 ( .A(n24249), .B(n24250), .Z(n24248) );
  XNOR U25272 ( .A(n24247), .B(n12126), .Z(n24250) );
  XNOR U25273 ( .A(n24243), .B(n24245), .Z(n12126) );
  NAND U25274 ( .A(n24251), .B(e_input[29]), .Z(n24245) );
  NAND U25275 ( .A(n12323), .B(e_input[29]), .Z(n24251) );
  XNOR U25276 ( .A(n24241), .B(n24252), .Z(n24243) );
  XOR U25277 ( .A(n24253), .B(n24254), .Z(n24241) );
  AND U25278 ( .A(n24255), .B(n24256), .Z(n24254) );
  XNOR U25279 ( .A(n24257), .B(n24253), .Z(n24256) );
  XOR U25280 ( .A(n24258), .B(e_input[29]), .Z(n24249) );
  IV U25281 ( .A(n24247), .Z(n24258) );
  XOR U25282 ( .A(n24259), .B(n24260), .Z(n24247) );
  AND U25283 ( .A(n24261), .B(n24262), .Z(n24260) );
  XNOR U25284 ( .A(n24259), .B(n12132), .Z(n24262) );
  XNOR U25285 ( .A(n24255), .B(n24257), .Z(n12132) );
  NAND U25286 ( .A(n24263), .B(e_input[28]), .Z(n24257) );
  NAND U25287 ( .A(n12323), .B(e_input[28]), .Z(n24263) );
  XNOR U25288 ( .A(n24253), .B(n24264), .Z(n24255) );
  XOR U25289 ( .A(n24265), .B(n24266), .Z(n24253) );
  AND U25290 ( .A(n24267), .B(n24268), .Z(n24266) );
  XNOR U25291 ( .A(n24269), .B(n24265), .Z(n24268) );
  XOR U25292 ( .A(n24270), .B(e_input[28]), .Z(n24261) );
  IV U25293 ( .A(n24259), .Z(n24270) );
  XOR U25294 ( .A(n24271), .B(n24272), .Z(n24259) );
  AND U25295 ( .A(n24273), .B(n24274), .Z(n24272) );
  XNOR U25296 ( .A(n24271), .B(n12138), .Z(n24274) );
  XNOR U25297 ( .A(n24267), .B(n24269), .Z(n12138) );
  NAND U25298 ( .A(n24275), .B(e_input[27]), .Z(n24269) );
  NAND U25299 ( .A(n12323), .B(e_input[27]), .Z(n24275) );
  XNOR U25300 ( .A(n24265), .B(n24276), .Z(n24267) );
  XOR U25301 ( .A(n24277), .B(n24278), .Z(n24265) );
  AND U25302 ( .A(n24279), .B(n24280), .Z(n24278) );
  XNOR U25303 ( .A(n24281), .B(n24277), .Z(n24280) );
  XOR U25304 ( .A(n24282), .B(e_input[27]), .Z(n24273) );
  IV U25305 ( .A(n24271), .Z(n24282) );
  XOR U25306 ( .A(n24283), .B(n24284), .Z(n24271) );
  AND U25307 ( .A(n24285), .B(n24286), .Z(n24284) );
  XNOR U25308 ( .A(n24283), .B(n12144), .Z(n24286) );
  XNOR U25309 ( .A(n24279), .B(n24281), .Z(n12144) );
  NAND U25310 ( .A(n24287), .B(e_input[26]), .Z(n24281) );
  NAND U25311 ( .A(n12323), .B(e_input[26]), .Z(n24287) );
  XNOR U25312 ( .A(n24277), .B(n24288), .Z(n24279) );
  XOR U25313 ( .A(n24289), .B(n24290), .Z(n24277) );
  AND U25314 ( .A(n24291), .B(n24292), .Z(n24290) );
  XNOR U25315 ( .A(n24293), .B(n24289), .Z(n24292) );
  XOR U25316 ( .A(n24294), .B(e_input[26]), .Z(n24285) );
  IV U25317 ( .A(n24283), .Z(n24294) );
  XOR U25318 ( .A(n24295), .B(n24296), .Z(n24283) );
  AND U25319 ( .A(n24297), .B(n24298), .Z(n24296) );
  XNOR U25320 ( .A(n24295), .B(n12150), .Z(n24298) );
  XNOR U25321 ( .A(n24291), .B(n24293), .Z(n12150) );
  NAND U25322 ( .A(n24299), .B(e_input[25]), .Z(n24293) );
  NAND U25323 ( .A(n12323), .B(e_input[25]), .Z(n24299) );
  XNOR U25324 ( .A(n24289), .B(n24300), .Z(n24291) );
  XOR U25325 ( .A(n24301), .B(n24302), .Z(n24289) );
  AND U25326 ( .A(n24303), .B(n24304), .Z(n24302) );
  XNOR U25327 ( .A(n24305), .B(n24301), .Z(n24304) );
  XOR U25328 ( .A(n24306), .B(e_input[25]), .Z(n24297) );
  IV U25329 ( .A(n24295), .Z(n24306) );
  XOR U25330 ( .A(n24307), .B(n24308), .Z(n24295) );
  AND U25331 ( .A(n24309), .B(n24310), .Z(n24308) );
  XNOR U25332 ( .A(n24307), .B(n12156), .Z(n24310) );
  XNOR U25333 ( .A(n24303), .B(n24305), .Z(n12156) );
  NAND U25334 ( .A(n24311), .B(e_input[24]), .Z(n24305) );
  NAND U25335 ( .A(n12323), .B(e_input[24]), .Z(n24311) );
  XNOR U25336 ( .A(n24301), .B(n24312), .Z(n24303) );
  XOR U25337 ( .A(n24313), .B(n24314), .Z(n24301) );
  AND U25338 ( .A(n24315), .B(n24316), .Z(n24314) );
  XNOR U25339 ( .A(n24317), .B(n24313), .Z(n24316) );
  XOR U25340 ( .A(n24318), .B(e_input[24]), .Z(n24309) );
  IV U25341 ( .A(n24307), .Z(n24318) );
  XOR U25342 ( .A(n24319), .B(n24320), .Z(n24307) );
  AND U25343 ( .A(n24321), .B(n24322), .Z(n24320) );
  XNOR U25344 ( .A(n24319), .B(n12162), .Z(n24322) );
  XNOR U25345 ( .A(n24315), .B(n24317), .Z(n12162) );
  NAND U25346 ( .A(n24323), .B(e_input[23]), .Z(n24317) );
  NAND U25347 ( .A(n12323), .B(e_input[23]), .Z(n24323) );
  XNOR U25348 ( .A(n24313), .B(n24324), .Z(n24315) );
  XOR U25349 ( .A(n24325), .B(n24326), .Z(n24313) );
  AND U25350 ( .A(n24327), .B(n24328), .Z(n24326) );
  XNOR U25351 ( .A(n24329), .B(n24325), .Z(n24328) );
  XOR U25352 ( .A(n24330), .B(e_input[23]), .Z(n24321) );
  IV U25353 ( .A(n24319), .Z(n24330) );
  XOR U25354 ( .A(n24331), .B(n24332), .Z(n24319) );
  AND U25355 ( .A(n24333), .B(n24334), .Z(n24332) );
  XNOR U25356 ( .A(n24331), .B(n12168), .Z(n24334) );
  XNOR U25357 ( .A(n24327), .B(n24329), .Z(n12168) );
  NAND U25358 ( .A(n24335), .B(e_input[22]), .Z(n24329) );
  NAND U25359 ( .A(n12323), .B(e_input[22]), .Z(n24335) );
  XNOR U25360 ( .A(n24325), .B(n24336), .Z(n24327) );
  XOR U25361 ( .A(n24337), .B(n24338), .Z(n24325) );
  AND U25362 ( .A(n24339), .B(n24340), .Z(n24338) );
  XNOR U25363 ( .A(n24341), .B(n24337), .Z(n24340) );
  XOR U25364 ( .A(n24342), .B(e_input[22]), .Z(n24333) );
  IV U25365 ( .A(n24331), .Z(n24342) );
  XOR U25366 ( .A(n24343), .B(n24344), .Z(n24331) );
  AND U25367 ( .A(n24345), .B(n24346), .Z(n24344) );
  XNOR U25368 ( .A(n24343), .B(n12174), .Z(n24346) );
  XNOR U25369 ( .A(n24339), .B(n24341), .Z(n12174) );
  NAND U25370 ( .A(n24347), .B(e_input[21]), .Z(n24341) );
  NAND U25371 ( .A(n12323), .B(e_input[21]), .Z(n24347) );
  XNOR U25372 ( .A(n24337), .B(n24348), .Z(n24339) );
  XOR U25373 ( .A(n24349), .B(n24350), .Z(n24337) );
  AND U25374 ( .A(n24351), .B(n24352), .Z(n24350) );
  XNOR U25375 ( .A(n24353), .B(n24349), .Z(n24352) );
  XOR U25376 ( .A(n24354), .B(e_input[21]), .Z(n24345) );
  IV U25377 ( .A(n24343), .Z(n24354) );
  XOR U25378 ( .A(n24355), .B(n24356), .Z(n24343) );
  AND U25379 ( .A(n24357), .B(n24358), .Z(n24356) );
  XNOR U25380 ( .A(n24355), .B(n12180), .Z(n24358) );
  XNOR U25381 ( .A(n24351), .B(n24353), .Z(n12180) );
  NAND U25382 ( .A(n24359), .B(e_input[20]), .Z(n24353) );
  NAND U25383 ( .A(n12323), .B(e_input[20]), .Z(n24359) );
  XNOR U25384 ( .A(n24349), .B(n24360), .Z(n24351) );
  XOR U25385 ( .A(n24361), .B(n24362), .Z(n24349) );
  AND U25386 ( .A(n24363), .B(n24364), .Z(n24362) );
  XNOR U25387 ( .A(n24365), .B(n24361), .Z(n24364) );
  XOR U25388 ( .A(n24366), .B(e_input[20]), .Z(n24357) );
  IV U25389 ( .A(n24355), .Z(n24366) );
  XOR U25390 ( .A(n24367), .B(n24368), .Z(n24355) );
  AND U25391 ( .A(n24369), .B(n24370), .Z(n24368) );
  XNOR U25392 ( .A(n24367), .B(n12186), .Z(n24370) );
  XNOR U25393 ( .A(n24363), .B(n24365), .Z(n12186) );
  NAND U25394 ( .A(n24371), .B(e_input[19]), .Z(n24365) );
  NAND U25395 ( .A(n12323), .B(e_input[19]), .Z(n24371) );
  XNOR U25396 ( .A(n24361), .B(n24372), .Z(n24363) );
  XOR U25397 ( .A(n24373), .B(n24374), .Z(n24361) );
  AND U25398 ( .A(n24375), .B(n24376), .Z(n24374) );
  XNOR U25399 ( .A(n24377), .B(n24373), .Z(n24376) );
  XOR U25400 ( .A(n24378), .B(e_input[19]), .Z(n24369) );
  IV U25401 ( .A(n24367), .Z(n24378) );
  XOR U25402 ( .A(n24379), .B(n24380), .Z(n24367) );
  AND U25403 ( .A(n24381), .B(n24382), .Z(n24380) );
  XNOR U25404 ( .A(n24379), .B(n12192), .Z(n24382) );
  XNOR U25405 ( .A(n24375), .B(n24377), .Z(n12192) );
  NAND U25406 ( .A(n24383), .B(e_input[18]), .Z(n24377) );
  NAND U25407 ( .A(n12323), .B(e_input[18]), .Z(n24383) );
  XNOR U25408 ( .A(n24373), .B(n24384), .Z(n24375) );
  XOR U25409 ( .A(n24385), .B(n24386), .Z(n24373) );
  AND U25410 ( .A(n24387), .B(n24388), .Z(n24386) );
  XNOR U25411 ( .A(n24389), .B(n24385), .Z(n24388) );
  XOR U25412 ( .A(n24390), .B(e_input[18]), .Z(n24381) );
  IV U25413 ( .A(n24379), .Z(n24390) );
  XOR U25414 ( .A(n24391), .B(n24392), .Z(n24379) );
  AND U25415 ( .A(n24393), .B(n24394), .Z(n24392) );
  XNOR U25416 ( .A(n24391), .B(n12198), .Z(n24394) );
  XNOR U25417 ( .A(n24387), .B(n24389), .Z(n12198) );
  NAND U25418 ( .A(n24395), .B(e_input[17]), .Z(n24389) );
  NAND U25419 ( .A(n12323), .B(e_input[17]), .Z(n24395) );
  XNOR U25420 ( .A(n24385), .B(n24396), .Z(n24387) );
  XOR U25421 ( .A(n24397), .B(n24398), .Z(n24385) );
  AND U25422 ( .A(n24399), .B(n24400), .Z(n24398) );
  XNOR U25423 ( .A(n24401), .B(n24397), .Z(n24400) );
  XOR U25424 ( .A(n24402), .B(e_input[17]), .Z(n24393) );
  IV U25425 ( .A(n24391), .Z(n24402) );
  XOR U25426 ( .A(n24403), .B(n24404), .Z(n24391) );
  AND U25427 ( .A(n24405), .B(n24406), .Z(n24404) );
  XNOR U25428 ( .A(n24403), .B(n12204), .Z(n24406) );
  XNOR U25429 ( .A(n24399), .B(n24401), .Z(n12204) );
  NAND U25430 ( .A(n24407), .B(e_input[16]), .Z(n24401) );
  NAND U25431 ( .A(n12323), .B(e_input[16]), .Z(n24407) );
  XNOR U25432 ( .A(n24397), .B(n24408), .Z(n24399) );
  XOR U25433 ( .A(n24409), .B(n24410), .Z(n24397) );
  AND U25434 ( .A(n24411), .B(n24412), .Z(n24410) );
  XNOR U25435 ( .A(n24413), .B(n24409), .Z(n24412) );
  XOR U25436 ( .A(n24414), .B(e_input[16]), .Z(n24405) );
  IV U25437 ( .A(n24403), .Z(n24414) );
  XOR U25438 ( .A(n24415), .B(n24416), .Z(n24403) );
  AND U25439 ( .A(n24417), .B(n24418), .Z(n24416) );
  XNOR U25440 ( .A(n24415), .B(n12210), .Z(n24418) );
  XNOR U25441 ( .A(n24411), .B(n24413), .Z(n12210) );
  NAND U25442 ( .A(n24419), .B(e_input[15]), .Z(n24413) );
  NAND U25443 ( .A(n12323), .B(e_input[15]), .Z(n24419) );
  XNOR U25444 ( .A(n24409), .B(n24420), .Z(n24411) );
  XOR U25445 ( .A(n24421), .B(n24422), .Z(n24409) );
  AND U25446 ( .A(n24423), .B(n24424), .Z(n24422) );
  XNOR U25447 ( .A(n24425), .B(n24421), .Z(n24424) );
  XOR U25448 ( .A(n24426), .B(e_input[15]), .Z(n24417) );
  IV U25449 ( .A(n24415), .Z(n24426) );
  XOR U25450 ( .A(n24427), .B(n24428), .Z(n24415) );
  AND U25451 ( .A(n24429), .B(n24430), .Z(n24428) );
  XNOR U25452 ( .A(n24427), .B(n12216), .Z(n24430) );
  XNOR U25453 ( .A(n24423), .B(n24425), .Z(n12216) );
  NAND U25454 ( .A(n24431), .B(e_input[14]), .Z(n24425) );
  NAND U25455 ( .A(n12323), .B(e_input[14]), .Z(n24431) );
  XNOR U25456 ( .A(n24421), .B(n24432), .Z(n24423) );
  XOR U25457 ( .A(n24433), .B(n24434), .Z(n24421) );
  AND U25458 ( .A(n24435), .B(n24436), .Z(n24434) );
  XNOR U25459 ( .A(n24437), .B(n24433), .Z(n24436) );
  XOR U25460 ( .A(n24438), .B(e_input[14]), .Z(n24429) );
  IV U25461 ( .A(n24427), .Z(n24438) );
  XOR U25462 ( .A(n24439), .B(n24440), .Z(n24427) );
  AND U25463 ( .A(n24441), .B(n24442), .Z(n24440) );
  XNOR U25464 ( .A(n24439), .B(n12222), .Z(n24442) );
  XNOR U25465 ( .A(n24435), .B(n24437), .Z(n12222) );
  NAND U25466 ( .A(n24443), .B(e_input[13]), .Z(n24437) );
  NAND U25467 ( .A(n12323), .B(e_input[13]), .Z(n24443) );
  XNOR U25468 ( .A(n24433), .B(n24444), .Z(n24435) );
  XOR U25469 ( .A(n24445), .B(n24446), .Z(n24433) );
  AND U25470 ( .A(n24447), .B(n24448), .Z(n24446) );
  XNOR U25471 ( .A(n24449), .B(n24445), .Z(n24448) );
  XOR U25472 ( .A(n24450), .B(e_input[13]), .Z(n24441) );
  IV U25473 ( .A(n24439), .Z(n24450) );
  XOR U25474 ( .A(n24451), .B(n24452), .Z(n24439) );
  AND U25475 ( .A(n24453), .B(n24454), .Z(n24452) );
  XNOR U25476 ( .A(n24451), .B(n12228), .Z(n24454) );
  XNOR U25477 ( .A(n24447), .B(n24449), .Z(n12228) );
  NAND U25478 ( .A(n24455), .B(e_input[12]), .Z(n24449) );
  NAND U25479 ( .A(n12323), .B(e_input[12]), .Z(n24455) );
  XNOR U25480 ( .A(n24445), .B(n24456), .Z(n24447) );
  XOR U25481 ( .A(n24457), .B(n24458), .Z(n24445) );
  AND U25482 ( .A(n24459), .B(n24460), .Z(n24458) );
  XNOR U25483 ( .A(n24461), .B(n24457), .Z(n24460) );
  XOR U25484 ( .A(n24462), .B(e_input[12]), .Z(n24453) );
  IV U25485 ( .A(n24451), .Z(n24462) );
  XOR U25486 ( .A(n24463), .B(n24464), .Z(n24451) );
  AND U25487 ( .A(n24465), .B(n24466), .Z(n24464) );
  XNOR U25488 ( .A(n24463), .B(n12234), .Z(n24466) );
  XNOR U25489 ( .A(n24459), .B(n24461), .Z(n12234) );
  NAND U25490 ( .A(n24467), .B(e_input[11]), .Z(n24461) );
  NAND U25491 ( .A(n12323), .B(e_input[11]), .Z(n24467) );
  XNOR U25492 ( .A(n24457), .B(n24468), .Z(n24459) );
  XOR U25493 ( .A(n24469), .B(n24470), .Z(n24457) );
  AND U25494 ( .A(n24471), .B(n24472), .Z(n24470) );
  XNOR U25495 ( .A(n24473), .B(n24469), .Z(n24472) );
  XOR U25496 ( .A(n24474), .B(e_input[11]), .Z(n24465) );
  IV U25497 ( .A(n24463), .Z(n24474) );
  XOR U25498 ( .A(n24475), .B(n24476), .Z(n24463) );
  AND U25499 ( .A(n24477), .B(n24478), .Z(n24476) );
  XNOR U25500 ( .A(n24475), .B(n12240), .Z(n24478) );
  XNOR U25501 ( .A(n24471), .B(n24473), .Z(n12240) );
  NAND U25502 ( .A(n24479), .B(e_input[10]), .Z(n24473) );
  NAND U25503 ( .A(n12323), .B(e_input[10]), .Z(n24479) );
  XNOR U25504 ( .A(n24469), .B(n24480), .Z(n24471) );
  XOR U25505 ( .A(n24481), .B(n24482), .Z(n24469) );
  AND U25506 ( .A(n24483), .B(n24484), .Z(n24482) );
  XNOR U25507 ( .A(n24485), .B(n24481), .Z(n24484) );
  XOR U25508 ( .A(n24486), .B(e_input[10]), .Z(n24477) );
  IV U25509 ( .A(n24475), .Z(n24486) );
  XOR U25510 ( .A(n24487), .B(n24488), .Z(n24475) );
  AND U25511 ( .A(n24489), .B(n24490), .Z(n24488) );
  XNOR U25512 ( .A(n12246), .B(n24487), .Z(n24490) );
  XNOR U25513 ( .A(n24483), .B(n24485), .Z(n12246) );
  NAND U25514 ( .A(n24491), .B(e_input[9]), .Z(n24485) );
  NAND U25515 ( .A(n12323), .B(e_input[9]), .Z(n24491) );
  XNOR U25516 ( .A(n24481), .B(n24492), .Z(n24483) );
  XOR U25517 ( .A(n24493), .B(n24494), .Z(n24481) );
  AND U25518 ( .A(n24495), .B(n24496), .Z(n24494) );
  XNOR U25519 ( .A(n24497), .B(n24493), .Z(n24496) );
  XOR U25520 ( .A(n24498), .B(e_input[9]), .Z(n24489) );
  IV U25521 ( .A(n24487), .Z(n24498) );
  XOR U25522 ( .A(n24499), .B(n24500), .Z(n24487) );
  AND U25523 ( .A(n24501), .B(n24502), .Z(n24500) );
  XNOR U25524 ( .A(n24499), .B(n12252), .Z(n24502) );
  XNOR U25525 ( .A(n24495), .B(n24497), .Z(n12252) );
  NAND U25526 ( .A(n24503), .B(e_input[8]), .Z(n24497) );
  NAND U25527 ( .A(n12323), .B(e_input[8]), .Z(n24503) );
  XNOR U25528 ( .A(n24493), .B(n24504), .Z(n24495) );
  XOR U25529 ( .A(n24505), .B(n24506), .Z(n24493) );
  AND U25530 ( .A(n24507), .B(n24508), .Z(n24506) );
  XNOR U25531 ( .A(n24509), .B(n24505), .Z(n24508) );
  XOR U25532 ( .A(n24510), .B(e_input[8]), .Z(n24501) );
  IV U25533 ( .A(n24499), .Z(n24510) );
  XOR U25534 ( .A(n24511), .B(n24512), .Z(n24499) );
  AND U25535 ( .A(n24513), .B(n24514), .Z(n24512) );
  XNOR U25536 ( .A(n24511), .B(n12258), .Z(n24514) );
  XNOR U25537 ( .A(n24507), .B(n24509), .Z(n12258) );
  NAND U25538 ( .A(n24515), .B(e_input[7]), .Z(n24509) );
  NAND U25539 ( .A(n12323), .B(e_input[7]), .Z(n24515) );
  XNOR U25540 ( .A(n24505), .B(n24516), .Z(n24507) );
  XOR U25541 ( .A(n24517), .B(n24518), .Z(n24505) );
  AND U25542 ( .A(n24519), .B(n24520), .Z(n24518) );
  XNOR U25543 ( .A(n24521), .B(n24517), .Z(n24520) );
  XOR U25544 ( .A(n24522), .B(e_input[7]), .Z(n24513) );
  IV U25545 ( .A(n24511), .Z(n24522) );
  XOR U25546 ( .A(n24523), .B(n24524), .Z(n24511) );
  AND U25547 ( .A(n24525), .B(n24526), .Z(n24524) );
  XNOR U25548 ( .A(n24523), .B(n12264), .Z(n24526) );
  XNOR U25549 ( .A(n24519), .B(n24521), .Z(n12264) );
  NAND U25550 ( .A(n24527), .B(e_input[6]), .Z(n24521) );
  NAND U25551 ( .A(n12323), .B(e_input[6]), .Z(n24527) );
  XNOR U25552 ( .A(n24517), .B(n24528), .Z(n24519) );
  XOR U25553 ( .A(n24529), .B(n24530), .Z(n24517) );
  AND U25554 ( .A(n24531), .B(n24532), .Z(n24530) );
  XNOR U25555 ( .A(n24533), .B(n24529), .Z(n24532) );
  XOR U25556 ( .A(n24534), .B(e_input[6]), .Z(n24525) );
  IV U25557 ( .A(n24523), .Z(n24534) );
  XOR U25558 ( .A(n24535), .B(n24536), .Z(n24523) );
  AND U25559 ( .A(n24537), .B(n24538), .Z(n24536) );
  XNOR U25560 ( .A(n24535), .B(n12270), .Z(n24538) );
  XNOR U25561 ( .A(n24531), .B(n24533), .Z(n12270) );
  NAND U25562 ( .A(n24539), .B(e_input[5]), .Z(n24533) );
  NAND U25563 ( .A(n12323), .B(e_input[5]), .Z(n24539) );
  XNOR U25564 ( .A(n24529), .B(n24540), .Z(n24531) );
  XOR U25565 ( .A(n24541), .B(n24542), .Z(n24529) );
  AND U25566 ( .A(n24543), .B(n24544), .Z(n24542) );
  XNOR U25567 ( .A(n24545), .B(n24541), .Z(n24544) );
  XOR U25568 ( .A(n24546), .B(e_input[5]), .Z(n24537) );
  IV U25569 ( .A(n24535), .Z(n24546) );
  XOR U25570 ( .A(n24547), .B(n24548), .Z(n24535) );
  AND U25571 ( .A(n24549), .B(n24550), .Z(n24548) );
  XNOR U25572 ( .A(n24547), .B(n12276), .Z(n24550) );
  XNOR U25573 ( .A(n24543), .B(n24545), .Z(n12276) );
  NAND U25574 ( .A(n24551), .B(e_input[4]), .Z(n24545) );
  NAND U25575 ( .A(n12323), .B(e_input[4]), .Z(n24551) );
  XNOR U25576 ( .A(n24541), .B(n24552), .Z(n24543) );
  XOR U25577 ( .A(n24553), .B(n24554), .Z(n24541) );
  AND U25578 ( .A(n24555), .B(n24556), .Z(n24554) );
  XNOR U25579 ( .A(n24557), .B(n24553), .Z(n24556) );
  XOR U25580 ( .A(n24558), .B(e_input[4]), .Z(n24549) );
  IV U25581 ( .A(n24547), .Z(n24558) );
  XOR U25582 ( .A(n24559), .B(n24560), .Z(n24547) );
  AND U25583 ( .A(n24561), .B(n24562), .Z(n24560) );
  XNOR U25584 ( .A(n24559), .B(n12282), .Z(n24562) );
  XNOR U25585 ( .A(n24555), .B(n24557), .Z(n12282) );
  NAND U25586 ( .A(n24563), .B(e_input[3]), .Z(n24557) );
  NAND U25587 ( .A(n12323), .B(e_input[3]), .Z(n24563) );
  XNOR U25588 ( .A(n24553), .B(n24564), .Z(n24555) );
  XOR U25589 ( .A(n24565), .B(n24566), .Z(n24553) );
  AND U25590 ( .A(n24567), .B(n24568), .Z(n24566) );
  XNOR U25591 ( .A(n24569), .B(n24565), .Z(n24568) );
  XOR U25592 ( .A(n24570), .B(e_input[3]), .Z(n24561) );
  IV U25593 ( .A(n24559), .Z(n24570) );
  XNOR U25594 ( .A(n24571), .B(n24572), .Z(n24559) );
  AND U25595 ( .A(n24573), .B(n24574), .Z(n24572) );
  XOR U25596 ( .A(n24571), .B(n12287), .Z(n24574) );
  XNOR U25597 ( .A(n24567), .B(n24569), .Z(n12287) );
  NAND U25598 ( .A(n24575), .B(e_input[2]), .Z(n24569) );
  NAND U25599 ( .A(n12323), .B(e_input[2]), .Z(n24575) );
  XOR U25600 ( .A(n24565), .B(n24576), .Z(n24567) );
  XOR U25601 ( .A(n24577), .B(n24578), .Z(n24565) );
  NANDN U25602 ( .B(n24579), .A(n24580), .Z(n24577) );
  XOR U25603 ( .A(n24578), .B(n24581), .Z(n24580) );
  XOR U25604 ( .A(n24571), .B(e_input[2]), .Z(n24573) );
  XOR U25605 ( .A(n24582), .B(n24583), .Z(n24571) );
  NAND U25606 ( .A(n24584), .B(n24585), .Z(n24582) );
  XOR U25607 ( .A(n24583), .B(n12294), .Z(n24585) );
  XNOR U25608 ( .A(n24579), .B(n24581), .Z(n12294) );
  NAND U25609 ( .A(n24586), .B(e_input[1]), .Z(n24581) );
  NAND U25610 ( .A(n12323), .B(e_input[1]), .Z(n24586) );
  XNOR U25611 ( .A(n24587), .B(n24578), .Z(n24579) );
  OR U25612 ( .A(n24588), .B(n24589), .Z(n24578) );
  XNOR U25613 ( .A(n24583), .B(e_input[1]), .Z(n24584) );
  NOR U25614 ( .A(e_input[0]), .B(n12295), .Z(n24583) );
  XOR U25615 ( .A(n24588), .B(n24589), .Z(n12295) );
  NAND U25616 ( .A(n24590), .B(e_input[0]), .Z(n24589) );
  NAND U25617 ( .A(n12323), .B(e_input[0]), .Z(n24590) );
  NAND U25618 ( .A(n24591), .B(n24592), .Z(n12323) );
  NAND U25619 ( .A(n24593), .B(n24592), .Z(n24591) );
  XOR U25620 ( .A(n12306), .B(n24592), .Z(n24593) );
  AND U25621 ( .A(n24594), .B(n24595), .Z(n24592) );
  NAND U25622 ( .A(n24596), .B(n24595), .Z(n24594) );
  XNOR U25623 ( .A(n12312), .B(n24595), .Z(n24596) );
  XOR U25624 ( .A(n24597), .B(n24598), .Z(n24595) );
  AND U25625 ( .A(n24599), .B(n24600), .Z(n24598) );
  XOR U25626 ( .A(e_input[1023]), .B(n24597), .Z(n24600) );
  XNOR U25627 ( .A(n12324), .B(n24597), .Z(n24599) );
  XOR U25628 ( .A(n24601), .B(n24602), .Z(n12324) );
  XOR U25629 ( .A(n24603), .B(n24604), .Z(n24597) );
  AND U25630 ( .A(n24605), .B(n24606), .Z(n24604) );
  XOR U25631 ( .A(e_input[1022]), .B(n24603), .Z(n24606) );
  XNOR U25632 ( .A(n12336), .B(n24603), .Z(n24605) );
  XOR U25633 ( .A(n24607), .B(n24608), .Z(n12336) );
  XOR U25634 ( .A(n24609), .B(n24610), .Z(n24603) );
  AND U25635 ( .A(n24611), .B(n24612), .Z(n24610) );
  XOR U25636 ( .A(e_input[1021]), .B(n24609), .Z(n24612) );
  XNOR U25637 ( .A(n12348), .B(n24609), .Z(n24611) );
  XOR U25638 ( .A(n24613), .B(n24614), .Z(n12348) );
  XOR U25639 ( .A(n24615), .B(n24616), .Z(n24609) );
  AND U25640 ( .A(n24617), .B(n24618), .Z(n24616) );
  XOR U25641 ( .A(e_input[1020]), .B(n24615), .Z(n24618) );
  XNOR U25642 ( .A(n12360), .B(n24615), .Z(n24617) );
  XOR U25643 ( .A(n24619), .B(n24620), .Z(n12360) );
  XOR U25644 ( .A(n24621), .B(n24622), .Z(n24615) );
  AND U25645 ( .A(n24623), .B(n24624), .Z(n24622) );
  XOR U25646 ( .A(e_input[1019]), .B(n24621), .Z(n24624) );
  XNOR U25647 ( .A(n12372), .B(n24621), .Z(n24623) );
  XOR U25648 ( .A(n24625), .B(n24626), .Z(n12372) );
  XOR U25649 ( .A(n24627), .B(n24628), .Z(n24621) );
  AND U25650 ( .A(n24629), .B(n24630), .Z(n24628) );
  XOR U25651 ( .A(e_input[1018]), .B(n24627), .Z(n24630) );
  XNOR U25652 ( .A(n12384), .B(n24627), .Z(n24629) );
  XOR U25653 ( .A(n24631), .B(n24632), .Z(n12384) );
  XOR U25654 ( .A(n24633), .B(n24634), .Z(n24627) );
  AND U25655 ( .A(n24635), .B(n24636), .Z(n24634) );
  XOR U25656 ( .A(e_input[1017]), .B(n24633), .Z(n24636) );
  XNOR U25657 ( .A(n12396), .B(n24633), .Z(n24635) );
  XOR U25658 ( .A(n24637), .B(n24638), .Z(n12396) );
  XOR U25659 ( .A(n24639), .B(n24640), .Z(n24633) );
  AND U25660 ( .A(n24641), .B(n24642), .Z(n24640) );
  XOR U25661 ( .A(e_input[1016]), .B(n24639), .Z(n24642) );
  XNOR U25662 ( .A(n12408), .B(n24639), .Z(n24641) );
  XOR U25663 ( .A(n24643), .B(n24644), .Z(n12408) );
  XOR U25664 ( .A(n24645), .B(n24646), .Z(n24639) );
  AND U25665 ( .A(n24647), .B(n24648), .Z(n24646) );
  XOR U25666 ( .A(e_input[1015]), .B(n24645), .Z(n24648) );
  XNOR U25667 ( .A(n12420), .B(n24645), .Z(n24647) );
  XOR U25668 ( .A(n24649), .B(n24650), .Z(n12420) );
  XOR U25669 ( .A(n24651), .B(n24652), .Z(n24645) );
  AND U25670 ( .A(n24653), .B(n24654), .Z(n24652) );
  XOR U25671 ( .A(e_input[1014]), .B(n24651), .Z(n24654) );
  XNOR U25672 ( .A(n12432), .B(n24651), .Z(n24653) );
  XOR U25673 ( .A(n24655), .B(n24656), .Z(n12432) );
  XOR U25674 ( .A(n24657), .B(n24658), .Z(n24651) );
  AND U25675 ( .A(n24659), .B(n24660), .Z(n24658) );
  XOR U25676 ( .A(e_input[1013]), .B(n24657), .Z(n24660) );
  XNOR U25677 ( .A(n12444), .B(n24657), .Z(n24659) );
  XOR U25678 ( .A(n24661), .B(n24662), .Z(n12444) );
  XOR U25679 ( .A(n24663), .B(n24664), .Z(n24657) );
  AND U25680 ( .A(n24665), .B(n24666), .Z(n24664) );
  XOR U25681 ( .A(e_input[1012]), .B(n24663), .Z(n24666) );
  XNOR U25682 ( .A(n12456), .B(n24663), .Z(n24665) );
  XOR U25683 ( .A(n24667), .B(n24668), .Z(n12456) );
  XOR U25684 ( .A(n24669), .B(n24670), .Z(n24663) );
  AND U25685 ( .A(n24671), .B(n24672), .Z(n24670) );
  XOR U25686 ( .A(e_input[1011]), .B(n24669), .Z(n24672) );
  XNOR U25687 ( .A(n12468), .B(n24669), .Z(n24671) );
  XOR U25688 ( .A(n24673), .B(n24674), .Z(n12468) );
  XOR U25689 ( .A(n24675), .B(n24676), .Z(n24669) );
  AND U25690 ( .A(n24677), .B(n24678), .Z(n24676) );
  XOR U25691 ( .A(e_input[1010]), .B(n24675), .Z(n24678) );
  XNOR U25692 ( .A(n12480), .B(n24675), .Z(n24677) );
  XOR U25693 ( .A(n24679), .B(n24680), .Z(n12480) );
  XOR U25694 ( .A(n24681), .B(n24682), .Z(n24675) );
  AND U25695 ( .A(n24683), .B(n24684), .Z(n24682) );
  XOR U25696 ( .A(e_input[1009]), .B(n24681), .Z(n24684) );
  XNOR U25697 ( .A(n12492), .B(n24681), .Z(n24683) );
  XOR U25698 ( .A(n24685), .B(n24686), .Z(n12492) );
  XOR U25699 ( .A(n24687), .B(n24688), .Z(n24681) );
  AND U25700 ( .A(n24689), .B(n24690), .Z(n24688) );
  XOR U25701 ( .A(e_input[1008]), .B(n24687), .Z(n24690) );
  XNOR U25702 ( .A(n12504), .B(n24687), .Z(n24689) );
  XOR U25703 ( .A(n24691), .B(n24692), .Z(n12504) );
  XOR U25704 ( .A(n24693), .B(n24694), .Z(n24687) );
  AND U25705 ( .A(n24695), .B(n24696), .Z(n24694) );
  XOR U25706 ( .A(e_input[1007]), .B(n24693), .Z(n24696) );
  XNOR U25707 ( .A(n12516), .B(n24693), .Z(n24695) );
  XOR U25708 ( .A(n24697), .B(n24698), .Z(n12516) );
  XOR U25709 ( .A(n24699), .B(n24700), .Z(n24693) );
  AND U25710 ( .A(n24701), .B(n24702), .Z(n24700) );
  XOR U25711 ( .A(e_input[1006]), .B(n24699), .Z(n24702) );
  XNOR U25712 ( .A(n12528), .B(n24699), .Z(n24701) );
  XOR U25713 ( .A(n24703), .B(n24704), .Z(n12528) );
  XOR U25714 ( .A(n24705), .B(n24706), .Z(n24699) );
  AND U25715 ( .A(n24707), .B(n24708), .Z(n24706) );
  XOR U25716 ( .A(e_input[1005]), .B(n24705), .Z(n24708) );
  XNOR U25717 ( .A(n12540), .B(n24705), .Z(n24707) );
  XOR U25718 ( .A(n24709), .B(n24710), .Z(n12540) );
  XOR U25719 ( .A(n24711), .B(n24712), .Z(n24705) );
  AND U25720 ( .A(n24713), .B(n24714), .Z(n24712) );
  XOR U25721 ( .A(e_input[1004]), .B(n24711), .Z(n24714) );
  XNOR U25722 ( .A(n12552), .B(n24711), .Z(n24713) );
  XOR U25723 ( .A(n24715), .B(n24716), .Z(n12552) );
  XOR U25724 ( .A(n24717), .B(n24718), .Z(n24711) );
  AND U25725 ( .A(n24719), .B(n24720), .Z(n24718) );
  XOR U25726 ( .A(e_input[1003]), .B(n24717), .Z(n24720) );
  XNOR U25727 ( .A(n12564), .B(n24717), .Z(n24719) );
  XOR U25728 ( .A(n24721), .B(n24722), .Z(n12564) );
  XOR U25729 ( .A(n24723), .B(n24724), .Z(n24717) );
  AND U25730 ( .A(n24725), .B(n24726), .Z(n24724) );
  XOR U25731 ( .A(e_input[1002]), .B(n24723), .Z(n24726) );
  XNOR U25732 ( .A(n12576), .B(n24723), .Z(n24725) );
  XOR U25733 ( .A(n24727), .B(n24728), .Z(n12576) );
  XOR U25734 ( .A(n24729), .B(n24730), .Z(n24723) );
  AND U25735 ( .A(n24731), .B(n24732), .Z(n24730) );
  XOR U25736 ( .A(e_input[1001]), .B(n24729), .Z(n24732) );
  XNOR U25737 ( .A(n12588), .B(n24729), .Z(n24731) );
  XOR U25738 ( .A(n24733), .B(n24734), .Z(n12588) );
  XOR U25739 ( .A(n24735), .B(n24736), .Z(n24729) );
  AND U25740 ( .A(n24737), .B(n24738), .Z(n24736) );
  XOR U25741 ( .A(e_input[1000]), .B(n24735), .Z(n24738) );
  XNOR U25742 ( .A(n12600), .B(n24735), .Z(n24737) );
  XOR U25743 ( .A(n24739), .B(n24740), .Z(n12600) );
  XOR U25744 ( .A(n24741), .B(n24742), .Z(n24735) );
  AND U25745 ( .A(n24743), .B(n24744), .Z(n24742) );
  XOR U25746 ( .A(e_input[999]), .B(n24741), .Z(n24744) );
  XNOR U25747 ( .A(n12612), .B(n24741), .Z(n24743) );
  XOR U25748 ( .A(n24745), .B(n24746), .Z(n12612) );
  XOR U25749 ( .A(n24747), .B(n24748), .Z(n24741) );
  AND U25750 ( .A(n24749), .B(n24750), .Z(n24748) );
  XOR U25751 ( .A(e_input[998]), .B(n24747), .Z(n24750) );
  XNOR U25752 ( .A(n12624), .B(n24747), .Z(n24749) );
  XOR U25753 ( .A(n24751), .B(n24752), .Z(n12624) );
  XOR U25754 ( .A(n24753), .B(n24754), .Z(n24747) );
  AND U25755 ( .A(n24755), .B(n24756), .Z(n24754) );
  XOR U25756 ( .A(e_input[997]), .B(n24753), .Z(n24756) );
  XNOR U25757 ( .A(n12636), .B(n24753), .Z(n24755) );
  XOR U25758 ( .A(n24757), .B(n24758), .Z(n12636) );
  XOR U25759 ( .A(n24759), .B(n24760), .Z(n24753) );
  AND U25760 ( .A(n24761), .B(n24762), .Z(n24760) );
  XOR U25761 ( .A(e_input[996]), .B(n24759), .Z(n24762) );
  XNOR U25762 ( .A(n12648), .B(n24759), .Z(n24761) );
  XOR U25763 ( .A(n24763), .B(n24764), .Z(n12648) );
  XOR U25764 ( .A(n24765), .B(n24766), .Z(n24759) );
  AND U25765 ( .A(n24767), .B(n24768), .Z(n24766) );
  XOR U25766 ( .A(e_input[995]), .B(n24765), .Z(n24768) );
  XNOR U25767 ( .A(n12660), .B(n24765), .Z(n24767) );
  XOR U25768 ( .A(n24769), .B(n24770), .Z(n12660) );
  XOR U25769 ( .A(n24771), .B(n24772), .Z(n24765) );
  AND U25770 ( .A(n24773), .B(n24774), .Z(n24772) );
  XOR U25771 ( .A(e_input[994]), .B(n24771), .Z(n24774) );
  XNOR U25772 ( .A(n12672), .B(n24771), .Z(n24773) );
  XOR U25773 ( .A(n24775), .B(n24776), .Z(n12672) );
  XOR U25774 ( .A(n24777), .B(n24778), .Z(n24771) );
  AND U25775 ( .A(n24779), .B(n24780), .Z(n24778) );
  XOR U25776 ( .A(e_input[993]), .B(n24777), .Z(n24780) );
  XNOR U25777 ( .A(n12684), .B(n24777), .Z(n24779) );
  XOR U25778 ( .A(n24781), .B(n24782), .Z(n12684) );
  XOR U25779 ( .A(n24783), .B(n24784), .Z(n24777) );
  AND U25780 ( .A(n24785), .B(n24786), .Z(n24784) );
  XOR U25781 ( .A(e_input[992]), .B(n24783), .Z(n24786) );
  XNOR U25782 ( .A(n12696), .B(n24783), .Z(n24785) );
  XOR U25783 ( .A(n24787), .B(n24788), .Z(n12696) );
  XOR U25784 ( .A(n24789), .B(n24790), .Z(n24783) );
  AND U25785 ( .A(n24791), .B(n24792), .Z(n24790) );
  XOR U25786 ( .A(e_input[991]), .B(n24789), .Z(n24792) );
  XNOR U25787 ( .A(n12708), .B(n24789), .Z(n24791) );
  XOR U25788 ( .A(n24793), .B(n24794), .Z(n12708) );
  XOR U25789 ( .A(n24795), .B(n24796), .Z(n24789) );
  AND U25790 ( .A(n24797), .B(n24798), .Z(n24796) );
  XOR U25791 ( .A(e_input[990]), .B(n24795), .Z(n24798) );
  XNOR U25792 ( .A(n12720), .B(n24795), .Z(n24797) );
  XOR U25793 ( .A(n24799), .B(n24800), .Z(n12720) );
  XOR U25794 ( .A(n24801), .B(n24802), .Z(n24795) );
  AND U25795 ( .A(n24803), .B(n24804), .Z(n24802) );
  XOR U25796 ( .A(e_input[989]), .B(n24801), .Z(n24804) );
  XNOR U25797 ( .A(n12732), .B(n24801), .Z(n24803) );
  XOR U25798 ( .A(n24805), .B(n24806), .Z(n12732) );
  XOR U25799 ( .A(n24807), .B(n24808), .Z(n24801) );
  AND U25800 ( .A(n24809), .B(n24810), .Z(n24808) );
  XOR U25801 ( .A(e_input[988]), .B(n24807), .Z(n24810) );
  XNOR U25802 ( .A(n12744), .B(n24807), .Z(n24809) );
  XOR U25803 ( .A(n24811), .B(n24812), .Z(n12744) );
  XOR U25804 ( .A(n24813), .B(n24814), .Z(n24807) );
  AND U25805 ( .A(n24815), .B(n24816), .Z(n24814) );
  XOR U25806 ( .A(e_input[987]), .B(n24813), .Z(n24816) );
  XNOR U25807 ( .A(n12756), .B(n24813), .Z(n24815) );
  XOR U25808 ( .A(n24817), .B(n24818), .Z(n12756) );
  XOR U25809 ( .A(n24819), .B(n24820), .Z(n24813) );
  AND U25810 ( .A(n24821), .B(n24822), .Z(n24820) );
  XOR U25811 ( .A(e_input[986]), .B(n24819), .Z(n24822) );
  XNOR U25812 ( .A(n12768), .B(n24819), .Z(n24821) );
  XOR U25813 ( .A(n24823), .B(n24824), .Z(n12768) );
  XOR U25814 ( .A(n24825), .B(n24826), .Z(n24819) );
  AND U25815 ( .A(n24827), .B(n24828), .Z(n24826) );
  XOR U25816 ( .A(e_input[985]), .B(n24825), .Z(n24828) );
  XNOR U25817 ( .A(n12780), .B(n24825), .Z(n24827) );
  XOR U25818 ( .A(n24829), .B(n24830), .Z(n12780) );
  XOR U25819 ( .A(n24831), .B(n24832), .Z(n24825) );
  AND U25820 ( .A(n24833), .B(n24834), .Z(n24832) );
  XOR U25821 ( .A(e_input[984]), .B(n24831), .Z(n24834) );
  XNOR U25822 ( .A(n12792), .B(n24831), .Z(n24833) );
  XOR U25823 ( .A(n24835), .B(n24836), .Z(n12792) );
  XOR U25824 ( .A(n24837), .B(n24838), .Z(n24831) );
  AND U25825 ( .A(n24839), .B(n24840), .Z(n24838) );
  XOR U25826 ( .A(e_input[983]), .B(n24837), .Z(n24840) );
  XNOR U25827 ( .A(n12804), .B(n24837), .Z(n24839) );
  XOR U25828 ( .A(n24841), .B(n24842), .Z(n12804) );
  XOR U25829 ( .A(n24843), .B(n24844), .Z(n24837) );
  AND U25830 ( .A(n24845), .B(n24846), .Z(n24844) );
  XOR U25831 ( .A(e_input[982]), .B(n24843), .Z(n24846) );
  XNOR U25832 ( .A(n12816), .B(n24843), .Z(n24845) );
  XOR U25833 ( .A(n24847), .B(n24848), .Z(n12816) );
  XOR U25834 ( .A(n24849), .B(n24850), .Z(n24843) );
  AND U25835 ( .A(n24851), .B(n24852), .Z(n24850) );
  XOR U25836 ( .A(e_input[981]), .B(n24849), .Z(n24852) );
  XNOR U25837 ( .A(n12828), .B(n24849), .Z(n24851) );
  XOR U25838 ( .A(n24853), .B(n24854), .Z(n12828) );
  XOR U25839 ( .A(n24855), .B(n24856), .Z(n24849) );
  AND U25840 ( .A(n24857), .B(n24858), .Z(n24856) );
  XOR U25841 ( .A(e_input[980]), .B(n24855), .Z(n24858) );
  XNOR U25842 ( .A(n12840), .B(n24855), .Z(n24857) );
  XOR U25843 ( .A(n24859), .B(n24860), .Z(n12840) );
  XOR U25844 ( .A(n24861), .B(n24862), .Z(n24855) );
  AND U25845 ( .A(n24863), .B(n24864), .Z(n24862) );
  XOR U25846 ( .A(e_input[979]), .B(n24861), .Z(n24864) );
  XNOR U25847 ( .A(n12852), .B(n24861), .Z(n24863) );
  XOR U25848 ( .A(n24865), .B(n24866), .Z(n12852) );
  XOR U25849 ( .A(n24867), .B(n24868), .Z(n24861) );
  AND U25850 ( .A(n24869), .B(n24870), .Z(n24868) );
  XOR U25851 ( .A(e_input[978]), .B(n24867), .Z(n24870) );
  XNOR U25852 ( .A(n12864), .B(n24867), .Z(n24869) );
  XOR U25853 ( .A(n24871), .B(n24872), .Z(n12864) );
  XOR U25854 ( .A(n24873), .B(n24874), .Z(n24867) );
  AND U25855 ( .A(n24875), .B(n24876), .Z(n24874) );
  XOR U25856 ( .A(e_input[977]), .B(n24873), .Z(n24876) );
  XNOR U25857 ( .A(n12876), .B(n24873), .Z(n24875) );
  XOR U25858 ( .A(n24877), .B(n24878), .Z(n12876) );
  XOR U25859 ( .A(n24879), .B(n24880), .Z(n24873) );
  AND U25860 ( .A(n24881), .B(n24882), .Z(n24880) );
  XOR U25861 ( .A(e_input[976]), .B(n24879), .Z(n24882) );
  XNOR U25862 ( .A(n12888), .B(n24879), .Z(n24881) );
  XOR U25863 ( .A(n24883), .B(n24884), .Z(n12888) );
  XOR U25864 ( .A(n24885), .B(n24886), .Z(n24879) );
  AND U25865 ( .A(n24887), .B(n24888), .Z(n24886) );
  XOR U25866 ( .A(e_input[975]), .B(n24885), .Z(n24888) );
  XNOR U25867 ( .A(n12900), .B(n24885), .Z(n24887) );
  XOR U25868 ( .A(n24889), .B(n24890), .Z(n12900) );
  XOR U25869 ( .A(n24891), .B(n24892), .Z(n24885) );
  AND U25870 ( .A(n24893), .B(n24894), .Z(n24892) );
  XOR U25871 ( .A(e_input[974]), .B(n24891), .Z(n24894) );
  XNOR U25872 ( .A(n12912), .B(n24891), .Z(n24893) );
  XOR U25873 ( .A(n24895), .B(n24896), .Z(n12912) );
  XOR U25874 ( .A(n24897), .B(n24898), .Z(n24891) );
  AND U25875 ( .A(n24899), .B(n24900), .Z(n24898) );
  XOR U25876 ( .A(e_input[973]), .B(n24897), .Z(n24900) );
  XNOR U25877 ( .A(n12924), .B(n24897), .Z(n24899) );
  XOR U25878 ( .A(n24901), .B(n24902), .Z(n12924) );
  XOR U25879 ( .A(n24903), .B(n24904), .Z(n24897) );
  AND U25880 ( .A(n24905), .B(n24906), .Z(n24904) );
  XOR U25881 ( .A(e_input[972]), .B(n24903), .Z(n24906) );
  XNOR U25882 ( .A(n12936), .B(n24903), .Z(n24905) );
  XOR U25883 ( .A(n24907), .B(n24908), .Z(n12936) );
  XOR U25884 ( .A(n24909), .B(n24910), .Z(n24903) );
  AND U25885 ( .A(n24911), .B(n24912), .Z(n24910) );
  XOR U25886 ( .A(e_input[971]), .B(n24909), .Z(n24912) );
  XNOR U25887 ( .A(n12948), .B(n24909), .Z(n24911) );
  XOR U25888 ( .A(n24913), .B(n24914), .Z(n12948) );
  XOR U25889 ( .A(n24915), .B(n24916), .Z(n24909) );
  AND U25890 ( .A(n24917), .B(n24918), .Z(n24916) );
  XOR U25891 ( .A(e_input[970]), .B(n24915), .Z(n24918) );
  XNOR U25892 ( .A(n12960), .B(n24915), .Z(n24917) );
  XOR U25893 ( .A(n24919), .B(n24920), .Z(n12960) );
  XOR U25894 ( .A(n24921), .B(n24922), .Z(n24915) );
  AND U25895 ( .A(n24923), .B(n24924), .Z(n24922) );
  XOR U25896 ( .A(e_input[969]), .B(n24921), .Z(n24924) );
  XNOR U25897 ( .A(n12972), .B(n24921), .Z(n24923) );
  XOR U25898 ( .A(n24925), .B(n24926), .Z(n12972) );
  XOR U25899 ( .A(n24927), .B(n24928), .Z(n24921) );
  AND U25900 ( .A(n24929), .B(n24930), .Z(n24928) );
  XOR U25901 ( .A(e_input[968]), .B(n24927), .Z(n24930) );
  XNOR U25902 ( .A(n12984), .B(n24927), .Z(n24929) );
  XOR U25903 ( .A(n24931), .B(n24932), .Z(n12984) );
  XOR U25904 ( .A(n24933), .B(n24934), .Z(n24927) );
  AND U25905 ( .A(n24935), .B(n24936), .Z(n24934) );
  XOR U25906 ( .A(e_input[967]), .B(n24933), .Z(n24936) );
  XNOR U25907 ( .A(n12996), .B(n24933), .Z(n24935) );
  XOR U25908 ( .A(n24937), .B(n24938), .Z(n12996) );
  XOR U25909 ( .A(n24939), .B(n24940), .Z(n24933) );
  AND U25910 ( .A(n24941), .B(n24942), .Z(n24940) );
  XOR U25911 ( .A(e_input[966]), .B(n24939), .Z(n24942) );
  XNOR U25912 ( .A(n13008), .B(n24939), .Z(n24941) );
  XOR U25913 ( .A(n24943), .B(n24944), .Z(n13008) );
  XOR U25914 ( .A(n24945), .B(n24946), .Z(n24939) );
  AND U25915 ( .A(n24947), .B(n24948), .Z(n24946) );
  XOR U25916 ( .A(e_input[965]), .B(n24945), .Z(n24948) );
  XNOR U25917 ( .A(n13020), .B(n24945), .Z(n24947) );
  XOR U25918 ( .A(n24949), .B(n24950), .Z(n13020) );
  XOR U25919 ( .A(n24951), .B(n24952), .Z(n24945) );
  AND U25920 ( .A(n24953), .B(n24954), .Z(n24952) );
  XOR U25921 ( .A(e_input[964]), .B(n24951), .Z(n24954) );
  XNOR U25922 ( .A(n13032), .B(n24951), .Z(n24953) );
  XOR U25923 ( .A(n24955), .B(n24956), .Z(n13032) );
  XOR U25924 ( .A(n24957), .B(n24958), .Z(n24951) );
  AND U25925 ( .A(n24959), .B(n24960), .Z(n24958) );
  XOR U25926 ( .A(e_input[963]), .B(n24957), .Z(n24960) );
  XNOR U25927 ( .A(n13044), .B(n24957), .Z(n24959) );
  XOR U25928 ( .A(n24961), .B(n24962), .Z(n13044) );
  XOR U25929 ( .A(n24963), .B(n24964), .Z(n24957) );
  AND U25930 ( .A(n24965), .B(n24966), .Z(n24964) );
  XOR U25931 ( .A(e_input[962]), .B(n24963), .Z(n24966) );
  XNOR U25932 ( .A(n13056), .B(n24963), .Z(n24965) );
  XOR U25933 ( .A(n24967), .B(n24968), .Z(n13056) );
  XOR U25934 ( .A(n24969), .B(n24970), .Z(n24963) );
  AND U25935 ( .A(n24971), .B(n24972), .Z(n24970) );
  XOR U25936 ( .A(e_input[961]), .B(n24969), .Z(n24972) );
  XNOR U25937 ( .A(n13068), .B(n24969), .Z(n24971) );
  XOR U25938 ( .A(n24973), .B(n24974), .Z(n13068) );
  XOR U25939 ( .A(n24975), .B(n24976), .Z(n24969) );
  AND U25940 ( .A(n24977), .B(n24978), .Z(n24976) );
  XOR U25941 ( .A(e_input[960]), .B(n24975), .Z(n24978) );
  XNOR U25942 ( .A(n13080), .B(n24975), .Z(n24977) );
  XOR U25943 ( .A(n24979), .B(n24980), .Z(n13080) );
  XOR U25944 ( .A(n24981), .B(n24982), .Z(n24975) );
  AND U25945 ( .A(n24983), .B(n24984), .Z(n24982) );
  XOR U25946 ( .A(e_input[959]), .B(n24981), .Z(n24984) );
  XNOR U25947 ( .A(n13092), .B(n24981), .Z(n24983) );
  XOR U25948 ( .A(n24985), .B(n24986), .Z(n13092) );
  XOR U25949 ( .A(n24987), .B(n24988), .Z(n24981) );
  AND U25950 ( .A(n24989), .B(n24990), .Z(n24988) );
  XOR U25951 ( .A(e_input[958]), .B(n24987), .Z(n24990) );
  XNOR U25952 ( .A(n13104), .B(n24987), .Z(n24989) );
  XOR U25953 ( .A(n24991), .B(n24992), .Z(n13104) );
  XOR U25954 ( .A(n24993), .B(n24994), .Z(n24987) );
  AND U25955 ( .A(n24995), .B(n24996), .Z(n24994) );
  XOR U25956 ( .A(e_input[957]), .B(n24993), .Z(n24996) );
  XNOR U25957 ( .A(n13116), .B(n24993), .Z(n24995) );
  XOR U25958 ( .A(n24997), .B(n24998), .Z(n13116) );
  XOR U25959 ( .A(n24999), .B(n25000), .Z(n24993) );
  AND U25960 ( .A(n25001), .B(n25002), .Z(n25000) );
  XOR U25961 ( .A(e_input[956]), .B(n24999), .Z(n25002) );
  XNOR U25962 ( .A(n13128), .B(n24999), .Z(n25001) );
  XOR U25963 ( .A(n25003), .B(n25004), .Z(n13128) );
  XOR U25964 ( .A(n25005), .B(n25006), .Z(n24999) );
  AND U25965 ( .A(n25007), .B(n25008), .Z(n25006) );
  XOR U25966 ( .A(e_input[955]), .B(n25005), .Z(n25008) );
  XNOR U25967 ( .A(n13140), .B(n25005), .Z(n25007) );
  XOR U25968 ( .A(n25009), .B(n25010), .Z(n13140) );
  XOR U25969 ( .A(n25011), .B(n25012), .Z(n25005) );
  AND U25970 ( .A(n25013), .B(n25014), .Z(n25012) );
  XOR U25971 ( .A(e_input[954]), .B(n25011), .Z(n25014) );
  XNOR U25972 ( .A(n13152), .B(n25011), .Z(n25013) );
  XOR U25973 ( .A(n25015), .B(n25016), .Z(n13152) );
  XOR U25974 ( .A(n25017), .B(n25018), .Z(n25011) );
  AND U25975 ( .A(n25019), .B(n25020), .Z(n25018) );
  XOR U25976 ( .A(e_input[953]), .B(n25017), .Z(n25020) );
  XNOR U25977 ( .A(n13164), .B(n25017), .Z(n25019) );
  XOR U25978 ( .A(n25021), .B(n25022), .Z(n13164) );
  XOR U25979 ( .A(n25023), .B(n25024), .Z(n25017) );
  AND U25980 ( .A(n25025), .B(n25026), .Z(n25024) );
  XOR U25981 ( .A(e_input[952]), .B(n25023), .Z(n25026) );
  XNOR U25982 ( .A(n13176), .B(n25023), .Z(n25025) );
  XOR U25983 ( .A(n25027), .B(n25028), .Z(n13176) );
  XOR U25984 ( .A(n25029), .B(n25030), .Z(n25023) );
  AND U25985 ( .A(n25031), .B(n25032), .Z(n25030) );
  XOR U25986 ( .A(e_input[951]), .B(n25029), .Z(n25032) );
  XNOR U25987 ( .A(n13188), .B(n25029), .Z(n25031) );
  XOR U25988 ( .A(n25033), .B(n25034), .Z(n13188) );
  XOR U25989 ( .A(n25035), .B(n25036), .Z(n25029) );
  AND U25990 ( .A(n25037), .B(n25038), .Z(n25036) );
  XOR U25991 ( .A(e_input[950]), .B(n25035), .Z(n25038) );
  XNOR U25992 ( .A(n13200), .B(n25035), .Z(n25037) );
  XOR U25993 ( .A(n25039), .B(n25040), .Z(n13200) );
  XOR U25994 ( .A(n25041), .B(n25042), .Z(n25035) );
  AND U25995 ( .A(n25043), .B(n25044), .Z(n25042) );
  XOR U25996 ( .A(e_input[949]), .B(n25041), .Z(n25044) );
  XNOR U25997 ( .A(n13212), .B(n25041), .Z(n25043) );
  XOR U25998 ( .A(n25045), .B(n25046), .Z(n13212) );
  XOR U25999 ( .A(n25047), .B(n25048), .Z(n25041) );
  AND U26000 ( .A(n25049), .B(n25050), .Z(n25048) );
  XOR U26001 ( .A(e_input[948]), .B(n25047), .Z(n25050) );
  XNOR U26002 ( .A(n13224), .B(n25047), .Z(n25049) );
  XOR U26003 ( .A(n25051), .B(n25052), .Z(n13224) );
  XOR U26004 ( .A(n25053), .B(n25054), .Z(n25047) );
  AND U26005 ( .A(n25055), .B(n25056), .Z(n25054) );
  XOR U26006 ( .A(e_input[947]), .B(n25053), .Z(n25056) );
  XNOR U26007 ( .A(n13236), .B(n25053), .Z(n25055) );
  XOR U26008 ( .A(n25057), .B(n25058), .Z(n13236) );
  XOR U26009 ( .A(n25059), .B(n25060), .Z(n25053) );
  AND U26010 ( .A(n25061), .B(n25062), .Z(n25060) );
  XOR U26011 ( .A(e_input[946]), .B(n25059), .Z(n25062) );
  XNOR U26012 ( .A(n13248), .B(n25059), .Z(n25061) );
  XOR U26013 ( .A(n25063), .B(n25064), .Z(n13248) );
  XOR U26014 ( .A(n25065), .B(n25066), .Z(n25059) );
  AND U26015 ( .A(n25067), .B(n25068), .Z(n25066) );
  XOR U26016 ( .A(e_input[945]), .B(n25065), .Z(n25068) );
  XNOR U26017 ( .A(n13260), .B(n25065), .Z(n25067) );
  XOR U26018 ( .A(n25069), .B(n25070), .Z(n13260) );
  XOR U26019 ( .A(n25071), .B(n25072), .Z(n25065) );
  AND U26020 ( .A(n25073), .B(n25074), .Z(n25072) );
  XOR U26021 ( .A(e_input[944]), .B(n25071), .Z(n25074) );
  XNOR U26022 ( .A(n13272), .B(n25071), .Z(n25073) );
  XOR U26023 ( .A(n25075), .B(n25076), .Z(n13272) );
  XOR U26024 ( .A(n25077), .B(n25078), .Z(n25071) );
  AND U26025 ( .A(n25079), .B(n25080), .Z(n25078) );
  XOR U26026 ( .A(e_input[943]), .B(n25077), .Z(n25080) );
  XNOR U26027 ( .A(n13284), .B(n25077), .Z(n25079) );
  XOR U26028 ( .A(n25081), .B(n25082), .Z(n13284) );
  XOR U26029 ( .A(n25083), .B(n25084), .Z(n25077) );
  AND U26030 ( .A(n25085), .B(n25086), .Z(n25084) );
  XOR U26031 ( .A(e_input[942]), .B(n25083), .Z(n25086) );
  XNOR U26032 ( .A(n13296), .B(n25083), .Z(n25085) );
  XOR U26033 ( .A(n25087), .B(n25088), .Z(n13296) );
  XOR U26034 ( .A(n25089), .B(n25090), .Z(n25083) );
  AND U26035 ( .A(n25091), .B(n25092), .Z(n25090) );
  XOR U26036 ( .A(e_input[941]), .B(n25089), .Z(n25092) );
  XNOR U26037 ( .A(n13308), .B(n25089), .Z(n25091) );
  XOR U26038 ( .A(n25093), .B(n25094), .Z(n13308) );
  XOR U26039 ( .A(n25095), .B(n25096), .Z(n25089) );
  AND U26040 ( .A(n25097), .B(n25098), .Z(n25096) );
  XOR U26041 ( .A(e_input[940]), .B(n25095), .Z(n25098) );
  XNOR U26042 ( .A(n13320), .B(n25095), .Z(n25097) );
  XOR U26043 ( .A(n25099), .B(n25100), .Z(n13320) );
  XOR U26044 ( .A(n25101), .B(n25102), .Z(n25095) );
  AND U26045 ( .A(n25103), .B(n25104), .Z(n25102) );
  XOR U26046 ( .A(e_input[939]), .B(n25101), .Z(n25104) );
  XNOR U26047 ( .A(n13332), .B(n25101), .Z(n25103) );
  XOR U26048 ( .A(n25105), .B(n25106), .Z(n13332) );
  XOR U26049 ( .A(n25107), .B(n25108), .Z(n25101) );
  AND U26050 ( .A(n25109), .B(n25110), .Z(n25108) );
  XOR U26051 ( .A(e_input[938]), .B(n25107), .Z(n25110) );
  XNOR U26052 ( .A(n13344), .B(n25107), .Z(n25109) );
  XOR U26053 ( .A(n25111), .B(n25112), .Z(n13344) );
  XOR U26054 ( .A(n25113), .B(n25114), .Z(n25107) );
  AND U26055 ( .A(n25115), .B(n25116), .Z(n25114) );
  XOR U26056 ( .A(e_input[937]), .B(n25113), .Z(n25116) );
  XNOR U26057 ( .A(n13356), .B(n25113), .Z(n25115) );
  XOR U26058 ( .A(n25117), .B(n25118), .Z(n13356) );
  XOR U26059 ( .A(n25119), .B(n25120), .Z(n25113) );
  AND U26060 ( .A(n25121), .B(n25122), .Z(n25120) );
  XOR U26061 ( .A(e_input[936]), .B(n25119), .Z(n25122) );
  XNOR U26062 ( .A(n13368), .B(n25119), .Z(n25121) );
  XOR U26063 ( .A(n25123), .B(n25124), .Z(n13368) );
  XOR U26064 ( .A(n25125), .B(n25126), .Z(n25119) );
  AND U26065 ( .A(n25127), .B(n25128), .Z(n25126) );
  XOR U26066 ( .A(e_input[935]), .B(n25125), .Z(n25128) );
  XNOR U26067 ( .A(n13380), .B(n25125), .Z(n25127) );
  XOR U26068 ( .A(n25129), .B(n25130), .Z(n13380) );
  XOR U26069 ( .A(n25131), .B(n25132), .Z(n25125) );
  AND U26070 ( .A(n25133), .B(n25134), .Z(n25132) );
  XOR U26071 ( .A(e_input[934]), .B(n25131), .Z(n25134) );
  XNOR U26072 ( .A(n13392), .B(n25131), .Z(n25133) );
  XOR U26073 ( .A(n25135), .B(n25136), .Z(n13392) );
  XOR U26074 ( .A(n25137), .B(n25138), .Z(n25131) );
  AND U26075 ( .A(n25139), .B(n25140), .Z(n25138) );
  XOR U26076 ( .A(e_input[933]), .B(n25137), .Z(n25140) );
  XNOR U26077 ( .A(n13404), .B(n25137), .Z(n25139) );
  XOR U26078 ( .A(n25141), .B(n25142), .Z(n13404) );
  XOR U26079 ( .A(n25143), .B(n25144), .Z(n25137) );
  AND U26080 ( .A(n25145), .B(n25146), .Z(n25144) );
  XOR U26081 ( .A(e_input[932]), .B(n25143), .Z(n25146) );
  XNOR U26082 ( .A(n13416), .B(n25143), .Z(n25145) );
  XOR U26083 ( .A(n25147), .B(n25148), .Z(n13416) );
  XOR U26084 ( .A(n25149), .B(n25150), .Z(n25143) );
  AND U26085 ( .A(n25151), .B(n25152), .Z(n25150) );
  XOR U26086 ( .A(e_input[931]), .B(n25149), .Z(n25152) );
  XNOR U26087 ( .A(n13428), .B(n25149), .Z(n25151) );
  XOR U26088 ( .A(n25153), .B(n25154), .Z(n13428) );
  XOR U26089 ( .A(n25155), .B(n25156), .Z(n25149) );
  AND U26090 ( .A(n25157), .B(n25158), .Z(n25156) );
  XOR U26091 ( .A(e_input[930]), .B(n25155), .Z(n25158) );
  XNOR U26092 ( .A(n13440), .B(n25155), .Z(n25157) );
  XOR U26093 ( .A(n25159), .B(n25160), .Z(n13440) );
  XOR U26094 ( .A(n25161), .B(n25162), .Z(n25155) );
  AND U26095 ( .A(n25163), .B(n25164), .Z(n25162) );
  XOR U26096 ( .A(e_input[929]), .B(n25161), .Z(n25164) );
  XNOR U26097 ( .A(n13452), .B(n25161), .Z(n25163) );
  XOR U26098 ( .A(n25165), .B(n25166), .Z(n13452) );
  XOR U26099 ( .A(n25167), .B(n25168), .Z(n25161) );
  AND U26100 ( .A(n25169), .B(n25170), .Z(n25168) );
  XOR U26101 ( .A(e_input[928]), .B(n25167), .Z(n25170) );
  XNOR U26102 ( .A(n13464), .B(n25167), .Z(n25169) );
  XOR U26103 ( .A(n25171), .B(n25172), .Z(n13464) );
  XOR U26104 ( .A(n25173), .B(n25174), .Z(n25167) );
  AND U26105 ( .A(n25175), .B(n25176), .Z(n25174) );
  XOR U26106 ( .A(e_input[927]), .B(n25173), .Z(n25176) );
  XNOR U26107 ( .A(n13476), .B(n25173), .Z(n25175) );
  XOR U26108 ( .A(n25177), .B(n25178), .Z(n13476) );
  XOR U26109 ( .A(n25179), .B(n25180), .Z(n25173) );
  AND U26110 ( .A(n25181), .B(n25182), .Z(n25180) );
  XOR U26111 ( .A(e_input[926]), .B(n25179), .Z(n25182) );
  XNOR U26112 ( .A(n13488), .B(n25179), .Z(n25181) );
  XOR U26113 ( .A(n25183), .B(n25184), .Z(n13488) );
  XOR U26114 ( .A(n25185), .B(n25186), .Z(n25179) );
  AND U26115 ( .A(n25187), .B(n25188), .Z(n25186) );
  XOR U26116 ( .A(e_input[925]), .B(n25185), .Z(n25188) );
  XNOR U26117 ( .A(n13500), .B(n25185), .Z(n25187) );
  XOR U26118 ( .A(n25189), .B(n25190), .Z(n13500) );
  XOR U26119 ( .A(n25191), .B(n25192), .Z(n25185) );
  AND U26120 ( .A(n25193), .B(n25194), .Z(n25192) );
  XOR U26121 ( .A(e_input[924]), .B(n25191), .Z(n25194) );
  XNOR U26122 ( .A(n13512), .B(n25191), .Z(n25193) );
  XOR U26123 ( .A(n25195), .B(n25196), .Z(n13512) );
  XOR U26124 ( .A(n25197), .B(n25198), .Z(n25191) );
  AND U26125 ( .A(n25199), .B(n25200), .Z(n25198) );
  XOR U26126 ( .A(e_input[923]), .B(n25197), .Z(n25200) );
  XNOR U26127 ( .A(n13524), .B(n25197), .Z(n25199) );
  XOR U26128 ( .A(n25201), .B(n25202), .Z(n13524) );
  XOR U26129 ( .A(n25203), .B(n25204), .Z(n25197) );
  AND U26130 ( .A(n25205), .B(n25206), .Z(n25204) );
  XOR U26131 ( .A(e_input[922]), .B(n25203), .Z(n25206) );
  XNOR U26132 ( .A(n13536), .B(n25203), .Z(n25205) );
  XOR U26133 ( .A(n25207), .B(n25208), .Z(n13536) );
  XOR U26134 ( .A(n25209), .B(n25210), .Z(n25203) );
  AND U26135 ( .A(n25211), .B(n25212), .Z(n25210) );
  XOR U26136 ( .A(e_input[921]), .B(n25209), .Z(n25212) );
  XNOR U26137 ( .A(n13548), .B(n25209), .Z(n25211) );
  XOR U26138 ( .A(n25213), .B(n25214), .Z(n13548) );
  XOR U26139 ( .A(n25215), .B(n25216), .Z(n25209) );
  AND U26140 ( .A(n25217), .B(n25218), .Z(n25216) );
  XOR U26141 ( .A(e_input[920]), .B(n25215), .Z(n25218) );
  XNOR U26142 ( .A(n13560), .B(n25215), .Z(n25217) );
  XOR U26143 ( .A(n25219), .B(n25220), .Z(n13560) );
  XOR U26144 ( .A(n25221), .B(n25222), .Z(n25215) );
  AND U26145 ( .A(n25223), .B(n25224), .Z(n25222) );
  XOR U26146 ( .A(e_input[919]), .B(n25221), .Z(n25224) );
  XNOR U26147 ( .A(n13572), .B(n25221), .Z(n25223) );
  XOR U26148 ( .A(n25225), .B(n25226), .Z(n13572) );
  XOR U26149 ( .A(n25227), .B(n25228), .Z(n25221) );
  AND U26150 ( .A(n25229), .B(n25230), .Z(n25228) );
  XOR U26151 ( .A(e_input[918]), .B(n25227), .Z(n25230) );
  XNOR U26152 ( .A(n13584), .B(n25227), .Z(n25229) );
  XOR U26153 ( .A(n25231), .B(n25232), .Z(n13584) );
  XOR U26154 ( .A(n25233), .B(n25234), .Z(n25227) );
  AND U26155 ( .A(n25235), .B(n25236), .Z(n25234) );
  XOR U26156 ( .A(e_input[917]), .B(n25233), .Z(n25236) );
  XNOR U26157 ( .A(n13596), .B(n25233), .Z(n25235) );
  XOR U26158 ( .A(n25237), .B(n25238), .Z(n13596) );
  XOR U26159 ( .A(n25239), .B(n25240), .Z(n25233) );
  AND U26160 ( .A(n25241), .B(n25242), .Z(n25240) );
  XOR U26161 ( .A(e_input[916]), .B(n25239), .Z(n25242) );
  XNOR U26162 ( .A(n13608), .B(n25239), .Z(n25241) );
  XOR U26163 ( .A(n25243), .B(n25244), .Z(n13608) );
  XOR U26164 ( .A(n25245), .B(n25246), .Z(n25239) );
  AND U26165 ( .A(n25247), .B(n25248), .Z(n25246) );
  XOR U26166 ( .A(e_input[915]), .B(n25245), .Z(n25248) );
  XNOR U26167 ( .A(n13620), .B(n25245), .Z(n25247) );
  XOR U26168 ( .A(n25249), .B(n25250), .Z(n13620) );
  XOR U26169 ( .A(n25251), .B(n25252), .Z(n25245) );
  AND U26170 ( .A(n25253), .B(n25254), .Z(n25252) );
  XOR U26171 ( .A(e_input[914]), .B(n25251), .Z(n25254) );
  XNOR U26172 ( .A(n13632), .B(n25251), .Z(n25253) );
  XOR U26173 ( .A(n25255), .B(n25256), .Z(n13632) );
  XOR U26174 ( .A(n25257), .B(n25258), .Z(n25251) );
  AND U26175 ( .A(n25259), .B(n25260), .Z(n25258) );
  XOR U26176 ( .A(e_input[913]), .B(n25257), .Z(n25260) );
  XNOR U26177 ( .A(n13644), .B(n25257), .Z(n25259) );
  XOR U26178 ( .A(n25261), .B(n25262), .Z(n13644) );
  XOR U26179 ( .A(n25263), .B(n25264), .Z(n25257) );
  AND U26180 ( .A(n25265), .B(n25266), .Z(n25264) );
  XOR U26181 ( .A(e_input[912]), .B(n25263), .Z(n25266) );
  XNOR U26182 ( .A(n13656), .B(n25263), .Z(n25265) );
  XOR U26183 ( .A(n25267), .B(n25268), .Z(n13656) );
  XOR U26184 ( .A(n25269), .B(n25270), .Z(n25263) );
  AND U26185 ( .A(n25271), .B(n25272), .Z(n25270) );
  XOR U26186 ( .A(e_input[911]), .B(n25269), .Z(n25272) );
  XNOR U26187 ( .A(n13668), .B(n25269), .Z(n25271) );
  XOR U26188 ( .A(n25273), .B(n25274), .Z(n13668) );
  XOR U26189 ( .A(n25275), .B(n25276), .Z(n25269) );
  AND U26190 ( .A(n25277), .B(n25278), .Z(n25276) );
  XOR U26191 ( .A(e_input[910]), .B(n25275), .Z(n25278) );
  XNOR U26192 ( .A(n13680), .B(n25275), .Z(n25277) );
  XOR U26193 ( .A(n25279), .B(n25280), .Z(n13680) );
  XOR U26194 ( .A(n25281), .B(n25282), .Z(n25275) );
  AND U26195 ( .A(n25283), .B(n25284), .Z(n25282) );
  XOR U26196 ( .A(e_input[909]), .B(n25281), .Z(n25284) );
  XNOR U26197 ( .A(n13692), .B(n25281), .Z(n25283) );
  XOR U26198 ( .A(n25285), .B(n25286), .Z(n13692) );
  XOR U26199 ( .A(n25287), .B(n25288), .Z(n25281) );
  AND U26200 ( .A(n25289), .B(n25290), .Z(n25288) );
  XOR U26201 ( .A(e_input[908]), .B(n25287), .Z(n25290) );
  XNOR U26202 ( .A(n13704), .B(n25287), .Z(n25289) );
  XOR U26203 ( .A(n25291), .B(n25292), .Z(n13704) );
  XOR U26204 ( .A(n25293), .B(n25294), .Z(n25287) );
  AND U26205 ( .A(n25295), .B(n25296), .Z(n25294) );
  XOR U26206 ( .A(e_input[907]), .B(n25293), .Z(n25296) );
  XNOR U26207 ( .A(n13716), .B(n25293), .Z(n25295) );
  XOR U26208 ( .A(n25297), .B(n25298), .Z(n13716) );
  XOR U26209 ( .A(n25299), .B(n25300), .Z(n25293) );
  AND U26210 ( .A(n25301), .B(n25302), .Z(n25300) );
  XOR U26211 ( .A(e_input[906]), .B(n25299), .Z(n25302) );
  XNOR U26212 ( .A(n13728), .B(n25299), .Z(n25301) );
  XOR U26213 ( .A(n25303), .B(n25304), .Z(n13728) );
  XOR U26214 ( .A(n25305), .B(n25306), .Z(n25299) );
  AND U26215 ( .A(n25307), .B(n25308), .Z(n25306) );
  XOR U26216 ( .A(e_input[905]), .B(n25305), .Z(n25308) );
  XNOR U26217 ( .A(n13740), .B(n25305), .Z(n25307) );
  XOR U26218 ( .A(n25309), .B(n25310), .Z(n13740) );
  XOR U26219 ( .A(n25311), .B(n25312), .Z(n25305) );
  AND U26220 ( .A(n25313), .B(n25314), .Z(n25312) );
  XOR U26221 ( .A(e_input[904]), .B(n25311), .Z(n25314) );
  XNOR U26222 ( .A(n13752), .B(n25311), .Z(n25313) );
  XOR U26223 ( .A(n25315), .B(n25316), .Z(n13752) );
  XOR U26224 ( .A(n25317), .B(n25318), .Z(n25311) );
  AND U26225 ( .A(n25319), .B(n25320), .Z(n25318) );
  XOR U26226 ( .A(e_input[903]), .B(n25317), .Z(n25320) );
  XNOR U26227 ( .A(n13764), .B(n25317), .Z(n25319) );
  XOR U26228 ( .A(n25321), .B(n25322), .Z(n13764) );
  XOR U26229 ( .A(n25323), .B(n25324), .Z(n25317) );
  AND U26230 ( .A(n25325), .B(n25326), .Z(n25324) );
  XOR U26231 ( .A(e_input[902]), .B(n25323), .Z(n25326) );
  XNOR U26232 ( .A(n13776), .B(n25323), .Z(n25325) );
  XOR U26233 ( .A(n25327), .B(n25328), .Z(n13776) );
  XOR U26234 ( .A(n25329), .B(n25330), .Z(n25323) );
  AND U26235 ( .A(n25331), .B(n25332), .Z(n25330) );
  XOR U26236 ( .A(e_input[901]), .B(n25329), .Z(n25332) );
  XNOR U26237 ( .A(n13788), .B(n25329), .Z(n25331) );
  XOR U26238 ( .A(n25333), .B(n25334), .Z(n13788) );
  XOR U26239 ( .A(n25335), .B(n25336), .Z(n25329) );
  AND U26240 ( .A(n25337), .B(n25338), .Z(n25336) );
  XOR U26241 ( .A(e_input[900]), .B(n25335), .Z(n25338) );
  XNOR U26242 ( .A(n13800), .B(n25335), .Z(n25337) );
  XOR U26243 ( .A(n25339), .B(n25340), .Z(n13800) );
  XOR U26244 ( .A(n25341), .B(n25342), .Z(n25335) );
  AND U26245 ( .A(n25343), .B(n25344), .Z(n25342) );
  XOR U26246 ( .A(e_input[899]), .B(n25341), .Z(n25344) );
  XNOR U26247 ( .A(n13812), .B(n25341), .Z(n25343) );
  XOR U26248 ( .A(n25345), .B(n25346), .Z(n13812) );
  XOR U26249 ( .A(n25347), .B(n25348), .Z(n25341) );
  AND U26250 ( .A(n25349), .B(n25350), .Z(n25348) );
  XOR U26251 ( .A(e_input[898]), .B(n25347), .Z(n25350) );
  XNOR U26252 ( .A(n13824), .B(n25347), .Z(n25349) );
  XOR U26253 ( .A(n25351), .B(n25352), .Z(n13824) );
  XOR U26254 ( .A(n25353), .B(n25354), .Z(n25347) );
  AND U26255 ( .A(n25355), .B(n25356), .Z(n25354) );
  XOR U26256 ( .A(e_input[897]), .B(n25353), .Z(n25356) );
  XNOR U26257 ( .A(n13836), .B(n25353), .Z(n25355) );
  XOR U26258 ( .A(n25357), .B(n25358), .Z(n13836) );
  XOR U26259 ( .A(n25359), .B(n25360), .Z(n25353) );
  AND U26260 ( .A(n25361), .B(n25362), .Z(n25360) );
  XOR U26261 ( .A(e_input[896]), .B(n25359), .Z(n25362) );
  XNOR U26262 ( .A(n13848), .B(n25359), .Z(n25361) );
  XOR U26263 ( .A(n25363), .B(n25364), .Z(n13848) );
  XOR U26264 ( .A(n25365), .B(n25366), .Z(n25359) );
  AND U26265 ( .A(n25367), .B(n25368), .Z(n25366) );
  XOR U26266 ( .A(e_input[895]), .B(n25365), .Z(n25368) );
  XNOR U26267 ( .A(n13860), .B(n25365), .Z(n25367) );
  XOR U26268 ( .A(n25369), .B(n25370), .Z(n13860) );
  XOR U26269 ( .A(n25371), .B(n25372), .Z(n25365) );
  AND U26270 ( .A(n25373), .B(n25374), .Z(n25372) );
  XOR U26271 ( .A(e_input[894]), .B(n25371), .Z(n25374) );
  XNOR U26272 ( .A(n13872), .B(n25371), .Z(n25373) );
  XOR U26273 ( .A(n25375), .B(n25376), .Z(n13872) );
  XOR U26274 ( .A(n25377), .B(n25378), .Z(n25371) );
  AND U26275 ( .A(n25379), .B(n25380), .Z(n25378) );
  XOR U26276 ( .A(e_input[893]), .B(n25377), .Z(n25380) );
  XNOR U26277 ( .A(n13884), .B(n25377), .Z(n25379) );
  XOR U26278 ( .A(n25381), .B(n25382), .Z(n13884) );
  XOR U26279 ( .A(n25383), .B(n25384), .Z(n25377) );
  AND U26280 ( .A(n25385), .B(n25386), .Z(n25384) );
  XOR U26281 ( .A(e_input[892]), .B(n25383), .Z(n25386) );
  XNOR U26282 ( .A(n13896), .B(n25383), .Z(n25385) );
  XOR U26283 ( .A(n25387), .B(n25388), .Z(n13896) );
  XOR U26284 ( .A(n25389), .B(n25390), .Z(n25383) );
  AND U26285 ( .A(n25391), .B(n25392), .Z(n25390) );
  XOR U26286 ( .A(e_input[891]), .B(n25389), .Z(n25392) );
  XNOR U26287 ( .A(n13908), .B(n25389), .Z(n25391) );
  XOR U26288 ( .A(n25393), .B(n25394), .Z(n13908) );
  XOR U26289 ( .A(n25395), .B(n25396), .Z(n25389) );
  AND U26290 ( .A(n25397), .B(n25398), .Z(n25396) );
  XOR U26291 ( .A(e_input[890]), .B(n25395), .Z(n25398) );
  XNOR U26292 ( .A(n13920), .B(n25395), .Z(n25397) );
  XOR U26293 ( .A(n25399), .B(n25400), .Z(n13920) );
  XOR U26294 ( .A(n25401), .B(n25402), .Z(n25395) );
  AND U26295 ( .A(n25403), .B(n25404), .Z(n25402) );
  XOR U26296 ( .A(e_input[889]), .B(n25401), .Z(n25404) );
  XNOR U26297 ( .A(n13932), .B(n25401), .Z(n25403) );
  XOR U26298 ( .A(n25405), .B(n25406), .Z(n13932) );
  XOR U26299 ( .A(n25407), .B(n25408), .Z(n25401) );
  AND U26300 ( .A(n25409), .B(n25410), .Z(n25408) );
  XOR U26301 ( .A(e_input[888]), .B(n25407), .Z(n25410) );
  XNOR U26302 ( .A(n13944), .B(n25407), .Z(n25409) );
  XOR U26303 ( .A(n25411), .B(n25412), .Z(n13944) );
  XOR U26304 ( .A(n25413), .B(n25414), .Z(n25407) );
  AND U26305 ( .A(n25415), .B(n25416), .Z(n25414) );
  XOR U26306 ( .A(e_input[887]), .B(n25413), .Z(n25416) );
  XNOR U26307 ( .A(n13956), .B(n25413), .Z(n25415) );
  XOR U26308 ( .A(n25417), .B(n25418), .Z(n13956) );
  XOR U26309 ( .A(n25419), .B(n25420), .Z(n25413) );
  AND U26310 ( .A(n25421), .B(n25422), .Z(n25420) );
  XOR U26311 ( .A(e_input[886]), .B(n25419), .Z(n25422) );
  XNOR U26312 ( .A(n13968), .B(n25419), .Z(n25421) );
  XOR U26313 ( .A(n25423), .B(n25424), .Z(n13968) );
  XOR U26314 ( .A(n25425), .B(n25426), .Z(n25419) );
  AND U26315 ( .A(n25427), .B(n25428), .Z(n25426) );
  XOR U26316 ( .A(e_input[885]), .B(n25425), .Z(n25428) );
  XNOR U26317 ( .A(n13980), .B(n25425), .Z(n25427) );
  XOR U26318 ( .A(n25429), .B(n25430), .Z(n13980) );
  XOR U26319 ( .A(n25431), .B(n25432), .Z(n25425) );
  AND U26320 ( .A(n25433), .B(n25434), .Z(n25432) );
  XOR U26321 ( .A(e_input[884]), .B(n25431), .Z(n25434) );
  XNOR U26322 ( .A(n13992), .B(n25431), .Z(n25433) );
  XOR U26323 ( .A(n25435), .B(n25436), .Z(n13992) );
  XOR U26324 ( .A(n25437), .B(n25438), .Z(n25431) );
  AND U26325 ( .A(n25439), .B(n25440), .Z(n25438) );
  XOR U26326 ( .A(e_input[883]), .B(n25437), .Z(n25440) );
  XNOR U26327 ( .A(n14004), .B(n25437), .Z(n25439) );
  XOR U26328 ( .A(n25441), .B(n25442), .Z(n14004) );
  XOR U26329 ( .A(n25443), .B(n25444), .Z(n25437) );
  AND U26330 ( .A(n25445), .B(n25446), .Z(n25444) );
  XOR U26331 ( .A(e_input[882]), .B(n25443), .Z(n25446) );
  XNOR U26332 ( .A(n14016), .B(n25443), .Z(n25445) );
  XOR U26333 ( .A(n25447), .B(n25448), .Z(n14016) );
  XOR U26334 ( .A(n25449), .B(n25450), .Z(n25443) );
  AND U26335 ( .A(n25451), .B(n25452), .Z(n25450) );
  XOR U26336 ( .A(e_input[881]), .B(n25449), .Z(n25452) );
  XNOR U26337 ( .A(n14028), .B(n25449), .Z(n25451) );
  XOR U26338 ( .A(n25453), .B(n25454), .Z(n14028) );
  XOR U26339 ( .A(n25455), .B(n25456), .Z(n25449) );
  AND U26340 ( .A(n25457), .B(n25458), .Z(n25456) );
  XOR U26341 ( .A(e_input[880]), .B(n25455), .Z(n25458) );
  XNOR U26342 ( .A(n14040), .B(n25455), .Z(n25457) );
  XOR U26343 ( .A(n25459), .B(n25460), .Z(n14040) );
  XOR U26344 ( .A(n25461), .B(n25462), .Z(n25455) );
  AND U26345 ( .A(n25463), .B(n25464), .Z(n25462) );
  XOR U26346 ( .A(e_input[879]), .B(n25461), .Z(n25464) );
  XNOR U26347 ( .A(n14052), .B(n25461), .Z(n25463) );
  XOR U26348 ( .A(n25465), .B(n25466), .Z(n14052) );
  XOR U26349 ( .A(n25467), .B(n25468), .Z(n25461) );
  AND U26350 ( .A(n25469), .B(n25470), .Z(n25468) );
  XOR U26351 ( .A(e_input[878]), .B(n25467), .Z(n25470) );
  XNOR U26352 ( .A(n14064), .B(n25467), .Z(n25469) );
  XOR U26353 ( .A(n25471), .B(n25472), .Z(n14064) );
  XOR U26354 ( .A(n25473), .B(n25474), .Z(n25467) );
  AND U26355 ( .A(n25475), .B(n25476), .Z(n25474) );
  XOR U26356 ( .A(e_input[877]), .B(n25473), .Z(n25476) );
  XNOR U26357 ( .A(n14076), .B(n25473), .Z(n25475) );
  XOR U26358 ( .A(n25477), .B(n25478), .Z(n14076) );
  XOR U26359 ( .A(n25479), .B(n25480), .Z(n25473) );
  AND U26360 ( .A(n25481), .B(n25482), .Z(n25480) );
  XOR U26361 ( .A(e_input[876]), .B(n25479), .Z(n25482) );
  XNOR U26362 ( .A(n14088), .B(n25479), .Z(n25481) );
  XOR U26363 ( .A(n25483), .B(n25484), .Z(n14088) );
  XOR U26364 ( .A(n25485), .B(n25486), .Z(n25479) );
  AND U26365 ( .A(n25487), .B(n25488), .Z(n25486) );
  XOR U26366 ( .A(e_input[875]), .B(n25485), .Z(n25488) );
  XNOR U26367 ( .A(n14100), .B(n25485), .Z(n25487) );
  XOR U26368 ( .A(n25489), .B(n25490), .Z(n14100) );
  XOR U26369 ( .A(n25491), .B(n25492), .Z(n25485) );
  AND U26370 ( .A(n25493), .B(n25494), .Z(n25492) );
  XOR U26371 ( .A(e_input[874]), .B(n25491), .Z(n25494) );
  XNOR U26372 ( .A(n14112), .B(n25491), .Z(n25493) );
  XOR U26373 ( .A(n25495), .B(n25496), .Z(n14112) );
  XOR U26374 ( .A(n25497), .B(n25498), .Z(n25491) );
  AND U26375 ( .A(n25499), .B(n25500), .Z(n25498) );
  XOR U26376 ( .A(e_input[873]), .B(n25497), .Z(n25500) );
  XNOR U26377 ( .A(n14124), .B(n25497), .Z(n25499) );
  XOR U26378 ( .A(n25501), .B(n25502), .Z(n14124) );
  XOR U26379 ( .A(n25503), .B(n25504), .Z(n25497) );
  AND U26380 ( .A(n25505), .B(n25506), .Z(n25504) );
  XOR U26381 ( .A(e_input[872]), .B(n25503), .Z(n25506) );
  XNOR U26382 ( .A(n14136), .B(n25503), .Z(n25505) );
  XOR U26383 ( .A(n25507), .B(n25508), .Z(n14136) );
  XOR U26384 ( .A(n25509), .B(n25510), .Z(n25503) );
  AND U26385 ( .A(n25511), .B(n25512), .Z(n25510) );
  XOR U26386 ( .A(e_input[871]), .B(n25509), .Z(n25512) );
  XNOR U26387 ( .A(n14148), .B(n25509), .Z(n25511) );
  XOR U26388 ( .A(n25513), .B(n25514), .Z(n14148) );
  XOR U26389 ( .A(n25515), .B(n25516), .Z(n25509) );
  AND U26390 ( .A(n25517), .B(n25518), .Z(n25516) );
  XOR U26391 ( .A(e_input[870]), .B(n25515), .Z(n25518) );
  XNOR U26392 ( .A(n14160), .B(n25515), .Z(n25517) );
  XOR U26393 ( .A(n25519), .B(n25520), .Z(n14160) );
  XOR U26394 ( .A(n25521), .B(n25522), .Z(n25515) );
  AND U26395 ( .A(n25523), .B(n25524), .Z(n25522) );
  XOR U26396 ( .A(e_input[869]), .B(n25521), .Z(n25524) );
  XNOR U26397 ( .A(n14172), .B(n25521), .Z(n25523) );
  XOR U26398 ( .A(n25525), .B(n25526), .Z(n14172) );
  XOR U26399 ( .A(n25527), .B(n25528), .Z(n25521) );
  AND U26400 ( .A(n25529), .B(n25530), .Z(n25528) );
  XOR U26401 ( .A(e_input[868]), .B(n25527), .Z(n25530) );
  XNOR U26402 ( .A(n14184), .B(n25527), .Z(n25529) );
  XOR U26403 ( .A(n25531), .B(n25532), .Z(n14184) );
  XOR U26404 ( .A(n25533), .B(n25534), .Z(n25527) );
  AND U26405 ( .A(n25535), .B(n25536), .Z(n25534) );
  XOR U26406 ( .A(e_input[867]), .B(n25533), .Z(n25536) );
  XNOR U26407 ( .A(n14196), .B(n25533), .Z(n25535) );
  XOR U26408 ( .A(n25537), .B(n25538), .Z(n14196) );
  XOR U26409 ( .A(n25539), .B(n25540), .Z(n25533) );
  AND U26410 ( .A(n25541), .B(n25542), .Z(n25540) );
  XOR U26411 ( .A(e_input[866]), .B(n25539), .Z(n25542) );
  XNOR U26412 ( .A(n14208), .B(n25539), .Z(n25541) );
  XOR U26413 ( .A(n25543), .B(n25544), .Z(n14208) );
  XOR U26414 ( .A(n25545), .B(n25546), .Z(n25539) );
  AND U26415 ( .A(n25547), .B(n25548), .Z(n25546) );
  XOR U26416 ( .A(e_input[865]), .B(n25545), .Z(n25548) );
  XNOR U26417 ( .A(n14220), .B(n25545), .Z(n25547) );
  XOR U26418 ( .A(n25549), .B(n25550), .Z(n14220) );
  XOR U26419 ( .A(n25551), .B(n25552), .Z(n25545) );
  AND U26420 ( .A(n25553), .B(n25554), .Z(n25552) );
  XOR U26421 ( .A(e_input[864]), .B(n25551), .Z(n25554) );
  XNOR U26422 ( .A(n14232), .B(n25551), .Z(n25553) );
  XOR U26423 ( .A(n25555), .B(n25556), .Z(n14232) );
  XOR U26424 ( .A(n25557), .B(n25558), .Z(n25551) );
  AND U26425 ( .A(n25559), .B(n25560), .Z(n25558) );
  XOR U26426 ( .A(e_input[863]), .B(n25557), .Z(n25560) );
  XNOR U26427 ( .A(n14244), .B(n25557), .Z(n25559) );
  XOR U26428 ( .A(n25561), .B(n25562), .Z(n14244) );
  XOR U26429 ( .A(n25563), .B(n25564), .Z(n25557) );
  AND U26430 ( .A(n25565), .B(n25566), .Z(n25564) );
  XOR U26431 ( .A(e_input[862]), .B(n25563), .Z(n25566) );
  XNOR U26432 ( .A(n14256), .B(n25563), .Z(n25565) );
  XOR U26433 ( .A(n25567), .B(n25568), .Z(n14256) );
  XOR U26434 ( .A(n25569), .B(n25570), .Z(n25563) );
  AND U26435 ( .A(n25571), .B(n25572), .Z(n25570) );
  XOR U26436 ( .A(e_input[861]), .B(n25569), .Z(n25572) );
  XNOR U26437 ( .A(n14268), .B(n25569), .Z(n25571) );
  XOR U26438 ( .A(n25573), .B(n25574), .Z(n14268) );
  XOR U26439 ( .A(n25575), .B(n25576), .Z(n25569) );
  AND U26440 ( .A(n25577), .B(n25578), .Z(n25576) );
  XOR U26441 ( .A(e_input[860]), .B(n25575), .Z(n25578) );
  XNOR U26442 ( .A(n14280), .B(n25575), .Z(n25577) );
  XOR U26443 ( .A(n25579), .B(n25580), .Z(n14280) );
  XOR U26444 ( .A(n25581), .B(n25582), .Z(n25575) );
  AND U26445 ( .A(n25583), .B(n25584), .Z(n25582) );
  XOR U26446 ( .A(e_input[859]), .B(n25581), .Z(n25584) );
  XNOR U26447 ( .A(n14292), .B(n25581), .Z(n25583) );
  XOR U26448 ( .A(n25585), .B(n25586), .Z(n14292) );
  XOR U26449 ( .A(n25587), .B(n25588), .Z(n25581) );
  AND U26450 ( .A(n25589), .B(n25590), .Z(n25588) );
  XOR U26451 ( .A(e_input[858]), .B(n25587), .Z(n25590) );
  XNOR U26452 ( .A(n14304), .B(n25587), .Z(n25589) );
  XOR U26453 ( .A(n25591), .B(n25592), .Z(n14304) );
  XOR U26454 ( .A(n25593), .B(n25594), .Z(n25587) );
  AND U26455 ( .A(n25595), .B(n25596), .Z(n25594) );
  XOR U26456 ( .A(e_input[857]), .B(n25593), .Z(n25596) );
  XNOR U26457 ( .A(n14316), .B(n25593), .Z(n25595) );
  XOR U26458 ( .A(n25597), .B(n25598), .Z(n14316) );
  XOR U26459 ( .A(n25599), .B(n25600), .Z(n25593) );
  AND U26460 ( .A(n25601), .B(n25602), .Z(n25600) );
  XOR U26461 ( .A(e_input[856]), .B(n25599), .Z(n25602) );
  XNOR U26462 ( .A(n14328), .B(n25599), .Z(n25601) );
  XOR U26463 ( .A(n25603), .B(n25604), .Z(n14328) );
  XOR U26464 ( .A(n25605), .B(n25606), .Z(n25599) );
  AND U26465 ( .A(n25607), .B(n25608), .Z(n25606) );
  XOR U26466 ( .A(e_input[855]), .B(n25605), .Z(n25608) );
  XNOR U26467 ( .A(n14340), .B(n25605), .Z(n25607) );
  XOR U26468 ( .A(n25609), .B(n25610), .Z(n14340) );
  XOR U26469 ( .A(n25611), .B(n25612), .Z(n25605) );
  AND U26470 ( .A(n25613), .B(n25614), .Z(n25612) );
  XOR U26471 ( .A(e_input[854]), .B(n25611), .Z(n25614) );
  XNOR U26472 ( .A(n14352), .B(n25611), .Z(n25613) );
  XOR U26473 ( .A(n25615), .B(n25616), .Z(n14352) );
  XOR U26474 ( .A(n25617), .B(n25618), .Z(n25611) );
  AND U26475 ( .A(n25619), .B(n25620), .Z(n25618) );
  XOR U26476 ( .A(e_input[853]), .B(n25617), .Z(n25620) );
  XNOR U26477 ( .A(n14364), .B(n25617), .Z(n25619) );
  XOR U26478 ( .A(n25621), .B(n25622), .Z(n14364) );
  XOR U26479 ( .A(n25623), .B(n25624), .Z(n25617) );
  AND U26480 ( .A(n25625), .B(n25626), .Z(n25624) );
  XOR U26481 ( .A(e_input[852]), .B(n25623), .Z(n25626) );
  XNOR U26482 ( .A(n14376), .B(n25623), .Z(n25625) );
  XOR U26483 ( .A(n25627), .B(n25628), .Z(n14376) );
  XOR U26484 ( .A(n25629), .B(n25630), .Z(n25623) );
  AND U26485 ( .A(n25631), .B(n25632), .Z(n25630) );
  XOR U26486 ( .A(e_input[851]), .B(n25629), .Z(n25632) );
  XNOR U26487 ( .A(n14388), .B(n25629), .Z(n25631) );
  XOR U26488 ( .A(n25633), .B(n25634), .Z(n14388) );
  XOR U26489 ( .A(n25635), .B(n25636), .Z(n25629) );
  AND U26490 ( .A(n25637), .B(n25638), .Z(n25636) );
  XOR U26491 ( .A(e_input[850]), .B(n25635), .Z(n25638) );
  XNOR U26492 ( .A(n14400), .B(n25635), .Z(n25637) );
  XOR U26493 ( .A(n25639), .B(n25640), .Z(n14400) );
  XOR U26494 ( .A(n25641), .B(n25642), .Z(n25635) );
  AND U26495 ( .A(n25643), .B(n25644), .Z(n25642) );
  XOR U26496 ( .A(e_input[849]), .B(n25641), .Z(n25644) );
  XNOR U26497 ( .A(n14412), .B(n25641), .Z(n25643) );
  XOR U26498 ( .A(n25645), .B(n25646), .Z(n14412) );
  XOR U26499 ( .A(n25647), .B(n25648), .Z(n25641) );
  AND U26500 ( .A(n25649), .B(n25650), .Z(n25648) );
  XOR U26501 ( .A(e_input[848]), .B(n25647), .Z(n25650) );
  XNOR U26502 ( .A(n14424), .B(n25647), .Z(n25649) );
  XOR U26503 ( .A(n25651), .B(n25652), .Z(n14424) );
  XOR U26504 ( .A(n25653), .B(n25654), .Z(n25647) );
  AND U26505 ( .A(n25655), .B(n25656), .Z(n25654) );
  XOR U26506 ( .A(e_input[847]), .B(n25653), .Z(n25656) );
  XNOR U26507 ( .A(n14436), .B(n25653), .Z(n25655) );
  XOR U26508 ( .A(n25657), .B(n25658), .Z(n14436) );
  XOR U26509 ( .A(n25659), .B(n25660), .Z(n25653) );
  AND U26510 ( .A(n25661), .B(n25662), .Z(n25660) );
  XOR U26511 ( .A(e_input[846]), .B(n25659), .Z(n25662) );
  XNOR U26512 ( .A(n14448), .B(n25659), .Z(n25661) );
  XOR U26513 ( .A(n25663), .B(n25664), .Z(n14448) );
  XOR U26514 ( .A(n25665), .B(n25666), .Z(n25659) );
  AND U26515 ( .A(n25667), .B(n25668), .Z(n25666) );
  XOR U26516 ( .A(e_input[845]), .B(n25665), .Z(n25668) );
  XNOR U26517 ( .A(n14460), .B(n25665), .Z(n25667) );
  XOR U26518 ( .A(n25669), .B(n25670), .Z(n14460) );
  XOR U26519 ( .A(n25671), .B(n25672), .Z(n25665) );
  AND U26520 ( .A(n25673), .B(n25674), .Z(n25672) );
  XOR U26521 ( .A(e_input[844]), .B(n25671), .Z(n25674) );
  XNOR U26522 ( .A(n14472), .B(n25671), .Z(n25673) );
  XOR U26523 ( .A(n25675), .B(n25676), .Z(n14472) );
  XOR U26524 ( .A(n25677), .B(n25678), .Z(n25671) );
  AND U26525 ( .A(n25679), .B(n25680), .Z(n25678) );
  XOR U26526 ( .A(e_input[843]), .B(n25677), .Z(n25680) );
  XNOR U26527 ( .A(n14484), .B(n25677), .Z(n25679) );
  XOR U26528 ( .A(n25681), .B(n25682), .Z(n14484) );
  XOR U26529 ( .A(n25683), .B(n25684), .Z(n25677) );
  AND U26530 ( .A(n25685), .B(n25686), .Z(n25684) );
  XOR U26531 ( .A(e_input[842]), .B(n25683), .Z(n25686) );
  XNOR U26532 ( .A(n14496), .B(n25683), .Z(n25685) );
  XOR U26533 ( .A(n25687), .B(n25688), .Z(n14496) );
  XOR U26534 ( .A(n25689), .B(n25690), .Z(n25683) );
  AND U26535 ( .A(n25691), .B(n25692), .Z(n25690) );
  XOR U26536 ( .A(e_input[841]), .B(n25689), .Z(n25692) );
  XNOR U26537 ( .A(n14508), .B(n25689), .Z(n25691) );
  XOR U26538 ( .A(n25693), .B(n25694), .Z(n14508) );
  XOR U26539 ( .A(n25695), .B(n25696), .Z(n25689) );
  AND U26540 ( .A(n25697), .B(n25698), .Z(n25696) );
  XOR U26541 ( .A(e_input[840]), .B(n25695), .Z(n25698) );
  XNOR U26542 ( .A(n14520), .B(n25695), .Z(n25697) );
  XOR U26543 ( .A(n25699), .B(n25700), .Z(n14520) );
  XOR U26544 ( .A(n25701), .B(n25702), .Z(n25695) );
  AND U26545 ( .A(n25703), .B(n25704), .Z(n25702) );
  XOR U26546 ( .A(e_input[839]), .B(n25701), .Z(n25704) );
  XNOR U26547 ( .A(n14532), .B(n25701), .Z(n25703) );
  XOR U26548 ( .A(n25705), .B(n25706), .Z(n14532) );
  XOR U26549 ( .A(n25707), .B(n25708), .Z(n25701) );
  AND U26550 ( .A(n25709), .B(n25710), .Z(n25708) );
  XOR U26551 ( .A(e_input[838]), .B(n25707), .Z(n25710) );
  XNOR U26552 ( .A(n14544), .B(n25707), .Z(n25709) );
  XOR U26553 ( .A(n25711), .B(n25712), .Z(n14544) );
  XOR U26554 ( .A(n25713), .B(n25714), .Z(n25707) );
  AND U26555 ( .A(n25715), .B(n25716), .Z(n25714) );
  XOR U26556 ( .A(e_input[837]), .B(n25713), .Z(n25716) );
  XNOR U26557 ( .A(n14556), .B(n25713), .Z(n25715) );
  XOR U26558 ( .A(n25717), .B(n25718), .Z(n14556) );
  XOR U26559 ( .A(n25719), .B(n25720), .Z(n25713) );
  AND U26560 ( .A(n25721), .B(n25722), .Z(n25720) );
  XOR U26561 ( .A(e_input[836]), .B(n25719), .Z(n25722) );
  XNOR U26562 ( .A(n14568), .B(n25719), .Z(n25721) );
  XOR U26563 ( .A(n25723), .B(n25724), .Z(n14568) );
  XOR U26564 ( .A(n25725), .B(n25726), .Z(n25719) );
  AND U26565 ( .A(n25727), .B(n25728), .Z(n25726) );
  XOR U26566 ( .A(e_input[835]), .B(n25725), .Z(n25728) );
  XNOR U26567 ( .A(n14580), .B(n25725), .Z(n25727) );
  XOR U26568 ( .A(n25729), .B(n25730), .Z(n14580) );
  XOR U26569 ( .A(n25731), .B(n25732), .Z(n25725) );
  AND U26570 ( .A(n25733), .B(n25734), .Z(n25732) );
  XOR U26571 ( .A(e_input[834]), .B(n25731), .Z(n25734) );
  XNOR U26572 ( .A(n14592), .B(n25731), .Z(n25733) );
  XOR U26573 ( .A(n25735), .B(n25736), .Z(n14592) );
  XOR U26574 ( .A(n25737), .B(n25738), .Z(n25731) );
  AND U26575 ( .A(n25739), .B(n25740), .Z(n25738) );
  XOR U26576 ( .A(e_input[833]), .B(n25737), .Z(n25740) );
  XNOR U26577 ( .A(n14604), .B(n25737), .Z(n25739) );
  XOR U26578 ( .A(n25741), .B(n25742), .Z(n14604) );
  XOR U26579 ( .A(n25743), .B(n25744), .Z(n25737) );
  AND U26580 ( .A(n25745), .B(n25746), .Z(n25744) );
  XOR U26581 ( .A(e_input[832]), .B(n25743), .Z(n25746) );
  XNOR U26582 ( .A(n14616), .B(n25743), .Z(n25745) );
  XOR U26583 ( .A(n25747), .B(n25748), .Z(n14616) );
  XOR U26584 ( .A(n25749), .B(n25750), .Z(n25743) );
  AND U26585 ( .A(n25751), .B(n25752), .Z(n25750) );
  XOR U26586 ( .A(e_input[831]), .B(n25749), .Z(n25752) );
  XNOR U26587 ( .A(n14628), .B(n25749), .Z(n25751) );
  XOR U26588 ( .A(n25753), .B(n25754), .Z(n14628) );
  XOR U26589 ( .A(n25755), .B(n25756), .Z(n25749) );
  AND U26590 ( .A(n25757), .B(n25758), .Z(n25756) );
  XOR U26591 ( .A(e_input[830]), .B(n25755), .Z(n25758) );
  XNOR U26592 ( .A(n14640), .B(n25755), .Z(n25757) );
  XOR U26593 ( .A(n25759), .B(n25760), .Z(n14640) );
  XOR U26594 ( .A(n25761), .B(n25762), .Z(n25755) );
  AND U26595 ( .A(n25763), .B(n25764), .Z(n25762) );
  XOR U26596 ( .A(e_input[829]), .B(n25761), .Z(n25764) );
  XNOR U26597 ( .A(n14652), .B(n25761), .Z(n25763) );
  XOR U26598 ( .A(n25765), .B(n25766), .Z(n14652) );
  XOR U26599 ( .A(n25767), .B(n25768), .Z(n25761) );
  AND U26600 ( .A(n25769), .B(n25770), .Z(n25768) );
  XOR U26601 ( .A(e_input[828]), .B(n25767), .Z(n25770) );
  XNOR U26602 ( .A(n14664), .B(n25767), .Z(n25769) );
  XOR U26603 ( .A(n25771), .B(n25772), .Z(n14664) );
  XOR U26604 ( .A(n25773), .B(n25774), .Z(n25767) );
  AND U26605 ( .A(n25775), .B(n25776), .Z(n25774) );
  XOR U26606 ( .A(e_input[827]), .B(n25773), .Z(n25776) );
  XNOR U26607 ( .A(n14676), .B(n25773), .Z(n25775) );
  XOR U26608 ( .A(n25777), .B(n25778), .Z(n14676) );
  XOR U26609 ( .A(n25779), .B(n25780), .Z(n25773) );
  AND U26610 ( .A(n25781), .B(n25782), .Z(n25780) );
  XOR U26611 ( .A(e_input[826]), .B(n25779), .Z(n25782) );
  XNOR U26612 ( .A(n14688), .B(n25779), .Z(n25781) );
  XOR U26613 ( .A(n25783), .B(n25784), .Z(n14688) );
  XOR U26614 ( .A(n25785), .B(n25786), .Z(n25779) );
  AND U26615 ( .A(n25787), .B(n25788), .Z(n25786) );
  XOR U26616 ( .A(e_input[825]), .B(n25785), .Z(n25788) );
  XNOR U26617 ( .A(n14700), .B(n25785), .Z(n25787) );
  XOR U26618 ( .A(n25789), .B(n25790), .Z(n14700) );
  XOR U26619 ( .A(n25791), .B(n25792), .Z(n25785) );
  AND U26620 ( .A(n25793), .B(n25794), .Z(n25792) );
  XOR U26621 ( .A(e_input[824]), .B(n25791), .Z(n25794) );
  XNOR U26622 ( .A(n14712), .B(n25791), .Z(n25793) );
  XOR U26623 ( .A(n25795), .B(n25796), .Z(n14712) );
  XOR U26624 ( .A(n25797), .B(n25798), .Z(n25791) );
  AND U26625 ( .A(n25799), .B(n25800), .Z(n25798) );
  XOR U26626 ( .A(e_input[823]), .B(n25797), .Z(n25800) );
  XNOR U26627 ( .A(n14724), .B(n25797), .Z(n25799) );
  XOR U26628 ( .A(n25801), .B(n25802), .Z(n14724) );
  XOR U26629 ( .A(n25803), .B(n25804), .Z(n25797) );
  AND U26630 ( .A(n25805), .B(n25806), .Z(n25804) );
  XOR U26631 ( .A(e_input[822]), .B(n25803), .Z(n25806) );
  XNOR U26632 ( .A(n14736), .B(n25803), .Z(n25805) );
  XOR U26633 ( .A(n25807), .B(n25808), .Z(n14736) );
  XOR U26634 ( .A(n25809), .B(n25810), .Z(n25803) );
  AND U26635 ( .A(n25811), .B(n25812), .Z(n25810) );
  XOR U26636 ( .A(e_input[821]), .B(n25809), .Z(n25812) );
  XNOR U26637 ( .A(n14748), .B(n25809), .Z(n25811) );
  XOR U26638 ( .A(n25813), .B(n25814), .Z(n14748) );
  XOR U26639 ( .A(n25815), .B(n25816), .Z(n25809) );
  AND U26640 ( .A(n25817), .B(n25818), .Z(n25816) );
  XOR U26641 ( .A(e_input[820]), .B(n25815), .Z(n25818) );
  XNOR U26642 ( .A(n14760), .B(n25815), .Z(n25817) );
  XOR U26643 ( .A(n25819), .B(n25820), .Z(n14760) );
  XOR U26644 ( .A(n25821), .B(n25822), .Z(n25815) );
  AND U26645 ( .A(n25823), .B(n25824), .Z(n25822) );
  XOR U26646 ( .A(e_input[819]), .B(n25821), .Z(n25824) );
  XNOR U26647 ( .A(n14772), .B(n25821), .Z(n25823) );
  XOR U26648 ( .A(n25825), .B(n25826), .Z(n14772) );
  XOR U26649 ( .A(n25827), .B(n25828), .Z(n25821) );
  AND U26650 ( .A(n25829), .B(n25830), .Z(n25828) );
  XOR U26651 ( .A(e_input[818]), .B(n25827), .Z(n25830) );
  XNOR U26652 ( .A(n14784), .B(n25827), .Z(n25829) );
  XOR U26653 ( .A(n25831), .B(n25832), .Z(n14784) );
  XOR U26654 ( .A(n25833), .B(n25834), .Z(n25827) );
  AND U26655 ( .A(n25835), .B(n25836), .Z(n25834) );
  XOR U26656 ( .A(e_input[817]), .B(n25833), .Z(n25836) );
  XNOR U26657 ( .A(n14796), .B(n25833), .Z(n25835) );
  XOR U26658 ( .A(n25837), .B(n25838), .Z(n14796) );
  XOR U26659 ( .A(n25839), .B(n25840), .Z(n25833) );
  AND U26660 ( .A(n25841), .B(n25842), .Z(n25840) );
  XOR U26661 ( .A(e_input[816]), .B(n25839), .Z(n25842) );
  XNOR U26662 ( .A(n14808), .B(n25839), .Z(n25841) );
  XOR U26663 ( .A(n25843), .B(n25844), .Z(n14808) );
  XOR U26664 ( .A(n25845), .B(n25846), .Z(n25839) );
  AND U26665 ( .A(n25847), .B(n25848), .Z(n25846) );
  XOR U26666 ( .A(e_input[815]), .B(n25845), .Z(n25848) );
  XNOR U26667 ( .A(n14820), .B(n25845), .Z(n25847) );
  XOR U26668 ( .A(n25849), .B(n25850), .Z(n14820) );
  XOR U26669 ( .A(n25851), .B(n25852), .Z(n25845) );
  AND U26670 ( .A(n25853), .B(n25854), .Z(n25852) );
  XOR U26671 ( .A(e_input[814]), .B(n25851), .Z(n25854) );
  XNOR U26672 ( .A(n14832), .B(n25851), .Z(n25853) );
  XOR U26673 ( .A(n25855), .B(n25856), .Z(n14832) );
  XOR U26674 ( .A(n25857), .B(n25858), .Z(n25851) );
  AND U26675 ( .A(n25859), .B(n25860), .Z(n25858) );
  XOR U26676 ( .A(e_input[813]), .B(n25857), .Z(n25860) );
  XNOR U26677 ( .A(n14844), .B(n25857), .Z(n25859) );
  XOR U26678 ( .A(n25861), .B(n25862), .Z(n14844) );
  XOR U26679 ( .A(n25863), .B(n25864), .Z(n25857) );
  AND U26680 ( .A(n25865), .B(n25866), .Z(n25864) );
  XOR U26681 ( .A(e_input[812]), .B(n25863), .Z(n25866) );
  XNOR U26682 ( .A(n14856), .B(n25863), .Z(n25865) );
  XOR U26683 ( .A(n25867), .B(n25868), .Z(n14856) );
  XOR U26684 ( .A(n25869), .B(n25870), .Z(n25863) );
  AND U26685 ( .A(n25871), .B(n25872), .Z(n25870) );
  XOR U26686 ( .A(e_input[811]), .B(n25869), .Z(n25872) );
  XNOR U26687 ( .A(n14868), .B(n25869), .Z(n25871) );
  XOR U26688 ( .A(n25873), .B(n25874), .Z(n14868) );
  XOR U26689 ( .A(n25875), .B(n25876), .Z(n25869) );
  AND U26690 ( .A(n25877), .B(n25878), .Z(n25876) );
  XOR U26691 ( .A(e_input[810]), .B(n25875), .Z(n25878) );
  XNOR U26692 ( .A(n14880), .B(n25875), .Z(n25877) );
  XOR U26693 ( .A(n25879), .B(n25880), .Z(n14880) );
  XOR U26694 ( .A(n25881), .B(n25882), .Z(n25875) );
  AND U26695 ( .A(n25883), .B(n25884), .Z(n25882) );
  XOR U26696 ( .A(e_input[809]), .B(n25881), .Z(n25884) );
  XNOR U26697 ( .A(n14892), .B(n25881), .Z(n25883) );
  XOR U26698 ( .A(n25885), .B(n25886), .Z(n14892) );
  XOR U26699 ( .A(n25887), .B(n25888), .Z(n25881) );
  AND U26700 ( .A(n25889), .B(n25890), .Z(n25888) );
  XOR U26701 ( .A(e_input[808]), .B(n25887), .Z(n25890) );
  XNOR U26702 ( .A(n14904), .B(n25887), .Z(n25889) );
  XOR U26703 ( .A(n25891), .B(n25892), .Z(n14904) );
  XOR U26704 ( .A(n25893), .B(n25894), .Z(n25887) );
  AND U26705 ( .A(n25895), .B(n25896), .Z(n25894) );
  XOR U26706 ( .A(e_input[807]), .B(n25893), .Z(n25896) );
  XNOR U26707 ( .A(n14916), .B(n25893), .Z(n25895) );
  XOR U26708 ( .A(n25897), .B(n25898), .Z(n14916) );
  XOR U26709 ( .A(n25899), .B(n25900), .Z(n25893) );
  AND U26710 ( .A(n25901), .B(n25902), .Z(n25900) );
  XOR U26711 ( .A(e_input[806]), .B(n25899), .Z(n25902) );
  XNOR U26712 ( .A(n14928), .B(n25899), .Z(n25901) );
  XOR U26713 ( .A(n25903), .B(n25904), .Z(n14928) );
  XOR U26714 ( .A(n25905), .B(n25906), .Z(n25899) );
  AND U26715 ( .A(n25907), .B(n25908), .Z(n25906) );
  XOR U26716 ( .A(e_input[805]), .B(n25905), .Z(n25908) );
  XNOR U26717 ( .A(n14940), .B(n25905), .Z(n25907) );
  XOR U26718 ( .A(n25909), .B(n25910), .Z(n14940) );
  XOR U26719 ( .A(n25911), .B(n25912), .Z(n25905) );
  AND U26720 ( .A(n25913), .B(n25914), .Z(n25912) );
  XOR U26721 ( .A(e_input[804]), .B(n25911), .Z(n25914) );
  XNOR U26722 ( .A(n14952), .B(n25911), .Z(n25913) );
  XOR U26723 ( .A(n25915), .B(n25916), .Z(n14952) );
  XOR U26724 ( .A(n25917), .B(n25918), .Z(n25911) );
  AND U26725 ( .A(n25919), .B(n25920), .Z(n25918) );
  XOR U26726 ( .A(e_input[803]), .B(n25917), .Z(n25920) );
  XNOR U26727 ( .A(n14964), .B(n25917), .Z(n25919) );
  XOR U26728 ( .A(n25921), .B(n25922), .Z(n14964) );
  XOR U26729 ( .A(n25923), .B(n25924), .Z(n25917) );
  AND U26730 ( .A(n25925), .B(n25926), .Z(n25924) );
  XOR U26731 ( .A(e_input[802]), .B(n25923), .Z(n25926) );
  XNOR U26732 ( .A(n14976), .B(n25923), .Z(n25925) );
  XOR U26733 ( .A(n25927), .B(n25928), .Z(n14976) );
  XOR U26734 ( .A(n25929), .B(n25930), .Z(n25923) );
  AND U26735 ( .A(n25931), .B(n25932), .Z(n25930) );
  XOR U26736 ( .A(e_input[801]), .B(n25929), .Z(n25932) );
  XNOR U26737 ( .A(n14988), .B(n25929), .Z(n25931) );
  XOR U26738 ( .A(n25933), .B(n25934), .Z(n14988) );
  XOR U26739 ( .A(n25935), .B(n25936), .Z(n25929) );
  AND U26740 ( .A(n25937), .B(n25938), .Z(n25936) );
  XOR U26741 ( .A(e_input[800]), .B(n25935), .Z(n25938) );
  XNOR U26742 ( .A(n15000), .B(n25935), .Z(n25937) );
  XOR U26743 ( .A(n25939), .B(n25940), .Z(n15000) );
  XOR U26744 ( .A(n25941), .B(n25942), .Z(n25935) );
  AND U26745 ( .A(n25943), .B(n25944), .Z(n25942) );
  XOR U26746 ( .A(e_input[799]), .B(n25941), .Z(n25944) );
  XNOR U26747 ( .A(n15012), .B(n25941), .Z(n25943) );
  XOR U26748 ( .A(n25945), .B(n25946), .Z(n15012) );
  XOR U26749 ( .A(n25947), .B(n25948), .Z(n25941) );
  AND U26750 ( .A(n25949), .B(n25950), .Z(n25948) );
  XOR U26751 ( .A(e_input[798]), .B(n25947), .Z(n25950) );
  XNOR U26752 ( .A(n15024), .B(n25947), .Z(n25949) );
  XOR U26753 ( .A(n25951), .B(n25952), .Z(n15024) );
  XOR U26754 ( .A(n25953), .B(n25954), .Z(n25947) );
  AND U26755 ( .A(n25955), .B(n25956), .Z(n25954) );
  XOR U26756 ( .A(e_input[797]), .B(n25953), .Z(n25956) );
  XNOR U26757 ( .A(n15036), .B(n25953), .Z(n25955) );
  XOR U26758 ( .A(n25957), .B(n25958), .Z(n15036) );
  XOR U26759 ( .A(n25959), .B(n25960), .Z(n25953) );
  AND U26760 ( .A(n25961), .B(n25962), .Z(n25960) );
  XOR U26761 ( .A(e_input[796]), .B(n25959), .Z(n25962) );
  XNOR U26762 ( .A(n15048), .B(n25959), .Z(n25961) );
  XOR U26763 ( .A(n25963), .B(n25964), .Z(n15048) );
  XOR U26764 ( .A(n25965), .B(n25966), .Z(n25959) );
  AND U26765 ( .A(n25967), .B(n25968), .Z(n25966) );
  XOR U26766 ( .A(e_input[795]), .B(n25965), .Z(n25968) );
  XNOR U26767 ( .A(n15060), .B(n25965), .Z(n25967) );
  XOR U26768 ( .A(n25969), .B(n25970), .Z(n15060) );
  XOR U26769 ( .A(n25971), .B(n25972), .Z(n25965) );
  AND U26770 ( .A(n25973), .B(n25974), .Z(n25972) );
  XOR U26771 ( .A(e_input[794]), .B(n25971), .Z(n25974) );
  XNOR U26772 ( .A(n15072), .B(n25971), .Z(n25973) );
  XOR U26773 ( .A(n25975), .B(n25976), .Z(n15072) );
  XOR U26774 ( .A(n25977), .B(n25978), .Z(n25971) );
  AND U26775 ( .A(n25979), .B(n25980), .Z(n25978) );
  XOR U26776 ( .A(e_input[793]), .B(n25977), .Z(n25980) );
  XNOR U26777 ( .A(n15084), .B(n25977), .Z(n25979) );
  XOR U26778 ( .A(n25981), .B(n25982), .Z(n15084) );
  XOR U26779 ( .A(n25983), .B(n25984), .Z(n25977) );
  AND U26780 ( .A(n25985), .B(n25986), .Z(n25984) );
  XOR U26781 ( .A(e_input[792]), .B(n25983), .Z(n25986) );
  XNOR U26782 ( .A(n15096), .B(n25983), .Z(n25985) );
  XOR U26783 ( .A(n25987), .B(n25988), .Z(n15096) );
  XOR U26784 ( .A(n25989), .B(n25990), .Z(n25983) );
  AND U26785 ( .A(n25991), .B(n25992), .Z(n25990) );
  XOR U26786 ( .A(e_input[791]), .B(n25989), .Z(n25992) );
  XNOR U26787 ( .A(n15108), .B(n25989), .Z(n25991) );
  XOR U26788 ( .A(n25993), .B(n25994), .Z(n15108) );
  XOR U26789 ( .A(n25995), .B(n25996), .Z(n25989) );
  AND U26790 ( .A(n25997), .B(n25998), .Z(n25996) );
  XOR U26791 ( .A(e_input[790]), .B(n25995), .Z(n25998) );
  XNOR U26792 ( .A(n15120), .B(n25995), .Z(n25997) );
  XOR U26793 ( .A(n25999), .B(n26000), .Z(n15120) );
  XOR U26794 ( .A(n26001), .B(n26002), .Z(n25995) );
  AND U26795 ( .A(n26003), .B(n26004), .Z(n26002) );
  XOR U26796 ( .A(e_input[789]), .B(n26001), .Z(n26004) );
  XNOR U26797 ( .A(n15132), .B(n26001), .Z(n26003) );
  XOR U26798 ( .A(n26005), .B(n26006), .Z(n15132) );
  XOR U26799 ( .A(n26007), .B(n26008), .Z(n26001) );
  AND U26800 ( .A(n26009), .B(n26010), .Z(n26008) );
  XOR U26801 ( .A(e_input[788]), .B(n26007), .Z(n26010) );
  XNOR U26802 ( .A(n15144), .B(n26007), .Z(n26009) );
  XOR U26803 ( .A(n26011), .B(n26012), .Z(n15144) );
  XOR U26804 ( .A(n26013), .B(n26014), .Z(n26007) );
  AND U26805 ( .A(n26015), .B(n26016), .Z(n26014) );
  XOR U26806 ( .A(e_input[787]), .B(n26013), .Z(n26016) );
  XNOR U26807 ( .A(n15156), .B(n26013), .Z(n26015) );
  XOR U26808 ( .A(n26017), .B(n26018), .Z(n15156) );
  XOR U26809 ( .A(n26019), .B(n26020), .Z(n26013) );
  AND U26810 ( .A(n26021), .B(n26022), .Z(n26020) );
  XOR U26811 ( .A(e_input[786]), .B(n26019), .Z(n26022) );
  XNOR U26812 ( .A(n15168), .B(n26019), .Z(n26021) );
  XOR U26813 ( .A(n26023), .B(n26024), .Z(n15168) );
  XOR U26814 ( .A(n26025), .B(n26026), .Z(n26019) );
  AND U26815 ( .A(n26027), .B(n26028), .Z(n26026) );
  XOR U26816 ( .A(e_input[785]), .B(n26025), .Z(n26028) );
  XNOR U26817 ( .A(n15180), .B(n26025), .Z(n26027) );
  XOR U26818 ( .A(n26029), .B(n26030), .Z(n15180) );
  XOR U26819 ( .A(n26031), .B(n26032), .Z(n26025) );
  AND U26820 ( .A(n26033), .B(n26034), .Z(n26032) );
  XOR U26821 ( .A(e_input[784]), .B(n26031), .Z(n26034) );
  XNOR U26822 ( .A(n15192), .B(n26031), .Z(n26033) );
  XOR U26823 ( .A(n26035), .B(n26036), .Z(n15192) );
  XOR U26824 ( .A(n26037), .B(n26038), .Z(n26031) );
  AND U26825 ( .A(n26039), .B(n26040), .Z(n26038) );
  XOR U26826 ( .A(e_input[783]), .B(n26037), .Z(n26040) );
  XNOR U26827 ( .A(n15204), .B(n26037), .Z(n26039) );
  XOR U26828 ( .A(n26041), .B(n26042), .Z(n15204) );
  XOR U26829 ( .A(n26043), .B(n26044), .Z(n26037) );
  AND U26830 ( .A(n26045), .B(n26046), .Z(n26044) );
  XOR U26831 ( .A(e_input[782]), .B(n26043), .Z(n26046) );
  XNOR U26832 ( .A(n15216), .B(n26043), .Z(n26045) );
  XOR U26833 ( .A(n26047), .B(n26048), .Z(n15216) );
  XOR U26834 ( .A(n26049), .B(n26050), .Z(n26043) );
  AND U26835 ( .A(n26051), .B(n26052), .Z(n26050) );
  XOR U26836 ( .A(e_input[781]), .B(n26049), .Z(n26052) );
  XNOR U26837 ( .A(n15228), .B(n26049), .Z(n26051) );
  XOR U26838 ( .A(n26053), .B(n26054), .Z(n15228) );
  XOR U26839 ( .A(n26055), .B(n26056), .Z(n26049) );
  AND U26840 ( .A(n26057), .B(n26058), .Z(n26056) );
  XOR U26841 ( .A(e_input[780]), .B(n26055), .Z(n26058) );
  XNOR U26842 ( .A(n15240), .B(n26055), .Z(n26057) );
  XOR U26843 ( .A(n26059), .B(n26060), .Z(n15240) );
  XOR U26844 ( .A(n26061), .B(n26062), .Z(n26055) );
  AND U26845 ( .A(n26063), .B(n26064), .Z(n26062) );
  XOR U26846 ( .A(e_input[779]), .B(n26061), .Z(n26064) );
  XNOR U26847 ( .A(n15252), .B(n26061), .Z(n26063) );
  XOR U26848 ( .A(n26065), .B(n26066), .Z(n15252) );
  XOR U26849 ( .A(n26067), .B(n26068), .Z(n26061) );
  AND U26850 ( .A(n26069), .B(n26070), .Z(n26068) );
  XOR U26851 ( .A(e_input[778]), .B(n26067), .Z(n26070) );
  XNOR U26852 ( .A(n15264), .B(n26067), .Z(n26069) );
  XOR U26853 ( .A(n26071), .B(n26072), .Z(n15264) );
  XOR U26854 ( .A(n26073), .B(n26074), .Z(n26067) );
  AND U26855 ( .A(n26075), .B(n26076), .Z(n26074) );
  XOR U26856 ( .A(e_input[777]), .B(n26073), .Z(n26076) );
  XNOR U26857 ( .A(n15276), .B(n26073), .Z(n26075) );
  XOR U26858 ( .A(n26077), .B(n26078), .Z(n15276) );
  XOR U26859 ( .A(n26079), .B(n26080), .Z(n26073) );
  AND U26860 ( .A(n26081), .B(n26082), .Z(n26080) );
  XOR U26861 ( .A(e_input[776]), .B(n26079), .Z(n26082) );
  XNOR U26862 ( .A(n15288), .B(n26079), .Z(n26081) );
  XOR U26863 ( .A(n26083), .B(n26084), .Z(n15288) );
  XOR U26864 ( .A(n26085), .B(n26086), .Z(n26079) );
  AND U26865 ( .A(n26087), .B(n26088), .Z(n26086) );
  XOR U26866 ( .A(e_input[775]), .B(n26085), .Z(n26088) );
  XNOR U26867 ( .A(n15300), .B(n26085), .Z(n26087) );
  XOR U26868 ( .A(n26089), .B(n26090), .Z(n15300) );
  XOR U26869 ( .A(n26091), .B(n26092), .Z(n26085) );
  AND U26870 ( .A(n26093), .B(n26094), .Z(n26092) );
  XOR U26871 ( .A(e_input[774]), .B(n26091), .Z(n26094) );
  XNOR U26872 ( .A(n15312), .B(n26091), .Z(n26093) );
  XOR U26873 ( .A(n26095), .B(n26096), .Z(n15312) );
  XOR U26874 ( .A(n26097), .B(n26098), .Z(n26091) );
  AND U26875 ( .A(n26099), .B(n26100), .Z(n26098) );
  XOR U26876 ( .A(e_input[773]), .B(n26097), .Z(n26100) );
  XNOR U26877 ( .A(n15324), .B(n26097), .Z(n26099) );
  XOR U26878 ( .A(n26101), .B(n26102), .Z(n15324) );
  XOR U26879 ( .A(n26103), .B(n26104), .Z(n26097) );
  AND U26880 ( .A(n26105), .B(n26106), .Z(n26104) );
  XOR U26881 ( .A(e_input[772]), .B(n26103), .Z(n26106) );
  XNOR U26882 ( .A(n15336), .B(n26103), .Z(n26105) );
  XOR U26883 ( .A(n26107), .B(n26108), .Z(n15336) );
  XOR U26884 ( .A(n26109), .B(n26110), .Z(n26103) );
  AND U26885 ( .A(n26111), .B(n26112), .Z(n26110) );
  XOR U26886 ( .A(e_input[771]), .B(n26109), .Z(n26112) );
  XNOR U26887 ( .A(n15348), .B(n26109), .Z(n26111) );
  XOR U26888 ( .A(n26113), .B(n26114), .Z(n15348) );
  XOR U26889 ( .A(n26115), .B(n26116), .Z(n26109) );
  AND U26890 ( .A(n26117), .B(n26118), .Z(n26116) );
  XOR U26891 ( .A(e_input[770]), .B(n26115), .Z(n26118) );
  XNOR U26892 ( .A(n15360), .B(n26115), .Z(n26117) );
  XOR U26893 ( .A(n26119), .B(n26120), .Z(n15360) );
  XOR U26894 ( .A(n26121), .B(n26122), .Z(n26115) );
  AND U26895 ( .A(n26123), .B(n26124), .Z(n26122) );
  XOR U26896 ( .A(e_input[769]), .B(n26121), .Z(n26124) );
  XNOR U26897 ( .A(n15372), .B(n26121), .Z(n26123) );
  XOR U26898 ( .A(n26125), .B(n26126), .Z(n15372) );
  XOR U26899 ( .A(n26127), .B(n26128), .Z(n26121) );
  AND U26900 ( .A(n26129), .B(n26130), .Z(n26128) );
  XOR U26901 ( .A(e_input[768]), .B(n26127), .Z(n26130) );
  XNOR U26902 ( .A(n15384), .B(n26127), .Z(n26129) );
  XOR U26903 ( .A(n26131), .B(n26132), .Z(n15384) );
  XOR U26904 ( .A(n26133), .B(n26134), .Z(n26127) );
  AND U26905 ( .A(n26135), .B(n26136), .Z(n26134) );
  XOR U26906 ( .A(e_input[767]), .B(n26133), .Z(n26136) );
  XNOR U26907 ( .A(n15396), .B(n26133), .Z(n26135) );
  XOR U26908 ( .A(n26137), .B(n26138), .Z(n15396) );
  XOR U26909 ( .A(n26139), .B(n26140), .Z(n26133) );
  AND U26910 ( .A(n26141), .B(n26142), .Z(n26140) );
  XOR U26911 ( .A(e_input[766]), .B(n26139), .Z(n26142) );
  XNOR U26912 ( .A(n15408), .B(n26139), .Z(n26141) );
  XOR U26913 ( .A(n26143), .B(n26144), .Z(n15408) );
  XOR U26914 ( .A(n26145), .B(n26146), .Z(n26139) );
  AND U26915 ( .A(n26147), .B(n26148), .Z(n26146) );
  XOR U26916 ( .A(e_input[765]), .B(n26145), .Z(n26148) );
  XNOR U26917 ( .A(n15420), .B(n26145), .Z(n26147) );
  XOR U26918 ( .A(n26149), .B(n26150), .Z(n15420) );
  XOR U26919 ( .A(n26151), .B(n26152), .Z(n26145) );
  AND U26920 ( .A(n26153), .B(n26154), .Z(n26152) );
  XOR U26921 ( .A(e_input[764]), .B(n26151), .Z(n26154) );
  XNOR U26922 ( .A(n15432), .B(n26151), .Z(n26153) );
  XOR U26923 ( .A(n26155), .B(n26156), .Z(n15432) );
  XOR U26924 ( .A(n26157), .B(n26158), .Z(n26151) );
  AND U26925 ( .A(n26159), .B(n26160), .Z(n26158) );
  XOR U26926 ( .A(e_input[763]), .B(n26157), .Z(n26160) );
  XNOR U26927 ( .A(n15444), .B(n26157), .Z(n26159) );
  XOR U26928 ( .A(n26161), .B(n26162), .Z(n15444) );
  XOR U26929 ( .A(n26163), .B(n26164), .Z(n26157) );
  AND U26930 ( .A(n26165), .B(n26166), .Z(n26164) );
  XOR U26931 ( .A(e_input[762]), .B(n26163), .Z(n26166) );
  XNOR U26932 ( .A(n15456), .B(n26163), .Z(n26165) );
  XOR U26933 ( .A(n26167), .B(n26168), .Z(n15456) );
  XOR U26934 ( .A(n26169), .B(n26170), .Z(n26163) );
  AND U26935 ( .A(n26171), .B(n26172), .Z(n26170) );
  XOR U26936 ( .A(e_input[761]), .B(n26169), .Z(n26172) );
  XNOR U26937 ( .A(n15468), .B(n26169), .Z(n26171) );
  XOR U26938 ( .A(n26173), .B(n26174), .Z(n15468) );
  XOR U26939 ( .A(n26175), .B(n26176), .Z(n26169) );
  AND U26940 ( .A(n26177), .B(n26178), .Z(n26176) );
  XOR U26941 ( .A(e_input[760]), .B(n26175), .Z(n26178) );
  XNOR U26942 ( .A(n15480), .B(n26175), .Z(n26177) );
  XOR U26943 ( .A(n26179), .B(n26180), .Z(n15480) );
  XOR U26944 ( .A(n26181), .B(n26182), .Z(n26175) );
  AND U26945 ( .A(n26183), .B(n26184), .Z(n26182) );
  XOR U26946 ( .A(e_input[759]), .B(n26181), .Z(n26184) );
  XNOR U26947 ( .A(n15492), .B(n26181), .Z(n26183) );
  XOR U26948 ( .A(n26185), .B(n26186), .Z(n15492) );
  XOR U26949 ( .A(n26187), .B(n26188), .Z(n26181) );
  AND U26950 ( .A(n26189), .B(n26190), .Z(n26188) );
  XOR U26951 ( .A(e_input[758]), .B(n26187), .Z(n26190) );
  XNOR U26952 ( .A(n15504), .B(n26187), .Z(n26189) );
  XOR U26953 ( .A(n26191), .B(n26192), .Z(n15504) );
  XOR U26954 ( .A(n26193), .B(n26194), .Z(n26187) );
  AND U26955 ( .A(n26195), .B(n26196), .Z(n26194) );
  XOR U26956 ( .A(e_input[757]), .B(n26193), .Z(n26196) );
  XNOR U26957 ( .A(n15516), .B(n26193), .Z(n26195) );
  XOR U26958 ( .A(n26197), .B(n26198), .Z(n15516) );
  XOR U26959 ( .A(n26199), .B(n26200), .Z(n26193) );
  AND U26960 ( .A(n26201), .B(n26202), .Z(n26200) );
  XOR U26961 ( .A(e_input[756]), .B(n26199), .Z(n26202) );
  XNOR U26962 ( .A(n15528), .B(n26199), .Z(n26201) );
  XOR U26963 ( .A(n26203), .B(n26204), .Z(n15528) );
  XOR U26964 ( .A(n26205), .B(n26206), .Z(n26199) );
  AND U26965 ( .A(n26207), .B(n26208), .Z(n26206) );
  XOR U26966 ( .A(e_input[755]), .B(n26205), .Z(n26208) );
  XNOR U26967 ( .A(n15540), .B(n26205), .Z(n26207) );
  XOR U26968 ( .A(n26209), .B(n26210), .Z(n15540) );
  XOR U26969 ( .A(n26211), .B(n26212), .Z(n26205) );
  AND U26970 ( .A(n26213), .B(n26214), .Z(n26212) );
  XOR U26971 ( .A(e_input[754]), .B(n26211), .Z(n26214) );
  XNOR U26972 ( .A(n15552), .B(n26211), .Z(n26213) );
  XOR U26973 ( .A(n26215), .B(n26216), .Z(n15552) );
  XOR U26974 ( .A(n26217), .B(n26218), .Z(n26211) );
  AND U26975 ( .A(n26219), .B(n26220), .Z(n26218) );
  XOR U26976 ( .A(e_input[753]), .B(n26217), .Z(n26220) );
  XNOR U26977 ( .A(n15564), .B(n26217), .Z(n26219) );
  XOR U26978 ( .A(n26221), .B(n26222), .Z(n15564) );
  XOR U26979 ( .A(n26223), .B(n26224), .Z(n26217) );
  AND U26980 ( .A(n26225), .B(n26226), .Z(n26224) );
  XOR U26981 ( .A(e_input[752]), .B(n26223), .Z(n26226) );
  XNOR U26982 ( .A(n15576), .B(n26223), .Z(n26225) );
  XOR U26983 ( .A(n26227), .B(n26228), .Z(n15576) );
  XOR U26984 ( .A(n26229), .B(n26230), .Z(n26223) );
  AND U26985 ( .A(n26231), .B(n26232), .Z(n26230) );
  XOR U26986 ( .A(e_input[751]), .B(n26229), .Z(n26232) );
  XNOR U26987 ( .A(n15588), .B(n26229), .Z(n26231) );
  XOR U26988 ( .A(n26233), .B(n26234), .Z(n15588) );
  XOR U26989 ( .A(n26235), .B(n26236), .Z(n26229) );
  AND U26990 ( .A(n26237), .B(n26238), .Z(n26236) );
  XOR U26991 ( .A(e_input[750]), .B(n26235), .Z(n26238) );
  XNOR U26992 ( .A(n15600), .B(n26235), .Z(n26237) );
  XOR U26993 ( .A(n26239), .B(n26240), .Z(n15600) );
  XOR U26994 ( .A(n26241), .B(n26242), .Z(n26235) );
  AND U26995 ( .A(n26243), .B(n26244), .Z(n26242) );
  XOR U26996 ( .A(e_input[749]), .B(n26241), .Z(n26244) );
  XNOR U26997 ( .A(n15612), .B(n26241), .Z(n26243) );
  XOR U26998 ( .A(n26245), .B(n26246), .Z(n15612) );
  XOR U26999 ( .A(n26247), .B(n26248), .Z(n26241) );
  AND U27000 ( .A(n26249), .B(n26250), .Z(n26248) );
  XOR U27001 ( .A(e_input[748]), .B(n26247), .Z(n26250) );
  XNOR U27002 ( .A(n15624), .B(n26247), .Z(n26249) );
  XOR U27003 ( .A(n26251), .B(n26252), .Z(n15624) );
  XOR U27004 ( .A(n26253), .B(n26254), .Z(n26247) );
  AND U27005 ( .A(n26255), .B(n26256), .Z(n26254) );
  XOR U27006 ( .A(e_input[747]), .B(n26253), .Z(n26256) );
  XNOR U27007 ( .A(n15636), .B(n26253), .Z(n26255) );
  XOR U27008 ( .A(n26257), .B(n26258), .Z(n15636) );
  XOR U27009 ( .A(n26259), .B(n26260), .Z(n26253) );
  AND U27010 ( .A(n26261), .B(n26262), .Z(n26260) );
  XOR U27011 ( .A(e_input[746]), .B(n26259), .Z(n26262) );
  XNOR U27012 ( .A(n15648), .B(n26259), .Z(n26261) );
  XOR U27013 ( .A(n26263), .B(n26264), .Z(n15648) );
  XOR U27014 ( .A(n26265), .B(n26266), .Z(n26259) );
  AND U27015 ( .A(n26267), .B(n26268), .Z(n26266) );
  XOR U27016 ( .A(e_input[745]), .B(n26265), .Z(n26268) );
  XNOR U27017 ( .A(n15660), .B(n26265), .Z(n26267) );
  XOR U27018 ( .A(n26269), .B(n26270), .Z(n15660) );
  XOR U27019 ( .A(n26271), .B(n26272), .Z(n26265) );
  AND U27020 ( .A(n26273), .B(n26274), .Z(n26272) );
  XOR U27021 ( .A(e_input[744]), .B(n26271), .Z(n26274) );
  XNOR U27022 ( .A(n15672), .B(n26271), .Z(n26273) );
  XOR U27023 ( .A(n26275), .B(n26276), .Z(n15672) );
  XOR U27024 ( .A(n26277), .B(n26278), .Z(n26271) );
  AND U27025 ( .A(n26279), .B(n26280), .Z(n26278) );
  XOR U27026 ( .A(e_input[743]), .B(n26277), .Z(n26280) );
  XNOR U27027 ( .A(n15684), .B(n26277), .Z(n26279) );
  XOR U27028 ( .A(n26281), .B(n26282), .Z(n15684) );
  XOR U27029 ( .A(n26283), .B(n26284), .Z(n26277) );
  AND U27030 ( .A(n26285), .B(n26286), .Z(n26284) );
  XOR U27031 ( .A(e_input[742]), .B(n26283), .Z(n26286) );
  XNOR U27032 ( .A(n15696), .B(n26283), .Z(n26285) );
  XOR U27033 ( .A(n26287), .B(n26288), .Z(n15696) );
  XOR U27034 ( .A(n26289), .B(n26290), .Z(n26283) );
  AND U27035 ( .A(n26291), .B(n26292), .Z(n26290) );
  XOR U27036 ( .A(e_input[741]), .B(n26289), .Z(n26292) );
  XNOR U27037 ( .A(n15708), .B(n26289), .Z(n26291) );
  XOR U27038 ( .A(n26293), .B(n26294), .Z(n15708) );
  XOR U27039 ( .A(n26295), .B(n26296), .Z(n26289) );
  AND U27040 ( .A(n26297), .B(n26298), .Z(n26296) );
  XOR U27041 ( .A(e_input[740]), .B(n26295), .Z(n26298) );
  XNOR U27042 ( .A(n15720), .B(n26295), .Z(n26297) );
  XOR U27043 ( .A(n26299), .B(n26300), .Z(n15720) );
  XOR U27044 ( .A(n26301), .B(n26302), .Z(n26295) );
  AND U27045 ( .A(n26303), .B(n26304), .Z(n26302) );
  XOR U27046 ( .A(e_input[739]), .B(n26301), .Z(n26304) );
  XNOR U27047 ( .A(n15732), .B(n26301), .Z(n26303) );
  XOR U27048 ( .A(n26305), .B(n26306), .Z(n15732) );
  XOR U27049 ( .A(n26307), .B(n26308), .Z(n26301) );
  AND U27050 ( .A(n26309), .B(n26310), .Z(n26308) );
  XOR U27051 ( .A(e_input[738]), .B(n26307), .Z(n26310) );
  XNOR U27052 ( .A(n15744), .B(n26307), .Z(n26309) );
  XOR U27053 ( .A(n26311), .B(n26312), .Z(n15744) );
  XOR U27054 ( .A(n26313), .B(n26314), .Z(n26307) );
  AND U27055 ( .A(n26315), .B(n26316), .Z(n26314) );
  XOR U27056 ( .A(e_input[737]), .B(n26313), .Z(n26316) );
  XNOR U27057 ( .A(n15756), .B(n26313), .Z(n26315) );
  XOR U27058 ( .A(n26317), .B(n26318), .Z(n15756) );
  XOR U27059 ( .A(n26319), .B(n26320), .Z(n26313) );
  AND U27060 ( .A(n26321), .B(n26322), .Z(n26320) );
  XOR U27061 ( .A(e_input[736]), .B(n26319), .Z(n26322) );
  XNOR U27062 ( .A(n15768), .B(n26319), .Z(n26321) );
  XOR U27063 ( .A(n26323), .B(n26324), .Z(n15768) );
  XOR U27064 ( .A(n26325), .B(n26326), .Z(n26319) );
  AND U27065 ( .A(n26327), .B(n26328), .Z(n26326) );
  XOR U27066 ( .A(e_input[735]), .B(n26325), .Z(n26328) );
  XNOR U27067 ( .A(n15780), .B(n26325), .Z(n26327) );
  XOR U27068 ( .A(n26329), .B(n26330), .Z(n15780) );
  XOR U27069 ( .A(n26331), .B(n26332), .Z(n26325) );
  AND U27070 ( .A(n26333), .B(n26334), .Z(n26332) );
  XOR U27071 ( .A(e_input[734]), .B(n26331), .Z(n26334) );
  XNOR U27072 ( .A(n15792), .B(n26331), .Z(n26333) );
  XOR U27073 ( .A(n26335), .B(n26336), .Z(n15792) );
  XOR U27074 ( .A(n26337), .B(n26338), .Z(n26331) );
  AND U27075 ( .A(n26339), .B(n26340), .Z(n26338) );
  XOR U27076 ( .A(e_input[733]), .B(n26337), .Z(n26340) );
  XNOR U27077 ( .A(n15804), .B(n26337), .Z(n26339) );
  XOR U27078 ( .A(n26341), .B(n26342), .Z(n15804) );
  XOR U27079 ( .A(n26343), .B(n26344), .Z(n26337) );
  AND U27080 ( .A(n26345), .B(n26346), .Z(n26344) );
  XOR U27081 ( .A(e_input[732]), .B(n26343), .Z(n26346) );
  XNOR U27082 ( .A(n15816), .B(n26343), .Z(n26345) );
  XOR U27083 ( .A(n26347), .B(n26348), .Z(n15816) );
  XOR U27084 ( .A(n26349), .B(n26350), .Z(n26343) );
  AND U27085 ( .A(n26351), .B(n26352), .Z(n26350) );
  XOR U27086 ( .A(e_input[731]), .B(n26349), .Z(n26352) );
  XNOR U27087 ( .A(n15828), .B(n26349), .Z(n26351) );
  XOR U27088 ( .A(n26353), .B(n26354), .Z(n15828) );
  XOR U27089 ( .A(n26355), .B(n26356), .Z(n26349) );
  AND U27090 ( .A(n26357), .B(n26358), .Z(n26356) );
  XOR U27091 ( .A(e_input[730]), .B(n26355), .Z(n26358) );
  XNOR U27092 ( .A(n15840), .B(n26355), .Z(n26357) );
  XOR U27093 ( .A(n26359), .B(n26360), .Z(n15840) );
  XOR U27094 ( .A(n26361), .B(n26362), .Z(n26355) );
  AND U27095 ( .A(n26363), .B(n26364), .Z(n26362) );
  XOR U27096 ( .A(e_input[729]), .B(n26361), .Z(n26364) );
  XNOR U27097 ( .A(n15852), .B(n26361), .Z(n26363) );
  XOR U27098 ( .A(n26365), .B(n26366), .Z(n15852) );
  XOR U27099 ( .A(n26367), .B(n26368), .Z(n26361) );
  AND U27100 ( .A(n26369), .B(n26370), .Z(n26368) );
  XOR U27101 ( .A(e_input[728]), .B(n26367), .Z(n26370) );
  XNOR U27102 ( .A(n15864), .B(n26367), .Z(n26369) );
  XOR U27103 ( .A(n26371), .B(n26372), .Z(n15864) );
  XOR U27104 ( .A(n26373), .B(n26374), .Z(n26367) );
  AND U27105 ( .A(n26375), .B(n26376), .Z(n26374) );
  XOR U27106 ( .A(e_input[727]), .B(n26373), .Z(n26376) );
  XNOR U27107 ( .A(n15876), .B(n26373), .Z(n26375) );
  XOR U27108 ( .A(n26377), .B(n26378), .Z(n15876) );
  XOR U27109 ( .A(n26379), .B(n26380), .Z(n26373) );
  AND U27110 ( .A(n26381), .B(n26382), .Z(n26380) );
  XOR U27111 ( .A(e_input[726]), .B(n26379), .Z(n26382) );
  XNOR U27112 ( .A(n15888), .B(n26379), .Z(n26381) );
  XOR U27113 ( .A(n26383), .B(n26384), .Z(n15888) );
  XOR U27114 ( .A(n26385), .B(n26386), .Z(n26379) );
  AND U27115 ( .A(n26387), .B(n26388), .Z(n26386) );
  XOR U27116 ( .A(e_input[725]), .B(n26385), .Z(n26388) );
  XNOR U27117 ( .A(n15900), .B(n26385), .Z(n26387) );
  XOR U27118 ( .A(n26389), .B(n26390), .Z(n15900) );
  XOR U27119 ( .A(n26391), .B(n26392), .Z(n26385) );
  AND U27120 ( .A(n26393), .B(n26394), .Z(n26392) );
  XOR U27121 ( .A(e_input[724]), .B(n26391), .Z(n26394) );
  XNOR U27122 ( .A(n15912), .B(n26391), .Z(n26393) );
  XOR U27123 ( .A(n26395), .B(n26396), .Z(n15912) );
  XOR U27124 ( .A(n26397), .B(n26398), .Z(n26391) );
  AND U27125 ( .A(n26399), .B(n26400), .Z(n26398) );
  XOR U27126 ( .A(e_input[723]), .B(n26397), .Z(n26400) );
  XNOR U27127 ( .A(n15924), .B(n26397), .Z(n26399) );
  XOR U27128 ( .A(n26401), .B(n26402), .Z(n15924) );
  XOR U27129 ( .A(n26403), .B(n26404), .Z(n26397) );
  AND U27130 ( .A(n26405), .B(n26406), .Z(n26404) );
  XOR U27131 ( .A(e_input[722]), .B(n26403), .Z(n26406) );
  XNOR U27132 ( .A(n15936), .B(n26403), .Z(n26405) );
  XOR U27133 ( .A(n26407), .B(n26408), .Z(n15936) );
  XOR U27134 ( .A(n26409), .B(n26410), .Z(n26403) );
  AND U27135 ( .A(n26411), .B(n26412), .Z(n26410) );
  XOR U27136 ( .A(e_input[721]), .B(n26409), .Z(n26412) );
  XNOR U27137 ( .A(n15948), .B(n26409), .Z(n26411) );
  XOR U27138 ( .A(n26413), .B(n26414), .Z(n15948) );
  XOR U27139 ( .A(n26415), .B(n26416), .Z(n26409) );
  AND U27140 ( .A(n26417), .B(n26418), .Z(n26416) );
  XOR U27141 ( .A(e_input[720]), .B(n26415), .Z(n26418) );
  XNOR U27142 ( .A(n15960), .B(n26415), .Z(n26417) );
  XOR U27143 ( .A(n26419), .B(n26420), .Z(n15960) );
  XOR U27144 ( .A(n26421), .B(n26422), .Z(n26415) );
  AND U27145 ( .A(n26423), .B(n26424), .Z(n26422) );
  XOR U27146 ( .A(e_input[719]), .B(n26421), .Z(n26424) );
  XNOR U27147 ( .A(n15972), .B(n26421), .Z(n26423) );
  XOR U27148 ( .A(n26425), .B(n26426), .Z(n15972) );
  XOR U27149 ( .A(n26427), .B(n26428), .Z(n26421) );
  AND U27150 ( .A(n26429), .B(n26430), .Z(n26428) );
  XOR U27151 ( .A(e_input[718]), .B(n26427), .Z(n26430) );
  XNOR U27152 ( .A(n15984), .B(n26427), .Z(n26429) );
  XOR U27153 ( .A(n26431), .B(n26432), .Z(n15984) );
  XOR U27154 ( .A(n26433), .B(n26434), .Z(n26427) );
  AND U27155 ( .A(n26435), .B(n26436), .Z(n26434) );
  XOR U27156 ( .A(e_input[717]), .B(n26433), .Z(n26436) );
  XNOR U27157 ( .A(n15996), .B(n26433), .Z(n26435) );
  XOR U27158 ( .A(n26437), .B(n26438), .Z(n15996) );
  XOR U27159 ( .A(n26439), .B(n26440), .Z(n26433) );
  AND U27160 ( .A(n26441), .B(n26442), .Z(n26440) );
  XOR U27161 ( .A(e_input[716]), .B(n26439), .Z(n26442) );
  XNOR U27162 ( .A(n16008), .B(n26439), .Z(n26441) );
  XOR U27163 ( .A(n26443), .B(n26444), .Z(n16008) );
  XOR U27164 ( .A(n26445), .B(n26446), .Z(n26439) );
  AND U27165 ( .A(n26447), .B(n26448), .Z(n26446) );
  XOR U27166 ( .A(e_input[715]), .B(n26445), .Z(n26448) );
  XNOR U27167 ( .A(n16020), .B(n26445), .Z(n26447) );
  XOR U27168 ( .A(n26449), .B(n26450), .Z(n16020) );
  XOR U27169 ( .A(n26451), .B(n26452), .Z(n26445) );
  AND U27170 ( .A(n26453), .B(n26454), .Z(n26452) );
  XOR U27171 ( .A(e_input[714]), .B(n26451), .Z(n26454) );
  XNOR U27172 ( .A(n16032), .B(n26451), .Z(n26453) );
  XOR U27173 ( .A(n26455), .B(n26456), .Z(n16032) );
  XOR U27174 ( .A(n26457), .B(n26458), .Z(n26451) );
  AND U27175 ( .A(n26459), .B(n26460), .Z(n26458) );
  XOR U27176 ( .A(e_input[713]), .B(n26457), .Z(n26460) );
  XNOR U27177 ( .A(n16044), .B(n26457), .Z(n26459) );
  XOR U27178 ( .A(n26461), .B(n26462), .Z(n16044) );
  XOR U27179 ( .A(n26463), .B(n26464), .Z(n26457) );
  AND U27180 ( .A(n26465), .B(n26466), .Z(n26464) );
  XOR U27181 ( .A(e_input[712]), .B(n26463), .Z(n26466) );
  XNOR U27182 ( .A(n16056), .B(n26463), .Z(n26465) );
  XOR U27183 ( .A(n26467), .B(n26468), .Z(n16056) );
  XOR U27184 ( .A(n26469), .B(n26470), .Z(n26463) );
  AND U27185 ( .A(n26471), .B(n26472), .Z(n26470) );
  XOR U27186 ( .A(e_input[711]), .B(n26469), .Z(n26472) );
  XNOR U27187 ( .A(n16068), .B(n26469), .Z(n26471) );
  XOR U27188 ( .A(n26473), .B(n26474), .Z(n16068) );
  XOR U27189 ( .A(n26475), .B(n26476), .Z(n26469) );
  AND U27190 ( .A(n26477), .B(n26478), .Z(n26476) );
  XOR U27191 ( .A(e_input[710]), .B(n26475), .Z(n26478) );
  XNOR U27192 ( .A(n16080), .B(n26475), .Z(n26477) );
  XOR U27193 ( .A(n26479), .B(n26480), .Z(n16080) );
  XOR U27194 ( .A(n26481), .B(n26482), .Z(n26475) );
  AND U27195 ( .A(n26483), .B(n26484), .Z(n26482) );
  XOR U27196 ( .A(e_input[709]), .B(n26481), .Z(n26484) );
  XNOR U27197 ( .A(n16092), .B(n26481), .Z(n26483) );
  XOR U27198 ( .A(n26485), .B(n26486), .Z(n16092) );
  XOR U27199 ( .A(n26487), .B(n26488), .Z(n26481) );
  AND U27200 ( .A(n26489), .B(n26490), .Z(n26488) );
  XOR U27201 ( .A(e_input[708]), .B(n26487), .Z(n26490) );
  XNOR U27202 ( .A(n16104), .B(n26487), .Z(n26489) );
  XOR U27203 ( .A(n26491), .B(n26492), .Z(n16104) );
  XOR U27204 ( .A(n26493), .B(n26494), .Z(n26487) );
  AND U27205 ( .A(n26495), .B(n26496), .Z(n26494) );
  XOR U27206 ( .A(e_input[707]), .B(n26493), .Z(n26496) );
  XNOR U27207 ( .A(n16116), .B(n26493), .Z(n26495) );
  XOR U27208 ( .A(n26497), .B(n26498), .Z(n16116) );
  XOR U27209 ( .A(n26499), .B(n26500), .Z(n26493) );
  AND U27210 ( .A(n26501), .B(n26502), .Z(n26500) );
  XOR U27211 ( .A(e_input[706]), .B(n26499), .Z(n26502) );
  XNOR U27212 ( .A(n16128), .B(n26499), .Z(n26501) );
  XOR U27213 ( .A(n26503), .B(n26504), .Z(n16128) );
  XOR U27214 ( .A(n26505), .B(n26506), .Z(n26499) );
  AND U27215 ( .A(n26507), .B(n26508), .Z(n26506) );
  XOR U27216 ( .A(e_input[705]), .B(n26505), .Z(n26508) );
  XNOR U27217 ( .A(n16140), .B(n26505), .Z(n26507) );
  XOR U27218 ( .A(n26509), .B(n26510), .Z(n16140) );
  XOR U27219 ( .A(n26511), .B(n26512), .Z(n26505) );
  AND U27220 ( .A(n26513), .B(n26514), .Z(n26512) );
  XOR U27221 ( .A(e_input[704]), .B(n26511), .Z(n26514) );
  XNOR U27222 ( .A(n16152), .B(n26511), .Z(n26513) );
  XOR U27223 ( .A(n26515), .B(n26516), .Z(n16152) );
  XOR U27224 ( .A(n26517), .B(n26518), .Z(n26511) );
  AND U27225 ( .A(n26519), .B(n26520), .Z(n26518) );
  XOR U27226 ( .A(e_input[703]), .B(n26517), .Z(n26520) );
  XNOR U27227 ( .A(n16164), .B(n26517), .Z(n26519) );
  XOR U27228 ( .A(n26521), .B(n26522), .Z(n16164) );
  XOR U27229 ( .A(n26523), .B(n26524), .Z(n26517) );
  AND U27230 ( .A(n26525), .B(n26526), .Z(n26524) );
  XOR U27231 ( .A(e_input[702]), .B(n26523), .Z(n26526) );
  XNOR U27232 ( .A(n16176), .B(n26523), .Z(n26525) );
  XOR U27233 ( .A(n26527), .B(n26528), .Z(n16176) );
  XOR U27234 ( .A(n26529), .B(n26530), .Z(n26523) );
  AND U27235 ( .A(n26531), .B(n26532), .Z(n26530) );
  XOR U27236 ( .A(e_input[701]), .B(n26529), .Z(n26532) );
  XNOR U27237 ( .A(n16188), .B(n26529), .Z(n26531) );
  XOR U27238 ( .A(n26533), .B(n26534), .Z(n16188) );
  XOR U27239 ( .A(n26535), .B(n26536), .Z(n26529) );
  AND U27240 ( .A(n26537), .B(n26538), .Z(n26536) );
  XOR U27241 ( .A(e_input[700]), .B(n26535), .Z(n26538) );
  XNOR U27242 ( .A(n16200), .B(n26535), .Z(n26537) );
  XOR U27243 ( .A(n26539), .B(n26540), .Z(n16200) );
  XOR U27244 ( .A(n26541), .B(n26542), .Z(n26535) );
  AND U27245 ( .A(n26543), .B(n26544), .Z(n26542) );
  XOR U27246 ( .A(e_input[699]), .B(n26541), .Z(n26544) );
  XNOR U27247 ( .A(n16212), .B(n26541), .Z(n26543) );
  XOR U27248 ( .A(n26545), .B(n26546), .Z(n16212) );
  XOR U27249 ( .A(n26547), .B(n26548), .Z(n26541) );
  AND U27250 ( .A(n26549), .B(n26550), .Z(n26548) );
  XOR U27251 ( .A(e_input[698]), .B(n26547), .Z(n26550) );
  XNOR U27252 ( .A(n16224), .B(n26547), .Z(n26549) );
  XOR U27253 ( .A(n26551), .B(n26552), .Z(n16224) );
  XOR U27254 ( .A(n26553), .B(n26554), .Z(n26547) );
  AND U27255 ( .A(n26555), .B(n26556), .Z(n26554) );
  XOR U27256 ( .A(e_input[697]), .B(n26553), .Z(n26556) );
  XNOR U27257 ( .A(n16236), .B(n26553), .Z(n26555) );
  XOR U27258 ( .A(n26557), .B(n26558), .Z(n16236) );
  XOR U27259 ( .A(n26559), .B(n26560), .Z(n26553) );
  AND U27260 ( .A(n26561), .B(n26562), .Z(n26560) );
  XOR U27261 ( .A(e_input[696]), .B(n26559), .Z(n26562) );
  XNOR U27262 ( .A(n16248), .B(n26559), .Z(n26561) );
  XOR U27263 ( .A(n26563), .B(n26564), .Z(n16248) );
  XOR U27264 ( .A(n26565), .B(n26566), .Z(n26559) );
  AND U27265 ( .A(n26567), .B(n26568), .Z(n26566) );
  XOR U27266 ( .A(e_input[695]), .B(n26565), .Z(n26568) );
  XNOR U27267 ( .A(n16260), .B(n26565), .Z(n26567) );
  XOR U27268 ( .A(n26569), .B(n26570), .Z(n16260) );
  XOR U27269 ( .A(n26571), .B(n26572), .Z(n26565) );
  AND U27270 ( .A(n26573), .B(n26574), .Z(n26572) );
  XOR U27271 ( .A(e_input[694]), .B(n26571), .Z(n26574) );
  XNOR U27272 ( .A(n16272), .B(n26571), .Z(n26573) );
  XOR U27273 ( .A(n26575), .B(n26576), .Z(n16272) );
  XOR U27274 ( .A(n26577), .B(n26578), .Z(n26571) );
  AND U27275 ( .A(n26579), .B(n26580), .Z(n26578) );
  XOR U27276 ( .A(e_input[693]), .B(n26577), .Z(n26580) );
  XNOR U27277 ( .A(n16284), .B(n26577), .Z(n26579) );
  XOR U27278 ( .A(n26581), .B(n26582), .Z(n16284) );
  XOR U27279 ( .A(n26583), .B(n26584), .Z(n26577) );
  AND U27280 ( .A(n26585), .B(n26586), .Z(n26584) );
  XOR U27281 ( .A(e_input[692]), .B(n26583), .Z(n26586) );
  XNOR U27282 ( .A(n16296), .B(n26583), .Z(n26585) );
  XOR U27283 ( .A(n26587), .B(n26588), .Z(n16296) );
  XOR U27284 ( .A(n26589), .B(n26590), .Z(n26583) );
  AND U27285 ( .A(n26591), .B(n26592), .Z(n26590) );
  XOR U27286 ( .A(e_input[691]), .B(n26589), .Z(n26592) );
  XNOR U27287 ( .A(n16308), .B(n26589), .Z(n26591) );
  XOR U27288 ( .A(n26593), .B(n26594), .Z(n16308) );
  XOR U27289 ( .A(n26595), .B(n26596), .Z(n26589) );
  AND U27290 ( .A(n26597), .B(n26598), .Z(n26596) );
  XOR U27291 ( .A(e_input[690]), .B(n26595), .Z(n26598) );
  XNOR U27292 ( .A(n16320), .B(n26595), .Z(n26597) );
  XOR U27293 ( .A(n26599), .B(n26600), .Z(n16320) );
  XOR U27294 ( .A(n26601), .B(n26602), .Z(n26595) );
  AND U27295 ( .A(n26603), .B(n26604), .Z(n26602) );
  XOR U27296 ( .A(e_input[689]), .B(n26601), .Z(n26604) );
  XNOR U27297 ( .A(n16332), .B(n26601), .Z(n26603) );
  XOR U27298 ( .A(n26605), .B(n26606), .Z(n16332) );
  XOR U27299 ( .A(n26607), .B(n26608), .Z(n26601) );
  AND U27300 ( .A(n26609), .B(n26610), .Z(n26608) );
  XOR U27301 ( .A(e_input[688]), .B(n26607), .Z(n26610) );
  XNOR U27302 ( .A(n16344), .B(n26607), .Z(n26609) );
  XOR U27303 ( .A(n26611), .B(n26612), .Z(n16344) );
  XOR U27304 ( .A(n26613), .B(n26614), .Z(n26607) );
  AND U27305 ( .A(n26615), .B(n26616), .Z(n26614) );
  XOR U27306 ( .A(e_input[687]), .B(n26613), .Z(n26616) );
  XNOR U27307 ( .A(n16356), .B(n26613), .Z(n26615) );
  XOR U27308 ( .A(n26617), .B(n26618), .Z(n16356) );
  XOR U27309 ( .A(n26619), .B(n26620), .Z(n26613) );
  AND U27310 ( .A(n26621), .B(n26622), .Z(n26620) );
  XOR U27311 ( .A(e_input[686]), .B(n26619), .Z(n26622) );
  XNOR U27312 ( .A(n16368), .B(n26619), .Z(n26621) );
  XOR U27313 ( .A(n26623), .B(n26624), .Z(n16368) );
  XOR U27314 ( .A(n26625), .B(n26626), .Z(n26619) );
  AND U27315 ( .A(n26627), .B(n26628), .Z(n26626) );
  XOR U27316 ( .A(e_input[685]), .B(n26625), .Z(n26628) );
  XNOR U27317 ( .A(n16380), .B(n26625), .Z(n26627) );
  XOR U27318 ( .A(n26629), .B(n26630), .Z(n16380) );
  XOR U27319 ( .A(n26631), .B(n26632), .Z(n26625) );
  AND U27320 ( .A(n26633), .B(n26634), .Z(n26632) );
  XOR U27321 ( .A(e_input[684]), .B(n26631), .Z(n26634) );
  XNOR U27322 ( .A(n16392), .B(n26631), .Z(n26633) );
  XOR U27323 ( .A(n26635), .B(n26636), .Z(n16392) );
  XOR U27324 ( .A(n26637), .B(n26638), .Z(n26631) );
  AND U27325 ( .A(n26639), .B(n26640), .Z(n26638) );
  XOR U27326 ( .A(e_input[683]), .B(n26637), .Z(n26640) );
  XNOR U27327 ( .A(n16404), .B(n26637), .Z(n26639) );
  XOR U27328 ( .A(n26641), .B(n26642), .Z(n16404) );
  XOR U27329 ( .A(n26643), .B(n26644), .Z(n26637) );
  AND U27330 ( .A(n26645), .B(n26646), .Z(n26644) );
  XOR U27331 ( .A(e_input[682]), .B(n26643), .Z(n26646) );
  XNOR U27332 ( .A(n16416), .B(n26643), .Z(n26645) );
  XOR U27333 ( .A(n26647), .B(n26648), .Z(n16416) );
  XOR U27334 ( .A(n26649), .B(n26650), .Z(n26643) );
  AND U27335 ( .A(n26651), .B(n26652), .Z(n26650) );
  XOR U27336 ( .A(e_input[681]), .B(n26649), .Z(n26652) );
  XNOR U27337 ( .A(n16428), .B(n26649), .Z(n26651) );
  XOR U27338 ( .A(n26653), .B(n26654), .Z(n16428) );
  XOR U27339 ( .A(n26655), .B(n26656), .Z(n26649) );
  AND U27340 ( .A(n26657), .B(n26658), .Z(n26656) );
  XOR U27341 ( .A(e_input[680]), .B(n26655), .Z(n26658) );
  XNOR U27342 ( .A(n16440), .B(n26655), .Z(n26657) );
  XOR U27343 ( .A(n26659), .B(n26660), .Z(n16440) );
  XOR U27344 ( .A(n26661), .B(n26662), .Z(n26655) );
  AND U27345 ( .A(n26663), .B(n26664), .Z(n26662) );
  XOR U27346 ( .A(e_input[679]), .B(n26661), .Z(n26664) );
  XNOR U27347 ( .A(n16452), .B(n26661), .Z(n26663) );
  XOR U27348 ( .A(n26665), .B(n26666), .Z(n16452) );
  XOR U27349 ( .A(n26667), .B(n26668), .Z(n26661) );
  AND U27350 ( .A(n26669), .B(n26670), .Z(n26668) );
  XOR U27351 ( .A(e_input[678]), .B(n26667), .Z(n26670) );
  XNOR U27352 ( .A(n16464), .B(n26667), .Z(n26669) );
  XOR U27353 ( .A(n26671), .B(n26672), .Z(n16464) );
  XOR U27354 ( .A(n26673), .B(n26674), .Z(n26667) );
  AND U27355 ( .A(n26675), .B(n26676), .Z(n26674) );
  XOR U27356 ( .A(e_input[677]), .B(n26673), .Z(n26676) );
  XNOR U27357 ( .A(n16476), .B(n26673), .Z(n26675) );
  XOR U27358 ( .A(n26677), .B(n26678), .Z(n16476) );
  XOR U27359 ( .A(n26679), .B(n26680), .Z(n26673) );
  AND U27360 ( .A(n26681), .B(n26682), .Z(n26680) );
  XOR U27361 ( .A(e_input[676]), .B(n26679), .Z(n26682) );
  XNOR U27362 ( .A(n16488), .B(n26679), .Z(n26681) );
  XOR U27363 ( .A(n26683), .B(n26684), .Z(n16488) );
  XOR U27364 ( .A(n26685), .B(n26686), .Z(n26679) );
  AND U27365 ( .A(n26687), .B(n26688), .Z(n26686) );
  XOR U27366 ( .A(e_input[675]), .B(n26685), .Z(n26688) );
  XNOR U27367 ( .A(n16500), .B(n26685), .Z(n26687) );
  XOR U27368 ( .A(n26689), .B(n26690), .Z(n16500) );
  XOR U27369 ( .A(n26691), .B(n26692), .Z(n26685) );
  AND U27370 ( .A(n26693), .B(n26694), .Z(n26692) );
  XOR U27371 ( .A(e_input[674]), .B(n26691), .Z(n26694) );
  XNOR U27372 ( .A(n16512), .B(n26691), .Z(n26693) );
  XOR U27373 ( .A(n26695), .B(n26696), .Z(n16512) );
  XOR U27374 ( .A(n26697), .B(n26698), .Z(n26691) );
  AND U27375 ( .A(n26699), .B(n26700), .Z(n26698) );
  XOR U27376 ( .A(e_input[673]), .B(n26697), .Z(n26700) );
  XNOR U27377 ( .A(n16524), .B(n26697), .Z(n26699) );
  XOR U27378 ( .A(n26701), .B(n26702), .Z(n16524) );
  XOR U27379 ( .A(n26703), .B(n26704), .Z(n26697) );
  AND U27380 ( .A(n26705), .B(n26706), .Z(n26704) );
  XOR U27381 ( .A(e_input[672]), .B(n26703), .Z(n26706) );
  XNOR U27382 ( .A(n16536), .B(n26703), .Z(n26705) );
  XOR U27383 ( .A(n26707), .B(n26708), .Z(n16536) );
  XOR U27384 ( .A(n26709), .B(n26710), .Z(n26703) );
  AND U27385 ( .A(n26711), .B(n26712), .Z(n26710) );
  XOR U27386 ( .A(e_input[671]), .B(n26709), .Z(n26712) );
  XNOR U27387 ( .A(n16548), .B(n26709), .Z(n26711) );
  XOR U27388 ( .A(n26713), .B(n26714), .Z(n16548) );
  XOR U27389 ( .A(n26715), .B(n26716), .Z(n26709) );
  AND U27390 ( .A(n26717), .B(n26718), .Z(n26716) );
  XOR U27391 ( .A(e_input[670]), .B(n26715), .Z(n26718) );
  XNOR U27392 ( .A(n16560), .B(n26715), .Z(n26717) );
  XOR U27393 ( .A(n26719), .B(n26720), .Z(n16560) );
  XOR U27394 ( .A(n26721), .B(n26722), .Z(n26715) );
  AND U27395 ( .A(n26723), .B(n26724), .Z(n26722) );
  XOR U27396 ( .A(e_input[669]), .B(n26721), .Z(n26724) );
  XNOR U27397 ( .A(n16572), .B(n26721), .Z(n26723) );
  XOR U27398 ( .A(n26725), .B(n26726), .Z(n16572) );
  XOR U27399 ( .A(n26727), .B(n26728), .Z(n26721) );
  AND U27400 ( .A(n26729), .B(n26730), .Z(n26728) );
  XOR U27401 ( .A(e_input[668]), .B(n26727), .Z(n26730) );
  XNOR U27402 ( .A(n16584), .B(n26727), .Z(n26729) );
  XOR U27403 ( .A(n26731), .B(n26732), .Z(n16584) );
  XOR U27404 ( .A(n26733), .B(n26734), .Z(n26727) );
  AND U27405 ( .A(n26735), .B(n26736), .Z(n26734) );
  XOR U27406 ( .A(e_input[667]), .B(n26733), .Z(n26736) );
  XNOR U27407 ( .A(n16596), .B(n26733), .Z(n26735) );
  XOR U27408 ( .A(n26737), .B(n26738), .Z(n16596) );
  XOR U27409 ( .A(n26739), .B(n26740), .Z(n26733) );
  AND U27410 ( .A(n26741), .B(n26742), .Z(n26740) );
  XOR U27411 ( .A(e_input[666]), .B(n26739), .Z(n26742) );
  XNOR U27412 ( .A(n16608), .B(n26739), .Z(n26741) );
  XOR U27413 ( .A(n26743), .B(n26744), .Z(n16608) );
  XOR U27414 ( .A(n26745), .B(n26746), .Z(n26739) );
  AND U27415 ( .A(n26747), .B(n26748), .Z(n26746) );
  XOR U27416 ( .A(e_input[665]), .B(n26745), .Z(n26748) );
  XNOR U27417 ( .A(n16620), .B(n26745), .Z(n26747) );
  XOR U27418 ( .A(n26749), .B(n26750), .Z(n16620) );
  XOR U27419 ( .A(n26751), .B(n26752), .Z(n26745) );
  AND U27420 ( .A(n26753), .B(n26754), .Z(n26752) );
  XOR U27421 ( .A(e_input[664]), .B(n26751), .Z(n26754) );
  XNOR U27422 ( .A(n16632), .B(n26751), .Z(n26753) );
  XOR U27423 ( .A(n26755), .B(n26756), .Z(n16632) );
  XOR U27424 ( .A(n26757), .B(n26758), .Z(n26751) );
  AND U27425 ( .A(n26759), .B(n26760), .Z(n26758) );
  XOR U27426 ( .A(e_input[663]), .B(n26757), .Z(n26760) );
  XNOR U27427 ( .A(n16644), .B(n26757), .Z(n26759) );
  XOR U27428 ( .A(n26761), .B(n26762), .Z(n16644) );
  XOR U27429 ( .A(n26763), .B(n26764), .Z(n26757) );
  AND U27430 ( .A(n26765), .B(n26766), .Z(n26764) );
  XOR U27431 ( .A(e_input[662]), .B(n26763), .Z(n26766) );
  XNOR U27432 ( .A(n16656), .B(n26763), .Z(n26765) );
  XOR U27433 ( .A(n26767), .B(n26768), .Z(n16656) );
  XOR U27434 ( .A(n26769), .B(n26770), .Z(n26763) );
  AND U27435 ( .A(n26771), .B(n26772), .Z(n26770) );
  XOR U27436 ( .A(e_input[661]), .B(n26769), .Z(n26772) );
  XNOR U27437 ( .A(n16668), .B(n26769), .Z(n26771) );
  XOR U27438 ( .A(n26773), .B(n26774), .Z(n16668) );
  XOR U27439 ( .A(n26775), .B(n26776), .Z(n26769) );
  AND U27440 ( .A(n26777), .B(n26778), .Z(n26776) );
  XOR U27441 ( .A(e_input[660]), .B(n26775), .Z(n26778) );
  XNOR U27442 ( .A(n16680), .B(n26775), .Z(n26777) );
  XOR U27443 ( .A(n26779), .B(n26780), .Z(n16680) );
  XOR U27444 ( .A(n26781), .B(n26782), .Z(n26775) );
  AND U27445 ( .A(n26783), .B(n26784), .Z(n26782) );
  XOR U27446 ( .A(e_input[659]), .B(n26781), .Z(n26784) );
  XNOR U27447 ( .A(n16692), .B(n26781), .Z(n26783) );
  XOR U27448 ( .A(n26785), .B(n26786), .Z(n16692) );
  XOR U27449 ( .A(n26787), .B(n26788), .Z(n26781) );
  AND U27450 ( .A(n26789), .B(n26790), .Z(n26788) );
  XOR U27451 ( .A(e_input[658]), .B(n26787), .Z(n26790) );
  XNOR U27452 ( .A(n16704), .B(n26787), .Z(n26789) );
  XOR U27453 ( .A(n26791), .B(n26792), .Z(n16704) );
  XOR U27454 ( .A(n26793), .B(n26794), .Z(n26787) );
  AND U27455 ( .A(n26795), .B(n26796), .Z(n26794) );
  XOR U27456 ( .A(e_input[657]), .B(n26793), .Z(n26796) );
  XNOR U27457 ( .A(n16716), .B(n26793), .Z(n26795) );
  XOR U27458 ( .A(n26797), .B(n26798), .Z(n16716) );
  XOR U27459 ( .A(n26799), .B(n26800), .Z(n26793) );
  AND U27460 ( .A(n26801), .B(n26802), .Z(n26800) );
  XOR U27461 ( .A(e_input[656]), .B(n26799), .Z(n26802) );
  XNOR U27462 ( .A(n16728), .B(n26799), .Z(n26801) );
  XOR U27463 ( .A(n26803), .B(n26804), .Z(n16728) );
  XOR U27464 ( .A(n26805), .B(n26806), .Z(n26799) );
  AND U27465 ( .A(n26807), .B(n26808), .Z(n26806) );
  XOR U27466 ( .A(e_input[655]), .B(n26805), .Z(n26808) );
  XNOR U27467 ( .A(n16740), .B(n26805), .Z(n26807) );
  XOR U27468 ( .A(n26809), .B(n26810), .Z(n16740) );
  XOR U27469 ( .A(n26811), .B(n26812), .Z(n26805) );
  AND U27470 ( .A(n26813), .B(n26814), .Z(n26812) );
  XOR U27471 ( .A(e_input[654]), .B(n26811), .Z(n26814) );
  XNOR U27472 ( .A(n16752), .B(n26811), .Z(n26813) );
  XOR U27473 ( .A(n26815), .B(n26816), .Z(n16752) );
  XOR U27474 ( .A(n26817), .B(n26818), .Z(n26811) );
  AND U27475 ( .A(n26819), .B(n26820), .Z(n26818) );
  XOR U27476 ( .A(e_input[653]), .B(n26817), .Z(n26820) );
  XNOR U27477 ( .A(n16764), .B(n26817), .Z(n26819) );
  XOR U27478 ( .A(n26821), .B(n26822), .Z(n16764) );
  XOR U27479 ( .A(n26823), .B(n26824), .Z(n26817) );
  AND U27480 ( .A(n26825), .B(n26826), .Z(n26824) );
  XOR U27481 ( .A(e_input[652]), .B(n26823), .Z(n26826) );
  XNOR U27482 ( .A(n16776), .B(n26823), .Z(n26825) );
  XOR U27483 ( .A(n26827), .B(n26828), .Z(n16776) );
  XOR U27484 ( .A(n26829), .B(n26830), .Z(n26823) );
  AND U27485 ( .A(n26831), .B(n26832), .Z(n26830) );
  XOR U27486 ( .A(e_input[651]), .B(n26829), .Z(n26832) );
  XNOR U27487 ( .A(n16788), .B(n26829), .Z(n26831) );
  XOR U27488 ( .A(n26833), .B(n26834), .Z(n16788) );
  XOR U27489 ( .A(n26835), .B(n26836), .Z(n26829) );
  AND U27490 ( .A(n26837), .B(n26838), .Z(n26836) );
  XOR U27491 ( .A(e_input[650]), .B(n26835), .Z(n26838) );
  XNOR U27492 ( .A(n16800), .B(n26835), .Z(n26837) );
  XOR U27493 ( .A(n26839), .B(n26840), .Z(n16800) );
  XOR U27494 ( .A(n26841), .B(n26842), .Z(n26835) );
  AND U27495 ( .A(n26843), .B(n26844), .Z(n26842) );
  XOR U27496 ( .A(e_input[649]), .B(n26841), .Z(n26844) );
  XNOR U27497 ( .A(n16812), .B(n26841), .Z(n26843) );
  XOR U27498 ( .A(n26845), .B(n26846), .Z(n16812) );
  XOR U27499 ( .A(n26847), .B(n26848), .Z(n26841) );
  AND U27500 ( .A(n26849), .B(n26850), .Z(n26848) );
  XOR U27501 ( .A(e_input[648]), .B(n26847), .Z(n26850) );
  XNOR U27502 ( .A(n16824), .B(n26847), .Z(n26849) );
  XOR U27503 ( .A(n26851), .B(n26852), .Z(n16824) );
  XOR U27504 ( .A(n26853), .B(n26854), .Z(n26847) );
  AND U27505 ( .A(n26855), .B(n26856), .Z(n26854) );
  XOR U27506 ( .A(e_input[647]), .B(n26853), .Z(n26856) );
  XNOR U27507 ( .A(n16836), .B(n26853), .Z(n26855) );
  XOR U27508 ( .A(n26857), .B(n26858), .Z(n16836) );
  XOR U27509 ( .A(n26859), .B(n26860), .Z(n26853) );
  AND U27510 ( .A(n26861), .B(n26862), .Z(n26860) );
  XOR U27511 ( .A(e_input[646]), .B(n26859), .Z(n26862) );
  XNOR U27512 ( .A(n16848), .B(n26859), .Z(n26861) );
  XOR U27513 ( .A(n26863), .B(n26864), .Z(n16848) );
  XOR U27514 ( .A(n26865), .B(n26866), .Z(n26859) );
  AND U27515 ( .A(n26867), .B(n26868), .Z(n26866) );
  XOR U27516 ( .A(e_input[645]), .B(n26865), .Z(n26868) );
  XNOR U27517 ( .A(n16860), .B(n26865), .Z(n26867) );
  XOR U27518 ( .A(n26869), .B(n26870), .Z(n16860) );
  XOR U27519 ( .A(n26871), .B(n26872), .Z(n26865) );
  AND U27520 ( .A(n26873), .B(n26874), .Z(n26872) );
  XOR U27521 ( .A(e_input[644]), .B(n26871), .Z(n26874) );
  XNOR U27522 ( .A(n16872), .B(n26871), .Z(n26873) );
  XOR U27523 ( .A(n26875), .B(n26876), .Z(n16872) );
  XOR U27524 ( .A(n26877), .B(n26878), .Z(n26871) );
  AND U27525 ( .A(n26879), .B(n26880), .Z(n26878) );
  XOR U27526 ( .A(e_input[643]), .B(n26877), .Z(n26880) );
  XNOR U27527 ( .A(n16884), .B(n26877), .Z(n26879) );
  XOR U27528 ( .A(n26881), .B(n26882), .Z(n16884) );
  XOR U27529 ( .A(n26883), .B(n26884), .Z(n26877) );
  AND U27530 ( .A(n26885), .B(n26886), .Z(n26884) );
  XOR U27531 ( .A(e_input[642]), .B(n26883), .Z(n26886) );
  XNOR U27532 ( .A(n16896), .B(n26883), .Z(n26885) );
  XOR U27533 ( .A(n26887), .B(n26888), .Z(n16896) );
  XOR U27534 ( .A(n26889), .B(n26890), .Z(n26883) );
  AND U27535 ( .A(n26891), .B(n26892), .Z(n26890) );
  XOR U27536 ( .A(e_input[641]), .B(n26889), .Z(n26892) );
  XNOR U27537 ( .A(n16908), .B(n26889), .Z(n26891) );
  XOR U27538 ( .A(n26893), .B(n26894), .Z(n16908) );
  XOR U27539 ( .A(n26895), .B(n26896), .Z(n26889) );
  AND U27540 ( .A(n26897), .B(n26898), .Z(n26896) );
  XOR U27541 ( .A(e_input[640]), .B(n26895), .Z(n26898) );
  XNOR U27542 ( .A(n16920), .B(n26895), .Z(n26897) );
  XOR U27543 ( .A(n26899), .B(n26900), .Z(n16920) );
  XOR U27544 ( .A(n26901), .B(n26902), .Z(n26895) );
  AND U27545 ( .A(n26903), .B(n26904), .Z(n26902) );
  XOR U27546 ( .A(e_input[639]), .B(n26901), .Z(n26904) );
  XNOR U27547 ( .A(n16932), .B(n26901), .Z(n26903) );
  XOR U27548 ( .A(n26905), .B(n26906), .Z(n16932) );
  XOR U27549 ( .A(n26907), .B(n26908), .Z(n26901) );
  AND U27550 ( .A(n26909), .B(n26910), .Z(n26908) );
  XOR U27551 ( .A(e_input[638]), .B(n26907), .Z(n26910) );
  XNOR U27552 ( .A(n16944), .B(n26907), .Z(n26909) );
  XOR U27553 ( .A(n26911), .B(n26912), .Z(n16944) );
  XOR U27554 ( .A(n26913), .B(n26914), .Z(n26907) );
  AND U27555 ( .A(n26915), .B(n26916), .Z(n26914) );
  XOR U27556 ( .A(e_input[637]), .B(n26913), .Z(n26916) );
  XNOR U27557 ( .A(n16956), .B(n26913), .Z(n26915) );
  XOR U27558 ( .A(n26917), .B(n26918), .Z(n16956) );
  XOR U27559 ( .A(n26919), .B(n26920), .Z(n26913) );
  AND U27560 ( .A(n26921), .B(n26922), .Z(n26920) );
  XOR U27561 ( .A(e_input[636]), .B(n26919), .Z(n26922) );
  XNOR U27562 ( .A(n16968), .B(n26919), .Z(n26921) );
  XOR U27563 ( .A(n26923), .B(n26924), .Z(n16968) );
  XOR U27564 ( .A(n26925), .B(n26926), .Z(n26919) );
  AND U27565 ( .A(n26927), .B(n26928), .Z(n26926) );
  XOR U27566 ( .A(e_input[635]), .B(n26925), .Z(n26928) );
  XNOR U27567 ( .A(n16980), .B(n26925), .Z(n26927) );
  XOR U27568 ( .A(n26929), .B(n26930), .Z(n16980) );
  XOR U27569 ( .A(n26931), .B(n26932), .Z(n26925) );
  AND U27570 ( .A(n26933), .B(n26934), .Z(n26932) );
  XOR U27571 ( .A(e_input[634]), .B(n26931), .Z(n26934) );
  XNOR U27572 ( .A(n16992), .B(n26931), .Z(n26933) );
  XOR U27573 ( .A(n26935), .B(n26936), .Z(n16992) );
  XOR U27574 ( .A(n26937), .B(n26938), .Z(n26931) );
  AND U27575 ( .A(n26939), .B(n26940), .Z(n26938) );
  XOR U27576 ( .A(e_input[633]), .B(n26937), .Z(n26940) );
  XNOR U27577 ( .A(n17004), .B(n26937), .Z(n26939) );
  XOR U27578 ( .A(n26941), .B(n26942), .Z(n17004) );
  XOR U27579 ( .A(n26943), .B(n26944), .Z(n26937) );
  AND U27580 ( .A(n26945), .B(n26946), .Z(n26944) );
  XOR U27581 ( .A(e_input[632]), .B(n26943), .Z(n26946) );
  XNOR U27582 ( .A(n17016), .B(n26943), .Z(n26945) );
  XOR U27583 ( .A(n26947), .B(n26948), .Z(n17016) );
  XOR U27584 ( .A(n26949), .B(n26950), .Z(n26943) );
  AND U27585 ( .A(n26951), .B(n26952), .Z(n26950) );
  XOR U27586 ( .A(e_input[631]), .B(n26949), .Z(n26952) );
  XNOR U27587 ( .A(n17028), .B(n26949), .Z(n26951) );
  XOR U27588 ( .A(n26953), .B(n26954), .Z(n17028) );
  XOR U27589 ( .A(n26955), .B(n26956), .Z(n26949) );
  AND U27590 ( .A(n26957), .B(n26958), .Z(n26956) );
  XOR U27591 ( .A(e_input[630]), .B(n26955), .Z(n26958) );
  XNOR U27592 ( .A(n17040), .B(n26955), .Z(n26957) );
  XOR U27593 ( .A(n26959), .B(n26960), .Z(n17040) );
  XOR U27594 ( .A(n26961), .B(n26962), .Z(n26955) );
  AND U27595 ( .A(n26963), .B(n26964), .Z(n26962) );
  XOR U27596 ( .A(e_input[629]), .B(n26961), .Z(n26964) );
  XNOR U27597 ( .A(n17052), .B(n26961), .Z(n26963) );
  XOR U27598 ( .A(n26965), .B(n26966), .Z(n17052) );
  XOR U27599 ( .A(n26967), .B(n26968), .Z(n26961) );
  AND U27600 ( .A(n26969), .B(n26970), .Z(n26968) );
  XOR U27601 ( .A(e_input[628]), .B(n26967), .Z(n26970) );
  XNOR U27602 ( .A(n17064), .B(n26967), .Z(n26969) );
  XOR U27603 ( .A(n26971), .B(n26972), .Z(n17064) );
  XOR U27604 ( .A(n26973), .B(n26974), .Z(n26967) );
  AND U27605 ( .A(n26975), .B(n26976), .Z(n26974) );
  XOR U27606 ( .A(e_input[627]), .B(n26973), .Z(n26976) );
  XNOR U27607 ( .A(n17076), .B(n26973), .Z(n26975) );
  XOR U27608 ( .A(n26977), .B(n26978), .Z(n17076) );
  XOR U27609 ( .A(n26979), .B(n26980), .Z(n26973) );
  AND U27610 ( .A(n26981), .B(n26982), .Z(n26980) );
  XOR U27611 ( .A(e_input[626]), .B(n26979), .Z(n26982) );
  XNOR U27612 ( .A(n17088), .B(n26979), .Z(n26981) );
  XOR U27613 ( .A(n26983), .B(n26984), .Z(n17088) );
  XOR U27614 ( .A(n26985), .B(n26986), .Z(n26979) );
  AND U27615 ( .A(n26987), .B(n26988), .Z(n26986) );
  XOR U27616 ( .A(e_input[625]), .B(n26985), .Z(n26988) );
  XNOR U27617 ( .A(n17100), .B(n26985), .Z(n26987) );
  XOR U27618 ( .A(n26989), .B(n26990), .Z(n17100) );
  XOR U27619 ( .A(n26991), .B(n26992), .Z(n26985) );
  AND U27620 ( .A(n26993), .B(n26994), .Z(n26992) );
  XOR U27621 ( .A(e_input[624]), .B(n26991), .Z(n26994) );
  XNOR U27622 ( .A(n17112), .B(n26991), .Z(n26993) );
  XOR U27623 ( .A(n26995), .B(n26996), .Z(n17112) );
  XOR U27624 ( .A(n26997), .B(n26998), .Z(n26991) );
  AND U27625 ( .A(n26999), .B(n27000), .Z(n26998) );
  XOR U27626 ( .A(e_input[623]), .B(n26997), .Z(n27000) );
  XNOR U27627 ( .A(n17124), .B(n26997), .Z(n26999) );
  XOR U27628 ( .A(n27001), .B(n27002), .Z(n17124) );
  XOR U27629 ( .A(n27003), .B(n27004), .Z(n26997) );
  AND U27630 ( .A(n27005), .B(n27006), .Z(n27004) );
  XOR U27631 ( .A(e_input[622]), .B(n27003), .Z(n27006) );
  XNOR U27632 ( .A(n17136), .B(n27003), .Z(n27005) );
  XOR U27633 ( .A(n27007), .B(n27008), .Z(n17136) );
  XOR U27634 ( .A(n27009), .B(n27010), .Z(n27003) );
  AND U27635 ( .A(n27011), .B(n27012), .Z(n27010) );
  XOR U27636 ( .A(e_input[621]), .B(n27009), .Z(n27012) );
  XNOR U27637 ( .A(n17148), .B(n27009), .Z(n27011) );
  XOR U27638 ( .A(n27013), .B(n27014), .Z(n17148) );
  XOR U27639 ( .A(n27015), .B(n27016), .Z(n27009) );
  AND U27640 ( .A(n27017), .B(n27018), .Z(n27016) );
  XOR U27641 ( .A(e_input[620]), .B(n27015), .Z(n27018) );
  XNOR U27642 ( .A(n17160), .B(n27015), .Z(n27017) );
  XOR U27643 ( .A(n27019), .B(n27020), .Z(n17160) );
  XOR U27644 ( .A(n27021), .B(n27022), .Z(n27015) );
  AND U27645 ( .A(n27023), .B(n27024), .Z(n27022) );
  XOR U27646 ( .A(e_input[619]), .B(n27021), .Z(n27024) );
  XNOR U27647 ( .A(n17172), .B(n27021), .Z(n27023) );
  XOR U27648 ( .A(n27025), .B(n27026), .Z(n17172) );
  XOR U27649 ( .A(n27027), .B(n27028), .Z(n27021) );
  AND U27650 ( .A(n27029), .B(n27030), .Z(n27028) );
  XOR U27651 ( .A(e_input[618]), .B(n27027), .Z(n27030) );
  XNOR U27652 ( .A(n17184), .B(n27027), .Z(n27029) );
  XOR U27653 ( .A(n27031), .B(n27032), .Z(n17184) );
  XOR U27654 ( .A(n27033), .B(n27034), .Z(n27027) );
  AND U27655 ( .A(n27035), .B(n27036), .Z(n27034) );
  XOR U27656 ( .A(e_input[617]), .B(n27033), .Z(n27036) );
  XNOR U27657 ( .A(n17196), .B(n27033), .Z(n27035) );
  XOR U27658 ( .A(n27037), .B(n27038), .Z(n17196) );
  XOR U27659 ( .A(n27039), .B(n27040), .Z(n27033) );
  AND U27660 ( .A(n27041), .B(n27042), .Z(n27040) );
  XOR U27661 ( .A(e_input[616]), .B(n27039), .Z(n27042) );
  XNOR U27662 ( .A(n17208), .B(n27039), .Z(n27041) );
  XOR U27663 ( .A(n27043), .B(n27044), .Z(n17208) );
  XOR U27664 ( .A(n27045), .B(n27046), .Z(n27039) );
  AND U27665 ( .A(n27047), .B(n27048), .Z(n27046) );
  XOR U27666 ( .A(e_input[615]), .B(n27045), .Z(n27048) );
  XNOR U27667 ( .A(n17220), .B(n27045), .Z(n27047) );
  XOR U27668 ( .A(n27049), .B(n27050), .Z(n17220) );
  XOR U27669 ( .A(n27051), .B(n27052), .Z(n27045) );
  AND U27670 ( .A(n27053), .B(n27054), .Z(n27052) );
  XOR U27671 ( .A(e_input[614]), .B(n27051), .Z(n27054) );
  XNOR U27672 ( .A(n17232), .B(n27051), .Z(n27053) );
  XOR U27673 ( .A(n27055), .B(n27056), .Z(n17232) );
  XOR U27674 ( .A(n27057), .B(n27058), .Z(n27051) );
  AND U27675 ( .A(n27059), .B(n27060), .Z(n27058) );
  XOR U27676 ( .A(e_input[613]), .B(n27057), .Z(n27060) );
  XNOR U27677 ( .A(n17244), .B(n27057), .Z(n27059) );
  XOR U27678 ( .A(n27061), .B(n27062), .Z(n17244) );
  XOR U27679 ( .A(n27063), .B(n27064), .Z(n27057) );
  AND U27680 ( .A(n27065), .B(n27066), .Z(n27064) );
  XOR U27681 ( .A(e_input[612]), .B(n27063), .Z(n27066) );
  XNOR U27682 ( .A(n17256), .B(n27063), .Z(n27065) );
  XOR U27683 ( .A(n27067), .B(n27068), .Z(n17256) );
  XOR U27684 ( .A(n27069), .B(n27070), .Z(n27063) );
  AND U27685 ( .A(n27071), .B(n27072), .Z(n27070) );
  XOR U27686 ( .A(e_input[611]), .B(n27069), .Z(n27072) );
  XNOR U27687 ( .A(n17268), .B(n27069), .Z(n27071) );
  XOR U27688 ( .A(n27073), .B(n27074), .Z(n17268) );
  XOR U27689 ( .A(n27075), .B(n27076), .Z(n27069) );
  AND U27690 ( .A(n27077), .B(n27078), .Z(n27076) );
  XOR U27691 ( .A(e_input[610]), .B(n27075), .Z(n27078) );
  XNOR U27692 ( .A(n17280), .B(n27075), .Z(n27077) );
  XOR U27693 ( .A(n27079), .B(n27080), .Z(n17280) );
  XOR U27694 ( .A(n27081), .B(n27082), .Z(n27075) );
  AND U27695 ( .A(n27083), .B(n27084), .Z(n27082) );
  XOR U27696 ( .A(e_input[609]), .B(n27081), .Z(n27084) );
  XNOR U27697 ( .A(n17292), .B(n27081), .Z(n27083) );
  XOR U27698 ( .A(n27085), .B(n27086), .Z(n17292) );
  XOR U27699 ( .A(n27087), .B(n27088), .Z(n27081) );
  AND U27700 ( .A(n27089), .B(n27090), .Z(n27088) );
  XOR U27701 ( .A(e_input[608]), .B(n27087), .Z(n27090) );
  XNOR U27702 ( .A(n17304), .B(n27087), .Z(n27089) );
  XOR U27703 ( .A(n27091), .B(n27092), .Z(n17304) );
  XOR U27704 ( .A(n27093), .B(n27094), .Z(n27087) );
  AND U27705 ( .A(n27095), .B(n27096), .Z(n27094) );
  XOR U27706 ( .A(e_input[607]), .B(n27093), .Z(n27096) );
  XNOR U27707 ( .A(n17316), .B(n27093), .Z(n27095) );
  XOR U27708 ( .A(n27097), .B(n27098), .Z(n17316) );
  XOR U27709 ( .A(n27099), .B(n27100), .Z(n27093) );
  AND U27710 ( .A(n27101), .B(n27102), .Z(n27100) );
  XOR U27711 ( .A(e_input[606]), .B(n27099), .Z(n27102) );
  XNOR U27712 ( .A(n17328), .B(n27099), .Z(n27101) );
  XOR U27713 ( .A(n27103), .B(n27104), .Z(n17328) );
  XOR U27714 ( .A(n27105), .B(n27106), .Z(n27099) );
  AND U27715 ( .A(n27107), .B(n27108), .Z(n27106) );
  XOR U27716 ( .A(e_input[605]), .B(n27105), .Z(n27108) );
  XNOR U27717 ( .A(n17340), .B(n27105), .Z(n27107) );
  XOR U27718 ( .A(n27109), .B(n27110), .Z(n17340) );
  XOR U27719 ( .A(n27111), .B(n27112), .Z(n27105) );
  AND U27720 ( .A(n27113), .B(n27114), .Z(n27112) );
  XOR U27721 ( .A(e_input[604]), .B(n27111), .Z(n27114) );
  XNOR U27722 ( .A(n17352), .B(n27111), .Z(n27113) );
  XOR U27723 ( .A(n27115), .B(n27116), .Z(n17352) );
  XOR U27724 ( .A(n27117), .B(n27118), .Z(n27111) );
  AND U27725 ( .A(n27119), .B(n27120), .Z(n27118) );
  XOR U27726 ( .A(e_input[603]), .B(n27117), .Z(n27120) );
  XNOR U27727 ( .A(n17364), .B(n27117), .Z(n27119) );
  XOR U27728 ( .A(n27121), .B(n27122), .Z(n17364) );
  XOR U27729 ( .A(n27123), .B(n27124), .Z(n27117) );
  AND U27730 ( .A(n27125), .B(n27126), .Z(n27124) );
  XOR U27731 ( .A(e_input[602]), .B(n27123), .Z(n27126) );
  XNOR U27732 ( .A(n17376), .B(n27123), .Z(n27125) );
  XOR U27733 ( .A(n27127), .B(n27128), .Z(n17376) );
  XOR U27734 ( .A(n27129), .B(n27130), .Z(n27123) );
  AND U27735 ( .A(n27131), .B(n27132), .Z(n27130) );
  XOR U27736 ( .A(e_input[601]), .B(n27129), .Z(n27132) );
  XNOR U27737 ( .A(n17388), .B(n27129), .Z(n27131) );
  XOR U27738 ( .A(n27133), .B(n27134), .Z(n17388) );
  XOR U27739 ( .A(n27135), .B(n27136), .Z(n27129) );
  AND U27740 ( .A(n27137), .B(n27138), .Z(n27136) );
  XOR U27741 ( .A(e_input[600]), .B(n27135), .Z(n27138) );
  XNOR U27742 ( .A(n17400), .B(n27135), .Z(n27137) );
  XOR U27743 ( .A(n27139), .B(n27140), .Z(n17400) );
  XOR U27744 ( .A(n27141), .B(n27142), .Z(n27135) );
  AND U27745 ( .A(n27143), .B(n27144), .Z(n27142) );
  XOR U27746 ( .A(e_input[599]), .B(n27141), .Z(n27144) );
  XNOR U27747 ( .A(n17412), .B(n27141), .Z(n27143) );
  XOR U27748 ( .A(n27145), .B(n27146), .Z(n17412) );
  XOR U27749 ( .A(n27147), .B(n27148), .Z(n27141) );
  AND U27750 ( .A(n27149), .B(n27150), .Z(n27148) );
  XOR U27751 ( .A(e_input[598]), .B(n27147), .Z(n27150) );
  XNOR U27752 ( .A(n17424), .B(n27147), .Z(n27149) );
  XOR U27753 ( .A(n27151), .B(n27152), .Z(n17424) );
  XOR U27754 ( .A(n27153), .B(n27154), .Z(n27147) );
  AND U27755 ( .A(n27155), .B(n27156), .Z(n27154) );
  XOR U27756 ( .A(e_input[597]), .B(n27153), .Z(n27156) );
  XNOR U27757 ( .A(n17436), .B(n27153), .Z(n27155) );
  XOR U27758 ( .A(n27157), .B(n27158), .Z(n17436) );
  XOR U27759 ( .A(n27159), .B(n27160), .Z(n27153) );
  AND U27760 ( .A(n27161), .B(n27162), .Z(n27160) );
  XOR U27761 ( .A(e_input[596]), .B(n27159), .Z(n27162) );
  XNOR U27762 ( .A(n17448), .B(n27159), .Z(n27161) );
  XOR U27763 ( .A(n27163), .B(n27164), .Z(n17448) );
  XOR U27764 ( .A(n27165), .B(n27166), .Z(n27159) );
  AND U27765 ( .A(n27167), .B(n27168), .Z(n27166) );
  XOR U27766 ( .A(e_input[595]), .B(n27165), .Z(n27168) );
  XNOR U27767 ( .A(n17460), .B(n27165), .Z(n27167) );
  XOR U27768 ( .A(n27169), .B(n27170), .Z(n17460) );
  XOR U27769 ( .A(n27171), .B(n27172), .Z(n27165) );
  AND U27770 ( .A(n27173), .B(n27174), .Z(n27172) );
  XOR U27771 ( .A(e_input[594]), .B(n27171), .Z(n27174) );
  XNOR U27772 ( .A(n17472), .B(n27171), .Z(n27173) );
  XOR U27773 ( .A(n27175), .B(n27176), .Z(n17472) );
  XOR U27774 ( .A(n27177), .B(n27178), .Z(n27171) );
  AND U27775 ( .A(n27179), .B(n27180), .Z(n27178) );
  XOR U27776 ( .A(e_input[593]), .B(n27177), .Z(n27180) );
  XNOR U27777 ( .A(n17484), .B(n27177), .Z(n27179) );
  XOR U27778 ( .A(n27181), .B(n27182), .Z(n17484) );
  XOR U27779 ( .A(n27183), .B(n27184), .Z(n27177) );
  AND U27780 ( .A(n27185), .B(n27186), .Z(n27184) );
  XOR U27781 ( .A(e_input[592]), .B(n27183), .Z(n27186) );
  XNOR U27782 ( .A(n17496), .B(n27183), .Z(n27185) );
  XOR U27783 ( .A(n27187), .B(n27188), .Z(n17496) );
  XOR U27784 ( .A(n27189), .B(n27190), .Z(n27183) );
  AND U27785 ( .A(n27191), .B(n27192), .Z(n27190) );
  XOR U27786 ( .A(e_input[591]), .B(n27189), .Z(n27192) );
  XNOR U27787 ( .A(n17508), .B(n27189), .Z(n27191) );
  XOR U27788 ( .A(n27193), .B(n27194), .Z(n17508) );
  XOR U27789 ( .A(n27195), .B(n27196), .Z(n27189) );
  AND U27790 ( .A(n27197), .B(n27198), .Z(n27196) );
  XOR U27791 ( .A(e_input[590]), .B(n27195), .Z(n27198) );
  XNOR U27792 ( .A(n17520), .B(n27195), .Z(n27197) );
  XOR U27793 ( .A(n27199), .B(n27200), .Z(n17520) );
  XOR U27794 ( .A(n27201), .B(n27202), .Z(n27195) );
  AND U27795 ( .A(n27203), .B(n27204), .Z(n27202) );
  XOR U27796 ( .A(e_input[589]), .B(n27201), .Z(n27204) );
  XNOR U27797 ( .A(n17532), .B(n27201), .Z(n27203) );
  XOR U27798 ( .A(n27205), .B(n27206), .Z(n17532) );
  XOR U27799 ( .A(n27207), .B(n27208), .Z(n27201) );
  AND U27800 ( .A(n27209), .B(n27210), .Z(n27208) );
  XOR U27801 ( .A(e_input[588]), .B(n27207), .Z(n27210) );
  XNOR U27802 ( .A(n17544), .B(n27207), .Z(n27209) );
  XOR U27803 ( .A(n27211), .B(n27212), .Z(n17544) );
  XOR U27804 ( .A(n27213), .B(n27214), .Z(n27207) );
  AND U27805 ( .A(n27215), .B(n27216), .Z(n27214) );
  XOR U27806 ( .A(e_input[587]), .B(n27213), .Z(n27216) );
  XNOR U27807 ( .A(n17556), .B(n27213), .Z(n27215) );
  XOR U27808 ( .A(n27217), .B(n27218), .Z(n17556) );
  XOR U27809 ( .A(n27219), .B(n27220), .Z(n27213) );
  AND U27810 ( .A(n27221), .B(n27222), .Z(n27220) );
  XOR U27811 ( .A(e_input[586]), .B(n27219), .Z(n27222) );
  XNOR U27812 ( .A(n17568), .B(n27219), .Z(n27221) );
  XOR U27813 ( .A(n27223), .B(n27224), .Z(n17568) );
  XOR U27814 ( .A(n27225), .B(n27226), .Z(n27219) );
  AND U27815 ( .A(n27227), .B(n27228), .Z(n27226) );
  XOR U27816 ( .A(e_input[585]), .B(n27225), .Z(n27228) );
  XNOR U27817 ( .A(n17580), .B(n27225), .Z(n27227) );
  XOR U27818 ( .A(n27229), .B(n27230), .Z(n17580) );
  XOR U27819 ( .A(n27231), .B(n27232), .Z(n27225) );
  AND U27820 ( .A(n27233), .B(n27234), .Z(n27232) );
  XOR U27821 ( .A(e_input[584]), .B(n27231), .Z(n27234) );
  XNOR U27822 ( .A(n17592), .B(n27231), .Z(n27233) );
  XOR U27823 ( .A(n27235), .B(n27236), .Z(n17592) );
  XOR U27824 ( .A(n27237), .B(n27238), .Z(n27231) );
  AND U27825 ( .A(n27239), .B(n27240), .Z(n27238) );
  XOR U27826 ( .A(e_input[583]), .B(n27237), .Z(n27240) );
  XNOR U27827 ( .A(n17604), .B(n27237), .Z(n27239) );
  XOR U27828 ( .A(n27241), .B(n27242), .Z(n17604) );
  XOR U27829 ( .A(n27243), .B(n27244), .Z(n27237) );
  AND U27830 ( .A(n27245), .B(n27246), .Z(n27244) );
  XOR U27831 ( .A(e_input[582]), .B(n27243), .Z(n27246) );
  XNOR U27832 ( .A(n17616), .B(n27243), .Z(n27245) );
  XOR U27833 ( .A(n27247), .B(n27248), .Z(n17616) );
  XOR U27834 ( .A(n27249), .B(n27250), .Z(n27243) );
  AND U27835 ( .A(n27251), .B(n27252), .Z(n27250) );
  XOR U27836 ( .A(e_input[581]), .B(n27249), .Z(n27252) );
  XNOR U27837 ( .A(n17628), .B(n27249), .Z(n27251) );
  XOR U27838 ( .A(n27253), .B(n27254), .Z(n17628) );
  XOR U27839 ( .A(n27255), .B(n27256), .Z(n27249) );
  AND U27840 ( .A(n27257), .B(n27258), .Z(n27256) );
  XOR U27841 ( .A(e_input[580]), .B(n27255), .Z(n27258) );
  XNOR U27842 ( .A(n17640), .B(n27255), .Z(n27257) );
  XOR U27843 ( .A(n27259), .B(n27260), .Z(n17640) );
  XOR U27844 ( .A(n27261), .B(n27262), .Z(n27255) );
  AND U27845 ( .A(n27263), .B(n27264), .Z(n27262) );
  XOR U27846 ( .A(e_input[579]), .B(n27261), .Z(n27264) );
  XNOR U27847 ( .A(n17652), .B(n27261), .Z(n27263) );
  XOR U27848 ( .A(n27265), .B(n27266), .Z(n17652) );
  XOR U27849 ( .A(n27267), .B(n27268), .Z(n27261) );
  AND U27850 ( .A(n27269), .B(n27270), .Z(n27268) );
  XOR U27851 ( .A(e_input[578]), .B(n27267), .Z(n27270) );
  XNOR U27852 ( .A(n17664), .B(n27267), .Z(n27269) );
  XOR U27853 ( .A(n27271), .B(n27272), .Z(n17664) );
  XOR U27854 ( .A(n27273), .B(n27274), .Z(n27267) );
  AND U27855 ( .A(n27275), .B(n27276), .Z(n27274) );
  XOR U27856 ( .A(e_input[577]), .B(n27273), .Z(n27276) );
  XNOR U27857 ( .A(n17676), .B(n27273), .Z(n27275) );
  XOR U27858 ( .A(n27277), .B(n27278), .Z(n17676) );
  XOR U27859 ( .A(n27279), .B(n27280), .Z(n27273) );
  AND U27860 ( .A(n27281), .B(n27282), .Z(n27280) );
  XOR U27861 ( .A(e_input[576]), .B(n27279), .Z(n27282) );
  XNOR U27862 ( .A(n17688), .B(n27279), .Z(n27281) );
  XOR U27863 ( .A(n27283), .B(n27284), .Z(n17688) );
  XOR U27864 ( .A(n27285), .B(n27286), .Z(n27279) );
  AND U27865 ( .A(n27287), .B(n27288), .Z(n27286) );
  XOR U27866 ( .A(e_input[575]), .B(n27285), .Z(n27288) );
  XNOR U27867 ( .A(n17700), .B(n27285), .Z(n27287) );
  XOR U27868 ( .A(n27289), .B(n27290), .Z(n17700) );
  XOR U27869 ( .A(n27291), .B(n27292), .Z(n27285) );
  AND U27870 ( .A(n27293), .B(n27294), .Z(n27292) );
  XOR U27871 ( .A(e_input[574]), .B(n27291), .Z(n27294) );
  XNOR U27872 ( .A(n17712), .B(n27291), .Z(n27293) );
  XOR U27873 ( .A(n27295), .B(n27296), .Z(n17712) );
  XOR U27874 ( .A(n27297), .B(n27298), .Z(n27291) );
  AND U27875 ( .A(n27299), .B(n27300), .Z(n27298) );
  XOR U27876 ( .A(e_input[573]), .B(n27297), .Z(n27300) );
  XNOR U27877 ( .A(n17724), .B(n27297), .Z(n27299) );
  XOR U27878 ( .A(n27301), .B(n27302), .Z(n17724) );
  XOR U27879 ( .A(n27303), .B(n27304), .Z(n27297) );
  AND U27880 ( .A(n27305), .B(n27306), .Z(n27304) );
  XOR U27881 ( .A(e_input[572]), .B(n27303), .Z(n27306) );
  XNOR U27882 ( .A(n17736), .B(n27303), .Z(n27305) );
  XOR U27883 ( .A(n27307), .B(n27308), .Z(n17736) );
  XOR U27884 ( .A(n27309), .B(n27310), .Z(n27303) );
  AND U27885 ( .A(n27311), .B(n27312), .Z(n27310) );
  XOR U27886 ( .A(e_input[571]), .B(n27309), .Z(n27312) );
  XNOR U27887 ( .A(n17748), .B(n27309), .Z(n27311) );
  XOR U27888 ( .A(n27313), .B(n27314), .Z(n17748) );
  XOR U27889 ( .A(n27315), .B(n27316), .Z(n27309) );
  AND U27890 ( .A(n27317), .B(n27318), .Z(n27316) );
  XOR U27891 ( .A(e_input[570]), .B(n27315), .Z(n27318) );
  XNOR U27892 ( .A(n17760), .B(n27315), .Z(n27317) );
  XOR U27893 ( .A(n27319), .B(n27320), .Z(n17760) );
  XOR U27894 ( .A(n27321), .B(n27322), .Z(n27315) );
  AND U27895 ( .A(n27323), .B(n27324), .Z(n27322) );
  XOR U27896 ( .A(e_input[569]), .B(n27321), .Z(n27324) );
  XNOR U27897 ( .A(n17772), .B(n27321), .Z(n27323) );
  XOR U27898 ( .A(n27325), .B(n27326), .Z(n17772) );
  XOR U27899 ( .A(n27327), .B(n27328), .Z(n27321) );
  AND U27900 ( .A(n27329), .B(n27330), .Z(n27328) );
  XOR U27901 ( .A(e_input[568]), .B(n27327), .Z(n27330) );
  XNOR U27902 ( .A(n17784), .B(n27327), .Z(n27329) );
  XOR U27903 ( .A(n27331), .B(n27332), .Z(n17784) );
  XOR U27904 ( .A(n27333), .B(n27334), .Z(n27327) );
  AND U27905 ( .A(n27335), .B(n27336), .Z(n27334) );
  XOR U27906 ( .A(e_input[567]), .B(n27333), .Z(n27336) );
  XNOR U27907 ( .A(n17796), .B(n27333), .Z(n27335) );
  XOR U27908 ( .A(n27337), .B(n27338), .Z(n17796) );
  XOR U27909 ( .A(n27339), .B(n27340), .Z(n27333) );
  AND U27910 ( .A(n27341), .B(n27342), .Z(n27340) );
  XOR U27911 ( .A(e_input[566]), .B(n27339), .Z(n27342) );
  XNOR U27912 ( .A(n17808), .B(n27339), .Z(n27341) );
  XOR U27913 ( .A(n27343), .B(n27344), .Z(n17808) );
  XOR U27914 ( .A(n27345), .B(n27346), .Z(n27339) );
  AND U27915 ( .A(n27347), .B(n27348), .Z(n27346) );
  XOR U27916 ( .A(e_input[565]), .B(n27345), .Z(n27348) );
  XNOR U27917 ( .A(n17820), .B(n27345), .Z(n27347) );
  XOR U27918 ( .A(n27349), .B(n27350), .Z(n17820) );
  XOR U27919 ( .A(n27351), .B(n27352), .Z(n27345) );
  AND U27920 ( .A(n27353), .B(n27354), .Z(n27352) );
  XOR U27921 ( .A(e_input[564]), .B(n27351), .Z(n27354) );
  XNOR U27922 ( .A(n17832), .B(n27351), .Z(n27353) );
  XOR U27923 ( .A(n27355), .B(n27356), .Z(n17832) );
  XOR U27924 ( .A(n27357), .B(n27358), .Z(n27351) );
  AND U27925 ( .A(n27359), .B(n27360), .Z(n27358) );
  XOR U27926 ( .A(e_input[563]), .B(n27357), .Z(n27360) );
  XNOR U27927 ( .A(n17844), .B(n27357), .Z(n27359) );
  XOR U27928 ( .A(n27361), .B(n27362), .Z(n17844) );
  XOR U27929 ( .A(n27363), .B(n27364), .Z(n27357) );
  AND U27930 ( .A(n27365), .B(n27366), .Z(n27364) );
  XOR U27931 ( .A(e_input[562]), .B(n27363), .Z(n27366) );
  XNOR U27932 ( .A(n17856), .B(n27363), .Z(n27365) );
  XOR U27933 ( .A(n27367), .B(n27368), .Z(n17856) );
  XOR U27934 ( .A(n27369), .B(n27370), .Z(n27363) );
  AND U27935 ( .A(n27371), .B(n27372), .Z(n27370) );
  XOR U27936 ( .A(e_input[561]), .B(n27369), .Z(n27372) );
  XNOR U27937 ( .A(n17868), .B(n27369), .Z(n27371) );
  XOR U27938 ( .A(n27373), .B(n27374), .Z(n17868) );
  XOR U27939 ( .A(n27375), .B(n27376), .Z(n27369) );
  AND U27940 ( .A(n27377), .B(n27378), .Z(n27376) );
  XOR U27941 ( .A(e_input[560]), .B(n27375), .Z(n27378) );
  XNOR U27942 ( .A(n17880), .B(n27375), .Z(n27377) );
  XOR U27943 ( .A(n27379), .B(n27380), .Z(n17880) );
  XOR U27944 ( .A(n27381), .B(n27382), .Z(n27375) );
  AND U27945 ( .A(n27383), .B(n27384), .Z(n27382) );
  XOR U27946 ( .A(e_input[559]), .B(n27381), .Z(n27384) );
  XNOR U27947 ( .A(n17892), .B(n27381), .Z(n27383) );
  XOR U27948 ( .A(n27385), .B(n27386), .Z(n17892) );
  XOR U27949 ( .A(n27387), .B(n27388), .Z(n27381) );
  AND U27950 ( .A(n27389), .B(n27390), .Z(n27388) );
  XOR U27951 ( .A(e_input[558]), .B(n27387), .Z(n27390) );
  XNOR U27952 ( .A(n17904), .B(n27387), .Z(n27389) );
  XOR U27953 ( .A(n27391), .B(n27392), .Z(n17904) );
  XOR U27954 ( .A(n27393), .B(n27394), .Z(n27387) );
  AND U27955 ( .A(n27395), .B(n27396), .Z(n27394) );
  XOR U27956 ( .A(e_input[557]), .B(n27393), .Z(n27396) );
  XNOR U27957 ( .A(n17916), .B(n27393), .Z(n27395) );
  XOR U27958 ( .A(n27397), .B(n27398), .Z(n17916) );
  XOR U27959 ( .A(n27399), .B(n27400), .Z(n27393) );
  AND U27960 ( .A(n27401), .B(n27402), .Z(n27400) );
  XOR U27961 ( .A(e_input[556]), .B(n27399), .Z(n27402) );
  XNOR U27962 ( .A(n17928), .B(n27399), .Z(n27401) );
  XOR U27963 ( .A(n27403), .B(n27404), .Z(n17928) );
  XOR U27964 ( .A(n27405), .B(n27406), .Z(n27399) );
  AND U27965 ( .A(n27407), .B(n27408), .Z(n27406) );
  XOR U27966 ( .A(e_input[555]), .B(n27405), .Z(n27408) );
  XNOR U27967 ( .A(n17940), .B(n27405), .Z(n27407) );
  XOR U27968 ( .A(n27409), .B(n27410), .Z(n17940) );
  XOR U27969 ( .A(n27411), .B(n27412), .Z(n27405) );
  AND U27970 ( .A(n27413), .B(n27414), .Z(n27412) );
  XOR U27971 ( .A(e_input[554]), .B(n27411), .Z(n27414) );
  XNOR U27972 ( .A(n17952), .B(n27411), .Z(n27413) );
  XOR U27973 ( .A(n27415), .B(n27416), .Z(n17952) );
  XOR U27974 ( .A(n27417), .B(n27418), .Z(n27411) );
  AND U27975 ( .A(n27419), .B(n27420), .Z(n27418) );
  XOR U27976 ( .A(e_input[553]), .B(n27417), .Z(n27420) );
  XNOR U27977 ( .A(n17964), .B(n27417), .Z(n27419) );
  XOR U27978 ( .A(n27421), .B(n27422), .Z(n17964) );
  XOR U27979 ( .A(n27423), .B(n27424), .Z(n27417) );
  AND U27980 ( .A(n27425), .B(n27426), .Z(n27424) );
  XOR U27981 ( .A(e_input[552]), .B(n27423), .Z(n27426) );
  XNOR U27982 ( .A(n17976), .B(n27423), .Z(n27425) );
  XOR U27983 ( .A(n27427), .B(n27428), .Z(n17976) );
  XOR U27984 ( .A(n27429), .B(n27430), .Z(n27423) );
  AND U27985 ( .A(n27431), .B(n27432), .Z(n27430) );
  XOR U27986 ( .A(e_input[551]), .B(n27429), .Z(n27432) );
  XNOR U27987 ( .A(n17988), .B(n27429), .Z(n27431) );
  XOR U27988 ( .A(n27433), .B(n27434), .Z(n17988) );
  XOR U27989 ( .A(n27435), .B(n27436), .Z(n27429) );
  AND U27990 ( .A(n27437), .B(n27438), .Z(n27436) );
  XOR U27991 ( .A(e_input[550]), .B(n27435), .Z(n27438) );
  XNOR U27992 ( .A(n18000), .B(n27435), .Z(n27437) );
  XOR U27993 ( .A(n27439), .B(n27440), .Z(n18000) );
  XOR U27994 ( .A(n27441), .B(n27442), .Z(n27435) );
  AND U27995 ( .A(n27443), .B(n27444), .Z(n27442) );
  XOR U27996 ( .A(e_input[549]), .B(n27441), .Z(n27444) );
  XNOR U27997 ( .A(n18012), .B(n27441), .Z(n27443) );
  XOR U27998 ( .A(n27445), .B(n27446), .Z(n18012) );
  XOR U27999 ( .A(n27447), .B(n27448), .Z(n27441) );
  AND U28000 ( .A(n27449), .B(n27450), .Z(n27448) );
  XOR U28001 ( .A(e_input[548]), .B(n27447), .Z(n27450) );
  XNOR U28002 ( .A(n18024), .B(n27447), .Z(n27449) );
  XOR U28003 ( .A(n27451), .B(n27452), .Z(n18024) );
  XOR U28004 ( .A(n27453), .B(n27454), .Z(n27447) );
  AND U28005 ( .A(n27455), .B(n27456), .Z(n27454) );
  XOR U28006 ( .A(e_input[547]), .B(n27453), .Z(n27456) );
  XNOR U28007 ( .A(n18036), .B(n27453), .Z(n27455) );
  XOR U28008 ( .A(n27457), .B(n27458), .Z(n18036) );
  XOR U28009 ( .A(n27459), .B(n27460), .Z(n27453) );
  AND U28010 ( .A(n27461), .B(n27462), .Z(n27460) );
  XOR U28011 ( .A(e_input[546]), .B(n27459), .Z(n27462) );
  XNOR U28012 ( .A(n18048), .B(n27459), .Z(n27461) );
  XOR U28013 ( .A(n27463), .B(n27464), .Z(n18048) );
  XOR U28014 ( .A(n27465), .B(n27466), .Z(n27459) );
  AND U28015 ( .A(n27467), .B(n27468), .Z(n27466) );
  XOR U28016 ( .A(e_input[545]), .B(n27465), .Z(n27468) );
  XNOR U28017 ( .A(n18060), .B(n27465), .Z(n27467) );
  XOR U28018 ( .A(n27469), .B(n27470), .Z(n18060) );
  XOR U28019 ( .A(n27471), .B(n27472), .Z(n27465) );
  AND U28020 ( .A(n27473), .B(n27474), .Z(n27472) );
  XOR U28021 ( .A(e_input[544]), .B(n27471), .Z(n27474) );
  XNOR U28022 ( .A(n18072), .B(n27471), .Z(n27473) );
  XOR U28023 ( .A(n27475), .B(n27476), .Z(n18072) );
  XOR U28024 ( .A(n27477), .B(n27478), .Z(n27471) );
  AND U28025 ( .A(n27479), .B(n27480), .Z(n27478) );
  XOR U28026 ( .A(e_input[543]), .B(n27477), .Z(n27480) );
  XNOR U28027 ( .A(n18084), .B(n27477), .Z(n27479) );
  XOR U28028 ( .A(n27481), .B(n27482), .Z(n18084) );
  XOR U28029 ( .A(n27483), .B(n27484), .Z(n27477) );
  AND U28030 ( .A(n27485), .B(n27486), .Z(n27484) );
  XOR U28031 ( .A(e_input[542]), .B(n27483), .Z(n27486) );
  XNOR U28032 ( .A(n18096), .B(n27483), .Z(n27485) );
  XOR U28033 ( .A(n27487), .B(n27488), .Z(n18096) );
  XOR U28034 ( .A(n27489), .B(n27490), .Z(n27483) );
  AND U28035 ( .A(n27491), .B(n27492), .Z(n27490) );
  XOR U28036 ( .A(e_input[541]), .B(n27489), .Z(n27492) );
  XNOR U28037 ( .A(n18108), .B(n27489), .Z(n27491) );
  XOR U28038 ( .A(n27493), .B(n27494), .Z(n18108) );
  XOR U28039 ( .A(n27495), .B(n27496), .Z(n27489) );
  AND U28040 ( .A(n27497), .B(n27498), .Z(n27496) );
  XOR U28041 ( .A(e_input[540]), .B(n27495), .Z(n27498) );
  XNOR U28042 ( .A(n18120), .B(n27495), .Z(n27497) );
  XOR U28043 ( .A(n27499), .B(n27500), .Z(n18120) );
  XOR U28044 ( .A(n27501), .B(n27502), .Z(n27495) );
  AND U28045 ( .A(n27503), .B(n27504), .Z(n27502) );
  XOR U28046 ( .A(e_input[539]), .B(n27501), .Z(n27504) );
  XNOR U28047 ( .A(n18132), .B(n27501), .Z(n27503) );
  XOR U28048 ( .A(n27505), .B(n27506), .Z(n18132) );
  XOR U28049 ( .A(n27507), .B(n27508), .Z(n27501) );
  AND U28050 ( .A(n27509), .B(n27510), .Z(n27508) );
  XOR U28051 ( .A(e_input[538]), .B(n27507), .Z(n27510) );
  XNOR U28052 ( .A(n18144), .B(n27507), .Z(n27509) );
  XOR U28053 ( .A(n27511), .B(n27512), .Z(n18144) );
  XOR U28054 ( .A(n27513), .B(n27514), .Z(n27507) );
  AND U28055 ( .A(n27515), .B(n27516), .Z(n27514) );
  XOR U28056 ( .A(e_input[537]), .B(n27513), .Z(n27516) );
  XNOR U28057 ( .A(n18156), .B(n27513), .Z(n27515) );
  XOR U28058 ( .A(n27517), .B(n27518), .Z(n18156) );
  XOR U28059 ( .A(n27519), .B(n27520), .Z(n27513) );
  AND U28060 ( .A(n27521), .B(n27522), .Z(n27520) );
  XOR U28061 ( .A(e_input[536]), .B(n27519), .Z(n27522) );
  XNOR U28062 ( .A(n18168), .B(n27519), .Z(n27521) );
  XOR U28063 ( .A(n27523), .B(n27524), .Z(n18168) );
  XOR U28064 ( .A(n27525), .B(n27526), .Z(n27519) );
  AND U28065 ( .A(n27527), .B(n27528), .Z(n27526) );
  XOR U28066 ( .A(e_input[535]), .B(n27525), .Z(n27528) );
  XNOR U28067 ( .A(n18180), .B(n27525), .Z(n27527) );
  XOR U28068 ( .A(n27529), .B(n27530), .Z(n18180) );
  XOR U28069 ( .A(n27531), .B(n27532), .Z(n27525) );
  AND U28070 ( .A(n27533), .B(n27534), .Z(n27532) );
  XOR U28071 ( .A(e_input[534]), .B(n27531), .Z(n27534) );
  XNOR U28072 ( .A(n18192), .B(n27531), .Z(n27533) );
  XOR U28073 ( .A(n27535), .B(n27536), .Z(n18192) );
  XOR U28074 ( .A(n27537), .B(n27538), .Z(n27531) );
  AND U28075 ( .A(n27539), .B(n27540), .Z(n27538) );
  XOR U28076 ( .A(e_input[533]), .B(n27537), .Z(n27540) );
  XNOR U28077 ( .A(n18204), .B(n27537), .Z(n27539) );
  XOR U28078 ( .A(n27541), .B(n27542), .Z(n18204) );
  XOR U28079 ( .A(n27543), .B(n27544), .Z(n27537) );
  AND U28080 ( .A(n27545), .B(n27546), .Z(n27544) );
  XOR U28081 ( .A(e_input[532]), .B(n27543), .Z(n27546) );
  XNOR U28082 ( .A(n18216), .B(n27543), .Z(n27545) );
  XOR U28083 ( .A(n27547), .B(n27548), .Z(n18216) );
  XOR U28084 ( .A(n27549), .B(n27550), .Z(n27543) );
  AND U28085 ( .A(n27551), .B(n27552), .Z(n27550) );
  XOR U28086 ( .A(e_input[531]), .B(n27549), .Z(n27552) );
  XNOR U28087 ( .A(n18228), .B(n27549), .Z(n27551) );
  XOR U28088 ( .A(n27553), .B(n27554), .Z(n18228) );
  XOR U28089 ( .A(n27555), .B(n27556), .Z(n27549) );
  AND U28090 ( .A(n27557), .B(n27558), .Z(n27556) );
  XOR U28091 ( .A(e_input[530]), .B(n27555), .Z(n27558) );
  XNOR U28092 ( .A(n18240), .B(n27555), .Z(n27557) );
  XOR U28093 ( .A(n27559), .B(n27560), .Z(n18240) );
  XOR U28094 ( .A(n27561), .B(n27562), .Z(n27555) );
  AND U28095 ( .A(n27563), .B(n27564), .Z(n27562) );
  XOR U28096 ( .A(e_input[529]), .B(n27561), .Z(n27564) );
  XNOR U28097 ( .A(n18252), .B(n27561), .Z(n27563) );
  XOR U28098 ( .A(n27565), .B(n27566), .Z(n18252) );
  XOR U28099 ( .A(n27567), .B(n27568), .Z(n27561) );
  AND U28100 ( .A(n27569), .B(n27570), .Z(n27568) );
  XOR U28101 ( .A(e_input[528]), .B(n27567), .Z(n27570) );
  XNOR U28102 ( .A(n18264), .B(n27567), .Z(n27569) );
  XOR U28103 ( .A(n27571), .B(n27572), .Z(n18264) );
  XOR U28104 ( .A(n27573), .B(n27574), .Z(n27567) );
  AND U28105 ( .A(n27575), .B(n27576), .Z(n27574) );
  XOR U28106 ( .A(e_input[527]), .B(n27573), .Z(n27576) );
  XNOR U28107 ( .A(n18276), .B(n27573), .Z(n27575) );
  XOR U28108 ( .A(n27577), .B(n27578), .Z(n18276) );
  XOR U28109 ( .A(n27579), .B(n27580), .Z(n27573) );
  AND U28110 ( .A(n27581), .B(n27582), .Z(n27580) );
  XOR U28111 ( .A(e_input[526]), .B(n27579), .Z(n27582) );
  XNOR U28112 ( .A(n18288), .B(n27579), .Z(n27581) );
  XOR U28113 ( .A(n27583), .B(n27584), .Z(n18288) );
  XOR U28114 ( .A(n27585), .B(n27586), .Z(n27579) );
  AND U28115 ( .A(n27587), .B(n27588), .Z(n27586) );
  XOR U28116 ( .A(e_input[525]), .B(n27585), .Z(n27588) );
  XNOR U28117 ( .A(n18300), .B(n27585), .Z(n27587) );
  XOR U28118 ( .A(n27589), .B(n27590), .Z(n18300) );
  XOR U28119 ( .A(n27591), .B(n27592), .Z(n27585) );
  AND U28120 ( .A(n27593), .B(n27594), .Z(n27592) );
  XOR U28121 ( .A(e_input[524]), .B(n27591), .Z(n27594) );
  XNOR U28122 ( .A(n18312), .B(n27591), .Z(n27593) );
  XOR U28123 ( .A(n27595), .B(n27596), .Z(n18312) );
  XOR U28124 ( .A(n27597), .B(n27598), .Z(n27591) );
  AND U28125 ( .A(n27599), .B(n27600), .Z(n27598) );
  XOR U28126 ( .A(e_input[523]), .B(n27597), .Z(n27600) );
  XNOR U28127 ( .A(n18324), .B(n27597), .Z(n27599) );
  XOR U28128 ( .A(n27601), .B(n27602), .Z(n18324) );
  XOR U28129 ( .A(n27603), .B(n27604), .Z(n27597) );
  AND U28130 ( .A(n27605), .B(n27606), .Z(n27604) );
  XOR U28131 ( .A(e_input[522]), .B(n27603), .Z(n27606) );
  XNOR U28132 ( .A(n18336), .B(n27603), .Z(n27605) );
  XOR U28133 ( .A(n27607), .B(n27608), .Z(n18336) );
  XOR U28134 ( .A(n27609), .B(n27610), .Z(n27603) );
  AND U28135 ( .A(n27611), .B(n27612), .Z(n27610) );
  XOR U28136 ( .A(e_input[521]), .B(n27609), .Z(n27612) );
  XNOR U28137 ( .A(n18348), .B(n27609), .Z(n27611) );
  XOR U28138 ( .A(n27613), .B(n27614), .Z(n18348) );
  XOR U28139 ( .A(n27615), .B(n27616), .Z(n27609) );
  AND U28140 ( .A(n27617), .B(n27618), .Z(n27616) );
  XOR U28141 ( .A(e_input[520]), .B(n27615), .Z(n27618) );
  XNOR U28142 ( .A(n18360), .B(n27615), .Z(n27617) );
  XOR U28143 ( .A(n27619), .B(n27620), .Z(n18360) );
  XOR U28144 ( .A(n27621), .B(n27622), .Z(n27615) );
  AND U28145 ( .A(n27623), .B(n27624), .Z(n27622) );
  XOR U28146 ( .A(e_input[519]), .B(n27621), .Z(n27624) );
  XNOR U28147 ( .A(n18372), .B(n27621), .Z(n27623) );
  XOR U28148 ( .A(n27625), .B(n27626), .Z(n18372) );
  XOR U28149 ( .A(n27627), .B(n27628), .Z(n27621) );
  AND U28150 ( .A(n27629), .B(n27630), .Z(n27628) );
  XOR U28151 ( .A(e_input[518]), .B(n27627), .Z(n27630) );
  XNOR U28152 ( .A(n18384), .B(n27627), .Z(n27629) );
  XOR U28153 ( .A(n27631), .B(n27632), .Z(n18384) );
  XOR U28154 ( .A(n27633), .B(n27634), .Z(n27627) );
  AND U28155 ( .A(n27635), .B(n27636), .Z(n27634) );
  XOR U28156 ( .A(e_input[517]), .B(n27633), .Z(n27636) );
  XNOR U28157 ( .A(n18396), .B(n27633), .Z(n27635) );
  XOR U28158 ( .A(n27637), .B(n27638), .Z(n18396) );
  XOR U28159 ( .A(n27639), .B(n27640), .Z(n27633) );
  AND U28160 ( .A(n27641), .B(n27642), .Z(n27640) );
  XOR U28161 ( .A(e_input[516]), .B(n27639), .Z(n27642) );
  XNOR U28162 ( .A(n18408), .B(n27639), .Z(n27641) );
  XOR U28163 ( .A(n27643), .B(n27644), .Z(n18408) );
  XOR U28164 ( .A(n27645), .B(n27646), .Z(n27639) );
  AND U28165 ( .A(n27647), .B(n27648), .Z(n27646) );
  XOR U28166 ( .A(e_input[515]), .B(n27645), .Z(n27648) );
  XNOR U28167 ( .A(n18420), .B(n27645), .Z(n27647) );
  XOR U28168 ( .A(n27649), .B(n27650), .Z(n18420) );
  XOR U28169 ( .A(n27651), .B(n27652), .Z(n27645) );
  AND U28170 ( .A(n27653), .B(n27654), .Z(n27652) );
  XOR U28171 ( .A(e_input[514]), .B(n27651), .Z(n27654) );
  XNOR U28172 ( .A(n18432), .B(n27651), .Z(n27653) );
  XOR U28173 ( .A(n27655), .B(n27656), .Z(n18432) );
  XOR U28174 ( .A(n27657), .B(n27658), .Z(n27651) );
  AND U28175 ( .A(n27659), .B(n27660), .Z(n27658) );
  XOR U28176 ( .A(e_input[513]), .B(n27657), .Z(n27660) );
  XNOR U28177 ( .A(n18444), .B(n27657), .Z(n27659) );
  XOR U28178 ( .A(n27661), .B(n27662), .Z(n18444) );
  XOR U28179 ( .A(n27663), .B(n27664), .Z(n27657) );
  AND U28180 ( .A(n27665), .B(n27666), .Z(n27664) );
  XOR U28181 ( .A(e_input[512]), .B(n27663), .Z(n27666) );
  XNOR U28182 ( .A(n18456), .B(n27663), .Z(n27665) );
  XOR U28183 ( .A(n27667), .B(n27668), .Z(n18456) );
  XOR U28184 ( .A(n27669), .B(n27670), .Z(n27663) );
  AND U28185 ( .A(n27671), .B(n27672), .Z(n27670) );
  XOR U28186 ( .A(e_input[511]), .B(n27669), .Z(n27672) );
  XNOR U28187 ( .A(n18468), .B(n27669), .Z(n27671) );
  XOR U28188 ( .A(n27673), .B(n27674), .Z(n18468) );
  XOR U28189 ( .A(n27675), .B(n27676), .Z(n27669) );
  AND U28190 ( .A(n27677), .B(n27678), .Z(n27676) );
  XOR U28191 ( .A(e_input[510]), .B(n27675), .Z(n27678) );
  XNOR U28192 ( .A(n18480), .B(n27675), .Z(n27677) );
  XOR U28193 ( .A(n27679), .B(n27680), .Z(n18480) );
  XOR U28194 ( .A(n27681), .B(n27682), .Z(n27675) );
  AND U28195 ( .A(n27683), .B(n27684), .Z(n27682) );
  XOR U28196 ( .A(e_input[509]), .B(n27681), .Z(n27684) );
  XNOR U28197 ( .A(n18492), .B(n27681), .Z(n27683) );
  XOR U28198 ( .A(n27685), .B(n27686), .Z(n18492) );
  XOR U28199 ( .A(n27687), .B(n27688), .Z(n27681) );
  AND U28200 ( .A(n27689), .B(n27690), .Z(n27688) );
  XOR U28201 ( .A(e_input[508]), .B(n27687), .Z(n27690) );
  XNOR U28202 ( .A(n18504), .B(n27687), .Z(n27689) );
  XOR U28203 ( .A(n27691), .B(n27692), .Z(n18504) );
  XOR U28204 ( .A(n27693), .B(n27694), .Z(n27687) );
  AND U28205 ( .A(n27695), .B(n27696), .Z(n27694) );
  XOR U28206 ( .A(e_input[507]), .B(n27693), .Z(n27696) );
  XNOR U28207 ( .A(n18516), .B(n27693), .Z(n27695) );
  XOR U28208 ( .A(n27697), .B(n27698), .Z(n18516) );
  XOR U28209 ( .A(n27699), .B(n27700), .Z(n27693) );
  AND U28210 ( .A(n27701), .B(n27702), .Z(n27700) );
  XOR U28211 ( .A(e_input[506]), .B(n27699), .Z(n27702) );
  XNOR U28212 ( .A(n18528), .B(n27699), .Z(n27701) );
  XOR U28213 ( .A(n27703), .B(n27704), .Z(n18528) );
  XOR U28214 ( .A(n27705), .B(n27706), .Z(n27699) );
  AND U28215 ( .A(n27707), .B(n27708), .Z(n27706) );
  XOR U28216 ( .A(e_input[505]), .B(n27705), .Z(n27708) );
  XNOR U28217 ( .A(n18540), .B(n27705), .Z(n27707) );
  XOR U28218 ( .A(n27709), .B(n27710), .Z(n18540) );
  XOR U28219 ( .A(n27711), .B(n27712), .Z(n27705) );
  AND U28220 ( .A(n27713), .B(n27714), .Z(n27712) );
  XOR U28221 ( .A(e_input[504]), .B(n27711), .Z(n27714) );
  XNOR U28222 ( .A(n18552), .B(n27711), .Z(n27713) );
  XOR U28223 ( .A(n27715), .B(n27716), .Z(n18552) );
  XOR U28224 ( .A(n27717), .B(n27718), .Z(n27711) );
  AND U28225 ( .A(n27719), .B(n27720), .Z(n27718) );
  XOR U28226 ( .A(e_input[503]), .B(n27717), .Z(n27720) );
  XNOR U28227 ( .A(n18564), .B(n27717), .Z(n27719) );
  XOR U28228 ( .A(n27721), .B(n27722), .Z(n18564) );
  XOR U28229 ( .A(n27723), .B(n27724), .Z(n27717) );
  AND U28230 ( .A(n27725), .B(n27726), .Z(n27724) );
  XOR U28231 ( .A(e_input[502]), .B(n27723), .Z(n27726) );
  XNOR U28232 ( .A(n18576), .B(n27723), .Z(n27725) );
  XOR U28233 ( .A(n27727), .B(n27728), .Z(n18576) );
  XOR U28234 ( .A(n27729), .B(n27730), .Z(n27723) );
  AND U28235 ( .A(n27731), .B(n27732), .Z(n27730) );
  XOR U28236 ( .A(e_input[501]), .B(n27729), .Z(n27732) );
  XNOR U28237 ( .A(n18588), .B(n27729), .Z(n27731) );
  XOR U28238 ( .A(n27733), .B(n27734), .Z(n18588) );
  XOR U28239 ( .A(n27735), .B(n27736), .Z(n27729) );
  AND U28240 ( .A(n27737), .B(n27738), .Z(n27736) );
  XOR U28241 ( .A(e_input[500]), .B(n27735), .Z(n27738) );
  XNOR U28242 ( .A(n18600), .B(n27735), .Z(n27737) );
  XOR U28243 ( .A(n27739), .B(n27740), .Z(n18600) );
  XOR U28244 ( .A(n27741), .B(n27742), .Z(n27735) );
  AND U28245 ( .A(n27743), .B(n27744), .Z(n27742) );
  XOR U28246 ( .A(e_input[499]), .B(n27741), .Z(n27744) );
  XNOR U28247 ( .A(n18612), .B(n27741), .Z(n27743) );
  XOR U28248 ( .A(n27745), .B(n27746), .Z(n18612) );
  XOR U28249 ( .A(n27747), .B(n27748), .Z(n27741) );
  AND U28250 ( .A(n27749), .B(n27750), .Z(n27748) );
  XOR U28251 ( .A(e_input[498]), .B(n27747), .Z(n27750) );
  XNOR U28252 ( .A(n18624), .B(n27747), .Z(n27749) );
  XOR U28253 ( .A(n27751), .B(n27752), .Z(n18624) );
  XOR U28254 ( .A(n27753), .B(n27754), .Z(n27747) );
  AND U28255 ( .A(n27755), .B(n27756), .Z(n27754) );
  XOR U28256 ( .A(e_input[497]), .B(n27753), .Z(n27756) );
  XNOR U28257 ( .A(n18636), .B(n27753), .Z(n27755) );
  XOR U28258 ( .A(n27757), .B(n27758), .Z(n18636) );
  XOR U28259 ( .A(n27759), .B(n27760), .Z(n27753) );
  AND U28260 ( .A(n27761), .B(n27762), .Z(n27760) );
  XOR U28261 ( .A(e_input[496]), .B(n27759), .Z(n27762) );
  XNOR U28262 ( .A(n18648), .B(n27759), .Z(n27761) );
  XOR U28263 ( .A(n27763), .B(n27764), .Z(n18648) );
  XOR U28264 ( .A(n27765), .B(n27766), .Z(n27759) );
  AND U28265 ( .A(n27767), .B(n27768), .Z(n27766) );
  XOR U28266 ( .A(e_input[495]), .B(n27765), .Z(n27768) );
  XNOR U28267 ( .A(n18660), .B(n27765), .Z(n27767) );
  XOR U28268 ( .A(n27769), .B(n27770), .Z(n18660) );
  XOR U28269 ( .A(n27771), .B(n27772), .Z(n27765) );
  AND U28270 ( .A(n27773), .B(n27774), .Z(n27772) );
  XOR U28271 ( .A(e_input[494]), .B(n27771), .Z(n27774) );
  XNOR U28272 ( .A(n18672), .B(n27771), .Z(n27773) );
  XOR U28273 ( .A(n27775), .B(n27776), .Z(n18672) );
  XOR U28274 ( .A(n27777), .B(n27778), .Z(n27771) );
  AND U28275 ( .A(n27779), .B(n27780), .Z(n27778) );
  XOR U28276 ( .A(e_input[493]), .B(n27777), .Z(n27780) );
  XNOR U28277 ( .A(n18684), .B(n27777), .Z(n27779) );
  XOR U28278 ( .A(n27781), .B(n27782), .Z(n18684) );
  XOR U28279 ( .A(n27783), .B(n27784), .Z(n27777) );
  AND U28280 ( .A(n27785), .B(n27786), .Z(n27784) );
  XOR U28281 ( .A(e_input[492]), .B(n27783), .Z(n27786) );
  XNOR U28282 ( .A(n18696), .B(n27783), .Z(n27785) );
  XOR U28283 ( .A(n27787), .B(n27788), .Z(n18696) );
  XOR U28284 ( .A(n27789), .B(n27790), .Z(n27783) );
  AND U28285 ( .A(n27791), .B(n27792), .Z(n27790) );
  XOR U28286 ( .A(e_input[491]), .B(n27789), .Z(n27792) );
  XNOR U28287 ( .A(n18708), .B(n27789), .Z(n27791) );
  XOR U28288 ( .A(n27793), .B(n27794), .Z(n18708) );
  XOR U28289 ( .A(n27795), .B(n27796), .Z(n27789) );
  AND U28290 ( .A(n27797), .B(n27798), .Z(n27796) );
  XOR U28291 ( .A(e_input[490]), .B(n27795), .Z(n27798) );
  XNOR U28292 ( .A(n18720), .B(n27795), .Z(n27797) );
  XOR U28293 ( .A(n27799), .B(n27800), .Z(n18720) );
  XOR U28294 ( .A(n27801), .B(n27802), .Z(n27795) );
  AND U28295 ( .A(n27803), .B(n27804), .Z(n27802) );
  XOR U28296 ( .A(e_input[489]), .B(n27801), .Z(n27804) );
  XNOR U28297 ( .A(n18732), .B(n27801), .Z(n27803) );
  XOR U28298 ( .A(n27805), .B(n27806), .Z(n18732) );
  XOR U28299 ( .A(n27807), .B(n27808), .Z(n27801) );
  AND U28300 ( .A(n27809), .B(n27810), .Z(n27808) );
  XOR U28301 ( .A(e_input[488]), .B(n27807), .Z(n27810) );
  XNOR U28302 ( .A(n18744), .B(n27807), .Z(n27809) );
  XOR U28303 ( .A(n27811), .B(n27812), .Z(n18744) );
  XOR U28304 ( .A(n27813), .B(n27814), .Z(n27807) );
  AND U28305 ( .A(n27815), .B(n27816), .Z(n27814) );
  XOR U28306 ( .A(e_input[487]), .B(n27813), .Z(n27816) );
  XNOR U28307 ( .A(n18756), .B(n27813), .Z(n27815) );
  XOR U28308 ( .A(n27817), .B(n27818), .Z(n18756) );
  XOR U28309 ( .A(n27819), .B(n27820), .Z(n27813) );
  AND U28310 ( .A(n27821), .B(n27822), .Z(n27820) );
  XOR U28311 ( .A(e_input[486]), .B(n27819), .Z(n27822) );
  XNOR U28312 ( .A(n18768), .B(n27819), .Z(n27821) );
  XOR U28313 ( .A(n27823), .B(n27824), .Z(n18768) );
  XOR U28314 ( .A(n27825), .B(n27826), .Z(n27819) );
  AND U28315 ( .A(n27827), .B(n27828), .Z(n27826) );
  XOR U28316 ( .A(e_input[485]), .B(n27825), .Z(n27828) );
  XNOR U28317 ( .A(n18780), .B(n27825), .Z(n27827) );
  XOR U28318 ( .A(n27829), .B(n27830), .Z(n18780) );
  XOR U28319 ( .A(n27831), .B(n27832), .Z(n27825) );
  AND U28320 ( .A(n27833), .B(n27834), .Z(n27832) );
  XOR U28321 ( .A(e_input[484]), .B(n27831), .Z(n27834) );
  XNOR U28322 ( .A(n18792), .B(n27831), .Z(n27833) );
  XOR U28323 ( .A(n27835), .B(n27836), .Z(n18792) );
  XOR U28324 ( .A(n27837), .B(n27838), .Z(n27831) );
  AND U28325 ( .A(n27839), .B(n27840), .Z(n27838) );
  XOR U28326 ( .A(e_input[483]), .B(n27837), .Z(n27840) );
  XNOR U28327 ( .A(n18804), .B(n27837), .Z(n27839) );
  XOR U28328 ( .A(n27841), .B(n27842), .Z(n18804) );
  XOR U28329 ( .A(n27843), .B(n27844), .Z(n27837) );
  AND U28330 ( .A(n27845), .B(n27846), .Z(n27844) );
  XOR U28331 ( .A(e_input[482]), .B(n27843), .Z(n27846) );
  XNOR U28332 ( .A(n18816), .B(n27843), .Z(n27845) );
  XOR U28333 ( .A(n27847), .B(n27848), .Z(n18816) );
  XOR U28334 ( .A(n27849), .B(n27850), .Z(n27843) );
  AND U28335 ( .A(n27851), .B(n27852), .Z(n27850) );
  XOR U28336 ( .A(e_input[481]), .B(n27849), .Z(n27852) );
  XNOR U28337 ( .A(n18828), .B(n27849), .Z(n27851) );
  XOR U28338 ( .A(n27853), .B(n27854), .Z(n18828) );
  XOR U28339 ( .A(n27855), .B(n27856), .Z(n27849) );
  AND U28340 ( .A(n27857), .B(n27858), .Z(n27856) );
  XOR U28341 ( .A(e_input[480]), .B(n27855), .Z(n27858) );
  XNOR U28342 ( .A(n18840), .B(n27855), .Z(n27857) );
  XOR U28343 ( .A(n27859), .B(n27860), .Z(n18840) );
  XOR U28344 ( .A(n27861), .B(n27862), .Z(n27855) );
  AND U28345 ( .A(n27863), .B(n27864), .Z(n27862) );
  XOR U28346 ( .A(e_input[479]), .B(n27861), .Z(n27864) );
  XNOR U28347 ( .A(n18852), .B(n27861), .Z(n27863) );
  XOR U28348 ( .A(n27865), .B(n27866), .Z(n18852) );
  XOR U28349 ( .A(n27867), .B(n27868), .Z(n27861) );
  AND U28350 ( .A(n27869), .B(n27870), .Z(n27868) );
  XOR U28351 ( .A(e_input[478]), .B(n27867), .Z(n27870) );
  XNOR U28352 ( .A(n18864), .B(n27867), .Z(n27869) );
  XOR U28353 ( .A(n27871), .B(n27872), .Z(n18864) );
  XOR U28354 ( .A(n27873), .B(n27874), .Z(n27867) );
  AND U28355 ( .A(n27875), .B(n27876), .Z(n27874) );
  XOR U28356 ( .A(e_input[477]), .B(n27873), .Z(n27876) );
  XNOR U28357 ( .A(n18876), .B(n27873), .Z(n27875) );
  XOR U28358 ( .A(n27877), .B(n27878), .Z(n18876) );
  XOR U28359 ( .A(n27879), .B(n27880), .Z(n27873) );
  AND U28360 ( .A(n27881), .B(n27882), .Z(n27880) );
  XOR U28361 ( .A(e_input[476]), .B(n27879), .Z(n27882) );
  XNOR U28362 ( .A(n18888), .B(n27879), .Z(n27881) );
  XOR U28363 ( .A(n27883), .B(n27884), .Z(n18888) );
  XOR U28364 ( .A(n27885), .B(n27886), .Z(n27879) );
  AND U28365 ( .A(n27887), .B(n27888), .Z(n27886) );
  XOR U28366 ( .A(e_input[475]), .B(n27885), .Z(n27888) );
  XNOR U28367 ( .A(n18900), .B(n27885), .Z(n27887) );
  XOR U28368 ( .A(n27889), .B(n27890), .Z(n18900) );
  XOR U28369 ( .A(n27891), .B(n27892), .Z(n27885) );
  AND U28370 ( .A(n27893), .B(n27894), .Z(n27892) );
  XOR U28371 ( .A(e_input[474]), .B(n27891), .Z(n27894) );
  XNOR U28372 ( .A(n18912), .B(n27891), .Z(n27893) );
  XOR U28373 ( .A(n27895), .B(n27896), .Z(n18912) );
  XOR U28374 ( .A(n27897), .B(n27898), .Z(n27891) );
  AND U28375 ( .A(n27899), .B(n27900), .Z(n27898) );
  XOR U28376 ( .A(e_input[473]), .B(n27897), .Z(n27900) );
  XNOR U28377 ( .A(n18924), .B(n27897), .Z(n27899) );
  XOR U28378 ( .A(n27901), .B(n27902), .Z(n18924) );
  XOR U28379 ( .A(n27903), .B(n27904), .Z(n27897) );
  AND U28380 ( .A(n27905), .B(n27906), .Z(n27904) );
  XOR U28381 ( .A(e_input[472]), .B(n27903), .Z(n27906) );
  XNOR U28382 ( .A(n18936), .B(n27903), .Z(n27905) );
  XOR U28383 ( .A(n27907), .B(n27908), .Z(n18936) );
  XOR U28384 ( .A(n27909), .B(n27910), .Z(n27903) );
  AND U28385 ( .A(n27911), .B(n27912), .Z(n27910) );
  XOR U28386 ( .A(e_input[471]), .B(n27909), .Z(n27912) );
  XNOR U28387 ( .A(n18948), .B(n27909), .Z(n27911) );
  XOR U28388 ( .A(n27913), .B(n27914), .Z(n18948) );
  XOR U28389 ( .A(n27915), .B(n27916), .Z(n27909) );
  AND U28390 ( .A(n27917), .B(n27918), .Z(n27916) );
  XOR U28391 ( .A(e_input[470]), .B(n27915), .Z(n27918) );
  XNOR U28392 ( .A(n18960), .B(n27915), .Z(n27917) );
  XOR U28393 ( .A(n27919), .B(n27920), .Z(n18960) );
  XOR U28394 ( .A(n27921), .B(n27922), .Z(n27915) );
  AND U28395 ( .A(n27923), .B(n27924), .Z(n27922) );
  XOR U28396 ( .A(e_input[469]), .B(n27921), .Z(n27924) );
  XNOR U28397 ( .A(n18972), .B(n27921), .Z(n27923) );
  XOR U28398 ( .A(n27925), .B(n27926), .Z(n18972) );
  XOR U28399 ( .A(n27927), .B(n27928), .Z(n27921) );
  AND U28400 ( .A(n27929), .B(n27930), .Z(n27928) );
  XOR U28401 ( .A(e_input[468]), .B(n27927), .Z(n27930) );
  XNOR U28402 ( .A(n18984), .B(n27927), .Z(n27929) );
  XOR U28403 ( .A(n27931), .B(n27932), .Z(n18984) );
  XOR U28404 ( .A(n27933), .B(n27934), .Z(n27927) );
  AND U28405 ( .A(n27935), .B(n27936), .Z(n27934) );
  XOR U28406 ( .A(e_input[467]), .B(n27933), .Z(n27936) );
  XNOR U28407 ( .A(n18996), .B(n27933), .Z(n27935) );
  XOR U28408 ( .A(n27937), .B(n27938), .Z(n18996) );
  XOR U28409 ( .A(n27939), .B(n27940), .Z(n27933) );
  AND U28410 ( .A(n27941), .B(n27942), .Z(n27940) );
  XOR U28411 ( .A(e_input[466]), .B(n27939), .Z(n27942) );
  XNOR U28412 ( .A(n19008), .B(n27939), .Z(n27941) );
  XOR U28413 ( .A(n27943), .B(n27944), .Z(n19008) );
  XOR U28414 ( .A(n27945), .B(n27946), .Z(n27939) );
  AND U28415 ( .A(n27947), .B(n27948), .Z(n27946) );
  XOR U28416 ( .A(e_input[465]), .B(n27945), .Z(n27948) );
  XNOR U28417 ( .A(n19020), .B(n27945), .Z(n27947) );
  XOR U28418 ( .A(n27949), .B(n27950), .Z(n19020) );
  XOR U28419 ( .A(n27951), .B(n27952), .Z(n27945) );
  AND U28420 ( .A(n27953), .B(n27954), .Z(n27952) );
  XOR U28421 ( .A(e_input[464]), .B(n27951), .Z(n27954) );
  XNOR U28422 ( .A(n19032), .B(n27951), .Z(n27953) );
  XOR U28423 ( .A(n27955), .B(n27956), .Z(n19032) );
  XOR U28424 ( .A(n27957), .B(n27958), .Z(n27951) );
  AND U28425 ( .A(n27959), .B(n27960), .Z(n27958) );
  XOR U28426 ( .A(e_input[463]), .B(n27957), .Z(n27960) );
  XNOR U28427 ( .A(n19044), .B(n27957), .Z(n27959) );
  XOR U28428 ( .A(n27961), .B(n27962), .Z(n19044) );
  XOR U28429 ( .A(n27963), .B(n27964), .Z(n27957) );
  AND U28430 ( .A(n27965), .B(n27966), .Z(n27964) );
  XOR U28431 ( .A(e_input[462]), .B(n27963), .Z(n27966) );
  XNOR U28432 ( .A(n19056), .B(n27963), .Z(n27965) );
  XOR U28433 ( .A(n27967), .B(n27968), .Z(n19056) );
  XOR U28434 ( .A(n27969), .B(n27970), .Z(n27963) );
  AND U28435 ( .A(n27971), .B(n27972), .Z(n27970) );
  XOR U28436 ( .A(e_input[461]), .B(n27969), .Z(n27972) );
  XNOR U28437 ( .A(n19068), .B(n27969), .Z(n27971) );
  XOR U28438 ( .A(n27973), .B(n27974), .Z(n19068) );
  XOR U28439 ( .A(n27975), .B(n27976), .Z(n27969) );
  AND U28440 ( .A(n27977), .B(n27978), .Z(n27976) );
  XOR U28441 ( .A(e_input[460]), .B(n27975), .Z(n27978) );
  XNOR U28442 ( .A(n19080), .B(n27975), .Z(n27977) );
  XOR U28443 ( .A(n27979), .B(n27980), .Z(n19080) );
  XOR U28444 ( .A(n27981), .B(n27982), .Z(n27975) );
  AND U28445 ( .A(n27983), .B(n27984), .Z(n27982) );
  XOR U28446 ( .A(e_input[459]), .B(n27981), .Z(n27984) );
  XNOR U28447 ( .A(n19092), .B(n27981), .Z(n27983) );
  XOR U28448 ( .A(n27985), .B(n27986), .Z(n19092) );
  XOR U28449 ( .A(n27987), .B(n27988), .Z(n27981) );
  AND U28450 ( .A(n27989), .B(n27990), .Z(n27988) );
  XOR U28451 ( .A(e_input[458]), .B(n27987), .Z(n27990) );
  XNOR U28452 ( .A(n19104), .B(n27987), .Z(n27989) );
  XOR U28453 ( .A(n27991), .B(n27992), .Z(n19104) );
  XOR U28454 ( .A(n27993), .B(n27994), .Z(n27987) );
  AND U28455 ( .A(n27995), .B(n27996), .Z(n27994) );
  XOR U28456 ( .A(e_input[457]), .B(n27993), .Z(n27996) );
  XNOR U28457 ( .A(n19116), .B(n27993), .Z(n27995) );
  XOR U28458 ( .A(n27997), .B(n27998), .Z(n19116) );
  XOR U28459 ( .A(n27999), .B(n28000), .Z(n27993) );
  AND U28460 ( .A(n28001), .B(n28002), .Z(n28000) );
  XOR U28461 ( .A(e_input[456]), .B(n27999), .Z(n28002) );
  XNOR U28462 ( .A(n19128), .B(n27999), .Z(n28001) );
  XOR U28463 ( .A(n28003), .B(n28004), .Z(n19128) );
  XOR U28464 ( .A(n28005), .B(n28006), .Z(n27999) );
  AND U28465 ( .A(n28007), .B(n28008), .Z(n28006) );
  XOR U28466 ( .A(e_input[455]), .B(n28005), .Z(n28008) );
  XNOR U28467 ( .A(n19140), .B(n28005), .Z(n28007) );
  XOR U28468 ( .A(n28009), .B(n28010), .Z(n19140) );
  XOR U28469 ( .A(n28011), .B(n28012), .Z(n28005) );
  AND U28470 ( .A(n28013), .B(n28014), .Z(n28012) );
  XOR U28471 ( .A(e_input[454]), .B(n28011), .Z(n28014) );
  XNOR U28472 ( .A(n19152), .B(n28011), .Z(n28013) );
  XOR U28473 ( .A(n28015), .B(n28016), .Z(n19152) );
  XOR U28474 ( .A(n28017), .B(n28018), .Z(n28011) );
  AND U28475 ( .A(n28019), .B(n28020), .Z(n28018) );
  XOR U28476 ( .A(e_input[453]), .B(n28017), .Z(n28020) );
  XNOR U28477 ( .A(n19164), .B(n28017), .Z(n28019) );
  XOR U28478 ( .A(n28021), .B(n28022), .Z(n19164) );
  XOR U28479 ( .A(n28023), .B(n28024), .Z(n28017) );
  AND U28480 ( .A(n28025), .B(n28026), .Z(n28024) );
  XOR U28481 ( .A(e_input[452]), .B(n28023), .Z(n28026) );
  XNOR U28482 ( .A(n19176), .B(n28023), .Z(n28025) );
  XOR U28483 ( .A(n28027), .B(n28028), .Z(n19176) );
  XOR U28484 ( .A(n28029), .B(n28030), .Z(n28023) );
  AND U28485 ( .A(n28031), .B(n28032), .Z(n28030) );
  XOR U28486 ( .A(e_input[451]), .B(n28029), .Z(n28032) );
  XNOR U28487 ( .A(n19188), .B(n28029), .Z(n28031) );
  XOR U28488 ( .A(n28033), .B(n28034), .Z(n19188) );
  XOR U28489 ( .A(n28035), .B(n28036), .Z(n28029) );
  AND U28490 ( .A(n28037), .B(n28038), .Z(n28036) );
  XOR U28491 ( .A(e_input[450]), .B(n28035), .Z(n28038) );
  XNOR U28492 ( .A(n19200), .B(n28035), .Z(n28037) );
  XOR U28493 ( .A(n28039), .B(n28040), .Z(n19200) );
  XOR U28494 ( .A(n28041), .B(n28042), .Z(n28035) );
  AND U28495 ( .A(n28043), .B(n28044), .Z(n28042) );
  XOR U28496 ( .A(e_input[449]), .B(n28041), .Z(n28044) );
  XNOR U28497 ( .A(n19212), .B(n28041), .Z(n28043) );
  XOR U28498 ( .A(n28045), .B(n28046), .Z(n19212) );
  XOR U28499 ( .A(n28047), .B(n28048), .Z(n28041) );
  AND U28500 ( .A(n28049), .B(n28050), .Z(n28048) );
  XOR U28501 ( .A(e_input[448]), .B(n28047), .Z(n28050) );
  XNOR U28502 ( .A(n19224), .B(n28047), .Z(n28049) );
  XOR U28503 ( .A(n28051), .B(n28052), .Z(n19224) );
  XOR U28504 ( .A(n28053), .B(n28054), .Z(n28047) );
  AND U28505 ( .A(n28055), .B(n28056), .Z(n28054) );
  XOR U28506 ( .A(e_input[447]), .B(n28053), .Z(n28056) );
  XNOR U28507 ( .A(n19236), .B(n28053), .Z(n28055) );
  XOR U28508 ( .A(n28057), .B(n28058), .Z(n19236) );
  XOR U28509 ( .A(n28059), .B(n28060), .Z(n28053) );
  AND U28510 ( .A(n28061), .B(n28062), .Z(n28060) );
  XOR U28511 ( .A(e_input[446]), .B(n28059), .Z(n28062) );
  XNOR U28512 ( .A(n19248), .B(n28059), .Z(n28061) );
  XOR U28513 ( .A(n28063), .B(n28064), .Z(n19248) );
  XOR U28514 ( .A(n28065), .B(n28066), .Z(n28059) );
  AND U28515 ( .A(n28067), .B(n28068), .Z(n28066) );
  XOR U28516 ( .A(e_input[445]), .B(n28065), .Z(n28068) );
  XNOR U28517 ( .A(n19260), .B(n28065), .Z(n28067) );
  XOR U28518 ( .A(n28069), .B(n28070), .Z(n19260) );
  XOR U28519 ( .A(n28071), .B(n28072), .Z(n28065) );
  AND U28520 ( .A(n28073), .B(n28074), .Z(n28072) );
  XOR U28521 ( .A(e_input[444]), .B(n28071), .Z(n28074) );
  XNOR U28522 ( .A(n19272), .B(n28071), .Z(n28073) );
  XOR U28523 ( .A(n28075), .B(n28076), .Z(n19272) );
  XOR U28524 ( .A(n28077), .B(n28078), .Z(n28071) );
  AND U28525 ( .A(n28079), .B(n28080), .Z(n28078) );
  XOR U28526 ( .A(e_input[443]), .B(n28077), .Z(n28080) );
  XNOR U28527 ( .A(n19284), .B(n28077), .Z(n28079) );
  XOR U28528 ( .A(n28081), .B(n28082), .Z(n19284) );
  XOR U28529 ( .A(n28083), .B(n28084), .Z(n28077) );
  AND U28530 ( .A(n28085), .B(n28086), .Z(n28084) );
  XOR U28531 ( .A(e_input[442]), .B(n28083), .Z(n28086) );
  XNOR U28532 ( .A(n19296), .B(n28083), .Z(n28085) );
  XOR U28533 ( .A(n28087), .B(n28088), .Z(n19296) );
  XOR U28534 ( .A(n28089), .B(n28090), .Z(n28083) );
  AND U28535 ( .A(n28091), .B(n28092), .Z(n28090) );
  XOR U28536 ( .A(e_input[441]), .B(n28089), .Z(n28092) );
  XNOR U28537 ( .A(n19308), .B(n28089), .Z(n28091) );
  XOR U28538 ( .A(n28093), .B(n28094), .Z(n19308) );
  XOR U28539 ( .A(n28095), .B(n28096), .Z(n28089) );
  AND U28540 ( .A(n28097), .B(n28098), .Z(n28096) );
  XOR U28541 ( .A(e_input[440]), .B(n28095), .Z(n28098) );
  XNOR U28542 ( .A(n19320), .B(n28095), .Z(n28097) );
  XOR U28543 ( .A(n28099), .B(n28100), .Z(n19320) );
  XOR U28544 ( .A(n28101), .B(n28102), .Z(n28095) );
  AND U28545 ( .A(n28103), .B(n28104), .Z(n28102) );
  XOR U28546 ( .A(e_input[439]), .B(n28101), .Z(n28104) );
  XNOR U28547 ( .A(n19332), .B(n28101), .Z(n28103) );
  XOR U28548 ( .A(n28105), .B(n28106), .Z(n19332) );
  XOR U28549 ( .A(n28107), .B(n28108), .Z(n28101) );
  AND U28550 ( .A(n28109), .B(n28110), .Z(n28108) );
  XOR U28551 ( .A(e_input[438]), .B(n28107), .Z(n28110) );
  XNOR U28552 ( .A(n19344), .B(n28107), .Z(n28109) );
  XOR U28553 ( .A(n28111), .B(n28112), .Z(n19344) );
  XOR U28554 ( .A(n28113), .B(n28114), .Z(n28107) );
  AND U28555 ( .A(n28115), .B(n28116), .Z(n28114) );
  XOR U28556 ( .A(e_input[437]), .B(n28113), .Z(n28116) );
  XNOR U28557 ( .A(n19356), .B(n28113), .Z(n28115) );
  XOR U28558 ( .A(n28117), .B(n28118), .Z(n19356) );
  XOR U28559 ( .A(n28119), .B(n28120), .Z(n28113) );
  AND U28560 ( .A(n28121), .B(n28122), .Z(n28120) );
  XOR U28561 ( .A(e_input[436]), .B(n28119), .Z(n28122) );
  XNOR U28562 ( .A(n19368), .B(n28119), .Z(n28121) );
  XOR U28563 ( .A(n28123), .B(n28124), .Z(n19368) );
  XOR U28564 ( .A(n28125), .B(n28126), .Z(n28119) );
  AND U28565 ( .A(n28127), .B(n28128), .Z(n28126) );
  XOR U28566 ( .A(e_input[435]), .B(n28125), .Z(n28128) );
  XNOR U28567 ( .A(n19380), .B(n28125), .Z(n28127) );
  XOR U28568 ( .A(n28129), .B(n28130), .Z(n19380) );
  XOR U28569 ( .A(n28131), .B(n28132), .Z(n28125) );
  AND U28570 ( .A(n28133), .B(n28134), .Z(n28132) );
  XOR U28571 ( .A(e_input[434]), .B(n28131), .Z(n28134) );
  XNOR U28572 ( .A(n19392), .B(n28131), .Z(n28133) );
  XOR U28573 ( .A(n28135), .B(n28136), .Z(n19392) );
  XOR U28574 ( .A(n28137), .B(n28138), .Z(n28131) );
  AND U28575 ( .A(n28139), .B(n28140), .Z(n28138) );
  XOR U28576 ( .A(e_input[433]), .B(n28137), .Z(n28140) );
  XNOR U28577 ( .A(n19404), .B(n28137), .Z(n28139) );
  XOR U28578 ( .A(n28141), .B(n28142), .Z(n19404) );
  XOR U28579 ( .A(n28143), .B(n28144), .Z(n28137) );
  AND U28580 ( .A(n28145), .B(n28146), .Z(n28144) );
  XOR U28581 ( .A(e_input[432]), .B(n28143), .Z(n28146) );
  XNOR U28582 ( .A(n19416), .B(n28143), .Z(n28145) );
  XOR U28583 ( .A(n28147), .B(n28148), .Z(n19416) );
  XOR U28584 ( .A(n28149), .B(n28150), .Z(n28143) );
  AND U28585 ( .A(n28151), .B(n28152), .Z(n28150) );
  XOR U28586 ( .A(e_input[431]), .B(n28149), .Z(n28152) );
  XNOR U28587 ( .A(n19428), .B(n28149), .Z(n28151) );
  XOR U28588 ( .A(n28153), .B(n28154), .Z(n19428) );
  XOR U28589 ( .A(n28155), .B(n28156), .Z(n28149) );
  AND U28590 ( .A(n28157), .B(n28158), .Z(n28156) );
  XOR U28591 ( .A(e_input[430]), .B(n28155), .Z(n28158) );
  XNOR U28592 ( .A(n19440), .B(n28155), .Z(n28157) );
  XOR U28593 ( .A(n28159), .B(n28160), .Z(n19440) );
  XOR U28594 ( .A(n28161), .B(n28162), .Z(n28155) );
  AND U28595 ( .A(n28163), .B(n28164), .Z(n28162) );
  XOR U28596 ( .A(e_input[429]), .B(n28161), .Z(n28164) );
  XNOR U28597 ( .A(n19452), .B(n28161), .Z(n28163) );
  XOR U28598 ( .A(n28165), .B(n28166), .Z(n19452) );
  XOR U28599 ( .A(n28167), .B(n28168), .Z(n28161) );
  AND U28600 ( .A(n28169), .B(n28170), .Z(n28168) );
  XOR U28601 ( .A(e_input[428]), .B(n28167), .Z(n28170) );
  XNOR U28602 ( .A(n19464), .B(n28167), .Z(n28169) );
  XOR U28603 ( .A(n28171), .B(n28172), .Z(n19464) );
  XOR U28604 ( .A(n28173), .B(n28174), .Z(n28167) );
  AND U28605 ( .A(n28175), .B(n28176), .Z(n28174) );
  XOR U28606 ( .A(e_input[427]), .B(n28173), .Z(n28176) );
  XNOR U28607 ( .A(n19476), .B(n28173), .Z(n28175) );
  XOR U28608 ( .A(n28177), .B(n28178), .Z(n19476) );
  XOR U28609 ( .A(n28179), .B(n28180), .Z(n28173) );
  AND U28610 ( .A(n28181), .B(n28182), .Z(n28180) );
  XOR U28611 ( .A(e_input[426]), .B(n28179), .Z(n28182) );
  XNOR U28612 ( .A(n19488), .B(n28179), .Z(n28181) );
  XOR U28613 ( .A(n28183), .B(n28184), .Z(n19488) );
  XOR U28614 ( .A(n28185), .B(n28186), .Z(n28179) );
  AND U28615 ( .A(n28187), .B(n28188), .Z(n28186) );
  XOR U28616 ( .A(e_input[425]), .B(n28185), .Z(n28188) );
  XNOR U28617 ( .A(n19500), .B(n28185), .Z(n28187) );
  XOR U28618 ( .A(n28189), .B(n28190), .Z(n19500) );
  XOR U28619 ( .A(n28191), .B(n28192), .Z(n28185) );
  AND U28620 ( .A(n28193), .B(n28194), .Z(n28192) );
  XOR U28621 ( .A(e_input[424]), .B(n28191), .Z(n28194) );
  XNOR U28622 ( .A(n19512), .B(n28191), .Z(n28193) );
  XOR U28623 ( .A(n28195), .B(n28196), .Z(n19512) );
  XOR U28624 ( .A(n28197), .B(n28198), .Z(n28191) );
  AND U28625 ( .A(n28199), .B(n28200), .Z(n28198) );
  XOR U28626 ( .A(e_input[423]), .B(n28197), .Z(n28200) );
  XNOR U28627 ( .A(n19524), .B(n28197), .Z(n28199) );
  XOR U28628 ( .A(n28201), .B(n28202), .Z(n19524) );
  XOR U28629 ( .A(n28203), .B(n28204), .Z(n28197) );
  AND U28630 ( .A(n28205), .B(n28206), .Z(n28204) );
  XOR U28631 ( .A(e_input[422]), .B(n28203), .Z(n28206) );
  XNOR U28632 ( .A(n19536), .B(n28203), .Z(n28205) );
  XOR U28633 ( .A(n28207), .B(n28208), .Z(n19536) );
  XOR U28634 ( .A(n28209), .B(n28210), .Z(n28203) );
  AND U28635 ( .A(n28211), .B(n28212), .Z(n28210) );
  XOR U28636 ( .A(e_input[421]), .B(n28209), .Z(n28212) );
  XNOR U28637 ( .A(n19548), .B(n28209), .Z(n28211) );
  XOR U28638 ( .A(n28213), .B(n28214), .Z(n19548) );
  XOR U28639 ( .A(n28215), .B(n28216), .Z(n28209) );
  AND U28640 ( .A(n28217), .B(n28218), .Z(n28216) );
  XOR U28641 ( .A(e_input[420]), .B(n28215), .Z(n28218) );
  XNOR U28642 ( .A(n19560), .B(n28215), .Z(n28217) );
  XOR U28643 ( .A(n28219), .B(n28220), .Z(n19560) );
  XOR U28644 ( .A(n28221), .B(n28222), .Z(n28215) );
  AND U28645 ( .A(n28223), .B(n28224), .Z(n28222) );
  XOR U28646 ( .A(e_input[419]), .B(n28221), .Z(n28224) );
  XNOR U28647 ( .A(n19572), .B(n28221), .Z(n28223) );
  XOR U28648 ( .A(n28225), .B(n28226), .Z(n19572) );
  XOR U28649 ( .A(n28227), .B(n28228), .Z(n28221) );
  AND U28650 ( .A(n28229), .B(n28230), .Z(n28228) );
  XOR U28651 ( .A(e_input[418]), .B(n28227), .Z(n28230) );
  XNOR U28652 ( .A(n19584), .B(n28227), .Z(n28229) );
  XOR U28653 ( .A(n28231), .B(n28232), .Z(n19584) );
  XOR U28654 ( .A(n28233), .B(n28234), .Z(n28227) );
  AND U28655 ( .A(n28235), .B(n28236), .Z(n28234) );
  XOR U28656 ( .A(e_input[417]), .B(n28233), .Z(n28236) );
  XNOR U28657 ( .A(n19596), .B(n28233), .Z(n28235) );
  XOR U28658 ( .A(n28237), .B(n28238), .Z(n19596) );
  XOR U28659 ( .A(n28239), .B(n28240), .Z(n28233) );
  AND U28660 ( .A(n28241), .B(n28242), .Z(n28240) );
  XOR U28661 ( .A(e_input[416]), .B(n28239), .Z(n28242) );
  XNOR U28662 ( .A(n19608), .B(n28239), .Z(n28241) );
  XOR U28663 ( .A(n28243), .B(n28244), .Z(n19608) );
  XOR U28664 ( .A(n28245), .B(n28246), .Z(n28239) );
  AND U28665 ( .A(n28247), .B(n28248), .Z(n28246) );
  XOR U28666 ( .A(e_input[415]), .B(n28245), .Z(n28248) );
  XNOR U28667 ( .A(n19620), .B(n28245), .Z(n28247) );
  XOR U28668 ( .A(n28249), .B(n28250), .Z(n19620) );
  XOR U28669 ( .A(n28251), .B(n28252), .Z(n28245) );
  AND U28670 ( .A(n28253), .B(n28254), .Z(n28252) );
  XOR U28671 ( .A(e_input[414]), .B(n28251), .Z(n28254) );
  XNOR U28672 ( .A(n19632), .B(n28251), .Z(n28253) );
  XOR U28673 ( .A(n28255), .B(n28256), .Z(n19632) );
  XOR U28674 ( .A(n28257), .B(n28258), .Z(n28251) );
  AND U28675 ( .A(n28259), .B(n28260), .Z(n28258) );
  XOR U28676 ( .A(e_input[413]), .B(n28257), .Z(n28260) );
  XNOR U28677 ( .A(n19644), .B(n28257), .Z(n28259) );
  XOR U28678 ( .A(n28261), .B(n28262), .Z(n19644) );
  XOR U28679 ( .A(n28263), .B(n28264), .Z(n28257) );
  AND U28680 ( .A(n28265), .B(n28266), .Z(n28264) );
  XOR U28681 ( .A(e_input[412]), .B(n28263), .Z(n28266) );
  XNOR U28682 ( .A(n19656), .B(n28263), .Z(n28265) );
  XOR U28683 ( .A(n28267), .B(n28268), .Z(n19656) );
  XOR U28684 ( .A(n28269), .B(n28270), .Z(n28263) );
  AND U28685 ( .A(n28271), .B(n28272), .Z(n28270) );
  XOR U28686 ( .A(e_input[411]), .B(n28269), .Z(n28272) );
  XNOR U28687 ( .A(n19668), .B(n28269), .Z(n28271) );
  XOR U28688 ( .A(n28273), .B(n28274), .Z(n19668) );
  XOR U28689 ( .A(n28275), .B(n28276), .Z(n28269) );
  AND U28690 ( .A(n28277), .B(n28278), .Z(n28276) );
  XOR U28691 ( .A(e_input[410]), .B(n28275), .Z(n28278) );
  XNOR U28692 ( .A(n19680), .B(n28275), .Z(n28277) );
  XOR U28693 ( .A(n28279), .B(n28280), .Z(n19680) );
  XOR U28694 ( .A(n28281), .B(n28282), .Z(n28275) );
  AND U28695 ( .A(n28283), .B(n28284), .Z(n28282) );
  XOR U28696 ( .A(e_input[409]), .B(n28281), .Z(n28284) );
  XNOR U28697 ( .A(n19692), .B(n28281), .Z(n28283) );
  XOR U28698 ( .A(n28285), .B(n28286), .Z(n19692) );
  XOR U28699 ( .A(n28287), .B(n28288), .Z(n28281) );
  AND U28700 ( .A(n28289), .B(n28290), .Z(n28288) );
  XOR U28701 ( .A(e_input[408]), .B(n28287), .Z(n28290) );
  XNOR U28702 ( .A(n19704), .B(n28287), .Z(n28289) );
  XOR U28703 ( .A(n28291), .B(n28292), .Z(n19704) );
  XOR U28704 ( .A(n28293), .B(n28294), .Z(n28287) );
  AND U28705 ( .A(n28295), .B(n28296), .Z(n28294) );
  XOR U28706 ( .A(e_input[407]), .B(n28293), .Z(n28296) );
  XNOR U28707 ( .A(n19716), .B(n28293), .Z(n28295) );
  XOR U28708 ( .A(n28297), .B(n28298), .Z(n19716) );
  XOR U28709 ( .A(n28299), .B(n28300), .Z(n28293) );
  AND U28710 ( .A(n28301), .B(n28302), .Z(n28300) );
  XOR U28711 ( .A(e_input[406]), .B(n28299), .Z(n28302) );
  XNOR U28712 ( .A(n19728), .B(n28299), .Z(n28301) );
  XOR U28713 ( .A(n28303), .B(n28304), .Z(n19728) );
  XOR U28714 ( .A(n28305), .B(n28306), .Z(n28299) );
  AND U28715 ( .A(n28307), .B(n28308), .Z(n28306) );
  XOR U28716 ( .A(e_input[405]), .B(n28305), .Z(n28308) );
  XNOR U28717 ( .A(n19740), .B(n28305), .Z(n28307) );
  XOR U28718 ( .A(n28309), .B(n28310), .Z(n19740) );
  XOR U28719 ( .A(n28311), .B(n28312), .Z(n28305) );
  AND U28720 ( .A(n28313), .B(n28314), .Z(n28312) );
  XOR U28721 ( .A(e_input[404]), .B(n28311), .Z(n28314) );
  XNOR U28722 ( .A(n19752), .B(n28311), .Z(n28313) );
  XOR U28723 ( .A(n28315), .B(n28316), .Z(n19752) );
  XOR U28724 ( .A(n28317), .B(n28318), .Z(n28311) );
  AND U28725 ( .A(n28319), .B(n28320), .Z(n28318) );
  XOR U28726 ( .A(e_input[403]), .B(n28317), .Z(n28320) );
  XNOR U28727 ( .A(n19764), .B(n28317), .Z(n28319) );
  XOR U28728 ( .A(n28321), .B(n28322), .Z(n19764) );
  XOR U28729 ( .A(n28323), .B(n28324), .Z(n28317) );
  AND U28730 ( .A(n28325), .B(n28326), .Z(n28324) );
  XOR U28731 ( .A(e_input[402]), .B(n28323), .Z(n28326) );
  XNOR U28732 ( .A(n19776), .B(n28323), .Z(n28325) );
  XOR U28733 ( .A(n28327), .B(n28328), .Z(n19776) );
  XOR U28734 ( .A(n28329), .B(n28330), .Z(n28323) );
  AND U28735 ( .A(n28331), .B(n28332), .Z(n28330) );
  XOR U28736 ( .A(e_input[401]), .B(n28329), .Z(n28332) );
  XNOR U28737 ( .A(n19788), .B(n28329), .Z(n28331) );
  XOR U28738 ( .A(n28333), .B(n28334), .Z(n19788) );
  XOR U28739 ( .A(n28335), .B(n28336), .Z(n28329) );
  AND U28740 ( .A(n28337), .B(n28338), .Z(n28336) );
  XOR U28741 ( .A(e_input[400]), .B(n28335), .Z(n28338) );
  XNOR U28742 ( .A(n19800), .B(n28335), .Z(n28337) );
  XOR U28743 ( .A(n28339), .B(n28340), .Z(n19800) );
  XOR U28744 ( .A(n28341), .B(n28342), .Z(n28335) );
  AND U28745 ( .A(n28343), .B(n28344), .Z(n28342) );
  XOR U28746 ( .A(e_input[399]), .B(n28341), .Z(n28344) );
  XNOR U28747 ( .A(n19812), .B(n28341), .Z(n28343) );
  XOR U28748 ( .A(n28345), .B(n28346), .Z(n19812) );
  XOR U28749 ( .A(n28347), .B(n28348), .Z(n28341) );
  AND U28750 ( .A(n28349), .B(n28350), .Z(n28348) );
  XOR U28751 ( .A(e_input[398]), .B(n28347), .Z(n28350) );
  XNOR U28752 ( .A(n19824), .B(n28347), .Z(n28349) );
  XOR U28753 ( .A(n28351), .B(n28352), .Z(n19824) );
  XOR U28754 ( .A(n28353), .B(n28354), .Z(n28347) );
  AND U28755 ( .A(n28355), .B(n28356), .Z(n28354) );
  XOR U28756 ( .A(e_input[397]), .B(n28353), .Z(n28356) );
  XNOR U28757 ( .A(n19836), .B(n28353), .Z(n28355) );
  XOR U28758 ( .A(n28357), .B(n28358), .Z(n19836) );
  XOR U28759 ( .A(n28359), .B(n28360), .Z(n28353) );
  AND U28760 ( .A(n28361), .B(n28362), .Z(n28360) );
  XOR U28761 ( .A(e_input[396]), .B(n28359), .Z(n28362) );
  XNOR U28762 ( .A(n19848), .B(n28359), .Z(n28361) );
  XOR U28763 ( .A(n28363), .B(n28364), .Z(n19848) );
  XOR U28764 ( .A(n28365), .B(n28366), .Z(n28359) );
  AND U28765 ( .A(n28367), .B(n28368), .Z(n28366) );
  XOR U28766 ( .A(e_input[395]), .B(n28365), .Z(n28368) );
  XNOR U28767 ( .A(n19860), .B(n28365), .Z(n28367) );
  XOR U28768 ( .A(n28369), .B(n28370), .Z(n19860) );
  XOR U28769 ( .A(n28371), .B(n28372), .Z(n28365) );
  AND U28770 ( .A(n28373), .B(n28374), .Z(n28372) );
  XOR U28771 ( .A(e_input[394]), .B(n28371), .Z(n28374) );
  XNOR U28772 ( .A(n19872), .B(n28371), .Z(n28373) );
  XOR U28773 ( .A(n28375), .B(n28376), .Z(n19872) );
  XOR U28774 ( .A(n28377), .B(n28378), .Z(n28371) );
  AND U28775 ( .A(n28379), .B(n28380), .Z(n28378) );
  XOR U28776 ( .A(e_input[393]), .B(n28377), .Z(n28380) );
  XNOR U28777 ( .A(n19884), .B(n28377), .Z(n28379) );
  XOR U28778 ( .A(n28381), .B(n28382), .Z(n19884) );
  XOR U28779 ( .A(n28383), .B(n28384), .Z(n28377) );
  AND U28780 ( .A(n28385), .B(n28386), .Z(n28384) );
  XOR U28781 ( .A(e_input[392]), .B(n28383), .Z(n28386) );
  XNOR U28782 ( .A(n19896), .B(n28383), .Z(n28385) );
  XOR U28783 ( .A(n28387), .B(n28388), .Z(n19896) );
  XOR U28784 ( .A(n28389), .B(n28390), .Z(n28383) );
  AND U28785 ( .A(n28391), .B(n28392), .Z(n28390) );
  XOR U28786 ( .A(e_input[391]), .B(n28389), .Z(n28392) );
  XNOR U28787 ( .A(n19908), .B(n28389), .Z(n28391) );
  XOR U28788 ( .A(n28393), .B(n28394), .Z(n19908) );
  XOR U28789 ( .A(n28395), .B(n28396), .Z(n28389) );
  AND U28790 ( .A(n28397), .B(n28398), .Z(n28396) );
  XOR U28791 ( .A(e_input[390]), .B(n28395), .Z(n28398) );
  XNOR U28792 ( .A(n19920), .B(n28395), .Z(n28397) );
  XOR U28793 ( .A(n28399), .B(n28400), .Z(n19920) );
  XOR U28794 ( .A(n28401), .B(n28402), .Z(n28395) );
  AND U28795 ( .A(n28403), .B(n28404), .Z(n28402) );
  XOR U28796 ( .A(e_input[389]), .B(n28401), .Z(n28404) );
  XNOR U28797 ( .A(n19932), .B(n28401), .Z(n28403) );
  XOR U28798 ( .A(n28405), .B(n28406), .Z(n19932) );
  XOR U28799 ( .A(n28407), .B(n28408), .Z(n28401) );
  AND U28800 ( .A(n28409), .B(n28410), .Z(n28408) );
  XOR U28801 ( .A(e_input[388]), .B(n28407), .Z(n28410) );
  XNOR U28802 ( .A(n19944), .B(n28407), .Z(n28409) );
  XOR U28803 ( .A(n28411), .B(n28412), .Z(n19944) );
  XOR U28804 ( .A(n28413), .B(n28414), .Z(n28407) );
  AND U28805 ( .A(n28415), .B(n28416), .Z(n28414) );
  XOR U28806 ( .A(e_input[387]), .B(n28413), .Z(n28416) );
  XNOR U28807 ( .A(n19956), .B(n28413), .Z(n28415) );
  XOR U28808 ( .A(n28417), .B(n28418), .Z(n19956) );
  XOR U28809 ( .A(n28419), .B(n28420), .Z(n28413) );
  AND U28810 ( .A(n28421), .B(n28422), .Z(n28420) );
  XOR U28811 ( .A(e_input[386]), .B(n28419), .Z(n28422) );
  XNOR U28812 ( .A(n19968), .B(n28419), .Z(n28421) );
  XOR U28813 ( .A(n28423), .B(n28424), .Z(n19968) );
  XOR U28814 ( .A(n28425), .B(n28426), .Z(n28419) );
  AND U28815 ( .A(n28427), .B(n28428), .Z(n28426) );
  XOR U28816 ( .A(e_input[385]), .B(n28425), .Z(n28428) );
  XNOR U28817 ( .A(n19980), .B(n28425), .Z(n28427) );
  XOR U28818 ( .A(n28429), .B(n28430), .Z(n19980) );
  XOR U28819 ( .A(n28431), .B(n28432), .Z(n28425) );
  AND U28820 ( .A(n28433), .B(n28434), .Z(n28432) );
  XOR U28821 ( .A(e_input[384]), .B(n28431), .Z(n28434) );
  XNOR U28822 ( .A(n19992), .B(n28431), .Z(n28433) );
  XOR U28823 ( .A(n28435), .B(n28436), .Z(n19992) );
  XOR U28824 ( .A(n28437), .B(n28438), .Z(n28431) );
  AND U28825 ( .A(n28439), .B(n28440), .Z(n28438) );
  XOR U28826 ( .A(e_input[383]), .B(n28437), .Z(n28440) );
  XNOR U28827 ( .A(n20004), .B(n28437), .Z(n28439) );
  XOR U28828 ( .A(n28441), .B(n28442), .Z(n20004) );
  XOR U28829 ( .A(n28443), .B(n28444), .Z(n28437) );
  AND U28830 ( .A(n28445), .B(n28446), .Z(n28444) );
  XOR U28831 ( .A(e_input[382]), .B(n28443), .Z(n28446) );
  XNOR U28832 ( .A(n20016), .B(n28443), .Z(n28445) );
  XOR U28833 ( .A(n28447), .B(n28448), .Z(n20016) );
  XOR U28834 ( .A(n28449), .B(n28450), .Z(n28443) );
  AND U28835 ( .A(n28451), .B(n28452), .Z(n28450) );
  XOR U28836 ( .A(e_input[381]), .B(n28449), .Z(n28452) );
  XNOR U28837 ( .A(n20028), .B(n28449), .Z(n28451) );
  XOR U28838 ( .A(n28453), .B(n28454), .Z(n20028) );
  XOR U28839 ( .A(n28455), .B(n28456), .Z(n28449) );
  AND U28840 ( .A(n28457), .B(n28458), .Z(n28456) );
  XOR U28841 ( .A(e_input[380]), .B(n28455), .Z(n28458) );
  XNOR U28842 ( .A(n20040), .B(n28455), .Z(n28457) );
  XOR U28843 ( .A(n28459), .B(n28460), .Z(n20040) );
  XOR U28844 ( .A(n28461), .B(n28462), .Z(n28455) );
  AND U28845 ( .A(n28463), .B(n28464), .Z(n28462) );
  XOR U28846 ( .A(e_input[379]), .B(n28461), .Z(n28464) );
  XNOR U28847 ( .A(n20052), .B(n28461), .Z(n28463) );
  XOR U28848 ( .A(n28465), .B(n28466), .Z(n20052) );
  XOR U28849 ( .A(n28467), .B(n28468), .Z(n28461) );
  AND U28850 ( .A(n28469), .B(n28470), .Z(n28468) );
  XOR U28851 ( .A(e_input[378]), .B(n28467), .Z(n28470) );
  XNOR U28852 ( .A(n20064), .B(n28467), .Z(n28469) );
  XOR U28853 ( .A(n28471), .B(n28472), .Z(n20064) );
  XOR U28854 ( .A(n28473), .B(n28474), .Z(n28467) );
  AND U28855 ( .A(n28475), .B(n28476), .Z(n28474) );
  XOR U28856 ( .A(e_input[377]), .B(n28473), .Z(n28476) );
  XNOR U28857 ( .A(n20076), .B(n28473), .Z(n28475) );
  XOR U28858 ( .A(n28477), .B(n28478), .Z(n20076) );
  XOR U28859 ( .A(n28479), .B(n28480), .Z(n28473) );
  AND U28860 ( .A(n28481), .B(n28482), .Z(n28480) );
  XOR U28861 ( .A(e_input[376]), .B(n28479), .Z(n28482) );
  XNOR U28862 ( .A(n20088), .B(n28479), .Z(n28481) );
  XOR U28863 ( .A(n28483), .B(n28484), .Z(n20088) );
  XOR U28864 ( .A(n28485), .B(n28486), .Z(n28479) );
  AND U28865 ( .A(n28487), .B(n28488), .Z(n28486) );
  XOR U28866 ( .A(e_input[375]), .B(n28485), .Z(n28488) );
  XNOR U28867 ( .A(n20100), .B(n28485), .Z(n28487) );
  XOR U28868 ( .A(n28489), .B(n28490), .Z(n20100) );
  XOR U28869 ( .A(n28491), .B(n28492), .Z(n28485) );
  AND U28870 ( .A(n28493), .B(n28494), .Z(n28492) );
  XOR U28871 ( .A(e_input[374]), .B(n28491), .Z(n28494) );
  XNOR U28872 ( .A(n20112), .B(n28491), .Z(n28493) );
  XOR U28873 ( .A(n28495), .B(n28496), .Z(n20112) );
  XOR U28874 ( .A(n28497), .B(n28498), .Z(n28491) );
  AND U28875 ( .A(n28499), .B(n28500), .Z(n28498) );
  XOR U28876 ( .A(e_input[373]), .B(n28497), .Z(n28500) );
  XNOR U28877 ( .A(n20124), .B(n28497), .Z(n28499) );
  XOR U28878 ( .A(n28501), .B(n28502), .Z(n20124) );
  XOR U28879 ( .A(n28503), .B(n28504), .Z(n28497) );
  AND U28880 ( .A(n28505), .B(n28506), .Z(n28504) );
  XOR U28881 ( .A(e_input[372]), .B(n28503), .Z(n28506) );
  XNOR U28882 ( .A(n20136), .B(n28503), .Z(n28505) );
  XOR U28883 ( .A(n28507), .B(n28508), .Z(n20136) );
  XOR U28884 ( .A(n28509), .B(n28510), .Z(n28503) );
  AND U28885 ( .A(n28511), .B(n28512), .Z(n28510) );
  XOR U28886 ( .A(e_input[371]), .B(n28509), .Z(n28512) );
  XNOR U28887 ( .A(n20148), .B(n28509), .Z(n28511) );
  XOR U28888 ( .A(n28513), .B(n28514), .Z(n20148) );
  XOR U28889 ( .A(n28515), .B(n28516), .Z(n28509) );
  AND U28890 ( .A(n28517), .B(n28518), .Z(n28516) );
  XOR U28891 ( .A(e_input[370]), .B(n28515), .Z(n28518) );
  XNOR U28892 ( .A(n20160), .B(n28515), .Z(n28517) );
  XOR U28893 ( .A(n28519), .B(n28520), .Z(n20160) );
  XOR U28894 ( .A(n28521), .B(n28522), .Z(n28515) );
  AND U28895 ( .A(n28523), .B(n28524), .Z(n28522) );
  XOR U28896 ( .A(e_input[369]), .B(n28521), .Z(n28524) );
  XNOR U28897 ( .A(n20172), .B(n28521), .Z(n28523) );
  XOR U28898 ( .A(n28525), .B(n28526), .Z(n20172) );
  XOR U28899 ( .A(n28527), .B(n28528), .Z(n28521) );
  AND U28900 ( .A(n28529), .B(n28530), .Z(n28528) );
  XOR U28901 ( .A(e_input[368]), .B(n28527), .Z(n28530) );
  XNOR U28902 ( .A(n20184), .B(n28527), .Z(n28529) );
  XOR U28903 ( .A(n28531), .B(n28532), .Z(n20184) );
  XOR U28904 ( .A(n28533), .B(n28534), .Z(n28527) );
  AND U28905 ( .A(n28535), .B(n28536), .Z(n28534) );
  XOR U28906 ( .A(e_input[367]), .B(n28533), .Z(n28536) );
  XNOR U28907 ( .A(n20196), .B(n28533), .Z(n28535) );
  XOR U28908 ( .A(n28537), .B(n28538), .Z(n20196) );
  XOR U28909 ( .A(n28539), .B(n28540), .Z(n28533) );
  AND U28910 ( .A(n28541), .B(n28542), .Z(n28540) );
  XOR U28911 ( .A(e_input[366]), .B(n28539), .Z(n28542) );
  XNOR U28912 ( .A(n20208), .B(n28539), .Z(n28541) );
  XOR U28913 ( .A(n28543), .B(n28544), .Z(n20208) );
  XOR U28914 ( .A(n28545), .B(n28546), .Z(n28539) );
  AND U28915 ( .A(n28547), .B(n28548), .Z(n28546) );
  XOR U28916 ( .A(e_input[365]), .B(n28545), .Z(n28548) );
  XNOR U28917 ( .A(n20220), .B(n28545), .Z(n28547) );
  XOR U28918 ( .A(n28549), .B(n28550), .Z(n20220) );
  XOR U28919 ( .A(n28551), .B(n28552), .Z(n28545) );
  AND U28920 ( .A(n28553), .B(n28554), .Z(n28552) );
  XOR U28921 ( .A(e_input[364]), .B(n28551), .Z(n28554) );
  XNOR U28922 ( .A(n20232), .B(n28551), .Z(n28553) );
  XOR U28923 ( .A(n28555), .B(n28556), .Z(n20232) );
  XOR U28924 ( .A(n28557), .B(n28558), .Z(n28551) );
  AND U28925 ( .A(n28559), .B(n28560), .Z(n28558) );
  XOR U28926 ( .A(e_input[363]), .B(n28557), .Z(n28560) );
  XNOR U28927 ( .A(n20244), .B(n28557), .Z(n28559) );
  XOR U28928 ( .A(n28561), .B(n28562), .Z(n20244) );
  XOR U28929 ( .A(n28563), .B(n28564), .Z(n28557) );
  AND U28930 ( .A(n28565), .B(n28566), .Z(n28564) );
  XOR U28931 ( .A(e_input[362]), .B(n28563), .Z(n28566) );
  XNOR U28932 ( .A(n20256), .B(n28563), .Z(n28565) );
  XOR U28933 ( .A(n28567), .B(n28568), .Z(n20256) );
  XOR U28934 ( .A(n28569), .B(n28570), .Z(n28563) );
  AND U28935 ( .A(n28571), .B(n28572), .Z(n28570) );
  XOR U28936 ( .A(e_input[361]), .B(n28569), .Z(n28572) );
  XNOR U28937 ( .A(n20268), .B(n28569), .Z(n28571) );
  XOR U28938 ( .A(n28573), .B(n28574), .Z(n20268) );
  XOR U28939 ( .A(n28575), .B(n28576), .Z(n28569) );
  AND U28940 ( .A(n28577), .B(n28578), .Z(n28576) );
  XOR U28941 ( .A(e_input[360]), .B(n28575), .Z(n28578) );
  XNOR U28942 ( .A(n20280), .B(n28575), .Z(n28577) );
  XOR U28943 ( .A(n28579), .B(n28580), .Z(n20280) );
  XOR U28944 ( .A(n28581), .B(n28582), .Z(n28575) );
  AND U28945 ( .A(n28583), .B(n28584), .Z(n28582) );
  XOR U28946 ( .A(e_input[359]), .B(n28581), .Z(n28584) );
  XNOR U28947 ( .A(n20292), .B(n28581), .Z(n28583) );
  XOR U28948 ( .A(n28585), .B(n28586), .Z(n20292) );
  XOR U28949 ( .A(n28587), .B(n28588), .Z(n28581) );
  AND U28950 ( .A(n28589), .B(n28590), .Z(n28588) );
  XOR U28951 ( .A(e_input[358]), .B(n28587), .Z(n28590) );
  XNOR U28952 ( .A(n20304), .B(n28587), .Z(n28589) );
  XOR U28953 ( .A(n28591), .B(n28592), .Z(n20304) );
  XOR U28954 ( .A(n28593), .B(n28594), .Z(n28587) );
  AND U28955 ( .A(n28595), .B(n28596), .Z(n28594) );
  XOR U28956 ( .A(e_input[357]), .B(n28593), .Z(n28596) );
  XNOR U28957 ( .A(n20316), .B(n28593), .Z(n28595) );
  XOR U28958 ( .A(n28597), .B(n28598), .Z(n20316) );
  XOR U28959 ( .A(n28599), .B(n28600), .Z(n28593) );
  AND U28960 ( .A(n28601), .B(n28602), .Z(n28600) );
  XOR U28961 ( .A(e_input[356]), .B(n28599), .Z(n28602) );
  XNOR U28962 ( .A(n20328), .B(n28599), .Z(n28601) );
  XOR U28963 ( .A(n28603), .B(n28604), .Z(n20328) );
  XOR U28964 ( .A(n28605), .B(n28606), .Z(n28599) );
  AND U28965 ( .A(n28607), .B(n28608), .Z(n28606) );
  XOR U28966 ( .A(e_input[355]), .B(n28605), .Z(n28608) );
  XNOR U28967 ( .A(n20340), .B(n28605), .Z(n28607) );
  XOR U28968 ( .A(n28609), .B(n28610), .Z(n20340) );
  XOR U28969 ( .A(n28611), .B(n28612), .Z(n28605) );
  AND U28970 ( .A(n28613), .B(n28614), .Z(n28612) );
  XOR U28971 ( .A(e_input[354]), .B(n28611), .Z(n28614) );
  XNOR U28972 ( .A(n20352), .B(n28611), .Z(n28613) );
  XOR U28973 ( .A(n28615), .B(n28616), .Z(n20352) );
  XOR U28974 ( .A(n28617), .B(n28618), .Z(n28611) );
  AND U28975 ( .A(n28619), .B(n28620), .Z(n28618) );
  XOR U28976 ( .A(e_input[353]), .B(n28617), .Z(n28620) );
  XNOR U28977 ( .A(n20364), .B(n28617), .Z(n28619) );
  XOR U28978 ( .A(n28621), .B(n28622), .Z(n20364) );
  XOR U28979 ( .A(n28623), .B(n28624), .Z(n28617) );
  AND U28980 ( .A(n28625), .B(n28626), .Z(n28624) );
  XOR U28981 ( .A(e_input[352]), .B(n28623), .Z(n28626) );
  XNOR U28982 ( .A(n20376), .B(n28623), .Z(n28625) );
  XOR U28983 ( .A(n28627), .B(n28628), .Z(n20376) );
  XOR U28984 ( .A(n28629), .B(n28630), .Z(n28623) );
  AND U28985 ( .A(n28631), .B(n28632), .Z(n28630) );
  XOR U28986 ( .A(e_input[351]), .B(n28629), .Z(n28632) );
  XNOR U28987 ( .A(n20388), .B(n28629), .Z(n28631) );
  XOR U28988 ( .A(n28633), .B(n28634), .Z(n20388) );
  XOR U28989 ( .A(n28635), .B(n28636), .Z(n28629) );
  AND U28990 ( .A(n28637), .B(n28638), .Z(n28636) );
  XOR U28991 ( .A(e_input[350]), .B(n28635), .Z(n28638) );
  XNOR U28992 ( .A(n20400), .B(n28635), .Z(n28637) );
  XOR U28993 ( .A(n28639), .B(n28640), .Z(n20400) );
  XOR U28994 ( .A(n28641), .B(n28642), .Z(n28635) );
  AND U28995 ( .A(n28643), .B(n28644), .Z(n28642) );
  XOR U28996 ( .A(e_input[349]), .B(n28641), .Z(n28644) );
  XNOR U28997 ( .A(n20412), .B(n28641), .Z(n28643) );
  XOR U28998 ( .A(n28645), .B(n28646), .Z(n20412) );
  XOR U28999 ( .A(n28647), .B(n28648), .Z(n28641) );
  AND U29000 ( .A(n28649), .B(n28650), .Z(n28648) );
  XOR U29001 ( .A(e_input[348]), .B(n28647), .Z(n28650) );
  XNOR U29002 ( .A(n20424), .B(n28647), .Z(n28649) );
  XOR U29003 ( .A(n28651), .B(n28652), .Z(n20424) );
  XOR U29004 ( .A(n28653), .B(n28654), .Z(n28647) );
  AND U29005 ( .A(n28655), .B(n28656), .Z(n28654) );
  XOR U29006 ( .A(e_input[347]), .B(n28653), .Z(n28656) );
  XNOR U29007 ( .A(n20436), .B(n28653), .Z(n28655) );
  XOR U29008 ( .A(n28657), .B(n28658), .Z(n20436) );
  XOR U29009 ( .A(n28659), .B(n28660), .Z(n28653) );
  AND U29010 ( .A(n28661), .B(n28662), .Z(n28660) );
  XOR U29011 ( .A(e_input[346]), .B(n28659), .Z(n28662) );
  XNOR U29012 ( .A(n20448), .B(n28659), .Z(n28661) );
  XOR U29013 ( .A(n28663), .B(n28664), .Z(n20448) );
  XOR U29014 ( .A(n28665), .B(n28666), .Z(n28659) );
  AND U29015 ( .A(n28667), .B(n28668), .Z(n28666) );
  XOR U29016 ( .A(e_input[345]), .B(n28665), .Z(n28668) );
  XNOR U29017 ( .A(n20460), .B(n28665), .Z(n28667) );
  XOR U29018 ( .A(n28669), .B(n28670), .Z(n20460) );
  XOR U29019 ( .A(n28671), .B(n28672), .Z(n28665) );
  AND U29020 ( .A(n28673), .B(n28674), .Z(n28672) );
  XOR U29021 ( .A(e_input[344]), .B(n28671), .Z(n28674) );
  XNOR U29022 ( .A(n20472), .B(n28671), .Z(n28673) );
  XOR U29023 ( .A(n28675), .B(n28676), .Z(n20472) );
  XOR U29024 ( .A(n28677), .B(n28678), .Z(n28671) );
  AND U29025 ( .A(n28679), .B(n28680), .Z(n28678) );
  XOR U29026 ( .A(e_input[343]), .B(n28677), .Z(n28680) );
  XNOR U29027 ( .A(n20484), .B(n28677), .Z(n28679) );
  XOR U29028 ( .A(n28681), .B(n28682), .Z(n20484) );
  XOR U29029 ( .A(n28683), .B(n28684), .Z(n28677) );
  AND U29030 ( .A(n28685), .B(n28686), .Z(n28684) );
  XOR U29031 ( .A(e_input[342]), .B(n28683), .Z(n28686) );
  XNOR U29032 ( .A(n20496), .B(n28683), .Z(n28685) );
  XOR U29033 ( .A(n28687), .B(n28688), .Z(n20496) );
  XOR U29034 ( .A(n28689), .B(n28690), .Z(n28683) );
  AND U29035 ( .A(n28691), .B(n28692), .Z(n28690) );
  XOR U29036 ( .A(e_input[341]), .B(n28689), .Z(n28692) );
  XNOR U29037 ( .A(n20508), .B(n28689), .Z(n28691) );
  XOR U29038 ( .A(n28693), .B(n28694), .Z(n20508) );
  XOR U29039 ( .A(n28695), .B(n28696), .Z(n28689) );
  AND U29040 ( .A(n28697), .B(n28698), .Z(n28696) );
  XOR U29041 ( .A(e_input[340]), .B(n28695), .Z(n28698) );
  XNOR U29042 ( .A(n20520), .B(n28695), .Z(n28697) );
  XOR U29043 ( .A(n28699), .B(n28700), .Z(n20520) );
  XOR U29044 ( .A(n28701), .B(n28702), .Z(n28695) );
  AND U29045 ( .A(n28703), .B(n28704), .Z(n28702) );
  XOR U29046 ( .A(e_input[339]), .B(n28701), .Z(n28704) );
  XNOR U29047 ( .A(n20532), .B(n28701), .Z(n28703) );
  XOR U29048 ( .A(n28705), .B(n28706), .Z(n20532) );
  XOR U29049 ( .A(n28707), .B(n28708), .Z(n28701) );
  AND U29050 ( .A(n28709), .B(n28710), .Z(n28708) );
  XOR U29051 ( .A(e_input[338]), .B(n28707), .Z(n28710) );
  XNOR U29052 ( .A(n20544), .B(n28707), .Z(n28709) );
  XOR U29053 ( .A(n28711), .B(n28712), .Z(n20544) );
  XOR U29054 ( .A(n28713), .B(n28714), .Z(n28707) );
  AND U29055 ( .A(n28715), .B(n28716), .Z(n28714) );
  XOR U29056 ( .A(e_input[337]), .B(n28713), .Z(n28716) );
  XNOR U29057 ( .A(n20556), .B(n28713), .Z(n28715) );
  XOR U29058 ( .A(n28717), .B(n28718), .Z(n20556) );
  XOR U29059 ( .A(n28719), .B(n28720), .Z(n28713) );
  AND U29060 ( .A(n28721), .B(n28722), .Z(n28720) );
  XOR U29061 ( .A(e_input[336]), .B(n28719), .Z(n28722) );
  XNOR U29062 ( .A(n20568), .B(n28719), .Z(n28721) );
  XOR U29063 ( .A(n28723), .B(n28724), .Z(n20568) );
  XOR U29064 ( .A(n28725), .B(n28726), .Z(n28719) );
  AND U29065 ( .A(n28727), .B(n28728), .Z(n28726) );
  XOR U29066 ( .A(e_input[335]), .B(n28725), .Z(n28728) );
  XNOR U29067 ( .A(n20580), .B(n28725), .Z(n28727) );
  XOR U29068 ( .A(n28729), .B(n28730), .Z(n20580) );
  XOR U29069 ( .A(n28731), .B(n28732), .Z(n28725) );
  AND U29070 ( .A(n28733), .B(n28734), .Z(n28732) );
  XOR U29071 ( .A(e_input[334]), .B(n28731), .Z(n28734) );
  XNOR U29072 ( .A(n20592), .B(n28731), .Z(n28733) );
  XOR U29073 ( .A(n28735), .B(n28736), .Z(n20592) );
  XOR U29074 ( .A(n28737), .B(n28738), .Z(n28731) );
  AND U29075 ( .A(n28739), .B(n28740), .Z(n28738) );
  XOR U29076 ( .A(e_input[333]), .B(n28737), .Z(n28740) );
  XNOR U29077 ( .A(n20604), .B(n28737), .Z(n28739) );
  XOR U29078 ( .A(n28741), .B(n28742), .Z(n20604) );
  XOR U29079 ( .A(n28743), .B(n28744), .Z(n28737) );
  AND U29080 ( .A(n28745), .B(n28746), .Z(n28744) );
  XOR U29081 ( .A(e_input[332]), .B(n28743), .Z(n28746) );
  XNOR U29082 ( .A(n20616), .B(n28743), .Z(n28745) );
  XOR U29083 ( .A(n28747), .B(n28748), .Z(n20616) );
  XOR U29084 ( .A(n28749), .B(n28750), .Z(n28743) );
  AND U29085 ( .A(n28751), .B(n28752), .Z(n28750) );
  XOR U29086 ( .A(e_input[331]), .B(n28749), .Z(n28752) );
  XNOR U29087 ( .A(n20628), .B(n28749), .Z(n28751) );
  XOR U29088 ( .A(n28753), .B(n28754), .Z(n20628) );
  XOR U29089 ( .A(n28755), .B(n28756), .Z(n28749) );
  AND U29090 ( .A(n28757), .B(n28758), .Z(n28756) );
  XOR U29091 ( .A(e_input[330]), .B(n28755), .Z(n28758) );
  XNOR U29092 ( .A(n20640), .B(n28755), .Z(n28757) );
  XOR U29093 ( .A(n28759), .B(n28760), .Z(n20640) );
  XOR U29094 ( .A(n28761), .B(n28762), .Z(n28755) );
  AND U29095 ( .A(n28763), .B(n28764), .Z(n28762) );
  XOR U29096 ( .A(e_input[329]), .B(n28761), .Z(n28764) );
  XNOR U29097 ( .A(n20652), .B(n28761), .Z(n28763) );
  XOR U29098 ( .A(n28765), .B(n28766), .Z(n20652) );
  XOR U29099 ( .A(n28767), .B(n28768), .Z(n28761) );
  AND U29100 ( .A(n28769), .B(n28770), .Z(n28768) );
  XOR U29101 ( .A(e_input[328]), .B(n28767), .Z(n28770) );
  XNOR U29102 ( .A(n20664), .B(n28767), .Z(n28769) );
  XOR U29103 ( .A(n28771), .B(n28772), .Z(n20664) );
  XOR U29104 ( .A(n28773), .B(n28774), .Z(n28767) );
  AND U29105 ( .A(n28775), .B(n28776), .Z(n28774) );
  XOR U29106 ( .A(e_input[327]), .B(n28773), .Z(n28776) );
  XNOR U29107 ( .A(n20676), .B(n28773), .Z(n28775) );
  XOR U29108 ( .A(n28777), .B(n28778), .Z(n20676) );
  XOR U29109 ( .A(n28779), .B(n28780), .Z(n28773) );
  AND U29110 ( .A(n28781), .B(n28782), .Z(n28780) );
  XOR U29111 ( .A(e_input[326]), .B(n28779), .Z(n28782) );
  XNOR U29112 ( .A(n20688), .B(n28779), .Z(n28781) );
  XOR U29113 ( .A(n28783), .B(n28784), .Z(n20688) );
  XOR U29114 ( .A(n28785), .B(n28786), .Z(n28779) );
  AND U29115 ( .A(n28787), .B(n28788), .Z(n28786) );
  XOR U29116 ( .A(e_input[325]), .B(n28785), .Z(n28788) );
  XNOR U29117 ( .A(n20700), .B(n28785), .Z(n28787) );
  XOR U29118 ( .A(n28789), .B(n28790), .Z(n20700) );
  XOR U29119 ( .A(n28791), .B(n28792), .Z(n28785) );
  AND U29120 ( .A(n28793), .B(n28794), .Z(n28792) );
  XOR U29121 ( .A(e_input[324]), .B(n28791), .Z(n28794) );
  XNOR U29122 ( .A(n20712), .B(n28791), .Z(n28793) );
  XOR U29123 ( .A(n28795), .B(n28796), .Z(n20712) );
  XOR U29124 ( .A(n28797), .B(n28798), .Z(n28791) );
  AND U29125 ( .A(n28799), .B(n28800), .Z(n28798) );
  XOR U29126 ( .A(e_input[323]), .B(n28797), .Z(n28800) );
  XNOR U29127 ( .A(n20724), .B(n28797), .Z(n28799) );
  XOR U29128 ( .A(n28801), .B(n28802), .Z(n20724) );
  XOR U29129 ( .A(n28803), .B(n28804), .Z(n28797) );
  AND U29130 ( .A(n28805), .B(n28806), .Z(n28804) );
  XOR U29131 ( .A(e_input[322]), .B(n28803), .Z(n28806) );
  XNOR U29132 ( .A(n20736), .B(n28803), .Z(n28805) );
  XOR U29133 ( .A(n28807), .B(n28808), .Z(n20736) );
  XOR U29134 ( .A(n28809), .B(n28810), .Z(n28803) );
  AND U29135 ( .A(n28811), .B(n28812), .Z(n28810) );
  XOR U29136 ( .A(e_input[321]), .B(n28809), .Z(n28812) );
  XNOR U29137 ( .A(n20748), .B(n28809), .Z(n28811) );
  XOR U29138 ( .A(n28813), .B(n28814), .Z(n20748) );
  XOR U29139 ( .A(n28815), .B(n28816), .Z(n28809) );
  AND U29140 ( .A(n28817), .B(n28818), .Z(n28816) );
  XOR U29141 ( .A(e_input[320]), .B(n28815), .Z(n28818) );
  XNOR U29142 ( .A(n20760), .B(n28815), .Z(n28817) );
  XOR U29143 ( .A(n28819), .B(n28820), .Z(n20760) );
  XOR U29144 ( .A(n28821), .B(n28822), .Z(n28815) );
  AND U29145 ( .A(n28823), .B(n28824), .Z(n28822) );
  XOR U29146 ( .A(e_input[319]), .B(n28821), .Z(n28824) );
  XNOR U29147 ( .A(n20772), .B(n28821), .Z(n28823) );
  XOR U29148 ( .A(n28825), .B(n28826), .Z(n20772) );
  XOR U29149 ( .A(n28827), .B(n28828), .Z(n28821) );
  AND U29150 ( .A(n28829), .B(n28830), .Z(n28828) );
  XOR U29151 ( .A(e_input[318]), .B(n28827), .Z(n28830) );
  XNOR U29152 ( .A(n20784), .B(n28827), .Z(n28829) );
  XOR U29153 ( .A(n28831), .B(n28832), .Z(n20784) );
  XOR U29154 ( .A(n28833), .B(n28834), .Z(n28827) );
  AND U29155 ( .A(n28835), .B(n28836), .Z(n28834) );
  XOR U29156 ( .A(e_input[317]), .B(n28833), .Z(n28836) );
  XNOR U29157 ( .A(n20796), .B(n28833), .Z(n28835) );
  XOR U29158 ( .A(n28837), .B(n28838), .Z(n20796) );
  XOR U29159 ( .A(n28839), .B(n28840), .Z(n28833) );
  AND U29160 ( .A(n28841), .B(n28842), .Z(n28840) );
  XOR U29161 ( .A(e_input[316]), .B(n28839), .Z(n28842) );
  XNOR U29162 ( .A(n20808), .B(n28839), .Z(n28841) );
  XOR U29163 ( .A(n28843), .B(n28844), .Z(n20808) );
  XOR U29164 ( .A(n28845), .B(n28846), .Z(n28839) );
  AND U29165 ( .A(n28847), .B(n28848), .Z(n28846) );
  XOR U29166 ( .A(e_input[315]), .B(n28845), .Z(n28848) );
  XNOR U29167 ( .A(n20820), .B(n28845), .Z(n28847) );
  XOR U29168 ( .A(n28849), .B(n28850), .Z(n20820) );
  XOR U29169 ( .A(n28851), .B(n28852), .Z(n28845) );
  AND U29170 ( .A(n28853), .B(n28854), .Z(n28852) );
  XOR U29171 ( .A(e_input[314]), .B(n28851), .Z(n28854) );
  XNOR U29172 ( .A(n20832), .B(n28851), .Z(n28853) );
  XOR U29173 ( .A(n28855), .B(n28856), .Z(n20832) );
  XOR U29174 ( .A(n28857), .B(n28858), .Z(n28851) );
  AND U29175 ( .A(n28859), .B(n28860), .Z(n28858) );
  XOR U29176 ( .A(e_input[313]), .B(n28857), .Z(n28860) );
  XNOR U29177 ( .A(n20844), .B(n28857), .Z(n28859) );
  XOR U29178 ( .A(n28861), .B(n28862), .Z(n20844) );
  XOR U29179 ( .A(n28863), .B(n28864), .Z(n28857) );
  AND U29180 ( .A(n28865), .B(n28866), .Z(n28864) );
  XOR U29181 ( .A(e_input[312]), .B(n28863), .Z(n28866) );
  XNOR U29182 ( .A(n20856), .B(n28863), .Z(n28865) );
  XOR U29183 ( .A(n28867), .B(n28868), .Z(n20856) );
  XOR U29184 ( .A(n28869), .B(n28870), .Z(n28863) );
  AND U29185 ( .A(n28871), .B(n28872), .Z(n28870) );
  XOR U29186 ( .A(e_input[311]), .B(n28869), .Z(n28872) );
  XNOR U29187 ( .A(n20868), .B(n28869), .Z(n28871) );
  XOR U29188 ( .A(n28873), .B(n28874), .Z(n20868) );
  XOR U29189 ( .A(n28875), .B(n28876), .Z(n28869) );
  AND U29190 ( .A(n28877), .B(n28878), .Z(n28876) );
  XOR U29191 ( .A(e_input[310]), .B(n28875), .Z(n28878) );
  XNOR U29192 ( .A(n20880), .B(n28875), .Z(n28877) );
  XOR U29193 ( .A(n28879), .B(n28880), .Z(n20880) );
  XOR U29194 ( .A(n28881), .B(n28882), .Z(n28875) );
  AND U29195 ( .A(n28883), .B(n28884), .Z(n28882) );
  XOR U29196 ( .A(e_input[309]), .B(n28881), .Z(n28884) );
  XNOR U29197 ( .A(n20892), .B(n28881), .Z(n28883) );
  XOR U29198 ( .A(n28885), .B(n28886), .Z(n20892) );
  XOR U29199 ( .A(n28887), .B(n28888), .Z(n28881) );
  AND U29200 ( .A(n28889), .B(n28890), .Z(n28888) );
  XOR U29201 ( .A(e_input[308]), .B(n28887), .Z(n28890) );
  XNOR U29202 ( .A(n20904), .B(n28887), .Z(n28889) );
  XOR U29203 ( .A(n28891), .B(n28892), .Z(n20904) );
  XOR U29204 ( .A(n28893), .B(n28894), .Z(n28887) );
  AND U29205 ( .A(n28895), .B(n28896), .Z(n28894) );
  XOR U29206 ( .A(e_input[307]), .B(n28893), .Z(n28896) );
  XNOR U29207 ( .A(n20916), .B(n28893), .Z(n28895) );
  XOR U29208 ( .A(n28897), .B(n28898), .Z(n20916) );
  XOR U29209 ( .A(n28899), .B(n28900), .Z(n28893) );
  AND U29210 ( .A(n28901), .B(n28902), .Z(n28900) );
  XOR U29211 ( .A(e_input[306]), .B(n28899), .Z(n28902) );
  XNOR U29212 ( .A(n20928), .B(n28899), .Z(n28901) );
  XOR U29213 ( .A(n28903), .B(n28904), .Z(n20928) );
  XOR U29214 ( .A(n28905), .B(n28906), .Z(n28899) );
  AND U29215 ( .A(n28907), .B(n28908), .Z(n28906) );
  XOR U29216 ( .A(e_input[305]), .B(n28905), .Z(n28908) );
  XNOR U29217 ( .A(n20940), .B(n28905), .Z(n28907) );
  XOR U29218 ( .A(n28909), .B(n28910), .Z(n20940) );
  XOR U29219 ( .A(n28911), .B(n28912), .Z(n28905) );
  AND U29220 ( .A(n28913), .B(n28914), .Z(n28912) );
  XOR U29221 ( .A(e_input[304]), .B(n28911), .Z(n28914) );
  XNOR U29222 ( .A(n20952), .B(n28911), .Z(n28913) );
  XOR U29223 ( .A(n28915), .B(n28916), .Z(n20952) );
  XOR U29224 ( .A(n28917), .B(n28918), .Z(n28911) );
  AND U29225 ( .A(n28919), .B(n28920), .Z(n28918) );
  XOR U29226 ( .A(e_input[303]), .B(n28917), .Z(n28920) );
  XNOR U29227 ( .A(n20964), .B(n28917), .Z(n28919) );
  XOR U29228 ( .A(n28921), .B(n28922), .Z(n20964) );
  XOR U29229 ( .A(n28923), .B(n28924), .Z(n28917) );
  AND U29230 ( .A(n28925), .B(n28926), .Z(n28924) );
  XOR U29231 ( .A(e_input[302]), .B(n28923), .Z(n28926) );
  XNOR U29232 ( .A(n20976), .B(n28923), .Z(n28925) );
  XOR U29233 ( .A(n28927), .B(n28928), .Z(n20976) );
  XOR U29234 ( .A(n28929), .B(n28930), .Z(n28923) );
  AND U29235 ( .A(n28931), .B(n28932), .Z(n28930) );
  XOR U29236 ( .A(e_input[301]), .B(n28929), .Z(n28932) );
  XNOR U29237 ( .A(n20988), .B(n28929), .Z(n28931) );
  XOR U29238 ( .A(n28933), .B(n28934), .Z(n20988) );
  XOR U29239 ( .A(n28935), .B(n28936), .Z(n28929) );
  AND U29240 ( .A(n28937), .B(n28938), .Z(n28936) );
  XOR U29241 ( .A(e_input[300]), .B(n28935), .Z(n28938) );
  XNOR U29242 ( .A(n21000), .B(n28935), .Z(n28937) );
  XOR U29243 ( .A(n28939), .B(n28940), .Z(n21000) );
  XOR U29244 ( .A(n28941), .B(n28942), .Z(n28935) );
  AND U29245 ( .A(n28943), .B(n28944), .Z(n28942) );
  XOR U29246 ( .A(e_input[299]), .B(n28941), .Z(n28944) );
  XNOR U29247 ( .A(n21012), .B(n28941), .Z(n28943) );
  XOR U29248 ( .A(n28945), .B(n28946), .Z(n21012) );
  XOR U29249 ( .A(n28947), .B(n28948), .Z(n28941) );
  AND U29250 ( .A(n28949), .B(n28950), .Z(n28948) );
  XOR U29251 ( .A(e_input[298]), .B(n28947), .Z(n28950) );
  XNOR U29252 ( .A(n21024), .B(n28947), .Z(n28949) );
  XOR U29253 ( .A(n28951), .B(n28952), .Z(n21024) );
  XOR U29254 ( .A(n28953), .B(n28954), .Z(n28947) );
  AND U29255 ( .A(n28955), .B(n28956), .Z(n28954) );
  XOR U29256 ( .A(e_input[297]), .B(n28953), .Z(n28956) );
  XNOR U29257 ( .A(n21036), .B(n28953), .Z(n28955) );
  XOR U29258 ( .A(n28957), .B(n28958), .Z(n21036) );
  XOR U29259 ( .A(n28959), .B(n28960), .Z(n28953) );
  AND U29260 ( .A(n28961), .B(n28962), .Z(n28960) );
  XOR U29261 ( .A(e_input[296]), .B(n28959), .Z(n28962) );
  XNOR U29262 ( .A(n21048), .B(n28959), .Z(n28961) );
  XOR U29263 ( .A(n28963), .B(n28964), .Z(n21048) );
  XOR U29264 ( .A(n28965), .B(n28966), .Z(n28959) );
  AND U29265 ( .A(n28967), .B(n28968), .Z(n28966) );
  XOR U29266 ( .A(e_input[295]), .B(n28965), .Z(n28968) );
  XNOR U29267 ( .A(n21060), .B(n28965), .Z(n28967) );
  XOR U29268 ( .A(n28969), .B(n28970), .Z(n21060) );
  XOR U29269 ( .A(n28971), .B(n28972), .Z(n28965) );
  AND U29270 ( .A(n28973), .B(n28974), .Z(n28972) );
  XOR U29271 ( .A(e_input[294]), .B(n28971), .Z(n28974) );
  XNOR U29272 ( .A(n21072), .B(n28971), .Z(n28973) );
  XOR U29273 ( .A(n28975), .B(n28976), .Z(n21072) );
  XOR U29274 ( .A(n28977), .B(n28978), .Z(n28971) );
  AND U29275 ( .A(n28979), .B(n28980), .Z(n28978) );
  XOR U29276 ( .A(e_input[293]), .B(n28977), .Z(n28980) );
  XNOR U29277 ( .A(n21084), .B(n28977), .Z(n28979) );
  XOR U29278 ( .A(n28981), .B(n28982), .Z(n21084) );
  XOR U29279 ( .A(n28983), .B(n28984), .Z(n28977) );
  AND U29280 ( .A(n28985), .B(n28986), .Z(n28984) );
  XOR U29281 ( .A(e_input[292]), .B(n28983), .Z(n28986) );
  XNOR U29282 ( .A(n21096), .B(n28983), .Z(n28985) );
  XOR U29283 ( .A(n28987), .B(n28988), .Z(n21096) );
  XOR U29284 ( .A(n28989), .B(n28990), .Z(n28983) );
  AND U29285 ( .A(n28991), .B(n28992), .Z(n28990) );
  XOR U29286 ( .A(e_input[291]), .B(n28989), .Z(n28992) );
  XNOR U29287 ( .A(n21108), .B(n28989), .Z(n28991) );
  XOR U29288 ( .A(n28993), .B(n28994), .Z(n21108) );
  XOR U29289 ( .A(n28995), .B(n28996), .Z(n28989) );
  AND U29290 ( .A(n28997), .B(n28998), .Z(n28996) );
  XOR U29291 ( .A(e_input[290]), .B(n28995), .Z(n28998) );
  XNOR U29292 ( .A(n21120), .B(n28995), .Z(n28997) );
  XOR U29293 ( .A(n28999), .B(n29000), .Z(n21120) );
  XOR U29294 ( .A(n29001), .B(n29002), .Z(n28995) );
  AND U29295 ( .A(n29003), .B(n29004), .Z(n29002) );
  XOR U29296 ( .A(e_input[289]), .B(n29001), .Z(n29004) );
  XNOR U29297 ( .A(n21132), .B(n29001), .Z(n29003) );
  XOR U29298 ( .A(n29005), .B(n29006), .Z(n21132) );
  XOR U29299 ( .A(n29007), .B(n29008), .Z(n29001) );
  AND U29300 ( .A(n29009), .B(n29010), .Z(n29008) );
  XOR U29301 ( .A(e_input[288]), .B(n29007), .Z(n29010) );
  XNOR U29302 ( .A(n21144), .B(n29007), .Z(n29009) );
  XOR U29303 ( .A(n29011), .B(n29012), .Z(n21144) );
  XOR U29304 ( .A(n29013), .B(n29014), .Z(n29007) );
  AND U29305 ( .A(n29015), .B(n29016), .Z(n29014) );
  XOR U29306 ( .A(e_input[287]), .B(n29013), .Z(n29016) );
  XNOR U29307 ( .A(n21156), .B(n29013), .Z(n29015) );
  XOR U29308 ( .A(n29017), .B(n29018), .Z(n21156) );
  XOR U29309 ( .A(n29019), .B(n29020), .Z(n29013) );
  AND U29310 ( .A(n29021), .B(n29022), .Z(n29020) );
  XOR U29311 ( .A(e_input[286]), .B(n29019), .Z(n29022) );
  XNOR U29312 ( .A(n21168), .B(n29019), .Z(n29021) );
  XOR U29313 ( .A(n29023), .B(n29024), .Z(n21168) );
  XOR U29314 ( .A(n29025), .B(n29026), .Z(n29019) );
  AND U29315 ( .A(n29027), .B(n29028), .Z(n29026) );
  XOR U29316 ( .A(e_input[285]), .B(n29025), .Z(n29028) );
  XNOR U29317 ( .A(n21180), .B(n29025), .Z(n29027) );
  XOR U29318 ( .A(n29029), .B(n29030), .Z(n21180) );
  XOR U29319 ( .A(n29031), .B(n29032), .Z(n29025) );
  AND U29320 ( .A(n29033), .B(n29034), .Z(n29032) );
  XOR U29321 ( .A(e_input[284]), .B(n29031), .Z(n29034) );
  XNOR U29322 ( .A(n21192), .B(n29031), .Z(n29033) );
  XOR U29323 ( .A(n29035), .B(n29036), .Z(n21192) );
  XOR U29324 ( .A(n29037), .B(n29038), .Z(n29031) );
  AND U29325 ( .A(n29039), .B(n29040), .Z(n29038) );
  XOR U29326 ( .A(e_input[283]), .B(n29037), .Z(n29040) );
  XNOR U29327 ( .A(n21204), .B(n29037), .Z(n29039) );
  XOR U29328 ( .A(n29041), .B(n29042), .Z(n21204) );
  XOR U29329 ( .A(n29043), .B(n29044), .Z(n29037) );
  AND U29330 ( .A(n29045), .B(n29046), .Z(n29044) );
  XOR U29331 ( .A(e_input[282]), .B(n29043), .Z(n29046) );
  XNOR U29332 ( .A(n21216), .B(n29043), .Z(n29045) );
  XOR U29333 ( .A(n29047), .B(n29048), .Z(n21216) );
  XOR U29334 ( .A(n29049), .B(n29050), .Z(n29043) );
  AND U29335 ( .A(n29051), .B(n29052), .Z(n29050) );
  XOR U29336 ( .A(e_input[281]), .B(n29049), .Z(n29052) );
  XNOR U29337 ( .A(n21228), .B(n29049), .Z(n29051) );
  XOR U29338 ( .A(n29053), .B(n29054), .Z(n21228) );
  XOR U29339 ( .A(n29055), .B(n29056), .Z(n29049) );
  AND U29340 ( .A(n29057), .B(n29058), .Z(n29056) );
  XOR U29341 ( .A(e_input[280]), .B(n29055), .Z(n29058) );
  XNOR U29342 ( .A(n21240), .B(n29055), .Z(n29057) );
  XOR U29343 ( .A(n29059), .B(n29060), .Z(n21240) );
  XOR U29344 ( .A(n29061), .B(n29062), .Z(n29055) );
  AND U29345 ( .A(n29063), .B(n29064), .Z(n29062) );
  XOR U29346 ( .A(e_input[279]), .B(n29061), .Z(n29064) );
  XNOR U29347 ( .A(n21252), .B(n29061), .Z(n29063) );
  XOR U29348 ( .A(n29065), .B(n29066), .Z(n21252) );
  XOR U29349 ( .A(n29067), .B(n29068), .Z(n29061) );
  AND U29350 ( .A(n29069), .B(n29070), .Z(n29068) );
  XOR U29351 ( .A(e_input[278]), .B(n29067), .Z(n29070) );
  XNOR U29352 ( .A(n21264), .B(n29067), .Z(n29069) );
  XOR U29353 ( .A(n29071), .B(n29072), .Z(n21264) );
  XOR U29354 ( .A(n29073), .B(n29074), .Z(n29067) );
  AND U29355 ( .A(n29075), .B(n29076), .Z(n29074) );
  XOR U29356 ( .A(e_input[277]), .B(n29073), .Z(n29076) );
  XNOR U29357 ( .A(n21276), .B(n29073), .Z(n29075) );
  XOR U29358 ( .A(n29077), .B(n29078), .Z(n21276) );
  XOR U29359 ( .A(n29079), .B(n29080), .Z(n29073) );
  AND U29360 ( .A(n29081), .B(n29082), .Z(n29080) );
  XOR U29361 ( .A(e_input[276]), .B(n29079), .Z(n29082) );
  XNOR U29362 ( .A(n21288), .B(n29079), .Z(n29081) );
  XOR U29363 ( .A(n29083), .B(n29084), .Z(n21288) );
  XOR U29364 ( .A(n29085), .B(n29086), .Z(n29079) );
  AND U29365 ( .A(n29087), .B(n29088), .Z(n29086) );
  XOR U29366 ( .A(e_input[275]), .B(n29085), .Z(n29088) );
  XNOR U29367 ( .A(n21300), .B(n29085), .Z(n29087) );
  XOR U29368 ( .A(n29089), .B(n29090), .Z(n21300) );
  XOR U29369 ( .A(n29091), .B(n29092), .Z(n29085) );
  AND U29370 ( .A(n29093), .B(n29094), .Z(n29092) );
  XOR U29371 ( .A(e_input[274]), .B(n29091), .Z(n29094) );
  XNOR U29372 ( .A(n21312), .B(n29091), .Z(n29093) );
  XOR U29373 ( .A(n29095), .B(n29096), .Z(n21312) );
  XOR U29374 ( .A(n29097), .B(n29098), .Z(n29091) );
  AND U29375 ( .A(n29099), .B(n29100), .Z(n29098) );
  XOR U29376 ( .A(e_input[273]), .B(n29097), .Z(n29100) );
  XNOR U29377 ( .A(n21324), .B(n29097), .Z(n29099) );
  XOR U29378 ( .A(n29101), .B(n29102), .Z(n21324) );
  XOR U29379 ( .A(n29103), .B(n29104), .Z(n29097) );
  AND U29380 ( .A(n29105), .B(n29106), .Z(n29104) );
  XOR U29381 ( .A(e_input[272]), .B(n29103), .Z(n29106) );
  XNOR U29382 ( .A(n21336), .B(n29103), .Z(n29105) );
  XOR U29383 ( .A(n29107), .B(n29108), .Z(n21336) );
  XOR U29384 ( .A(n29109), .B(n29110), .Z(n29103) );
  AND U29385 ( .A(n29111), .B(n29112), .Z(n29110) );
  XOR U29386 ( .A(e_input[271]), .B(n29109), .Z(n29112) );
  XNOR U29387 ( .A(n21348), .B(n29109), .Z(n29111) );
  XOR U29388 ( .A(n29113), .B(n29114), .Z(n21348) );
  XOR U29389 ( .A(n29115), .B(n29116), .Z(n29109) );
  AND U29390 ( .A(n29117), .B(n29118), .Z(n29116) );
  XOR U29391 ( .A(e_input[270]), .B(n29115), .Z(n29118) );
  XNOR U29392 ( .A(n21360), .B(n29115), .Z(n29117) );
  XOR U29393 ( .A(n29119), .B(n29120), .Z(n21360) );
  XOR U29394 ( .A(n29121), .B(n29122), .Z(n29115) );
  AND U29395 ( .A(n29123), .B(n29124), .Z(n29122) );
  XOR U29396 ( .A(e_input[269]), .B(n29121), .Z(n29124) );
  XNOR U29397 ( .A(n21372), .B(n29121), .Z(n29123) );
  XOR U29398 ( .A(n29125), .B(n29126), .Z(n21372) );
  XOR U29399 ( .A(n29127), .B(n29128), .Z(n29121) );
  AND U29400 ( .A(n29129), .B(n29130), .Z(n29128) );
  XOR U29401 ( .A(e_input[268]), .B(n29127), .Z(n29130) );
  XNOR U29402 ( .A(n21384), .B(n29127), .Z(n29129) );
  XOR U29403 ( .A(n29131), .B(n29132), .Z(n21384) );
  XOR U29404 ( .A(n29133), .B(n29134), .Z(n29127) );
  AND U29405 ( .A(n29135), .B(n29136), .Z(n29134) );
  XOR U29406 ( .A(e_input[267]), .B(n29133), .Z(n29136) );
  XNOR U29407 ( .A(n21396), .B(n29133), .Z(n29135) );
  XOR U29408 ( .A(n29137), .B(n29138), .Z(n21396) );
  XOR U29409 ( .A(n29139), .B(n29140), .Z(n29133) );
  AND U29410 ( .A(n29141), .B(n29142), .Z(n29140) );
  XOR U29411 ( .A(e_input[266]), .B(n29139), .Z(n29142) );
  XNOR U29412 ( .A(n21408), .B(n29139), .Z(n29141) );
  XOR U29413 ( .A(n29143), .B(n29144), .Z(n21408) );
  XOR U29414 ( .A(n29145), .B(n29146), .Z(n29139) );
  AND U29415 ( .A(n29147), .B(n29148), .Z(n29146) );
  XOR U29416 ( .A(e_input[265]), .B(n29145), .Z(n29148) );
  XNOR U29417 ( .A(n21420), .B(n29145), .Z(n29147) );
  XOR U29418 ( .A(n29149), .B(n29150), .Z(n21420) );
  XOR U29419 ( .A(n29151), .B(n29152), .Z(n29145) );
  AND U29420 ( .A(n29153), .B(n29154), .Z(n29152) );
  XOR U29421 ( .A(e_input[264]), .B(n29151), .Z(n29154) );
  XNOR U29422 ( .A(n21432), .B(n29151), .Z(n29153) );
  XOR U29423 ( .A(n29155), .B(n29156), .Z(n21432) );
  XOR U29424 ( .A(n29157), .B(n29158), .Z(n29151) );
  AND U29425 ( .A(n29159), .B(n29160), .Z(n29158) );
  XOR U29426 ( .A(e_input[263]), .B(n29157), .Z(n29160) );
  XNOR U29427 ( .A(n21444), .B(n29157), .Z(n29159) );
  XOR U29428 ( .A(n29161), .B(n29162), .Z(n21444) );
  XOR U29429 ( .A(n29163), .B(n29164), .Z(n29157) );
  AND U29430 ( .A(n29165), .B(n29166), .Z(n29164) );
  XOR U29431 ( .A(e_input[262]), .B(n29163), .Z(n29166) );
  XNOR U29432 ( .A(n21456), .B(n29163), .Z(n29165) );
  XOR U29433 ( .A(n29167), .B(n29168), .Z(n21456) );
  XOR U29434 ( .A(n29169), .B(n29170), .Z(n29163) );
  AND U29435 ( .A(n29171), .B(n29172), .Z(n29170) );
  XOR U29436 ( .A(e_input[261]), .B(n29169), .Z(n29172) );
  XNOR U29437 ( .A(n21468), .B(n29169), .Z(n29171) );
  XOR U29438 ( .A(n29173), .B(n29174), .Z(n21468) );
  XOR U29439 ( .A(n29175), .B(n29176), .Z(n29169) );
  AND U29440 ( .A(n29177), .B(n29178), .Z(n29176) );
  XOR U29441 ( .A(e_input[260]), .B(n29175), .Z(n29178) );
  XNOR U29442 ( .A(n21480), .B(n29175), .Z(n29177) );
  XOR U29443 ( .A(n29179), .B(n29180), .Z(n21480) );
  XOR U29444 ( .A(n29181), .B(n29182), .Z(n29175) );
  AND U29445 ( .A(n29183), .B(n29184), .Z(n29182) );
  XOR U29446 ( .A(e_input[259]), .B(n29181), .Z(n29184) );
  XNOR U29447 ( .A(n21492), .B(n29181), .Z(n29183) );
  XOR U29448 ( .A(n29185), .B(n29186), .Z(n21492) );
  XOR U29449 ( .A(n29187), .B(n29188), .Z(n29181) );
  AND U29450 ( .A(n29189), .B(n29190), .Z(n29188) );
  XOR U29451 ( .A(e_input[258]), .B(n29187), .Z(n29190) );
  XNOR U29452 ( .A(n21504), .B(n29187), .Z(n29189) );
  XOR U29453 ( .A(n29191), .B(n29192), .Z(n21504) );
  XOR U29454 ( .A(n29193), .B(n29194), .Z(n29187) );
  AND U29455 ( .A(n29195), .B(n29196), .Z(n29194) );
  XOR U29456 ( .A(e_input[257]), .B(n29193), .Z(n29196) );
  XNOR U29457 ( .A(n21516), .B(n29193), .Z(n29195) );
  XOR U29458 ( .A(n29197), .B(n29198), .Z(n21516) );
  XOR U29459 ( .A(n29199), .B(n29200), .Z(n29193) );
  AND U29460 ( .A(n29201), .B(n29202), .Z(n29200) );
  XOR U29461 ( .A(e_input[256]), .B(n29199), .Z(n29202) );
  XNOR U29462 ( .A(n21528), .B(n29199), .Z(n29201) );
  XOR U29463 ( .A(n29203), .B(n29204), .Z(n21528) );
  XOR U29464 ( .A(n29205), .B(n29206), .Z(n29199) );
  AND U29465 ( .A(n29207), .B(n29208), .Z(n29206) );
  XOR U29466 ( .A(e_input[255]), .B(n29205), .Z(n29208) );
  XNOR U29467 ( .A(n21540), .B(n29205), .Z(n29207) );
  XOR U29468 ( .A(n29209), .B(n29210), .Z(n21540) );
  XOR U29469 ( .A(n29211), .B(n29212), .Z(n29205) );
  AND U29470 ( .A(n29213), .B(n29214), .Z(n29212) );
  XOR U29471 ( .A(e_input[254]), .B(n29211), .Z(n29214) );
  XNOR U29472 ( .A(n21552), .B(n29211), .Z(n29213) );
  XOR U29473 ( .A(n29215), .B(n29216), .Z(n21552) );
  XOR U29474 ( .A(n29217), .B(n29218), .Z(n29211) );
  AND U29475 ( .A(n29219), .B(n29220), .Z(n29218) );
  XOR U29476 ( .A(e_input[253]), .B(n29217), .Z(n29220) );
  XNOR U29477 ( .A(n21564), .B(n29217), .Z(n29219) );
  XOR U29478 ( .A(n29221), .B(n29222), .Z(n21564) );
  XOR U29479 ( .A(n29223), .B(n29224), .Z(n29217) );
  AND U29480 ( .A(n29225), .B(n29226), .Z(n29224) );
  XOR U29481 ( .A(e_input[252]), .B(n29223), .Z(n29226) );
  XNOR U29482 ( .A(n21576), .B(n29223), .Z(n29225) );
  XOR U29483 ( .A(n29227), .B(n29228), .Z(n21576) );
  XOR U29484 ( .A(n29229), .B(n29230), .Z(n29223) );
  AND U29485 ( .A(n29231), .B(n29232), .Z(n29230) );
  XOR U29486 ( .A(e_input[251]), .B(n29229), .Z(n29232) );
  XNOR U29487 ( .A(n21588), .B(n29229), .Z(n29231) );
  XOR U29488 ( .A(n29233), .B(n29234), .Z(n21588) );
  XOR U29489 ( .A(n29235), .B(n29236), .Z(n29229) );
  AND U29490 ( .A(n29237), .B(n29238), .Z(n29236) );
  XOR U29491 ( .A(e_input[250]), .B(n29235), .Z(n29238) );
  XNOR U29492 ( .A(n21600), .B(n29235), .Z(n29237) );
  XOR U29493 ( .A(n29239), .B(n29240), .Z(n21600) );
  XOR U29494 ( .A(n29241), .B(n29242), .Z(n29235) );
  AND U29495 ( .A(n29243), .B(n29244), .Z(n29242) );
  XOR U29496 ( .A(e_input[249]), .B(n29241), .Z(n29244) );
  XNOR U29497 ( .A(n21612), .B(n29241), .Z(n29243) );
  XOR U29498 ( .A(n29245), .B(n29246), .Z(n21612) );
  XOR U29499 ( .A(n29247), .B(n29248), .Z(n29241) );
  AND U29500 ( .A(n29249), .B(n29250), .Z(n29248) );
  XOR U29501 ( .A(e_input[248]), .B(n29247), .Z(n29250) );
  XNOR U29502 ( .A(n21624), .B(n29247), .Z(n29249) );
  XOR U29503 ( .A(n29251), .B(n29252), .Z(n21624) );
  XOR U29504 ( .A(n29253), .B(n29254), .Z(n29247) );
  AND U29505 ( .A(n29255), .B(n29256), .Z(n29254) );
  XOR U29506 ( .A(e_input[247]), .B(n29253), .Z(n29256) );
  XNOR U29507 ( .A(n21636), .B(n29253), .Z(n29255) );
  XOR U29508 ( .A(n29257), .B(n29258), .Z(n21636) );
  XOR U29509 ( .A(n29259), .B(n29260), .Z(n29253) );
  AND U29510 ( .A(n29261), .B(n29262), .Z(n29260) );
  XOR U29511 ( .A(e_input[246]), .B(n29259), .Z(n29262) );
  XNOR U29512 ( .A(n21648), .B(n29259), .Z(n29261) );
  XOR U29513 ( .A(n29263), .B(n29264), .Z(n21648) );
  XOR U29514 ( .A(n29265), .B(n29266), .Z(n29259) );
  AND U29515 ( .A(n29267), .B(n29268), .Z(n29266) );
  XOR U29516 ( .A(e_input[245]), .B(n29265), .Z(n29268) );
  XNOR U29517 ( .A(n21660), .B(n29265), .Z(n29267) );
  XOR U29518 ( .A(n29269), .B(n29270), .Z(n21660) );
  XOR U29519 ( .A(n29271), .B(n29272), .Z(n29265) );
  AND U29520 ( .A(n29273), .B(n29274), .Z(n29272) );
  XOR U29521 ( .A(e_input[244]), .B(n29271), .Z(n29274) );
  XNOR U29522 ( .A(n21672), .B(n29271), .Z(n29273) );
  XOR U29523 ( .A(n29275), .B(n29276), .Z(n21672) );
  XOR U29524 ( .A(n29277), .B(n29278), .Z(n29271) );
  AND U29525 ( .A(n29279), .B(n29280), .Z(n29278) );
  XOR U29526 ( .A(e_input[243]), .B(n29277), .Z(n29280) );
  XNOR U29527 ( .A(n21684), .B(n29277), .Z(n29279) );
  XOR U29528 ( .A(n29281), .B(n29282), .Z(n21684) );
  XOR U29529 ( .A(n29283), .B(n29284), .Z(n29277) );
  AND U29530 ( .A(n29285), .B(n29286), .Z(n29284) );
  XOR U29531 ( .A(e_input[242]), .B(n29283), .Z(n29286) );
  XNOR U29532 ( .A(n21696), .B(n29283), .Z(n29285) );
  XOR U29533 ( .A(n29287), .B(n29288), .Z(n21696) );
  XOR U29534 ( .A(n29289), .B(n29290), .Z(n29283) );
  AND U29535 ( .A(n29291), .B(n29292), .Z(n29290) );
  XOR U29536 ( .A(e_input[241]), .B(n29289), .Z(n29292) );
  XNOR U29537 ( .A(n21708), .B(n29289), .Z(n29291) );
  XOR U29538 ( .A(n29293), .B(n29294), .Z(n21708) );
  XOR U29539 ( .A(n29295), .B(n29296), .Z(n29289) );
  AND U29540 ( .A(n29297), .B(n29298), .Z(n29296) );
  XOR U29541 ( .A(e_input[240]), .B(n29295), .Z(n29298) );
  XNOR U29542 ( .A(n21720), .B(n29295), .Z(n29297) );
  XOR U29543 ( .A(n29299), .B(n29300), .Z(n21720) );
  XOR U29544 ( .A(n29301), .B(n29302), .Z(n29295) );
  AND U29545 ( .A(n29303), .B(n29304), .Z(n29302) );
  XOR U29546 ( .A(e_input[239]), .B(n29301), .Z(n29304) );
  XNOR U29547 ( .A(n21732), .B(n29301), .Z(n29303) );
  XOR U29548 ( .A(n29305), .B(n29306), .Z(n21732) );
  XOR U29549 ( .A(n29307), .B(n29308), .Z(n29301) );
  AND U29550 ( .A(n29309), .B(n29310), .Z(n29308) );
  XOR U29551 ( .A(e_input[238]), .B(n29307), .Z(n29310) );
  XNOR U29552 ( .A(n21744), .B(n29307), .Z(n29309) );
  XOR U29553 ( .A(n29311), .B(n29312), .Z(n21744) );
  XOR U29554 ( .A(n29313), .B(n29314), .Z(n29307) );
  AND U29555 ( .A(n29315), .B(n29316), .Z(n29314) );
  XOR U29556 ( .A(e_input[237]), .B(n29313), .Z(n29316) );
  XNOR U29557 ( .A(n21756), .B(n29313), .Z(n29315) );
  XOR U29558 ( .A(n29317), .B(n29318), .Z(n21756) );
  XOR U29559 ( .A(n29319), .B(n29320), .Z(n29313) );
  AND U29560 ( .A(n29321), .B(n29322), .Z(n29320) );
  XOR U29561 ( .A(e_input[236]), .B(n29319), .Z(n29322) );
  XNOR U29562 ( .A(n21768), .B(n29319), .Z(n29321) );
  XOR U29563 ( .A(n29323), .B(n29324), .Z(n21768) );
  XOR U29564 ( .A(n29325), .B(n29326), .Z(n29319) );
  AND U29565 ( .A(n29327), .B(n29328), .Z(n29326) );
  XOR U29566 ( .A(e_input[235]), .B(n29325), .Z(n29328) );
  XNOR U29567 ( .A(n21780), .B(n29325), .Z(n29327) );
  XOR U29568 ( .A(n29329), .B(n29330), .Z(n21780) );
  XOR U29569 ( .A(n29331), .B(n29332), .Z(n29325) );
  AND U29570 ( .A(n29333), .B(n29334), .Z(n29332) );
  XOR U29571 ( .A(e_input[234]), .B(n29331), .Z(n29334) );
  XNOR U29572 ( .A(n21792), .B(n29331), .Z(n29333) );
  XOR U29573 ( .A(n29335), .B(n29336), .Z(n21792) );
  XOR U29574 ( .A(n29337), .B(n29338), .Z(n29331) );
  AND U29575 ( .A(n29339), .B(n29340), .Z(n29338) );
  XOR U29576 ( .A(e_input[233]), .B(n29337), .Z(n29340) );
  XNOR U29577 ( .A(n21804), .B(n29337), .Z(n29339) );
  XOR U29578 ( .A(n29341), .B(n29342), .Z(n21804) );
  XOR U29579 ( .A(n29343), .B(n29344), .Z(n29337) );
  AND U29580 ( .A(n29345), .B(n29346), .Z(n29344) );
  XOR U29581 ( .A(e_input[232]), .B(n29343), .Z(n29346) );
  XNOR U29582 ( .A(n21816), .B(n29343), .Z(n29345) );
  XOR U29583 ( .A(n29347), .B(n29348), .Z(n21816) );
  XOR U29584 ( .A(n29349), .B(n29350), .Z(n29343) );
  AND U29585 ( .A(n29351), .B(n29352), .Z(n29350) );
  XOR U29586 ( .A(e_input[231]), .B(n29349), .Z(n29352) );
  XNOR U29587 ( .A(n21828), .B(n29349), .Z(n29351) );
  XOR U29588 ( .A(n29353), .B(n29354), .Z(n21828) );
  XOR U29589 ( .A(n29355), .B(n29356), .Z(n29349) );
  AND U29590 ( .A(n29357), .B(n29358), .Z(n29356) );
  XOR U29591 ( .A(e_input[230]), .B(n29355), .Z(n29358) );
  XNOR U29592 ( .A(n21840), .B(n29355), .Z(n29357) );
  XOR U29593 ( .A(n29359), .B(n29360), .Z(n21840) );
  XOR U29594 ( .A(n29361), .B(n29362), .Z(n29355) );
  AND U29595 ( .A(n29363), .B(n29364), .Z(n29362) );
  XOR U29596 ( .A(e_input[229]), .B(n29361), .Z(n29364) );
  XNOR U29597 ( .A(n21852), .B(n29361), .Z(n29363) );
  XOR U29598 ( .A(n29365), .B(n29366), .Z(n21852) );
  XOR U29599 ( .A(n29367), .B(n29368), .Z(n29361) );
  AND U29600 ( .A(n29369), .B(n29370), .Z(n29368) );
  XOR U29601 ( .A(e_input[228]), .B(n29367), .Z(n29370) );
  XNOR U29602 ( .A(n21864), .B(n29367), .Z(n29369) );
  XOR U29603 ( .A(n29371), .B(n29372), .Z(n21864) );
  XOR U29604 ( .A(n29373), .B(n29374), .Z(n29367) );
  AND U29605 ( .A(n29375), .B(n29376), .Z(n29374) );
  XOR U29606 ( .A(e_input[227]), .B(n29373), .Z(n29376) );
  XNOR U29607 ( .A(n21876), .B(n29373), .Z(n29375) );
  XOR U29608 ( .A(n29377), .B(n29378), .Z(n21876) );
  XOR U29609 ( .A(n29379), .B(n29380), .Z(n29373) );
  AND U29610 ( .A(n29381), .B(n29382), .Z(n29380) );
  XOR U29611 ( .A(e_input[226]), .B(n29379), .Z(n29382) );
  XNOR U29612 ( .A(n21888), .B(n29379), .Z(n29381) );
  XOR U29613 ( .A(n29383), .B(n29384), .Z(n21888) );
  XOR U29614 ( .A(n29385), .B(n29386), .Z(n29379) );
  AND U29615 ( .A(n29387), .B(n29388), .Z(n29386) );
  XOR U29616 ( .A(e_input[225]), .B(n29385), .Z(n29388) );
  XNOR U29617 ( .A(n21900), .B(n29385), .Z(n29387) );
  XOR U29618 ( .A(n29389), .B(n29390), .Z(n21900) );
  XOR U29619 ( .A(n29391), .B(n29392), .Z(n29385) );
  AND U29620 ( .A(n29393), .B(n29394), .Z(n29392) );
  XOR U29621 ( .A(e_input[224]), .B(n29391), .Z(n29394) );
  XNOR U29622 ( .A(n21912), .B(n29391), .Z(n29393) );
  XOR U29623 ( .A(n29395), .B(n29396), .Z(n21912) );
  XOR U29624 ( .A(n29397), .B(n29398), .Z(n29391) );
  AND U29625 ( .A(n29399), .B(n29400), .Z(n29398) );
  XOR U29626 ( .A(e_input[223]), .B(n29397), .Z(n29400) );
  XNOR U29627 ( .A(n21924), .B(n29397), .Z(n29399) );
  XOR U29628 ( .A(n29401), .B(n29402), .Z(n21924) );
  XOR U29629 ( .A(n29403), .B(n29404), .Z(n29397) );
  AND U29630 ( .A(n29405), .B(n29406), .Z(n29404) );
  XOR U29631 ( .A(e_input[222]), .B(n29403), .Z(n29406) );
  XNOR U29632 ( .A(n21936), .B(n29403), .Z(n29405) );
  XOR U29633 ( .A(n29407), .B(n29408), .Z(n21936) );
  XOR U29634 ( .A(n29409), .B(n29410), .Z(n29403) );
  AND U29635 ( .A(n29411), .B(n29412), .Z(n29410) );
  XOR U29636 ( .A(e_input[221]), .B(n29409), .Z(n29412) );
  XNOR U29637 ( .A(n21948), .B(n29409), .Z(n29411) );
  XOR U29638 ( .A(n29413), .B(n29414), .Z(n21948) );
  XOR U29639 ( .A(n29415), .B(n29416), .Z(n29409) );
  AND U29640 ( .A(n29417), .B(n29418), .Z(n29416) );
  XOR U29641 ( .A(e_input[220]), .B(n29415), .Z(n29418) );
  XNOR U29642 ( .A(n21960), .B(n29415), .Z(n29417) );
  XOR U29643 ( .A(n29419), .B(n29420), .Z(n21960) );
  XOR U29644 ( .A(n29421), .B(n29422), .Z(n29415) );
  AND U29645 ( .A(n29423), .B(n29424), .Z(n29422) );
  XOR U29646 ( .A(e_input[219]), .B(n29421), .Z(n29424) );
  XNOR U29647 ( .A(n21972), .B(n29421), .Z(n29423) );
  XOR U29648 ( .A(n29425), .B(n29426), .Z(n21972) );
  XOR U29649 ( .A(n29427), .B(n29428), .Z(n29421) );
  AND U29650 ( .A(n29429), .B(n29430), .Z(n29428) );
  XOR U29651 ( .A(e_input[218]), .B(n29427), .Z(n29430) );
  XNOR U29652 ( .A(n21984), .B(n29427), .Z(n29429) );
  XOR U29653 ( .A(n29431), .B(n29432), .Z(n21984) );
  XOR U29654 ( .A(n29433), .B(n29434), .Z(n29427) );
  AND U29655 ( .A(n29435), .B(n29436), .Z(n29434) );
  XOR U29656 ( .A(e_input[217]), .B(n29433), .Z(n29436) );
  XNOR U29657 ( .A(n21996), .B(n29433), .Z(n29435) );
  XOR U29658 ( .A(n29437), .B(n29438), .Z(n21996) );
  XOR U29659 ( .A(n29439), .B(n29440), .Z(n29433) );
  AND U29660 ( .A(n29441), .B(n29442), .Z(n29440) );
  XOR U29661 ( .A(e_input[216]), .B(n29439), .Z(n29442) );
  XNOR U29662 ( .A(n22008), .B(n29439), .Z(n29441) );
  XOR U29663 ( .A(n29443), .B(n29444), .Z(n22008) );
  XOR U29664 ( .A(n29445), .B(n29446), .Z(n29439) );
  AND U29665 ( .A(n29447), .B(n29448), .Z(n29446) );
  XOR U29666 ( .A(e_input[215]), .B(n29445), .Z(n29448) );
  XNOR U29667 ( .A(n22020), .B(n29445), .Z(n29447) );
  XOR U29668 ( .A(n29449), .B(n29450), .Z(n22020) );
  XOR U29669 ( .A(n29451), .B(n29452), .Z(n29445) );
  AND U29670 ( .A(n29453), .B(n29454), .Z(n29452) );
  XOR U29671 ( .A(e_input[214]), .B(n29451), .Z(n29454) );
  XNOR U29672 ( .A(n22032), .B(n29451), .Z(n29453) );
  XOR U29673 ( .A(n29455), .B(n29456), .Z(n22032) );
  XOR U29674 ( .A(n29457), .B(n29458), .Z(n29451) );
  AND U29675 ( .A(n29459), .B(n29460), .Z(n29458) );
  XOR U29676 ( .A(e_input[213]), .B(n29457), .Z(n29460) );
  XNOR U29677 ( .A(n22044), .B(n29457), .Z(n29459) );
  XOR U29678 ( .A(n29461), .B(n29462), .Z(n22044) );
  XOR U29679 ( .A(n29463), .B(n29464), .Z(n29457) );
  AND U29680 ( .A(n29465), .B(n29466), .Z(n29464) );
  XOR U29681 ( .A(e_input[212]), .B(n29463), .Z(n29466) );
  XNOR U29682 ( .A(n22056), .B(n29463), .Z(n29465) );
  XOR U29683 ( .A(n29467), .B(n29468), .Z(n22056) );
  XOR U29684 ( .A(n29469), .B(n29470), .Z(n29463) );
  AND U29685 ( .A(n29471), .B(n29472), .Z(n29470) );
  XOR U29686 ( .A(e_input[211]), .B(n29469), .Z(n29472) );
  XNOR U29687 ( .A(n22068), .B(n29469), .Z(n29471) );
  XOR U29688 ( .A(n29473), .B(n29474), .Z(n22068) );
  XOR U29689 ( .A(n29475), .B(n29476), .Z(n29469) );
  AND U29690 ( .A(n29477), .B(n29478), .Z(n29476) );
  XOR U29691 ( .A(e_input[210]), .B(n29475), .Z(n29478) );
  XNOR U29692 ( .A(n22080), .B(n29475), .Z(n29477) );
  XOR U29693 ( .A(n29479), .B(n29480), .Z(n22080) );
  XOR U29694 ( .A(n29481), .B(n29482), .Z(n29475) );
  AND U29695 ( .A(n29483), .B(n29484), .Z(n29482) );
  XOR U29696 ( .A(e_input[209]), .B(n29481), .Z(n29484) );
  XNOR U29697 ( .A(n22092), .B(n29481), .Z(n29483) );
  XOR U29698 ( .A(n29485), .B(n29486), .Z(n22092) );
  XOR U29699 ( .A(n29487), .B(n29488), .Z(n29481) );
  AND U29700 ( .A(n29489), .B(n29490), .Z(n29488) );
  XOR U29701 ( .A(e_input[208]), .B(n29487), .Z(n29490) );
  XNOR U29702 ( .A(n22104), .B(n29487), .Z(n29489) );
  XOR U29703 ( .A(n29491), .B(n29492), .Z(n22104) );
  XOR U29704 ( .A(n29493), .B(n29494), .Z(n29487) );
  AND U29705 ( .A(n29495), .B(n29496), .Z(n29494) );
  XOR U29706 ( .A(e_input[207]), .B(n29493), .Z(n29496) );
  XNOR U29707 ( .A(n22116), .B(n29493), .Z(n29495) );
  XOR U29708 ( .A(n29497), .B(n29498), .Z(n22116) );
  XOR U29709 ( .A(n29499), .B(n29500), .Z(n29493) );
  AND U29710 ( .A(n29501), .B(n29502), .Z(n29500) );
  XOR U29711 ( .A(e_input[206]), .B(n29499), .Z(n29502) );
  XNOR U29712 ( .A(n22128), .B(n29499), .Z(n29501) );
  XOR U29713 ( .A(n29503), .B(n29504), .Z(n22128) );
  XOR U29714 ( .A(n29505), .B(n29506), .Z(n29499) );
  AND U29715 ( .A(n29507), .B(n29508), .Z(n29506) );
  XOR U29716 ( .A(e_input[205]), .B(n29505), .Z(n29508) );
  XNOR U29717 ( .A(n22140), .B(n29505), .Z(n29507) );
  XOR U29718 ( .A(n29509), .B(n29510), .Z(n22140) );
  XOR U29719 ( .A(n29511), .B(n29512), .Z(n29505) );
  AND U29720 ( .A(n29513), .B(n29514), .Z(n29512) );
  XOR U29721 ( .A(e_input[204]), .B(n29511), .Z(n29514) );
  XNOR U29722 ( .A(n22152), .B(n29511), .Z(n29513) );
  XOR U29723 ( .A(n29515), .B(n29516), .Z(n22152) );
  XOR U29724 ( .A(n29517), .B(n29518), .Z(n29511) );
  AND U29725 ( .A(n29519), .B(n29520), .Z(n29518) );
  XOR U29726 ( .A(e_input[203]), .B(n29517), .Z(n29520) );
  XNOR U29727 ( .A(n22164), .B(n29517), .Z(n29519) );
  XOR U29728 ( .A(n29521), .B(n29522), .Z(n22164) );
  XOR U29729 ( .A(n29523), .B(n29524), .Z(n29517) );
  AND U29730 ( .A(n29525), .B(n29526), .Z(n29524) );
  XOR U29731 ( .A(e_input[202]), .B(n29523), .Z(n29526) );
  XNOR U29732 ( .A(n22176), .B(n29523), .Z(n29525) );
  XOR U29733 ( .A(n29527), .B(n29528), .Z(n22176) );
  XOR U29734 ( .A(n29529), .B(n29530), .Z(n29523) );
  AND U29735 ( .A(n29531), .B(n29532), .Z(n29530) );
  XOR U29736 ( .A(e_input[201]), .B(n29529), .Z(n29532) );
  XNOR U29737 ( .A(n22188), .B(n29529), .Z(n29531) );
  XOR U29738 ( .A(n29533), .B(n29534), .Z(n22188) );
  XOR U29739 ( .A(n29535), .B(n29536), .Z(n29529) );
  AND U29740 ( .A(n29537), .B(n29538), .Z(n29536) );
  XOR U29741 ( .A(e_input[200]), .B(n29535), .Z(n29538) );
  XNOR U29742 ( .A(n22200), .B(n29535), .Z(n29537) );
  XOR U29743 ( .A(n29539), .B(n29540), .Z(n22200) );
  XOR U29744 ( .A(n29541), .B(n29542), .Z(n29535) );
  AND U29745 ( .A(n29543), .B(n29544), .Z(n29542) );
  XOR U29746 ( .A(e_input[199]), .B(n29541), .Z(n29544) );
  XNOR U29747 ( .A(n22212), .B(n29541), .Z(n29543) );
  XOR U29748 ( .A(n29545), .B(n29546), .Z(n22212) );
  XOR U29749 ( .A(n29547), .B(n29548), .Z(n29541) );
  AND U29750 ( .A(n29549), .B(n29550), .Z(n29548) );
  XOR U29751 ( .A(e_input[198]), .B(n29547), .Z(n29550) );
  XNOR U29752 ( .A(n22224), .B(n29547), .Z(n29549) );
  XOR U29753 ( .A(n29551), .B(n29552), .Z(n22224) );
  XOR U29754 ( .A(n29553), .B(n29554), .Z(n29547) );
  AND U29755 ( .A(n29555), .B(n29556), .Z(n29554) );
  XOR U29756 ( .A(e_input[197]), .B(n29553), .Z(n29556) );
  XNOR U29757 ( .A(n22236), .B(n29553), .Z(n29555) );
  XOR U29758 ( .A(n29557), .B(n29558), .Z(n22236) );
  XOR U29759 ( .A(n29559), .B(n29560), .Z(n29553) );
  AND U29760 ( .A(n29561), .B(n29562), .Z(n29560) );
  XOR U29761 ( .A(e_input[196]), .B(n29559), .Z(n29562) );
  XNOR U29762 ( .A(n22248), .B(n29559), .Z(n29561) );
  XOR U29763 ( .A(n29563), .B(n29564), .Z(n22248) );
  XOR U29764 ( .A(n29565), .B(n29566), .Z(n29559) );
  AND U29765 ( .A(n29567), .B(n29568), .Z(n29566) );
  XOR U29766 ( .A(e_input[195]), .B(n29565), .Z(n29568) );
  XNOR U29767 ( .A(n22260), .B(n29565), .Z(n29567) );
  XOR U29768 ( .A(n29569), .B(n29570), .Z(n22260) );
  XOR U29769 ( .A(n29571), .B(n29572), .Z(n29565) );
  AND U29770 ( .A(n29573), .B(n29574), .Z(n29572) );
  XOR U29771 ( .A(e_input[194]), .B(n29571), .Z(n29574) );
  XNOR U29772 ( .A(n22272), .B(n29571), .Z(n29573) );
  XOR U29773 ( .A(n29575), .B(n29576), .Z(n22272) );
  XOR U29774 ( .A(n29577), .B(n29578), .Z(n29571) );
  AND U29775 ( .A(n29579), .B(n29580), .Z(n29578) );
  XOR U29776 ( .A(e_input[193]), .B(n29577), .Z(n29580) );
  XNOR U29777 ( .A(n22284), .B(n29577), .Z(n29579) );
  XOR U29778 ( .A(n29581), .B(n29582), .Z(n22284) );
  XOR U29779 ( .A(n29583), .B(n29584), .Z(n29577) );
  AND U29780 ( .A(n29585), .B(n29586), .Z(n29584) );
  XOR U29781 ( .A(e_input[192]), .B(n29583), .Z(n29586) );
  XNOR U29782 ( .A(n22296), .B(n29583), .Z(n29585) );
  XOR U29783 ( .A(n29587), .B(n29588), .Z(n22296) );
  XOR U29784 ( .A(n29589), .B(n29590), .Z(n29583) );
  AND U29785 ( .A(n29591), .B(n29592), .Z(n29590) );
  XOR U29786 ( .A(e_input[191]), .B(n29589), .Z(n29592) );
  XNOR U29787 ( .A(n22308), .B(n29589), .Z(n29591) );
  XOR U29788 ( .A(n29593), .B(n29594), .Z(n22308) );
  XOR U29789 ( .A(n29595), .B(n29596), .Z(n29589) );
  AND U29790 ( .A(n29597), .B(n29598), .Z(n29596) );
  XOR U29791 ( .A(e_input[190]), .B(n29595), .Z(n29598) );
  XNOR U29792 ( .A(n22320), .B(n29595), .Z(n29597) );
  XOR U29793 ( .A(n29599), .B(n29600), .Z(n22320) );
  XOR U29794 ( .A(n29601), .B(n29602), .Z(n29595) );
  AND U29795 ( .A(n29603), .B(n29604), .Z(n29602) );
  XOR U29796 ( .A(e_input[189]), .B(n29601), .Z(n29604) );
  XNOR U29797 ( .A(n22332), .B(n29601), .Z(n29603) );
  XOR U29798 ( .A(n29605), .B(n29606), .Z(n22332) );
  XOR U29799 ( .A(n29607), .B(n29608), .Z(n29601) );
  AND U29800 ( .A(n29609), .B(n29610), .Z(n29608) );
  XOR U29801 ( .A(e_input[188]), .B(n29607), .Z(n29610) );
  XNOR U29802 ( .A(n22344), .B(n29607), .Z(n29609) );
  XOR U29803 ( .A(n29611), .B(n29612), .Z(n22344) );
  XOR U29804 ( .A(n29613), .B(n29614), .Z(n29607) );
  AND U29805 ( .A(n29615), .B(n29616), .Z(n29614) );
  XOR U29806 ( .A(e_input[187]), .B(n29613), .Z(n29616) );
  XNOR U29807 ( .A(n22356), .B(n29613), .Z(n29615) );
  XOR U29808 ( .A(n29617), .B(n29618), .Z(n22356) );
  XOR U29809 ( .A(n29619), .B(n29620), .Z(n29613) );
  AND U29810 ( .A(n29621), .B(n29622), .Z(n29620) );
  XOR U29811 ( .A(e_input[186]), .B(n29619), .Z(n29622) );
  XNOR U29812 ( .A(n22368), .B(n29619), .Z(n29621) );
  XOR U29813 ( .A(n29623), .B(n29624), .Z(n22368) );
  XOR U29814 ( .A(n29625), .B(n29626), .Z(n29619) );
  AND U29815 ( .A(n29627), .B(n29628), .Z(n29626) );
  XOR U29816 ( .A(e_input[185]), .B(n29625), .Z(n29628) );
  XNOR U29817 ( .A(n22380), .B(n29625), .Z(n29627) );
  XOR U29818 ( .A(n29629), .B(n29630), .Z(n22380) );
  XOR U29819 ( .A(n29631), .B(n29632), .Z(n29625) );
  AND U29820 ( .A(n29633), .B(n29634), .Z(n29632) );
  XOR U29821 ( .A(e_input[184]), .B(n29631), .Z(n29634) );
  XNOR U29822 ( .A(n22392), .B(n29631), .Z(n29633) );
  XOR U29823 ( .A(n29635), .B(n29636), .Z(n22392) );
  XOR U29824 ( .A(n29637), .B(n29638), .Z(n29631) );
  AND U29825 ( .A(n29639), .B(n29640), .Z(n29638) );
  XOR U29826 ( .A(e_input[183]), .B(n29637), .Z(n29640) );
  XNOR U29827 ( .A(n22404), .B(n29637), .Z(n29639) );
  XOR U29828 ( .A(n29641), .B(n29642), .Z(n22404) );
  XOR U29829 ( .A(n29643), .B(n29644), .Z(n29637) );
  AND U29830 ( .A(n29645), .B(n29646), .Z(n29644) );
  XOR U29831 ( .A(e_input[182]), .B(n29643), .Z(n29646) );
  XNOR U29832 ( .A(n22416), .B(n29643), .Z(n29645) );
  XOR U29833 ( .A(n29647), .B(n29648), .Z(n22416) );
  XOR U29834 ( .A(n29649), .B(n29650), .Z(n29643) );
  AND U29835 ( .A(n29651), .B(n29652), .Z(n29650) );
  XOR U29836 ( .A(e_input[181]), .B(n29649), .Z(n29652) );
  XNOR U29837 ( .A(n22428), .B(n29649), .Z(n29651) );
  XOR U29838 ( .A(n29653), .B(n29654), .Z(n22428) );
  XOR U29839 ( .A(n29655), .B(n29656), .Z(n29649) );
  AND U29840 ( .A(n29657), .B(n29658), .Z(n29656) );
  XOR U29841 ( .A(e_input[180]), .B(n29655), .Z(n29658) );
  XNOR U29842 ( .A(n22440), .B(n29655), .Z(n29657) );
  XOR U29843 ( .A(n29659), .B(n29660), .Z(n22440) );
  XOR U29844 ( .A(n29661), .B(n29662), .Z(n29655) );
  AND U29845 ( .A(n29663), .B(n29664), .Z(n29662) );
  XOR U29846 ( .A(e_input[179]), .B(n29661), .Z(n29664) );
  XNOR U29847 ( .A(n22452), .B(n29661), .Z(n29663) );
  XOR U29848 ( .A(n29665), .B(n29666), .Z(n22452) );
  XOR U29849 ( .A(n29667), .B(n29668), .Z(n29661) );
  AND U29850 ( .A(n29669), .B(n29670), .Z(n29668) );
  XOR U29851 ( .A(e_input[178]), .B(n29667), .Z(n29670) );
  XNOR U29852 ( .A(n22464), .B(n29667), .Z(n29669) );
  XOR U29853 ( .A(n29671), .B(n29672), .Z(n22464) );
  XOR U29854 ( .A(n29673), .B(n29674), .Z(n29667) );
  AND U29855 ( .A(n29675), .B(n29676), .Z(n29674) );
  XOR U29856 ( .A(e_input[177]), .B(n29673), .Z(n29676) );
  XNOR U29857 ( .A(n22476), .B(n29673), .Z(n29675) );
  XOR U29858 ( .A(n29677), .B(n29678), .Z(n22476) );
  XOR U29859 ( .A(n29679), .B(n29680), .Z(n29673) );
  AND U29860 ( .A(n29681), .B(n29682), .Z(n29680) );
  XOR U29861 ( .A(e_input[176]), .B(n29679), .Z(n29682) );
  XNOR U29862 ( .A(n22488), .B(n29679), .Z(n29681) );
  XOR U29863 ( .A(n29683), .B(n29684), .Z(n22488) );
  XOR U29864 ( .A(n29685), .B(n29686), .Z(n29679) );
  AND U29865 ( .A(n29687), .B(n29688), .Z(n29686) );
  XOR U29866 ( .A(e_input[175]), .B(n29685), .Z(n29688) );
  XNOR U29867 ( .A(n22500), .B(n29685), .Z(n29687) );
  XOR U29868 ( .A(n29689), .B(n29690), .Z(n22500) );
  XOR U29869 ( .A(n29691), .B(n29692), .Z(n29685) );
  AND U29870 ( .A(n29693), .B(n29694), .Z(n29692) );
  XOR U29871 ( .A(e_input[174]), .B(n29691), .Z(n29694) );
  XNOR U29872 ( .A(n22512), .B(n29691), .Z(n29693) );
  XOR U29873 ( .A(n29695), .B(n29696), .Z(n22512) );
  XOR U29874 ( .A(n29697), .B(n29698), .Z(n29691) );
  AND U29875 ( .A(n29699), .B(n29700), .Z(n29698) );
  XOR U29876 ( .A(e_input[173]), .B(n29697), .Z(n29700) );
  XNOR U29877 ( .A(n22524), .B(n29697), .Z(n29699) );
  XOR U29878 ( .A(n29701), .B(n29702), .Z(n22524) );
  XOR U29879 ( .A(n29703), .B(n29704), .Z(n29697) );
  AND U29880 ( .A(n29705), .B(n29706), .Z(n29704) );
  XOR U29881 ( .A(e_input[172]), .B(n29703), .Z(n29706) );
  XNOR U29882 ( .A(n22536), .B(n29703), .Z(n29705) );
  XOR U29883 ( .A(n29707), .B(n29708), .Z(n22536) );
  XOR U29884 ( .A(n29709), .B(n29710), .Z(n29703) );
  AND U29885 ( .A(n29711), .B(n29712), .Z(n29710) );
  XOR U29886 ( .A(e_input[171]), .B(n29709), .Z(n29712) );
  XNOR U29887 ( .A(n22548), .B(n29709), .Z(n29711) );
  XOR U29888 ( .A(n29713), .B(n29714), .Z(n22548) );
  XOR U29889 ( .A(n29715), .B(n29716), .Z(n29709) );
  AND U29890 ( .A(n29717), .B(n29718), .Z(n29716) );
  XOR U29891 ( .A(e_input[170]), .B(n29715), .Z(n29718) );
  XNOR U29892 ( .A(n22560), .B(n29715), .Z(n29717) );
  XOR U29893 ( .A(n29719), .B(n29720), .Z(n22560) );
  XOR U29894 ( .A(n29721), .B(n29722), .Z(n29715) );
  AND U29895 ( .A(n29723), .B(n29724), .Z(n29722) );
  XOR U29896 ( .A(e_input[169]), .B(n29721), .Z(n29724) );
  XNOR U29897 ( .A(n22572), .B(n29721), .Z(n29723) );
  XOR U29898 ( .A(n29725), .B(n29726), .Z(n22572) );
  XOR U29899 ( .A(n29727), .B(n29728), .Z(n29721) );
  AND U29900 ( .A(n29729), .B(n29730), .Z(n29728) );
  XOR U29901 ( .A(e_input[168]), .B(n29727), .Z(n29730) );
  XNOR U29902 ( .A(n22584), .B(n29727), .Z(n29729) );
  XOR U29903 ( .A(n29731), .B(n29732), .Z(n22584) );
  XOR U29904 ( .A(n29733), .B(n29734), .Z(n29727) );
  AND U29905 ( .A(n29735), .B(n29736), .Z(n29734) );
  XOR U29906 ( .A(e_input[167]), .B(n29733), .Z(n29736) );
  XNOR U29907 ( .A(n22596), .B(n29733), .Z(n29735) );
  XOR U29908 ( .A(n29737), .B(n29738), .Z(n22596) );
  XOR U29909 ( .A(n29739), .B(n29740), .Z(n29733) );
  AND U29910 ( .A(n29741), .B(n29742), .Z(n29740) );
  XOR U29911 ( .A(e_input[166]), .B(n29739), .Z(n29742) );
  XNOR U29912 ( .A(n22608), .B(n29739), .Z(n29741) );
  XOR U29913 ( .A(n29743), .B(n29744), .Z(n22608) );
  XOR U29914 ( .A(n29745), .B(n29746), .Z(n29739) );
  AND U29915 ( .A(n29747), .B(n29748), .Z(n29746) );
  XOR U29916 ( .A(e_input[165]), .B(n29745), .Z(n29748) );
  XNOR U29917 ( .A(n22620), .B(n29745), .Z(n29747) );
  XOR U29918 ( .A(n29749), .B(n29750), .Z(n22620) );
  XOR U29919 ( .A(n29751), .B(n29752), .Z(n29745) );
  AND U29920 ( .A(n29753), .B(n29754), .Z(n29752) );
  XOR U29921 ( .A(e_input[164]), .B(n29751), .Z(n29754) );
  XNOR U29922 ( .A(n22632), .B(n29751), .Z(n29753) );
  XOR U29923 ( .A(n29755), .B(n29756), .Z(n22632) );
  XOR U29924 ( .A(n29757), .B(n29758), .Z(n29751) );
  AND U29925 ( .A(n29759), .B(n29760), .Z(n29758) );
  XOR U29926 ( .A(e_input[163]), .B(n29757), .Z(n29760) );
  XNOR U29927 ( .A(n22644), .B(n29757), .Z(n29759) );
  XOR U29928 ( .A(n29761), .B(n29762), .Z(n22644) );
  XOR U29929 ( .A(n29763), .B(n29764), .Z(n29757) );
  AND U29930 ( .A(n29765), .B(n29766), .Z(n29764) );
  XOR U29931 ( .A(e_input[162]), .B(n29763), .Z(n29766) );
  XNOR U29932 ( .A(n22656), .B(n29763), .Z(n29765) );
  XOR U29933 ( .A(n29767), .B(n29768), .Z(n22656) );
  XOR U29934 ( .A(n29769), .B(n29770), .Z(n29763) );
  AND U29935 ( .A(n29771), .B(n29772), .Z(n29770) );
  XOR U29936 ( .A(e_input[161]), .B(n29769), .Z(n29772) );
  XNOR U29937 ( .A(n22668), .B(n29769), .Z(n29771) );
  XOR U29938 ( .A(n29773), .B(n29774), .Z(n22668) );
  XOR U29939 ( .A(n29775), .B(n29776), .Z(n29769) );
  AND U29940 ( .A(n29777), .B(n29778), .Z(n29776) );
  XOR U29941 ( .A(e_input[160]), .B(n29775), .Z(n29778) );
  XNOR U29942 ( .A(n22680), .B(n29775), .Z(n29777) );
  XOR U29943 ( .A(n29779), .B(n29780), .Z(n22680) );
  XOR U29944 ( .A(n29781), .B(n29782), .Z(n29775) );
  AND U29945 ( .A(n29783), .B(n29784), .Z(n29782) );
  XOR U29946 ( .A(e_input[159]), .B(n29781), .Z(n29784) );
  XNOR U29947 ( .A(n22692), .B(n29781), .Z(n29783) );
  XOR U29948 ( .A(n29785), .B(n29786), .Z(n22692) );
  XOR U29949 ( .A(n29787), .B(n29788), .Z(n29781) );
  AND U29950 ( .A(n29789), .B(n29790), .Z(n29788) );
  XOR U29951 ( .A(e_input[158]), .B(n29787), .Z(n29790) );
  XNOR U29952 ( .A(n22704), .B(n29787), .Z(n29789) );
  XOR U29953 ( .A(n29791), .B(n29792), .Z(n22704) );
  XOR U29954 ( .A(n29793), .B(n29794), .Z(n29787) );
  AND U29955 ( .A(n29795), .B(n29796), .Z(n29794) );
  XOR U29956 ( .A(e_input[157]), .B(n29793), .Z(n29796) );
  XNOR U29957 ( .A(n22716), .B(n29793), .Z(n29795) );
  XOR U29958 ( .A(n29797), .B(n29798), .Z(n22716) );
  XOR U29959 ( .A(n29799), .B(n29800), .Z(n29793) );
  AND U29960 ( .A(n29801), .B(n29802), .Z(n29800) );
  XOR U29961 ( .A(e_input[156]), .B(n29799), .Z(n29802) );
  XNOR U29962 ( .A(n22728), .B(n29799), .Z(n29801) );
  XOR U29963 ( .A(n29803), .B(n29804), .Z(n22728) );
  XOR U29964 ( .A(n29805), .B(n29806), .Z(n29799) );
  AND U29965 ( .A(n29807), .B(n29808), .Z(n29806) );
  XOR U29966 ( .A(e_input[155]), .B(n29805), .Z(n29808) );
  XNOR U29967 ( .A(n22740), .B(n29805), .Z(n29807) );
  XOR U29968 ( .A(n29809), .B(n29810), .Z(n22740) );
  XOR U29969 ( .A(n29811), .B(n29812), .Z(n29805) );
  AND U29970 ( .A(n29813), .B(n29814), .Z(n29812) );
  XOR U29971 ( .A(e_input[154]), .B(n29811), .Z(n29814) );
  XNOR U29972 ( .A(n22752), .B(n29811), .Z(n29813) );
  XOR U29973 ( .A(n29815), .B(n29816), .Z(n22752) );
  XOR U29974 ( .A(n29817), .B(n29818), .Z(n29811) );
  AND U29975 ( .A(n29819), .B(n29820), .Z(n29818) );
  XOR U29976 ( .A(e_input[153]), .B(n29817), .Z(n29820) );
  XNOR U29977 ( .A(n22764), .B(n29817), .Z(n29819) );
  XOR U29978 ( .A(n29821), .B(n29822), .Z(n22764) );
  XOR U29979 ( .A(n29823), .B(n29824), .Z(n29817) );
  AND U29980 ( .A(n29825), .B(n29826), .Z(n29824) );
  XOR U29981 ( .A(e_input[152]), .B(n29823), .Z(n29826) );
  XNOR U29982 ( .A(n22776), .B(n29823), .Z(n29825) );
  XOR U29983 ( .A(n29827), .B(n29828), .Z(n22776) );
  XOR U29984 ( .A(n29829), .B(n29830), .Z(n29823) );
  AND U29985 ( .A(n29831), .B(n29832), .Z(n29830) );
  XOR U29986 ( .A(e_input[151]), .B(n29829), .Z(n29832) );
  XNOR U29987 ( .A(n22788), .B(n29829), .Z(n29831) );
  XOR U29988 ( .A(n29833), .B(n29834), .Z(n22788) );
  XOR U29989 ( .A(n29835), .B(n29836), .Z(n29829) );
  AND U29990 ( .A(n29837), .B(n29838), .Z(n29836) );
  XOR U29991 ( .A(e_input[150]), .B(n29835), .Z(n29838) );
  XNOR U29992 ( .A(n22800), .B(n29835), .Z(n29837) );
  XOR U29993 ( .A(n29839), .B(n29840), .Z(n22800) );
  XOR U29994 ( .A(n29841), .B(n29842), .Z(n29835) );
  AND U29995 ( .A(n29843), .B(n29844), .Z(n29842) );
  XOR U29996 ( .A(e_input[149]), .B(n29841), .Z(n29844) );
  XNOR U29997 ( .A(n22812), .B(n29841), .Z(n29843) );
  XOR U29998 ( .A(n29845), .B(n29846), .Z(n22812) );
  XOR U29999 ( .A(n29847), .B(n29848), .Z(n29841) );
  AND U30000 ( .A(n29849), .B(n29850), .Z(n29848) );
  XOR U30001 ( .A(e_input[148]), .B(n29847), .Z(n29850) );
  XNOR U30002 ( .A(n22824), .B(n29847), .Z(n29849) );
  XOR U30003 ( .A(n29851), .B(n29852), .Z(n22824) );
  XOR U30004 ( .A(n29853), .B(n29854), .Z(n29847) );
  AND U30005 ( .A(n29855), .B(n29856), .Z(n29854) );
  XOR U30006 ( .A(e_input[147]), .B(n29853), .Z(n29856) );
  XNOR U30007 ( .A(n22836), .B(n29853), .Z(n29855) );
  XOR U30008 ( .A(n29857), .B(n29858), .Z(n22836) );
  XOR U30009 ( .A(n29859), .B(n29860), .Z(n29853) );
  AND U30010 ( .A(n29861), .B(n29862), .Z(n29860) );
  XOR U30011 ( .A(e_input[146]), .B(n29859), .Z(n29862) );
  XNOR U30012 ( .A(n22848), .B(n29859), .Z(n29861) );
  XOR U30013 ( .A(n29863), .B(n29864), .Z(n22848) );
  XOR U30014 ( .A(n29865), .B(n29866), .Z(n29859) );
  AND U30015 ( .A(n29867), .B(n29868), .Z(n29866) );
  XOR U30016 ( .A(e_input[145]), .B(n29865), .Z(n29868) );
  XNOR U30017 ( .A(n22860), .B(n29865), .Z(n29867) );
  XOR U30018 ( .A(n29869), .B(n29870), .Z(n22860) );
  XOR U30019 ( .A(n29871), .B(n29872), .Z(n29865) );
  AND U30020 ( .A(n29873), .B(n29874), .Z(n29872) );
  XOR U30021 ( .A(e_input[144]), .B(n29871), .Z(n29874) );
  XNOR U30022 ( .A(n22872), .B(n29871), .Z(n29873) );
  XOR U30023 ( .A(n29875), .B(n29876), .Z(n22872) );
  XOR U30024 ( .A(n29877), .B(n29878), .Z(n29871) );
  AND U30025 ( .A(n29879), .B(n29880), .Z(n29878) );
  XOR U30026 ( .A(e_input[143]), .B(n29877), .Z(n29880) );
  XNOR U30027 ( .A(n22884), .B(n29877), .Z(n29879) );
  XOR U30028 ( .A(n29881), .B(n29882), .Z(n22884) );
  XOR U30029 ( .A(n29883), .B(n29884), .Z(n29877) );
  AND U30030 ( .A(n29885), .B(n29886), .Z(n29884) );
  XOR U30031 ( .A(e_input[142]), .B(n29883), .Z(n29886) );
  XNOR U30032 ( .A(n22896), .B(n29883), .Z(n29885) );
  XOR U30033 ( .A(n29887), .B(n29888), .Z(n22896) );
  XOR U30034 ( .A(n29889), .B(n29890), .Z(n29883) );
  AND U30035 ( .A(n29891), .B(n29892), .Z(n29890) );
  XOR U30036 ( .A(e_input[141]), .B(n29889), .Z(n29892) );
  XNOR U30037 ( .A(n22908), .B(n29889), .Z(n29891) );
  XOR U30038 ( .A(n29893), .B(n29894), .Z(n22908) );
  XOR U30039 ( .A(n29895), .B(n29896), .Z(n29889) );
  AND U30040 ( .A(n29897), .B(n29898), .Z(n29896) );
  XOR U30041 ( .A(e_input[140]), .B(n29895), .Z(n29898) );
  XNOR U30042 ( .A(n22920), .B(n29895), .Z(n29897) );
  XOR U30043 ( .A(n29899), .B(n29900), .Z(n22920) );
  XOR U30044 ( .A(n29901), .B(n29902), .Z(n29895) );
  AND U30045 ( .A(n29903), .B(n29904), .Z(n29902) );
  XOR U30046 ( .A(e_input[139]), .B(n29901), .Z(n29904) );
  XNOR U30047 ( .A(n22932), .B(n29901), .Z(n29903) );
  XOR U30048 ( .A(n29905), .B(n29906), .Z(n22932) );
  XOR U30049 ( .A(n29907), .B(n29908), .Z(n29901) );
  AND U30050 ( .A(n29909), .B(n29910), .Z(n29908) );
  XOR U30051 ( .A(e_input[138]), .B(n29907), .Z(n29910) );
  XNOR U30052 ( .A(n22944), .B(n29907), .Z(n29909) );
  XOR U30053 ( .A(n29911), .B(n29912), .Z(n22944) );
  XOR U30054 ( .A(n29913), .B(n29914), .Z(n29907) );
  AND U30055 ( .A(n29915), .B(n29916), .Z(n29914) );
  XOR U30056 ( .A(e_input[137]), .B(n29913), .Z(n29916) );
  XNOR U30057 ( .A(n22956), .B(n29913), .Z(n29915) );
  XOR U30058 ( .A(n29917), .B(n29918), .Z(n22956) );
  XOR U30059 ( .A(n29919), .B(n29920), .Z(n29913) );
  AND U30060 ( .A(n29921), .B(n29922), .Z(n29920) );
  XOR U30061 ( .A(e_input[136]), .B(n29919), .Z(n29922) );
  XNOR U30062 ( .A(n22968), .B(n29919), .Z(n29921) );
  XOR U30063 ( .A(n29923), .B(n29924), .Z(n22968) );
  XOR U30064 ( .A(n29925), .B(n29926), .Z(n29919) );
  AND U30065 ( .A(n29927), .B(n29928), .Z(n29926) );
  XOR U30066 ( .A(e_input[135]), .B(n29925), .Z(n29928) );
  XNOR U30067 ( .A(n22980), .B(n29925), .Z(n29927) );
  XOR U30068 ( .A(n29929), .B(n29930), .Z(n22980) );
  XOR U30069 ( .A(n29931), .B(n29932), .Z(n29925) );
  AND U30070 ( .A(n29933), .B(n29934), .Z(n29932) );
  XOR U30071 ( .A(e_input[134]), .B(n29931), .Z(n29934) );
  XNOR U30072 ( .A(n22992), .B(n29931), .Z(n29933) );
  XOR U30073 ( .A(n29935), .B(n29936), .Z(n22992) );
  XOR U30074 ( .A(n29937), .B(n29938), .Z(n29931) );
  AND U30075 ( .A(n29939), .B(n29940), .Z(n29938) );
  XOR U30076 ( .A(e_input[133]), .B(n29937), .Z(n29940) );
  XNOR U30077 ( .A(n23004), .B(n29937), .Z(n29939) );
  XOR U30078 ( .A(n29941), .B(n29942), .Z(n23004) );
  XOR U30079 ( .A(n29943), .B(n29944), .Z(n29937) );
  AND U30080 ( .A(n29945), .B(n29946), .Z(n29944) );
  XOR U30081 ( .A(e_input[132]), .B(n29943), .Z(n29946) );
  XNOR U30082 ( .A(n23016), .B(n29943), .Z(n29945) );
  XOR U30083 ( .A(n29947), .B(n29948), .Z(n23016) );
  XOR U30084 ( .A(n29949), .B(n29950), .Z(n29943) );
  AND U30085 ( .A(n29951), .B(n29952), .Z(n29950) );
  XOR U30086 ( .A(e_input[131]), .B(n29949), .Z(n29952) );
  XNOR U30087 ( .A(n23028), .B(n29949), .Z(n29951) );
  XOR U30088 ( .A(n29953), .B(n29954), .Z(n23028) );
  XOR U30089 ( .A(n29955), .B(n29956), .Z(n29949) );
  AND U30090 ( .A(n29957), .B(n29958), .Z(n29956) );
  XOR U30091 ( .A(e_input[130]), .B(n29955), .Z(n29958) );
  XNOR U30092 ( .A(n23040), .B(n29955), .Z(n29957) );
  XOR U30093 ( .A(n29959), .B(n29960), .Z(n23040) );
  XOR U30094 ( .A(n29961), .B(n29962), .Z(n29955) );
  AND U30095 ( .A(n29963), .B(n29964), .Z(n29962) );
  XOR U30096 ( .A(e_input[129]), .B(n29961), .Z(n29964) );
  XNOR U30097 ( .A(n23052), .B(n29961), .Z(n29963) );
  XOR U30098 ( .A(n29965), .B(n29966), .Z(n23052) );
  XOR U30099 ( .A(n29967), .B(n29968), .Z(n29961) );
  AND U30100 ( .A(n29969), .B(n29970), .Z(n29968) );
  XOR U30101 ( .A(e_input[128]), .B(n29967), .Z(n29970) );
  XNOR U30102 ( .A(n23064), .B(n29967), .Z(n29969) );
  XOR U30103 ( .A(n29971), .B(n29972), .Z(n23064) );
  XOR U30104 ( .A(n29973), .B(n29974), .Z(n29967) );
  AND U30105 ( .A(n29975), .B(n29976), .Z(n29974) );
  XOR U30106 ( .A(e_input[127]), .B(n29973), .Z(n29976) );
  XNOR U30107 ( .A(n23076), .B(n29973), .Z(n29975) );
  XOR U30108 ( .A(n29977), .B(n29978), .Z(n23076) );
  XOR U30109 ( .A(n29979), .B(n29980), .Z(n29973) );
  AND U30110 ( .A(n29981), .B(n29982), .Z(n29980) );
  XOR U30111 ( .A(e_input[126]), .B(n29979), .Z(n29982) );
  XNOR U30112 ( .A(n23088), .B(n29979), .Z(n29981) );
  XOR U30113 ( .A(n29983), .B(n29984), .Z(n23088) );
  XOR U30114 ( .A(n29985), .B(n29986), .Z(n29979) );
  AND U30115 ( .A(n29987), .B(n29988), .Z(n29986) );
  XOR U30116 ( .A(e_input[125]), .B(n29985), .Z(n29988) );
  XNOR U30117 ( .A(n23100), .B(n29985), .Z(n29987) );
  XOR U30118 ( .A(n29989), .B(n29990), .Z(n23100) );
  XOR U30119 ( .A(n29991), .B(n29992), .Z(n29985) );
  AND U30120 ( .A(n29993), .B(n29994), .Z(n29992) );
  XOR U30121 ( .A(e_input[124]), .B(n29991), .Z(n29994) );
  XNOR U30122 ( .A(n23112), .B(n29991), .Z(n29993) );
  XOR U30123 ( .A(n29995), .B(n29996), .Z(n23112) );
  XOR U30124 ( .A(n29997), .B(n29998), .Z(n29991) );
  AND U30125 ( .A(n29999), .B(n30000), .Z(n29998) );
  XOR U30126 ( .A(e_input[123]), .B(n29997), .Z(n30000) );
  XNOR U30127 ( .A(n23124), .B(n29997), .Z(n29999) );
  XOR U30128 ( .A(n30001), .B(n30002), .Z(n23124) );
  XOR U30129 ( .A(n30003), .B(n30004), .Z(n29997) );
  AND U30130 ( .A(n30005), .B(n30006), .Z(n30004) );
  XOR U30131 ( .A(e_input[122]), .B(n30003), .Z(n30006) );
  XNOR U30132 ( .A(n23136), .B(n30003), .Z(n30005) );
  XOR U30133 ( .A(n30007), .B(n30008), .Z(n23136) );
  XOR U30134 ( .A(n30009), .B(n30010), .Z(n30003) );
  AND U30135 ( .A(n30011), .B(n30012), .Z(n30010) );
  XOR U30136 ( .A(e_input[121]), .B(n30009), .Z(n30012) );
  XNOR U30137 ( .A(n23148), .B(n30009), .Z(n30011) );
  XOR U30138 ( .A(n30013), .B(n30014), .Z(n23148) );
  XOR U30139 ( .A(n30015), .B(n30016), .Z(n30009) );
  AND U30140 ( .A(n30017), .B(n30018), .Z(n30016) );
  XOR U30141 ( .A(e_input[120]), .B(n30015), .Z(n30018) );
  XNOR U30142 ( .A(n23160), .B(n30015), .Z(n30017) );
  XOR U30143 ( .A(n30019), .B(n30020), .Z(n23160) );
  XOR U30144 ( .A(n30021), .B(n30022), .Z(n30015) );
  AND U30145 ( .A(n30023), .B(n30024), .Z(n30022) );
  XOR U30146 ( .A(e_input[119]), .B(n30021), .Z(n30024) );
  XNOR U30147 ( .A(n23172), .B(n30021), .Z(n30023) );
  XOR U30148 ( .A(n30025), .B(n30026), .Z(n23172) );
  XOR U30149 ( .A(n30027), .B(n30028), .Z(n30021) );
  AND U30150 ( .A(n30029), .B(n30030), .Z(n30028) );
  XOR U30151 ( .A(e_input[118]), .B(n30027), .Z(n30030) );
  XNOR U30152 ( .A(n23184), .B(n30027), .Z(n30029) );
  XOR U30153 ( .A(n30031), .B(n30032), .Z(n23184) );
  XOR U30154 ( .A(n30033), .B(n30034), .Z(n30027) );
  AND U30155 ( .A(n30035), .B(n30036), .Z(n30034) );
  XOR U30156 ( .A(e_input[117]), .B(n30033), .Z(n30036) );
  XNOR U30157 ( .A(n23196), .B(n30033), .Z(n30035) );
  XOR U30158 ( .A(n30037), .B(n30038), .Z(n23196) );
  XOR U30159 ( .A(n30039), .B(n30040), .Z(n30033) );
  AND U30160 ( .A(n30041), .B(n30042), .Z(n30040) );
  XOR U30161 ( .A(e_input[116]), .B(n30039), .Z(n30042) );
  XNOR U30162 ( .A(n23208), .B(n30039), .Z(n30041) );
  XOR U30163 ( .A(n30043), .B(n30044), .Z(n23208) );
  XOR U30164 ( .A(n30045), .B(n30046), .Z(n30039) );
  AND U30165 ( .A(n30047), .B(n30048), .Z(n30046) );
  XOR U30166 ( .A(e_input[115]), .B(n30045), .Z(n30048) );
  XNOR U30167 ( .A(n23220), .B(n30045), .Z(n30047) );
  XOR U30168 ( .A(n30049), .B(n30050), .Z(n23220) );
  XOR U30169 ( .A(n30051), .B(n30052), .Z(n30045) );
  AND U30170 ( .A(n30053), .B(n30054), .Z(n30052) );
  XOR U30171 ( .A(e_input[114]), .B(n30051), .Z(n30054) );
  XNOR U30172 ( .A(n23232), .B(n30051), .Z(n30053) );
  XOR U30173 ( .A(n30055), .B(n30056), .Z(n23232) );
  XOR U30174 ( .A(n30057), .B(n30058), .Z(n30051) );
  AND U30175 ( .A(n30059), .B(n30060), .Z(n30058) );
  XOR U30176 ( .A(e_input[113]), .B(n30057), .Z(n30060) );
  XNOR U30177 ( .A(n23244), .B(n30057), .Z(n30059) );
  XOR U30178 ( .A(n30061), .B(n30062), .Z(n23244) );
  XOR U30179 ( .A(n30063), .B(n30064), .Z(n30057) );
  AND U30180 ( .A(n30065), .B(n30066), .Z(n30064) );
  XOR U30181 ( .A(e_input[112]), .B(n30063), .Z(n30066) );
  XNOR U30182 ( .A(n23256), .B(n30063), .Z(n30065) );
  XOR U30183 ( .A(n30067), .B(n30068), .Z(n23256) );
  XOR U30184 ( .A(n30069), .B(n30070), .Z(n30063) );
  AND U30185 ( .A(n30071), .B(n30072), .Z(n30070) );
  XOR U30186 ( .A(e_input[111]), .B(n30069), .Z(n30072) );
  XNOR U30187 ( .A(n23268), .B(n30069), .Z(n30071) );
  XOR U30188 ( .A(n30073), .B(n30074), .Z(n23268) );
  XOR U30189 ( .A(n30075), .B(n30076), .Z(n30069) );
  AND U30190 ( .A(n30077), .B(n30078), .Z(n30076) );
  XOR U30191 ( .A(e_input[110]), .B(n30075), .Z(n30078) );
  XNOR U30192 ( .A(n23280), .B(n30075), .Z(n30077) );
  XOR U30193 ( .A(n30079), .B(n30080), .Z(n23280) );
  XOR U30194 ( .A(n30081), .B(n30082), .Z(n30075) );
  AND U30195 ( .A(n30083), .B(n30084), .Z(n30082) );
  XOR U30196 ( .A(e_input[109]), .B(n30081), .Z(n30084) );
  XNOR U30197 ( .A(n23292), .B(n30081), .Z(n30083) );
  XOR U30198 ( .A(n30085), .B(n30086), .Z(n23292) );
  XOR U30199 ( .A(n30087), .B(n30088), .Z(n30081) );
  AND U30200 ( .A(n30089), .B(n30090), .Z(n30088) );
  XOR U30201 ( .A(e_input[108]), .B(n30087), .Z(n30090) );
  XNOR U30202 ( .A(n23304), .B(n30087), .Z(n30089) );
  XOR U30203 ( .A(n30091), .B(n30092), .Z(n23304) );
  XOR U30204 ( .A(n30093), .B(n30094), .Z(n30087) );
  AND U30205 ( .A(n30095), .B(n30096), .Z(n30094) );
  XOR U30206 ( .A(e_input[107]), .B(n30093), .Z(n30096) );
  XNOR U30207 ( .A(n23316), .B(n30093), .Z(n30095) );
  XOR U30208 ( .A(n30097), .B(n30098), .Z(n23316) );
  XOR U30209 ( .A(n30099), .B(n30100), .Z(n30093) );
  AND U30210 ( .A(n30101), .B(n30102), .Z(n30100) );
  XOR U30211 ( .A(e_input[106]), .B(n30099), .Z(n30102) );
  XNOR U30212 ( .A(n23328), .B(n30099), .Z(n30101) );
  XOR U30213 ( .A(n30103), .B(n30104), .Z(n23328) );
  XOR U30214 ( .A(n30105), .B(n30106), .Z(n30099) );
  AND U30215 ( .A(n30107), .B(n30108), .Z(n30106) );
  XOR U30216 ( .A(e_input[105]), .B(n30105), .Z(n30108) );
  XNOR U30217 ( .A(n23340), .B(n30105), .Z(n30107) );
  XOR U30218 ( .A(n30109), .B(n30110), .Z(n23340) );
  XOR U30219 ( .A(n30111), .B(n30112), .Z(n30105) );
  AND U30220 ( .A(n30113), .B(n30114), .Z(n30112) );
  XOR U30221 ( .A(e_input[104]), .B(n30111), .Z(n30114) );
  XNOR U30222 ( .A(n23352), .B(n30111), .Z(n30113) );
  XOR U30223 ( .A(n30115), .B(n30116), .Z(n23352) );
  XOR U30224 ( .A(n30117), .B(n30118), .Z(n30111) );
  AND U30225 ( .A(n30119), .B(n30120), .Z(n30118) );
  XOR U30226 ( .A(e_input[103]), .B(n30117), .Z(n30120) );
  XNOR U30227 ( .A(n23364), .B(n30117), .Z(n30119) );
  XOR U30228 ( .A(n30121), .B(n30122), .Z(n23364) );
  XOR U30229 ( .A(n30123), .B(n30124), .Z(n30117) );
  AND U30230 ( .A(n30125), .B(n30126), .Z(n30124) );
  XOR U30231 ( .A(e_input[102]), .B(n30123), .Z(n30126) );
  XNOR U30232 ( .A(n23376), .B(n30123), .Z(n30125) );
  XOR U30233 ( .A(n30127), .B(n30128), .Z(n23376) );
  XOR U30234 ( .A(n30129), .B(n30130), .Z(n30123) );
  AND U30235 ( .A(n30131), .B(n30132), .Z(n30130) );
  XOR U30236 ( .A(e_input[101]), .B(n30129), .Z(n30132) );
  XNOR U30237 ( .A(n23388), .B(n30129), .Z(n30131) );
  XOR U30238 ( .A(n30133), .B(n30134), .Z(n23388) );
  XOR U30239 ( .A(n30135), .B(n30136), .Z(n30129) );
  AND U30240 ( .A(n30137), .B(n30138), .Z(n30136) );
  XOR U30241 ( .A(e_input[100]), .B(n30135), .Z(n30138) );
  XNOR U30242 ( .A(n23400), .B(n30135), .Z(n30137) );
  XOR U30243 ( .A(n30139), .B(n30140), .Z(n23400) );
  XOR U30244 ( .A(n30141), .B(n30142), .Z(n30135) );
  AND U30245 ( .A(n30143), .B(n30144), .Z(n30142) );
  XOR U30246 ( .A(e_input[99]), .B(n30141), .Z(n30144) );
  XNOR U30247 ( .A(n23412), .B(n30141), .Z(n30143) );
  XOR U30248 ( .A(n30145), .B(n30146), .Z(n23412) );
  XOR U30249 ( .A(n30147), .B(n30148), .Z(n30141) );
  AND U30250 ( .A(n30149), .B(n30150), .Z(n30148) );
  XOR U30251 ( .A(e_input[98]), .B(n30147), .Z(n30150) );
  XNOR U30252 ( .A(n23424), .B(n30147), .Z(n30149) );
  XOR U30253 ( .A(n30151), .B(n30152), .Z(n23424) );
  XOR U30254 ( .A(n30153), .B(n30154), .Z(n30147) );
  AND U30255 ( .A(n30155), .B(n30156), .Z(n30154) );
  XOR U30256 ( .A(e_input[97]), .B(n30153), .Z(n30156) );
  XNOR U30257 ( .A(n23436), .B(n30153), .Z(n30155) );
  XOR U30258 ( .A(n30157), .B(n30158), .Z(n23436) );
  XOR U30259 ( .A(n30159), .B(n30160), .Z(n30153) );
  AND U30260 ( .A(n30161), .B(n30162), .Z(n30160) );
  XOR U30261 ( .A(e_input[96]), .B(n30159), .Z(n30162) );
  XNOR U30262 ( .A(n23448), .B(n30159), .Z(n30161) );
  XOR U30263 ( .A(n30163), .B(n30164), .Z(n23448) );
  XOR U30264 ( .A(n30165), .B(n30166), .Z(n30159) );
  AND U30265 ( .A(n30167), .B(n30168), .Z(n30166) );
  XOR U30266 ( .A(e_input[95]), .B(n30165), .Z(n30168) );
  XNOR U30267 ( .A(n23460), .B(n30165), .Z(n30167) );
  XOR U30268 ( .A(n30169), .B(n30170), .Z(n23460) );
  XOR U30269 ( .A(n30171), .B(n30172), .Z(n30165) );
  AND U30270 ( .A(n30173), .B(n30174), .Z(n30172) );
  XOR U30271 ( .A(e_input[94]), .B(n30171), .Z(n30174) );
  XNOR U30272 ( .A(n23472), .B(n30171), .Z(n30173) );
  XOR U30273 ( .A(n30175), .B(n30176), .Z(n23472) );
  XOR U30274 ( .A(n30177), .B(n30178), .Z(n30171) );
  AND U30275 ( .A(n30179), .B(n30180), .Z(n30178) );
  XOR U30276 ( .A(e_input[93]), .B(n30177), .Z(n30180) );
  XNOR U30277 ( .A(n23484), .B(n30177), .Z(n30179) );
  XOR U30278 ( .A(n30181), .B(n30182), .Z(n23484) );
  XOR U30279 ( .A(n30183), .B(n30184), .Z(n30177) );
  AND U30280 ( .A(n30185), .B(n30186), .Z(n30184) );
  XOR U30281 ( .A(e_input[92]), .B(n30183), .Z(n30186) );
  XNOR U30282 ( .A(n23496), .B(n30183), .Z(n30185) );
  XOR U30283 ( .A(n30187), .B(n30188), .Z(n23496) );
  XOR U30284 ( .A(n30189), .B(n30190), .Z(n30183) );
  AND U30285 ( .A(n30191), .B(n30192), .Z(n30190) );
  XOR U30286 ( .A(e_input[91]), .B(n30189), .Z(n30192) );
  XNOR U30287 ( .A(n23508), .B(n30189), .Z(n30191) );
  XOR U30288 ( .A(n30193), .B(n30194), .Z(n23508) );
  XOR U30289 ( .A(n30195), .B(n30196), .Z(n30189) );
  AND U30290 ( .A(n30197), .B(n30198), .Z(n30196) );
  XOR U30291 ( .A(e_input[90]), .B(n30195), .Z(n30198) );
  XNOR U30292 ( .A(n23520), .B(n30195), .Z(n30197) );
  XOR U30293 ( .A(n30199), .B(n30200), .Z(n23520) );
  XOR U30294 ( .A(n30201), .B(n30202), .Z(n30195) );
  AND U30295 ( .A(n30203), .B(n30204), .Z(n30202) );
  XOR U30296 ( .A(e_input[89]), .B(n30201), .Z(n30204) );
  XNOR U30297 ( .A(n23532), .B(n30201), .Z(n30203) );
  XOR U30298 ( .A(n30205), .B(n30206), .Z(n23532) );
  XOR U30299 ( .A(n30207), .B(n30208), .Z(n30201) );
  AND U30300 ( .A(n30209), .B(n30210), .Z(n30208) );
  XOR U30301 ( .A(e_input[88]), .B(n30207), .Z(n30210) );
  XNOR U30302 ( .A(n23544), .B(n30207), .Z(n30209) );
  XOR U30303 ( .A(n30211), .B(n30212), .Z(n23544) );
  XOR U30304 ( .A(n30213), .B(n30214), .Z(n30207) );
  AND U30305 ( .A(n30215), .B(n30216), .Z(n30214) );
  XOR U30306 ( .A(e_input[87]), .B(n30213), .Z(n30216) );
  XNOR U30307 ( .A(n23556), .B(n30213), .Z(n30215) );
  XOR U30308 ( .A(n30217), .B(n30218), .Z(n23556) );
  XOR U30309 ( .A(n30219), .B(n30220), .Z(n30213) );
  AND U30310 ( .A(n30221), .B(n30222), .Z(n30220) );
  XOR U30311 ( .A(e_input[86]), .B(n30219), .Z(n30222) );
  XNOR U30312 ( .A(n23568), .B(n30219), .Z(n30221) );
  XOR U30313 ( .A(n30223), .B(n30224), .Z(n23568) );
  XOR U30314 ( .A(n30225), .B(n30226), .Z(n30219) );
  AND U30315 ( .A(n30227), .B(n30228), .Z(n30226) );
  XOR U30316 ( .A(e_input[85]), .B(n30225), .Z(n30228) );
  XNOR U30317 ( .A(n23580), .B(n30225), .Z(n30227) );
  XOR U30318 ( .A(n30229), .B(n30230), .Z(n23580) );
  XOR U30319 ( .A(n30231), .B(n30232), .Z(n30225) );
  AND U30320 ( .A(n30233), .B(n30234), .Z(n30232) );
  XOR U30321 ( .A(e_input[84]), .B(n30231), .Z(n30234) );
  XNOR U30322 ( .A(n23592), .B(n30231), .Z(n30233) );
  XOR U30323 ( .A(n30235), .B(n30236), .Z(n23592) );
  XOR U30324 ( .A(n30237), .B(n30238), .Z(n30231) );
  AND U30325 ( .A(n30239), .B(n30240), .Z(n30238) );
  XOR U30326 ( .A(e_input[83]), .B(n30237), .Z(n30240) );
  XNOR U30327 ( .A(n23604), .B(n30237), .Z(n30239) );
  XOR U30328 ( .A(n30241), .B(n30242), .Z(n23604) );
  XOR U30329 ( .A(n30243), .B(n30244), .Z(n30237) );
  AND U30330 ( .A(n30245), .B(n30246), .Z(n30244) );
  XOR U30331 ( .A(e_input[82]), .B(n30243), .Z(n30246) );
  XNOR U30332 ( .A(n23616), .B(n30243), .Z(n30245) );
  XOR U30333 ( .A(n30247), .B(n30248), .Z(n23616) );
  XOR U30334 ( .A(n30249), .B(n30250), .Z(n30243) );
  AND U30335 ( .A(n30251), .B(n30252), .Z(n30250) );
  XOR U30336 ( .A(e_input[81]), .B(n30249), .Z(n30252) );
  XNOR U30337 ( .A(n23628), .B(n30249), .Z(n30251) );
  XOR U30338 ( .A(n30253), .B(n30254), .Z(n23628) );
  XOR U30339 ( .A(n30255), .B(n30256), .Z(n30249) );
  AND U30340 ( .A(n30257), .B(n30258), .Z(n30256) );
  XOR U30341 ( .A(e_input[80]), .B(n30255), .Z(n30258) );
  XNOR U30342 ( .A(n23640), .B(n30255), .Z(n30257) );
  XOR U30343 ( .A(n30259), .B(n30260), .Z(n23640) );
  XOR U30344 ( .A(n30261), .B(n30262), .Z(n30255) );
  AND U30345 ( .A(n30263), .B(n30264), .Z(n30262) );
  XOR U30346 ( .A(e_input[79]), .B(n30261), .Z(n30264) );
  XNOR U30347 ( .A(n23652), .B(n30261), .Z(n30263) );
  XOR U30348 ( .A(n30265), .B(n30266), .Z(n23652) );
  XOR U30349 ( .A(n30267), .B(n30268), .Z(n30261) );
  AND U30350 ( .A(n30269), .B(n30270), .Z(n30268) );
  XOR U30351 ( .A(e_input[78]), .B(n30267), .Z(n30270) );
  XNOR U30352 ( .A(n23664), .B(n30267), .Z(n30269) );
  XOR U30353 ( .A(n30271), .B(n30272), .Z(n23664) );
  XOR U30354 ( .A(n30273), .B(n30274), .Z(n30267) );
  AND U30355 ( .A(n30275), .B(n30276), .Z(n30274) );
  XOR U30356 ( .A(e_input[77]), .B(n30273), .Z(n30276) );
  XNOR U30357 ( .A(n23676), .B(n30273), .Z(n30275) );
  XOR U30358 ( .A(n30277), .B(n30278), .Z(n23676) );
  XOR U30359 ( .A(n30279), .B(n30280), .Z(n30273) );
  AND U30360 ( .A(n30281), .B(n30282), .Z(n30280) );
  XOR U30361 ( .A(e_input[76]), .B(n30279), .Z(n30282) );
  XNOR U30362 ( .A(n23688), .B(n30279), .Z(n30281) );
  XOR U30363 ( .A(n30283), .B(n30284), .Z(n23688) );
  XOR U30364 ( .A(n30285), .B(n30286), .Z(n30279) );
  AND U30365 ( .A(n30287), .B(n30288), .Z(n30286) );
  XOR U30366 ( .A(e_input[75]), .B(n30285), .Z(n30288) );
  XNOR U30367 ( .A(n23700), .B(n30285), .Z(n30287) );
  XOR U30368 ( .A(n30289), .B(n30290), .Z(n23700) );
  XOR U30369 ( .A(n30291), .B(n30292), .Z(n30285) );
  AND U30370 ( .A(n30293), .B(n30294), .Z(n30292) );
  XOR U30371 ( .A(e_input[74]), .B(n30291), .Z(n30294) );
  XNOR U30372 ( .A(n23712), .B(n30291), .Z(n30293) );
  XOR U30373 ( .A(n30295), .B(n30296), .Z(n23712) );
  XOR U30374 ( .A(n30297), .B(n30298), .Z(n30291) );
  AND U30375 ( .A(n30299), .B(n30300), .Z(n30298) );
  XOR U30376 ( .A(e_input[73]), .B(n30297), .Z(n30300) );
  XNOR U30377 ( .A(n23724), .B(n30297), .Z(n30299) );
  XOR U30378 ( .A(n30301), .B(n30302), .Z(n23724) );
  XOR U30379 ( .A(n30303), .B(n30304), .Z(n30297) );
  AND U30380 ( .A(n30305), .B(n30306), .Z(n30304) );
  XOR U30381 ( .A(e_input[72]), .B(n30303), .Z(n30306) );
  XNOR U30382 ( .A(n23736), .B(n30303), .Z(n30305) );
  XOR U30383 ( .A(n30307), .B(n30308), .Z(n23736) );
  XOR U30384 ( .A(n30309), .B(n30310), .Z(n30303) );
  AND U30385 ( .A(n30311), .B(n30312), .Z(n30310) );
  XOR U30386 ( .A(e_input[71]), .B(n30309), .Z(n30312) );
  XNOR U30387 ( .A(n23748), .B(n30309), .Z(n30311) );
  XOR U30388 ( .A(n30313), .B(n30314), .Z(n23748) );
  XOR U30389 ( .A(n30315), .B(n30316), .Z(n30309) );
  AND U30390 ( .A(n30317), .B(n30318), .Z(n30316) );
  XOR U30391 ( .A(e_input[70]), .B(n30315), .Z(n30318) );
  XNOR U30392 ( .A(n23760), .B(n30315), .Z(n30317) );
  XOR U30393 ( .A(n30319), .B(n30320), .Z(n23760) );
  XOR U30394 ( .A(n30321), .B(n30322), .Z(n30315) );
  AND U30395 ( .A(n30323), .B(n30324), .Z(n30322) );
  XOR U30396 ( .A(e_input[69]), .B(n30321), .Z(n30324) );
  XNOR U30397 ( .A(n23772), .B(n30321), .Z(n30323) );
  XOR U30398 ( .A(n30325), .B(n30326), .Z(n23772) );
  XOR U30399 ( .A(n30327), .B(n30328), .Z(n30321) );
  AND U30400 ( .A(n30329), .B(n30330), .Z(n30328) );
  XOR U30401 ( .A(e_input[68]), .B(n30327), .Z(n30330) );
  XNOR U30402 ( .A(n23784), .B(n30327), .Z(n30329) );
  XOR U30403 ( .A(n30331), .B(n30332), .Z(n23784) );
  XOR U30404 ( .A(n30333), .B(n30334), .Z(n30327) );
  AND U30405 ( .A(n30335), .B(n30336), .Z(n30334) );
  XOR U30406 ( .A(e_input[67]), .B(n30333), .Z(n30336) );
  XNOR U30407 ( .A(n23796), .B(n30333), .Z(n30335) );
  XOR U30408 ( .A(n30337), .B(n30338), .Z(n23796) );
  XOR U30409 ( .A(n30339), .B(n30340), .Z(n30333) );
  AND U30410 ( .A(n30341), .B(n30342), .Z(n30340) );
  XOR U30411 ( .A(e_input[66]), .B(n30339), .Z(n30342) );
  XNOR U30412 ( .A(n23808), .B(n30339), .Z(n30341) );
  XOR U30413 ( .A(n30343), .B(n30344), .Z(n23808) );
  XOR U30414 ( .A(n30345), .B(n30346), .Z(n30339) );
  AND U30415 ( .A(n30347), .B(n30348), .Z(n30346) );
  XOR U30416 ( .A(e_input[65]), .B(n30345), .Z(n30348) );
  XNOR U30417 ( .A(n23820), .B(n30345), .Z(n30347) );
  XOR U30418 ( .A(n30349), .B(n30350), .Z(n23820) );
  XOR U30419 ( .A(n30351), .B(n30352), .Z(n30345) );
  AND U30420 ( .A(n30353), .B(n30354), .Z(n30352) );
  XOR U30421 ( .A(e_input[64]), .B(n30351), .Z(n30354) );
  XNOR U30422 ( .A(n23832), .B(n30351), .Z(n30353) );
  XOR U30423 ( .A(n30355), .B(n30356), .Z(n23832) );
  XOR U30424 ( .A(n30357), .B(n30358), .Z(n30351) );
  AND U30425 ( .A(n30359), .B(n30360), .Z(n30358) );
  XOR U30426 ( .A(e_input[63]), .B(n30357), .Z(n30360) );
  XNOR U30427 ( .A(n23844), .B(n30357), .Z(n30359) );
  XOR U30428 ( .A(n30361), .B(n30362), .Z(n23844) );
  XOR U30429 ( .A(n30363), .B(n30364), .Z(n30357) );
  AND U30430 ( .A(n30365), .B(n30366), .Z(n30364) );
  XOR U30431 ( .A(e_input[62]), .B(n30363), .Z(n30366) );
  XNOR U30432 ( .A(n23856), .B(n30363), .Z(n30365) );
  XOR U30433 ( .A(n30367), .B(n30368), .Z(n23856) );
  XOR U30434 ( .A(n30369), .B(n30370), .Z(n30363) );
  AND U30435 ( .A(n30371), .B(n30372), .Z(n30370) );
  XOR U30436 ( .A(e_input[61]), .B(n30369), .Z(n30372) );
  XNOR U30437 ( .A(n23868), .B(n30369), .Z(n30371) );
  XOR U30438 ( .A(n30373), .B(n30374), .Z(n23868) );
  XOR U30439 ( .A(n30375), .B(n30376), .Z(n30369) );
  AND U30440 ( .A(n30377), .B(n30378), .Z(n30376) );
  XOR U30441 ( .A(e_input[60]), .B(n30375), .Z(n30378) );
  XNOR U30442 ( .A(n23880), .B(n30375), .Z(n30377) );
  XOR U30443 ( .A(n30379), .B(n30380), .Z(n23880) );
  XOR U30444 ( .A(n30381), .B(n30382), .Z(n30375) );
  AND U30445 ( .A(n30383), .B(n30384), .Z(n30382) );
  XOR U30446 ( .A(e_input[59]), .B(n30381), .Z(n30384) );
  XNOR U30447 ( .A(n23892), .B(n30381), .Z(n30383) );
  XOR U30448 ( .A(n30385), .B(n30386), .Z(n23892) );
  XOR U30449 ( .A(n30387), .B(n30388), .Z(n30381) );
  AND U30450 ( .A(n30389), .B(n30390), .Z(n30388) );
  XOR U30451 ( .A(e_input[58]), .B(n30387), .Z(n30390) );
  XNOR U30452 ( .A(n23904), .B(n30387), .Z(n30389) );
  XOR U30453 ( .A(n30391), .B(n30392), .Z(n23904) );
  XOR U30454 ( .A(n30393), .B(n30394), .Z(n30387) );
  AND U30455 ( .A(n30395), .B(n30396), .Z(n30394) );
  XOR U30456 ( .A(e_input[57]), .B(n30393), .Z(n30396) );
  XNOR U30457 ( .A(n23916), .B(n30393), .Z(n30395) );
  XOR U30458 ( .A(n30397), .B(n30398), .Z(n23916) );
  XOR U30459 ( .A(n30399), .B(n30400), .Z(n30393) );
  AND U30460 ( .A(n30401), .B(n30402), .Z(n30400) );
  XOR U30461 ( .A(e_input[56]), .B(n30399), .Z(n30402) );
  XNOR U30462 ( .A(n23928), .B(n30399), .Z(n30401) );
  XOR U30463 ( .A(n30403), .B(n30404), .Z(n23928) );
  XOR U30464 ( .A(n30405), .B(n30406), .Z(n30399) );
  AND U30465 ( .A(n30407), .B(n30408), .Z(n30406) );
  XOR U30466 ( .A(e_input[55]), .B(n30405), .Z(n30408) );
  XNOR U30467 ( .A(n23940), .B(n30405), .Z(n30407) );
  XOR U30468 ( .A(n30409), .B(n30410), .Z(n23940) );
  XOR U30469 ( .A(n30411), .B(n30412), .Z(n30405) );
  AND U30470 ( .A(n30413), .B(n30414), .Z(n30412) );
  XOR U30471 ( .A(e_input[54]), .B(n30411), .Z(n30414) );
  XNOR U30472 ( .A(n23952), .B(n30411), .Z(n30413) );
  XOR U30473 ( .A(n30415), .B(n30416), .Z(n23952) );
  XOR U30474 ( .A(n30417), .B(n30418), .Z(n30411) );
  AND U30475 ( .A(n30419), .B(n30420), .Z(n30418) );
  XOR U30476 ( .A(e_input[53]), .B(n30417), .Z(n30420) );
  XNOR U30477 ( .A(n23964), .B(n30417), .Z(n30419) );
  XOR U30478 ( .A(n30421), .B(n30422), .Z(n23964) );
  XOR U30479 ( .A(n30423), .B(n30424), .Z(n30417) );
  AND U30480 ( .A(n30425), .B(n30426), .Z(n30424) );
  XOR U30481 ( .A(e_input[52]), .B(n30423), .Z(n30426) );
  XNOR U30482 ( .A(n23976), .B(n30423), .Z(n30425) );
  XOR U30483 ( .A(n30427), .B(n30428), .Z(n23976) );
  XOR U30484 ( .A(n30429), .B(n30430), .Z(n30423) );
  AND U30485 ( .A(n30431), .B(n30432), .Z(n30430) );
  XOR U30486 ( .A(e_input[51]), .B(n30429), .Z(n30432) );
  XNOR U30487 ( .A(n23988), .B(n30429), .Z(n30431) );
  XOR U30488 ( .A(n30433), .B(n30434), .Z(n23988) );
  XOR U30489 ( .A(n30435), .B(n30436), .Z(n30429) );
  AND U30490 ( .A(n30437), .B(n30438), .Z(n30436) );
  XOR U30491 ( .A(e_input[50]), .B(n30435), .Z(n30438) );
  XNOR U30492 ( .A(n24000), .B(n30435), .Z(n30437) );
  XOR U30493 ( .A(n30439), .B(n30440), .Z(n24000) );
  XOR U30494 ( .A(n30441), .B(n30442), .Z(n30435) );
  AND U30495 ( .A(n30443), .B(n30444), .Z(n30442) );
  XOR U30496 ( .A(e_input[49]), .B(n30441), .Z(n30444) );
  XNOR U30497 ( .A(n24012), .B(n30441), .Z(n30443) );
  XOR U30498 ( .A(n30445), .B(n30446), .Z(n24012) );
  XOR U30499 ( .A(n30447), .B(n30448), .Z(n30441) );
  AND U30500 ( .A(n30449), .B(n30450), .Z(n30448) );
  XOR U30501 ( .A(e_input[48]), .B(n30447), .Z(n30450) );
  XNOR U30502 ( .A(n24024), .B(n30447), .Z(n30449) );
  XOR U30503 ( .A(n30451), .B(n30452), .Z(n24024) );
  XOR U30504 ( .A(n30453), .B(n30454), .Z(n30447) );
  AND U30505 ( .A(n30455), .B(n30456), .Z(n30454) );
  XOR U30506 ( .A(e_input[47]), .B(n30453), .Z(n30456) );
  XNOR U30507 ( .A(n24036), .B(n30453), .Z(n30455) );
  XOR U30508 ( .A(n30457), .B(n30458), .Z(n24036) );
  XOR U30509 ( .A(n30459), .B(n30460), .Z(n30453) );
  AND U30510 ( .A(n30461), .B(n30462), .Z(n30460) );
  XOR U30511 ( .A(e_input[46]), .B(n30459), .Z(n30462) );
  XNOR U30512 ( .A(n24048), .B(n30459), .Z(n30461) );
  XOR U30513 ( .A(n30463), .B(n30464), .Z(n24048) );
  XOR U30514 ( .A(n30465), .B(n30466), .Z(n30459) );
  AND U30515 ( .A(n30467), .B(n30468), .Z(n30466) );
  XOR U30516 ( .A(e_input[45]), .B(n30465), .Z(n30468) );
  XNOR U30517 ( .A(n24060), .B(n30465), .Z(n30467) );
  XOR U30518 ( .A(n30469), .B(n30470), .Z(n24060) );
  XOR U30519 ( .A(n30471), .B(n30472), .Z(n30465) );
  AND U30520 ( .A(n30473), .B(n30474), .Z(n30472) );
  XOR U30521 ( .A(e_input[44]), .B(n30471), .Z(n30474) );
  XNOR U30522 ( .A(n24072), .B(n30471), .Z(n30473) );
  XOR U30523 ( .A(n30475), .B(n30476), .Z(n24072) );
  XOR U30524 ( .A(n30477), .B(n30478), .Z(n30471) );
  AND U30525 ( .A(n30479), .B(n30480), .Z(n30478) );
  XOR U30526 ( .A(e_input[43]), .B(n30477), .Z(n30480) );
  XNOR U30527 ( .A(n24084), .B(n30477), .Z(n30479) );
  XOR U30528 ( .A(n30481), .B(n30482), .Z(n24084) );
  XOR U30529 ( .A(n30483), .B(n30484), .Z(n30477) );
  AND U30530 ( .A(n30485), .B(n30486), .Z(n30484) );
  XOR U30531 ( .A(e_input[42]), .B(n30483), .Z(n30486) );
  XNOR U30532 ( .A(n24096), .B(n30483), .Z(n30485) );
  XOR U30533 ( .A(n30487), .B(n30488), .Z(n24096) );
  XOR U30534 ( .A(n30489), .B(n30490), .Z(n30483) );
  AND U30535 ( .A(n30491), .B(n30492), .Z(n30490) );
  XOR U30536 ( .A(e_input[41]), .B(n30489), .Z(n30492) );
  XNOR U30537 ( .A(n24108), .B(n30489), .Z(n30491) );
  XOR U30538 ( .A(n30493), .B(n30494), .Z(n24108) );
  XOR U30539 ( .A(n30495), .B(n30496), .Z(n30489) );
  AND U30540 ( .A(n30497), .B(n30498), .Z(n30496) );
  XOR U30541 ( .A(e_input[40]), .B(n30495), .Z(n30498) );
  XNOR U30542 ( .A(n24120), .B(n30495), .Z(n30497) );
  XOR U30543 ( .A(n30499), .B(n30500), .Z(n24120) );
  XOR U30544 ( .A(n30501), .B(n30502), .Z(n30495) );
  AND U30545 ( .A(n30503), .B(n30504), .Z(n30502) );
  XOR U30546 ( .A(e_input[39]), .B(n30501), .Z(n30504) );
  XNOR U30547 ( .A(n24132), .B(n30501), .Z(n30503) );
  XOR U30548 ( .A(n30505), .B(n30506), .Z(n24132) );
  XOR U30549 ( .A(n30507), .B(n30508), .Z(n30501) );
  AND U30550 ( .A(n30509), .B(n30510), .Z(n30508) );
  XOR U30551 ( .A(e_input[38]), .B(n30507), .Z(n30510) );
  XNOR U30552 ( .A(n24144), .B(n30507), .Z(n30509) );
  XOR U30553 ( .A(n30511), .B(n30512), .Z(n24144) );
  XOR U30554 ( .A(n30513), .B(n30514), .Z(n30507) );
  AND U30555 ( .A(n30515), .B(n30516), .Z(n30514) );
  XOR U30556 ( .A(e_input[37]), .B(n30513), .Z(n30516) );
  XNOR U30557 ( .A(n24156), .B(n30513), .Z(n30515) );
  XOR U30558 ( .A(n30517), .B(n30518), .Z(n24156) );
  XOR U30559 ( .A(n30519), .B(n30520), .Z(n30513) );
  AND U30560 ( .A(n30521), .B(n30522), .Z(n30520) );
  XOR U30561 ( .A(e_input[36]), .B(n30519), .Z(n30522) );
  XNOR U30562 ( .A(n24168), .B(n30519), .Z(n30521) );
  XOR U30563 ( .A(n30523), .B(n30524), .Z(n24168) );
  XOR U30564 ( .A(n30525), .B(n30526), .Z(n30519) );
  AND U30565 ( .A(n30527), .B(n30528), .Z(n30526) );
  XOR U30566 ( .A(e_input[35]), .B(n30525), .Z(n30528) );
  XNOR U30567 ( .A(n24180), .B(n30525), .Z(n30527) );
  XOR U30568 ( .A(n30529), .B(n30530), .Z(n24180) );
  XOR U30569 ( .A(n30531), .B(n30532), .Z(n30525) );
  AND U30570 ( .A(n30533), .B(n30534), .Z(n30532) );
  XOR U30571 ( .A(e_input[34]), .B(n30531), .Z(n30534) );
  XNOR U30572 ( .A(n24192), .B(n30531), .Z(n30533) );
  XOR U30573 ( .A(n30535), .B(n30536), .Z(n24192) );
  XOR U30574 ( .A(n30537), .B(n30538), .Z(n30531) );
  AND U30575 ( .A(n30539), .B(n30540), .Z(n30538) );
  XOR U30576 ( .A(e_input[33]), .B(n30537), .Z(n30540) );
  XNOR U30577 ( .A(n24204), .B(n30537), .Z(n30539) );
  XOR U30578 ( .A(n30541), .B(n30542), .Z(n24204) );
  XOR U30579 ( .A(n30543), .B(n30544), .Z(n30537) );
  AND U30580 ( .A(n30545), .B(n30546), .Z(n30544) );
  XOR U30581 ( .A(e_input[32]), .B(n30543), .Z(n30546) );
  XNOR U30582 ( .A(n24216), .B(n30543), .Z(n30545) );
  XOR U30583 ( .A(n30547), .B(n30548), .Z(n24216) );
  XOR U30584 ( .A(n30549), .B(n30550), .Z(n30543) );
  AND U30585 ( .A(n30551), .B(n30552), .Z(n30550) );
  XOR U30586 ( .A(e_input[31]), .B(n30549), .Z(n30552) );
  XNOR U30587 ( .A(n24228), .B(n30549), .Z(n30551) );
  XOR U30588 ( .A(n30553), .B(n30554), .Z(n24228) );
  XOR U30589 ( .A(n30555), .B(n30556), .Z(n30549) );
  AND U30590 ( .A(n30557), .B(n30558), .Z(n30556) );
  XOR U30591 ( .A(e_input[30]), .B(n30555), .Z(n30558) );
  XNOR U30592 ( .A(n24240), .B(n30555), .Z(n30557) );
  XOR U30593 ( .A(n30559), .B(n30560), .Z(n24240) );
  XOR U30594 ( .A(n30561), .B(n30562), .Z(n30555) );
  AND U30595 ( .A(n30563), .B(n30564), .Z(n30562) );
  XOR U30596 ( .A(e_input[29]), .B(n30561), .Z(n30564) );
  XNOR U30597 ( .A(n24252), .B(n30561), .Z(n30563) );
  XOR U30598 ( .A(n30565), .B(n30566), .Z(n24252) );
  XOR U30599 ( .A(n30567), .B(n30568), .Z(n30561) );
  AND U30600 ( .A(n30569), .B(n30570), .Z(n30568) );
  XOR U30601 ( .A(e_input[28]), .B(n30567), .Z(n30570) );
  XNOR U30602 ( .A(n24264), .B(n30567), .Z(n30569) );
  XOR U30603 ( .A(n30571), .B(n30572), .Z(n24264) );
  XOR U30604 ( .A(n30573), .B(n30574), .Z(n30567) );
  AND U30605 ( .A(n30575), .B(n30576), .Z(n30574) );
  XOR U30606 ( .A(e_input[27]), .B(n30573), .Z(n30576) );
  XNOR U30607 ( .A(n24276), .B(n30573), .Z(n30575) );
  XOR U30608 ( .A(n30577), .B(n30578), .Z(n24276) );
  XOR U30609 ( .A(n30579), .B(n30580), .Z(n30573) );
  AND U30610 ( .A(n30581), .B(n30582), .Z(n30580) );
  XOR U30611 ( .A(e_input[26]), .B(n30579), .Z(n30582) );
  XNOR U30612 ( .A(n24288), .B(n30579), .Z(n30581) );
  XOR U30613 ( .A(n30583), .B(n30584), .Z(n24288) );
  XOR U30614 ( .A(n30585), .B(n30586), .Z(n30579) );
  AND U30615 ( .A(n30587), .B(n30588), .Z(n30586) );
  XOR U30616 ( .A(e_input[25]), .B(n30585), .Z(n30588) );
  XNOR U30617 ( .A(n24300), .B(n30585), .Z(n30587) );
  XOR U30618 ( .A(n30589), .B(n30590), .Z(n24300) );
  XOR U30619 ( .A(n30591), .B(n30592), .Z(n30585) );
  AND U30620 ( .A(n30593), .B(n30594), .Z(n30592) );
  XOR U30621 ( .A(e_input[24]), .B(n30591), .Z(n30594) );
  XNOR U30622 ( .A(n24312), .B(n30591), .Z(n30593) );
  XOR U30623 ( .A(n30595), .B(n30596), .Z(n24312) );
  XOR U30624 ( .A(n30597), .B(n30598), .Z(n30591) );
  AND U30625 ( .A(n30599), .B(n30600), .Z(n30598) );
  XOR U30626 ( .A(e_input[23]), .B(n30597), .Z(n30600) );
  XNOR U30627 ( .A(n24324), .B(n30597), .Z(n30599) );
  XOR U30628 ( .A(n30601), .B(n30602), .Z(n24324) );
  XOR U30629 ( .A(n30603), .B(n30604), .Z(n30597) );
  AND U30630 ( .A(n30605), .B(n30606), .Z(n30604) );
  XOR U30631 ( .A(e_input[22]), .B(n30603), .Z(n30606) );
  XNOR U30632 ( .A(n24336), .B(n30603), .Z(n30605) );
  XOR U30633 ( .A(n30607), .B(n30608), .Z(n24336) );
  XOR U30634 ( .A(n30609), .B(n30610), .Z(n30603) );
  AND U30635 ( .A(n30611), .B(n30612), .Z(n30610) );
  XOR U30636 ( .A(e_input[21]), .B(n30609), .Z(n30612) );
  XNOR U30637 ( .A(n24348), .B(n30609), .Z(n30611) );
  XOR U30638 ( .A(n30613), .B(n30614), .Z(n24348) );
  XOR U30639 ( .A(n30615), .B(n30616), .Z(n30609) );
  AND U30640 ( .A(n30617), .B(n30618), .Z(n30616) );
  XOR U30641 ( .A(e_input[20]), .B(n30615), .Z(n30618) );
  XNOR U30642 ( .A(n24360), .B(n30615), .Z(n30617) );
  XOR U30643 ( .A(n30619), .B(n30620), .Z(n24360) );
  XOR U30644 ( .A(n30621), .B(n30622), .Z(n30615) );
  AND U30645 ( .A(n30623), .B(n30624), .Z(n30622) );
  XOR U30646 ( .A(e_input[19]), .B(n30621), .Z(n30624) );
  XNOR U30647 ( .A(n24372), .B(n30621), .Z(n30623) );
  XOR U30648 ( .A(n30625), .B(n30626), .Z(n24372) );
  XOR U30649 ( .A(n30627), .B(n30628), .Z(n30621) );
  AND U30650 ( .A(n30629), .B(n30630), .Z(n30628) );
  XOR U30651 ( .A(e_input[18]), .B(n30627), .Z(n30630) );
  XNOR U30652 ( .A(n24384), .B(n30627), .Z(n30629) );
  XOR U30653 ( .A(n30631), .B(n30632), .Z(n24384) );
  XOR U30654 ( .A(n30633), .B(n30634), .Z(n30627) );
  AND U30655 ( .A(n30635), .B(n30636), .Z(n30634) );
  XOR U30656 ( .A(e_input[17]), .B(n30633), .Z(n30636) );
  XNOR U30657 ( .A(n24396), .B(n30633), .Z(n30635) );
  XOR U30658 ( .A(n30637), .B(n30638), .Z(n24396) );
  XOR U30659 ( .A(n30639), .B(n30640), .Z(n30633) );
  AND U30660 ( .A(n30641), .B(n30642), .Z(n30640) );
  XOR U30661 ( .A(e_input[16]), .B(n30639), .Z(n30642) );
  XNOR U30662 ( .A(n24408), .B(n30639), .Z(n30641) );
  XOR U30663 ( .A(n30643), .B(n30644), .Z(n24408) );
  XOR U30664 ( .A(n30645), .B(n30646), .Z(n30639) );
  AND U30665 ( .A(n30647), .B(n30648), .Z(n30646) );
  XOR U30666 ( .A(e_input[15]), .B(n30645), .Z(n30648) );
  XNOR U30667 ( .A(n24420), .B(n30645), .Z(n30647) );
  XOR U30668 ( .A(n30649), .B(n30650), .Z(n24420) );
  XOR U30669 ( .A(n30651), .B(n30652), .Z(n30645) );
  AND U30670 ( .A(n30653), .B(n30654), .Z(n30652) );
  XOR U30671 ( .A(e_input[14]), .B(n30651), .Z(n30654) );
  XNOR U30672 ( .A(n24432), .B(n30651), .Z(n30653) );
  XOR U30673 ( .A(n30655), .B(n30656), .Z(n24432) );
  XOR U30674 ( .A(n30657), .B(n30658), .Z(n30651) );
  AND U30675 ( .A(n30659), .B(n30660), .Z(n30658) );
  XOR U30676 ( .A(e_input[13]), .B(n30657), .Z(n30660) );
  XNOR U30677 ( .A(n24444), .B(n30657), .Z(n30659) );
  XOR U30678 ( .A(n30661), .B(n30662), .Z(n24444) );
  XOR U30679 ( .A(n30663), .B(n30664), .Z(n30657) );
  AND U30680 ( .A(n30665), .B(n30666), .Z(n30664) );
  XOR U30681 ( .A(e_input[12]), .B(n30663), .Z(n30666) );
  XNOR U30682 ( .A(n24456), .B(n30663), .Z(n30665) );
  XOR U30683 ( .A(n30667), .B(n30668), .Z(n24456) );
  XOR U30684 ( .A(n30669), .B(n30670), .Z(n30663) );
  AND U30685 ( .A(n30671), .B(n30672), .Z(n30670) );
  XOR U30686 ( .A(e_input[11]), .B(n30669), .Z(n30672) );
  XNOR U30687 ( .A(n24468), .B(n30669), .Z(n30671) );
  XOR U30688 ( .A(n30673), .B(n30674), .Z(n24468) );
  XOR U30689 ( .A(n30675), .B(n30676), .Z(n30669) );
  AND U30690 ( .A(n30677), .B(n30678), .Z(n30676) );
  XOR U30691 ( .A(e_input[10]), .B(n30675), .Z(n30678) );
  XNOR U30692 ( .A(n24480), .B(n30675), .Z(n30677) );
  XOR U30693 ( .A(n30679), .B(n30680), .Z(n24480) );
  XOR U30694 ( .A(n30681), .B(n30682), .Z(n30675) );
  AND U30695 ( .A(n30683), .B(n30684), .Z(n30682) );
  XOR U30696 ( .A(e_input[9]), .B(n30681), .Z(n30684) );
  XNOR U30697 ( .A(n24492), .B(n30681), .Z(n30683) );
  XOR U30698 ( .A(n30685), .B(n30686), .Z(n24492) );
  XOR U30699 ( .A(n30687), .B(n30688), .Z(n30681) );
  AND U30700 ( .A(n30689), .B(n30690), .Z(n30688) );
  XOR U30701 ( .A(e_input[8]), .B(n30687), .Z(n30690) );
  XNOR U30702 ( .A(n24504), .B(n30687), .Z(n30689) );
  XOR U30703 ( .A(n30691), .B(n30692), .Z(n24504) );
  XOR U30704 ( .A(n30693), .B(n30694), .Z(n30687) );
  AND U30705 ( .A(n30695), .B(n30696), .Z(n30694) );
  XOR U30706 ( .A(e_input[7]), .B(n30693), .Z(n30696) );
  XNOR U30707 ( .A(n24516), .B(n30693), .Z(n30695) );
  XOR U30708 ( .A(n30697), .B(n30698), .Z(n24516) );
  XOR U30709 ( .A(n30699), .B(n30700), .Z(n30693) );
  AND U30710 ( .A(n30701), .B(n30702), .Z(n30700) );
  XOR U30711 ( .A(e_input[6]), .B(n30699), .Z(n30702) );
  XNOR U30712 ( .A(n24528), .B(n30699), .Z(n30701) );
  XOR U30713 ( .A(n30703), .B(n30704), .Z(n24528) );
  XOR U30714 ( .A(n30705), .B(n30706), .Z(n30699) );
  AND U30715 ( .A(n30707), .B(n30708), .Z(n30706) );
  XOR U30716 ( .A(e_input[5]), .B(n30705), .Z(n30708) );
  XNOR U30717 ( .A(n24540), .B(n30705), .Z(n30707) );
  XOR U30718 ( .A(n30709), .B(n30710), .Z(n24540) );
  XOR U30719 ( .A(n30711), .B(n30712), .Z(n30705) );
  AND U30720 ( .A(n30713), .B(n30714), .Z(n30712) );
  XOR U30721 ( .A(e_input[4]), .B(n30711), .Z(n30714) );
  XNOR U30722 ( .A(n24552), .B(n30711), .Z(n30713) );
  XOR U30723 ( .A(n30715), .B(n30716), .Z(n24552) );
  XOR U30724 ( .A(n30717), .B(n30718), .Z(n30711) );
  AND U30725 ( .A(n30719), .B(n30720), .Z(n30718) );
  XOR U30726 ( .A(e_input[3]), .B(n30717), .Z(n30720) );
  XNOR U30727 ( .A(n24564), .B(n30717), .Z(n30719) );
  XOR U30728 ( .A(n30721), .B(n30722), .Z(n24564) );
  XNOR U30729 ( .A(n30723), .B(n30724), .Z(n30717) );
  AND U30730 ( .A(n30725), .B(n30726), .Z(n30724) );
  XNOR U30731 ( .A(e_input[2]), .B(n30723), .Z(n30726) );
  XNOR U30732 ( .A(n24576), .B(n30723), .Z(n30725) );
  XOR U30733 ( .A(n30727), .B(n30728), .Z(n24576) );
  XOR U30734 ( .A(n30729), .B(n30730), .Z(n30723) );
  NAND U30735 ( .A(n30731), .B(n30732), .Z(n30729) );
  XNOR U30736 ( .A(e_input[1]), .B(n30733), .Z(n30732) );
  IV U30737 ( .A(n30730), .Z(n30733) );
  XNOR U30738 ( .A(n24587), .B(n30730), .Z(n30731) );
  ANDN U30739 ( .A(e_input[0]), .B(n24588), .Z(n30730) );
  XNOR U30740 ( .A(n30734), .B(\modmult_1/zin[0][0] ), .Z(n24587) );
  XOR U30741 ( .A(n30735), .B(n30736), .Z(n12306) );
  XOR U30742 ( .A(n30737), .B(\modmult_1/zin[0][1024] ), .Z(n30735) );
  NAND U30743 ( .A(n30736), .B(n12312), .Z(n30737) );
  XNOR U30744 ( .A(n30738), .B(\modmult_1/zin[0][1023] ), .Z(n12312) );
  IV U30745 ( .A(n30736), .Z(n30738) );
  XOR U30746 ( .A(n30739), .B(n30740), .Z(n30736) );
  ANDN U30747 ( .A(n30741), .B(n24602), .Z(n30740) );
  XOR U30748 ( .A(n30742), .B(\modmult_1/zin[0][1022] ), .Z(n24602) );
  IV U30749 ( .A(n30739), .Z(n30742) );
  XNOR U30750 ( .A(n30739), .B(n24601), .Z(n30741) );
  XOR U30751 ( .A(n30743), .B(n30744), .Z(n24601) );
  ANDN U30752 ( .A(\modmult_1/xin[1023] ), .B(n30743), .Z(n30744) );
  XOR U30753 ( .A(n30745), .B(g_input[1023]), .Z(n30743) );
  NAND U30754 ( .A(n30746), .B(mul_pow), .Z(n30745) );
  XOR U30755 ( .A(g_input[1023]), .B(creg[1023]), .Z(n30746) );
  XOR U30756 ( .A(n30747), .B(n30748), .Z(n30739) );
  ANDN U30757 ( .A(n30749), .B(n24608), .Z(n30748) );
  XOR U30758 ( .A(n30750), .B(\modmult_1/zin[0][1021] ), .Z(n24608) );
  IV U30759 ( .A(n30747), .Z(n30750) );
  XNOR U30760 ( .A(n30747), .B(n24607), .Z(n30749) );
  XOR U30761 ( .A(n30751), .B(n30752), .Z(n24607) );
  AND U30762 ( .A(\modmult_1/xin[1023] ), .B(n30753), .Z(n30752) );
  IV U30763 ( .A(n30751), .Z(n30753) );
  XOR U30764 ( .A(n30754), .B(g_input[1022]), .Z(n30751) );
  NAND U30765 ( .A(n30755), .B(mul_pow), .Z(n30754) );
  XOR U30766 ( .A(g_input[1022]), .B(creg[1022]), .Z(n30755) );
  XOR U30767 ( .A(n30756), .B(n30757), .Z(n30747) );
  ANDN U30768 ( .A(n30758), .B(n24614), .Z(n30757) );
  XOR U30769 ( .A(n30759), .B(\modmult_1/zin[0][1020] ), .Z(n24614) );
  IV U30770 ( .A(n30756), .Z(n30759) );
  XNOR U30771 ( .A(n30756), .B(n24613), .Z(n30758) );
  XOR U30772 ( .A(n30760), .B(n30761), .Z(n24613) );
  AND U30773 ( .A(\modmult_1/xin[1023] ), .B(n30762), .Z(n30761) );
  IV U30774 ( .A(n30760), .Z(n30762) );
  XOR U30775 ( .A(n30763), .B(g_input[1021]), .Z(n30760) );
  NAND U30776 ( .A(n30764), .B(mul_pow), .Z(n30763) );
  XOR U30777 ( .A(g_input[1021]), .B(creg[1021]), .Z(n30764) );
  XOR U30778 ( .A(n30765), .B(n30766), .Z(n30756) );
  ANDN U30779 ( .A(n30767), .B(n24620), .Z(n30766) );
  XOR U30780 ( .A(n30768), .B(\modmult_1/zin[0][1019] ), .Z(n24620) );
  IV U30781 ( .A(n30765), .Z(n30768) );
  XNOR U30782 ( .A(n30765), .B(n24619), .Z(n30767) );
  XOR U30783 ( .A(n30769), .B(n30770), .Z(n24619) );
  AND U30784 ( .A(\modmult_1/xin[1023] ), .B(n30771), .Z(n30770) );
  IV U30785 ( .A(n30769), .Z(n30771) );
  XOR U30786 ( .A(n30772), .B(g_input[1020]), .Z(n30769) );
  NAND U30787 ( .A(n30773), .B(mul_pow), .Z(n30772) );
  XOR U30788 ( .A(g_input[1020]), .B(creg[1020]), .Z(n30773) );
  XOR U30789 ( .A(n30774), .B(n30775), .Z(n30765) );
  ANDN U30790 ( .A(n30776), .B(n24626), .Z(n30775) );
  XOR U30791 ( .A(n30777), .B(\modmult_1/zin[0][1018] ), .Z(n24626) );
  IV U30792 ( .A(n30774), .Z(n30777) );
  XNOR U30793 ( .A(n30774), .B(n24625), .Z(n30776) );
  XOR U30794 ( .A(n30778), .B(n30779), .Z(n24625) );
  AND U30795 ( .A(\modmult_1/xin[1023] ), .B(n30780), .Z(n30779) );
  IV U30796 ( .A(n30778), .Z(n30780) );
  XOR U30797 ( .A(n30781), .B(g_input[1019]), .Z(n30778) );
  NAND U30798 ( .A(n30782), .B(mul_pow), .Z(n30781) );
  XOR U30799 ( .A(g_input[1019]), .B(creg[1019]), .Z(n30782) );
  XOR U30800 ( .A(n30783), .B(n30784), .Z(n30774) );
  ANDN U30801 ( .A(n30785), .B(n24632), .Z(n30784) );
  XOR U30802 ( .A(n30786), .B(\modmult_1/zin[0][1017] ), .Z(n24632) );
  IV U30803 ( .A(n30783), .Z(n30786) );
  XNOR U30804 ( .A(n30783), .B(n24631), .Z(n30785) );
  XOR U30805 ( .A(n30787), .B(n30788), .Z(n24631) );
  AND U30806 ( .A(\modmult_1/xin[1023] ), .B(n30789), .Z(n30788) );
  IV U30807 ( .A(n30787), .Z(n30789) );
  XOR U30808 ( .A(n30790), .B(g_input[1018]), .Z(n30787) );
  NAND U30809 ( .A(n30791), .B(mul_pow), .Z(n30790) );
  XOR U30810 ( .A(g_input[1018]), .B(creg[1018]), .Z(n30791) );
  XOR U30811 ( .A(n30792), .B(n30793), .Z(n30783) );
  ANDN U30812 ( .A(n30794), .B(n24638), .Z(n30793) );
  XOR U30813 ( .A(n30795), .B(\modmult_1/zin[0][1016] ), .Z(n24638) );
  IV U30814 ( .A(n30792), .Z(n30795) );
  XNOR U30815 ( .A(n30792), .B(n24637), .Z(n30794) );
  XOR U30816 ( .A(n30796), .B(n30797), .Z(n24637) );
  AND U30817 ( .A(\modmult_1/xin[1023] ), .B(n30798), .Z(n30797) );
  IV U30818 ( .A(n30796), .Z(n30798) );
  XOR U30819 ( .A(n30799), .B(g_input[1017]), .Z(n30796) );
  NAND U30820 ( .A(n30800), .B(mul_pow), .Z(n30799) );
  XOR U30821 ( .A(g_input[1017]), .B(creg[1017]), .Z(n30800) );
  XOR U30822 ( .A(n30801), .B(n30802), .Z(n30792) );
  ANDN U30823 ( .A(n30803), .B(n24644), .Z(n30802) );
  XOR U30824 ( .A(n30804), .B(\modmult_1/zin[0][1015] ), .Z(n24644) );
  IV U30825 ( .A(n30801), .Z(n30804) );
  XNOR U30826 ( .A(n30801), .B(n24643), .Z(n30803) );
  XOR U30827 ( .A(n30805), .B(n30806), .Z(n24643) );
  AND U30828 ( .A(\modmult_1/xin[1023] ), .B(n30807), .Z(n30806) );
  IV U30829 ( .A(n30805), .Z(n30807) );
  XOR U30830 ( .A(n30808), .B(g_input[1016]), .Z(n30805) );
  NAND U30831 ( .A(n30809), .B(mul_pow), .Z(n30808) );
  XOR U30832 ( .A(g_input[1016]), .B(creg[1016]), .Z(n30809) );
  XOR U30833 ( .A(n30810), .B(n30811), .Z(n30801) );
  ANDN U30834 ( .A(n30812), .B(n24650), .Z(n30811) );
  XOR U30835 ( .A(n30813), .B(\modmult_1/zin[0][1014] ), .Z(n24650) );
  IV U30836 ( .A(n30810), .Z(n30813) );
  XNOR U30837 ( .A(n30810), .B(n24649), .Z(n30812) );
  XOR U30838 ( .A(n30814), .B(n30815), .Z(n24649) );
  AND U30839 ( .A(\modmult_1/xin[1023] ), .B(n30816), .Z(n30815) );
  IV U30840 ( .A(n30814), .Z(n30816) );
  XOR U30841 ( .A(n30817), .B(g_input[1015]), .Z(n30814) );
  NAND U30842 ( .A(n30818), .B(mul_pow), .Z(n30817) );
  XOR U30843 ( .A(g_input[1015]), .B(creg[1015]), .Z(n30818) );
  XOR U30844 ( .A(n30819), .B(n30820), .Z(n30810) );
  ANDN U30845 ( .A(n30821), .B(n24656), .Z(n30820) );
  XOR U30846 ( .A(n30822), .B(\modmult_1/zin[0][1013] ), .Z(n24656) );
  IV U30847 ( .A(n30819), .Z(n30822) );
  XNOR U30848 ( .A(n30819), .B(n24655), .Z(n30821) );
  XOR U30849 ( .A(n30823), .B(n30824), .Z(n24655) );
  AND U30850 ( .A(\modmult_1/xin[1023] ), .B(n30825), .Z(n30824) );
  IV U30851 ( .A(n30823), .Z(n30825) );
  XOR U30852 ( .A(n30826), .B(g_input[1014]), .Z(n30823) );
  NAND U30853 ( .A(n30827), .B(mul_pow), .Z(n30826) );
  XOR U30854 ( .A(g_input[1014]), .B(creg[1014]), .Z(n30827) );
  XOR U30855 ( .A(n30828), .B(n30829), .Z(n30819) );
  ANDN U30856 ( .A(n30830), .B(n24662), .Z(n30829) );
  XOR U30857 ( .A(n30831), .B(\modmult_1/zin[0][1012] ), .Z(n24662) );
  IV U30858 ( .A(n30828), .Z(n30831) );
  XNOR U30859 ( .A(n30828), .B(n24661), .Z(n30830) );
  XOR U30860 ( .A(n30832), .B(n30833), .Z(n24661) );
  AND U30861 ( .A(\modmult_1/xin[1023] ), .B(n30834), .Z(n30833) );
  IV U30862 ( .A(n30832), .Z(n30834) );
  XOR U30863 ( .A(n30835), .B(g_input[1013]), .Z(n30832) );
  NAND U30864 ( .A(n30836), .B(mul_pow), .Z(n30835) );
  XOR U30865 ( .A(g_input[1013]), .B(creg[1013]), .Z(n30836) );
  XOR U30866 ( .A(n30837), .B(n30838), .Z(n30828) );
  ANDN U30867 ( .A(n30839), .B(n24668), .Z(n30838) );
  XOR U30868 ( .A(n30840), .B(\modmult_1/zin[0][1011] ), .Z(n24668) );
  IV U30869 ( .A(n30837), .Z(n30840) );
  XNOR U30870 ( .A(n30837), .B(n24667), .Z(n30839) );
  XOR U30871 ( .A(n30841), .B(n30842), .Z(n24667) );
  AND U30872 ( .A(\modmult_1/xin[1023] ), .B(n30843), .Z(n30842) );
  IV U30873 ( .A(n30841), .Z(n30843) );
  XOR U30874 ( .A(n30844), .B(g_input[1012]), .Z(n30841) );
  NAND U30875 ( .A(n30845), .B(mul_pow), .Z(n30844) );
  XOR U30876 ( .A(g_input[1012]), .B(creg[1012]), .Z(n30845) );
  XOR U30877 ( .A(n30846), .B(n30847), .Z(n30837) );
  ANDN U30878 ( .A(n30848), .B(n24674), .Z(n30847) );
  XOR U30879 ( .A(n30849), .B(\modmult_1/zin[0][1010] ), .Z(n24674) );
  IV U30880 ( .A(n30846), .Z(n30849) );
  XNOR U30881 ( .A(n30846), .B(n24673), .Z(n30848) );
  XOR U30882 ( .A(n30850), .B(n30851), .Z(n24673) );
  AND U30883 ( .A(\modmult_1/xin[1023] ), .B(n30852), .Z(n30851) );
  IV U30884 ( .A(n30850), .Z(n30852) );
  XOR U30885 ( .A(n30853), .B(g_input[1011]), .Z(n30850) );
  NAND U30886 ( .A(n30854), .B(mul_pow), .Z(n30853) );
  XOR U30887 ( .A(g_input[1011]), .B(creg[1011]), .Z(n30854) );
  XOR U30888 ( .A(n30855), .B(n30856), .Z(n30846) );
  ANDN U30889 ( .A(n30857), .B(n24680), .Z(n30856) );
  XOR U30890 ( .A(n30858), .B(\modmult_1/zin[0][1009] ), .Z(n24680) );
  IV U30891 ( .A(n30855), .Z(n30858) );
  XNOR U30892 ( .A(n30855), .B(n24679), .Z(n30857) );
  XOR U30893 ( .A(n30859), .B(n30860), .Z(n24679) );
  AND U30894 ( .A(\modmult_1/xin[1023] ), .B(n30861), .Z(n30860) );
  IV U30895 ( .A(n30859), .Z(n30861) );
  XOR U30896 ( .A(n30862), .B(g_input[1010]), .Z(n30859) );
  NAND U30897 ( .A(n30863), .B(mul_pow), .Z(n30862) );
  XOR U30898 ( .A(g_input[1010]), .B(creg[1010]), .Z(n30863) );
  XOR U30899 ( .A(n30864), .B(n30865), .Z(n30855) );
  ANDN U30900 ( .A(n30866), .B(n24686), .Z(n30865) );
  XOR U30901 ( .A(n30867), .B(\modmult_1/zin[0][1008] ), .Z(n24686) );
  IV U30902 ( .A(n30864), .Z(n30867) );
  XNOR U30903 ( .A(n30864), .B(n24685), .Z(n30866) );
  XOR U30904 ( .A(n30868), .B(n30869), .Z(n24685) );
  AND U30905 ( .A(\modmult_1/xin[1023] ), .B(n30870), .Z(n30869) );
  IV U30906 ( .A(n30868), .Z(n30870) );
  XOR U30907 ( .A(n30871), .B(g_input[1009]), .Z(n30868) );
  NAND U30908 ( .A(n30872), .B(mul_pow), .Z(n30871) );
  XOR U30909 ( .A(g_input[1009]), .B(creg[1009]), .Z(n30872) );
  XOR U30910 ( .A(n30873), .B(n30874), .Z(n30864) );
  ANDN U30911 ( .A(n30875), .B(n24692), .Z(n30874) );
  XOR U30912 ( .A(n30876), .B(\modmult_1/zin[0][1007] ), .Z(n24692) );
  IV U30913 ( .A(n30873), .Z(n30876) );
  XNOR U30914 ( .A(n30873), .B(n24691), .Z(n30875) );
  XOR U30915 ( .A(n30877), .B(n30878), .Z(n24691) );
  AND U30916 ( .A(\modmult_1/xin[1023] ), .B(n30879), .Z(n30878) );
  IV U30917 ( .A(n30877), .Z(n30879) );
  XOR U30918 ( .A(n30880), .B(g_input[1008]), .Z(n30877) );
  NAND U30919 ( .A(n30881), .B(mul_pow), .Z(n30880) );
  XOR U30920 ( .A(g_input[1008]), .B(creg[1008]), .Z(n30881) );
  XOR U30921 ( .A(n30882), .B(n30883), .Z(n30873) );
  ANDN U30922 ( .A(n30884), .B(n24698), .Z(n30883) );
  XOR U30923 ( .A(n30885), .B(\modmult_1/zin[0][1006] ), .Z(n24698) );
  IV U30924 ( .A(n30882), .Z(n30885) );
  XNOR U30925 ( .A(n30882), .B(n24697), .Z(n30884) );
  XOR U30926 ( .A(n30886), .B(n30887), .Z(n24697) );
  AND U30927 ( .A(\modmult_1/xin[1023] ), .B(n30888), .Z(n30887) );
  IV U30928 ( .A(n30886), .Z(n30888) );
  XOR U30929 ( .A(n30889), .B(g_input[1007]), .Z(n30886) );
  NAND U30930 ( .A(n30890), .B(mul_pow), .Z(n30889) );
  XOR U30931 ( .A(g_input[1007]), .B(creg[1007]), .Z(n30890) );
  XOR U30932 ( .A(n30891), .B(n30892), .Z(n30882) );
  ANDN U30933 ( .A(n30893), .B(n24704), .Z(n30892) );
  XOR U30934 ( .A(n30894), .B(\modmult_1/zin[0][1005] ), .Z(n24704) );
  IV U30935 ( .A(n30891), .Z(n30894) );
  XNOR U30936 ( .A(n30891), .B(n24703), .Z(n30893) );
  XOR U30937 ( .A(n30895), .B(n30896), .Z(n24703) );
  AND U30938 ( .A(\modmult_1/xin[1023] ), .B(n30897), .Z(n30896) );
  IV U30939 ( .A(n30895), .Z(n30897) );
  XOR U30940 ( .A(n30898), .B(g_input[1006]), .Z(n30895) );
  NAND U30941 ( .A(n30899), .B(mul_pow), .Z(n30898) );
  XOR U30942 ( .A(g_input[1006]), .B(creg[1006]), .Z(n30899) );
  XOR U30943 ( .A(n30900), .B(n30901), .Z(n30891) );
  ANDN U30944 ( .A(n30902), .B(n24710), .Z(n30901) );
  XOR U30945 ( .A(n30903), .B(\modmult_1/zin[0][1004] ), .Z(n24710) );
  IV U30946 ( .A(n30900), .Z(n30903) );
  XNOR U30947 ( .A(n30900), .B(n24709), .Z(n30902) );
  XOR U30948 ( .A(n30904), .B(n30905), .Z(n24709) );
  AND U30949 ( .A(\modmult_1/xin[1023] ), .B(n30906), .Z(n30905) );
  IV U30950 ( .A(n30904), .Z(n30906) );
  XOR U30951 ( .A(n30907), .B(g_input[1005]), .Z(n30904) );
  NAND U30952 ( .A(n30908), .B(mul_pow), .Z(n30907) );
  XOR U30953 ( .A(g_input[1005]), .B(creg[1005]), .Z(n30908) );
  XOR U30954 ( .A(n30909), .B(n30910), .Z(n30900) );
  ANDN U30955 ( .A(n30911), .B(n24716), .Z(n30910) );
  XOR U30956 ( .A(n30912), .B(\modmult_1/zin[0][1003] ), .Z(n24716) );
  IV U30957 ( .A(n30909), .Z(n30912) );
  XNOR U30958 ( .A(n30909), .B(n24715), .Z(n30911) );
  XOR U30959 ( .A(n30913), .B(n30914), .Z(n24715) );
  AND U30960 ( .A(\modmult_1/xin[1023] ), .B(n30915), .Z(n30914) );
  IV U30961 ( .A(n30913), .Z(n30915) );
  XOR U30962 ( .A(n30916), .B(g_input[1004]), .Z(n30913) );
  NAND U30963 ( .A(n30917), .B(mul_pow), .Z(n30916) );
  XOR U30964 ( .A(g_input[1004]), .B(creg[1004]), .Z(n30917) );
  XOR U30965 ( .A(n30918), .B(n30919), .Z(n30909) );
  ANDN U30966 ( .A(n30920), .B(n24722), .Z(n30919) );
  XOR U30967 ( .A(n30921), .B(\modmult_1/zin[0][1002] ), .Z(n24722) );
  IV U30968 ( .A(n30918), .Z(n30921) );
  XNOR U30969 ( .A(n30918), .B(n24721), .Z(n30920) );
  XOR U30970 ( .A(n30922), .B(n30923), .Z(n24721) );
  AND U30971 ( .A(\modmult_1/xin[1023] ), .B(n30924), .Z(n30923) );
  IV U30972 ( .A(n30922), .Z(n30924) );
  XOR U30973 ( .A(n30925), .B(g_input[1003]), .Z(n30922) );
  NAND U30974 ( .A(n30926), .B(mul_pow), .Z(n30925) );
  XOR U30975 ( .A(g_input[1003]), .B(creg[1003]), .Z(n30926) );
  XOR U30976 ( .A(n30927), .B(n30928), .Z(n30918) );
  ANDN U30977 ( .A(n30929), .B(n24728), .Z(n30928) );
  XOR U30978 ( .A(n30930), .B(\modmult_1/zin[0][1001] ), .Z(n24728) );
  IV U30979 ( .A(n30927), .Z(n30930) );
  XNOR U30980 ( .A(n30927), .B(n24727), .Z(n30929) );
  XOR U30981 ( .A(n30931), .B(n30932), .Z(n24727) );
  AND U30982 ( .A(\modmult_1/xin[1023] ), .B(n30933), .Z(n30932) );
  IV U30983 ( .A(n30931), .Z(n30933) );
  XOR U30984 ( .A(n30934), .B(g_input[1002]), .Z(n30931) );
  NAND U30985 ( .A(n30935), .B(mul_pow), .Z(n30934) );
  XOR U30986 ( .A(g_input[1002]), .B(creg[1002]), .Z(n30935) );
  XOR U30987 ( .A(n30936), .B(n30937), .Z(n30927) );
  ANDN U30988 ( .A(n30938), .B(n24734), .Z(n30937) );
  XOR U30989 ( .A(n30939), .B(\modmult_1/zin[0][1000] ), .Z(n24734) );
  IV U30990 ( .A(n30936), .Z(n30939) );
  XNOR U30991 ( .A(n30936), .B(n24733), .Z(n30938) );
  XOR U30992 ( .A(n30940), .B(n30941), .Z(n24733) );
  AND U30993 ( .A(\modmult_1/xin[1023] ), .B(n30942), .Z(n30941) );
  IV U30994 ( .A(n30940), .Z(n30942) );
  XOR U30995 ( .A(n30943), .B(g_input[1001]), .Z(n30940) );
  NAND U30996 ( .A(n30944), .B(mul_pow), .Z(n30943) );
  XOR U30997 ( .A(g_input[1001]), .B(creg[1001]), .Z(n30944) );
  XOR U30998 ( .A(n30945), .B(n30946), .Z(n30936) );
  ANDN U30999 ( .A(n30947), .B(n24740), .Z(n30946) );
  XOR U31000 ( .A(n30948), .B(\modmult_1/zin[0][999] ), .Z(n24740) );
  IV U31001 ( .A(n30945), .Z(n30948) );
  XNOR U31002 ( .A(n30945), .B(n24739), .Z(n30947) );
  XOR U31003 ( .A(n30949), .B(n30950), .Z(n24739) );
  AND U31004 ( .A(\modmult_1/xin[1023] ), .B(n30951), .Z(n30950) );
  IV U31005 ( .A(n30949), .Z(n30951) );
  XOR U31006 ( .A(n30952), .B(g_input[1000]), .Z(n30949) );
  NAND U31007 ( .A(n30953), .B(mul_pow), .Z(n30952) );
  XOR U31008 ( .A(g_input[1000]), .B(creg[1000]), .Z(n30953) );
  XOR U31009 ( .A(n30954), .B(n30955), .Z(n30945) );
  ANDN U31010 ( .A(n30956), .B(n24746), .Z(n30955) );
  XOR U31011 ( .A(n30957), .B(\modmult_1/zin[0][998] ), .Z(n24746) );
  IV U31012 ( .A(n30954), .Z(n30957) );
  XNOR U31013 ( .A(n30954), .B(n24745), .Z(n30956) );
  XOR U31014 ( .A(n30958), .B(n30959), .Z(n24745) );
  AND U31015 ( .A(\modmult_1/xin[1023] ), .B(n30960), .Z(n30959) );
  IV U31016 ( .A(n30958), .Z(n30960) );
  XOR U31017 ( .A(n30961), .B(g_input[999]), .Z(n30958) );
  NAND U31018 ( .A(n30962), .B(mul_pow), .Z(n30961) );
  XOR U31019 ( .A(g_input[999]), .B(creg[999]), .Z(n30962) );
  XOR U31020 ( .A(n30963), .B(n30964), .Z(n30954) );
  ANDN U31021 ( .A(n30965), .B(n24752), .Z(n30964) );
  XOR U31022 ( .A(n30966), .B(\modmult_1/zin[0][997] ), .Z(n24752) );
  IV U31023 ( .A(n30963), .Z(n30966) );
  XNOR U31024 ( .A(n30963), .B(n24751), .Z(n30965) );
  XOR U31025 ( .A(n30967), .B(n30968), .Z(n24751) );
  AND U31026 ( .A(\modmult_1/xin[1023] ), .B(n30969), .Z(n30968) );
  IV U31027 ( .A(n30967), .Z(n30969) );
  XOR U31028 ( .A(n30970), .B(g_input[998]), .Z(n30967) );
  NAND U31029 ( .A(n30971), .B(mul_pow), .Z(n30970) );
  XOR U31030 ( .A(g_input[998]), .B(creg[998]), .Z(n30971) );
  XOR U31031 ( .A(n30972), .B(n30973), .Z(n30963) );
  ANDN U31032 ( .A(n30974), .B(n24758), .Z(n30973) );
  XOR U31033 ( .A(n30975), .B(\modmult_1/zin[0][996] ), .Z(n24758) );
  IV U31034 ( .A(n30972), .Z(n30975) );
  XNOR U31035 ( .A(n30972), .B(n24757), .Z(n30974) );
  XOR U31036 ( .A(n30976), .B(n30977), .Z(n24757) );
  AND U31037 ( .A(\modmult_1/xin[1023] ), .B(n30978), .Z(n30977) );
  IV U31038 ( .A(n30976), .Z(n30978) );
  XOR U31039 ( .A(n30979), .B(g_input[997]), .Z(n30976) );
  NAND U31040 ( .A(n30980), .B(mul_pow), .Z(n30979) );
  XOR U31041 ( .A(g_input[997]), .B(creg[997]), .Z(n30980) );
  XOR U31042 ( .A(n30981), .B(n30982), .Z(n30972) );
  ANDN U31043 ( .A(n30983), .B(n24764), .Z(n30982) );
  XOR U31044 ( .A(n30984), .B(\modmult_1/zin[0][995] ), .Z(n24764) );
  IV U31045 ( .A(n30981), .Z(n30984) );
  XNOR U31046 ( .A(n30981), .B(n24763), .Z(n30983) );
  XOR U31047 ( .A(n30985), .B(n30986), .Z(n24763) );
  AND U31048 ( .A(\modmult_1/xin[1023] ), .B(n30987), .Z(n30986) );
  IV U31049 ( .A(n30985), .Z(n30987) );
  XOR U31050 ( .A(n30988), .B(g_input[996]), .Z(n30985) );
  NAND U31051 ( .A(n30989), .B(mul_pow), .Z(n30988) );
  XOR U31052 ( .A(g_input[996]), .B(creg[996]), .Z(n30989) );
  XOR U31053 ( .A(n30990), .B(n30991), .Z(n30981) );
  ANDN U31054 ( .A(n30992), .B(n24770), .Z(n30991) );
  XOR U31055 ( .A(n30993), .B(\modmult_1/zin[0][994] ), .Z(n24770) );
  IV U31056 ( .A(n30990), .Z(n30993) );
  XNOR U31057 ( .A(n30990), .B(n24769), .Z(n30992) );
  XOR U31058 ( .A(n30994), .B(n30995), .Z(n24769) );
  AND U31059 ( .A(\modmult_1/xin[1023] ), .B(n30996), .Z(n30995) );
  IV U31060 ( .A(n30994), .Z(n30996) );
  XOR U31061 ( .A(n30997), .B(g_input[995]), .Z(n30994) );
  NAND U31062 ( .A(n30998), .B(mul_pow), .Z(n30997) );
  XOR U31063 ( .A(g_input[995]), .B(creg[995]), .Z(n30998) );
  XOR U31064 ( .A(n30999), .B(n31000), .Z(n30990) );
  ANDN U31065 ( .A(n31001), .B(n24776), .Z(n31000) );
  XOR U31066 ( .A(n31002), .B(\modmult_1/zin[0][993] ), .Z(n24776) );
  IV U31067 ( .A(n30999), .Z(n31002) );
  XNOR U31068 ( .A(n30999), .B(n24775), .Z(n31001) );
  XOR U31069 ( .A(n31003), .B(n31004), .Z(n24775) );
  AND U31070 ( .A(\modmult_1/xin[1023] ), .B(n31005), .Z(n31004) );
  IV U31071 ( .A(n31003), .Z(n31005) );
  XOR U31072 ( .A(n31006), .B(g_input[994]), .Z(n31003) );
  NAND U31073 ( .A(n31007), .B(mul_pow), .Z(n31006) );
  XOR U31074 ( .A(g_input[994]), .B(creg[994]), .Z(n31007) );
  XOR U31075 ( .A(n31008), .B(n31009), .Z(n30999) );
  ANDN U31076 ( .A(n31010), .B(n24782), .Z(n31009) );
  XOR U31077 ( .A(n31011), .B(\modmult_1/zin[0][992] ), .Z(n24782) );
  IV U31078 ( .A(n31008), .Z(n31011) );
  XNOR U31079 ( .A(n31008), .B(n24781), .Z(n31010) );
  XOR U31080 ( .A(n31012), .B(n31013), .Z(n24781) );
  AND U31081 ( .A(\modmult_1/xin[1023] ), .B(n31014), .Z(n31013) );
  IV U31082 ( .A(n31012), .Z(n31014) );
  XOR U31083 ( .A(n31015), .B(g_input[993]), .Z(n31012) );
  NAND U31084 ( .A(n31016), .B(mul_pow), .Z(n31015) );
  XOR U31085 ( .A(g_input[993]), .B(creg[993]), .Z(n31016) );
  XOR U31086 ( .A(n31017), .B(n31018), .Z(n31008) );
  ANDN U31087 ( .A(n31019), .B(n24788), .Z(n31018) );
  XOR U31088 ( .A(n31020), .B(\modmult_1/zin[0][991] ), .Z(n24788) );
  IV U31089 ( .A(n31017), .Z(n31020) );
  XNOR U31090 ( .A(n31017), .B(n24787), .Z(n31019) );
  XOR U31091 ( .A(n31021), .B(n31022), .Z(n24787) );
  AND U31092 ( .A(\modmult_1/xin[1023] ), .B(n31023), .Z(n31022) );
  IV U31093 ( .A(n31021), .Z(n31023) );
  XOR U31094 ( .A(n31024), .B(g_input[992]), .Z(n31021) );
  NAND U31095 ( .A(n31025), .B(mul_pow), .Z(n31024) );
  XOR U31096 ( .A(g_input[992]), .B(creg[992]), .Z(n31025) );
  XOR U31097 ( .A(n31026), .B(n31027), .Z(n31017) );
  ANDN U31098 ( .A(n31028), .B(n24794), .Z(n31027) );
  XOR U31099 ( .A(n31029), .B(\modmult_1/zin[0][990] ), .Z(n24794) );
  IV U31100 ( .A(n31026), .Z(n31029) );
  XNOR U31101 ( .A(n31026), .B(n24793), .Z(n31028) );
  XOR U31102 ( .A(n31030), .B(n31031), .Z(n24793) );
  AND U31103 ( .A(\modmult_1/xin[1023] ), .B(n31032), .Z(n31031) );
  IV U31104 ( .A(n31030), .Z(n31032) );
  XOR U31105 ( .A(n31033), .B(g_input[991]), .Z(n31030) );
  NAND U31106 ( .A(n31034), .B(mul_pow), .Z(n31033) );
  XOR U31107 ( .A(g_input[991]), .B(creg[991]), .Z(n31034) );
  XOR U31108 ( .A(n31035), .B(n31036), .Z(n31026) );
  ANDN U31109 ( .A(n31037), .B(n24800), .Z(n31036) );
  XOR U31110 ( .A(n31038), .B(\modmult_1/zin[0][989] ), .Z(n24800) );
  IV U31111 ( .A(n31035), .Z(n31038) );
  XNOR U31112 ( .A(n31035), .B(n24799), .Z(n31037) );
  XOR U31113 ( .A(n31039), .B(n31040), .Z(n24799) );
  AND U31114 ( .A(\modmult_1/xin[1023] ), .B(n31041), .Z(n31040) );
  IV U31115 ( .A(n31039), .Z(n31041) );
  XOR U31116 ( .A(n31042), .B(g_input[990]), .Z(n31039) );
  NAND U31117 ( .A(n31043), .B(mul_pow), .Z(n31042) );
  XOR U31118 ( .A(g_input[990]), .B(creg[990]), .Z(n31043) );
  XOR U31119 ( .A(n31044), .B(n31045), .Z(n31035) );
  ANDN U31120 ( .A(n31046), .B(n24806), .Z(n31045) );
  XOR U31121 ( .A(n31047), .B(\modmult_1/zin[0][988] ), .Z(n24806) );
  IV U31122 ( .A(n31044), .Z(n31047) );
  XNOR U31123 ( .A(n31044), .B(n24805), .Z(n31046) );
  XOR U31124 ( .A(n31048), .B(n31049), .Z(n24805) );
  AND U31125 ( .A(\modmult_1/xin[1023] ), .B(n31050), .Z(n31049) );
  IV U31126 ( .A(n31048), .Z(n31050) );
  XOR U31127 ( .A(n31051), .B(g_input[989]), .Z(n31048) );
  NAND U31128 ( .A(n31052), .B(mul_pow), .Z(n31051) );
  XOR U31129 ( .A(g_input[989]), .B(creg[989]), .Z(n31052) );
  XOR U31130 ( .A(n31053), .B(n31054), .Z(n31044) );
  ANDN U31131 ( .A(n31055), .B(n24812), .Z(n31054) );
  XOR U31132 ( .A(n31056), .B(\modmult_1/zin[0][987] ), .Z(n24812) );
  IV U31133 ( .A(n31053), .Z(n31056) );
  XNOR U31134 ( .A(n31053), .B(n24811), .Z(n31055) );
  XOR U31135 ( .A(n31057), .B(n31058), .Z(n24811) );
  AND U31136 ( .A(\modmult_1/xin[1023] ), .B(n31059), .Z(n31058) );
  IV U31137 ( .A(n31057), .Z(n31059) );
  XOR U31138 ( .A(n31060), .B(g_input[988]), .Z(n31057) );
  NAND U31139 ( .A(n31061), .B(mul_pow), .Z(n31060) );
  XOR U31140 ( .A(g_input[988]), .B(creg[988]), .Z(n31061) );
  XOR U31141 ( .A(n31062), .B(n31063), .Z(n31053) );
  ANDN U31142 ( .A(n31064), .B(n24818), .Z(n31063) );
  XOR U31143 ( .A(n31065), .B(\modmult_1/zin[0][986] ), .Z(n24818) );
  IV U31144 ( .A(n31062), .Z(n31065) );
  XNOR U31145 ( .A(n31062), .B(n24817), .Z(n31064) );
  XOR U31146 ( .A(n31066), .B(n31067), .Z(n24817) );
  AND U31147 ( .A(\modmult_1/xin[1023] ), .B(n31068), .Z(n31067) );
  IV U31148 ( .A(n31066), .Z(n31068) );
  XOR U31149 ( .A(n31069), .B(g_input[987]), .Z(n31066) );
  NAND U31150 ( .A(n31070), .B(mul_pow), .Z(n31069) );
  XOR U31151 ( .A(g_input[987]), .B(creg[987]), .Z(n31070) );
  XOR U31152 ( .A(n31071), .B(n31072), .Z(n31062) );
  ANDN U31153 ( .A(n31073), .B(n24824), .Z(n31072) );
  XOR U31154 ( .A(n31074), .B(\modmult_1/zin[0][985] ), .Z(n24824) );
  IV U31155 ( .A(n31071), .Z(n31074) );
  XNOR U31156 ( .A(n31071), .B(n24823), .Z(n31073) );
  XOR U31157 ( .A(n31075), .B(n31076), .Z(n24823) );
  AND U31158 ( .A(\modmult_1/xin[1023] ), .B(n31077), .Z(n31076) );
  IV U31159 ( .A(n31075), .Z(n31077) );
  XOR U31160 ( .A(n31078), .B(g_input[986]), .Z(n31075) );
  NAND U31161 ( .A(n31079), .B(mul_pow), .Z(n31078) );
  XOR U31162 ( .A(g_input[986]), .B(creg[986]), .Z(n31079) );
  XOR U31163 ( .A(n31080), .B(n31081), .Z(n31071) );
  ANDN U31164 ( .A(n31082), .B(n24830), .Z(n31081) );
  XOR U31165 ( .A(n31083), .B(\modmult_1/zin[0][984] ), .Z(n24830) );
  IV U31166 ( .A(n31080), .Z(n31083) );
  XNOR U31167 ( .A(n31080), .B(n24829), .Z(n31082) );
  XOR U31168 ( .A(n31084), .B(n31085), .Z(n24829) );
  AND U31169 ( .A(\modmult_1/xin[1023] ), .B(n31086), .Z(n31085) );
  IV U31170 ( .A(n31084), .Z(n31086) );
  XOR U31171 ( .A(n31087), .B(g_input[985]), .Z(n31084) );
  NAND U31172 ( .A(n31088), .B(mul_pow), .Z(n31087) );
  XOR U31173 ( .A(g_input[985]), .B(creg[985]), .Z(n31088) );
  XOR U31174 ( .A(n31089), .B(n31090), .Z(n31080) );
  ANDN U31175 ( .A(n31091), .B(n24836), .Z(n31090) );
  XOR U31176 ( .A(n31092), .B(\modmult_1/zin[0][983] ), .Z(n24836) );
  IV U31177 ( .A(n31089), .Z(n31092) );
  XNOR U31178 ( .A(n31089), .B(n24835), .Z(n31091) );
  XOR U31179 ( .A(n31093), .B(n31094), .Z(n24835) );
  AND U31180 ( .A(\modmult_1/xin[1023] ), .B(n31095), .Z(n31094) );
  IV U31181 ( .A(n31093), .Z(n31095) );
  XOR U31182 ( .A(n31096), .B(g_input[984]), .Z(n31093) );
  NAND U31183 ( .A(n31097), .B(mul_pow), .Z(n31096) );
  XOR U31184 ( .A(g_input[984]), .B(creg[984]), .Z(n31097) );
  XOR U31185 ( .A(n31098), .B(n31099), .Z(n31089) );
  ANDN U31186 ( .A(n31100), .B(n24842), .Z(n31099) );
  XOR U31187 ( .A(n31101), .B(\modmult_1/zin[0][982] ), .Z(n24842) );
  IV U31188 ( .A(n31098), .Z(n31101) );
  XNOR U31189 ( .A(n31098), .B(n24841), .Z(n31100) );
  XOR U31190 ( .A(n31102), .B(n31103), .Z(n24841) );
  AND U31191 ( .A(\modmult_1/xin[1023] ), .B(n31104), .Z(n31103) );
  IV U31192 ( .A(n31102), .Z(n31104) );
  XOR U31193 ( .A(n31105), .B(g_input[983]), .Z(n31102) );
  NAND U31194 ( .A(n31106), .B(mul_pow), .Z(n31105) );
  XOR U31195 ( .A(g_input[983]), .B(creg[983]), .Z(n31106) );
  XOR U31196 ( .A(n31107), .B(n31108), .Z(n31098) );
  ANDN U31197 ( .A(n31109), .B(n24848), .Z(n31108) );
  XOR U31198 ( .A(n31110), .B(\modmult_1/zin[0][981] ), .Z(n24848) );
  IV U31199 ( .A(n31107), .Z(n31110) );
  XNOR U31200 ( .A(n31107), .B(n24847), .Z(n31109) );
  XOR U31201 ( .A(n31111), .B(n31112), .Z(n24847) );
  AND U31202 ( .A(\modmult_1/xin[1023] ), .B(n31113), .Z(n31112) );
  IV U31203 ( .A(n31111), .Z(n31113) );
  XOR U31204 ( .A(n31114), .B(g_input[982]), .Z(n31111) );
  NAND U31205 ( .A(n31115), .B(mul_pow), .Z(n31114) );
  XOR U31206 ( .A(g_input[982]), .B(creg[982]), .Z(n31115) );
  XOR U31207 ( .A(n31116), .B(n31117), .Z(n31107) );
  ANDN U31208 ( .A(n31118), .B(n24854), .Z(n31117) );
  XOR U31209 ( .A(n31119), .B(\modmult_1/zin[0][980] ), .Z(n24854) );
  IV U31210 ( .A(n31116), .Z(n31119) );
  XNOR U31211 ( .A(n31116), .B(n24853), .Z(n31118) );
  XOR U31212 ( .A(n31120), .B(n31121), .Z(n24853) );
  AND U31213 ( .A(\modmult_1/xin[1023] ), .B(n31122), .Z(n31121) );
  IV U31214 ( .A(n31120), .Z(n31122) );
  XOR U31215 ( .A(n31123), .B(g_input[981]), .Z(n31120) );
  NAND U31216 ( .A(n31124), .B(mul_pow), .Z(n31123) );
  XOR U31217 ( .A(g_input[981]), .B(creg[981]), .Z(n31124) );
  XOR U31218 ( .A(n31125), .B(n31126), .Z(n31116) );
  ANDN U31219 ( .A(n31127), .B(n24860), .Z(n31126) );
  XOR U31220 ( .A(n31128), .B(\modmult_1/zin[0][979] ), .Z(n24860) );
  IV U31221 ( .A(n31125), .Z(n31128) );
  XNOR U31222 ( .A(n31125), .B(n24859), .Z(n31127) );
  XOR U31223 ( .A(n31129), .B(n31130), .Z(n24859) );
  AND U31224 ( .A(\modmult_1/xin[1023] ), .B(n31131), .Z(n31130) );
  IV U31225 ( .A(n31129), .Z(n31131) );
  XOR U31226 ( .A(n31132), .B(g_input[980]), .Z(n31129) );
  NAND U31227 ( .A(n31133), .B(mul_pow), .Z(n31132) );
  XOR U31228 ( .A(g_input[980]), .B(creg[980]), .Z(n31133) );
  XOR U31229 ( .A(n31134), .B(n31135), .Z(n31125) );
  ANDN U31230 ( .A(n31136), .B(n24866), .Z(n31135) );
  XOR U31231 ( .A(n31137), .B(\modmult_1/zin[0][978] ), .Z(n24866) );
  IV U31232 ( .A(n31134), .Z(n31137) );
  XNOR U31233 ( .A(n31134), .B(n24865), .Z(n31136) );
  XOR U31234 ( .A(n31138), .B(n31139), .Z(n24865) );
  AND U31235 ( .A(\modmult_1/xin[1023] ), .B(n31140), .Z(n31139) );
  IV U31236 ( .A(n31138), .Z(n31140) );
  XOR U31237 ( .A(n31141), .B(g_input[979]), .Z(n31138) );
  NAND U31238 ( .A(n31142), .B(mul_pow), .Z(n31141) );
  XOR U31239 ( .A(g_input[979]), .B(creg[979]), .Z(n31142) );
  XOR U31240 ( .A(n31143), .B(n31144), .Z(n31134) );
  ANDN U31241 ( .A(n31145), .B(n24872), .Z(n31144) );
  XOR U31242 ( .A(n31146), .B(\modmult_1/zin[0][977] ), .Z(n24872) );
  IV U31243 ( .A(n31143), .Z(n31146) );
  XNOR U31244 ( .A(n31143), .B(n24871), .Z(n31145) );
  XOR U31245 ( .A(n31147), .B(n31148), .Z(n24871) );
  AND U31246 ( .A(\modmult_1/xin[1023] ), .B(n31149), .Z(n31148) );
  IV U31247 ( .A(n31147), .Z(n31149) );
  XOR U31248 ( .A(n31150), .B(g_input[978]), .Z(n31147) );
  NAND U31249 ( .A(n31151), .B(mul_pow), .Z(n31150) );
  XOR U31250 ( .A(g_input[978]), .B(creg[978]), .Z(n31151) );
  XOR U31251 ( .A(n31152), .B(n31153), .Z(n31143) );
  ANDN U31252 ( .A(n31154), .B(n24878), .Z(n31153) );
  XOR U31253 ( .A(n31155), .B(\modmult_1/zin[0][976] ), .Z(n24878) );
  IV U31254 ( .A(n31152), .Z(n31155) );
  XNOR U31255 ( .A(n31152), .B(n24877), .Z(n31154) );
  XOR U31256 ( .A(n31156), .B(n31157), .Z(n24877) );
  AND U31257 ( .A(\modmult_1/xin[1023] ), .B(n31158), .Z(n31157) );
  IV U31258 ( .A(n31156), .Z(n31158) );
  XOR U31259 ( .A(n31159), .B(g_input[977]), .Z(n31156) );
  NAND U31260 ( .A(n31160), .B(mul_pow), .Z(n31159) );
  XOR U31261 ( .A(g_input[977]), .B(creg[977]), .Z(n31160) );
  XOR U31262 ( .A(n31161), .B(n31162), .Z(n31152) );
  ANDN U31263 ( .A(n31163), .B(n24884), .Z(n31162) );
  XOR U31264 ( .A(n31164), .B(\modmult_1/zin[0][975] ), .Z(n24884) );
  IV U31265 ( .A(n31161), .Z(n31164) );
  XNOR U31266 ( .A(n31161), .B(n24883), .Z(n31163) );
  XOR U31267 ( .A(n31165), .B(n31166), .Z(n24883) );
  AND U31268 ( .A(\modmult_1/xin[1023] ), .B(n31167), .Z(n31166) );
  IV U31269 ( .A(n31165), .Z(n31167) );
  XOR U31270 ( .A(n31168), .B(g_input[976]), .Z(n31165) );
  NAND U31271 ( .A(n31169), .B(mul_pow), .Z(n31168) );
  XOR U31272 ( .A(g_input[976]), .B(creg[976]), .Z(n31169) );
  XOR U31273 ( .A(n31170), .B(n31171), .Z(n31161) );
  ANDN U31274 ( .A(n31172), .B(n24890), .Z(n31171) );
  XOR U31275 ( .A(n31173), .B(\modmult_1/zin[0][974] ), .Z(n24890) );
  IV U31276 ( .A(n31170), .Z(n31173) );
  XNOR U31277 ( .A(n31170), .B(n24889), .Z(n31172) );
  XOR U31278 ( .A(n31174), .B(n31175), .Z(n24889) );
  AND U31279 ( .A(\modmult_1/xin[1023] ), .B(n31176), .Z(n31175) );
  IV U31280 ( .A(n31174), .Z(n31176) );
  XOR U31281 ( .A(n31177), .B(g_input[975]), .Z(n31174) );
  NAND U31282 ( .A(n31178), .B(mul_pow), .Z(n31177) );
  XOR U31283 ( .A(g_input[975]), .B(creg[975]), .Z(n31178) );
  XOR U31284 ( .A(n31179), .B(n31180), .Z(n31170) );
  ANDN U31285 ( .A(n31181), .B(n24896), .Z(n31180) );
  XOR U31286 ( .A(n31182), .B(\modmult_1/zin[0][973] ), .Z(n24896) );
  IV U31287 ( .A(n31179), .Z(n31182) );
  XNOR U31288 ( .A(n31179), .B(n24895), .Z(n31181) );
  XOR U31289 ( .A(n31183), .B(n31184), .Z(n24895) );
  AND U31290 ( .A(\modmult_1/xin[1023] ), .B(n31185), .Z(n31184) );
  IV U31291 ( .A(n31183), .Z(n31185) );
  XOR U31292 ( .A(n31186), .B(g_input[974]), .Z(n31183) );
  NAND U31293 ( .A(n31187), .B(mul_pow), .Z(n31186) );
  XOR U31294 ( .A(g_input[974]), .B(creg[974]), .Z(n31187) );
  XOR U31295 ( .A(n31188), .B(n31189), .Z(n31179) );
  ANDN U31296 ( .A(n31190), .B(n24902), .Z(n31189) );
  XOR U31297 ( .A(n31191), .B(\modmult_1/zin[0][972] ), .Z(n24902) );
  IV U31298 ( .A(n31188), .Z(n31191) );
  XNOR U31299 ( .A(n31188), .B(n24901), .Z(n31190) );
  XOR U31300 ( .A(n31192), .B(n31193), .Z(n24901) );
  AND U31301 ( .A(\modmult_1/xin[1023] ), .B(n31194), .Z(n31193) );
  IV U31302 ( .A(n31192), .Z(n31194) );
  XOR U31303 ( .A(n31195), .B(g_input[973]), .Z(n31192) );
  NAND U31304 ( .A(n31196), .B(mul_pow), .Z(n31195) );
  XOR U31305 ( .A(g_input[973]), .B(creg[973]), .Z(n31196) );
  XOR U31306 ( .A(n31197), .B(n31198), .Z(n31188) );
  ANDN U31307 ( .A(n31199), .B(n24908), .Z(n31198) );
  XOR U31308 ( .A(n31200), .B(\modmult_1/zin[0][971] ), .Z(n24908) );
  IV U31309 ( .A(n31197), .Z(n31200) );
  XNOR U31310 ( .A(n31197), .B(n24907), .Z(n31199) );
  XOR U31311 ( .A(n31201), .B(n31202), .Z(n24907) );
  AND U31312 ( .A(\modmult_1/xin[1023] ), .B(n31203), .Z(n31202) );
  IV U31313 ( .A(n31201), .Z(n31203) );
  XOR U31314 ( .A(n31204), .B(g_input[972]), .Z(n31201) );
  NAND U31315 ( .A(n31205), .B(mul_pow), .Z(n31204) );
  XOR U31316 ( .A(g_input[972]), .B(creg[972]), .Z(n31205) );
  XOR U31317 ( .A(n31206), .B(n31207), .Z(n31197) );
  ANDN U31318 ( .A(n31208), .B(n24914), .Z(n31207) );
  XOR U31319 ( .A(n31209), .B(\modmult_1/zin[0][970] ), .Z(n24914) );
  IV U31320 ( .A(n31206), .Z(n31209) );
  XNOR U31321 ( .A(n31206), .B(n24913), .Z(n31208) );
  XOR U31322 ( .A(n31210), .B(n31211), .Z(n24913) );
  AND U31323 ( .A(\modmult_1/xin[1023] ), .B(n31212), .Z(n31211) );
  IV U31324 ( .A(n31210), .Z(n31212) );
  XOR U31325 ( .A(n31213), .B(g_input[971]), .Z(n31210) );
  NAND U31326 ( .A(n31214), .B(mul_pow), .Z(n31213) );
  XOR U31327 ( .A(g_input[971]), .B(creg[971]), .Z(n31214) );
  XOR U31328 ( .A(n31215), .B(n31216), .Z(n31206) );
  ANDN U31329 ( .A(n31217), .B(n24920), .Z(n31216) );
  XOR U31330 ( .A(n31218), .B(\modmult_1/zin[0][969] ), .Z(n24920) );
  IV U31331 ( .A(n31215), .Z(n31218) );
  XNOR U31332 ( .A(n31215), .B(n24919), .Z(n31217) );
  XOR U31333 ( .A(n31219), .B(n31220), .Z(n24919) );
  AND U31334 ( .A(\modmult_1/xin[1023] ), .B(n31221), .Z(n31220) );
  IV U31335 ( .A(n31219), .Z(n31221) );
  XOR U31336 ( .A(n31222), .B(g_input[970]), .Z(n31219) );
  NAND U31337 ( .A(n31223), .B(mul_pow), .Z(n31222) );
  XOR U31338 ( .A(g_input[970]), .B(creg[970]), .Z(n31223) );
  XOR U31339 ( .A(n31224), .B(n31225), .Z(n31215) );
  ANDN U31340 ( .A(n31226), .B(n24926), .Z(n31225) );
  XOR U31341 ( .A(n31227), .B(\modmult_1/zin[0][968] ), .Z(n24926) );
  IV U31342 ( .A(n31224), .Z(n31227) );
  XNOR U31343 ( .A(n31224), .B(n24925), .Z(n31226) );
  XOR U31344 ( .A(n31228), .B(n31229), .Z(n24925) );
  AND U31345 ( .A(\modmult_1/xin[1023] ), .B(n31230), .Z(n31229) );
  IV U31346 ( .A(n31228), .Z(n31230) );
  XOR U31347 ( .A(n31231), .B(g_input[969]), .Z(n31228) );
  NAND U31348 ( .A(n31232), .B(mul_pow), .Z(n31231) );
  XOR U31349 ( .A(g_input[969]), .B(creg[969]), .Z(n31232) );
  XOR U31350 ( .A(n31233), .B(n31234), .Z(n31224) );
  ANDN U31351 ( .A(n31235), .B(n24932), .Z(n31234) );
  XOR U31352 ( .A(n31236), .B(\modmult_1/zin[0][967] ), .Z(n24932) );
  IV U31353 ( .A(n31233), .Z(n31236) );
  XNOR U31354 ( .A(n31233), .B(n24931), .Z(n31235) );
  XOR U31355 ( .A(n31237), .B(n31238), .Z(n24931) );
  AND U31356 ( .A(\modmult_1/xin[1023] ), .B(n31239), .Z(n31238) );
  IV U31357 ( .A(n31237), .Z(n31239) );
  XOR U31358 ( .A(n31240), .B(g_input[968]), .Z(n31237) );
  NAND U31359 ( .A(n31241), .B(mul_pow), .Z(n31240) );
  XOR U31360 ( .A(g_input[968]), .B(creg[968]), .Z(n31241) );
  XOR U31361 ( .A(n31242), .B(n31243), .Z(n31233) );
  ANDN U31362 ( .A(n31244), .B(n24938), .Z(n31243) );
  XOR U31363 ( .A(n31245), .B(\modmult_1/zin[0][966] ), .Z(n24938) );
  IV U31364 ( .A(n31242), .Z(n31245) );
  XNOR U31365 ( .A(n31242), .B(n24937), .Z(n31244) );
  XOR U31366 ( .A(n31246), .B(n31247), .Z(n24937) );
  AND U31367 ( .A(\modmult_1/xin[1023] ), .B(n31248), .Z(n31247) );
  IV U31368 ( .A(n31246), .Z(n31248) );
  XOR U31369 ( .A(n31249), .B(g_input[967]), .Z(n31246) );
  NAND U31370 ( .A(n31250), .B(mul_pow), .Z(n31249) );
  XOR U31371 ( .A(g_input[967]), .B(creg[967]), .Z(n31250) );
  XOR U31372 ( .A(n31251), .B(n31252), .Z(n31242) );
  ANDN U31373 ( .A(n31253), .B(n24944), .Z(n31252) );
  XOR U31374 ( .A(n31254), .B(\modmult_1/zin[0][965] ), .Z(n24944) );
  IV U31375 ( .A(n31251), .Z(n31254) );
  XNOR U31376 ( .A(n31251), .B(n24943), .Z(n31253) );
  XOR U31377 ( .A(n31255), .B(n31256), .Z(n24943) );
  AND U31378 ( .A(\modmult_1/xin[1023] ), .B(n31257), .Z(n31256) );
  IV U31379 ( .A(n31255), .Z(n31257) );
  XOR U31380 ( .A(n31258), .B(g_input[966]), .Z(n31255) );
  NAND U31381 ( .A(n31259), .B(mul_pow), .Z(n31258) );
  XOR U31382 ( .A(g_input[966]), .B(creg[966]), .Z(n31259) );
  XOR U31383 ( .A(n31260), .B(n31261), .Z(n31251) );
  ANDN U31384 ( .A(n31262), .B(n24950), .Z(n31261) );
  XOR U31385 ( .A(n31263), .B(\modmult_1/zin[0][964] ), .Z(n24950) );
  IV U31386 ( .A(n31260), .Z(n31263) );
  XNOR U31387 ( .A(n31260), .B(n24949), .Z(n31262) );
  XOR U31388 ( .A(n31264), .B(n31265), .Z(n24949) );
  AND U31389 ( .A(\modmult_1/xin[1023] ), .B(n31266), .Z(n31265) );
  IV U31390 ( .A(n31264), .Z(n31266) );
  XOR U31391 ( .A(n31267), .B(g_input[965]), .Z(n31264) );
  NAND U31392 ( .A(n31268), .B(mul_pow), .Z(n31267) );
  XOR U31393 ( .A(g_input[965]), .B(creg[965]), .Z(n31268) );
  XOR U31394 ( .A(n31269), .B(n31270), .Z(n31260) );
  ANDN U31395 ( .A(n31271), .B(n24956), .Z(n31270) );
  XOR U31396 ( .A(n31272), .B(\modmult_1/zin[0][963] ), .Z(n24956) );
  IV U31397 ( .A(n31269), .Z(n31272) );
  XNOR U31398 ( .A(n31269), .B(n24955), .Z(n31271) );
  XOR U31399 ( .A(n31273), .B(n31274), .Z(n24955) );
  AND U31400 ( .A(\modmult_1/xin[1023] ), .B(n31275), .Z(n31274) );
  IV U31401 ( .A(n31273), .Z(n31275) );
  XOR U31402 ( .A(n31276), .B(g_input[964]), .Z(n31273) );
  NAND U31403 ( .A(n31277), .B(mul_pow), .Z(n31276) );
  XOR U31404 ( .A(g_input[964]), .B(creg[964]), .Z(n31277) );
  XOR U31405 ( .A(n31278), .B(n31279), .Z(n31269) );
  ANDN U31406 ( .A(n31280), .B(n24962), .Z(n31279) );
  XOR U31407 ( .A(n31281), .B(\modmult_1/zin[0][962] ), .Z(n24962) );
  IV U31408 ( .A(n31278), .Z(n31281) );
  XNOR U31409 ( .A(n31278), .B(n24961), .Z(n31280) );
  XOR U31410 ( .A(n31282), .B(n31283), .Z(n24961) );
  AND U31411 ( .A(\modmult_1/xin[1023] ), .B(n31284), .Z(n31283) );
  IV U31412 ( .A(n31282), .Z(n31284) );
  XOR U31413 ( .A(n31285), .B(g_input[963]), .Z(n31282) );
  NAND U31414 ( .A(n31286), .B(mul_pow), .Z(n31285) );
  XOR U31415 ( .A(g_input[963]), .B(creg[963]), .Z(n31286) );
  XOR U31416 ( .A(n31287), .B(n31288), .Z(n31278) );
  ANDN U31417 ( .A(n31289), .B(n24968), .Z(n31288) );
  XOR U31418 ( .A(n31290), .B(\modmult_1/zin[0][961] ), .Z(n24968) );
  IV U31419 ( .A(n31287), .Z(n31290) );
  XNOR U31420 ( .A(n31287), .B(n24967), .Z(n31289) );
  XOR U31421 ( .A(n31291), .B(n31292), .Z(n24967) );
  AND U31422 ( .A(\modmult_1/xin[1023] ), .B(n31293), .Z(n31292) );
  IV U31423 ( .A(n31291), .Z(n31293) );
  XOR U31424 ( .A(n31294), .B(g_input[962]), .Z(n31291) );
  NAND U31425 ( .A(n31295), .B(mul_pow), .Z(n31294) );
  XOR U31426 ( .A(g_input[962]), .B(creg[962]), .Z(n31295) );
  XOR U31427 ( .A(n31296), .B(n31297), .Z(n31287) );
  ANDN U31428 ( .A(n31298), .B(n24974), .Z(n31297) );
  XOR U31429 ( .A(n31299), .B(\modmult_1/zin[0][960] ), .Z(n24974) );
  IV U31430 ( .A(n31296), .Z(n31299) );
  XNOR U31431 ( .A(n31296), .B(n24973), .Z(n31298) );
  XOR U31432 ( .A(n31300), .B(n31301), .Z(n24973) );
  AND U31433 ( .A(\modmult_1/xin[1023] ), .B(n31302), .Z(n31301) );
  IV U31434 ( .A(n31300), .Z(n31302) );
  XOR U31435 ( .A(n31303), .B(g_input[961]), .Z(n31300) );
  NAND U31436 ( .A(n31304), .B(mul_pow), .Z(n31303) );
  XOR U31437 ( .A(g_input[961]), .B(creg[961]), .Z(n31304) );
  XOR U31438 ( .A(n31305), .B(n31306), .Z(n31296) );
  ANDN U31439 ( .A(n31307), .B(n24980), .Z(n31306) );
  XOR U31440 ( .A(n31308), .B(\modmult_1/zin[0][959] ), .Z(n24980) );
  IV U31441 ( .A(n31305), .Z(n31308) );
  XNOR U31442 ( .A(n31305), .B(n24979), .Z(n31307) );
  XOR U31443 ( .A(n31309), .B(n31310), .Z(n24979) );
  AND U31444 ( .A(\modmult_1/xin[1023] ), .B(n31311), .Z(n31310) );
  IV U31445 ( .A(n31309), .Z(n31311) );
  XOR U31446 ( .A(n31312), .B(g_input[960]), .Z(n31309) );
  NAND U31447 ( .A(n31313), .B(mul_pow), .Z(n31312) );
  XOR U31448 ( .A(g_input[960]), .B(creg[960]), .Z(n31313) );
  XOR U31449 ( .A(n31314), .B(n31315), .Z(n31305) );
  ANDN U31450 ( .A(n31316), .B(n24986), .Z(n31315) );
  XOR U31451 ( .A(n31317), .B(\modmult_1/zin[0][958] ), .Z(n24986) );
  IV U31452 ( .A(n31314), .Z(n31317) );
  XNOR U31453 ( .A(n31314), .B(n24985), .Z(n31316) );
  XOR U31454 ( .A(n31318), .B(n31319), .Z(n24985) );
  AND U31455 ( .A(\modmult_1/xin[1023] ), .B(n31320), .Z(n31319) );
  IV U31456 ( .A(n31318), .Z(n31320) );
  XOR U31457 ( .A(n31321), .B(g_input[959]), .Z(n31318) );
  NAND U31458 ( .A(n31322), .B(mul_pow), .Z(n31321) );
  XOR U31459 ( .A(g_input[959]), .B(creg[959]), .Z(n31322) );
  XOR U31460 ( .A(n31323), .B(n31324), .Z(n31314) );
  ANDN U31461 ( .A(n31325), .B(n24992), .Z(n31324) );
  XOR U31462 ( .A(n31326), .B(\modmult_1/zin[0][957] ), .Z(n24992) );
  IV U31463 ( .A(n31323), .Z(n31326) );
  XNOR U31464 ( .A(n31323), .B(n24991), .Z(n31325) );
  XOR U31465 ( .A(n31327), .B(n31328), .Z(n24991) );
  AND U31466 ( .A(\modmult_1/xin[1023] ), .B(n31329), .Z(n31328) );
  IV U31467 ( .A(n31327), .Z(n31329) );
  XOR U31468 ( .A(n31330), .B(g_input[958]), .Z(n31327) );
  NAND U31469 ( .A(n31331), .B(mul_pow), .Z(n31330) );
  XOR U31470 ( .A(g_input[958]), .B(creg[958]), .Z(n31331) );
  XOR U31471 ( .A(n31332), .B(n31333), .Z(n31323) );
  ANDN U31472 ( .A(n31334), .B(n24998), .Z(n31333) );
  XOR U31473 ( .A(n31335), .B(\modmult_1/zin[0][956] ), .Z(n24998) );
  IV U31474 ( .A(n31332), .Z(n31335) );
  XNOR U31475 ( .A(n31332), .B(n24997), .Z(n31334) );
  XOR U31476 ( .A(n31336), .B(n31337), .Z(n24997) );
  AND U31477 ( .A(\modmult_1/xin[1023] ), .B(n31338), .Z(n31337) );
  IV U31478 ( .A(n31336), .Z(n31338) );
  XOR U31479 ( .A(n31339), .B(g_input[957]), .Z(n31336) );
  NAND U31480 ( .A(n31340), .B(mul_pow), .Z(n31339) );
  XOR U31481 ( .A(g_input[957]), .B(creg[957]), .Z(n31340) );
  XOR U31482 ( .A(n31341), .B(n31342), .Z(n31332) );
  ANDN U31483 ( .A(n31343), .B(n25004), .Z(n31342) );
  XOR U31484 ( .A(n31344), .B(\modmult_1/zin[0][955] ), .Z(n25004) );
  IV U31485 ( .A(n31341), .Z(n31344) );
  XNOR U31486 ( .A(n31341), .B(n25003), .Z(n31343) );
  XOR U31487 ( .A(n31345), .B(n31346), .Z(n25003) );
  AND U31488 ( .A(\modmult_1/xin[1023] ), .B(n31347), .Z(n31346) );
  IV U31489 ( .A(n31345), .Z(n31347) );
  XOR U31490 ( .A(n31348), .B(g_input[956]), .Z(n31345) );
  NAND U31491 ( .A(n31349), .B(mul_pow), .Z(n31348) );
  XOR U31492 ( .A(g_input[956]), .B(creg[956]), .Z(n31349) );
  XOR U31493 ( .A(n31350), .B(n31351), .Z(n31341) );
  ANDN U31494 ( .A(n31352), .B(n25010), .Z(n31351) );
  XOR U31495 ( .A(n31353), .B(\modmult_1/zin[0][954] ), .Z(n25010) );
  IV U31496 ( .A(n31350), .Z(n31353) );
  XNOR U31497 ( .A(n31350), .B(n25009), .Z(n31352) );
  XOR U31498 ( .A(n31354), .B(n31355), .Z(n25009) );
  AND U31499 ( .A(\modmult_1/xin[1023] ), .B(n31356), .Z(n31355) );
  IV U31500 ( .A(n31354), .Z(n31356) );
  XOR U31501 ( .A(n31357), .B(g_input[955]), .Z(n31354) );
  NAND U31502 ( .A(n31358), .B(mul_pow), .Z(n31357) );
  XOR U31503 ( .A(g_input[955]), .B(creg[955]), .Z(n31358) );
  XOR U31504 ( .A(n31359), .B(n31360), .Z(n31350) );
  ANDN U31505 ( .A(n31361), .B(n25016), .Z(n31360) );
  XOR U31506 ( .A(n31362), .B(\modmult_1/zin[0][953] ), .Z(n25016) );
  IV U31507 ( .A(n31359), .Z(n31362) );
  XNOR U31508 ( .A(n31359), .B(n25015), .Z(n31361) );
  XOR U31509 ( .A(n31363), .B(n31364), .Z(n25015) );
  AND U31510 ( .A(\modmult_1/xin[1023] ), .B(n31365), .Z(n31364) );
  IV U31511 ( .A(n31363), .Z(n31365) );
  XOR U31512 ( .A(n31366), .B(g_input[954]), .Z(n31363) );
  NAND U31513 ( .A(n31367), .B(mul_pow), .Z(n31366) );
  XOR U31514 ( .A(g_input[954]), .B(creg[954]), .Z(n31367) );
  XOR U31515 ( .A(n31368), .B(n31369), .Z(n31359) );
  ANDN U31516 ( .A(n31370), .B(n25022), .Z(n31369) );
  XOR U31517 ( .A(n31371), .B(\modmult_1/zin[0][952] ), .Z(n25022) );
  IV U31518 ( .A(n31368), .Z(n31371) );
  XNOR U31519 ( .A(n31368), .B(n25021), .Z(n31370) );
  XOR U31520 ( .A(n31372), .B(n31373), .Z(n25021) );
  AND U31521 ( .A(\modmult_1/xin[1023] ), .B(n31374), .Z(n31373) );
  IV U31522 ( .A(n31372), .Z(n31374) );
  XOR U31523 ( .A(n31375), .B(g_input[953]), .Z(n31372) );
  NAND U31524 ( .A(n31376), .B(mul_pow), .Z(n31375) );
  XOR U31525 ( .A(g_input[953]), .B(creg[953]), .Z(n31376) );
  XOR U31526 ( .A(n31377), .B(n31378), .Z(n31368) );
  ANDN U31527 ( .A(n31379), .B(n25028), .Z(n31378) );
  XOR U31528 ( .A(n31380), .B(\modmult_1/zin[0][951] ), .Z(n25028) );
  IV U31529 ( .A(n31377), .Z(n31380) );
  XNOR U31530 ( .A(n31377), .B(n25027), .Z(n31379) );
  XOR U31531 ( .A(n31381), .B(n31382), .Z(n25027) );
  AND U31532 ( .A(\modmult_1/xin[1023] ), .B(n31383), .Z(n31382) );
  IV U31533 ( .A(n31381), .Z(n31383) );
  XOR U31534 ( .A(n31384), .B(g_input[952]), .Z(n31381) );
  NAND U31535 ( .A(n31385), .B(mul_pow), .Z(n31384) );
  XOR U31536 ( .A(g_input[952]), .B(creg[952]), .Z(n31385) );
  XOR U31537 ( .A(n31386), .B(n31387), .Z(n31377) );
  ANDN U31538 ( .A(n31388), .B(n25034), .Z(n31387) );
  XOR U31539 ( .A(n31389), .B(\modmult_1/zin[0][950] ), .Z(n25034) );
  IV U31540 ( .A(n31386), .Z(n31389) );
  XNOR U31541 ( .A(n31386), .B(n25033), .Z(n31388) );
  XOR U31542 ( .A(n31390), .B(n31391), .Z(n25033) );
  AND U31543 ( .A(\modmult_1/xin[1023] ), .B(n31392), .Z(n31391) );
  IV U31544 ( .A(n31390), .Z(n31392) );
  XOR U31545 ( .A(n31393), .B(g_input[951]), .Z(n31390) );
  NAND U31546 ( .A(n31394), .B(mul_pow), .Z(n31393) );
  XOR U31547 ( .A(g_input[951]), .B(creg[951]), .Z(n31394) );
  XOR U31548 ( .A(n31395), .B(n31396), .Z(n31386) );
  ANDN U31549 ( .A(n31397), .B(n25040), .Z(n31396) );
  XOR U31550 ( .A(n31398), .B(\modmult_1/zin[0][949] ), .Z(n25040) );
  IV U31551 ( .A(n31395), .Z(n31398) );
  XNOR U31552 ( .A(n31395), .B(n25039), .Z(n31397) );
  XOR U31553 ( .A(n31399), .B(n31400), .Z(n25039) );
  AND U31554 ( .A(\modmult_1/xin[1023] ), .B(n31401), .Z(n31400) );
  IV U31555 ( .A(n31399), .Z(n31401) );
  XOR U31556 ( .A(n31402), .B(g_input[950]), .Z(n31399) );
  NAND U31557 ( .A(n31403), .B(mul_pow), .Z(n31402) );
  XOR U31558 ( .A(g_input[950]), .B(creg[950]), .Z(n31403) );
  XOR U31559 ( .A(n31404), .B(n31405), .Z(n31395) );
  ANDN U31560 ( .A(n31406), .B(n25046), .Z(n31405) );
  XOR U31561 ( .A(n31407), .B(\modmult_1/zin[0][948] ), .Z(n25046) );
  IV U31562 ( .A(n31404), .Z(n31407) );
  XNOR U31563 ( .A(n31404), .B(n25045), .Z(n31406) );
  XOR U31564 ( .A(n31408), .B(n31409), .Z(n25045) );
  AND U31565 ( .A(\modmult_1/xin[1023] ), .B(n31410), .Z(n31409) );
  IV U31566 ( .A(n31408), .Z(n31410) );
  XOR U31567 ( .A(n31411), .B(g_input[949]), .Z(n31408) );
  NAND U31568 ( .A(n31412), .B(mul_pow), .Z(n31411) );
  XOR U31569 ( .A(g_input[949]), .B(creg[949]), .Z(n31412) );
  XOR U31570 ( .A(n31413), .B(n31414), .Z(n31404) );
  ANDN U31571 ( .A(n31415), .B(n25052), .Z(n31414) );
  XOR U31572 ( .A(n31416), .B(\modmult_1/zin[0][947] ), .Z(n25052) );
  IV U31573 ( .A(n31413), .Z(n31416) );
  XNOR U31574 ( .A(n31413), .B(n25051), .Z(n31415) );
  XOR U31575 ( .A(n31417), .B(n31418), .Z(n25051) );
  AND U31576 ( .A(\modmult_1/xin[1023] ), .B(n31419), .Z(n31418) );
  IV U31577 ( .A(n31417), .Z(n31419) );
  XOR U31578 ( .A(n31420), .B(g_input[948]), .Z(n31417) );
  NAND U31579 ( .A(n31421), .B(mul_pow), .Z(n31420) );
  XOR U31580 ( .A(g_input[948]), .B(creg[948]), .Z(n31421) );
  XOR U31581 ( .A(n31422), .B(n31423), .Z(n31413) );
  ANDN U31582 ( .A(n31424), .B(n25058), .Z(n31423) );
  XOR U31583 ( .A(n31425), .B(\modmult_1/zin[0][946] ), .Z(n25058) );
  IV U31584 ( .A(n31422), .Z(n31425) );
  XNOR U31585 ( .A(n31422), .B(n25057), .Z(n31424) );
  XOR U31586 ( .A(n31426), .B(n31427), .Z(n25057) );
  AND U31587 ( .A(\modmult_1/xin[1023] ), .B(n31428), .Z(n31427) );
  IV U31588 ( .A(n31426), .Z(n31428) );
  XOR U31589 ( .A(n31429), .B(g_input[947]), .Z(n31426) );
  NAND U31590 ( .A(n31430), .B(mul_pow), .Z(n31429) );
  XOR U31591 ( .A(g_input[947]), .B(creg[947]), .Z(n31430) );
  XOR U31592 ( .A(n31431), .B(n31432), .Z(n31422) );
  ANDN U31593 ( .A(n31433), .B(n25064), .Z(n31432) );
  XOR U31594 ( .A(n31434), .B(\modmult_1/zin[0][945] ), .Z(n25064) );
  IV U31595 ( .A(n31431), .Z(n31434) );
  XNOR U31596 ( .A(n31431), .B(n25063), .Z(n31433) );
  XOR U31597 ( .A(n31435), .B(n31436), .Z(n25063) );
  AND U31598 ( .A(\modmult_1/xin[1023] ), .B(n31437), .Z(n31436) );
  IV U31599 ( .A(n31435), .Z(n31437) );
  XOR U31600 ( .A(n31438), .B(g_input[946]), .Z(n31435) );
  NAND U31601 ( .A(n31439), .B(mul_pow), .Z(n31438) );
  XOR U31602 ( .A(g_input[946]), .B(creg[946]), .Z(n31439) );
  XOR U31603 ( .A(n31440), .B(n31441), .Z(n31431) );
  ANDN U31604 ( .A(n31442), .B(n25070), .Z(n31441) );
  XOR U31605 ( .A(n31443), .B(\modmult_1/zin[0][944] ), .Z(n25070) );
  IV U31606 ( .A(n31440), .Z(n31443) );
  XNOR U31607 ( .A(n31440), .B(n25069), .Z(n31442) );
  XOR U31608 ( .A(n31444), .B(n31445), .Z(n25069) );
  AND U31609 ( .A(\modmult_1/xin[1023] ), .B(n31446), .Z(n31445) );
  IV U31610 ( .A(n31444), .Z(n31446) );
  XOR U31611 ( .A(n31447), .B(g_input[945]), .Z(n31444) );
  NAND U31612 ( .A(n31448), .B(mul_pow), .Z(n31447) );
  XOR U31613 ( .A(g_input[945]), .B(creg[945]), .Z(n31448) );
  XOR U31614 ( .A(n31449), .B(n31450), .Z(n31440) );
  ANDN U31615 ( .A(n31451), .B(n25076), .Z(n31450) );
  XOR U31616 ( .A(n31452), .B(\modmult_1/zin[0][943] ), .Z(n25076) );
  IV U31617 ( .A(n31449), .Z(n31452) );
  XNOR U31618 ( .A(n31449), .B(n25075), .Z(n31451) );
  XOR U31619 ( .A(n31453), .B(n31454), .Z(n25075) );
  AND U31620 ( .A(\modmult_1/xin[1023] ), .B(n31455), .Z(n31454) );
  IV U31621 ( .A(n31453), .Z(n31455) );
  XOR U31622 ( .A(n31456), .B(g_input[944]), .Z(n31453) );
  NAND U31623 ( .A(n31457), .B(mul_pow), .Z(n31456) );
  XOR U31624 ( .A(g_input[944]), .B(creg[944]), .Z(n31457) );
  XOR U31625 ( .A(n31458), .B(n31459), .Z(n31449) );
  ANDN U31626 ( .A(n31460), .B(n25082), .Z(n31459) );
  XOR U31627 ( .A(n31461), .B(\modmult_1/zin[0][942] ), .Z(n25082) );
  IV U31628 ( .A(n31458), .Z(n31461) );
  XNOR U31629 ( .A(n31458), .B(n25081), .Z(n31460) );
  XOR U31630 ( .A(n31462), .B(n31463), .Z(n25081) );
  AND U31631 ( .A(\modmult_1/xin[1023] ), .B(n31464), .Z(n31463) );
  IV U31632 ( .A(n31462), .Z(n31464) );
  XOR U31633 ( .A(n31465), .B(g_input[943]), .Z(n31462) );
  NAND U31634 ( .A(n31466), .B(mul_pow), .Z(n31465) );
  XOR U31635 ( .A(g_input[943]), .B(creg[943]), .Z(n31466) );
  XOR U31636 ( .A(n31467), .B(n31468), .Z(n31458) );
  ANDN U31637 ( .A(n31469), .B(n25088), .Z(n31468) );
  XOR U31638 ( .A(n31470), .B(\modmult_1/zin[0][941] ), .Z(n25088) );
  IV U31639 ( .A(n31467), .Z(n31470) );
  XNOR U31640 ( .A(n31467), .B(n25087), .Z(n31469) );
  XOR U31641 ( .A(n31471), .B(n31472), .Z(n25087) );
  AND U31642 ( .A(\modmult_1/xin[1023] ), .B(n31473), .Z(n31472) );
  IV U31643 ( .A(n31471), .Z(n31473) );
  XOR U31644 ( .A(n31474), .B(g_input[942]), .Z(n31471) );
  NAND U31645 ( .A(n31475), .B(mul_pow), .Z(n31474) );
  XOR U31646 ( .A(g_input[942]), .B(creg[942]), .Z(n31475) );
  XOR U31647 ( .A(n31476), .B(n31477), .Z(n31467) );
  ANDN U31648 ( .A(n31478), .B(n25094), .Z(n31477) );
  XOR U31649 ( .A(n31479), .B(\modmult_1/zin[0][940] ), .Z(n25094) );
  IV U31650 ( .A(n31476), .Z(n31479) );
  XNOR U31651 ( .A(n31476), .B(n25093), .Z(n31478) );
  XOR U31652 ( .A(n31480), .B(n31481), .Z(n25093) );
  AND U31653 ( .A(\modmult_1/xin[1023] ), .B(n31482), .Z(n31481) );
  IV U31654 ( .A(n31480), .Z(n31482) );
  XOR U31655 ( .A(n31483), .B(g_input[941]), .Z(n31480) );
  NAND U31656 ( .A(n31484), .B(mul_pow), .Z(n31483) );
  XOR U31657 ( .A(g_input[941]), .B(creg[941]), .Z(n31484) );
  XOR U31658 ( .A(n31485), .B(n31486), .Z(n31476) );
  ANDN U31659 ( .A(n31487), .B(n25100), .Z(n31486) );
  XOR U31660 ( .A(n31488), .B(\modmult_1/zin[0][939] ), .Z(n25100) );
  IV U31661 ( .A(n31485), .Z(n31488) );
  XNOR U31662 ( .A(n31485), .B(n25099), .Z(n31487) );
  XOR U31663 ( .A(n31489), .B(n31490), .Z(n25099) );
  AND U31664 ( .A(\modmult_1/xin[1023] ), .B(n31491), .Z(n31490) );
  IV U31665 ( .A(n31489), .Z(n31491) );
  XOR U31666 ( .A(n31492), .B(g_input[940]), .Z(n31489) );
  NAND U31667 ( .A(n31493), .B(mul_pow), .Z(n31492) );
  XOR U31668 ( .A(g_input[940]), .B(creg[940]), .Z(n31493) );
  XOR U31669 ( .A(n31494), .B(n31495), .Z(n31485) );
  ANDN U31670 ( .A(n31496), .B(n25106), .Z(n31495) );
  XOR U31671 ( .A(n31497), .B(\modmult_1/zin[0][938] ), .Z(n25106) );
  IV U31672 ( .A(n31494), .Z(n31497) );
  XNOR U31673 ( .A(n31494), .B(n25105), .Z(n31496) );
  XOR U31674 ( .A(n31498), .B(n31499), .Z(n25105) );
  AND U31675 ( .A(\modmult_1/xin[1023] ), .B(n31500), .Z(n31499) );
  IV U31676 ( .A(n31498), .Z(n31500) );
  XOR U31677 ( .A(n31501), .B(g_input[939]), .Z(n31498) );
  NAND U31678 ( .A(n31502), .B(mul_pow), .Z(n31501) );
  XOR U31679 ( .A(g_input[939]), .B(creg[939]), .Z(n31502) );
  XOR U31680 ( .A(n31503), .B(n31504), .Z(n31494) );
  ANDN U31681 ( .A(n31505), .B(n25112), .Z(n31504) );
  XOR U31682 ( .A(n31506), .B(\modmult_1/zin[0][937] ), .Z(n25112) );
  IV U31683 ( .A(n31503), .Z(n31506) );
  XNOR U31684 ( .A(n31503), .B(n25111), .Z(n31505) );
  XOR U31685 ( .A(n31507), .B(n31508), .Z(n25111) );
  AND U31686 ( .A(\modmult_1/xin[1023] ), .B(n31509), .Z(n31508) );
  IV U31687 ( .A(n31507), .Z(n31509) );
  XOR U31688 ( .A(n31510), .B(g_input[938]), .Z(n31507) );
  NAND U31689 ( .A(n31511), .B(mul_pow), .Z(n31510) );
  XOR U31690 ( .A(g_input[938]), .B(creg[938]), .Z(n31511) );
  XOR U31691 ( .A(n31512), .B(n31513), .Z(n31503) );
  ANDN U31692 ( .A(n31514), .B(n25118), .Z(n31513) );
  XOR U31693 ( .A(n31515), .B(\modmult_1/zin[0][936] ), .Z(n25118) );
  IV U31694 ( .A(n31512), .Z(n31515) );
  XNOR U31695 ( .A(n31512), .B(n25117), .Z(n31514) );
  XOR U31696 ( .A(n31516), .B(n31517), .Z(n25117) );
  AND U31697 ( .A(\modmult_1/xin[1023] ), .B(n31518), .Z(n31517) );
  IV U31698 ( .A(n31516), .Z(n31518) );
  XOR U31699 ( .A(n31519), .B(g_input[937]), .Z(n31516) );
  NAND U31700 ( .A(n31520), .B(mul_pow), .Z(n31519) );
  XOR U31701 ( .A(g_input[937]), .B(creg[937]), .Z(n31520) );
  XOR U31702 ( .A(n31521), .B(n31522), .Z(n31512) );
  ANDN U31703 ( .A(n31523), .B(n25124), .Z(n31522) );
  XOR U31704 ( .A(n31524), .B(\modmult_1/zin[0][935] ), .Z(n25124) );
  IV U31705 ( .A(n31521), .Z(n31524) );
  XNOR U31706 ( .A(n31521), .B(n25123), .Z(n31523) );
  XOR U31707 ( .A(n31525), .B(n31526), .Z(n25123) );
  AND U31708 ( .A(\modmult_1/xin[1023] ), .B(n31527), .Z(n31526) );
  IV U31709 ( .A(n31525), .Z(n31527) );
  XOR U31710 ( .A(n31528), .B(g_input[936]), .Z(n31525) );
  NAND U31711 ( .A(n31529), .B(mul_pow), .Z(n31528) );
  XOR U31712 ( .A(g_input[936]), .B(creg[936]), .Z(n31529) );
  XOR U31713 ( .A(n31530), .B(n31531), .Z(n31521) );
  ANDN U31714 ( .A(n31532), .B(n25130), .Z(n31531) );
  XOR U31715 ( .A(n31533), .B(\modmult_1/zin[0][934] ), .Z(n25130) );
  IV U31716 ( .A(n31530), .Z(n31533) );
  XNOR U31717 ( .A(n31530), .B(n25129), .Z(n31532) );
  XOR U31718 ( .A(n31534), .B(n31535), .Z(n25129) );
  AND U31719 ( .A(\modmult_1/xin[1023] ), .B(n31536), .Z(n31535) );
  IV U31720 ( .A(n31534), .Z(n31536) );
  XOR U31721 ( .A(n31537), .B(g_input[935]), .Z(n31534) );
  NAND U31722 ( .A(n31538), .B(mul_pow), .Z(n31537) );
  XOR U31723 ( .A(g_input[935]), .B(creg[935]), .Z(n31538) );
  XOR U31724 ( .A(n31539), .B(n31540), .Z(n31530) );
  ANDN U31725 ( .A(n31541), .B(n25136), .Z(n31540) );
  XOR U31726 ( .A(n31542), .B(\modmult_1/zin[0][933] ), .Z(n25136) );
  IV U31727 ( .A(n31539), .Z(n31542) );
  XNOR U31728 ( .A(n31539), .B(n25135), .Z(n31541) );
  XOR U31729 ( .A(n31543), .B(n31544), .Z(n25135) );
  AND U31730 ( .A(\modmult_1/xin[1023] ), .B(n31545), .Z(n31544) );
  IV U31731 ( .A(n31543), .Z(n31545) );
  XOR U31732 ( .A(n31546), .B(g_input[934]), .Z(n31543) );
  NAND U31733 ( .A(n31547), .B(mul_pow), .Z(n31546) );
  XOR U31734 ( .A(g_input[934]), .B(creg[934]), .Z(n31547) );
  XOR U31735 ( .A(n31548), .B(n31549), .Z(n31539) );
  ANDN U31736 ( .A(n31550), .B(n25142), .Z(n31549) );
  XOR U31737 ( .A(n31551), .B(\modmult_1/zin[0][932] ), .Z(n25142) );
  IV U31738 ( .A(n31548), .Z(n31551) );
  XNOR U31739 ( .A(n31548), .B(n25141), .Z(n31550) );
  XOR U31740 ( .A(n31552), .B(n31553), .Z(n25141) );
  AND U31741 ( .A(\modmult_1/xin[1023] ), .B(n31554), .Z(n31553) );
  IV U31742 ( .A(n31552), .Z(n31554) );
  XOR U31743 ( .A(n31555), .B(g_input[933]), .Z(n31552) );
  NAND U31744 ( .A(n31556), .B(mul_pow), .Z(n31555) );
  XOR U31745 ( .A(g_input[933]), .B(creg[933]), .Z(n31556) );
  XOR U31746 ( .A(n31557), .B(n31558), .Z(n31548) );
  ANDN U31747 ( .A(n31559), .B(n25148), .Z(n31558) );
  XOR U31748 ( .A(n31560), .B(\modmult_1/zin[0][931] ), .Z(n25148) );
  IV U31749 ( .A(n31557), .Z(n31560) );
  XNOR U31750 ( .A(n31557), .B(n25147), .Z(n31559) );
  XOR U31751 ( .A(n31561), .B(n31562), .Z(n25147) );
  AND U31752 ( .A(\modmult_1/xin[1023] ), .B(n31563), .Z(n31562) );
  IV U31753 ( .A(n31561), .Z(n31563) );
  XOR U31754 ( .A(n31564), .B(g_input[932]), .Z(n31561) );
  NAND U31755 ( .A(n31565), .B(mul_pow), .Z(n31564) );
  XOR U31756 ( .A(g_input[932]), .B(creg[932]), .Z(n31565) );
  XOR U31757 ( .A(n31566), .B(n31567), .Z(n31557) );
  ANDN U31758 ( .A(n31568), .B(n25154), .Z(n31567) );
  XOR U31759 ( .A(n31569), .B(\modmult_1/zin[0][930] ), .Z(n25154) );
  IV U31760 ( .A(n31566), .Z(n31569) );
  XNOR U31761 ( .A(n31566), .B(n25153), .Z(n31568) );
  XOR U31762 ( .A(n31570), .B(n31571), .Z(n25153) );
  AND U31763 ( .A(\modmult_1/xin[1023] ), .B(n31572), .Z(n31571) );
  IV U31764 ( .A(n31570), .Z(n31572) );
  XOR U31765 ( .A(n31573), .B(g_input[931]), .Z(n31570) );
  NAND U31766 ( .A(n31574), .B(mul_pow), .Z(n31573) );
  XOR U31767 ( .A(g_input[931]), .B(creg[931]), .Z(n31574) );
  XOR U31768 ( .A(n31575), .B(n31576), .Z(n31566) );
  ANDN U31769 ( .A(n31577), .B(n25160), .Z(n31576) );
  XOR U31770 ( .A(n31578), .B(\modmult_1/zin[0][929] ), .Z(n25160) );
  IV U31771 ( .A(n31575), .Z(n31578) );
  XNOR U31772 ( .A(n31575), .B(n25159), .Z(n31577) );
  XOR U31773 ( .A(n31579), .B(n31580), .Z(n25159) );
  AND U31774 ( .A(\modmult_1/xin[1023] ), .B(n31581), .Z(n31580) );
  IV U31775 ( .A(n31579), .Z(n31581) );
  XOR U31776 ( .A(n31582), .B(g_input[930]), .Z(n31579) );
  NAND U31777 ( .A(n31583), .B(mul_pow), .Z(n31582) );
  XOR U31778 ( .A(g_input[930]), .B(creg[930]), .Z(n31583) );
  XOR U31779 ( .A(n31584), .B(n31585), .Z(n31575) );
  ANDN U31780 ( .A(n31586), .B(n25166), .Z(n31585) );
  XOR U31781 ( .A(n31587), .B(\modmult_1/zin[0][928] ), .Z(n25166) );
  IV U31782 ( .A(n31584), .Z(n31587) );
  XNOR U31783 ( .A(n31584), .B(n25165), .Z(n31586) );
  XOR U31784 ( .A(n31588), .B(n31589), .Z(n25165) );
  AND U31785 ( .A(\modmult_1/xin[1023] ), .B(n31590), .Z(n31589) );
  IV U31786 ( .A(n31588), .Z(n31590) );
  XOR U31787 ( .A(n31591), .B(g_input[929]), .Z(n31588) );
  NAND U31788 ( .A(n31592), .B(mul_pow), .Z(n31591) );
  XOR U31789 ( .A(g_input[929]), .B(creg[929]), .Z(n31592) );
  XOR U31790 ( .A(n31593), .B(n31594), .Z(n31584) );
  ANDN U31791 ( .A(n31595), .B(n25172), .Z(n31594) );
  XOR U31792 ( .A(n31596), .B(\modmult_1/zin[0][927] ), .Z(n25172) );
  IV U31793 ( .A(n31593), .Z(n31596) );
  XNOR U31794 ( .A(n31593), .B(n25171), .Z(n31595) );
  XOR U31795 ( .A(n31597), .B(n31598), .Z(n25171) );
  AND U31796 ( .A(\modmult_1/xin[1023] ), .B(n31599), .Z(n31598) );
  IV U31797 ( .A(n31597), .Z(n31599) );
  XOR U31798 ( .A(n31600), .B(g_input[928]), .Z(n31597) );
  NAND U31799 ( .A(n31601), .B(mul_pow), .Z(n31600) );
  XOR U31800 ( .A(g_input[928]), .B(creg[928]), .Z(n31601) );
  XOR U31801 ( .A(n31602), .B(n31603), .Z(n31593) );
  ANDN U31802 ( .A(n31604), .B(n25178), .Z(n31603) );
  XOR U31803 ( .A(n31605), .B(\modmult_1/zin[0][926] ), .Z(n25178) );
  IV U31804 ( .A(n31602), .Z(n31605) );
  XNOR U31805 ( .A(n31602), .B(n25177), .Z(n31604) );
  XOR U31806 ( .A(n31606), .B(n31607), .Z(n25177) );
  AND U31807 ( .A(\modmult_1/xin[1023] ), .B(n31608), .Z(n31607) );
  IV U31808 ( .A(n31606), .Z(n31608) );
  XOR U31809 ( .A(n31609), .B(g_input[927]), .Z(n31606) );
  NAND U31810 ( .A(n31610), .B(mul_pow), .Z(n31609) );
  XOR U31811 ( .A(g_input[927]), .B(creg[927]), .Z(n31610) );
  XOR U31812 ( .A(n31611), .B(n31612), .Z(n31602) );
  ANDN U31813 ( .A(n31613), .B(n25184), .Z(n31612) );
  XOR U31814 ( .A(n31614), .B(\modmult_1/zin[0][925] ), .Z(n25184) );
  IV U31815 ( .A(n31611), .Z(n31614) );
  XNOR U31816 ( .A(n31611), .B(n25183), .Z(n31613) );
  XOR U31817 ( .A(n31615), .B(n31616), .Z(n25183) );
  AND U31818 ( .A(\modmult_1/xin[1023] ), .B(n31617), .Z(n31616) );
  IV U31819 ( .A(n31615), .Z(n31617) );
  XOR U31820 ( .A(n31618), .B(g_input[926]), .Z(n31615) );
  NAND U31821 ( .A(n31619), .B(mul_pow), .Z(n31618) );
  XOR U31822 ( .A(g_input[926]), .B(creg[926]), .Z(n31619) );
  XOR U31823 ( .A(n31620), .B(n31621), .Z(n31611) );
  ANDN U31824 ( .A(n31622), .B(n25190), .Z(n31621) );
  XOR U31825 ( .A(n31623), .B(\modmult_1/zin[0][924] ), .Z(n25190) );
  IV U31826 ( .A(n31620), .Z(n31623) );
  XNOR U31827 ( .A(n31620), .B(n25189), .Z(n31622) );
  XOR U31828 ( .A(n31624), .B(n31625), .Z(n25189) );
  AND U31829 ( .A(\modmult_1/xin[1023] ), .B(n31626), .Z(n31625) );
  IV U31830 ( .A(n31624), .Z(n31626) );
  XOR U31831 ( .A(n31627), .B(g_input[925]), .Z(n31624) );
  NAND U31832 ( .A(n31628), .B(mul_pow), .Z(n31627) );
  XOR U31833 ( .A(g_input[925]), .B(creg[925]), .Z(n31628) );
  XOR U31834 ( .A(n31629), .B(n31630), .Z(n31620) );
  ANDN U31835 ( .A(n31631), .B(n25196), .Z(n31630) );
  XOR U31836 ( .A(n31632), .B(\modmult_1/zin[0][923] ), .Z(n25196) );
  IV U31837 ( .A(n31629), .Z(n31632) );
  XNOR U31838 ( .A(n31629), .B(n25195), .Z(n31631) );
  XOR U31839 ( .A(n31633), .B(n31634), .Z(n25195) );
  AND U31840 ( .A(\modmult_1/xin[1023] ), .B(n31635), .Z(n31634) );
  IV U31841 ( .A(n31633), .Z(n31635) );
  XOR U31842 ( .A(n31636), .B(g_input[924]), .Z(n31633) );
  NAND U31843 ( .A(n31637), .B(mul_pow), .Z(n31636) );
  XOR U31844 ( .A(g_input[924]), .B(creg[924]), .Z(n31637) );
  XOR U31845 ( .A(n31638), .B(n31639), .Z(n31629) );
  ANDN U31846 ( .A(n31640), .B(n25202), .Z(n31639) );
  XOR U31847 ( .A(n31641), .B(\modmult_1/zin[0][922] ), .Z(n25202) );
  IV U31848 ( .A(n31638), .Z(n31641) );
  XNOR U31849 ( .A(n31638), .B(n25201), .Z(n31640) );
  XOR U31850 ( .A(n31642), .B(n31643), .Z(n25201) );
  AND U31851 ( .A(\modmult_1/xin[1023] ), .B(n31644), .Z(n31643) );
  IV U31852 ( .A(n31642), .Z(n31644) );
  XOR U31853 ( .A(n31645), .B(g_input[923]), .Z(n31642) );
  NAND U31854 ( .A(n31646), .B(mul_pow), .Z(n31645) );
  XOR U31855 ( .A(g_input[923]), .B(creg[923]), .Z(n31646) );
  XOR U31856 ( .A(n31647), .B(n31648), .Z(n31638) );
  ANDN U31857 ( .A(n31649), .B(n25208), .Z(n31648) );
  XOR U31858 ( .A(n31650), .B(\modmult_1/zin[0][921] ), .Z(n25208) );
  IV U31859 ( .A(n31647), .Z(n31650) );
  XNOR U31860 ( .A(n31647), .B(n25207), .Z(n31649) );
  XOR U31861 ( .A(n31651), .B(n31652), .Z(n25207) );
  AND U31862 ( .A(\modmult_1/xin[1023] ), .B(n31653), .Z(n31652) );
  IV U31863 ( .A(n31651), .Z(n31653) );
  XOR U31864 ( .A(n31654), .B(g_input[922]), .Z(n31651) );
  NAND U31865 ( .A(n31655), .B(mul_pow), .Z(n31654) );
  XOR U31866 ( .A(g_input[922]), .B(creg[922]), .Z(n31655) );
  XOR U31867 ( .A(n31656), .B(n31657), .Z(n31647) );
  ANDN U31868 ( .A(n31658), .B(n25214), .Z(n31657) );
  XOR U31869 ( .A(n31659), .B(\modmult_1/zin[0][920] ), .Z(n25214) );
  IV U31870 ( .A(n31656), .Z(n31659) );
  XNOR U31871 ( .A(n31656), .B(n25213), .Z(n31658) );
  XOR U31872 ( .A(n31660), .B(n31661), .Z(n25213) );
  AND U31873 ( .A(\modmult_1/xin[1023] ), .B(n31662), .Z(n31661) );
  IV U31874 ( .A(n31660), .Z(n31662) );
  XOR U31875 ( .A(n31663), .B(g_input[921]), .Z(n31660) );
  NAND U31876 ( .A(n31664), .B(mul_pow), .Z(n31663) );
  XOR U31877 ( .A(g_input[921]), .B(creg[921]), .Z(n31664) );
  XOR U31878 ( .A(n31665), .B(n31666), .Z(n31656) );
  ANDN U31879 ( .A(n31667), .B(n25220), .Z(n31666) );
  XOR U31880 ( .A(n31668), .B(\modmult_1/zin[0][919] ), .Z(n25220) );
  IV U31881 ( .A(n31665), .Z(n31668) );
  XNOR U31882 ( .A(n31665), .B(n25219), .Z(n31667) );
  XOR U31883 ( .A(n31669), .B(n31670), .Z(n25219) );
  AND U31884 ( .A(\modmult_1/xin[1023] ), .B(n31671), .Z(n31670) );
  IV U31885 ( .A(n31669), .Z(n31671) );
  XOR U31886 ( .A(n31672), .B(g_input[920]), .Z(n31669) );
  NAND U31887 ( .A(n31673), .B(mul_pow), .Z(n31672) );
  XOR U31888 ( .A(g_input[920]), .B(creg[920]), .Z(n31673) );
  XOR U31889 ( .A(n31674), .B(n31675), .Z(n31665) );
  ANDN U31890 ( .A(n31676), .B(n25226), .Z(n31675) );
  XOR U31891 ( .A(n31677), .B(\modmult_1/zin[0][918] ), .Z(n25226) );
  IV U31892 ( .A(n31674), .Z(n31677) );
  XNOR U31893 ( .A(n31674), .B(n25225), .Z(n31676) );
  XOR U31894 ( .A(n31678), .B(n31679), .Z(n25225) );
  AND U31895 ( .A(\modmult_1/xin[1023] ), .B(n31680), .Z(n31679) );
  IV U31896 ( .A(n31678), .Z(n31680) );
  XOR U31897 ( .A(n31681), .B(g_input[919]), .Z(n31678) );
  NAND U31898 ( .A(n31682), .B(mul_pow), .Z(n31681) );
  XOR U31899 ( .A(g_input[919]), .B(creg[919]), .Z(n31682) );
  XOR U31900 ( .A(n31683), .B(n31684), .Z(n31674) );
  ANDN U31901 ( .A(n31685), .B(n25232), .Z(n31684) );
  XOR U31902 ( .A(n31686), .B(\modmult_1/zin[0][917] ), .Z(n25232) );
  IV U31903 ( .A(n31683), .Z(n31686) );
  XNOR U31904 ( .A(n31683), .B(n25231), .Z(n31685) );
  XOR U31905 ( .A(n31687), .B(n31688), .Z(n25231) );
  AND U31906 ( .A(\modmult_1/xin[1023] ), .B(n31689), .Z(n31688) );
  IV U31907 ( .A(n31687), .Z(n31689) );
  XOR U31908 ( .A(n31690), .B(g_input[918]), .Z(n31687) );
  NAND U31909 ( .A(n31691), .B(mul_pow), .Z(n31690) );
  XOR U31910 ( .A(g_input[918]), .B(creg[918]), .Z(n31691) );
  XOR U31911 ( .A(n31692), .B(n31693), .Z(n31683) );
  ANDN U31912 ( .A(n31694), .B(n25238), .Z(n31693) );
  XOR U31913 ( .A(n31695), .B(\modmult_1/zin[0][916] ), .Z(n25238) );
  IV U31914 ( .A(n31692), .Z(n31695) );
  XNOR U31915 ( .A(n31692), .B(n25237), .Z(n31694) );
  XOR U31916 ( .A(n31696), .B(n31697), .Z(n25237) );
  AND U31917 ( .A(\modmult_1/xin[1023] ), .B(n31698), .Z(n31697) );
  IV U31918 ( .A(n31696), .Z(n31698) );
  XOR U31919 ( .A(n31699), .B(g_input[917]), .Z(n31696) );
  NAND U31920 ( .A(n31700), .B(mul_pow), .Z(n31699) );
  XOR U31921 ( .A(g_input[917]), .B(creg[917]), .Z(n31700) );
  XOR U31922 ( .A(n31701), .B(n31702), .Z(n31692) );
  ANDN U31923 ( .A(n31703), .B(n25244), .Z(n31702) );
  XOR U31924 ( .A(n31704), .B(\modmult_1/zin[0][915] ), .Z(n25244) );
  IV U31925 ( .A(n31701), .Z(n31704) );
  XNOR U31926 ( .A(n31701), .B(n25243), .Z(n31703) );
  XOR U31927 ( .A(n31705), .B(n31706), .Z(n25243) );
  AND U31928 ( .A(\modmult_1/xin[1023] ), .B(n31707), .Z(n31706) );
  IV U31929 ( .A(n31705), .Z(n31707) );
  XOR U31930 ( .A(n31708), .B(g_input[916]), .Z(n31705) );
  NAND U31931 ( .A(n31709), .B(mul_pow), .Z(n31708) );
  XOR U31932 ( .A(g_input[916]), .B(creg[916]), .Z(n31709) );
  XOR U31933 ( .A(n31710), .B(n31711), .Z(n31701) );
  ANDN U31934 ( .A(n31712), .B(n25250), .Z(n31711) );
  XOR U31935 ( .A(n31713), .B(\modmult_1/zin[0][914] ), .Z(n25250) );
  IV U31936 ( .A(n31710), .Z(n31713) );
  XNOR U31937 ( .A(n31710), .B(n25249), .Z(n31712) );
  XOR U31938 ( .A(n31714), .B(n31715), .Z(n25249) );
  AND U31939 ( .A(\modmult_1/xin[1023] ), .B(n31716), .Z(n31715) );
  IV U31940 ( .A(n31714), .Z(n31716) );
  XOR U31941 ( .A(n31717), .B(g_input[915]), .Z(n31714) );
  NAND U31942 ( .A(n31718), .B(mul_pow), .Z(n31717) );
  XOR U31943 ( .A(g_input[915]), .B(creg[915]), .Z(n31718) );
  XOR U31944 ( .A(n31719), .B(n31720), .Z(n31710) );
  ANDN U31945 ( .A(n31721), .B(n25256), .Z(n31720) );
  XOR U31946 ( .A(n31722), .B(\modmult_1/zin[0][913] ), .Z(n25256) );
  IV U31947 ( .A(n31719), .Z(n31722) );
  XNOR U31948 ( .A(n31719), .B(n25255), .Z(n31721) );
  XOR U31949 ( .A(n31723), .B(n31724), .Z(n25255) );
  AND U31950 ( .A(\modmult_1/xin[1023] ), .B(n31725), .Z(n31724) );
  IV U31951 ( .A(n31723), .Z(n31725) );
  XOR U31952 ( .A(n31726), .B(g_input[914]), .Z(n31723) );
  NAND U31953 ( .A(n31727), .B(mul_pow), .Z(n31726) );
  XOR U31954 ( .A(g_input[914]), .B(creg[914]), .Z(n31727) );
  XOR U31955 ( .A(n31728), .B(n31729), .Z(n31719) );
  ANDN U31956 ( .A(n31730), .B(n25262), .Z(n31729) );
  XOR U31957 ( .A(n31731), .B(\modmult_1/zin[0][912] ), .Z(n25262) );
  IV U31958 ( .A(n31728), .Z(n31731) );
  XNOR U31959 ( .A(n31728), .B(n25261), .Z(n31730) );
  XOR U31960 ( .A(n31732), .B(n31733), .Z(n25261) );
  AND U31961 ( .A(\modmult_1/xin[1023] ), .B(n31734), .Z(n31733) );
  IV U31962 ( .A(n31732), .Z(n31734) );
  XOR U31963 ( .A(n31735), .B(g_input[913]), .Z(n31732) );
  NAND U31964 ( .A(n31736), .B(mul_pow), .Z(n31735) );
  XOR U31965 ( .A(g_input[913]), .B(creg[913]), .Z(n31736) );
  XOR U31966 ( .A(n31737), .B(n31738), .Z(n31728) );
  ANDN U31967 ( .A(n31739), .B(n25268), .Z(n31738) );
  XOR U31968 ( .A(n31740), .B(\modmult_1/zin[0][911] ), .Z(n25268) );
  IV U31969 ( .A(n31737), .Z(n31740) );
  XNOR U31970 ( .A(n31737), .B(n25267), .Z(n31739) );
  XOR U31971 ( .A(n31741), .B(n31742), .Z(n25267) );
  AND U31972 ( .A(\modmult_1/xin[1023] ), .B(n31743), .Z(n31742) );
  IV U31973 ( .A(n31741), .Z(n31743) );
  XOR U31974 ( .A(n31744), .B(g_input[912]), .Z(n31741) );
  NAND U31975 ( .A(n31745), .B(mul_pow), .Z(n31744) );
  XOR U31976 ( .A(g_input[912]), .B(creg[912]), .Z(n31745) );
  XOR U31977 ( .A(n31746), .B(n31747), .Z(n31737) );
  ANDN U31978 ( .A(n31748), .B(n25274), .Z(n31747) );
  XOR U31979 ( .A(n31749), .B(\modmult_1/zin[0][910] ), .Z(n25274) );
  IV U31980 ( .A(n31746), .Z(n31749) );
  XNOR U31981 ( .A(n31746), .B(n25273), .Z(n31748) );
  XOR U31982 ( .A(n31750), .B(n31751), .Z(n25273) );
  AND U31983 ( .A(\modmult_1/xin[1023] ), .B(n31752), .Z(n31751) );
  IV U31984 ( .A(n31750), .Z(n31752) );
  XOR U31985 ( .A(n31753), .B(g_input[911]), .Z(n31750) );
  NAND U31986 ( .A(n31754), .B(mul_pow), .Z(n31753) );
  XOR U31987 ( .A(g_input[911]), .B(creg[911]), .Z(n31754) );
  XOR U31988 ( .A(n31755), .B(n31756), .Z(n31746) );
  ANDN U31989 ( .A(n31757), .B(n25280), .Z(n31756) );
  XOR U31990 ( .A(n31758), .B(\modmult_1/zin[0][909] ), .Z(n25280) );
  IV U31991 ( .A(n31755), .Z(n31758) );
  XNOR U31992 ( .A(n31755), .B(n25279), .Z(n31757) );
  XOR U31993 ( .A(n31759), .B(n31760), .Z(n25279) );
  AND U31994 ( .A(\modmult_1/xin[1023] ), .B(n31761), .Z(n31760) );
  IV U31995 ( .A(n31759), .Z(n31761) );
  XOR U31996 ( .A(n31762), .B(g_input[910]), .Z(n31759) );
  NAND U31997 ( .A(n31763), .B(mul_pow), .Z(n31762) );
  XOR U31998 ( .A(g_input[910]), .B(creg[910]), .Z(n31763) );
  XOR U31999 ( .A(n31764), .B(n31765), .Z(n31755) );
  ANDN U32000 ( .A(n31766), .B(n25286), .Z(n31765) );
  XOR U32001 ( .A(n31767), .B(\modmult_1/zin[0][908] ), .Z(n25286) );
  IV U32002 ( .A(n31764), .Z(n31767) );
  XNOR U32003 ( .A(n31764), .B(n25285), .Z(n31766) );
  XOR U32004 ( .A(n31768), .B(n31769), .Z(n25285) );
  AND U32005 ( .A(\modmult_1/xin[1023] ), .B(n31770), .Z(n31769) );
  IV U32006 ( .A(n31768), .Z(n31770) );
  XOR U32007 ( .A(n31771), .B(g_input[909]), .Z(n31768) );
  NAND U32008 ( .A(n31772), .B(mul_pow), .Z(n31771) );
  XOR U32009 ( .A(g_input[909]), .B(creg[909]), .Z(n31772) );
  XOR U32010 ( .A(n31773), .B(n31774), .Z(n31764) );
  ANDN U32011 ( .A(n31775), .B(n25292), .Z(n31774) );
  XOR U32012 ( .A(n31776), .B(\modmult_1/zin[0][907] ), .Z(n25292) );
  IV U32013 ( .A(n31773), .Z(n31776) );
  XNOR U32014 ( .A(n31773), .B(n25291), .Z(n31775) );
  XOR U32015 ( .A(n31777), .B(n31778), .Z(n25291) );
  AND U32016 ( .A(\modmult_1/xin[1023] ), .B(n31779), .Z(n31778) );
  IV U32017 ( .A(n31777), .Z(n31779) );
  XOR U32018 ( .A(n31780), .B(g_input[908]), .Z(n31777) );
  NAND U32019 ( .A(n31781), .B(mul_pow), .Z(n31780) );
  XOR U32020 ( .A(g_input[908]), .B(creg[908]), .Z(n31781) );
  XOR U32021 ( .A(n31782), .B(n31783), .Z(n31773) );
  ANDN U32022 ( .A(n31784), .B(n25298), .Z(n31783) );
  XOR U32023 ( .A(n31785), .B(\modmult_1/zin[0][906] ), .Z(n25298) );
  IV U32024 ( .A(n31782), .Z(n31785) );
  XNOR U32025 ( .A(n31782), .B(n25297), .Z(n31784) );
  XOR U32026 ( .A(n31786), .B(n31787), .Z(n25297) );
  AND U32027 ( .A(\modmult_1/xin[1023] ), .B(n31788), .Z(n31787) );
  IV U32028 ( .A(n31786), .Z(n31788) );
  XOR U32029 ( .A(n31789), .B(g_input[907]), .Z(n31786) );
  NAND U32030 ( .A(n31790), .B(mul_pow), .Z(n31789) );
  XOR U32031 ( .A(g_input[907]), .B(creg[907]), .Z(n31790) );
  XOR U32032 ( .A(n31791), .B(n31792), .Z(n31782) );
  ANDN U32033 ( .A(n31793), .B(n25304), .Z(n31792) );
  XOR U32034 ( .A(n31794), .B(\modmult_1/zin[0][905] ), .Z(n25304) );
  IV U32035 ( .A(n31791), .Z(n31794) );
  XNOR U32036 ( .A(n31791), .B(n25303), .Z(n31793) );
  XOR U32037 ( .A(n31795), .B(n31796), .Z(n25303) );
  AND U32038 ( .A(\modmult_1/xin[1023] ), .B(n31797), .Z(n31796) );
  IV U32039 ( .A(n31795), .Z(n31797) );
  XOR U32040 ( .A(n31798), .B(g_input[906]), .Z(n31795) );
  NAND U32041 ( .A(n31799), .B(mul_pow), .Z(n31798) );
  XOR U32042 ( .A(g_input[906]), .B(creg[906]), .Z(n31799) );
  XOR U32043 ( .A(n31800), .B(n31801), .Z(n31791) );
  ANDN U32044 ( .A(n31802), .B(n25310), .Z(n31801) );
  XOR U32045 ( .A(n31803), .B(\modmult_1/zin[0][904] ), .Z(n25310) );
  IV U32046 ( .A(n31800), .Z(n31803) );
  XNOR U32047 ( .A(n31800), .B(n25309), .Z(n31802) );
  XOR U32048 ( .A(n31804), .B(n31805), .Z(n25309) );
  AND U32049 ( .A(\modmult_1/xin[1023] ), .B(n31806), .Z(n31805) );
  IV U32050 ( .A(n31804), .Z(n31806) );
  XOR U32051 ( .A(n31807), .B(g_input[905]), .Z(n31804) );
  NAND U32052 ( .A(n31808), .B(mul_pow), .Z(n31807) );
  XOR U32053 ( .A(g_input[905]), .B(creg[905]), .Z(n31808) );
  XOR U32054 ( .A(n31809), .B(n31810), .Z(n31800) );
  ANDN U32055 ( .A(n31811), .B(n25316), .Z(n31810) );
  XOR U32056 ( .A(n31812), .B(\modmult_1/zin[0][903] ), .Z(n25316) );
  IV U32057 ( .A(n31809), .Z(n31812) );
  XNOR U32058 ( .A(n31809), .B(n25315), .Z(n31811) );
  XOR U32059 ( .A(n31813), .B(n31814), .Z(n25315) );
  AND U32060 ( .A(\modmult_1/xin[1023] ), .B(n31815), .Z(n31814) );
  IV U32061 ( .A(n31813), .Z(n31815) );
  XOR U32062 ( .A(n31816), .B(g_input[904]), .Z(n31813) );
  NAND U32063 ( .A(n31817), .B(mul_pow), .Z(n31816) );
  XOR U32064 ( .A(g_input[904]), .B(creg[904]), .Z(n31817) );
  XOR U32065 ( .A(n31818), .B(n31819), .Z(n31809) );
  ANDN U32066 ( .A(n31820), .B(n25322), .Z(n31819) );
  XOR U32067 ( .A(n31821), .B(\modmult_1/zin[0][902] ), .Z(n25322) );
  IV U32068 ( .A(n31818), .Z(n31821) );
  XNOR U32069 ( .A(n31818), .B(n25321), .Z(n31820) );
  XOR U32070 ( .A(n31822), .B(n31823), .Z(n25321) );
  AND U32071 ( .A(\modmult_1/xin[1023] ), .B(n31824), .Z(n31823) );
  IV U32072 ( .A(n31822), .Z(n31824) );
  XOR U32073 ( .A(n31825), .B(g_input[903]), .Z(n31822) );
  NAND U32074 ( .A(n31826), .B(mul_pow), .Z(n31825) );
  XOR U32075 ( .A(g_input[903]), .B(creg[903]), .Z(n31826) );
  XOR U32076 ( .A(n31827), .B(n31828), .Z(n31818) );
  ANDN U32077 ( .A(n31829), .B(n25328), .Z(n31828) );
  XOR U32078 ( .A(n31830), .B(\modmult_1/zin[0][901] ), .Z(n25328) );
  IV U32079 ( .A(n31827), .Z(n31830) );
  XNOR U32080 ( .A(n31827), .B(n25327), .Z(n31829) );
  XOR U32081 ( .A(n31831), .B(n31832), .Z(n25327) );
  AND U32082 ( .A(\modmult_1/xin[1023] ), .B(n31833), .Z(n31832) );
  IV U32083 ( .A(n31831), .Z(n31833) );
  XOR U32084 ( .A(n31834), .B(g_input[902]), .Z(n31831) );
  NAND U32085 ( .A(n31835), .B(mul_pow), .Z(n31834) );
  XOR U32086 ( .A(g_input[902]), .B(creg[902]), .Z(n31835) );
  XOR U32087 ( .A(n31836), .B(n31837), .Z(n31827) );
  ANDN U32088 ( .A(n31838), .B(n25334), .Z(n31837) );
  XOR U32089 ( .A(n31839), .B(\modmult_1/zin[0][900] ), .Z(n25334) );
  IV U32090 ( .A(n31836), .Z(n31839) );
  XNOR U32091 ( .A(n31836), .B(n25333), .Z(n31838) );
  XOR U32092 ( .A(n31840), .B(n31841), .Z(n25333) );
  AND U32093 ( .A(\modmult_1/xin[1023] ), .B(n31842), .Z(n31841) );
  IV U32094 ( .A(n31840), .Z(n31842) );
  XOR U32095 ( .A(n31843), .B(g_input[901]), .Z(n31840) );
  NAND U32096 ( .A(n31844), .B(mul_pow), .Z(n31843) );
  XOR U32097 ( .A(g_input[901]), .B(creg[901]), .Z(n31844) );
  XOR U32098 ( .A(n31845), .B(n31846), .Z(n31836) );
  ANDN U32099 ( .A(n31847), .B(n25340), .Z(n31846) );
  XOR U32100 ( .A(n31848), .B(\modmult_1/zin[0][899] ), .Z(n25340) );
  IV U32101 ( .A(n31845), .Z(n31848) );
  XNOR U32102 ( .A(n31845), .B(n25339), .Z(n31847) );
  XOR U32103 ( .A(n31849), .B(n31850), .Z(n25339) );
  AND U32104 ( .A(\modmult_1/xin[1023] ), .B(n31851), .Z(n31850) );
  IV U32105 ( .A(n31849), .Z(n31851) );
  XOR U32106 ( .A(n31852), .B(g_input[900]), .Z(n31849) );
  NAND U32107 ( .A(n31853), .B(mul_pow), .Z(n31852) );
  XOR U32108 ( .A(g_input[900]), .B(creg[900]), .Z(n31853) );
  XOR U32109 ( .A(n31854), .B(n31855), .Z(n31845) );
  ANDN U32110 ( .A(n31856), .B(n25346), .Z(n31855) );
  XOR U32111 ( .A(n31857), .B(\modmult_1/zin[0][898] ), .Z(n25346) );
  IV U32112 ( .A(n31854), .Z(n31857) );
  XNOR U32113 ( .A(n31854), .B(n25345), .Z(n31856) );
  XOR U32114 ( .A(n31858), .B(n31859), .Z(n25345) );
  AND U32115 ( .A(\modmult_1/xin[1023] ), .B(n31860), .Z(n31859) );
  IV U32116 ( .A(n31858), .Z(n31860) );
  XOR U32117 ( .A(n31861), .B(g_input[899]), .Z(n31858) );
  NAND U32118 ( .A(n31862), .B(mul_pow), .Z(n31861) );
  XOR U32119 ( .A(g_input[899]), .B(creg[899]), .Z(n31862) );
  XOR U32120 ( .A(n31863), .B(n31864), .Z(n31854) );
  ANDN U32121 ( .A(n31865), .B(n25352), .Z(n31864) );
  XOR U32122 ( .A(n31866), .B(\modmult_1/zin[0][897] ), .Z(n25352) );
  IV U32123 ( .A(n31863), .Z(n31866) );
  XNOR U32124 ( .A(n31863), .B(n25351), .Z(n31865) );
  XOR U32125 ( .A(n31867), .B(n31868), .Z(n25351) );
  AND U32126 ( .A(\modmult_1/xin[1023] ), .B(n31869), .Z(n31868) );
  IV U32127 ( .A(n31867), .Z(n31869) );
  XOR U32128 ( .A(n31870), .B(g_input[898]), .Z(n31867) );
  NAND U32129 ( .A(n31871), .B(mul_pow), .Z(n31870) );
  XOR U32130 ( .A(g_input[898]), .B(creg[898]), .Z(n31871) );
  XOR U32131 ( .A(n31872), .B(n31873), .Z(n31863) );
  ANDN U32132 ( .A(n31874), .B(n25358), .Z(n31873) );
  XOR U32133 ( .A(n31875), .B(\modmult_1/zin[0][896] ), .Z(n25358) );
  IV U32134 ( .A(n31872), .Z(n31875) );
  XNOR U32135 ( .A(n31872), .B(n25357), .Z(n31874) );
  XOR U32136 ( .A(n31876), .B(n31877), .Z(n25357) );
  AND U32137 ( .A(\modmult_1/xin[1023] ), .B(n31878), .Z(n31877) );
  IV U32138 ( .A(n31876), .Z(n31878) );
  XOR U32139 ( .A(n31879), .B(g_input[897]), .Z(n31876) );
  NAND U32140 ( .A(n31880), .B(mul_pow), .Z(n31879) );
  XOR U32141 ( .A(g_input[897]), .B(creg[897]), .Z(n31880) );
  XOR U32142 ( .A(n31881), .B(n31882), .Z(n31872) );
  ANDN U32143 ( .A(n31883), .B(n25364), .Z(n31882) );
  XOR U32144 ( .A(n31884), .B(\modmult_1/zin[0][895] ), .Z(n25364) );
  IV U32145 ( .A(n31881), .Z(n31884) );
  XNOR U32146 ( .A(n31881), .B(n25363), .Z(n31883) );
  XOR U32147 ( .A(n31885), .B(n31886), .Z(n25363) );
  AND U32148 ( .A(\modmult_1/xin[1023] ), .B(n31887), .Z(n31886) );
  IV U32149 ( .A(n31885), .Z(n31887) );
  XOR U32150 ( .A(n31888), .B(g_input[896]), .Z(n31885) );
  NAND U32151 ( .A(n31889), .B(mul_pow), .Z(n31888) );
  XOR U32152 ( .A(g_input[896]), .B(creg[896]), .Z(n31889) );
  XOR U32153 ( .A(n31890), .B(n31891), .Z(n31881) );
  ANDN U32154 ( .A(n31892), .B(n25370), .Z(n31891) );
  XOR U32155 ( .A(n31893), .B(\modmult_1/zin[0][894] ), .Z(n25370) );
  IV U32156 ( .A(n31890), .Z(n31893) );
  XNOR U32157 ( .A(n31890), .B(n25369), .Z(n31892) );
  XOR U32158 ( .A(n31894), .B(n31895), .Z(n25369) );
  AND U32159 ( .A(\modmult_1/xin[1023] ), .B(n31896), .Z(n31895) );
  IV U32160 ( .A(n31894), .Z(n31896) );
  XOR U32161 ( .A(n31897), .B(g_input[895]), .Z(n31894) );
  NAND U32162 ( .A(n31898), .B(mul_pow), .Z(n31897) );
  XOR U32163 ( .A(g_input[895]), .B(creg[895]), .Z(n31898) );
  XOR U32164 ( .A(n31899), .B(n31900), .Z(n31890) );
  ANDN U32165 ( .A(n31901), .B(n25376), .Z(n31900) );
  XOR U32166 ( .A(n31902), .B(\modmult_1/zin[0][893] ), .Z(n25376) );
  IV U32167 ( .A(n31899), .Z(n31902) );
  XNOR U32168 ( .A(n31899), .B(n25375), .Z(n31901) );
  XOR U32169 ( .A(n31903), .B(n31904), .Z(n25375) );
  AND U32170 ( .A(\modmult_1/xin[1023] ), .B(n31905), .Z(n31904) );
  IV U32171 ( .A(n31903), .Z(n31905) );
  XOR U32172 ( .A(n31906), .B(g_input[894]), .Z(n31903) );
  NAND U32173 ( .A(n31907), .B(mul_pow), .Z(n31906) );
  XOR U32174 ( .A(g_input[894]), .B(creg[894]), .Z(n31907) );
  XOR U32175 ( .A(n31908), .B(n31909), .Z(n31899) );
  ANDN U32176 ( .A(n31910), .B(n25382), .Z(n31909) );
  XOR U32177 ( .A(n31911), .B(\modmult_1/zin[0][892] ), .Z(n25382) );
  IV U32178 ( .A(n31908), .Z(n31911) );
  XNOR U32179 ( .A(n31908), .B(n25381), .Z(n31910) );
  XOR U32180 ( .A(n31912), .B(n31913), .Z(n25381) );
  AND U32181 ( .A(\modmult_1/xin[1023] ), .B(n31914), .Z(n31913) );
  IV U32182 ( .A(n31912), .Z(n31914) );
  XOR U32183 ( .A(n31915), .B(g_input[893]), .Z(n31912) );
  NAND U32184 ( .A(n31916), .B(mul_pow), .Z(n31915) );
  XOR U32185 ( .A(g_input[893]), .B(creg[893]), .Z(n31916) );
  XOR U32186 ( .A(n31917), .B(n31918), .Z(n31908) );
  ANDN U32187 ( .A(n31919), .B(n25388), .Z(n31918) );
  XOR U32188 ( .A(n31920), .B(\modmult_1/zin[0][891] ), .Z(n25388) );
  IV U32189 ( .A(n31917), .Z(n31920) );
  XNOR U32190 ( .A(n31917), .B(n25387), .Z(n31919) );
  XOR U32191 ( .A(n31921), .B(n31922), .Z(n25387) );
  AND U32192 ( .A(\modmult_1/xin[1023] ), .B(n31923), .Z(n31922) );
  IV U32193 ( .A(n31921), .Z(n31923) );
  XOR U32194 ( .A(n31924), .B(g_input[892]), .Z(n31921) );
  NAND U32195 ( .A(n31925), .B(mul_pow), .Z(n31924) );
  XOR U32196 ( .A(g_input[892]), .B(creg[892]), .Z(n31925) );
  XOR U32197 ( .A(n31926), .B(n31927), .Z(n31917) );
  ANDN U32198 ( .A(n31928), .B(n25394), .Z(n31927) );
  XOR U32199 ( .A(n31929), .B(\modmult_1/zin[0][890] ), .Z(n25394) );
  IV U32200 ( .A(n31926), .Z(n31929) );
  XNOR U32201 ( .A(n31926), .B(n25393), .Z(n31928) );
  XOR U32202 ( .A(n31930), .B(n31931), .Z(n25393) );
  AND U32203 ( .A(\modmult_1/xin[1023] ), .B(n31932), .Z(n31931) );
  IV U32204 ( .A(n31930), .Z(n31932) );
  XOR U32205 ( .A(n31933), .B(g_input[891]), .Z(n31930) );
  NAND U32206 ( .A(n31934), .B(mul_pow), .Z(n31933) );
  XOR U32207 ( .A(g_input[891]), .B(creg[891]), .Z(n31934) );
  XOR U32208 ( .A(n31935), .B(n31936), .Z(n31926) );
  ANDN U32209 ( .A(n31937), .B(n25400), .Z(n31936) );
  XOR U32210 ( .A(n31938), .B(\modmult_1/zin[0][889] ), .Z(n25400) );
  IV U32211 ( .A(n31935), .Z(n31938) );
  XNOR U32212 ( .A(n31935), .B(n25399), .Z(n31937) );
  XOR U32213 ( .A(n31939), .B(n31940), .Z(n25399) );
  AND U32214 ( .A(\modmult_1/xin[1023] ), .B(n31941), .Z(n31940) );
  IV U32215 ( .A(n31939), .Z(n31941) );
  XOR U32216 ( .A(n31942), .B(g_input[890]), .Z(n31939) );
  NAND U32217 ( .A(n31943), .B(mul_pow), .Z(n31942) );
  XOR U32218 ( .A(g_input[890]), .B(creg[890]), .Z(n31943) );
  XOR U32219 ( .A(n31944), .B(n31945), .Z(n31935) );
  ANDN U32220 ( .A(n31946), .B(n25406), .Z(n31945) );
  XOR U32221 ( .A(n31947), .B(\modmult_1/zin[0][888] ), .Z(n25406) );
  IV U32222 ( .A(n31944), .Z(n31947) );
  XNOR U32223 ( .A(n31944), .B(n25405), .Z(n31946) );
  XOR U32224 ( .A(n31948), .B(n31949), .Z(n25405) );
  AND U32225 ( .A(\modmult_1/xin[1023] ), .B(n31950), .Z(n31949) );
  IV U32226 ( .A(n31948), .Z(n31950) );
  XOR U32227 ( .A(n31951), .B(g_input[889]), .Z(n31948) );
  NAND U32228 ( .A(n31952), .B(mul_pow), .Z(n31951) );
  XOR U32229 ( .A(g_input[889]), .B(creg[889]), .Z(n31952) );
  XOR U32230 ( .A(n31953), .B(n31954), .Z(n31944) );
  ANDN U32231 ( .A(n31955), .B(n25412), .Z(n31954) );
  XOR U32232 ( .A(n31956), .B(\modmult_1/zin[0][887] ), .Z(n25412) );
  IV U32233 ( .A(n31953), .Z(n31956) );
  XNOR U32234 ( .A(n31953), .B(n25411), .Z(n31955) );
  XOR U32235 ( .A(n31957), .B(n31958), .Z(n25411) );
  AND U32236 ( .A(\modmult_1/xin[1023] ), .B(n31959), .Z(n31958) );
  IV U32237 ( .A(n31957), .Z(n31959) );
  XOR U32238 ( .A(n31960), .B(g_input[888]), .Z(n31957) );
  NAND U32239 ( .A(n31961), .B(mul_pow), .Z(n31960) );
  XOR U32240 ( .A(g_input[888]), .B(creg[888]), .Z(n31961) );
  XOR U32241 ( .A(n31962), .B(n31963), .Z(n31953) );
  ANDN U32242 ( .A(n31964), .B(n25418), .Z(n31963) );
  XOR U32243 ( .A(n31965), .B(\modmult_1/zin[0][886] ), .Z(n25418) );
  IV U32244 ( .A(n31962), .Z(n31965) );
  XNOR U32245 ( .A(n31962), .B(n25417), .Z(n31964) );
  XOR U32246 ( .A(n31966), .B(n31967), .Z(n25417) );
  AND U32247 ( .A(\modmult_1/xin[1023] ), .B(n31968), .Z(n31967) );
  IV U32248 ( .A(n31966), .Z(n31968) );
  XOR U32249 ( .A(n31969), .B(g_input[887]), .Z(n31966) );
  NAND U32250 ( .A(n31970), .B(mul_pow), .Z(n31969) );
  XOR U32251 ( .A(g_input[887]), .B(creg[887]), .Z(n31970) );
  XOR U32252 ( .A(n31971), .B(n31972), .Z(n31962) );
  ANDN U32253 ( .A(n31973), .B(n25424), .Z(n31972) );
  XOR U32254 ( .A(n31974), .B(\modmult_1/zin[0][885] ), .Z(n25424) );
  IV U32255 ( .A(n31971), .Z(n31974) );
  XNOR U32256 ( .A(n31971), .B(n25423), .Z(n31973) );
  XOR U32257 ( .A(n31975), .B(n31976), .Z(n25423) );
  AND U32258 ( .A(\modmult_1/xin[1023] ), .B(n31977), .Z(n31976) );
  IV U32259 ( .A(n31975), .Z(n31977) );
  XOR U32260 ( .A(n31978), .B(g_input[886]), .Z(n31975) );
  NAND U32261 ( .A(n31979), .B(mul_pow), .Z(n31978) );
  XOR U32262 ( .A(g_input[886]), .B(creg[886]), .Z(n31979) );
  XOR U32263 ( .A(n31980), .B(n31981), .Z(n31971) );
  ANDN U32264 ( .A(n31982), .B(n25430), .Z(n31981) );
  XOR U32265 ( .A(n31983), .B(\modmult_1/zin[0][884] ), .Z(n25430) );
  IV U32266 ( .A(n31980), .Z(n31983) );
  XNOR U32267 ( .A(n31980), .B(n25429), .Z(n31982) );
  XOR U32268 ( .A(n31984), .B(n31985), .Z(n25429) );
  AND U32269 ( .A(\modmult_1/xin[1023] ), .B(n31986), .Z(n31985) );
  IV U32270 ( .A(n31984), .Z(n31986) );
  XOR U32271 ( .A(n31987), .B(g_input[885]), .Z(n31984) );
  NAND U32272 ( .A(n31988), .B(mul_pow), .Z(n31987) );
  XOR U32273 ( .A(g_input[885]), .B(creg[885]), .Z(n31988) );
  XOR U32274 ( .A(n31989), .B(n31990), .Z(n31980) );
  ANDN U32275 ( .A(n31991), .B(n25436), .Z(n31990) );
  XOR U32276 ( .A(n31992), .B(\modmult_1/zin[0][883] ), .Z(n25436) );
  IV U32277 ( .A(n31989), .Z(n31992) );
  XNOR U32278 ( .A(n31989), .B(n25435), .Z(n31991) );
  XOR U32279 ( .A(n31993), .B(n31994), .Z(n25435) );
  AND U32280 ( .A(\modmult_1/xin[1023] ), .B(n31995), .Z(n31994) );
  IV U32281 ( .A(n31993), .Z(n31995) );
  XOR U32282 ( .A(n31996), .B(g_input[884]), .Z(n31993) );
  NAND U32283 ( .A(n31997), .B(mul_pow), .Z(n31996) );
  XOR U32284 ( .A(g_input[884]), .B(creg[884]), .Z(n31997) );
  XOR U32285 ( .A(n31998), .B(n31999), .Z(n31989) );
  ANDN U32286 ( .A(n32000), .B(n25442), .Z(n31999) );
  XOR U32287 ( .A(n32001), .B(\modmult_1/zin[0][882] ), .Z(n25442) );
  IV U32288 ( .A(n31998), .Z(n32001) );
  XNOR U32289 ( .A(n31998), .B(n25441), .Z(n32000) );
  XOR U32290 ( .A(n32002), .B(n32003), .Z(n25441) );
  AND U32291 ( .A(\modmult_1/xin[1023] ), .B(n32004), .Z(n32003) );
  IV U32292 ( .A(n32002), .Z(n32004) );
  XOR U32293 ( .A(n32005), .B(g_input[883]), .Z(n32002) );
  NAND U32294 ( .A(n32006), .B(mul_pow), .Z(n32005) );
  XOR U32295 ( .A(g_input[883]), .B(creg[883]), .Z(n32006) );
  XOR U32296 ( .A(n32007), .B(n32008), .Z(n31998) );
  ANDN U32297 ( .A(n32009), .B(n25448), .Z(n32008) );
  XOR U32298 ( .A(n32010), .B(\modmult_1/zin[0][881] ), .Z(n25448) );
  IV U32299 ( .A(n32007), .Z(n32010) );
  XNOR U32300 ( .A(n32007), .B(n25447), .Z(n32009) );
  XOR U32301 ( .A(n32011), .B(n32012), .Z(n25447) );
  AND U32302 ( .A(\modmult_1/xin[1023] ), .B(n32013), .Z(n32012) );
  IV U32303 ( .A(n32011), .Z(n32013) );
  XOR U32304 ( .A(n32014), .B(g_input[882]), .Z(n32011) );
  NAND U32305 ( .A(n32015), .B(mul_pow), .Z(n32014) );
  XOR U32306 ( .A(g_input[882]), .B(creg[882]), .Z(n32015) );
  XOR U32307 ( .A(n32016), .B(n32017), .Z(n32007) );
  ANDN U32308 ( .A(n32018), .B(n25454), .Z(n32017) );
  XOR U32309 ( .A(n32019), .B(\modmult_1/zin[0][880] ), .Z(n25454) );
  IV U32310 ( .A(n32016), .Z(n32019) );
  XNOR U32311 ( .A(n32016), .B(n25453), .Z(n32018) );
  XOR U32312 ( .A(n32020), .B(n32021), .Z(n25453) );
  AND U32313 ( .A(\modmult_1/xin[1023] ), .B(n32022), .Z(n32021) );
  IV U32314 ( .A(n32020), .Z(n32022) );
  XOR U32315 ( .A(n32023), .B(g_input[881]), .Z(n32020) );
  NAND U32316 ( .A(n32024), .B(mul_pow), .Z(n32023) );
  XOR U32317 ( .A(g_input[881]), .B(creg[881]), .Z(n32024) );
  XOR U32318 ( .A(n32025), .B(n32026), .Z(n32016) );
  ANDN U32319 ( .A(n32027), .B(n25460), .Z(n32026) );
  XOR U32320 ( .A(n32028), .B(\modmult_1/zin[0][879] ), .Z(n25460) );
  IV U32321 ( .A(n32025), .Z(n32028) );
  XNOR U32322 ( .A(n32025), .B(n25459), .Z(n32027) );
  XOR U32323 ( .A(n32029), .B(n32030), .Z(n25459) );
  AND U32324 ( .A(\modmult_1/xin[1023] ), .B(n32031), .Z(n32030) );
  IV U32325 ( .A(n32029), .Z(n32031) );
  XOR U32326 ( .A(n32032), .B(g_input[880]), .Z(n32029) );
  NAND U32327 ( .A(n32033), .B(mul_pow), .Z(n32032) );
  XOR U32328 ( .A(g_input[880]), .B(creg[880]), .Z(n32033) );
  XOR U32329 ( .A(n32034), .B(n32035), .Z(n32025) );
  ANDN U32330 ( .A(n32036), .B(n25466), .Z(n32035) );
  XOR U32331 ( .A(n32037), .B(\modmult_1/zin[0][878] ), .Z(n25466) );
  IV U32332 ( .A(n32034), .Z(n32037) );
  XNOR U32333 ( .A(n32034), .B(n25465), .Z(n32036) );
  XOR U32334 ( .A(n32038), .B(n32039), .Z(n25465) );
  AND U32335 ( .A(\modmult_1/xin[1023] ), .B(n32040), .Z(n32039) );
  IV U32336 ( .A(n32038), .Z(n32040) );
  XOR U32337 ( .A(n32041), .B(g_input[879]), .Z(n32038) );
  NAND U32338 ( .A(n32042), .B(mul_pow), .Z(n32041) );
  XOR U32339 ( .A(g_input[879]), .B(creg[879]), .Z(n32042) );
  XOR U32340 ( .A(n32043), .B(n32044), .Z(n32034) );
  ANDN U32341 ( .A(n32045), .B(n25472), .Z(n32044) );
  XOR U32342 ( .A(n32046), .B(\modmult_1/zin[0][877] ), .Z(n25472) );
  IV U32343 ( .A(n32043), .Z(n32046) );
  XNOR U32344 ( .A(n32043), .B(n25471), .Z(n32045) );
  XOR U32345 ( .A(n32047), .B(n32048), .Z(n25471) );
  AND U32346 ( .A(\modmult_1/xin[1023] ), .B(n32049), .Z(n32048) );
  IV U32347 ( .A(n32047), .Z(n32049) );
  XOR U32348 ( .A(n32050), .B(g_input[878]), .Z(n32047) );
  NAND U32349 ( .A(n32051), .B(mul_pow), .Z(n32050) );
  XOR U32350 ( .A(g_input[878]), .B(creg[878]), .Z(n32051) );
  XOR U32351 ( .A(n32052), .B(n32053), .Z(n32043) );
  ANDN U32352 ( .A(n32054), .B(n25478), .Z(n32053) );
  XOR U32353 ( .A(n32055), .B(\modmult_1/zin[0][876] ), .Z(n25478) );
  IV U32354 ( .A(n32052), .Z(n32055) );
  XNOR U32355 ( .A(n32052), .B(n25477), .Z(n32054) );
  XOR U32356 ( .A(n32056), .B(n32057), .Z(n25477) );
  AND U32357 ( .A(\modmult_1/xin[1023] ), .B(n32058), .Z(n32057) );
  IV U32358 ( .A(n32056), .Z(n32058) );
  XOR U32359 ( .A(n32059), .B(g_input[877]), .Z(n32056) );
  NAND U32360 ( .A(n32060), .B(mul_pow), .Z(n32059) );
  XOR U32361 ( .A(g_input[877]), .B(creg[877]), .Z(n32060) );
  XOR U32362 ( .A(n32061), .B(n32062), .Z(n32052) );
  ANDN U32363 ( .A(n32063), .B(n25484), .Z(n32062) );
  XOR U32364 ( .A(n32064), .B(\modmult_1/zin[0][875] ), .Z(n25484) );
  IV U32365 ( .A(n32061), .Z(n32064) );
  XNOR U32366 ( .A(n32061), .B(n25483), .Z(n32063) );
  XOR U32367 ( .A(n32065), .B(n32066), .Z(n25483) );
  AND U32368 ( .A(\modmult_1/xin[1023] ), .B(n32067), .Z(n32066) );
  IV U32369 ( .A(n32065), .Z(n32067) );
  XOR U32370 ( .A(n32068), .B(g_input[876]), .Z(n32065) );
  NAND U32371 ( .A(n32069), .B(mul_pow), .Z(n32068) );
  XOR U32372 ( .A(g_input[876]), .B(creg[876]), .Z(n32069) );
  XOR U32373 ( .A(n32070), .B(n32071), .Z(n32061) );
  ANDN U32374 ( .A(n32072), .B(n25490), .Z(n32071) );
  XOR U32375 ( .A(n32073), .B(\modmult_1/zin[0][874] ), .Z(n25490) );
  IV U32376 ( .A(n32070), .Z(n32073) );
  XNOR U32377 ( .A(n32070), .B(n25489), .Z(n32072) );
  XOR U32378 ( .A(n32074), .B(n32075), .Z(n25489) );
  AND U32379 ( .A(\modmult_1/xin[1023] ), .B(n32076), .Z(n32075) );
  IV U32380 ( .A(n32074), .Z(n32076) );
  XOR U32381 ( .A(n32077), .B(g_input[875]), .Z(n32074) );
  NAND U32382 ( .A(n32078), .B(mul_pow), .Z(n32077) );
  XOR U32383 ( .A(g_input[875]), .B(creg[875]), .Z(n32078) );
  XOR U32384 ( .A(n32079), .B(n32080), .Z(n32070) );
  ANDN U32385 ( .A(n32081), .B(n25496), .Z(n32080) );
  XOR U32386 ( .A(n32082), .B(\modmult_1/zin[0][873] ), .Z(n25496) );
  IV U32387 ( .A(n32079), .Z(n32082) );
  XNOR U32388 ( .A(n32079), .B(n25495), .Z(n32081) );
  XOR U32389 ( .A(n32083), .B(n32084), .Z(n25495) );
  AND U32390 ( .A(\modmult_1/xin[1023] ), .B(n32085), .Z(n32084) );
  IV U32391 ( .A(n32083), .Z(n32085) );
  XOR U32392 ( .A(n32086), .B(g_input[874]), .Z(n32083) );
  NAND U32393 ( .A(n32087), .B(mul_pow), .Z(n32086) );
  XOR U32394 ( .A(g_input[874]), .B(creg[874]), .Z(n32087) );
  XOR U32395 ( .A(n32088), .B(n32089), .Z(n32079) );
  ANDN U32396 ( .A(n32090), .B(n25502), .Z(n32089) );
  XOR U32397 ( .A(n32091), .B(\modmult_1/zin[0][872] ), .Z(n25502) );
  IV U32398 ( .A(n32088), .Z(n32091) );
  XNOR U32399 ( .A(n32088), .B(n25501), .Z(n32090) );
  XOR U32400 ( .A(n32092), .B(n32093), .Z(n25501) );
  AND U32401 ( .A(\modmult_1/xin[1023] ), .B(n32094), .Z(n32093) );
  IV U32402 ( .A(n32092), .Z(n32094) );
  XOR U32403 ( .A(n32095), .B(g_input[873]), .Z(n32092) );
  NAND U32404 ( .A(n32096), .B(mul_pow), .Z(n32095) );
  XOR U32405 ( .A(g_input[873]), .B(creg[873]), .Z(n32096) );
  XOR U32406 ( .A(n32097), .B(n32098), .Z(n32088) );
  ANDN U32407 ( .A(n32099), .B(n25508), .Z(n32098) );
  XOR U32408 ( .A(n32100), .B(\modmult_1/zin[0][871] ), .Z(n25508) );
  IV U32409 ( .A(n32097), .Z(n32100) );
  XNOR U32410 ( .A(n32097), .B(n25507), .Z(n32099) );
  XOR U32411 ( .A(n32101), .B(n32102), .Z(n25507) );
  AND U32412 ( .A(\modmult_1/xin[1023] ), .B(n32103), .Z(n32102) );
  IV U32413 ( .A(n32101), .Z(n32103) );
  XOR U32414 ( .A(n32104), .B(g_input[872]), .Z(n32101) );
  NAND U32415 ( .A(n32105), .B(mul_pow), .Z(n32104) );
  XOR U32416 ( .A(g_input[872]), .B(creg[872]), .Z(n32105) );
  XOR U32417 ( .A(n32106), .B(n32107), .Z(n32097) );
  ANDN U32418 ( .A(n32108), .B(n25514), .Z(n32107) );
  XOR U32419 ( .A(n32109), .B(\modmult_1/zin[0][870] ), .Z(n25514) );
  IV U32420 ( .A(n32106), .Z(n32109) );
  XNOR U32421 ( .A(n32106), .B(n25513), .Z(n32108) );
  XOR U32422 ( .A(n32110), .B(n32111), .Z(n25513) );
  AND U32423 ( .A(\modmult_1/xin[1023] ), .B(n32112), .Z(n32111) );
  IV U32424 ( .A(n32110), .Z(n32112) );
  XOR U32425 ( .A(n32113), .B(g_input[871]), .Z(n32110) );
  NAND U32426 ( .A(n32114), .B(mul_pow), .Z(n32113) );
  XOR U32427 ( .A(g_input[871]), .B(creg[871]), .Z(n32114) );
  XOR U32428 ( .A(n32115), .B(n32116), .Z(n32106) );
  ANDN U32429 ( .A(n32117), .B(n25520), .Z(n32116) );
  XOR U32430 ( .A(n32118), .B(\modmult_1/zin[0][869] ), .Z(n25520) );
  IV U32431 ( .A(n32115), .Z(n32118) );
  XNOR U32432 ( .A(n32115), .B(n25519), .Z(n32117) );
  XOR U32433 ( .A(n32119), .B(n32120), .Z(n25519) );
  AND U32434 ( .A(\modmult_1/xin[1023] ), .B(n32121), .Z(n32120) );
  IV U32435 ( .A(n32119), .Z(n32121) );
  XOR U32436 ( .A(n32122), .B(g_input[870]), .Z(n32119) );
  NAND U32437 ( .A(n32123), .B(mul_pow), .Z(n32122) );
  XOR U32438 ( .A(g_input[870]), .B(creg[870]), .Z(n32123) );
  XOR U32439 ( .A(n32124), .B(n32125), .Z(n32115) );
  ANDN U32440 ( .A(n32126), .B(n25526), .Z(n32125) );
  XOR U32441 ( .A(n32127), .B(\modmult_1/zin[0][868] ), .Z(n25526) );
  IV U32442 ( .A(n32124), .Z(n32127) );
  XNOR U32443 ( .A(n32124), .B(n25525), .Z(n32126) );
  XOR U32444 ( .A(n32128), .B(n32129), .Z(n25525) );
  AND U32445 ( .A(\modmult_1/xin[1023] ), .B(n32130), .Z(n32129) );
  IV U32446 ( .A(n32128), .Z(n32130) );
  XOR U32447 ( .A(n32131), .B(g_input[869]), .Z(n32128) );
  NAND U32448 ( .A(n32132), .B(mul_pow), .Z(n32131) );
  XOR U32449 ( .A(g_input[869]), .B(creg[869]), .Z(n32132) );
  XOR U32450 ( .A(n32133), .B(n32134), .Z(n32124) );
  ANDN U32451 ( .A(n32135), .B(n25532), .Z(n32134) );
  XOR U32452 ( .A(n32136), .B(\modmult_1/zin[0][867] ), .Z(n25532) );
  IV U32453 ( .A(n32133), .Z(n32136) );
  XNOR U32454 ( .A(n32133), .B(n25531), .Z(n32135) );
  XOR U32455 ( .A(n32137), .B(n32138), .Z(n25531) );
  AND U32456 ( .A(\modmult_1/xin[1023] ), .B(n32139), .Z(n32138) );
  IV U32457 ( .A(n32137), .Z(n32139) );
  XOR U32458 ( .A(n32140), .B(g_input[868]), .Z(n32137) );
  NAND U32459 ( .A(n32141), .B(mul_pow), .Z(n32140) );
  XOR U32460 ( .A(g_input[868]), .B(creg[868]), .Z(n32141) );
  XOR U32461 ( .A(n32142), .B(n32143), .Z(n32133) );
  ANDN U32462 ( .A(n32144), .B(n25538), .Z(n32143) );
  XOR U32463 ( .A(n32145), .B(\modmult_1/zin[0][866] ), .Z(n25538) );
  IV U32464 ( .A(n32142), .Z(n32145) );
  XNOR U32465 ( .A(n32142), .B(n25537), .Z(n32144) );
  XOR U32466 ( .A(n32146), .B(n32147), .Z(n25537) );
  AND U32467 ( .A(\modmult_1/xin[1023] ), .B(n32148), .Z(n32147) );
  IV U32468 ( .A(n32146), .Z(n32148) );
  XOR U32469 ( .A(n32149), .B(g_input[867]), .Z(n32146) );
  NAND U32470 ( .A(n32150), .B(mul_pow), .Z(n32149) );
  XOR U32471 ( .A(g_input[867]), .B(creg[867]), .Z(n32150) );
  XOR U32472 ( .A(n32151), .B(n32152), .Z(n32142) );
  ANDN U32473 ( .A(n32153), .B(n25544), .Z(n32152) );
  XOR U32474 ( .A(n32154), .B(\modmult_1/zin[0][865] ), .Z(n25544) );
  IV U32475 ( .A(n32151), .Z(n32154) );
  XNOR U32476 ( .A(n32151), .B(n25543), .Z(n32153) );
  XOR U32477 ( .A(n32155), .B(n32156), .Z(n25543) );
  AND U32478 ( .A(\modmult_1/xin[1023] ), .B(n32157), .Z(n32156) );
  IV U32479 ( .A(n32155), .Z(n32157) );
  XOR U32480 ( .A(n32158), .B(g_input[866]), .Z(n32155) );
  NAND U32481 ( .A(n32159), .B(mul_pow), .Z(n32158) );
  XOR U32482 ( .A(g_input[866]), .B(creg[866]), .Z(n32159) );
  XOR U32483 ( .A(n32160), .B(n32161), .Z(n32151) );
  ANDN U32484 ( .A(n32162), .B(n25550), .Z(n32161) );
  XOR U32485 ( .A(n32163), .B(\modmult_1/zin[0][864] ), .Z(n25550) );
  IV U32486 ( .A(n32160), .Z(n32163) );
  XNOR U32487 ( .A(n32160), .B(n25549), .Z(n32162) );
  XOR U32488 ( .A(n32164), .B(n32165), .Z(n25549) );
  AND U32489 ( .A(\modmult_1/xin[1023] ), .B(n32166), .Z(n32165) );
  IV U32490 ( .A(n32164), .Z(n32166) );
  XOR U32491 ( .A(n32167), .B(g_input[865]), .Z(n32164) );
  NAND U32492 ( .A(n32168), .B(mul_pow), .Z(n32167) );
  XOR U32493 ( .A(g_input[865]), .B(creg[865]), .Z(n32168) );
  XOR U32494 ( .A(n32169), .B(n32170), .Z(n32160) );
  ANDN U32495 ( .A(n32171), .B(n25556), .Z(n32170) );
  XOR U32496 ( .A(n32172), .B(\modmult_1/zin[0][863] ), .Z(n25556) );
  IV U32497 ( .A(n32169), .Z(n32172) );
  XNOR U32498 ( .A(n32169), .B(n25555), .Z(n32171) );
  XOR U32499 ( .A(n32173), .B(n32174), .Z(n25555) );
  AND U32500 ( .A(\modmult_1/xin[1023] ), .B(n32175), .Z(n32174) );
  IV U32501 ( .A(n32173), .Z(n32175) );
  XOR U32502 ( .A(n32176), .B(g_input[864]), .Z(n32173) );
  NAND U32503 ( .A(n32177), .B(mul_pow), .Z(n32176) );
  XOR U32504 ( .A(g_input[864]), .B(creg[864]), .Z(n32177) );
  XOR U32505 ( .A(n32178), .B(n32179), .Z(n32169) );
  ANDN U32506 ( .A(n32180), .B(n25562), .Z(n32179) );
  XOR U32507 ( .A(n32181), .B(\modmult_1/zin[0][862] ), .Z(n25562) );
  IV U32508 ( .A(n32178), .Z(n32181) );
  XNOR U32509 ( .A(n32178), .B(n25561), .Z(n32180) );
  XOR U32510 ( .A(n32182), .B(n32183), .Z(n25561) );
  AND U32511 ( .A(\modmult_1/xin[1023] ), .B(n32184), .Z(n32183) );
  IV U32512 ( .A(n32182), .Z(n32184) );
  XOR U32513 ( .A(n32185), .B(g_input[863]), .Z(n32182) );
  NAND U32514 ( .A(n32186), .B(mul_pow), .Z(n32185) );
  XOR U32515 ( .A(g_input[863]), .B(creg[863]), .Z(n32186) );
  XOR U32516 ( .A(n32187), .B(n32188), .Z(n32178) );
  ANDN U32517 ( .A(n32189), .B(n25568), .Z(n32188) );
  XOR U32518 ( .A(n32190), .B(\modmult_1/zin[0][861] ), .Z(n25568) );
  IV U32519 ( .A(n32187), .Z(n32190) );
  XNOR U32520 ( .A(n32187), .B(n25567), .Z(n32189) );
  XOR U32521 ( .A(n32191), .B(n32192), .Z(n25567) );
  AND U32522 ( .A(\modmult_1/xin[1023] ), .B(n32193), .Z(n32192) );
  IV U32523 ( .A(n32191), .Z(n32193) );
  XOR U32524 ( .A(n32194), .B(g_input[862]), .Z(n32191) );
  NAND U32525 ( .A(n32195), .B(mul_pow), .Z(n32194) );
  XOR U32526 ( .A(g_input[862]), .B(creg[862]), .Z(n32195) );
  XOR U32527 ( .A(n32196), .B(n32197), .Z(n32187) );
  ANDN U32528 ( .A(n32198), .B(n25574), .Z(n32197) );
  XOR U32529 ( .A(n32199), .B(\modmult_1/zin[0][860] ), .Z(n25574) );
  IV U32530 ( .A(n32196), .Z(n32199) );
  XNOR U32531 ( .A(n32196), .B(n25573), .Z(n32198) );
  XOR U32532 ( .A(n32200), .B(n32201), .Z(n25573) );
  AND U32533 ( .A(\modmult_1/xin[1023] ), .B(n32202), .Z(n32201) );
  IV U32534 ( .A(n32200), .Z(n32202) );
  XOR U32535 ( .A(n32203), .B(g_input[861]), .Z(n32200) );
  NAND U32536 ( .A(n32204), .B(mul_pow), .Z(n32203) );
  XOR U32537 ( .A(g_input[861]), .B(creg[861]), .Z(n32204) );
  XOR U32538 ( .A(n32205), .B(n32206), .Z(n32196) );
  ANDN U32539 ( .A(n32207), .B(n25580), .Z(n32206) );
  XOR U32540 ( .A(n32208), .B(\modmult_1/zin[0][859] ), .Z(n25580) );
  IV U32541 ( .A(n32205), .Z(n32208) );
  XNOR U32542 ( .A(n32205), .B(n25579), .Z(n32207) );
  XOR U32543 ( .A(n32209), .B(n32210), .Z(n25579) );
  AND U32544 ( .A(\modmult_1/xin[1023] ), .B(n32211), .Z(n32210) );
  IV U32545 ( .A(n32209), .Z(n32211) );
  XOR U32546 ( .A(n32212), .B(g_input[860]), .Z(n32209) );
  NAND U32547 ( .A(n32213), .B(mul_pow), .Z(n32212) );
  XOR U32548 ( .A(g_input[860]), .B(creg[860]), .Z(n32213) );
  XOR U32549 ( .A(n32214), .B(n32215), .Z(n32205) );
  ANDN U32550 ( .A(n32216), .B(n25586), .Z(n32215) );
  XOR U32551 ( .A(n32217), .B(\modmult_1/zin[0][858] ), .Z(n25586) );
  IV U32552 ( .A(n32214), .Z(n32217) );
  XNOR U32553 ( .A(n32214), .B(n25585), .Z(n32216) );
  XOR U32554 ( .A(n32218), .B(n32219), .Z(n25585) );
  AND U32555 ( .A(\modmult_1/xin[1023] ), .B(n32220), .Z(n32219) );
  IV U32556 ( .A(n32218), .Z(n32220) );
  XOR U32557 ( .A(n32221), .B(g_input[859]), .Z(n32218) );
  NAND U32558 ( .A(n32222), .B(mul_pow), .Z(n32221) );
  XOR U32559 ( .A(g_input[859]), .B(creg[859]), .Z(n32222) );
  XOR U32560 ( .A(n32223), .B(n32224), .Z(n32214) );
  ANDN U32561 ( .A(n32225), .B(n25592), .Z(n32224) );
  XOR U32562 ( .A(n32226), .B(\modmult_1/zin[0][857] ), .Z(n25592) );
  IV U32563 ( .A(n32223), .Z(n32226) );
  XNOR U32564 ( .A(n32223), .B(n25591), .Z(n32225) );
  XOR U32565 ( .A(n32227), .B(n32228), .Z(n25591) );
  AND U32566 ( .A(\modmult_1/xin[1023] ), .B(n32229), .Z(n32228) );
  IV U32567 ( .A(n32227), .Z(n32229) );
  XOR U32568 ( .A(n32230), .B(g_input[858]), .Z(n32227) );
  NAND U32569 ( .A(n32231), .B(mul_pow), .Z(n32230) );
  XOR U32570 ( .A(g_input[858]), .B(creg[858]), .Z(n32231) );
  XOR U32571 ( .A(n32232), .B(n32233), .Z(n32223) );
  ANDN U32572 ( .A(n32234), .B(n25598), .Z(n32233) );
  XOR U32573 ( .A(n32235), .B(\modmult_1/zin[0][856] ), .Z(n25598) );
  IV U32574 ( .A(n32232), .Z(n32235) );
  XNOR U32575 ( .A(n32232), .B(n25597), .Z(n32234) );
  XOR U32576 ( .A(n32236), .B(n32237), .Z(n25597) );
  AND U32577 ( .A(\modmult_1/xin[1023] ), .B(n32238), .Z(n32237) );
  IV U32578 ( .A(n32236), .Z(n32238) );
  XOR U32579 ( .A(n32239), .B(g_input[857]), .Z(n32236) );
  NAND U32580 ( .A(n32240), .B(mul_pow), .Z(n32239) );
  XOR U32581 ( .A(g_input[857]), .B(creg[857]), .Z(n32240) );
  XOR U32582 ( .A(n32241), .B(n32242), .Z(n32232) );
  ANDN U32583 ( .A(n32243), .B(n25604), .Z(n32242) );
  XOR U32584 ( .A(n32244), .B(\modmult_1/zin[0][855] ), .Z(n25604) );
  IV U32585 ( .A(n32241), .Z(n32244) );
  XNOR U32586 ( .A(n32241), .B(n25603), .Z(n32243) );
  XOR U32587 ( .A(n32245), .B(n32246), .Z(n25603) );
  AND U32588 ( .A(\modmult_1/xin[1023] ), .B(n32247), .Z(n32246) );
  IV U32589 ( .A(n32245), .Z(n32247) );
  XOR U32590 ( .A(n32248), .B(g_input[856]), .Z(n32245) );
  NAND U32591 ( .A(n32249), .B(mul_pow), .Z(n32248) );
  XOR U32592 ( .A(g_input[856]), .B(creg[856]), .Z(n32249) );
  XOR U32593 ( .A(n32250), .B(n32251), .Z(n32241) );
  ANDN U32594 ( .A(n32252), .B(n25610), .Z(n32251) );
  XOR U32595 ( .A(n32253), .B(\modmult_1/zin[0][854] ), .Z(n25610) );
  IV U32596 ( .A(n32250), .Z(n32253) );
  XNOR U32597 ( .A(n32250), .B(n25609), .Z(n32252) );
  XOR U32598 ( .A(n32254), .B(n32255), .Z(n25609) );
  AND U32599 ( .A(\modmult_1/xin[1023] ), .B(n32256), .Z(n32255) );
  IV U32600 ( .A(n32254), .Z(n32256) );
  XOR U32601 ( .A(n32257), .B(g_input[855]), .Z(n32254) );
  NAND U32602 ( .A(n32258), .B(mul_pow), .Z(n32257) );
  XOR U32603 ( .A(g_input[855]), .B(creg[855]), .Z(n32258) );
  XOR U32604 ( .A(n32259), .B(n32260), .Z(n32250) );
  ANDN U32605 ( .A(n32261), .B(n25616), .Z(n32260) );
  XOR U32606 ( .A(n32262), .B(\modmult_1/zin[0][853] ), .Z(n25616) );
  IV U32607 ( .A(n32259), .Z(n32262) );
  XNOR U32608 ( .A(n32259), .B(n25615), .Z(n32261) );
  XOR U32609 ( .A(n32263), .B(n32264), .Z(n25615) );
  AND U32610 ( .A(\modmult_1/xin[1023] ), .B(n32265), .Z(n32264) );
  IV U32611 ( .A(n32263), .Z(n32265) );
  XOR U32612 ( .A(n32266), .B(g_input[854]), .Z(n32263) );
  NAND U32613 ( .A(n32267), .B(mul_pow), .Z(n32266) );
  XOR U32614 ( .A(g_input[854]), .B(creg[854]), .Z(n32267) );
  XOR U32615 ( .A(n32268), .B(n32269), .Z(n32259) );
  ANDN U32616 ( .A(n32270), .B(n25622), .Z(n32269) );
  XOR U32617 ( .A(n32271), .B(\modmult_1/zin[0][852] ), .Z(n25622) );
  IV U32618 ( .A(n32268), .Z(n32271) );
  XNOR U32619 ( .A(n32268), .B(n25621), .Z(n32270) );
  XOR U32620 ( .A(n32272), .B(n32273), .Z(n25621) );
  AND U32621 ( .A(\modmult_1/xin[1023] ), .B(n32274), .Z(n32273) );
  IV U32622 ( .A(n32272), .Z(n32274) );
  XOR U32623 ( .A(n32275), .B(g_input[853]), .Z(n32272) );
  NAND U32624 ( .A(n32276), .B(mul_pow), .Z(n32275) );
  XOR U32625 ( .A(g_input[853]), .B(creg[853]), .Z(n32276) );
  XOR U32626 ( .A(n32277), .B(n32278), .Z(n32268) );
  ANDN U32627 ( .A(n32279), .B(n25628), .Z(n32278) );
  XOR U32628 ( .A(n32280), .B(\modmult_1/zin[0][851] ), .Z(n25628) );
  IV U32629 ( .A(n32277), .Z(n32280) );
  XNOR U32630 ( .A(n32277), .B(n25627), .Z(n32279) );
  XOR U32631 ( .A(n32281), .B(n32282), .Z(n25627) );
  AND U32632 ( .A(\modmult_1/xin[1023] ), .B(n32283), .Z(n32282) );
  IV U32633 ( .A(n32281), .Z(n32283) );
  XOR U32634 ( .A(n32284), .B(g_input[852]), .Z(n32281) );
  NAND U32635 ( .A(n32285), .B(mul_pow), .Z(n32284) );
  XOR U32636 ( .A(g_input[852]), .B(creg[852]), .Z(n32285) );
  XOR U32637 ( .A(n32286), .B(n32287), .Z(n32277) );
  ANDN U32638 ( .A(n32288), .B(n25634), .Z(n32287) );
  XOR U32639 ( .A(n32289), .B(\modmult_1/zin[0][850] ), .Z(n25634) );
  IV U32640 ( .A(n32286), .Z(n32289) );
  XNOR U32641 ( .A(n32286), .B(n25633), .Z(n32288) );
  XOR U32642 ( .A(n32290), .B(n32291), .Z(n25633) );
  AND U32643 ( .A(\modmult_1/xin[1023] ), .B(n32292), .Z(n32291) );
  IV U32644 ( .A(n32290), .Z(n32292) );
  XOR U32645 ( .A(n32293), .B(g_input[851]), .Z(n32290) );
  NAND U32646 ( .A(n32294), .B(mul_pow), .Z(n32293) );
  XOR U32647 ( .A(g_input[851]), .B(creg[851]), .Z(n32294) );
  XOR U32648 ( .A(n32295), .B(n32296), .Z(n32286) );
  ANDN U32649 ( .A(n32297), .B(n25640), .Z(n32296) );
  XOR U32650 ( .A(n32298), .B(\modmult_1/zin[0][849] ), .Z(n25640) );
  IV U32651 ( .A(n32295), .Z(n32298) );
  XNOR U32652 ( .A(n32295), .B(n25639), .Z(n32297) );
  XOR U32653 ( .A(n32299), .B(n32300), .Z(n25639) );
  AND U32654 ( .A(\modmult_1/xin[1023] ), .B(n32301), .Z(n32300) );
  IV U32655 ( .A(n32299), .Z(n32301) );
  XOR U32656 ( .A(n32302), .B(g_input[850]), .Z(n32299) );
  NAND U32657 ( .A(n32303), .B(mul_pow), .Z(n32302) );
  XOR U32658 ( .A(g_input[850]), .B(creg[850]), .Z(n32303) );
  XOR U32659 ( .A(n32304), .B(n32305), .Z(n32295) );
  ANDN U32660 ( .A(n32306), .B(n25646), .Z(n32305) );
  XOR U32661 ( .A(n32307), .B(\modmult_1/zin[0][848] ), .Z(n25646) );
  IV U32662 ( .A(n32304), .Z(n32307) );
  XNOR U32663 ( .A(n32304), .B(n25645), .Z(n32306) );
  XOR U32664 ( .A(n32308), .B(n32309), .Z(n25645) );
  AND U32665 ( .A(\modmult_1/xin[1023] ), .B(n32310), .Z(n32309) );
  IV U32666 ( .A(n32308), .Z(n32310) );
  XOR U32667 ( .A(n32311), .B(g_input[849]), .Z(n32308) );
  NAND U32668 ( .A(n32312), .B(mul_pow), .Z(n32311) );
  XOR U32669 ( .A(g_input[849]), .B(creg[849]), .Z(n32312) );
  XOR U32670 ( .A(n32313), .B(n32314), .Z(n32304) );
  ANDN U32671 ( .A(n32315), .B(n25652), .Z(n32314) );
  XOR U32672 ( .A(n32316), .B(\modmult_1/zin[0][847] ), .Z(n25652) );
  IV U32673 ( .A(n32313), .Z(n32316) );
  XNOR U32674 ( .A(n32313), .B(n25651), .Z(n32315) );
  XOR U32675 ( .A(n32317), .B(n32318), .Z(n25651) );
  AND U32676 ( .A(\modmult_1/xin[1023] ), .B(n32319), .Z(n32318) );
  IV U32677 ( .A(n32317), .Z(n32319) );
  XOR U32678 ( .A(n32320), .B(g_input[848]), .Z(n32317) );
  NAND U32679 ( .A(n32321), .B(mul_pow), .Z(n32320) );
  XOR U32680 ( .A(g_input[848]), .B(creg[848]), .Z(n32321) );
  XOR U32681 ( .A(n32322), .B(n32323), .Z(n32313) );
  ANDN U32682 ( .A(n32324), .B(n25658), .Z(n32323) );
  XOR U32683 ( .A(n32325), .B(\modmult_1/zin[0][846] ), .Z(n25658) );
  IV U32684 ( .A(n32322), .Z(n32325) );
  XNOR U32685 ( .A(n32322), .B(n25657), .Z(n32324) );
  XOR U32686 ( .A(n32326), .B(n32327), .Z(n25657) );
  AND U32687 ( .A(\modmult_1/xin[1023] ), .B(n32328), .Z(n32327) );
  IV U32688 ( .A(n32326), .Z(n32328) );
  XOR U32689 ( .A(n32329), .B(g_input[847]), .Z(n32326) );
  NAND U32690 ( .A(n32330), .B(mul_pow), .Z(n32329) );
  XOR U32691 ( .A(g_input[847]), .B(creg[847]), .Z(n32330) );
  XOR U32692 ( .A(n32331), .B(n32332), .Z(n32322) );
  ANDN U32693 ( .A(n32333), .B(n25664), .Z(n32332) );
  XOR U32694 ( .A(n32334), .B(\modmult_1/zin[0][845] ), .Z(n25664) );
  IV U32695 ( .A(n32331), .Z(n32334) );
  XNOR U32696 ( .A(n32331), .B(n25663), .Z(n32333) );
  XOR U32697 ( .A(n32335), .B(n32336), .Z(n25663) );
  AND U32698 ( .A(\modmult_1/xin[1023] ), .B(n32337), .Z(n32336) );
  IV U32699 ( .A(n32335), .Z(n32337) );
  XOR U32700 ( .A(n32338), .B(g_input[846]), .Z(n32335) );
  NAND U32701 ( .A(n32339), .B(mul_pow), .Z(n32338) );
  XOR U32702 ( .A(g_input[846]), .B(creg[846]), .Z(n32339) );
  XOR U32703 ( .A(n32340), .B(n32341), .Z(n32331) );
  ANDN U32704 ( .A(n32342), .B(n25670), .Z(n32341) );
  XOR U32705 ( .A(n32343), .B(\modmult_1/zin[0][844] ), .Z(n25670) );
  IV U32706 ( .A(n32340), .Z(n32343) );
  XNOR U32707 ( .A(n32340), .B(n25669), .Z(n32342) );
  XOR U32708 ( .A(n32344), .B(n32345), .Z(n25669) );
  AND U32709 ( .A(\modmult_1/xin[1023] ), .B(n32346), .Z(n32345) );
  IV U32710 ( .A(n32344), .Z(n32346) );
  XOR U32711 ( .A(n32347), .B(g_input[845]), .Z(n32344) );
  NAND U32712 ( .A(n32348), .B(mul_pow), .Z(n32347) );
  XOR U32713 ( .A(g_input[845]), .B(creg[845]), .Z(n32348) );
  XOR U32714 ( .A(n32349), .B(n32350), .Z(n32340) );
  ANDN U32715 ( .A(n32351), .B(n25676), .Z(n32350) );
  XOR U32716 ( .A(n32352), .B(\modmult_1/zin[0][843] ), .Z(n25676) );
  IV U32717 ( .A(n32349), .Z(n32352) );
  XNOR U32718 ( .A(n32349), .B(n25675), .Z(n32351) );
  XOR U32719 ( .A(n32353), .B(n32354), .Z(n25675) );
  AND U32720 ( .A(\modmult_1/xin[1023] ), .B(n32355), .Z(n32354) );
  IV U32721 ( .A(n32353), .Z(n32355) );
  XOR U32722 ( .A(n32356), .B(g_input[844]), .Z(n32353) );
  NAND U32723 ( .A(n32357), .B(mul_pow), .Z(n32356) );
  XOR U32724 ( .A(g_input[844]), .B(creg[844]), .Z(n32357) );
  XOR U32725 ( .A(n32358), .B(n32359), .Z(n32349) );
  ANDN U32726 ( .A(n32360), .B(n25682), .Z(n32359) );
  XOR U32727 ( .A(n32361), .B(\modmult_1/zin[0][842] ), .Z(n25682) );
  IV U32728 ( .A(n32358), .Z(n32361) );
  XNOR U32729 ( .A(n32358), .B(n25681), .Z(n32360) );
  XOR U32730 ( .A(n32362), .B(n32363), .Z(n25681) );
  AND U32731 ( .A(\modmult_1/xin[1023] ), .B(n32364), .Z(n32363) );
  IV U32732 ( .A(n32362), .Z(n32364) );
  XOR U32733 ( .A(n32365), .B(g_input[843]), .Z(n32362) );
  NAND U32734 ( .A(n32366), .B(mul_pow), .Z(n32365) );
  XOR U32735 ( .A(g_input[843]), .B(creg[843]), .Z(n32366) );
  XOR U32736 ( .A(n32367), .B(n32368), .Z(n32358) );
  ANDN U32737 ( .A(n32369), .B(n25688), .Z(n32368) );
  XOR U32738 ( .A(n32370), .B(\modmult_1/zin[0][841] ), .Z(n25688) );
  IV U32739 ( .A(n32367), .Z(n32370) );
  XNOR U32740 ( .A(n32367), .B(n25687), .Z(n32369) );
  XOR U32741 ( .A(n32371), .B(n32372), .Z(n25687) );
  AND U32742 ( .A(\modmult_1/xin[1023] ), .B(n32373), .Z(n32372) );
  IV U32743 ( .A(n32371), .Z(n32373) );
  XOR U32744 ( .A(n32374), .B(g_input[842]), .Z(n32371) );
  NAND U32745 ( .A(n32375), .B(mul_pow), .Z(n32374) );
  XOR U32746 ( .A(g_input[842]), .B(creg[842]), .Z(n32375) );
  XOR U32747 ( .A(n32376), .B(n32377), .Z(n32367) );
  ANDN U32748 ( .A(n32378), .B(n25694), .Z(n32377) );
  XOR U32749 ( .A(n32379), .B(\modmult_1/zin[0][840] ), .Z(n25694) );
  IV U32750 ( .A(n32376), .Z(n32379) );
  XNOR U32751 ( .A(n32376), .B(n25693), .Z(n32378) );
  XOR U32752 ( .A(n32380), .B(n32381), .Z(n25693) );
  AND U32753 ( .A(\modmult_1/xin[1023] ), .B(n32382), .Z(n32381) );
  IV U32754 ( .A(n32380), .Z(n32382) );
  XOR U32755 ( .A(n32383), .B(g_input[841]), .Z(n32380) );
  NAND U32756 ( .A(n32384), .B(mul_pow), .Z(n32383) );
  XOR U32757 ( .A(g_input[841]), .B(creg[841]), .Z(n32384) );
  XOR U32758 ( .A(n32385), .B(n32386), .Z(n32376) );
  ANDN U32759 ( .A(n32387), .B(n25700), .Z(n32386) );
  XOR U32760 ( .A(n32388), .B(\modmult_1/zin[0][839] ), .Z(n25700) );
  IV U32761 ( .A(n32385), .Z(n32388) );
  XNOR U32762 ( .A(n32385), .B(n25699), .Z(n32387) );
  XOR U32763 ( .A(n32389), .B(n32390), .Z(n25699) );
  AND U32764 ( .A(\modmult_1/xin[1023] ), .B(n32391), .Z(n32390) );
  IV U32765 ( .A(n32389), .Z(n32391) );
  XOR U32766 ( .A(n32392), .B(g_input[840]), .Z(n32389) );
  NAND U32767 ( .A(n32393), .B(mul_pow), .Z(n32392) );
  XOR U32768 ( .A(g_input[840]), .B(creg[840]), .Z(n32393) );
  XOR U32769 ( .A(n32394), .B(n32395), .Z(n32385) );
  ANDN U32770 ( .A(n32396), .B(n25706), .Z(n32395) );
  XOR U32771 ( .A(n32397), .B(\modmult_1/zin[0][838] ), .Z(n25706) );
  IV U32772 ( .A(n32394), .Z(n32397) );
  XNOR U32773 ( .A(n32394), .B(n25705), .Z(n32396) );
  XOR U32774 ( .A(n32398), .B(n32399), .Z(n25705) );
  AND U32775 ( .A(\modmult_1/xin[1023] ), .B(n32400), .Z(n32399) );
  IV U32776 ( .A(n32398), .Z(n32400) );
  XOR U32777 ( .A(n32401), .B(g_input[839]), .Z(n32398) );
  NAND U32778 ( .A(n32402), .B(mul_pow), .Z(n32401) );
  XOR U32779 ( .A(g_input[839]), .B(creg[839]), .Z(n32402) );
  XOR U32780 ( .A(n32403), .B(n32404), .Z(n32394) );
  ANDN U32781 ( .A(n32405), .B(n25712), .Z(n32404) );
  XOR U32782 ( .A(n32406), .B(\modmult_1/zin[0][837] ), .Z(n25712) );
  IV U32783 ( .A(n32403), .Z(n32406) );
  XNOR U32784 ( .A(n32403), .B(n25711), .Z(n32405) );
  XOR U32785 ( .A(n32407), .B(n32408), .Z(n25711) );
  AND U32786 ( .A(\modmult_1/xin[1023] ), .B(n32409), .Z(n32408) );
  IV U32787 ( .A(n32407), .Z(n32409) );
  XOR U32788 ( .A(n32410), .B(g_input[838]), .Z(n32407) );
  NAND U32789 ( .A(n32411), .B(mul_pow), .Z(n32410) );
  XOR U32790 ( .A(g_input[838]), .B(creg[838]), .Z(n32411) );
  XOR U32791 ( .A(n32412), .B(n32413), .Z(n32403) );
  ANDN U32792 ( .A(n32414), .B(n25718), .Z(n32413) );
  XOR U32793 ( .A(n32415), .B(\modmult_1/zin[0][836] ), .Z(n25718) );
  IV U32794 ( .A(n32412), .Z(n32415) );
  XNOR U32795 ( .A(n32412), .B(n25717), .Z(n32414) );
  XOR U32796 ( .A(n32416), .B(n32417), .Z(n25717) );
  AND U32797 ( .A(\modmult_1/xin[1023] ), .B(n32418), .Z(n32417) );
  IV U32798 ( .A(n32416), .Z(n32418) );
  XOR U32799 ( .A(n32419), .B(g_input[837]), .Z(n32416) );
  NAND U32800 ( .A(n32420), .B(mul_pow), .Z(n32419) );
  XOR U32801 ( .A(g_input[837]), .B(creg[837]), .Z(n32420) );
  XOR U32802 ( .A(n32421), .B(n32422), .Z(n32412) );
  ANDN U32803 ( .A(n32423), .B(n25724), .Z(n32422) );
  XOR U32804 ( .A(n32424), .B(\modmult_1/zin[0][835] ), .Z(n25724) );
  IV U32805 ( .A(n32421), .Z(n32424) );
  XNOR U32806 ( .A(n32421), .B(n25723), .Z(n32423) );
  XOR U32807 ( .A(n32425), .B(n32426), .Z(n25723) );
  AND U32808 ( .A(\modmult_1/xin[1023] ), .B(n32427), .Z(n32426) );
  IV U32809 ( .A(n32425), .Z(n32427) );
  XOR U32810 ( .A(n32428), .B(g_input[836]), .Z(n32425) );
  NAND U32811 ( .A(n32429), .B(mul_pow), .Z(n32428) );
  XOR U32812 ( .A(g_input[836]), .B(creg[836]), .Z(n32429) );
  XOR U32813 ( .A(n32430), .B(n32431), .Z(n32421) );
  ANDN U32814 ( .A(n32432), .B(n25730), .Z(n32431) );
  XOR U32815 ( .A(n32433), .B(\modmult_1/zin[0][834] ), .Z(n25730) );
  IV U32816 ( .A(n32430), .Z(n32433) );
  XNOR U32817 ( .A(n32430), .B(n25729), .Z(n32432) );
  XOR U32818 ( .A(n32434), .B(n32435), .Z(n25729) );
  AND U32819 ( .A(\modmult_1/xin[1023] ), .B(n32436), .Z(n32435) );
  IV U32820 ( .A(n32434), .Z(n32436) );
  XOR U32821 ( .A(n32437), .B(g_input[835]), .Z(n32434) );
  NAND U32822 ( .A(n32438), .B(mul_pow), .Z(n32437) );
  XOR U32823 ( .A(g_input[835]), .B(creg[835]), .Z(n32438) );
  XOR U32824 ( .A(n32439), .B(n32440), .Z(n32430) );
  ANDN U32825 ( .A(n32441), .B(n25736), .Z(n32440) );
  XOR U32826 ( .A(n32442), .B(\modmult_1/zin[0][833] ), .Z(n25736) );
  IV U32827 ( .A(n32439), .Z(n32442) );
  XNOR U32828 ( .A(n32439), .B(n25735), .Z(n32441) );
  XOR U32829 ( .A(n32443), .B(n32444), .Z(n25735) );
  AND U32830 ( .A(\modmult_1/xin[1023] ), .B(n32445), .Z(n32444) );
  IV U32831 ( .A(n32443), .Z(n32445) );
  XOR U32832 ( .A(n32446), .B(g_input[834]), .Z(n32443) );
  NAND U32833 ( .A(n32447), .B(mul_pow), .Z(n32446) );
  XOR U32834 ( .A(g_input[834]), .B(creg[834]), .Z(n32447) );
  XOR U32835 ( .A(n32448), .B(n32449), .Z(n32439) );
  ANDN U32836 ( .A(n32450), .B(n25742), .Z(n32449) );
  XOR U32837 ( .A(n32451), .B(\modmult_1/zin[0][832] ), .Z(n25742) );
  IV U32838 ( .A(n32448), .Z(n32451) );
  XNOR U32839 ( .A(n32448), .B(n25741), .Z(n32450) );
  XOR U32840 ( .A(n32452), .B(n32453), .Z(n25741) );
  AND U32841 ( .A(\modmult_1/xin[1023] ), .B(n32454), .Z(n32453) );
  IV U32842 ( .A(n32452), .Z(n32454) );
  XOR U32843 ( .A(n32455), .B(g_input[833]), .Z(n32452) );
  NAND U32844 ( .A(n32456), .B(mul_pow), .Z(n32455) );
  XOR U32845 ( .A(g_input[833]), .B(creg[833]), .Z(n32456) );
  XOR U32846 ( .A(n32457), .B(n32458), .Z(n32448) );
  ANDN U32847 ( .A(n32459), .B(n25748), .Z(n32458) );
  XOR U32848 ( .A(n32460), .B(\modmult_1/zin[0][831] ), .Z(n25748) );
  IV U32849 ( .A(n32457), .Z(n32460) );
  XNOR U32850 ( .A(n32457), .B(n25747), .Z(n32459) );
  XOR U32851 ( .A(n32461), .B(n32462), .Z(n25747) );
  AND U32852 ( .A(\modmult_1/xin[1023] ), .B(n32463), .Z(n32462) );
  IV U32853 ( .A(n32461), .Z(n32463) );
  XOR U32854 ( .A(n32464), .B(g_input[832]), .Z(n32461) );
  NAND U32855 ( .A(n32465), .B(mul_pow), .Z(n32464) );
  XOR U32856 ( .A(g_input[832]), .B(creg[832]), .Z(n32465) );
  XOR U32857 ( .A(n32466), .B(n32467), .Z(n32457) );
  ANDN U32858 ( .A(n32468), .B(n25754), .Z(n32467) );
  XOR U32859 ( .A(n32469), .B(\modmult_1/zin[0][830] ), .Z(n25754) );
  IV U32860 ( .A(n32466), .Z(n32469) );
  XNOR U32861 ( .A(n32466), .B(n25753), .Z(n32468) );
  XOR U32862 ( .A(n32470), .B(n32471), .Z(n25753) );
  AND U32863 ( .A(\modmult_1/xin[1023] ), .B(n32472), .Z(n32471) );
  IV U32864 ( .A(n32470), .Z(n32472) );
  XOR U32865 ( .A(n32473), .B(g_input[831]), .Z(n32470) );
  NAND U32866 ( .A(n32474), .B(mul_pow), .Z(n32473) );
  XOR U32867 ( .A(g_input[831]), .B(creg[831]), .Z(n32474) );
  XOR U32868 ( .A(n32475), .B(n32476), .Z(n32466) );
  ANDN U32869 ( .A(n32477), .B(n25760), .Z(n32476) );
  XOR U32870 ( .A(n32478), .B(\modmult_1/zin[0][829] ), .Z(n25760) );
  IV U32871 ( .A(n32475), .Z(n32478) );
  XNOR U32872 ( .A(n32475), .B(n25759), .Z(n32477) );
  XOR U32873 ( .A(n32479), .B(n32480), .Z(n25759) );
  AND U32874 ( .A(\modmult_1/xin[1023] ), .B(n32481), .Z(n32480) );
  IV U32875 ( .A(n32479), .Z(n32481) );
  XOR U32876 ( .A(n32482), .B(g_input[830]), .Z(n32479) );
  NAND U32877 ( .A(n32483), .B(mul_pow), .Z(n32482) );
  XOR U32878 ( .A(g_input[830]), .B(creg[830]), .Z(n32483) );
  XOR U32879 ( .A(n32484), .B(n32485), .Z(n32475) );
  ANDN U32880 ( .A(n32486), .B(n25766), .Z(n32485) );
  XOR U32881 ( .A(n32487), .B(\modmult_1/zin[0][828] ), .Z(n25766) );
  IV U32882 ( .A(n32484), .Z(n32487) );
  XNOR U32883 ( .A(n32484), .B(n25765), .Z(n32486) );
  XOR U32884 ( .A(n32488), .B(n32489), .Z(n25765) );
  AND U32885 ( .A(\modmult_1/xin[1023] ), .B(n32490), .Z(n32489) );
  IV U32886 ( .A(n32488), .Z(n32490) );
  XOR U32887 ( .A(n32491), .B(g_input[829]), .Z(n32488) );
  NAND U32888 ( .A(n32492), .B(mul_pow), .Z(n32491) );
  XOR U32889 ( .A(g_input[829]), .B(creg[829]), .Z(n32492) );
  XOR U32890 ( .A(n32493), .B(n32494), .Z(n32484) );
  ANDN U32891 ( .A(n32495), .B(n25772), .Z(n32494) );
  XOR U32892 ( .A(n32496), .B(\modmult_1/zin[0][827] ), .Z(n25772) );
  IV U32893 ( .A(n32493), .Z(n32496) );
  XNOR U32894 ( .A(n32493), .B(n25771), .Z(n32495) );
  XOR U32895 ( .A(n32497), .B(n32498), .Z(n25771) );
  AND U32896 ( .A(\modmult_1/xin[1023] ), .B(n32499), .Z(n32498) );
  IV U32897 ( .A(n32497), .Z(n32499) );
  XOR U32898 ( .A(n32500), .B(g_input[828]), .Z(n32497) );
  NAND U32899 ( .A(n32501), .B(mul_pow), .Z(n32500) );
  XOR U32900 ( .A(g_input[828]), .B(creg[828]), .Z(n32501) );
  XOR U32901 ( .A(n32502), .B(n32503), .Z(n32493) );
  ANDN U32902 ( .A(n32504), .B(n25778), .Z(n32503) );
  XOR U32903 ( .A(n32505), .B(\modmult_1/zin[0][826] ), .Z(n25778) );
  IV U32904 ( .A(n32502), .Z(n32505) );
  XNOR U32905 ( .A(n32502), .B(n25777), .Z(n32504) );
  XOR U32906 ( .A(n32506), .B(n32507), .Z(n25777) );
  AND U32907 ( .A(\modmult_1/xin[1023] ), .B(n32508), .Z(n32507) );
  IV U32908 ( .A(n32506), .Z(n32508) );
  XOR U32909 ( .A(n32509), .B(g_input[827]), .Z(n32506) );
  NAND U32910 ( .A(n32510), .B(mul_pow), .Z(n32509) );
  XOR U32911 ( .A(g_input[827]), .B(creg[827]), .Z(n32510) );
  XOR U32912 ( .A(n32511), .B(n32512), .Z(n32502) );
  ANDN U32913 ( .A(n32513), .B(n25784), .Z(n32512) );
  XOR U32914 ( .A(n32514), .B(\modmult_1/zin[0][825] ), .Z(n25784) );
  IV U32915 ( .A(n32511), .Z(n32514) );
  XNOR U32916 ( .A(n32511), .B(n25783), .Z(n32513) );
  XOR U32917 ( .A(n32515), .B(n32516), .Z(n25783) );
  AND U32918 ( .A(\modmult_1/xin[1023] ), .B(n32517), .Z(n32516) );
  IV U32919 ( .A(n32515), .Z(n32517) );
  XOR U32920 ( .A(n32518), .B(g_input[826]), .Z(n32515) );
  NAND U32921 ( .A(n32519), .B(mul_pow), .Z(n32518) );
  XOR U32922 ( .A(g_input[826]), .B(creg[826]), .Z(n32519) );
  XOR U32923 ( .A(n32520), .B(n32521), .Z(n32511) );
  ANDN U32924 ( .A(n32522), .B(n25790), .Z(n32521) );
  XOR U32925 ( .A(n32523), .B(\modmult_1/zin[0][824] ), .Z(n25790) );
  IV U32926 ( .A(n32520), .Z(n32523) );
  XNOR U32927 ( .A(n32520), .B(n25789), .Z(n32522) );
  XOR U32928 ( .A(n32524), .B(n32525), .Z(n25789) );
  AND U32929 ( .A(\modmult_1/xin[1023] ), .B(n32526), .Z(n32525) );
  IV U32930 ( .A(n32524), .Z(n32526) );
  XOR U32931 ( .A(n32527), .B(g_input[825]), .Z(n32524) );
  NAND U32932 ( .A(n32528), .B(mul_pow), .Z(n32527) );
  XOR U32933 ( .A(g_input[825]), .B(creg[825]), .Z(n32528) );
  XOR U32934 ( .A(n32529), .B(n32530), .Z(n32520) );
  ANDN U32935 ( .A(n32531), .B(n25796), .Z(n32530) );
  XOR U32936 ( .A(n32532), .B(\modmult_1/zin[0][823] ), .Z(n25796) );
  IV U32937 ( .A(n32529), .Z(n32532) );
  XNOR U32938 ( .A(n32529), .B(n25795), .Z(n32531) );
  XOR U32939 ( .A(n32533), .B(n32534), .Z(n25795) );
  AND U32940 ( .A(\modmult_1/xin[1023] ), .B(n32535), .Z(n32534) );
  IV U32941 ( .A(n32533), .Z(n32535) );
  XOR U32942 ( .A(n32536), .B(g_input[824]), .Z(n32533) );
  NAND U32943 ( .A(n32537), .B(mul_pow), .Z(n32536) );
  XOR U32944 ( .A(g_input[824]), .B(creg[824]), .Z(n32537) );
  XOR U32945 ( .A(n32538), .B(n32539), .Z(n32529) );
  ANDN U32946 ( .A(n32540), .B(n25802), .Z(n32539) );
  XOR U32947 ( .A(n32541), .B(\modmult_1/zin[0][822] ), .Z(n25802) );
  IV U32948 ( .A(n32538), .Z(n32541) );
  XNOR U32949 ( .A(n32538), .B(n25801), .Z(n32540) );
  XOR U32950 ( .A(n32542), .B(n32543), .Z(n25801) );
  AND U32951 ( .A(\modmult_1/xin[1023] ), .B(n32544), .Z(n32543) );
  IV U32952 ( .A(n32542), .Z(n32544) );
  XOR U32953 ( .A(n32545), .B(g_input[823]), .Z(n32542) );
  NAND U32954 ( .A(n32546), .B(mul_pow), .Z(n32545) );
  XOR U32955 ( .A(g_input[823]), .B(creg[823]), .Z(n32546) );
  XOR U32956 ( .A(n32547), .B(n32548), .Z(n32538) );
  ANDN U32957 ( .A(n32549), .B(n25808), .Z(n32548) );
  XOR U32958 ( .A(n32550), .B(\modmult_1/zin[0][821] ), .Z(n25808) );
  IV U32959 ( .A(n32547), .Z(n32550) );
  XNOR U32960 ( .A(n32547), .B(n25807), .Z(n32549) );
  XOR U32961 ( .A(n32551), .B(n32552), .Z(n25807) );
  AND U32962 ( .A(\modmult_1/xin[1023] ), .B(n32553), .Z(n32552) );
  IV U32963 ( .A(n32551), .Z(n32553) );
  XOR U32964 ( .A(n32554), .B(g_input[822]), .Z(n32551) );
  NAND U32965 ( .A(n32555), .B(mul_pow), .Z(n32554) );
  XOR U32966 ( .A(g_input[822]), .B(creg[822]), .Z(n32555) );
  XOR U32967 ( .A(n32556), .B(n32557), .Z(n32547) );
  ANDN U32968 ( .A(n32558), .B(n25814), .Z(n32557) );
  XOR U32969 ( .A(n32559), .B(\modmult_1/zin[0][820] ), .Z(n25814) );
  IV U32970 ( .A(n32556), .Z(n32559) );
  XNOR U32971 ( .A(n32556), .B(n25813), .Z(n32558) );
  XOR U32972 ( .A(n32560), .B(n32561), .Z(n25813) );
  AND U32973 ( .A(\modmult_1/xin[1023] ), .B(n32562), .Z(n32561) );
  IV U32974 ( .A(n32560), .Z(n32562) );
  XOR U32975 ( .A(n32563), .B(g_input[821]), .Z(n32560) );
  NAND U32976 ( .A(n32564), .B(mul_pow), .Z(n32563) );
  XOR U32977 ( .A(g_input[821]), .B(creg[821]), .Z(n32564) );
  XOR U32978 ( .A(n32565), .B(n32566), .Z(n32556) );
  ANDN U32979 ( .A(n32567), .B(n25820), .Z(n32566) );
  XOR U32980 ( .A(n32568), .B(\modmult_1/zin[0][819] ), .Z(n25820) );
  IV U32981 ( .A(n32565), .Z(n32568) );
  XNOR U32982 ( .A(n32565), .B(n25819), .Z(n32567) );
  XOR U32983 ( .A(n32569), .B(n32570), .Z(n25819) );
  AND U32984 ( .A(\modmult_1/xin[1023] ), .B(n32571), .Z(n32570) );
  IV U32985 ( .A(n32569), .Z(n32571) );
  XOR U32986 ( .A(n32572), .B(g_input[820]), .Z(n32569) );
  NAND U32987 ( .A(n32573), .B(mul_pow), .Z(n32572) );
  XOR U32988 ( .A(g_input[820]), .B(creg[820]), .Z(n32573) );
  XOR U32989 ( .A(n32574), .B(n32575), .Z(n32565) );
  ANDN U32990 ( .A(n32576), .B(n25826), .Z(n32575) );
  XOR U32991 ( .A(n32577), .B(\modmult_1/zin[0][818] ), .Z(n25826) );
  IV U32992 ( .A(n32574), .Z(n32577) );
  XNOR U32993 ( .A(n32574), .B(n25825), .Z(n32576) );
  XOR U32994 ( .A(n32578), .B(n32579), .Z(n25825) );
  AND U32995 ( .A(\modmult_1/xin[1023] ), .B(n32580), .Z(n32579) );
  IV U32996 ( .A(n32578), .Z(n32580) );
  XOR U32997 ( .A(n32581), .B(g_input[819]), .Z(n32578) );
  NAND U32998 ( .A(n32582), .B(mul_pow), .Z(n32581) );
  XOR U32999 ( .A(g_input[819]), .B(creg[819]), .Z(n32582) );
  XOR U33000 ( .A(n32583), .B(n32584), .Z(n32574) );
  ANDN U33001 ( .A(n32585), .B(n25832), .Z(n32584) );
  XOR U33002 ( .A(n32586), .B(\modmult_1/zin[0][817] ), .Z(n25832) );
  IV U33003 ( .A(n32583), .Z(n32586) );
  XNOR U33004 ( .A(n32583), .B(n25831), .Z(n32585) );
  XOR U33005 ( .A(n32587), .B(n32588), .Z(n25831) );
  AND U33006 ( .A(\modmult_1/xin[1023] ), .B(n32589), .Z(n32588) );
  IV U33007 ( .A(n32587), .Z(n32589) );
  XOR U33008 ( .A(n32590), .B(g_input[818]), .Z(n32587) );
  NAND U33009 ( .A(n32591), .B(mul_pow), .Z(n32590) );
  XOR U33010 ( .A(g_input[818]), .B(creg[818]), .Z(n32591) );
  XOR U33011 ( .A(n32592), .B(n32593), .Z(n32583) );
  ANDN U33012 ( .A(n32594), .B(n25838), .Z(n32593) );
  XOR U33013 ( .A(n32595), .B(\modmult_1/zin[0][816] ), .Z(n25838) );
  IV U33014 ( .A(n32592), .Z(n32595) );
  XNOR U33015 ( .A(n32592), .B(n25837), .Z(n32594) );
  XOR U33016 ( .A(n32596), .B(n32597), .Z(n25837) );
  AND U33017 ( .A(\modmult_1/xin[1023] ), .B(n32598), .Z(n32597) );
  IV U33018 ( .A(n32596), .Z(n32598) );
  XOR U33019 ( .A(n32599), .B(g_input[817]), .Z(n32596) );
  NAND U33020 ( .A(n32600), .B(mul_pow), .Z(n32599) );
  XOR U33021 ( .A(g_input[817]), .B(creg[817]), .Z(n32600) );
  XOR U33022 ( .A(n32601), .B(n32602), .Z(n32592) );
  ANDN U33023 ( .A(n32603), .B(n25844), .Z(n32602) );
  XOR U33024 ( .A(n32604), .B(\modmult_1/zin[0][815] ), .Z(n25844) );
  IV U33025 ( .A(n32601), .Z(n32604) );
  XNOR U33026 ( .A(n32601), .B(n25843), .Z(n32603) );
  XOR U33027 ( .A(n32605), .B(n32606), .Z(n25843) );
  AND U33028 ( .A(\modmult_1/xin[1023] ), .B(n32607), .Z(n32606) );
  IV U33029 ( .A(n32605), .Z(n32607) );
  XOR U33030 ( .A(n32608), .B(g_input[816]), .Z(n32605) );
  NAND U33031 ( .A(n32609), .B(mul_pow), .Z(n32608) );
  XOR U33032 ( .A(g_input[816]), .B(creg[816]), .Z(n32609) );
  XOR U33033 ( .A(n32610), .B(n32611), .Z(n32601) );
  ANDN U33034 ( .A(n32612), .B(n25850), .Z(n32611) );
  XOR U33035 ( .A(n32613), .B(\modmult_1/zin[0][814] ), .Z(n25850) );
  IV U33036 ( .A(n32610), .Z(n32613) );
  XNOR U33037 ( .A(n32610), .B(n25849), .Z(n32612) );
  XOR U33038 ( .A(n32614), .B(n32615), .Z(n25849) );
  AND U33039 ( .A(\modmult_1/xin[1023] ), .B(n32616), .Z(n32615) );
  IV U33040 ( .A(n32614), .Z(n32616) );
  XOR U33041 ( .A(n32617), .B(g_input[815]), .Z(n32614) );
  NAND U33042 ( .A(n32618), .B(mul_pow), .Z(n32617) );
  XOR U33043 ( .A(g_input[815]), .B(creg[815]), .Z(n32618) );
  XOR U33044 ( .A(n32619), .B(n32620), .Z(n32610) );
  ANDN U33045 ( .A(n32621), .B(n25856), .Z(n32620) );
  XOR U33046 ( .A(n32622), .B(\modmult_1/zin[0][813] ), .Z(n25856) );
  IV U33047 ( .A(n32619), .Z(n32622) );
  XNOR U33048 ( .A(n32619), .B(n25855), .Z(n32621) );
  XOR U33049 ( .A(n32623), .B(n32624), .Z(n25855) );
  AND U33050 ( .A(\modmult_1/xin[1023] ), .B(n32625), .Z(n32624) );
  IV U33051 ( .A(n32623), .Z(n32625) );
  XOR U33052 ( .A(n32626), .B(g_input[814]), .Z(n32623) );
  NAND U33053 ( .A(n32627), .B(mul_pow), .Z(n32626) );
  XOR U33054 ( .A(g_input[814]), .B(creg[814]), .Z(n32627) );
  XOR U33055 ( .A(n32628), .B(n32629), .Z(n32619) );
  ANDN U33056 ( .A(n32630), .B(n25862), .Z(n32629) );
  XOR U33057 ( .A(n32631), .B(\modmult_1/zin[0][812] ), .Z(n25862) );
  IV U33058 ( .A(n32628), .Z(n32631) );
  XNOR U33059 ( .A(n32628), .B(n25861), .Z(n32630) );
  XOR U33060 ( .A(n32632), .B(n32633), .Z(n25861) );
  AND U33061 ( .A(\modmult_1/xin[1023] ), .B(n32634), .Z(n32633) );
  IV U33062 ( .A(n32632), .Z(n32634) );
  XOR U33063 ( .A(n32635), .B(g_input[813]), .Z(n32632) );
  NAND U33064 ( .A(n32636), .B(mul_pow), .Z(n32635) );
  XOR U33065 ( .A(g_input[813]), .B(creg[813]), .Z(n32636) );
  XOR U33066 ( .A(n32637), .B(n32638), .Z(n32628) );
  ANDN U33067 ( .A(n32639), .B(n25868), .Z(n32638) );
  XOR U33068 ( .A(n32640), .B(\modmult_1/zin[0][811] ), .Z(n25868) );
  IV U33069 ( .A(n32637), .Z(n32640) );
  XNOR U33070 ( .A(n32637), .B(n25867), .Z(n32639) );
  XOR U33071 ( .A(n32641), .B(n32642), .Z(n25867) );
  AND U33072 ( .A(\modmult_1/xin[1023] ), .B(n32643), .Z(n32642) );
  IV U33073 ( .A(n32641), .Z(n32643) );
  XOR U33074 ( .A(n32644), .B(g_input[812]), .Z(n32641) );
  NAND U33075 ( .A(n32645), .B(mul_pow), .Z(n32644) );
  XOR U33076 ( .A(g_input[812]), .B(creg[812]), .Z(n32645) );
  XOR U33077 ( .A(n32646), .B(n32647), .Z(n32637) );
  ANDN U33078 ( .A(n32648), .B(n25874), .Z(n32647) );
  XOR U33079 ( .A(n32649), .B(\modmult_1/zin[0][810] ), .Z(n25874) );
  IV U33080 ( .A(n32646), .Z(n32649) );
  XNOR U33081 ( .A(n32646), .B(n25873), .Z(n32648) );
  XOR U33082 ( .A(n32650), .B(n32651), .Z(n25873) );
  AND U33083 ( .A(\modmult_1/xin[1023] ), .B(n32652), .Z(n32651) );
  IV U33084 ( .A(n32650), .Z(n32652) );
  XOR U33085 ( .A(n32653), .B(g_input[811]), .Z(n32650) );
  NAND U33086 ( .A(n32654), .B(mul_pow), .Z(n32653) );
  XOR U33087 ( .A(g_input[811]), .B(creg[811]), .Z(n32654) );
  XOR U33088 ( .A(n32655), .B(n32656), .Z(n32646) );
  ANDN U33089 ( .A(n32657), .B(n25880), .Z(n32656) );
  XOR U33090 ( .A(n32658), .B(\modmult_1/zin[0][809] ), .Z(n25880) );
  IV U33091 ( .A(n32655), .Z(n32658) );
  XNOR U33092 ( .A(n32655), .B(n25879), .Z(n32657) );
  XOR U33093 ( .A(n32659), .B(n32660), .Z(n25879) );
  AND U33094 ( .A(\modmult_1/xin[1023] ), .B(n32661), .Z(n32660) );
  IV U33095 ( .A(n32659), .Z(n32661) );
  XOR U33096 ( .A(n32662), .B(g_input[810]), .Z(n32659) );
  NAND U33097 ( .A(n32663), .B(mul_pow), .Z(n32662) );
  XOR U33098 ( .A(g_input[810]), .B(creg[810]), .Z(n32663) );
  XOR U33099 ( .A(n32664), .B(n32665), .Z(n32655) );
  ANDN U33100 ( .A(n32666), .B(n25886), .Z(n32665) );
  XOR U33101 ( .A(n32667), .B(\modmult_1/zin[0][808] ), .Z(n25886) );
  IV U33102 ( .A(n32664), .Z(n32667) );
  XNOR U33103 ( .A(n32664), .B(n25885), .Z(n32666) );
  XOR U33104 ( .A(n32668), .B(n32669), .Z(n25885) );
  AND U33105 ( .A(\modmult_1/xin[1023] ), .B(n32670), .Z(n32669) );
  IV U33106 ( .A(n32668), .Z(n32670) );
  XOR U33107 ( .A(n32671), .B(g_input[809]), .Z(n32668) );
  NAND U33108 ( .A(n32672), .B(mul_pow), .Z(n32671) );
  XOR U33109 ( .A(g_input[809]), .B(creg[809]), .Z(n32672) );
  XOR U33110 ( .A(n32673), .B(n32674), .Z(n32664) );
  ANDN U33111 ( .A(n32675), .B(n25892), .Z(n32674) );
  XOR U33112 ( .A(n32676), .B(\modmult_1/zin[0][807] ), .Z(n25892) );
  IV U33113 ( .A(n32673), .Z(n32676) );
  XNOR U33114 ( .A(n32673), .B(n25891), .Z(n32675) );
  XOR U33115 ( .A(n32677), .B(n32678), .Z(n25891) );
  AND U33116 ( .A(\modmult_1/xin[1023] ), .B(n32679), .Z(n32678) );
  IV U33117 ( .A(n32677), .Z(n32679) );
  XOR U33118 ( .A(n32680), .B(g_input[808]), .Z(n32677) );
  NAND U33119 ( .A(n32681), .B(mul_pow), .Z(n32680) );
  XOR U33120 ( .A(g_input[808]), .B(creg[808]), .Z(n32681) );
  XOR U33121 ( .A(n32682), .B(n32683), .Z(n32673) );
  ANDN U33122 ( .A(n32684), .B(n25898), .Z(n32683) );
  XOR U33123 ( .A(n32685), .B(\modmult_1/zin[0][806] ), .Z(n25898) );
  IV U33124 ( .A(n32682), .Z(n32685) );
  XNOR U33125 ( .A(n32682), .B(n25897), .Z(n32684) );
  XOR U33126 ( .A(n32686), .B(n32687), .Z(n25897) );
  AND U33127 ( .A(\modmult_1/xin[1023] ), .B(n32688), .Z(n32687) );
  IV U33128 ( .A(n32686), .Z(n32688) );
  XOR U33129 ( .A(n32689), .B(g_input[807]), .Z(n32686) );
  NAND U33130 ( .A(n32690), .B(mul_pow), .Z(n32689) );
  XOR U33131 ( .A(g_input[807]), .B(creg[807]), .Z(n32690) );
  XOR U33132 ( .A(n32691), .B(n32692), .Z(n32682) );
  ANDN U33133 ( .A(n32693), .B(n25904), .Z(n32692) );
  XOR U33134 ( .A(n32694), .B(\modmult_1/zin[0][805] ), .Z(n25904) );
  IV U33135 ( .A(n32691), .Z(n32694) );
  XNOR U33136 ( .A(n32691), .B(n25903), .Z(n32693) );
  XOR U33137 ( .A(n32695), .B(n32696), .Z(n25903) );
  AND U33138 ( .A(\modmult_1/xin[1023] ), .B(n32697), .Z(n32696) );
  IV U33139 ( .A(n32695), .Z(n32697) );
  XOR U33140 ( .A(n32698), .B(g_input[806]), .Z(n32695) );
  NAND U33141 ( .A(n32699), .B(mul_pow), .Z(n32698) );
  XOR U33142 ( .A(g_input[806]), .B(creg[806]), .Z(n32699) );
  XOR U33143 ( .A(n32700), .B(n32701), .Z(n32691) );
  ANDN U33144 ( .A(n32702), .B(n25910), .Z(n32701) );
  XOR U33145 ( .A(n32703), .B(\modmult_1/zin[0][804] ), .Z(n25910) );
  IV U33146 ( .A(n32700), .Z(n32703) );
  XNOR U33147 ( .A(n32700), .B(n25909), .Z(n32702) );
  XOR U33148 ( .A(n32704), .B(n32705), .Z(n25909) );
  AND U33149 ( .A(\modmult_1/xin[1023] ), .B(n32706), .Z(n32705) );
  IV U33150 ( .A(n32704), .Z(n32706) );
  XOR U33151 ( .A(n32707), .B(g_input[805]), .Z(n32704) );
  NAND U33152 ( .A(n32708), .B(mul_pow), .Z(n32707) );
  XOR U33153 ( .A(g_input[805]), .B(creg[805]), .Z(n32708) );
  XOR U33154 ( .A(n32709), .B(n32710), .Z(n32700) );
  ANDN U33155 ( .A(n32711), .B(n25916), .Z(n32710) );
  XOR U33156 ( .A(n32712), .B(\modmult_1/zin[0][803] ), .Z(n25916) );
  IV U33157 ( .A(n32709), .Z(n32712) );
  XNOR U33158 ( .A(n32709), .B(n25915), .Z(n32711) );
  XOR U33159 ( .A(n32713), .B(n32714), .Z(n25915) );
  AND U33160 ( .A(\modmult_1/xin[1023] ), .B(n32715), .Z(n32714) );
  IV U33161 ( .A(n32713), .Z(n32715) );
  XOR U33162 ( .A(n32716), .B(g_input[804]), .Z(n32713) );
  NAND U33163 ( .A(n32717), .B(mul_pow), .Z(n32716) );
  XOR U33164 ( .A(g_input[804]), .B(creg[804]), .Z(n32717) );
  XOR U33165 ( .A(n32718), .B(n32719), .Z(n32709) );
  ANDN U33166 ( .A(n32720), .B(n25922), .Z(n32719) );
  XOR U33167 ( .A(n32721), .B(\modmult_1/zin[0][802] ), .Z(n25922) );
  IV U33168 ( .A(n32718), .Z(n32721) );
  XNOR U33169 ( .A(n32718), .B(n25921), .Z(n32720) );
  XOR U33170 ( .A(n32722), .B(n32723), .Z(n25921) );
  AND U33171 ( .A(\modmult_1/xin[1023] ), .B(n32724), .Z(n32723) );
  IV U33172 ( .A(n32722), .Z(n32724) );
  XOR U33173 ( .A(n32725), .B(g_input[803]), .Z(n32722) );
  NAND U33174 ( .A(n32726), .B(mul_pow), .Z(n32725) );
  XOR U33175 ( .A(g_input[803]), .B(creg[803]), .Z(n32726) );
  XOR U33176 ( .A(n32727), .B(n32728), .Z(n32718) );
  ANDN U33177 ( .A(n32729), .B(n25928), .Z(n32728) );
  XOR U33178 ( .A(n32730), .B(\modmult_1/zin[0][801] ), .Z(n25928) );
  IV U33179 ( .A(n32727), .Z(n32730) );
  XNOR U33180 ( .A(n32727), .B(n25927), .Z(n32729) );
  XOR U33181 ( .A(n32731), .B(n32732), .Z(n25927) );
  AND U33182 ( .A(\modmult_1/xin[1023] ), .B(n32733), .Z(n32732) );
  IV U33183 ( .A(n32731), .Z(n32733) );
  XOR U33184 ( .A(n32734), .B(g_input[802]), .Z(n32731) );
  NAND U33185 ( .A(n32735), .B(mul_pow), .Z(n32734) );
  XOR U33186 ( .A(g_input[802]), .B(creg[802]), .Z(n32735) );
  XOR U33187 ( .A(n32736), .B(n32737), .Z(n32727) );
  ANDN U33188 ( .A(n32738), .B(n25934), .Z(n32737) );
  XOR U33189 ( .A(n32739), .B(\modmult_1/zin[0][800] ), .Z(n25934) );
  IV U33190 ( .A(n32736), .Z(n32739) );
  XNOR U33191 ( .A(n32736), .B(n25933), .Z(n32738) );
  XOR U33192 ( .A(n32740), .B(n32741), .Z(n25933) );
  AND U33193 ( .A(\modmult_1/xin[1023] ), .B(n32742), .Z(n32741) );
  IV U33194 ( .A(n32740), .Z(n32742) );
  XOR U33195 ( .A(n32743), .B(g_input[801]), .Z(n32740) );
  NAND U33196 ( .A(n32744), .B(mul_pow), .Z(n32743) );
  XOR U33197 ( .A(g_input[801]), .B(creg[801]), .Z(n32744) );
  XOR U33198 ( .A(n32745), .B(n32746), .Z(n32736) );
  ANDN U33199 ( .A(n32747), .B(n25940), .Z(n32746) );
  XOR U33200 ( .A(n32748), .B(\modmult_1/zin[0][799] ), .Z(n25940) );
  IV U33201 ( .A(n32745), .Z(n32748) );
  XNOR U33202 ( .A(n32745), .B(n25939), .Z(n32747) );
  XOR U33203 ( .A(n32749), .B(n32750), .Z(n25939) );
  AND U33204 ( .A(\modmult_1/xin[1023] ), .B(n32751), .Z(n32750) );
  IV U33205 ( .A(n32749), .Z(n32751) );
  XOR U33206 ( .A(n32752), .B(g_input[800]), .Z(n32749) );
  NAND U33207 ( .A(n32753), .B(mul_pow), .Z(n32752) );
  XOR U33208 ( .A(g_input[800]), .B(creg[800]), .Z(n32753) );
  XOR U33209 ( .A(n32754), .B(n32755), .Z(n32745) );
  ANDN U33210 ( .A(n32756), .B(n25946), .Z(n32755) );
  XOR U33211 ( .A(n32757), .B(\modmult_1/zin[0][798] ), .Z(n25946) );
  IV U33212 ( .A(n32754), .Z(n32757) );
  XNOR U33213 ( .A(n32754), .B(n25945), .Z(n32756) );
  XOR U33214 ( .A(n32758), .B(n32759), .Z(n25945) );
  AND U33215 ( .A(\modmult_1/xin[1023] ), .B(n32760), .Z(n32759) );
  IV U33216 ( .A(n32758), .Z(n32760) );
  XOR U33217 ( .A(n32761), .B(g_input[799]), .Z(n32758) );
  NAND U33218 ( .A(n32762), .B(mul_pow), .Z(n32761) );
  XOR U33219 ( .A(g_input[799]), .B(creg[799]), .Z(n32762) );
  XOR U33220 ( .A(n32763), .B(n32764), .Z(n32754) );
  ANDN U33221 ( .A(n32765), .B(n25952), .Z(n32764) );
  XOR U33222 ( .A(n32766), .B(\modmult_1/zin[0][797] ), .Z(n25952) );
  IV U33223 ( .A(n32763), .Z(n32766) );
  XNOR U33224 ( .A(n32763), .B(n25951), .Z(n32765) );
  XOR U33225 ( .A(n32767), .B(n32768), .Z(n25951) );
  AND U33226 ( .A(\modmult_1/xin[1023] ), .B(n32769), .Z(n32768) );
  IV U33227 ( .A(n32767), .Z(n32769) );
  XOR U33228 ( .A(n32770), .B(g_input[798]), .Z(n32767) );
  NAND U33229 ( .A(n32771), .B(mul_pow), .Z(n32770) );
  XOR U33230 ( .A(g_input[798]), .B(creg[798]), .Z(n32771) );
  XOR U33231 ( .A(n32772), .B(n32773), .Z(n32763) );
  ANDN U33232 ( .A(n32774), .B(n25958), .Z(n32773) );
  XOR U33233 ( .A(n32775), .B(\modmult_1/zin[0][796] ), .Z(n25958) );
  IV U33234 ( .A(n32772), .Z(n32775) );
  XNOR U33235 ( .A(n32772), .B(n25957), .Z(n32774) );
  XOR U33236 ( .A(n32776), .B(n32777), .Z(n25957) );
  AND U33237 ( .A(\modmult_1/xin[1023] ), .B(n32778), .Z(n32777) );
  IV U33238 ( .A(n32776), .Z(n32778) );
  XOR U33239 ( .A(n32779), .B(g_input[797]), .Z(n32776) );
  NAND U33240 ( .A(n32780), .B(mul_pow), .Z(n32779) );
  XOR U33241 ( .A(g_input[797]), .B(creg[797]), .Z(n32780) );
  XOR U33242 ( .A(n32781), .B(n32782), .Z(n32772) );
  ANDN U33243 ( .A(n32783), .B(n25964), .Z(n32782) );
  XOR U33244 ( .A(n32784), .B(\modmult_1/zin[0][795] ), .Z(n25964) );
  IV U33245 ( .A(n32781), .Z(n32784) );
  XNOR U33246 ( .A(n32781), .B(n25963), .Z(n32783) );
  XOR U33247 ( .A(n32785), .B(n32786), .Z(n25963) );
  AND U33248 ( .A(\modmult_1/xin[1023] ), .B(n32787), .Z(n32786) );
  IV U33249 ( .A(n32785), .Z(n32787) );
  XOR U33250 ( .A(n32788), .B(g_input[796]), .Z(n32785) );
  NAND U33251 ( .A(n32789), .B(mul_pow), .Z(n32788) );
  XOR U33252 ( .A(g_input[796]), .B(creg[796]), .Z(n32789) );
  XOR U33253 ( .A(n32790), .B(n32791), .Z(n32781) );
  ANDN U33254 ( .A(n32792), .B(n25970), .Z(n32791) );
  XOR U33255 ( .A(n32793), .B(\modmult_1/zin[0][794] ), .Z(n25970) );
  IV U33256 ( .A(n32790), .Z(n32793) );
  XNOR U33257 ( .A(n32790), .B(n25969), .Z(n32792) );
  XOR U33258 ( .A(n32794), .B(n32795), .Z(n25969) );
  AND U33259 ( .A(\modmult_1/xin[1023] ), .B(n32796), .Z(n32795) );
  IV U33260 ( .A(n32794), .Z(n32796) );
  XOR U33261 ( .A(n32797), .B(g_input[795]), .Z(n32794) );
  NAND U33262 ( .A(n32798), .B(mul_pow), .Z(n32797) );
  XOR U33263 ( .A(g_input[795]), .B(creg[795]), .Z(n32798) );
  XOR U33264 ( .A(n32799), .B(n32800), .Z(n32790) );
  ANDN U33265 ( .A(n32801), .B(n25976), .Z(n32800) );
  XOR U33266 ( .A(n32802), .B(\modmult_1/zin[0][793] ), .Z(n25976) );
  IV U33267 ( .A(n32799), .Z(n32802) );
  XNOR U33268 ( .A(n32799), .B(n25975), .Z(n32801) );
  XOR U33269 ( .A(n32803), .B(n32804), .Z(n25975) );
  AND U33270 ( .A(\modmult_1/xin[1023] ), .B(n32805), .Z(n32804) );
  IV U33271 ( .A(n32803), .Z(n32805) );
  XOR U33272 ( .A(n32806), .B(g_input[794]), .Z(n32803) );
  NAND U33273 ( .A(n32807), .B(mul_pow), .Z(n32806) );
  XOR U33274 ( .A(g_input[794]), .B(creg[794]), .Z(n32807) );
  XOR U33275 ( .A(n32808), .B(n32809), .Z(n32799) );
  ANDN U33276 ( .A(n32810), .B(n25982), .Z(n32809) );
  XOR U33277 ( .A(n32811), .B(\modmult_1/zin[0][792] ), .Z(n25982) );
  IV U33278 ( .A(n32808), .Z(n32811) );
  XNOR U33279 ( .A(n32808), .B(n25981), .Z(n32810) );
  XOR U33280 ( .A(n32812), .B(n32813), .Z(n25981) );
  AND U33281 ( .A(\modmult_1/xin[1023] ), .B(n32814), .Z(n32813) );
  IV U33282 ( .A(n32812), .Z(n32814) );
  XOR U33283 ( .A(n32815), .B(g_input[793]), .Z(n32812) );
  NAND U33284 ( .A(n32816), .B(mul_pow), .Z(n32815) );
  XOR U33285 ( .A(g_input[793]), .B(creg[793]), .Z(n32816) );
  XOR U33286 ( .A(n32817), .B(n32818), .Z(n32808) );
  ANDN U33287 ( .A(n32819), .B(n25988), .Z(n32818) );
  XOR U33288 ( .A(n32820), .B(\modmult_1/zin[0][791] ), .Z(n25988) );
  IV U33289 ( .A(n32817), .Z(n32820) );
  XNOR U33290 ( .A(n32817), .B(n25987), .Z(n32819) );
  XOR U33291 ( .A(n32821), .B(n32822), .Z(n25987) );
  AND U33292 ( .A(\modmult_1/xin[1023] ), .B(n32823), .Z(n32822) );
  IV U33293 ( .A(n32821), .Z(n32823) );
  XOR U33294 ( .A(n32824), .B(g_input[792]), .Z(n32821) );
  NAND U33295 ( .A(n32825), .B(mul_pow), .Z(n32824) );
  XOR U33296 ( .A(g_input[792]), .B(creg[792]), .Z(n32825) );
  XOR U33297 ( .A(n32826), .B(n32827), .Z(n32817) );
  ANDN U33298 ( .A(n32828), .B(n25994), .Z(n32827) );
  XOR U33299 ( .A(n32829), .B(\modmult_1/zin[0][790] ), .Z(n25994) );
  IV U33300 ( .A(n32826), .Z(n32829) );
  XNOR U33301 ( .A(n32826), .B(n25993), .Z(n32828) );
  XOR U33302 ( .A(n32830), .B(n32831), .Z(n25993) );
  AND U33303 ( .A(\modmult_1/xin[1023] ), .B(n32832), .Z(n32831) );
  IV U33304 ( .A(n32830), .Z(n32832) );
  XOR U33305 ( .A(n32833), .B(g_input[791]), .Z(n32830) );
  NAND U33306 ( .A(n32834), .B(mul_pow), .Z(n32833) );
  XOR U33307 ( .A(g_input[791]), .B(creg[791]), .Z(n32834) );
  XOR U33308 ( .A(n32835), .B(n32836), .Z(n32826) );
  ANDN U33309 ( .A(n32837), .B(n26000), .Z(n32836) );
  XOR U33310 ( .A(n32838), .B(\modmult_1/zin[0][789] ), .Z(n26000) );
  IV U33311 ( .A(n32835), .Z(n32838) );
  XNOR U33312 ( .A(n32835), .B(n25999), .Z(n32837) );
  XOR U33313 ( .A(n32839), .B(n32840), .Z(n25999) );
  AND U33314 ( .A(\modmult_1/xin[1023] ), .B(n32841), .Z(n32840) );
  IV U33315 ( .A(n32839), .Z(n32841) );
  XOR U33316 ( .A(n32842), .B(g_input[790]), .Z(n32839) );
  NAND U33317 ( .A(n32843), .B(mul_pow), .Z(n32842) );
  XOR U33318 ( .A(g_input[790]), .B(creg[790]), .Z(n32843) );
  XOR U33319 ( .A(n32844), .B(n32845), .Z(n32835) );
  ANDN U33320 ( .A(n32846), .B(n26006), .Z(n32845) );
  XOR U33321 ( .A(n32847), .B(\modmult_1/zin[0][788] ), .Z(n26006) );
  IV U33322 ( .A(n32844), .Z(n32847) );
  XNOR U33323 ( .A(n32844), .B(n26005), .Z(n32846) );
  XOR U33324 ( .A(n32848), .B(n32849), .Z(n26005) );
  AND U33325 ( .A(\modmult_1/xin[1023] ), .B(n32850), .Z(n32849) );
  IV U33326 ( .A(n32848), .Z(n32850) );
  XOR U33327 ( .A(n32851), .B(g_input[789]), .Z(n32848) );
  NAND U33328 ( .A(n32852), .B(mul_pow), .Z(n32851) );
  XOR U33329 ( .A(g_input[789]), .B(creg[789]), .Z(n32852) );
  XOR U33330 ( .A(n32853), .B(n32854), .Z(n32844) );
  ANDN U33331 ( .A(n32855), .B(n26012), .Z(n32854) );
  XOR U33332 ( .A(n32856), .B(\modmult_1/zin[0][787] ), .Z(n26012) );
  IV U33333 ( .A(n32853), .Z(n32856) );
  XNOR U33334 ( .A(n32853), .B(n26011), .Z(n32855) );
  XOR U33335 ( .A(n32857), .B(n32858), .Z(n26011) );
  AND U33336 ( .A(\modmult_1/xin[1023] ), .B(n32859), .Z(n32858) );
  IV U33337 ( .A(n32857), .Z(n32859) );
  XOR U33338 ( .A(n32860), .B(g_input[788]), .Z(n32857) );
  NAND U33339 ( .A(n32861), .B(mul_pow), .Z(n32860) );
  XOR U33340 ( .A(g_input[788]), .B(creg[788]), .Z(n32861) );
  XOR U33341 ( .A(n32862), .B(n32863), .Z(n32853) );
  ANDN U33342 ( .A(n32864), .B(n26018), .Z(n32863) );
  XOR U33343 ( .A(n32865), .B(\modmult_1/zin[0][786] ), .Z(n26018) );
  IV U33344 ( .A(n32862), .Z(n32865) );
  XNOR U33345 ( .A(n32862), .B(n26017), .Z(n32864) );
  XOR U33346 ( .A(n32866), .B(n32867), .Z(n26017) );
  AND U33347 ( .A(\modmult_1/xin[1023] ), .B(n32868), .Z(n32867) );
  IV U33348 ( .A(n32866), .Z(n32868) );
  XOR U33349 ( .A(n32869), .B(g_input[787]), .Z(n32866) );
  NAND U33350 ( .A(n32870), .B(mul_pow), .Z(n32869) );
  XOR U33351 ( .A(g_input[787]), .B(creg[787]), .Z(n32870) );
  XOR U33352 ( .A(n32871), .B(n32872), .Z(n32862) );
  ANDN U33353 ( .A(n32873), .B(n26024), .Z(n32872) );
  XOR U33354 ( .A(n32874), .B(\modmult_1/zin[0][785] ), .Z(n26024) );
  IV U33355 ( .A(n32871), .Z(n32874) );
  XNOR U33356 ( .A(n32871), .B(n26023), .Z(n32873) );
  XOR U33357 ( .A(n32875), .B(n32876), .Z(n26023) );
  AND U33358 ( .A(\modmult_1/xin[1023] ), .B(n32877), .Z(n32876) );
  IV U33359 ( .A(n32875), .Z(n32877) );
  XOR U33360 ( .A(n32878), .B(g_input[786]), .Z(n32875) );
  NAND U33361 ( .A(n32879), .B(mul_pow), .Z(n32878) );
  XOR U33362 ( .A(g_input[786]), .B(creg[786]), .Z(n32879) );
  XOR U33363 ( .A(n32880), .B(n32881), .Z(n32871) );
  ANDN U33364 ( .A(n32882), .B(n26030), .Z(n32881) );
  XOR U33365 ( .A(n32883), .B(\modmult_1/zin[0][784] ), .Z(n26030) );
  IV U33366 ( .A(n32880), .Z(n32883) );
  XNOR U33367 ( .A(n32880), .B(n26029), .Z(n32882) );
  XOR U33368 ( .A(n32884), .B(n32885), .Z(n26029) );
  AND U33369 ( .A(\modmult_1/xin[1023] ), .B(n32886), .Z(n32885) );
  IV U33370 ( .A(n32884), .Z(n32886) );
  XOR U33371 ( .A(n32887), .B(g_input[785]), .Z(n32884) );
  NAND U33372 ( .A(n32888), .B(mul_pow), .Z(n32887) );
  XOR U33373 ( .A(g_input[785]), .B(creg[785]), .Z(n32888) );
  XOR U33374 ( .A(n32889), .B(n32890), .Z(n32880) );
  ANDN U33375 ( .A(n32891), .B(n26036), .Z(n32890) );
  XOR U33376 ( .A(n32892), .B(\modmult_1/zin[0][783] ), .Z(n26036) );
  IV U33377 ( .A(n32889), .Z(n32892) );
  XNOR U33378 ( .A(n32889), .B(n26035), .Z(n32891) );
  XOR U33379 ( .A(n32893), .B(n32894), .Z(n26035) );
  AND U33380 ( .A(\modmult_1/xin[1023] ), .B(n32895), .Z(n32894) );
  IV U33381 ( .A(n32893), .Z(n32895) );
  XOR U33382 ( .A(n32896), .B(g_input[784]), .Z(n32893) );
  NAND U33383 ( .A(n32897), .B(mul_pow), .Z(n32896) );
  XOR U33384 ( .A(g_input[784]), .B(creg[784]), .Z(n32897) );
  XOR U33385 ( .A(n32898), .B(n32899), .Z(n32889) );
  ANDN U33386 ( .A(n32900), .B(n26042), .Z(n32899) );
  XOR U33387 ( .A(n32901), .B(\modmult_1/zin[0][782] ), .Z(n26042) );
  IV U33388 ( .A(n32898), .Z(n32901) );
  XNOR U33389 ( .A(n32898), .B(n26041), .Z(n32900) );
  XOR U33390 ( .A(n32902), .B(n32903), .Z(n26041) );
  AND U33391 ( .A(\modmult_1/xin[1023] ), .B(n32904), .Z(n32903) );
  IV U33392 ( .A(n32902), .Z(n32904) );
  XOR U33393 ( .A(n32905), .B(g_input[783]), .Z(n32902) );
  NAND U33394 ( .A(n32906), .B(mul_pow), .Z(n32905) );
  XOR U33395 ( .A(g_input[783]), .B(creg[783]), .Z(n32906) );
  XOR U33396 ( .A(n32907), .B(n32908), .Z(n32898) );
  ANDN U33397 ( .A(n32909), .B(n26048), .Z(n32908) );
  XOR U33398 ( .A(n32910), .B(\modmult_1/zin[0][781] ), .Z(n26048) );
  IV U33399 ( .A(n32907), .Z(n32910) );
  XNOR U33400 ( .A(n32907), .B(n26047), .Z(n32909) );
  XOR U33401 ( .A(n32911), .B(n32912), .Z(n26047) );
  AND U33402 ( .A(\modmult_1/xin[1023] ), .B(n32913), .Z(n32912) );
  IV U33403 ( .A(n32911), .Z(n32913) );
  XOR U33404 ( .A(n32914), .B(g_input[782]), .Z(n32911) );
  NAND U33405 ( .A(n32915), .B(mul_pow), .Z(n32914) );
  XOR U33406 ( .A(g_input[782]), .B(creg[782]), .Z(n32915) );
  XOR U33407 ( .A(n32916), .B(n32917), .Z(n32907) );
  ANDN U33408 ( .A(n32918), .B(n26054), .Z(n32917) );
  XOR U33409 ( .A(n32919), .B(\modmult_1/zin[0][780] ), .Z(n26054) );
  IV U33410 ( .A(n32916), .Z(n32919) );
  XNOR U33411 ( .A(n32916), .B(n26053), .Z(n32918) );
  XOR U33412 ( .A(n32920), .B(n32921), .Z(n26053) );
  AND U33413 ( .A(\modmult_1/xin[1023] ), .B(n32922), .Z(n32921) );
  IV U33414 ( .A(n32920), .Z(n32922) );
  XOR U33415 ( .A(n32923), .B(g_input[781]), .Z(n32920) );
  NAND U33416 ( .A(n32924), .B(mul_pow), .Z(n32923) );
  XOR U33417 ( .A(g_input[781]), .B(creg[781]), .Z(n32924) );
  XOR U33418 ( .A(n32925), .B(n32926), .Z(n32916) );
  ANDN U33419 ( .A(n32927), .B(n26060), .Z(n32926) );
  XOR U33420 ( .A(n32928), .B(\modmult_1/zin[0][779] ), .Z(n26060) );
  IV U33421 ( .A(n32925), .Z(n32928) );
  XNOR U33422 ( .A(n32925), .B(n26059), .Z(n32927) );
  XOR U33423 ( .A(n32929), .B(n32930), .Z(n26059) );
  AND U33424 ( .A(\modmult_1/xin[1023] ), .B(n32931), .Z(n32930) );
  IV U33425 ( .A(n32929), .Z(n32931) );
  XOR U33426 ( .A(n32932), .B(g_input[780]), .Z(n32929) );
  NAND U33427 ( .A(n32933), .B(mul_pow), .Z(n32932) );
  XOR U33428 ( .A(g_input[780]), .B(creg[780]), .Z(n32933) );
  XOR U33429 ( .A(n32934), .B(n32935), .Z(n32925) );
  ANDN U33430 ( .A(n32936), .B(n26066), .Z(n32935) );
  XOR U33431 ( .A(n32937), .B(\modmult_1/zin[0][778] ), .Z(n26066) );
  IV U33432 ( .A(n32934), .Z(n32937) );
  XNOR U33433 ( .A(n32934), .B(n26065), .Z(n32936) );
  XOR U33434 ( .A(n32938), .B(n32939), .Z(n26065) );
  AND U33435 ( .A(\modmult_1/xin[1023] ), .B(n32940), .Z(n32939) );
  IV U33436 ( .A(n32938), .Z(n32940) );
  XOR U33437 ( .A(n32941), .B(g_input[779]), .Z(n32938) );
  NAND U33438 ( .A(n32942), .B(mul_pow), .Z(n32941) );
  XOR U33439 ( .A(g_input[779]), .B(creg[779]), .Z(n32942) );
  XOR U33440 ( .A(n32943), .B(n32944), .Z(n32934) );
  ANDN U33441 ( .A(n32945), .B(n26072), .Z(n32944) );
  XOR U33442 ( .A(n32946), .B(\modmult_1/zin[0][777] ), .Z(n26072) );
  IV U33443 ( .A(n32943), .Z(n32946) );
  XNOR U33444 ( .A(n32943), .B(n26071), .Z(n32945) );
  XOR U33445 ( .A(n32947), .B(n32948), .Z(n26071) );
  AND U33446 ( .A(\modmult_1/xin[1023] ), .B(n32949), .Z(n32948) );
  IV U33447 ( .A(n32947), .Z(n32949) );
  XOR U33448 ( .A(n32950), .B(g_input[778]), .Z(n32947) );
  NAND U33449 ( .A(n32951), .B(mul_pow), .Z(n32950) );
  XOR U33450 ( .A(g_input[778]), .B(creg[778]), .Z(n32951) );
  XOR U33451 ( .A(n32952), .B(n32953), .Z(n32943) );
  ANDN U33452 ( .A(n32954), .B(n26078), .Z(n32953) );
  XOR U33453 ( .A(n32955), .B(\modmult_1/zin[0][776] ), .Z(n26078) );
  IV U33454 ( .A(n32952), .Z(n32955) );
  XNOR U33455 ( .A(n32952), .B(n26077), .Z(n32954) );
  XOR U33456 ( .A(n32956), .B(n32957), .Z(n26077) );
  AND U33457 ( .A(\modmult_1/xin[1023] ), .B(n32958), .Z(n32957) );
  IV U33458 ( .A(n32956), .Z(n32958) );
  XOR U33459 ( .A(n32959), .B(g_input[777]), .Z(n32956) );
  NAND U33460 ( .A(n32960), .B(mul_pow), .Z(n32959) );
  XOR U33461 ( .A(g_input[777]), .B(creg[777]), .Z(n32960) );
  XOR U33462 ( .A(n32961), .B(n32962), .Z(n32952) );
  ANDN U33463 ( .A(n32963), .B(n26084), .Z(n32962) );
  XOR U33464 ( .A(n32964), .B(\modmult_1/zin[0][775] ), .Z(n26084) );
  IV U33465 ( .A(n32961), .Z(n32964) );
  XNOR U33466 ( .A(n32961), .B(n26083), .Z(n32963) );
  XOR U33467 ( .A(n32965), .B(n32966), .Z(n26083) );
  AND U33468 ( .A(\modmult_1/xin[1023] ), .B(n32967), .Z(n32966) );
  IV U33469 ( .A(n32965), .Z(n32967) );
  XOR U33470 ( .A(n32968), .B(g_input[776]), .Z(n32965) );
  NAND U33471 ( .A(n32969), .B(mul_pow), .Z(n32968) );
  XOR U33472 ( .A(g_input[776]), .B(creg[776]), .Z(n32969) );
  XOR U33473 ( .A(n32970), .B(n32971), .Z(n32961) );
  ANDN U33474 ( .A(n32972), .B(n26090), .Z(n32971) );
  XOR U33475 ( .A(n32973), .B(\modmult_1/zin[0][774] ), .Z(n26090) );
  IV U33476 ( .A(n32970), .Z(n32973) );
  XNOR U33477 ( .A(n32970), .B(n26089), .Z(n32972) );
  XOR U33478 ( .A(n32974), .B(n32975), .Z(n26089) );
  AND U33479 ( .A(\modmult_1/xin[1023] ), .B(n32976), .Z(n32975) );
  IV U33480 ( .A(n32974), .Z(n32976) );
  XOR U33481 ( .A(n32977), .B(g_input[775]), .Z(n32974) );
  NAND U33482 ( .A(n32978), .B(mul_pow), .Z(n32977) );
  XOR U33483 ( .A(g_input[775]), .B(creg[775]), .Z(n32978) );
  XOR U33484 ( .A(n32979), .B(n32980), .Z(n32970) );
  ANDN U33485 ( .A(n32981), .B(n26096), .Z(n32980) );
  XOR U33486 ( .A(n32982), .B(\modmult_1/zin[0][773] ), .Z(n26096) );
  IV U33487 ( .A(n32979), .Z(n32982) );
  XNOR U33488 ( .A(n32979), .B(n26095), .Z(n32981) );
  XOR U33489 ( .A(n32983), .B(n32984), .Z(n26095) );
  AND U33490 ( .A(\modmult_1/xin[1023] ), .B(n32985), .Z(n32984) );
  IV U33491 ( .A(n32983), .Z(n32985) );
  XOR U33492 ( .A(n32986), .B(g_input[774]), .Z(n32983) );
  NAND U33493 ( .A(n32987), .B(mul_pow), .Z(n32986) );
  XOR U33494 ( .A(g_input[774]), .B(creg[774]), .Z(n32987) );
  XOR U33495 ( .A(n32988), .B(n32989), .Z(n32979) );
  ANDN U33496 ( .A(n32990), .B(n26102), .Z(n32989) );
  XOR U33497 ( .A(n32991), .B(\modmult_1/zin[0][772] ), .Z(n26102) );
  IV U33498 ( .A(n32988), .Z(n32991) );
  XNOR U33499 ( .A(n32988), .B(n26101), .Z(n32990) );
  XOR U33500 ( .A(n32992), .B(n32993), .Z(n26101) );
  AND U33501 ( .A(\modmult_1/xin[1023] ), .B(n32994), .Z(n32993) );
  IV U33502 ( .A(n32992), .Z(n32994) );
  XOR U33503 ( .A(n32995), .B(g_input[773]), .Z(n32992) );
  NAND U33504 ( .A(n32996), .B(mul_pow), .Z(n32995) );
  XOR U33505 ( .A(g_input[773]), .B(creg[773]), .Z(n32996) );
  XOR U33506 ( .A(n32997), .B(n32998), .Z(n32988) );
  ANDN U33507 ( .A(n32999), .B(n26108), .Z(n32998) );
  XOR U33508 ( .A(n33000), .B(\modmult_1/zin[0][771] ), .Z(n26108) );
  IV U33509 ( .A(n32997), .Z(n33000) );
  XNOR U33510 ( .A(n32997), .B(n26107), .Z(n32999) );
  XOR U33511 ( .A(n33001), .B(n33002), .Z(n26107) );
  AND U33512 ( .A(\modmult_1/xin[1023] ), .B(n33003), .Z(n33002) );
  IV U33513 ( .A(n33001), .Z(n33003) );
  XOR U33514 ( .A(n33004), .B(g_input[772]), .Z(n33001) );
  NAND U33515 ( .A(n33005), .B(mul_pow), .Z(n33004) );
  XOR U33516 ( .A(g_input[772]), .B(creg[772]), .Z(n33005) );
  XOR U33517 ( .A(n33006), .B(n33007), .Z(n32997) );
  ANDN U33518 ( .A(n33008), .B(n26114), .Z(n33007) );
  XOR U33519 ( .A(n33009), .B(\modmult_1/zin[0][770] ), .Z(n26114) );
  IV U33520 ( .A(n33006), .Z(n33009) );
  XNOR U33521 ( .A(n33006), .B(n26113), .Z(n33008) );
  XOR U33522 ( .A(n33010), .B(n33011), .Z(n26113) );
  AND U33523 ( .A(\modmult_1/xin[1023] ), .B(n33012), .Z(n33011) );
  IV U33524 ( .A(n33010), .Z(n33012) );
  XOR U33525 ( .A(n33013), .B(g_input[771]), .Z(n33010) );
  NAND U33526 ( .A(n33014), .B(mul_pow), .Z(n33013) );
  XOR U33527 ( .A(g_input[771]), .B(creg[771]), .Z(n33014) );
  XOR U33528 ( .A(n33015), .B(n33016), .Z(n33006) );
  ANDN U33529 ( .A(n33017), .B(n26120), .Z(n33016) );
  XOR U33530 ( .A(n33018), .B(\modmult_1/zin[0][769] ), .Z(n26120) );
  IV U33531 ( .A(n33015), .Z(n33018) );
  XNOR U33532 ( .A(n33015), .B(n26119), .Z(n33017) );
  XOR U33533 ( .A(n33019), .B(n33020), .Z(n26119) );
  AND U33534 ( .A(\modmult_1/xin[1023] ), .B(n33021), .Z(n33020) );
  IV U33535 ( .A(n33019), .Z(n33021) );
  XOR U33536 ( .A(n33022), .B(g_input[770]), .Z(n33019) );
  NAND U33537 ( .A(n33023), .B(mul_pow), .Z(n33022) );
  XOR U33538 ( .A(g_input[770]), .B(creg[770]), .Z(n33023) );
  XOR U33539 ( .A(n33024), .B(n33025), .Z(n33015) );
  ANDN U33540 ( .A(n33026), .B(n26126), .Z(n33025) );
  XOR U33541 ( .A(n33027), .B(\modmult_1/zin[0][768] ), .Z(n26126) );
  IV U33542 ( .A(n33024), .Z(n33027) );
  XNOR U33543 ( .A(n33024), .B(n26125), .Z(n33026) );
  XOR U33544 ( .A(n33028), .B(n33029), .Z(n26125) );
  AND U33545 ( .A(\modmult_1/xin[1023] ), .B(n33030), .Z(n33029) );
  IV U33546 ( .A(n33028), .Z(n33030) );
  XOR U33547 ( .A(n33031), .B(g_input[769]), .Z(n33028) );
  NAND U33548 ( .A(n33032), .B(mul_pow), .Z(n33031) );
  XOR U33549 ( .A(g_input[769]), .B(creg[769]), .Z(n33032) );
  XOR U33550 ( .A(n33033), .B(n33034), .Z(n33024) );
  ANDN U33551 ( .A(n33035), .B(n26132), .Z(n33034) );
  XOR U33552 ( .A(n33036), .B(\modmult_1/zin[0][767] ), .Z(n26132) );
  IV U33553 ( .A(n33033), .Z(n33036) );
  XNOR U33554 ( .A(n33033), .B(n26131), .Z(n33035) );
  XOR U33555 ( .A(n33037), .B(n33038), .Z(n26131) );
  AND U33556 ( .A(\modmult_1/xin[1023] ), .B(n33039), .Z(n33038) );
  IV U33557 ( .A(n33037), .Z(n33039) );
  XOR U33558 ( .A(n33040), .B(g_input[768]), .Z(n33037) );
  NAND U33559 ( .A(n33041), .B(mul_pow), .Z(n33040) );
  XOR U33560 ( .A(g_input[768]), .B(creg[768]), .Z(n33041) );
  XOR U33561 ( .A(n33042), .B(n33043), .Z(n33033) );
  ANDN U33562 ( .A(n33044), .B(n26138), .Z(n33043) );
  XOR U33563 ( .A(n33045), .B(\modmult_1/zin[0][766] ), .Z(n26138) );
  IV U33564 ( .A(n33042), .Z(n33045) );
  XNOR U33565 ( .A(n33042), .B(n26137), .Z(n33044) );
  XOR U33566 ( .A(n33046), .B(n33047), .Z(n26137) );
  AND U33567 ( .A(\modmult_1/xin[1023] ), .B(n33048), .Z(n33047) );
  IV U33568 ( .A(n33046), .Z(n33048) );
  XOR U33569 ( .A(n33049), .B(g_input[767]), .Z(n33046) );
  NAND U33570 ( .A(n33050), .B(mul_pow), .Z(n33049) );
  XOR U33571 ( .A(g_input[767]), .B(creg[767]), .Z(n33050) );
  XOR U33572 ( .A(n33051), .B(n33052), .Z(n33042) );
  ANDN U33573 ( .A(n33053), .B(n26144), .Z(n33052) );
  XOR U33574 ( .A(n33054), .B(\modmult_1/zin[0][765] ), .Z(n26144) );
  IV U33575 ( .A(n33051), .Z(n33054) );
  XNOR U33576 ( .A(n33051), .B(n26143), .Z(n33053) );
  XOR U33577 ( .A(n33055), .B(n33056), .Z(n26143) );
  AND U33578 ( .A(\modmult_1/xin[1023] ), .B(n33057), .Z(n33056) );
  IV U33579 ( .A(n33055), .Z(n33057) );
  XOR U33580 ( .A(n33058), .B(g_input[766]), .Z(n33055) );
  NAND U33581 ( .A(n33059), .B(mul_pow), .Z(n33058) );
  XOR U33582 ( .A(g_input[766]), .B(creg[766]), .Z(n33059) );
  XOR U33583 ( .A(n33060), .B(n33061), .Z(n33051) );
  ANDN U33584 ( .A(n33062), .B(n26150), .Z(n33061) );
  XOR U33585 ( .A(n33063), .B(\modmult_1/zin[0][764] ), .Z(n26150) );
  IV U33586 ( .A(n33060), .Z(n33063) );
  XNOR U33587 ( .A(n33060), .B(n26149), .Z(n33062) );
  XOR U33588 ( .A(n33064), .B(n33065), .Z(n26149) );
  AND U33589 ( .A(\modmult_1/xin[1023] ), .B(n33066), .Z(n33065) );
  IV U33590 ( .A(n33064), .Z(n33066) );
  XOR U33591 ( .A(n33067), .B(g_input[765]), .Z(n33064) );
  NAND U33592 ( .A(n33068), .B(mul_pow), .Z(n33067) );
  XOR U33593 ( .A(g_input[765]), .B(creg[765]), .Z(n33068) );
  XOR U33594 ( .A(n33069), .B(n33070), .Z(n33060) );
  ANDN U33595 ( .A(n33071), .B(n26156), .Z(n33070) );
  XOR U33596 ( .A(n33072), .B(\modmult_1/zin[0][763] ), .Z(n26156) );
  IV U33597 ( .A(n33069), .Z(n33072) );
  XNOR U33598 ( .A(n33069), .B(n26155), .Z(n33071) );
  XOR U33599 ( .A(n33073), .B(n33074), .Z(n26155) );
  AND U33600 ( .A(\modmult_1/xin[1023] ), .B(n33075), .Z(n33074) );
  IV U33601 ( .A(n33073), .Z(n33075) );
  XOR U33602 ( .A(n33076), .B(g_input[764]), .Z(n33073) );
  NAND U33603 ( .A(n33077), .B(mul_pow), .Z(n33076) );
  XOR U33604 ( .A(g_input[764]), .B(creg[764]), .Z(n33077) );
  XOR U33605 ( .A(n33078), .B(n33079), .Z(n33069) );
  ANDN U33606 ( .A(n33080), .B(n26162), .Z(n33079) );
  XOR U33607 ( .A(n33081), .B(\modmult_1/zin[0][762] ), .Z(n26162) );
  IV U33608 ( .A(n33078), .Z(n33081) );
  XNOR U33609 ( .A(n33078), .B(n26161), .Z(n33080) );
  XOR U33610 ( .A(n33082), .B(n33083), .Z(n26161) );
  AND U33611 ( .A(\modmult_1/xin[1023] ), .B(n33084), .Z(n33083) );
  IV U33612 ( .A(n33082), .Z(n33084) );
  XOR U33613 ( .A(n33085), .B(g_input[763]), .Z(n33082) );
  NAND U33614 ( .A(n33086), .B(mul_pow), .Z(n33085) );
  XOR U33615 ( .A(g_input[763]), .B(creg[763]), .Z(n33086) );
  XOR U33616 ( .A(n33087), .B(n33088), .Z(n33078) );
  ANDN U33617 ( .A(n33089), .B(n26168), .Z(n33088) );
  XOR U33618 ( .A(n33090), .B(\modmult_1/zin[0][761] ), .Z(n26168) );
  IV U33619 ( .A(n33087), .Z(n33090) );
  XNOR U33620 ( .A(n33087), .B(n26167), .Z(n33089) );
  XOR U33621 ( .A(n33091), .B(n33092), .Z(n26167) );
  AND U33622 ( .A(\modmult_1/xin[1023] ), .B(n33093), .Z(n33092) );
  IV U33623 ( .A(n33091), .Z(n33093) );
  XOR U33624 ( .A(n33094), .B(g_input[762]), .Z(n33091) );
  NAND U33625 ( .A(n33095), .B(mul_pow), .Z(n33094) );
  XOR U33626 ( .A(g_input[762]), .B(creg[762]), .Z(n33095) );
  XOR U33627 ( .A(n33096), .B(n33097), .Z(n33087) );
  ANDN U33628 ( .A(n33098), .B(n26174), .Z(n33097) );
  XOR U33629 ( .A(n33099), .B(\modmult_1/zin[0][760] ), .Z(n26174) );
  IV U33630 ( .A(n33096), .Z(n33099) );
  XNOR U33631 ( .A(n33096), .B(n26173), .Z(n33098) );
  XOR U33632 ( .A(n33100), .B(n33101), .Z(n26173) );
  AND U33633 ( .A(\modmult_1/xin[1023] ), .B(n33102), .Z(n33101) );
  IV U33634 ( .A(n33100), .Z(n33102) );
  XOR U33635 ( .A(n33103), .B(g_input[761]), .Z(n33100) );
  NAND U33636 ( .A(n33104), .B(mul_pow), .Z(n33103) );
  XOR U33637 ( .A(g_input[761]), .B(creg[761]), .Z(n33104) );
  XOR U33638 ( .A(n33105), .B(n33106), .Z(n33096) );
  ANDN U33639 ( .A(n33107), .B(n26180), .Z(n33106) );
  XOR U33640 ( .A(n33108), .B(\modmult_1/zin[0][759] ), .Z(n26180) );
  IV U33641 ( .A(n33105), .Z(n33108) );
  XNOR U33642 ( .A(n33105), .B(n26179), .Z(n33107) );
  XOR U33643 ( .A(n33109), .B(n33110), .Z(n26179) );
  AND U33644 ( .A(\modmult_1/xin[1023] ), .B(n33111), .Z(n33110) );
  IV U33645 ( .A(n33109), .Z(n33111) );
  XOR U33646 ( .A(n33112), .B(g_input[760]), .Z(n33109) );
  NAND U33647 ( .A(n33113), .B(mul_pow), .Z(n33112) );
  XOR U33648 ( .A(g_input[760]), .B(creg[760]), .Z(n33113) );
  XOR U33649 ( .A(n33114), .B(n33115), .Z(n33105) );
  ANDN U33650 ( .A(n33116), .B(n26186), .Z(n33115) );
  XOR U33651 ( .A(n33117), .B(\modmult_1/zin[0][758] ), .Z(n26186) );
  IV U33652 ( .A(n33114), .Z(n33117) );
  XNOR U33653 ( .A(n33114), .B(n26185), .Z(n33116) );
  XOR U33654 ( .A(n33118), .B(n33119), .Z(n26185) );
  AND U33655 ( .A(\modmult_1/xin[1023] ), .B(n33120), .Z(n33119) );
  IV U33656 ( .A(n33118), .Z(n33120) );
  XOR U33657 ( .A(n33121), .B(g_input[759]), .Z(n33118) );
  NAND U33658 ( .A(n33122), .B(mul_pow), .Z(n33121) );
  XOR U33659 ( .A(g_input[759]), .B(creg[759]), .Z(n33122) );
  XOR U33660 ( .A(n33123), .B(n33124), .Z(n33114) );
  ANDN U33661 ( .A(n33125), .B(n26192), .Z(n33124) );
  XOR U33662 ( .A(n33126), .B(\modmult_1/zin[0][757] ), .Z(n26192) );
  IV U33663 ( .A(n33123), .Z(n33126) );
  XNOR U33664 ( .A(n33123), .B(n26191), .Z(n33125) );
  XOR U33665 ( .A(n33127), .B(n33128), .Z(n26191) );
  AND U33666 ( .A(\modmult_1/xin[1023] ), .B(n33129), .Z(n33128) );
  IV U33667 ( .A(n33127), .Z(n33129) );
  XOR U33668 ( .A(n33130), .B(g_input[758]), .Z(n33127) );
  NAND U33669 ( .A(n33131), .B(mul_pow), .Z(n33130) );
  XOR U33670 ( .A(g_input[758]), .B(creg[758]), .Z(n33131) );
  XOR U33671 ( .A(n33132), .B(n33133), .Z(n33123) );
  ANDN U33672 ( .A(n33134), .B(n26198), .Z(n33133) );
  XOR U33673 ( .A(n33135), .B(\modmult_1/zin[0][756] ), .Z(n26198) );
  IV U33674 ( .A(n33132), .Z(n33135) );
  XNOR U33675 ( .A(n33132), .B(n26197), .Z(n33134) );
  XOR U33676 ( .A(n33136), .B(n33137), .Z(n26197) );
  AND U33677 ( .A(\modmult_1/xin[1023] ), .B(n33138), .Z(n33137) );
  IV U33678 ( .A(n33136), .Z(n33138) );
  XOR U33679 ( .A(n33139), .B(g_input[757]), .Z(n33136) );
  NAND U33680 ( .A(n33140), .B(mul_pow), .Z(n33139) );
  XOR U33681 ( .A(g_input[757]), .B(creg[757]), .Z(n33140) );
  XOR U33682 ( .A(n33141), .B(n33142), .Z(n33132) );
  ANDN U33683 ( .A(n33143), .B(n26204), .Z(n33142) );
  XOR U33684 ( .A(n33144), .B(\modmult_1/zin[0][755] ), .Z(n26204) );
  IV U33685 ( .A(n33141), .Z(n33144) );
  XNOR U33686 ( .A(n33141), .B(n26203), .Z(n33143) );
  XOR U33687 ( .A(n33145), .B(n33146), .Z(n26203) );
  AND U33688 ( .A(\modmult_1/xin[1023] ), .B(n33147), .Z(n33146) );
  IV U33689 ( .A(n33145), .Z(n33147) );
  XOR U33690 ( .A(n33148), .B(g_input[756]), .Z(n33145) );
  NAND U33691 ( .A(n33149), .B(mul_pow), .Z(n33148) );
  XOR U33692 ( .A(g_input[756]), .B(creg[756]), .Z(n33149) );
  XOR U33693 ( .A(n33150), .B(n33151), .Z(n33141) );
  ANDN U33694 ( .A(n33152), .B(n26210), .Z(n33151) );
  XOR U33695 ( .A(n33153), .B(\modmult_1/zin[0][754] ), .Z(n26210) );
  IV U33696 ( .A(n33150), .Z(n33153) );
  XNOR U33697 ( .A(n33150), .B(n26209), .Z(n33152) );
  XOR U33698 ( .A(n33154), .B(n33155), .Z(n26209) );
  AND U33699 ( .A(\modmult_1/xin[1023] ), .B(n33156), .Z(n33155) );
  IV U33700 ( .A(n33154), .Z(n33156) );
  XOR U33701 ( .A(n33157), .B(g_input[755]), .Z(n33154) );
  NAND U33702 ( .A(n33158), .B(mul_pow), .Z(n33157) );
  XOR U33703 ( .A(g_input[755]), .B(creg[755]), .Z(n33158) );
  XOR U33704 ( .A(n33159), .B(n33160), .Z(n33150) );
  ANDN U33705 ( .A(n33161), .B(n26216), .Z(n33160) );
  XOR U33706 ( .A(n33162), .B(\modmult_1/zin[0][753] ), .Z(n26216) );
  IV U33707 ( .A(n33159), .Z(n33162) );
  XNOR U33708 ( .A(n33159), .B(n26215), .Z(n33161) );
  XOR U33709 ( .A(n33163), .B(n33164), .Z(n26215) );
  AND U33710 ( .A(\modmult_1/xin[1023] ), .B(n33165), .Z(n33164) );
  IV U33711 ( .A(n33163), .Z(n33165) );
  XOR U33712 ( .A(n33166), .B(g_input[754]), .Z(n33163) );
  NAND U33713 ( .A(n33167), .B(mul_pow), .Z(n33166) );
  XOR U33714 ( .A(g_input[754]), .B(creg[754]), .Z(n33167) );
  XOR U33715 ( .A(n33168), .B(n33169), .Z(n33159) );
  ANDN U33716 ( .A(n33170), .B(n26222), .Z(n33169) );
  XOR U33717 ( .A(n33171), .B(\modmult_1/zin[0][752] ), .Z(n26222) );
  IV U33718 ( .A(n33168), .Z(n33171) );
  XNOR U33719 ( .A(n33168), .B(n26221), .Z(n33170) );
  XOR U33720 ( .A(n33172), .B(n33173), .Z(n26221) );
  AND U33721 ( .A(\modmult_1/xin[1023] ), .B(n33174), .Z(n33173) );
  IV U33722 ( .A(n33172), .Z(n33174) );
  XOR U33723 ( .A(n33175), .B(g_input[753]), .Z(n33172) );
  NAND U33724 ( .A(n33176), .B(mul_pow), .Z(n33175) );
  XOR U33725 ( .A(g_input[753]), .B(creg[753]), .Z(n33176) );
  XOR U33726 ( .A(n33177), .B(n33178), .Z(n33168) );
  ANDN U33727 ( .A(n33179), .B(n26228), .Z(n33178) );
  XOR U33728 ( .A(n33180), .B(\modmult_1/zin[0][751] ), .Z(n26228) );
  IV U33729 ( .A(n33177), .Z(n33180) );
  XNOR U33730 ( .A(n33177), .B(n26227), .Z(n33179) );
  XOR U33731 ( .A(n33181), .B(n33182), .Z(n26227) );
  AND U33732 ( .A(\modmult_1/xin[1023] ), .B(n33183), .Z(n33182) );
  IV U33733 ( .A(n33181), .Z(n33183) );
  XOR U33734 ( .A(n33184), .B(g_input[752]), .Z(n33181) );
  NAND U33735 ( .A(n33185), .B(mul_pow), .Z(n33184) );
  XOR U33736 ( .A(g_input[752]), .B(creg[752]), .Z(n33185) );
  XOR U33737 ( .A(n33186), .B(n33187), .Z(n33177) );
  ANDN U33738 ( .A(n33188), .B(n26234), .Z(n33187) );
  XOR U33739 ( .A(n33189), .B(\modmult_1/zin[0][750] ), .Z(n26234) );
  IV U33740 ( .A(n33186), .Z(n33189) );
  XNOR U33741 ( .A(n33186), .B(n26233), .Z(n33188) );
  XOR U33742 ( .A(n33190), .B(n33191), .Z(n26233) );
  AND U33743 ( .A(\modmult_1/xin[1023] ), .B(n33192), .Z(n33191) );
  IV U33744 ( .A(n33190), .Z(n33192) );
  XOR U33745 ( .A(n33193), .B(g_input[751]), .Z(n33190) );
  NAND U33746 ( .A(n33194), .B(mul_pow), .Z(n33193) );
  XOR U33747 ( .A(g_input[751]), .B(creg[751]), .Z(n33194) );
  XOR U33748 ( .A(n33195), .B(n33196), .Z(n33186) );
  ANDN U33749 ( .A(n33197), .B(n26240), .Z(n33196) );
  XOR U33750 ( .A(n33198), .B(\modmult_1/zin[0][749] ), .Z(n26240) );
  IV U33751 ( .A(n33195), .Z(n33198) );
  XNOR U33752 ( .A(n33195), .B(n26239), .Z(n33197) );
  XOR U33753 ( .A(n33199), .B(n33200), .Z(n26239) );
  AND U33754 ( .A(\modmult_1/xin[1023] ), .B(n33201), .Z(n33200) );
  IV U33755 ( .A(n33199), .Z(n33201) );
  XOR U33756 ( .A(n33202), .B(g_input[750]), .Z(n33199) );
  NAND U33757 ( .A(n33203), .B(mul_pow), .Z(n33202) );
  XOR U33758 ( .A(g_input[750]), .B(creg[750]), .Z(n33203) );
  XOR U33759 ( .A(n33204), .B(n33205), .Z(n33195) );
  ANDN U33760 ( .A(n33206), .B(n26246), .Z(n33205) );
  XOR U33761 ( .A(n33207), .B(\modmult_1/zin[0][748] ), .Z(n26246) );
  IV U33762 ( .A(n33204), .Z(n33207) );
  XNOR U33763 ( .A(n33204), .B(n26245), .Z(n33206) );
  XOR U33764 ( .A(n33208), .B(n33209), .Z(n26245) );
  AND U33765 ( .A(\modmult_1/xin[1023] ), .B(n33210), .Z(n33209) );
  IV U33766 ( .A(n33208), .Z(n33210) );
  XOR U33767 ( .A(n33211), .B(g_input[749]), .Z(n33208) );
  NAND U33768 ( .A(n33212), .B(mul_pow), .Z(n33211) );
  XOR U33769 ( .A(g_input[749]), .B(creg[749]), .Z(n33212) );
  XOR U33770 ( .A(n33213), .B(n33214), .Z(n33204) );
  ANDN U33771 ( .A(n33215), .B(n26252), .Z(n33214) );
  XOR U33772 ( .A(n33216), .B(\modmult_1/zin[0][747] ), .Z(n26252) );
  IV U33773 ( .A(n33213), .Z(n33216) );
  XNOR U33774 ( .A(n33213), .B(n26251), .Z(n33215) );
  XOR U33775 ( .A(n33217), .B(n33218), .Z(n26251) );
  AND U33776 ( .A(\modmult_1/xin[1023] ), .B(n33219), .Z(n33218) );
  IV U33777 ( .A(n33217), .Z(n33219) );
  XOR U33778 ( .A(n33220), .B(g_input[748]), .Z(n33217) );
  NAND U33779 ( .A(n33221), .B(mul_pow), .Z(n33220) );
  XOR U33780 ( .A(g_input[748]), .B(creg[748]), .Z(n33221) );
  XOR U33781 ( .A(n33222), .B(n33223), .Z(n33213) );
  ANDN U33782 ( .A(n33224), .B(n26258), .Z(n33223) );
  XOR U33783 ( .A(n33225), .B(\modmult_1/zin[0][746] ), .Z(n26258) );
  IV U33784 ( .A(n33222), .Z(n33225) );
  XNOR U33785 ( .A(n33222), .B(n26257), .Z(n33224) );
  XOR U33786 ( .A(n33226), .B(n33227), .Z(n26257) );
  AND U33787 ( .A(\modmult_1/xin[1023] ), .B(n33228), .Z(n33227) );
  IV U33788 ( .A(n33226), .Z(n33228) );
  XOR U33789 ( .A(n33229), .B(g_input[747]), .Z(n33226) );
  NAND U33790 ( .A(n33230), .B(mul_pow), .Z(n33229) );
  XOR U33791 ( .A(g_input[747]), .B(creg[747]), .Z(n33230) );
  XOR U33792 ( .A(n33231), .B(n33232), .Z(n33222) );
  ANDN U33793 ( .A(n33233), .B(n26264), .Z(n33232) );
  XOR U33794 ( .A(n33234), .B(\modmult_1/zin[0][745] ), .Z(n26264) );
  IV U33795 ( .A(n33231), .Z(n33234) );
  XNOR U33796 ( .A(n33231), .B(n26263), .Z(n33233) );
  XOR U33797 ( .A(n33235), .B(n33236), .Z(n26263) );
  AND U33798 ( .A(\modmult_1/xin[1023] ), .B(n33237), .Z(n33236) );
  IV U33799 ( .A(n33235), .Z(n33237) );
  XOR U33800 ( .A(n33238), .B(g_input[746]), .Z(n33235) );
  NAND U33801 ( .A(n33239), .B(mul_pow), .Z(n33238) );
  XOR U33802 ( .A(g_input[746]), .B(creg[746]), .Z(n33239) );
  XOR U33803 ( .A(n33240), .B(n33241), .Z(n33231) );
  ANDN U33804 ( .A(n33242), .B(n26270), .Z(n33241) );
  XOR U33805 ( .A(n33243), .B(\modmult_1/zin[0][744] ), .Z(n26270) );
  IV U33806 ( .A(n33240), .Z(n33243) );
  XNOR U33807 ( .A(n33240), .B(n26269), .Z(n33242) );
  XOR U33808 ( .A(n33244), .B(n33245), .Z(n26269) );
  AND U33809 ( .A(\modmult_1/xin[1023] ), .B(n33246), .Z(n33245) );
  IV U33810 ( .A(n33244), .Z(n33246) );
  XOR U33811 ( .A(n33247), .B(g_input[745]), .Z(n33244) );
  NAND U33812 ( .A(n33248), .B(mul_pow), .Z(n33247) );
  XOR U33813 ( .A(g_input[745]), .B(creg[745]), .Z(n33248) );
  XOR U33814 ( .A(n33249), .B(n33250), .Z(n33240) );
  ANDN U33815 ( .A(n33251), .B(n26276), .Z(n33250) );
  XOR U33816 ( .A(n33252), .B(\modmult_1/zin[0][743] ), .Z(n26276) );
  IV U33817 ( .A(n33249), .Z(n33252) );
  XNOR U33818 ( .A(n33249), .B(n26275), .Z(n33251) );
  XOR U33819 ( .A(n33253), .B(n33254), .Z(n26275) );
  AND U33820 ( .A(\modmult_1/xin[1023] ), .B(n33255), .Z(n33254) );
  IV U33821 ( .A(n33253), .Z(n33255) );
  XOR U33822 ( .A(n33256), .B(g_input[744]), .Z(n33253) );
  NAND U33823 ( .A(n33257), .B(mul_pow), .Z(n33256) );
  XOR U33824 ( .A(g_input[744]), .B(creg[744]), .Z(n33257) );
  XOR U33825 ( .A(n33258), .B(n33259), .Z(n33249) );
  ANDN U33826 ( .A(n33260), .B(n26282), .Z(n33259) );
  XOR U33827 ( .A(n33261), .B(\modmult_1/zin[0][742] ), .Z(n26282) );
  IV U33828 ( .A(n33258), .Z(n33261) );
  XNOR U33829 ( .A(n33258), .B(n26281), .Z(n33260) );
  XOR U33830 ( .A(n33262), .B(n33263), .Z(n26281) );
  AND U33831 ( .A(\modmult_1/xin[1023] ), .B(n33264), .Z(n33263) );
  IV U33832 ( .A(n33262), .Z(n33264) );
  XOR U33833 ( .A(n33265), .B(g_input[743]), .Z(n33262) );
  NAND U33834 ( .A(n33266), .B(mul_pow), .Z(n33265) );
  XOR U33835 ( .A(g_input[743]), .B(creg[743]), .Z(n33266) );
  XOR U33836 ( .A(n33267), .B(n33268), .Z(n33258) );
  ANDN U33837 ( .A(n33269), .B(n26288), .Z(n33268) );
  XOR U33838 ( .A(n33270), .B(\modmult_1/zin[0][741] ), .Z(n26288) );
  IV U33839 ( .A(n33267), .Z(n33270) );
  XNOR U33840 ( .A(n33267), .B(n26287), .Z(n33269) );
  XOR U33841 ( .A(n33271), .B(n33272), .Z(n26287) );
  AND U33842 ( .A(\modmult_1/xin[1023] ), .B(n33273), .Z(n33272) );
  IV U33843 ( .A(n33271), .Z(n33273) );
  XOR U33844 ( .A(n33274), .B(g_input[742]), .Z(n33271) );
  NAND U33845 ( .A(n33275), .B(mul_pow), .Z(n33274) );
  XOR U33846 ( .A(g_input[742]), .B(creg[742]), .Z(n33275) );
  XOR U33847 ( .A(n33276), .B(n33277), .Z(n33267) );
  ANDN U33848 ( .A(n33278), .B(n26294), .Z(n33277) );
  XOR U33849 ( .A(n33279), .B(\modmult_1/zin[0][740] ), .Z(n26294) );
  IV U33850 ( .A(n33276), .Z(n33279) );
  XNOR U33851 ( .A(n33276), .B(n26293), .Z(n33278) );
  XOR U33852 ( .A(n33280), .B(n33281), .Z(n26293) );
  AND U33853 ( .A(\modmult_1/xin[1023] ), .B(n33282), .Z(n33281) );
  IV U33854 ( .A(n33280), .Z(n33282) );
  XOR U33855 ( .A(n33283), .B(g_input[741]), .Z(n33280) );
  NAND U33856 ( .A(n33284), .B(mul_pow), .Z(n33283) );
  XOR U33857 ( .A(g_input[741]), .B(creg[741]), .Z(n33284) );
  XOR U33858 ( .A(n33285), .B(n33286), .Z(n33276) );
  ANDN U33859 ( .A(n33287), .B(n26300), .Z(n33286) );
  XOR U33860 ( .A(n33288), .B(\modmult_1/zin[0][739] ), .Z(n26300) );
  IV U33861 ( .A(n33285), .Z(n33288) );
  XNOR U33862 ( .A(n33285), .B(n26299), .Z(n33287) );
  XOR U33863 ( .A(n33289), .B(n33290), .Z(n26299) );
  AND U33864 ( .A(\modmult_1/xin[1023] ), .B(n33291), .Z(n33290) );
  IV U33865 ( .A(n33289), .Z(n33291) );
  XOR U33866 ( .A(n33292), .B(g_input[740]), .Z(n33289) );
  NAND U33867 ( .A(n33293), .B(mul_pow), .Z(n33292) );
  XOR U33868 ( .A(g_input[740]), .B(creg[740]), .Z(n33293) );
  XOR U33869 ( .A(n33294), .B(n33295), .Z(n33285) );
  ANDN U33870 ( .A(n33296), .B(n26306), .Z(n33295) );
  XOR U33871 ( .A(n33297), .B(\modmult_1/zin[0][738] ), .Z(n26306) );
  IV U33872 ( .A(n33294), .Z(n33297) );
  XNOR U33873 ( .A(n33294), .B(n26305), .Z(n33296) );
  XOR U33874 ( .A(n33298), .B(n33299), .Z(n26305) );
  AND U33875 ( .A(\modmult_1/xin[1023] ), .B(n33300), .Z(n33299) );
  IV U33876 ( .A(n33298), .Z(n33300) );
  XOR U33877 ( .A(n33301), .B(g_input[739]), .Z(n33298) );
  NAND U33878 ( .A(n33302), .B(mul_pow), .Z(n33301) );
  XOR U33879 ( .A(g_input[739]), .B(creg[739]), .Z(n33302) );
  XOR U33880 ( .A(n33303), .B(n33304), .Z(n33294) );
  ANDN U33881 ( .A(n33305), .B(n26312), .Z(n33304) );
  XOR U33882 ( .A(n33306), .B(\modmult_1/zin[0][737] ), .Z(n26312) );
  IV U33883 ( .A(n33303), .Z(n33306) );
  XNOR U33884 ( .A(n33303), .B(n26311), .Z(n33305) );
  XOR U33885 ( .A(n33307), .B(n33308), .Z(n26311) );
  AND U33886 ( .A(\modmult_1/xin[1023] ), .B(n33309), .Z(n33308) );
  IV U33887 ( .A(n33307), .Z(n33309) );
  XOR U33888 ( .A(n33310), .B(g_input[738]), .Z(n33307) );
  NAND U33889 ( .A(n33311), .B(mul_pow), .Z(n33310) );
  XOR U33890 ( .A(g_input[738]), .B(creg[738]), .Z(n33311) );
  XOR U33891 ( .A(n33312), .B(n33313), .Z(n33303) );
  ANDN U33892 ( .A(n33314), .B(n26318), .Z(n33313) );
  XOR U33893 ( .A(n33315), .B(\modmult_1/zin[0][736] ), .Z(n26318) );
  IV U33894 ( .A(n33312), .Z(n33315) );
  XNOR U33895 ( .A(n33312), .B(n26317), .Z(n33314) );
  XOR U33896 ( .A(n33316), .B(n33317), .Z(n26317) );
  AND U33897 ( .A(\modmult_1/xin[1023] ), .B(n33318), .Z(n33317) );
  IV U33898 ( .A(n33316), .Z(n33318) );
  XOR U33899 ( .A(n33319), .B(g_input[737]), .Z(n33316) );
  NAND U33900 ( .A(n33320), .B(mul_pow), .Z(n33319) );
  XOR U33901 ( .A(g_input[737]), .B(creg[737]), .Z(n33320) );
  XOR U33902 ( .A(n33321), .B(n33322), .Z(n33312) );
  ANDN U33903 ( .A(n33323), .B(n26324), .Z(n33322) );
  XOR U33904 ( .A(n33324), .B(\modmult_1/zin[0][735] ), .Z(n26324) );
  IV U33905 ( .A(n33321), .Z(n33324) );
  XNOR U33906 ( .A(n33321), .B(n26323), .Z(n33323) );
  XOR U33907 ( .A(n33325), .B(n33326), .Z(n26323) );
  AND U33908 ( .A(\modmult_1/xin[1023] ), .B(n33327), .Z(n33326) );
  IV U33909 ( .A(n33325), .Z(n33327) );
  XOR U33910 ( .A(n33328), .B(g_input[736]), .Z(n33325) );
  NAND U33911 ( .A(n33329), .B(mul_pow), .Z(n33328) );
  XOR U33912 ( .A(g_input[736]), .B(creg[736]), .Z(n33329) );
  XOR U33913 ( .A(n33330), .B(n33331), .Z(n33321) );
  ANDN U33914 ( .A(n33332), .B(n26330), .Z(n33331) );
  XOR U33915 ( .A(n33333), .B(\modmult_1/zin[0][734] ), .Z(n26330) );
  IV U33916 ( .A(n33330), .Z(n33333) );
  XNOR U33917 ( .A(n33330), .B(n26329), .Z(n33332) );
  XOR U33918 ( .A(n33334), .B(n33335), .Z(n26329) );
  AND U33919 ( .A(\modmult_1/xin[1023] ), .B(n33336), .Z(n33335) );
  IV U33920 ( .A(n33334), .Z(n33336) );
  XOR U33921 ( .A(n33337), .B(g_input[735]), .Z(n33334) );
  NAND U33922 ( .A(n33338), .B(mul_pow), .Z(n33337) );
  XOR U33923 ( .A(g_input[735]), .B(creg[735]), .Z(n33338) );
  XOR U33924 ( .A(n33339), .B(n33340), .Z(n33330) );
  ANDN U33925 ( .A(n33341), .B(n26336), .Z(n33340) );
  XOR U33926 ( .A(n33342), .B(\modmult_1/zin[0][733] ), .Z(n26336) );
  IV U33927 ( .A(n33339), .Z(n33342) );
  XNOR U33928 ( .A(n33339), .B(n26335), .Z(n33341) );
  XOR U33929 ( .A(n33343), .B(n33344), .Z(n26335) );
  AND U33930 ( .A(\modmult_1/xin[1023] ), .B(n33345), .Z(n33344) );
  IV U33931 ( .A(n33343), .Z(n33345) );
  XOR U33932 ( .A(n33346), .B(g_input[734]), .Z(n33343) );
  NAND U33933 ( .A(n33347), .B(mul_pow), .Z(n33346) );
  XOR U33934 ( .A(g_input[734]), .B(creg[734]), .Z(n33347) );
  XOR U33935 ( .A(n33348), .B(n33349), .Z(n33339) );
  ANDN U33936 ( .A(n33350), .B(n26342), .Z(n33349) );
  XOR U33937 ( .A(n33351), .B(\modmult_1/zin[0][732] ), .Z(n26342) );
  IV U33938 ( .A(n33348), .Z(n33351) );
  XNOR U33939 ( .A(n33348), .B(n26341), .Z(n33350) );
  XOR U33940 ( .A(n33352), .B(n33353), .Z(n26341) );
  AND U33941 ( .A(\modmult_1/xin[1023] ), .B(n33354), .Z(n33353) );
  IV U33942 ( .A(n33352), .Z(n33354) );
  XOR U33943 ( .A(n33355), .B(g_input[733]), .Z(n33352) );
  NAND U33944 ( .A(n33356), .B(mul_pow), .Z(n33355) );
  XOR U33945 ( .A(g_input[733]), .B(creg[733]), .Z(n33356) );
  XOR U33946 ( .A(n33357), .B(n33358), .Z(n33348) );
  ANDN U33947 ( .A(n33359), .B(n26348), .Z(n33358) );
  XOR U33948 ( .A(n33360), .B(\modmult_1/zin[0][731] ), .Z(n26348) );
  IV U33949 ( .A(n33357), .Z(n33360) );
  XNOR U33950 ( .A(n33357), .B(n26347), .Z(n33359) );
  XOR U33951 ( .A(n33361), .B(n33362), .Z(n26347) );
  AND U33952 ( .A(\modmult_1/xin[1023] ), .B(n33363), .Z(n33362) );
  IV U33953 ( .A(n33361), .Z(n33363) );
  XOR U33954 ( .A(n33364), .B(g_input[732]), .Z(n33361) );
  NAND U33955 ( .A(n33365), .B(mul_pow), .Z(n33364) );
  XOR U33956 ( .A(g_input[732]), .B(creg[732]), .Z(n33365) );
  XOR U33957 ( .A(n33366), .B(n33367), .Z(n33357) );
  ANDN U33958 ( .A(n33368), .B(n26354), .Z(n33367) );
  XOR U33959 ( .A(n33369), .B(\modmult_1/zin[0][730] ), .Z(n26354) );
  IV U33960 ( .A(n33366), .Z(n33369) );
  XNOR U33961 ( .A(n33366), .B(n26353), .Z(n33368) );
  XOR U33962 ( .A(n33370), .B(n33371), .Z(n26353) );
  AND U33963 ( .A(\modmult_1/xin[1023] ), .B(n33372), .Z(n33371) );
  IV U33964 ( .A(n33370), .Z(n33372) );
  XOR U33965 ( .A(n33373), .B(g_input[731]), .Z(n33370) );
  NAND U33966 ( .A(n33374), .B(mul_pow), .Z(n33373) );
  XOR U33967 ( .A(g_input[731]), .B(creg[731]), .Z(n33374) );
  XOR U33968 ( .A(n33375), .B(n33376), .Z(n33366) );
  ANDN U33969 ( .A(n33377), .B(n26360), .Z(n33376) );
  XOR U33970 ( .A(n33378), .B(\modmult_1/zin[0][729] ), .Z(n26360) );
  IV U33971 ( .A(n33375), .Z(n33378) );
  XNOR U33972 ( .A(n33375), .B(n26359), .Z(n33377) );
  XOR U33973 ( .A(n33379), .B(n33380), .Z(n26359) );
  AND U33974 ( .A(\modmult_1/xin[1023] ), .B(n33381), .Z(n33380) );
  IV U33975 ( .A(n33379), .Z(n33381) );
  XOR U33976 ( .A(n33382), .B(g_input[730]), .Z(n33379) );
  NAND U33977 ( .A(n33383), .B(mul_pow), .Z(n33382) );
  XOR U33978 ( .A(g_input[730]), .B(creg[730]), .Z(n33383) );
  XOR U33979 ( .A(n33384), .B(n33385), .Z(n33375) );
  ANDN U33980 ( .A(n33386), .B(n26366), .Z(n33385) );
  XOR U33981 ( .A(n33387), .B(\modmult_1/zin[0][728] ), .Z(n26366) );
  IV U33982 ( .A(n33384), .Z(n33387) );
  XNOR U33983 ( .A(n33384), .B(n26365), .Z(n33386) );
  XOR U33984 ( .A(n33388), .B(n33389), .Z(n26365) );
  AND U33985 ( .A(\modmult_1/xin[1023] ), .B(n33390), .Z(n33389) );
  IV U33986 ( .A(n33388), .Z(n33390) );
  XOR U33987 ( .A(n33391), .B(g_input[729]), .Z(n33388) );
  NAND U33988 ( .A(n33392), .B(mul_pow), .Z(n33391) );
  XOR U33989 ( .A(g_input[729]), .B(creg[729]), .Z(n33392) );
  XOR U33990 ( .A(n33393), .B(n33394), .Z(n33384) );
  ANDN U33991 ( .A(n33395), .B(n26372), .Z(n33394) );
  XOR U33992 ( .A(n33396), .B(\modmult_1/zin[0][727] ), .Z(n26372) );
  IV U33993 ( .A(n33393), .Z(n33396) );
  XNOR U33994 ( .A(n33393), .B(n26371), .Z(n33395) );
  XOR U33995 ( .A(n33397), .B(n33398), .Z(n26371) );
  AND U33996 ( .A(\modmult_1/xin[1023] ), .B(n33399), .Z(n33398) );
  IV U33997 ( .A(n33397), .Z(n33399) );
  XOR U33998 ( .A(n33400), .B(g_input[728]), .Z(n33397) );
  NAND U33999 ( .A(n33401), .B(mul_pow), .Z(n33400) );
  XOR U34000 ( .A(g_input[728]), .B(creg[728]), .Z(n33401) );
  XOR U34001 ( .A(n33402), .B(n33403), .Z(n33393) );
  ANDN U34002 ( .A(n33404), .B(n26378), .Z(n33403) );
  XOR U34003 ( .A(n33405), .B(\modmult_1/zin[0][726] ), .Z(n26378) );
  IV U34004 ( .A(n33402), .Z(n33405) );
  XNOR U34005 ( .A(n33402), .B(n26377), .Z(n33404) );
  XOR U34006 ( .A(n33406), .B(n33407), .Z(n26377) );
  AND U34007 ( .A(\modmult_1/xin[1023] ), .B(n33408), .Z(n33407) );
  IV U34008 ( .A(n33406), .Z(n33408) );
  XOR U34009 ( .A(n33409), .B(g_input[727]), .Z(n33406) );
  NAND U34010 ( .A(n33410), .B(mul_pow), .Z(n33409) );
  XOR U34011 ( .A(g_input[727]), .B(creg[727]), .Z(n33410) );
  XOR U34012 ( .A(n33411), .B(n33412), .Z(n33402) );
  ANDN U34013 ( .A(n33413), .B(n26384), .Z(n33412) );
  XOR U34014 ( .A(n33414), .B(\modmult_1/zin[0][725] ), .Z(n26384) );
  IV U34015 ( .A(n33411), .Z(n33414) );
  XNOR U34016 ( .A(n33411), .B(n26383), .Z(n33413) );
  XOR U34017 ( .A(n33415), .B(n33416), .Z(n26383) );
  AND U34018 ( .A(\modmult_1/xin[1023] ), .B(n33417), .Z(n33416) );
  IV U34019 ( .A(n33415), .Z(n33417) );
  XOR U34020 ( .A(n33418), .B(g_input[726]), .Z(n33415) );
  NAND U34021 ( .A(n33419), .B(mul_pow), .Z(n33418) );
  XOR U34022 ( .A(g_input[726]), .B(creg[726]), .Z(n33419) );
  XOR U34023 ( .A(n33420), .B(n33421), .Z(n33411) );
  ANDN U34024 ( .A(n33422), .B(n26390), .Z(n33421) );
  XOR U34025 ( .A(n33423), .B(\modmult_1/zin[0][724] ), .Z(n26390) );
  IV U34026 ( .A(n33420), .Z(n33423) );
  XNOR U34027 ( .A(n33420), .B(n26389), .Z(n33422) );
  XOR U34028 ( .A(n33424), .B(n33425), .Z(n26389) );
  AND U34029 ( .A(\modmult_1/xin[1023] ), .B(n33426), .Z(n33425) );
  IV U34030 ( .A(n33424), .Z(n33426) );
  XOR U34031 ( .A(n33427), .B(g_input[725]), .Z(n33424) );
  NAND U34032 ( .A(n33428), .B(mul_pow), .Z(n33427) );
  XOR U34033 ( .A(g_input[725]), .B(creg[725]), .Z(n33428) );
  XOR U34034 ( .A(n33429), .B(n33430), .Z(n33420) );
  ANDN U34035 ( .A(n33431), .B(n26396), .Z(n33430) );
  XOR U34036 ( .A(n33432), .B(\modmult_1/zin[0][723] ), .Z(n26396) );
  IV U34037 ( .A(n33429), .Z(n33432) );
  XNOR U34038 ( .A(n33429), .B(n26395), .Z(n33431) );
  XOR U34039 ( .A(n33433), .B(n33434), .Z(n26395) );
  AND U34040 ( .A(\modmult_1/xin[1023] ), .B(n33435), .Z(n33434) );
  IV U34041 ( .A(n33433), .Z(n33435) );
  XOR U34042 ( .A(n33436), .B(g_input[724]), .Z(n33433) );
  NAND U34043 ( .A(n33437), .B(mul_pow), .Z(n33436) );
  XOR U34044 ( .A(g_input[724]), .B(creg[724]), .Z(n33437) );
  XOR U34045 ( .A(n33438), .B(n33439), .Z(n33429) );
  ANDN U34046 ( .A(n33440), .B(n26402), .Z(n33439) );
  XOR U34047 ( .A(n33441), .B(\modmult_1/zin[0][722] ), .Z(n26402) );
  IV U34048 ( .A(n33438), .Z(n33441) );
  XNOR U34049 ( .A(n33438), .B(n26401), .Z(n33440) );
  XOR U34050 ( .A(n33442), .B(n33443), .Z(n26401) );
  AND U34051 ( .A(\modmult_1/xin[1023] ), .B(n33444), .Z(n33443) );
  IV U34052 ( .A(n33442), .Z(n33444) );
  XOR U34053 ( .A(n33445), .B(g_input[723]), .Z(n33442) );
  NAND U34054 ( .A(n33446), .B(mul_pow), .Z(n33445) );
  XOR U34055 ( .A(g_input[723]), .B(creg[723]), .Z(n33446) );
  XOR U34056 ( .A(n33447), .B(n33448), .Z(n33438) );
  ANDN U34057 ( .A(n33449), .B(n26408), .Z(n33448) );
  XOR U34058 ( .A(n33450), .B(\modmult_1/zin[0][721] ), .Z(n26408) );
  IV U34059 ( .A(n33447), .Z(n33450) );
  XNOR U34060 ( .A(n33447), .B(n26407), .Z(n33449) );
  XOR U34061 ( .A(n33451), .B(n33452), .Z(n26407) );
  AND U34062 ( .A(\modmult_1/xin[1023] ), .B(n33453), .Z(n33452) );
  IV U34063 ( .A(n33451), .Z(n33453) );
  XOR U34064 ( .A(n33454), .B(g_input[722]), .Z(n33451) );
  NAND U34065 ( .A(n33455), .B(mul_pow), .Z(n33454) );
  XOR U34066 ( .A(g_input[722]), .B(creg[722]), .Z(n33455) );
  XOR U34067 ( .A(n33456), .B(n33457), .Z(n33447) );
  ANDN U34068 ( .A(n33458), .B(n26414), .Z(n33457) );
  XOR U34069 ( .A(n33459), .B(\modmult_1/zin[0][720] ), .Z(n26414) );
  IV U34070 ( .A(n33456), .Z(n33459) );
  XNOR U34071 ( .A(n33456), .B(n26413), .Z(n33458) );
  XOR U34072 ( .A(n33460), .B(n33461), .Z(n26413) );
  AND U34073 ( .A(\modmult_1/xin[1023] ), .B(n33462), .Z(n33461) );
  IV U34074 ( .A(n33460), .Z(n33462) );
  XOR U34075 ( .A(n33463), .B(g_input[721]), .Z(n33460) );
  NAND U34076 ( .A(n33464), .B(mul_pow), .Z(n33463) );
  XOR U34077 ( .A(g_input[721]), .B(creg[721]), .Z(n33464) );
  XOR U34078 ( .A(n33465), .B(n33466), .Z(n33456) );
  ANDN U34079 ( .A(n33467), .B(n26420), .Z(n33466) );
  XOR U34080 ( .A(n33468), .B(\modmult_1/zin[0][719] ), .Z(n26420) );
  IV U34081 ( .A(n33465), .Z(n33468) );
  XNOR U34082 ( .A(n33465), .B(n26419), .Z(n33467) );
  XOR U34083 ( .A(n33469), .B(n33470), .Z(n26419) );
  AND U34084 ( .A(\modmult_1/xin[1023] ), .B(n33471), .Z(n33470) );
  IV U34085 ( .A(n33469), .Z(n33471) );
  XOR U34086 ( .A(n33472), .B(g_input[720]), .Z(n33469) );
  NAND U34087 ( .A(n33473), .B(mul_pow), .Z(n33472) );
  XOR U34088 ( .A(g_input[720]), .B(creg[720]), .Z(n33473) );
  XOR U34089 ( .A(n33474), .B(n33475), .Z(n33465) );
  ANDN U34090 ( .A(n33476), .B(n26426), .Z(n33475) );
  XOR U34091 ( .A(n33477), .B(\modmult_1/zin[0][718] ), .Z(n26426) );
  IV U34092 ( .A(n33474), .Z(n33477) );
  XNOR U34093 ( .A(n33474), .B(n26425), .Z(n33476) );
  XOR U34094 ( .A(n33478), .B(n33479), .Z(n26425) );
  AND U34095 ( .A(\modmult_1/xin[1023] ), .B(n33480), .Z(n33479) );
  IV U34096 ( .A(n33478), .Z(n33480) );
  XOR U34097 ( .A(n33481), .B(g_input[719]), .Z(n33478) );
  NAND U34098 ( .A(n33482), .B(mul_pow), .Z(n33481) );
  XOR U34099 ( .A(g_input[719]), .B(creg[719]), .Z(n33482) );
  XOR U34100 ( .A(n33483), .B(n33484), .Z(n33474) );
  ANDN U34101 ( .A(n33485), .B(n26432), .Z(n33484) );
  XOR U34102 ( .A(n33486), .B(\modmult_1/zin[0][717] ), .Z(n26432) );
  IV U34103 ( .A(n33483), .Z(n33486) );
  XNOR U34104 ( .A(n33483), .B(n26431), .Z(n33485) );
  XOR U34105 ( .A(n33487), .B(n33488), .Z(n26431) );
  AND U34106 ( .A(\modmult_1/xin[1023] ), .B(n33489), .Z(n33488) );
  IV U34107 ( .A(n33487), .Z(n33489) );
  XOR U34108 ( .A(n33490), .B(g_input[718]), .Z(n33487) );
  NAND U34109 ( .A(n33491), .B(mul_pow), .Z(n33490) );
  XOR U34110 ( .A(g_input[718]), .B(creg[718]), .Z(n33491) );
  XOR U34111 ( .A(n33492), .B(n33493), .Z(n33483) );
  ANDN U34112 ( .A(n33494), .B(n26438), .Z(n33493) );
  XOR U34113 ( .A(n33495), .B(\modmult_1/zin[0][716] ), .Z(n26438) );
  IV U34114 ( .A(n33492), .Z(n33495) );
  XNOR U34115 ( .A(n33492), .B(n26437), .Z(n33494) );
  XOR U34116 ( .A(n33496), .B(n33497), .Z(n26437) );
  AND U34117 ( .A(\modmult_1/xin[1023] ), .B(n33498), .Z(n33497) );
  IV U34118 ( .A(n33496), .Z(n33498) );
  XOR U34119 ( .A(n33499), .B(g_input[717]), .Z(n33496) );
  NAND U34120 ( .A(n33500), .B(mul_pow), .Z(n33499) );
  XOR U34121 ( .A(g_input[717]), .B(creg[717]), .Z(n33500) );
  XOR U34122 ( .A(n33501), .B(n33502), .Z(n33492) );
  ANDN U34123 ( .A(n33503), .B(n26444), .Z(n33502) );
  XOR U34124 ( .A(n33504), .B(\modmult_1/zin[0][715] ), .Z(n26444) );
  IV U34125 ( .A(n33501), .Z(n33504) );
  XNOR U34126 ( .A(n33501), .B(n26443), .Z(n33503) );
  XOR U34127 ( .A(n33505), .B(n33506), .Z(n26443) );
  AND U34128 ( .A(\modmult_1/xin[1023] ), .B(n33507), .Z(n33506) );
  IV U34129 ( .A(n33505), .Z(n33507) );
  XOR U34130 ( .A(n33508), .B(g_input[716]), .Z(n33505) );
  NAND U34131 ( .A(n33509), .B(mul_pow), .Z(n33508) );
  XOR U34132 ( .A(g_input[716]), .B(creg[716]), .Z(n33509) );
  XOR U34133 ( .A(n33510), .B(n33511), .Z(n33501) );
  ANDN U34134 ( .A(n33512), .B(n26450), .Z(n33511) );
  XOR U34135 ( .A(n33513), .B(\modmult_1/zin[0][714] ), .Z(n26450) );
  IV U34136 ( .A(n33510), .Z(n33513) );
  XNOR U34137 ( .A(n33510), .B(n26449), .Z(n33512) );
  XOR U34138 ( .A(n33514), .B(n33515), .Z(n26449) );
  AND U34139 ( .A(\modmult_1/xin[1023] ), .B(n33516), .Z(n33515) );
  IV U34140 ( .A(n33514), .Z(n33516) );
  XOR U34141 ( .A(n33517), .B(g_input[715]), .Z(n33514) );
  NAND U34142 ( .A(n33518), .B(mul_pow), .Z(n33517) );
  XOR U34143 ( .A(g_input[715]), .B(creg[715]), .Z(n33518) );
  XOR U34144 ( .A(n33519), .B(n33520), .Z(n33510) );
  ANDN U34145 ( .A(n33521), .B(n26456), .Z(n33520) );
  XOR U34146 ( .A(n33522), .B(\modmult_1/zin[0][713] ), .Z(n26456) );
  IV U34147 ( .A(n33519), .Z(n33522) );
  XNOR U34148 ( .A(n33519), .B(n26455), .Z(n33521) );
  XOR U34149 ( .A(n33523), .B(n33524), .Z(n26455) );
  AND U34150 ( .A(\modmult_1/xin[1023] ), .B(n33525), .Z(n33524) );
  IV U34151 ( .A(n33523), .Z(n33525) );
  XOR U34152 ( .A(n33526), .B(g_input[714]), .Z(n33523) );
  NAND U34153 ( .A(n33527), .B(mul_pow), .Z(n33526) );
  XOR U34154 ( .A(g_input[714]), .B(creg[714]), .Z(n33527) );
  XOR U34155 ( .A(n33528), .B(n33529), .Z(n33519) );
  ANDN U34156 ( .A(n33530), .B(n26462), .Z(n33529) );
  XOR U34157 ( .A(n33531), .B(\modmult_1/zin[0][712] ), .Z(n26462) );
  IV U34158 ( .A(n33528), .Z(n33531) );
  XNOR U34159 ( .A(n33528), .B(n26461), .Z(n33530) );
  XOR U34160 ( .A(n33532), .B(n33533), .Z(n26461) );
  AND U34161 ( .A(\modmult_1/xin[1023] ), .B(n33534), .Z(n33533) );
  IV U34162 ( .A(n33532), .Z(n33534) );
  XOR U34163 ( .A(n33535), .B(g_input[713]), .Z(n33532) );
  NAND U34164 ( .A(n33536), .B(mul_pow), .Z(n33535) );
  XOR U34165 ( .A(g_input[713]), .B(creg[713]), .Z(n33536) );
  XOR U34166 ( .A(n33537), .B(n33538), .Z(n33528) );
  ANDN U34167 ( .A(n33539), .B(n26468), .Z(n33538) );
  XOR U34168 ( .A(n33540), .B(\modmult_1/zin[0][711] ), .Z(n26468) );
  IV U34169 ( .A(n33537), .Z(n33540) );
  XNOR U34170 ( .A(n33537), .B(n26467), .Z(n33539) );
  XOR U34171 ( .A(n33541), .B(n33542), .Z(n26467) );
  AND U34172 ( .A(\modmult_1/xin[1023] ), .B(n33543), .Z(n33542) );
  IV U34173 ( .A(n33541), .Z(n33543) );
  XOR U34174 ( .A(n33544), .B(g_input[712]), .Z(n33541) );
  NAND U34175 ( .A(n33545), .B(mul_pow), .Z(n33544) );
  XOR U34176 ( .A(g_input[712]), .B(creg[712]), .Z(n33545) );
  XOR U34177 ( .A(n33546), .B(n33547), .Z(n33537) );
  ANDN U34178 ( .A(n33548), .B(n26474), .Z(n33547) );
  XOR U34179 ( .A(n33549), .B(\modmult_1/zin[0][710] ), .Z(n26474) );
  IV U34180 ( .A(n33546), .Z(n33549) );
  XNOR U34181 ( .A(n33546), .B(n26473), .Z(n33548) );
  XOR U34182 ( .A(n33550), .B(n33551), .Z(n26473) );
  AND U34183 ( .A(\modmult_1/xin[1023] ), .B(n33552), .Z(n33551) );
  IV U34184 ( .A(n33550), .Z(n33552) );
  XOR U34185 ( .A(n33553), .B(g_input[711]), .Z(n33550) );
  NAND U34186 ( .A(n33554), .B(mul_pow), .Z(n33553) );
  XOR U34187 ( .A(g_input[711]), .B(creg[711]), .Z(n33554) );
  XOR U34188 ( .A(n33555), .B(n33556), .Z(n33546) );
  ANDN U34189 ( .A(n33557), .B(n26480), .Z(n33556) );
  XOR U34190 ( .A(n33558), .B(\modmult_1/zin[0][709] ), .Z(n26480) );
  IV U34191 ( .A(n33555), .Z(n33558) );
  XNOR U34192 ( .A(n33555), .B(n26479), .Z(n33557) );
  XOR U34193 ( .A(n33559), .B(n33560), .Z(n26479) );
  AND U34194 ( .A(\modmult_1/xin[1023] ), .B(n33561), .Z(n33560) );
  IV U34195 ( .A(n33559), .Z(n33561) );
  XOR U34196 ( .A(n33562), .B(g_input[710]), .Z(n33559) );
  NAND U34197 ( .A(n33563), .B(mul_pow), .Z(n33562) );
  XOR U34198 ( .A(g_input[710]), .B(creg[710]), .Z(n33563) );
  XOR U34199 ( .A(n33564), .B(n33565), .Z(n33555) );
  ANDN U34200 ( .A(n33566), .B(n26486), .Z(n33565) );
  XOR U34201 ( .A(n33567), .B(\modmult_1/zin[0][708] ), .Z(n26486) );
  IV U34202 ( .A(n33564), .Z(n33567) );
  XNOR U34203 ( .A(n33564), .B(n26485), .Z(n33566) );
  XOR U34204 ( .A(n33568), .B(n33569), .Z(n26485) );
  AND U34205 ( .A(\modmult_1/xin[1023] ), .B(n33570), .Z(n33569) );
  IV U34206 ( .A(n33568), .Z(n33570) );
  XOR U34207 ( .A(n33571), .B(g_input[709]), .Z(n33568) );
  NAND U34208 ( .A(n33572), .B(mul_pow), .Z(n33571) );
  XOR U34209 ( .A(g_input[709]), .B(creg[709]), .Z(n33572) );
  XOR U34210 ( .A(n33573), .B(n33574), .Z(n33564) );
  ANDN U34211 ( .A(n33575), .B(n26492), .Z(n33574) );
  XOR U34212 ( .A(n33576), .B(\modmult_1/zin[0][707] ), .Z(n26492) );
  IV U34213 ( .A(n33573), .Z(n33576) );
  XNOR U34214 ( .A(n33573), .B(n26491), .Z(n33575) );
  XOR U34215 ( .A(n33577), .B(n33578), .Z(n26491) );
  AND U34216 ( .A(\modmult_1/xin[1023] ), .B(n33579), .Z(n33578) );
  IV U34217 ( .A(n33577), .Z(n33579) );
  XOR U34218 ( .A(n33580), .B(g_input[708]), .Z(n33577) );
  NAND U34219 ( .A(n33581), .B(mul_pow), .Z(n33580) );
  XOR U34220 ( .A(g_input[708]), .B(creg[708]), .Z(n33581) );
  XOR U34221 ( .A(n33582), .B(n33583), .Z(n33573) );
  ANDN U34222 ( .A(n33584), .B(n26498), .Z(n33583) );
  XOR U34223 ( .A(n33585), .B(\modmult_1/zin[0][706] ), .Z(n26498) );
  IV U34224 ( .A(n33582), .Z(n33585) );
  XNOR U34225 ( .A(n33582), .B(n26497), .Z(n33584) );
  XOR U34226 ( .A(n33586), .B(n33587), .Z(n26497) );
  AND U34227 ( .A(\modmult_1/xin[1023] ), .B(n33588), .Z(n33587) );
  IV U34228 ( .A(n33586), .Z(n33588) );
  XOR U34229 ( .A(n33589), .B(g_input[707]), .Z(n33586) );
  NAND U34230 ( .A(n33590), .B(mul_pow), .Z(n33589) );
  XOR U34231 ( .A(g_input[707]), .B(creg[707]), .Z(n33590) );
  XOR U34232 ( .A(n33591), .B(n33592), .Z(n33582) );
  ANDN U34233 ( .A(n33593), .B(n26504), .Z(n33592) );
  XOR U34234 ( .A(n33594), .B(\modmult_1/zin[0][705] ), .Z(n26504) );
  IV U34235 ( .A(n33591), .Z(n33594) );
  XNOR U34236 ( .A(n33591), .B(n26503), .Z(n33593) );
  XOR U34237 ( .A(n33595), .B(n33596), .Z(n26503) );
  AND U34238 ( .A(\modmult_1/xin[1023] ), .B(n33597), .Z(n33596) );
  IV U34239 ( .A(n33595), .Z(n33597) );
  XOR U34240 ( .A(n33598), .B(g_input[706]), .Z(n33595) );
  NAND U34241 ( .A(n33599), .B(mul_pow), .Z(n33598) );
  XOR U34242 ( .A(g_input[706]), .B(creg[706]), .Z(n33599) );
  XOR U34243 ( .A(n33600), .B(n33601), .Z(n33591) );
  ANDN U34244 ( .A(n33602), .B(n26510), .Z(n33601) );
  XOR U34245 ( .A(n33603), .B(\modmult_1/zin[0][704] ), .Z(n26510) );
  IV U34246 ( .A(n33600), .Z(n33603) );
  XNOR U34247 ( .A(n33600), .B(n26509), .Z(n33602) );
  XOR U34248 ( .A(n33604), .B(n33605), .Z(n26509) );
  AND U34249 ( .A(\modmult_1/xin[1023] ), .B(n33606), .Z(n33605) );
  IV U34250 ( .A(n33604), .Z(n33606) );
  XOR U34251 ( .A(n33607), .B(g_input[705]), .Z(n33604) );
  NAND U34252 ( .A(n33608), .B(mul_pow), .Z(n33607) );
  XOR U34253 ( .A(g_input[705]), .B(creg[705]), .Z(n33608) );
  XOR U34254 ( .A(n33609), .B(n33610), .Z(n33600) );
  ANDN U34255 ( .A(n33611), .B(n26516), .Z(n33610) );
  XOR U34256 ( .A(n33612), .B(\modmult_1/zin[0][703] ), .Z(n26516) );
  IV U34257 ( .A(n33609), .Z(n33612) );
  XNOR U34258 ( .A(n33609), .B(n26515), .Z(n33611) );
  XOR U34259 ( .A(n33613), .B(n33614), .Z(n26515) );
  AND U34260 ( .A(\modmult_1/xin[1023] ), .B(n33615), .Z(n33614) );
  IV U34261 ( .A(n33613), .Z(n33615) );
  XOR U34262 ( .A(n33616), .B(g_input[704]), .Z(n33613) );
  NAND U34263 ( .A(n33617), .B(mul_pow), .Z(n33616) );
  XOR U34264 ( .A(g_input[704]), .B(creg[704]), .Z(n33617) );
  XOR U34265 ( .A(n33618), .B(n33619), .Z(n33609) );
  ANDN U34266 ( .A(n33620), .B(n26522), .Z(n33619) );
  XOR U34267 ( .A(n33621), .B(\modmult_1/zin[0][702] ), .Z(n26522) );
  IV U34268 ( .A(n33618), .Z(n33621) );
  XNOR U34269 ( .A(n33618), .B(n26521), .Z(n33620) );
  XOR U34270 ( .A(n33622), .B(n33623), .Z(n26521) );
  AND U34271 ( .A(\modmult_1/xin[1023] ), .B(n33624), .Z(n33623) );
  IV U34272 ( .A(n33622), .Z(n33624) );
  XOR U34273 ( .A(n33625), .B(g_input[703]), .Z(n33622) );
  NAND U34274 ( .A(n33626), .B(mul_pow), .Z(n33625) );
  XOR U34275 ( .A(g_input[703]), .B(creg[703]), .Z(n33626) );
  XOR U34276 ( .A(n33627), .B(n33628), .Z(n33618) );
  ANDN U34277 ( .A(n33629), .B(n26528), .Z(n33628) );
  XOR U34278 ( .A(n33630), .B(\modmult_1/zin[0][701] ), .Z(n26528) );
  IV U34279 ( .A(n33627), .Z(n33630) );
  XNOR U34280 ( .A(n33627), .B(n26527), .Z(n33629) );
  XOR U34281 ( .A(n33631), .B(n33632), .Z(n26527) );
  AND U34282 ( .A(\modmult_1/xin[1023] ), .B(n33633), .Z(n33632) );
  IV U34283 ( .A(n33631), .Z(n33633) );
  XOR U34284 ( .A(n33634), .B(g_input[702]), .Z(n33631) );
  NAND U34285 ( .A(n33635), .B(mul_pow), .Z(n33634) );
  XOR U34286 ( .A(g_input[702]), .B(creg[702]), .Z(n33635) );
  XOR U34287 ( .A(n33636), .B(n33637), .Z(n33627) );
  ANDN U34288 ( .A(n33638), .B(n26534), .Z(n33637) );
  XOR U34289 ( .A(n33639), .B(\modmult_1/zin[0][700] ), .Z(n26534) );
  IV U34290 ( .A(n33636), .Z(n33639) );
  XNOR U34291 ( .A(n33636), .B(n26533), .Z(n33638) );
  XOR U34292 ( .A(n33640), .B(n33641), .Z(n26533) );
  AND U34293 ( .A(\modmult_1/xin[1023] ), .B(n33642), .Z(n33641) );
  IV U34294 ( .A(n33640), .Z(n33642) );
  XOR U34295 ( .A(n33643), .B(g_input[701]), .Z(n33640) );
  NAND U34296 ( .A(n33644), .B(mul_pow), .Z(n33643) );
  XOR U34297 ( .A(g_input[701]), .B(creg[701]), .Z(n33644) );
  XOR U34298 ( .A(n33645), .B(n33646), .Z(n33636) );
  ANDN U34299 ( .A(n33647), .B(n26540), .Z(n33646) );
  XOR U34300 ( .A(n33648), .B(\modmult_1/zin[0][699] ), .Z(n26540) );
  IV U34301 ( .A(n33645), .Z(n33648) );
  XNOR U34302 ( .A(n33645), .B(n26539), .Z(n33647) );
  XOR U34303 ( .A(n33649), .B(n33650), .Z(n26539) );
  AND U34304 ( .A(\modmult_1/xin[1023] ), .B(n33651), .Z(n33650) );
  IV U34305 ( .A(n33649), .Z(n33651) );
  XOR U34306 ( .A(n33652), .B(g_input[700]), .Z(n33649) );
  NAND U34307 ( .A(n33653), .B(mul_pow), .Z(n33652) );
  XOR U34308 ( .A(g_input[700]), .B(creg[700]), .Z(n33653) );
  XOR U34309 ( .A(n33654), .B(n33655), .Z(n33645) );
  ANDN U34310 ( .A(n33656), .B(n26546), .Z(n33655) );
  XOR U34311 ( .A(n33657), .B(\modmult_1/zin[0][698] ), .Z(n26546) );
  IV U34312 ( .A(n33654), .Z(n33657) );
  XNOR U34313 ( .A(n33654), .B(n26545), .Z(n33656) );
  XOR U34314 ( .A(n33658), .B(n33659), .Z(n26545) );
  AND U34315 ( .A(\modmult_1/xin[1023] ), .B(n33660), .Z(n33659) );
  IV U34316 ( .A(n33658), .Z(n33660) );
  XOR U34317 ( .A(n33661), .B(g_input[699]), .Z(n33658) );
  NAND U34318 ( .A(n33662), .B(mul_pow), .Z(n33661) );
  XOR U34319 ( .A(g_input[699]), .B(creg[699]), .Z(n33662) );
  XOR U34320 ( .A(n33663), .B(n33664), .Z(n33654) );
  ANDN U34321 ( .A(n33665), .B(n26552), .Z(n33664) );
  XOR U34322 ( .A(n33666), .B(\modmult_1/zin[0][697] ), .Z(n26552) );
  IV U34323 ( .A(n33663), .Z(n33666) );
  XNOR U34324 ( .A(n33663), .B(n26551), .Z(n33665) );
  XOR U34325 ( .A(n33667), .B(n33668), .Z(n26551) );
  AND U34326 ( .A(\modmult_1/xin[1023] ), .B(n33669), .Z(n33668) );
  IV U34327 ( .A(n33667), .Z(n33669) );
  XOR U34328 ( .A(n33670), .B(g_input[698]), .Z(n33667) );
  NAND U34329 ( .A(n33671), .B(mul_pow), .Z(n33670) );
  XOR U34330 ( .A(g_input[698]), .B(creg[698]), .Z(n33671) );
  XOR U34331 ( .A(n33672), .B(n33673), .Z(n33663) );
  ANDN U34332 ( .A(n33674), .B(n26558), .Z(n33673) );
  XOR U34333 ( .A(n33675), .B(\modmult_1/zin[0][696] ), .Z(n26558) );
  IV U34334 ( .A(n33672), .Z(n33675) );
  XNOR U34335 ( .A(n33672), .B(n26557), .Z(n33674) );
  XOR U34336 ( .A(n33676), .B(n33677), .Z(n26557) );
  AND U34337 ( .A(\modmult_1/xin[1023] ), .B(n33678), .Z(n33677) );
  IV U34338 ( .A(n33676), .Z(n33678) );
  XOR U34339 ( .A(n33679), .B(g_input[697]), .Z(n33676) );
  NAND U34340 ( .A(n33680), .B(mul_pow), .Z(n33679) );
  XOR U34341 ( .A(g_input[697]), .B(creg[697]), .Z(n33680) );
  XOR U34342 ( .A(n33681), .B(n33682), .Z(n33672) );
  ANDN U34343 ( .A(n33683), .B(n26564), .Z(n33682) );
  XOR U34344 ( .A(n33684), .B(\modmult_1/zin[0][695] ), .Z(n26564) );
  IV U34345 ( .A(n33681), .Z(n33684) );
  XNOR U34346 ( .A(n33681), .B(n26563), .Z(n33683) );
  XOR U34347 ( .A(n33685), .B(n33686), .Z(n26563) );
  AND U34348 ( .A(\modmult_1/xin[1023] ), .B(n33687), .Z(n33686) );
  IV U34349 ( .A(n33685), .Z(n33687) );
  XOR U34350 ( .A(n33688), .B(g_input[696]), .Z(n33685) );
  NAND U34351 ( .A(n33689), .B(mul_pow), .Z(n33688) );
  XOR U34352 ( .A(g_input[696]), .B(creg[696]), .Z(n33689) );
  XOR U34353 ( .A(n33690), .B(n33691), .Z(n33681) );
  ANDN U34354 ( .A(n33692), .B(n26570), .Z(n33691) );
  XOR U34355 ( .A(n33693), .B(\modmult_1/zin[0][694] ), .Z(n26570) );
  IV U34356 ( .A(n33690), .Z(n33693) );
  XNOR U34357 ( .A(n33690), .B(n26569), .Z(n33692) );
  XOR U34358 ( .A(n33694), .B(n33695), .Z(n26569) );
  AND U34359 ( .A(\modmult_1/xin[1023] ), .B(n33696), .Z(n33695) );
  IV U34360 ( .A(n33694), .Z(n33696) );
  XOR U34361 ( .A(n33697), .B(g_input[695]), .Z(n33694) );
  NAND U34362 ( .A(n33698), .B(mul_pow), .Z(n33697) );
  XOR U34363 ( .A(g_input[695]), .B(creg[695]), .Z(n33698) );
  XOR U34364 ( .A(n33699), .B(n33700), .Z(n33690) );
  ANDN U34365 ( .A(n33701), .B(n26576), .Z(n33700) );
  XOR U34366 ( .A(n33702), .B(\modmult_1/zin[0][693] ), .Z(n26576) );
  IV U34367 ( .A(n33699), .Z(n33702) );
  XNOR U34368 ( .A(n33699), .B(n26575), .Z(n33701) );
  XOR U34369 ( .A(n33703), .B(n33704), .Z(n26575) );
  AND U34370 ( .A(\modmult_1/xin[1023] ), .B(n33705), .Z(n33704) );
  IV U34371 ( .A(n33703), .Z(n33705) );
  XOR U34372 ( .A(n33706), .B(g_input[694]), .Z(n33703) );
  NAND U34373 ( .A(n33707), .B(mul_pow), .Z(n33706) );
  XOR U34374 ( .A(g_input[694]), .B(creg[694]), .Z(n33707) );
  XOR U34375 ( .A(n33708), .B(n33709), .Z(n33699) );
  ANDN U34376 ( .A(n33710), .B(n26582), .Z(n33709) );
  XOR U34377 ( .A(n33711), .B(\modmult_1/zin[0][692] ), .Z(n26582) );
  IV U34378 ( .A(n33708), .Z(n33711) );
  XNOR U34379 ( .A(n33708), .B(n26581), .Z(n33710) );
  XOR U34380 ( .A(n33712), .B(n33713), .Z(n26581) );
  AND U34381 ( .A(\modmult_1/xin[1023] ), .B(n33714), .Z(n33713) );
  IV U34382 ( .A(n33712), .Z(n33714) );
  XOR U34383 ( .A(n33715), .B(g_input[693]), .Z(n33712) );
  NAND U34384 ( .A(n33716), .B(mul_pow), .Z(n33715) );
  XOR U34385 ( .A(g_input[693]), .B(creg[693]), .Z(n33716) );
  XOR U34386 ( .A(n33717), .B(n33718), .Z(n33708) );
  ANDN U34387 ( .A(n33719), .B(n26588), .Z(n33718) );
  XOR U34388 ( .A(n33720), .B(\modmult_1/zin[0][691] ), .Z(n26588) );
  IV U34389 ( .A(n33717), .Z(n33720) );
  XNOR U34390 ( .A(n33717), .B(n26587), .Z(n33719) );
  XOR U34391 ( .A(n33721), .B(n33722), .Z(n26587) );
  AND U34392 ( .A(\modmult_1/xin[1023] ), .B(n33723), .Z(n33722) );
  IV U34393 ( .A(n33721), .Z(n33723) );
  XOR U34394 ( .A(n33724), .B(g_input[692]), .Z(n33721) );
  NAND U34395 ( .A(n33725), .B(mul_pow), .Z(n33724) );
  XOR U34396 ( .A(g_input[692]), .B(creg[692]), .Z(n33725) );
  XOR U34397 ( .A(n33726), .B(n33727), .Z(n33717) );
  ANDN U34398 ( .A(n33728), .B(n26594), .Z(n33727) );
  XOR U34399 ( .A(n33729), .B(\modmult_1/zin[0][690] ), .Z(n26594) );
  IV U34400 ( .A(n33726), .Z(n33729) );
  XNOR U34401 ( .A(n33726), .B(n26593), .Z(n33728) );
  XOR U34402 ( .A(n33730), .B(n33731), .Z(n26593) );
  AND U34403 ( .A(\modmult_1/xin[1023] ), .B(n33732), .Z(n33731) );
  IV U34404 ( .A(n33730), .Z(n33732) );
  XOR U34405 ( .A(n33733), .B(g_input[691]), .Z(n33730) );
  NAND U34406 ( .A(n33734), .B(mul_pow), .Z(n33733) );
  XOR U34407 ( .A(g_input[691]), .B(creg[691]), .Z(n33734) );
  XOR U34408 ( .A(n33735), .B(n33736), .Z(n33726) );
  ANDN U34409 ( .A(n33737), .B(n26600), .Z(n33736) );
  XOR U34410 ( .A(n33738), .B(\modmult_1/zin[0][689] ), .Z(n26600) );
  IV U34411 ( .A(n33735), .Z(n33738) );
  XNOR U34412 ( .A(n33735), .B(n26599), .Z(n33737) );
  XOR U34413 ( .A(n33739), .B(n33740), .Z(n26599) );
  AND U34414 ( .A(\modmult_1/xin[1023] ), .B(n33741), .Z(n33740) );
  IV U34415 ( .A(n33739), .Z(n33741) );
  XOR U34416 ( .A(n33742), .B(g_input[690]), .Z(n33739) );
  NAND U34417 ( .A(n33743), .B(mul_pow), .Z(n33742) );
  XOR U34418 ( .A(g_input[690]), .B(creg[690]), .Z(n33743) );
  XOR U34419 ( .A(n33744), .B(n33745), .Z(n33735) );
  ANDN U34420 ( .A(n33746), .B(n26606), .Z(n33745) );
  XOR U34421 ( .A(n33747), .B(\modmult_1/zin[0][688] ), .Z(n26606) );
  IV U34422 ( .A(n33744), .Z(n33747) );
  XNOR U34423 ( .A(n33744), .B(n26605), .Z(n33746) );
  XOR U34424 ( .A(n33748), .B(n33749), .Z(n26605) );
  AND U34425 ( .A(\modmult_1/xin[1023] ), .B(n33750), .Z(n33749) );
  IV U34426 ( .A(n33748), .Z(n33750) );
  XOR U34427 ( .A(n33751), .B(g_input[689]), .Z(n33748) );
  NAND U34428 ( .A(n33752), .B(mul_pow), .Z(n33751) );
  XOR U34429 ( .A(g_input[689]), .B(creg[689]), .Z(n33752) );
  XOR U34430 ( .A(n33753), .B(n33754), .Z(n33744) );
  ANDN U34431 ( .A(n33755), .B(n26612), .Z(n33754) );
  XOR U34432 ( .A(n33756), .B(\modmult_1/zin[0][687] ), .Z(n26612) );
  IV U34433 ( .A(n33753), .Z(n33756) );
  XNOR U34434 ( .A(n33753), .B(n26611), .Z(n33755) );
  XOR U34435 ( .A(n33757), .B(n33758), .Z(n26611) );
  AND U34436 ( .A(\modmult_1/xin[1023] ), .B(n33759), .Z(n33758) );
  IV U34437 ( .A(n33757), .Z(n33759) );
  XOR U34438 ( .A(n33760), .B(g_input[688]), .Z(n33757) );
  NAND U34439 ( .A(n33761), .B(mul_pow), .Z(n33760) );
  XOR U34440 ( .A(g_input[688]), .B(creg[688]), .Z(n33761) );
  XOR U34441 ( .A(n33762), .B(n33763), .Z(n33753) );
  ANDN U34442 ( .A(n33764), .B(n26618), .Z(n33763) );
  XOR U34443 ( .A(n33765), .B(\modmult_1/zin[0][686] ), .Z(n26618) );
  IV U34444 ( .A(n33762), .Z(n33765) );
  XNOR U34445 ( .A(n33762), .B(n26617), .Z(n33764) );
  XOR U34446 ( .A(n33766), .B(n33767), .Z(n26617) );
  AND U34447 ( .A(\modmult_1/xin[1023] ), .B(n33768), .Z(n33767) );
  IV U34448 ( .A(n33766), .Z(n33768) );
  XOR U34449 ( .A(n33769), .B(g_input[687]), .Z(n33766) );
  NAND U34450 ( .A(n33770), .B(mul_pow), .Z(n33769) );
  XOR U34451 ( .A(g_input[687]), .B(creg[687]), .Z(n33770) );
  XOR U34452 ( .A(n33771), .B(n33772), .Z(n33762) );
  ANDN U34453 ( .A(n33773), .B(n26624), .Z(n33772) );
  XOR U34454 ( .A(n33774), .B(\modmult_1/zin[0][685] ), .Z(n26624) );
  IV U34455 ( .A(n33771), .Z(n33774) );
  XNOR U34456 ( .A(n33771), .B(n26623), .Z(n33773) );
  XOR U34457 ( .A(n33775), .B(n33776), .Z(n26623) );
  AND U34458 ( .A(\modmult_1/xin[1023] ), .B(n33777), .Z(n33776) );
  IV U34459 ( .A(n33775), .Z(n33777) );
  XOR U34460 ( .A(n33778), .B(g_input[686]), .Z(n33775) );
  NAND U34461 ( .A(n33779), .B(mul_pow), .Z(n33778) );
  XOR U34462 ( .A(g_input[686]), .B(creg[686]), .Z(n33779) );
  XOR U34463 ( .A(n33780), .B(n33781), .Z(n33771) );
  ANDN U34464 ( .A(n33782), .B(n26630), .Z(n33781) );
  XOR U34465 ( .A(n33783), .B(\modmult_1/zin[0][684] ), .Z(n26630) );
  IV U34466 ( .A(n33780), .Z(n33783) );
  XNOR U34467 ( .A(n33780), .B(n26629), .Z(n33782) );
  XOR U34468 ( .A(n33784), .B(n33785), .Z(n26629) );
  AND U34469 ( .A(\modmult_1/xin[1023] ), .B(n33786), .Z(n33785) );
  IV U34470 ( .A(n33784), .Z(n33786) );
  XOR U34471 ( .A(n33787), .B(g_input[685]), .Z(n33784) );
  NAND U34472 ( .A(n33788), .B(mul_pow), .Z(n33787) );
  XOR U34473 ( .A(g_input[685]), .B(creg[685]), .Z(n33788) );
  XOR U34474 ( .A(n33789), .B(n33790), .Z(n33780) );
  ANDN U34475 ( .A(n33791), .B(n26636), .Z(n33790) );
  XOR U34476 ( .A(n33792), .B(\modmult_1/zin[0][683] ), .Z(n26636) );
  IV U34477 ( .A(n33789), .Z(n33792) );
  XNOR U34478 ( .A(n33789), .B(n26635), .Z(n33791) );
  XOR U34479 ( .A(n33793), .B(n33794), .Z(n26635) );
  AND U34480 ( .A(\modmult_1/xin[1023] ), .B(n33795), .Z(n33794) );
  IV U34481 ( .A(n33793), .Z(n33795) );
  XOR U34482 ( .A(n33796), .B(g_input[684]), .Z(n33793) );
  NAND U34483 ( .A(n33797), .B(mul_pow), .Z(n33796) );
  XOR U34484 ( .A(g_input[684]), .B(creg[684]), .Z(n33797) );
  XOR U34485 ( .A(n33798), .B(n33799), .Z(n33789) );
  ANDN U34486 ( .A(n33800), .B(n26642), .Z(n33799) );
  XOR U34487 ( .A(n33801), .B(\modmult_1/zin[0][682] ), .Z(n26642) );
  IV U34488 ( .A(n33798), .Z(n33801) );
  XNOR U34489 ( .A(n33798), .B(n26641), .Z(n33800) );
  XOR U34490 ( .A(n33802), .B(n33803), .Z(n26641) );
  AND U34491 ( .A(\modmult_1/xin[1023] ), .B(n33804), .Z(n33803) );
  IV U34492 ( .A(n33802), .Z(n33804) );
  XOR U34493 ( .A(n33805), .B(g_input[683]), .Z(n33802) );
  NAND U34494 ( .A(n33806), .B(mul_pow), .Z(n33805) );
  XOR U34495 ( .A(g_input[683]), .B(creg[683]), .Z(n33806) );
  XOR U34496 ( .A(n33807), .B(n33808), .Z(n33798) );
  ANDN U34497 ( .A(n33809), .B(n26648), .Z(n33808) );
  XOR U34498 ( .A(n33810), .B(\modmult_1/zin[0][681] ), .Z(n26648) );
  IV U34499 ( .A(n33807), .Z(n33810) );
  XNOR U34500 ( .A(n33807), .B(n26647), .Z(n33809) );
  XOR U34501 ( .A(n33811), .B(n33812), .Z(n26647) );
  AND U34502 ( .A(\modmult_1/xin[1023] ), .B(n33813), .Z(n33812) );
  IV U34503 ( .A(n33811), .Z(n33813) );
  XOR U34504 ( .A(n33814), .B(g_input[682]), .Z(n33811) );
  NAND U34505 ( .A(n33815), .B(mul_pow), .Z(n33814) );
  XOR U34506 ( .A(g_input[682]), .B(creg[682]), .Z(n33815) );
  XOR U34507 ( .A(n33816), .B(n33817), .Z(n33807) );
  ANDN U34508 ( .A(n33818), .B(n26654), .Z(n33817) );
  XOR U34509 ( .A(n33819), .B(\modmult_1/zin[0][680] ), .Z(n26654) );
  IV U34510 ( .A(n33816), .Z(n33819) );
  XNOR U34511 ( .A(n33816), .B(n26653), .Z(n33818) );
  XOR U34512 ( .A(n33820), .B(n33821), .Z(n26653) );
  AND U34513 ( .A(\modmult_1/xin[1023] ), .B(n33822), .Z(n33821) );
  IV U34514 ( .A(n33820), .Z(n33822) );
  XOR U34515 ( .A(n33823), .B(g_input[681]), .Z(n33820) );
  NAND U34516 ( .A(n33824), .B(mul_pow), .Z(n33823) );
  XOR U34517 ( .A(g_input[681]), .B(creg[681]), .Z(n33824) );
  XOR U34518 ( .A(n33825), .B(n33826), .Z(n33816) );
  ANDN U34519 ( .A(n33827), .B(n26660), .Z(n33826) );
  XOR U34520 ( .A(n33828), .B(\modmult_1/zin[0][679] ), .Z(n26660) );
  IV U34521 ( .A(n33825), .Z(n33828) );
  XNOR U34522 ( .A(n33825), .B(n26659), .Z(n33827) );
  XOR U34523 ( .A(n33829), .B(n33830), .Z(n26659) );
  AND U34524 ( .A(\modmult_1/xin[1023] ), .B(n33831), .Z(n33830) );
  IV U34525 ( .A(n33829), .Z(n33831) );
  XOR U34526 ( .A(n33832), .B(g_input[680]), .Z(n33829) );
  NAND U34527 ( .A(n33833), .B(mul_pow), .Z(n33832) );
  XOR U34528 ( .A(g_input[680]), .B(creg[680]), .Z(n33833) );
  XOR U34529 ( .A(n33834), .B(n33835), .Z(n33825) );
  ANDN U34530 ( .A(n33836), .B(n26666), .Z(n33835) );
  XOR U34531 ( .A(n33837), .B(\modmult_1/zin[0][678] ), .Z(n26666) );
  IV U34532 ( .A(n33834), .Z(n33837) );
  XNOR U34533 ( .A(n33834), .B(n26665), .Z(n33836) );
  XOR U34534 ( .A(n33838), .B(n33839), .Z(n26665) );
  AND U34535 ( .A(\modmult_1/xin[1023] ), .B(n33840), .Z(n33839) );
  IV U34536 ( .A(n33838), .Z(n33840) );
  XOR U34537 ( .A(n33841), .B(g_input[679]), .Z(n33838) );
  NAND U34538 ( .A(n33842), .B(mul_pow), .Z(n33841) );
  XOR U34539 ( .A(g_input[679]), .B(creg[679]), .Z(n33842) );
  XOR U34540 ( .A(n33843), .B(n33844), .Z(n33834) );
  ANDN U34541 ( .A(n33845), .B(n26672), .Z(n33844) );
  XOR U34542 ( .A(n33846), .B(\modmult_1/zin[0][677] ), .Z(n26672) );
  IV U34543 ( .A(n33843), .Z(n33846) );
  XNOR U34544 ( .A(n33843), .B(n26671), .Z(n33845) );
  XOR U34545 ( .A(n33847), .B(n33848), .Z(n26671) );
  AND U34546 ( .A(\modmult_1/xin[1023] ), .B(n33849), .Z(n33848) );
  IV U34547 ( .A(n33847), .Z(n33849) );
  XOR U34548 ( .A(n33850), .B(g_input[678]), .Z(n33847) );
  NAND U34549 ( .A(n33851), .B(mul_pow), .Z(n33850) );
  XOR U34550 ( .A(g_input[678]), .B(creg[678]), .Z(n33851) );
  XOR U34551 ( .A(n33852), .B(n33853), .Z(n33843) );
  ANDN U34552 ( .A(n33854), .B(n26678), .Z(n33853) );
  XOR U34553 ( .A(n33855), .B(\modmult_1/zin[0][676] ), .Z(n26678) );
  IV U34554 ( .A(n33852), .Z(n33855) );
  XNOR U34555 ( .A(n33852), .B(n26677), .Z(n33854) );
  XOR U34556 ( .A(n33856), .B(n33857), .Z(n26677) );
  AND U34557 ( .A(\modmult_1/xin[1023] ), .B(n33858), .Z(n33857) );
  IV U34558 ( .A(n33856), .Z(n33858) );
  XOR U34559 ( .A(n33859), .B(g_input[677]), .Z(n33856) );
  NAND U34560 ( .A(n33860), .B(mul_pow), .Z(n33859) );
  XOR U34561 ( .A(g_input[677]), .B(creg[677]), .Z(n33860) );
  XOR U34562 ( .A(n33861), .B(n33862), .Z(n33852) );
  ANDN U34563 ( .A(n33863), .B(n26684), .Z(n33862) );
  XOR U34564 ( .A(n33864), .B(\modmult_1/zin[0][675] ), .Z(n26684) );
  IV U34565 ( .A(n33861), .Z(n33864) );
  XNOR U34566 ( .A(n33861), .B(n26683), .Z(n33863) );
  XOR U34567 ( .A(n33865), .B(n33866), .Z(n26683) );
  AND U34568 ( .A(\modmult_1/xin[1023] ), .B(n33867), .Z(n33866) );
  IV U34569 ( .A(n33865), .Z(n33867) );
  XOR U34570 ( .A(n33868), .B(g_input[676]), .Z(n33865) );
  NAND U34571 ( .A(n33869), .B(mul_pow), .Z(n33868) );
  XOR U34572 ( .A(g_input[676]), .B(creg[676]), .Z(n33869) );
  XOR U34573 ( .A(n33870), .B(n33871), .Z(n33861) );
  ANDN U34574 ( .A(n33872), .B(n26690), .Z(n33871) );
  XOR U34575 ( .A(n33873), .B(\modmult_1/zin[0][674] ), .Z(n26690) );
  IV U34576 ( .A(n33870), .Z(n33873) );
  XNOR U34577 ( .A(n33870), .B(n26689), .Z(n33872) );
  XOR U34578 ( .A(n33874), .B(n33875), .Z(n26689) );
  AND U34579 ( .A(\modmult_1/xin[1023] ), .B(n33876), .Z(n33875) );
  IV U34580 ( .A(n33874), .Z(n33876) );
  XOR U34581 ( .A(n33877), .B(g_input[675]), .Z(n33874) );
  NAND U34582 ( .A(n33878), .B(mul_pow), .Z(n33877) );
  XOR U34583 ( .A(g_input[675]), .B(creg[675]), .Z(n33878) );
  XOR U34584 ( .A(n33879), .B(n33880), .Z(n33870) );
  ANDN U34585 ( .A(n33881), .B(n26696), .Z(n33880) );
  XOR U34586 ( .A(n33882), .B(\modmult_1/zin[0][673] ), .Z(n26696) );
  IV U34587 ( .A(n33879), .Z(n33882) );
  XNOR U34588 ( .A(n33879), .B(n26695), .Z(n33881) );
  XOR U34589 ( .A(n33883), .B(n33884), .Z(n26695) );
  AND U34590 ( .A(\modmult_1/xin[1023] ), .B(n33885), .Z(n33884) );
  IV U34591 ( .A(n33883), .Z(n33885) );
  XOR U34592 ( .A(n33886), .B(g_input[674]), .Z(n33883) );
  NAND U34593 ( .A(n33887), .B(mul_pow), .Z(n33886) );
  XOR U34594 ( .A(g_input[674]), .B(creg[674]), .Z(n33887) );
  XOR U34595 ( .A(n33888), .B(n33889), .Z(n33879) );
  ANDN U34596 ( .A(n33890), .B(n26702), .Z(n33889) );
  XOR U34597 ( .A(n33891), .B(\modmult_1/zin[0][672] ), .Z(n26702) );
  IV U34598 ( .A(n33888), .Z(n33891) );
  XNOR U34599 ( .A(n33888), .B(n26701), .Z(n33890) );
  XOR U34600 ( .A(n33892), .B(n33893), .Z(n26701) );
  AND U34601 ( .A(\modmult_1/xin[1023] ), .B(n33894), .Z(n33893) );
  IV U34602 ( .A(n33892), .Z(n33894) );
  XOR U34603 ( .A(n33895), .B(g_input[673]), .Z(n33892) );
  NAND U34604 ( .A(n33896), .B(mul_pow), .Z(n33895) );
  XOR U34605 ( .A(g_input[673]), .B(creg[673]), .Z(n33896) );
  XOR U34606 ( .A(n33897), .B(n33898), .Z(n33888) );
  ANDN U34607 ( .A(n33899), .B(n26708), .Z(n33898) );
  XOR U34608 ( .A(n33900), .B(\modmult_1/zin[0][671] ), .Z(n26708) );
  IV U34609 ( .A(n33897), .Z(n33900) );
  XNOR U34610 ( .A(n33897), .B(n26707), .Z(n33899) );
  XOR U34611 ( .A(n33901), .B(n33902), .Z(n26707) );
  AND U34612 ( .A(\modmult_1/xin[1023] ), .B(n33903), .Z(n33902) );
  IV U34613 ( .A(n33901), .Z(n33903) );
  XOR U34614 ( .A(n33904), .B(g_input[672]), .Z(n33901) );
  NAND U34615 ( .A(n33905), .B(mul_pow), .Z(n33904) );
  XOR U34616 ( .A(g_input[672]), .B(creg[672]), .Z(n33905) );
  XOR U34617 ( .A(n33906), .B(n33907), .Z(n33897) );
  ANDN U34618 ( .A(n33908), .B(n26714), .Z(n33907) );
  XOR U34619 ( .A(n33909), .B(\modmult_1/zin[0][670] ), .Z(n26714) );
  IV U34620 ( .A(n33906), .Z(n33909) );
  XNOR U34621 ( .A(n33906), .B(n26713), .Z(n33908) );
  XOR U34622 ( .A(n33910), .B(n33911), .Z(n26713) );
  AND U34623 ( .A(\modmult_1/xin[1023] ), .B(n33912), .Z(n33911) );
  IV U34624 ( .A(n33910), .Z(n33912) );
  XOR U34625 ( .A(n33913), .B(g_input[671]), .Z(n33910) );
  NAND U34626 ( .A(n33914), .B(mul_pow), .Z(n33913) );
  XOR U34627 ( .A(g_input[671]), .B(creg[671]), .Z(n33914) );
  XOR U34628 ( .A(n33915), .B(n33916), .Z(n33906) );
  ANDN U34629 ( .A(n33917), .B(n26720), .Z(n33916) );
  XOR U34630 ( .A(n33918), .B(\modmult_1/zin[0][669] ), .Z(n26720) );
  IV U34631 ( .A(n33915), .Z(n33918) );
  XNOR U34632 ( .A(n33915), .B(n26719), .Z(n33917) );
  XOR U34633 ( .A(n33919), .B(n33920), .Z(n26719) );
  AND U34634 ( .A(\modmult_1/xin[1023] ), .B(n33921), .Z(n33920) );
  IV U34635 ( .A(n33919), .Z(n33921) );
  XOR U34636 ( .A(n33922), .B(g_input[670]), .Z(n33919) );
  NAND U34637 ( .A(n33923), .B(mul_pow), .Z(n33922) );
  XOR U34638 ( .A(g_input[670]), .B(creg[670]), .Z(n33923) );
  XOR U34639 ( .A(n33924), .B(n33925), .Z(n33915) );
  ANDN U34640 ( .A(n33926), .B(n26726), .Z(n33925) );
  XOR U34641 ( .A(n33927), .B(\modmult_1/zin[0][668] ), .Z(n26726) );
  IV U34642 ( .A(n33924), .Z(n33927) );
  XNOR U34643 ( .A(n33924), .B(n26725), .Z(n33926) );
  XOR U34644 ( .A(n33928), .B(n33929), .Z(n26725) );
  AND U34645 ( .A(\modmult_1/xin[1023] ), .B(n33930), .Z(n33929) );
  IV U34646 ( .A(n33928), .Z(n33930) );
  XOR U34647 ( .A(n33931), .B(g_input[669]), .Z(n33928) );
  NAND U34648 ( .A(n33932), .B(mul_pow), .Z(n33931) );
  XOR U34649 ( .A(g_input[669]), .B(creg[669]), .Z(n33932) );
  XOR U34650 ( .A(n33933), .B(n33934), .Z(n33924) );
  ANDN U34651 ( .A(n33935), .B(n26732), .Z(n33934) );
  XOR U34652 ( .A(n33936), .B(\modmult_1/zin[0][667] ), .Z(n26732) );
  IV U34653 ( .A(n33933), .Z(n33936) );
  XNOR U34654 ( .A(n33933), .B(n26731), .Z(n33935) );
  XOR U34655 ( .A(n33937), .B(n33938), .Z(n26731) );
  AND U34656 ( .A(\modmult_1/xin[1023] ), .B(n33939), .Z(n33938) );
  IV U34657 ( .A(n33937), .Z(n33939) );
  XOR U34658 ( .A(n33940), .B(g_input[668]), .Z(n33937) );
  NAND U34659 ( .A(n33941), .B(mul_pow), .Z(n33940) );
  XOR U34660 ( .A(g_input[668]), .B(creg[668]), .Z(n33941) );
  XOR U34661 ( .A(n33942), .B(n33943), .Z(n33933) );
  ANDN U34662 ( .A(n33944), .B(n26738), .Z(n33943) );
  XOR U34663 ( .A(n33945), .B(\modmult_1/zin[0][666] ), .Z(n26738) );
  IV U34664 ( .A(n33942), .Z(n33945) );
  XNOR U34665 ( .A(n33942), .B(n26737), .Z(n33944) );
  XOR U34666 ( .A(n33946), .B(n33947), .Z(n26737) );
  AND U34667 ( .A(\modmult_1/xin[1023] ), .B(n33948), .Z(n33947) );
  IV U34668 ( .A(n33946), .Z(n33948) );
  XOR U34669 ( .A(n33949), .B(g_input[667]), .Z(n33946) );
  NAND U34670 ( .A(n33950), .B(mul_pow), .Z(n33949) );
  XOR U34671 ( .A(g_input[667]), .B(creg[667]), .Z(n33950) );
  XOR U34672 ( .A(n33951), .B(n33952), .Z(n33942) );
  ANDN U34673 ( .A(n33953), .B(n26744), .Z(n33952) );
  XOR U34674 ( .A(n33954), .B(\modmult_1/zin[0][665] ), .Z(n26744) );
  IV U34675 ( .A(n33951), .Z(n33954) );
  XNOR U34676 ( .A(n33951), .B(n26743), .Z(n33953) );
  XOR U34677 ( .A(n33955), .B(n33956), .Z(n26743) );
  AND U34678 ( .A(\modmult_1/xin[1023] ), .B(n33957), .Z(n33956) );
  IV U34679 ( .A(n33955), .Z(n33957) );
  XOR U34680 ( .A(n33958), .B(g_input[666]), .Z(n33955) );
  NAND U34681 ( .A(n33959), .B(mul_pow), .Z(n33958) );
  XOR U34682 ( .A(g_input[666]), .B(creg[666]), .Z(n33959) );
  XOR U34683 ( .A(n33960), .B(n33961), .Z(n33951) );
  ANDN U34684 ( .A(n33962), .B(n26750), .Z(n33961) );
  XOR U34685 ( .A(n33963), .B(\modmult_1/zin[0][664] ), .Z(n26750) );
  IV U34686 ( .A(n33960), .Z(n33963) );
  XNOR U34687 ( .A(n33960), .B(n26749), .Z(n33962) );
  XOR U34688 ( .A(n33964), .B(n33965), .Z(n26749) );
  AND U34689 ( .A(\modmult_1/xin[1023] ), .B(n33966), .Z(n33965) );
  IV U34690 ( .A(n33964), .Z(n33966) );
  XOR U34691 ( .A(n33967), .B(g_input[665]), .Z(n33964) );
  NAND U34692 ( .A(n33968), .B(mul_pow), .Z(n33967) );
  XOR U34693 ( .A(g_input[665]), .B(creg[665]), .Z(n33968) );
  XOR U34694 ( .A(n33969), .B(n33970), .Z(n33960) );
  ANDN U34695 ( .A(n33971), .B(n26756), .Z(n33970) );
  XOR U34696 ( .A(n33972), .B(\modmult_1/zin[0][663] ), .Z(n26756) );
  IV U34697 ( .A(n33969), .Z(n33972) );
  XNOR U34698 ( .A(n33969), .B(n26755), .Z(n33971) );
  XOR U34699 ( .A(n33973), .B(n33974), .Z(n26755) );
  AND U34700 ( .A(\modmult_1/xin[1023] ), .B(n33975), .Z(n33974) );
  IV U34701 ( .A(n33973), .Z(n33975) );
  XOR U34702 ( .A(n33976), .B(g_input[664]), .Z(n33973) );
  NAND U34703 ( .A(n33977), .B(mul_pow), .Z(n33976) );
  XOR U34704 ( .A(g_input[664]), .B(creg[664]), .Z(n33977) );
  XOR U34705 ( .A(n33978), .B(n33979), .Z(n33969) );
  ANDN U34706 ( .A(n33980), .B(n26762), .Z(n33979) );
  XOR U34707 ( .A(n33981), .B(\modmult_1/zin[0][662] ), .Z(n26762) );
  IV U34708 ( .A(n33978), .Z(n33981) );
  XNOR U34709 ( .A(n33978), .B(n26761), .Z(n33980) );
  XOR U34710 ( .A(n33982), .B(n33983), .Z(n26761) );
  AND U34711 ( .A(\modmult_1/xin[1023] ), .B(n33984), .Z(n33983) );
  IV U34712 ( .A(n33982), .Z(n33984) );
  XOR U34713 ( .A(n33985), .B(g_input[663]), .Z(n33982) );
  NAND U34714 ( .A(n33986), .B(mul_pow), .Z(n33985) );
  XOR U34715 ( .A(g_input[663]), .B(creg[663]), .Z(n33986) );
  XOR U34716 ( .A(n33987), .B(n33988), .Z(n33978) );
  ANDN U34717 ( .A(n33989), .B(n26768), .Z(n33988) );
  XOR U34718 ( .A(n33990), .B(\modmult_1/zin[0][661] ), .Z(n26768) );
  IV U34719 ( .A(n33987), .Z(n33990) );
  XNOR U34720 ( .A(n33987), .B(n26767), .Z(n33989) );
  XOR U34721 ( .A(n33991), .B(n33992), .Z(n26767) );
  AND U34722 ( .A(\modmult_1/xin[1023] ), .B(n33993), .Z(n33992) );
  IV U34723 ( .A(n33991), .Z(n33993) );
  XOR U34724 ( .A(n33994), .B(g_input[662]), .Z(n33991) );
  NAND U34725 ( .A(n33995), .B(mul_pow), .Z(n33994) );
  XOR U34726 ( .A(g_input[662]), .B(creg[662]), .Z(n33995) );
  XOR U34727 ( .A(n33996), .B(n33997), .Z(n33987) );
  ANDN U34728 ( .A(n33998), .B(n26774), .Z(n33997) );
  XOR U34729 ( .A(n33999), .B(\modmult_1/zin[0][660] ), .Z(n26774) );
  IV U34730 ( .A(n33996), .Z(n33999) );
  XNOR U34731 ( .A(n33996), .B(n26773), .Z(n33998) );
  XOR U34732 ( .A(n34000), .B(n34001), .Z(n26773) );
  AND U34733 ( .A(\modmult_1/xin[1023] ), .B(n34002), .Z(n34001) );
  IV U34734 ( .A(n34000), .Z(n34002) );
  XOR U34735 ( .A(n34003), .B(g_input[661]), .Z(n34000) );
  NAND U34736 ( .A(n34004), .B(mul_pow), .Z(n34003) );
  XOR U34737 ( .A(g_input[661]), .B(creg[661]), .Z(n34004) );
  XOR U34738 ( .A(n34005), .B(n34006), .Z(n33996) );
  ANDN U34739 ( .A(n34007), .B(n26780), .Z(n34006) );
  XOR U34740 ( .A(n34008), .B(\modmult_1/zin[0][659] ), .Z(n26780) );
  IV U34741 ( .A(n34005), .Z(n34008) );
  XNOR U34742 ( .A(n34005), .B(n26779), .Z(n34007) );
  XOR U34743 ( .A(n34009), .B(n34010), .Z(n26779) );
  AND U34744 ( .A(\modmult_1/xin[1023] ), .B(n34011), .Z(n34010) );
  IV U34745 ( .A(n34009), .Z(n34011) );
  XOR U34746 ( .A(n34012), .B(g_input[660]), .Z(n34009) );
  NAND U34747 ( .A(n34013), .B(mul_pow), .Z(n34012) );
  XOR U34748 ( .A(g_input[660]), .B(creg[660]), .Z(n34013) );
  XOR U34749 ( .A(n34014), .B(n34015), .Z(n34005) );
  ANDN U34750 ( .A(n34016), .B(n26786), .Z(n34015) );
  XOR U34751 ( .A(n34017), .B(\modmult_1/zin[0][658] ), .Z(n26786) );
  IV U34752 ( .A(n34014), .Z(n34017) );
  XNOR U34753 ( .A(n34014), .B(n26785), .Z(n34016) );
  XOR U34754 ( .A(n34018), .B(n34019), .Z(n26785) );
  AND U34755 ( .A(\modmult_1/xin[1023] ), .B(n34020), .Z(n34019) );
  IV U34756 ( .A(n34018), .Z(n34020) );
  XOR U34757 ( .A(n34021), .B(g_input[659]), .Z(n34018) );
  NAND U34758 ( .A(n34022), .B(mul_pow), .Z(n34021) );
  XOR U34759 ( .A(g_input[659]), .B(creg[659]), .Z(n34022) );
  XOR U34760 ( .A(n34023), .B(n34024), .Z(n34014) );
  ANDN U34761 ( .A(n34025), .B(n26792), .Z(n34024) );
  XOR U34762 ( .A(n34026), .B(\modmult_1/zin[0][657] ), .Z(n26792) );
  IV U34763 ( .A(n34023), .Z(n34026) );
  XNOR U34764 ( .A(n34023), .B(n26791), .Z(n34025) );
  XOR U34765 ( .A(n34027), .B(n34028), .Z(n26791) );
  AND U34766 ( .A(\modmult_1/xin[1023] ), .B(n34029), .Z(n34028) );
  IV U34767 ( .A(n34027), .Z(n34029) );
  XOR U34768 ( .A(n34030), .B(g_input[658]), .Z(n34027) );
  NAND U34769 ( .A(n34031), .B(mul_pow), .Z(n34030) );
  XOR U34770 ( .A(g_input[658]), .B(creg[658]), .Z(n34031) );
  XOR U34771 ( .A(n34032), .B(n34033), .Z(n34023) );
  ANDN U34772 ( .A(n34034), .B(n26798), .Z(n34033) );
  XOR U34773 ( .A(n34035), .B(\modmult_1/zin[0][656] ), .Z(n26798) );
  IV U34774 ( .A(n34032), .Z(n34035) );
  XNOR U34775 ( .A(n34032), .B(n26797), .Z(n34034) );
  XOR U34776 ( .A(n34036), .B(n34037), .Z(n26797) );
  AND U34777 ( .A(\modmult_1/xin[1023] ), .B(n34038), .Z(n34037) );
  IV U34778 ( .A(n34036), .Z(n34038) );
  XOR U34779 ( .A(n34039), .B(g_input[657]), .Z(n34036) );
  NAND U34780 ( .A(n34040), .B(mul_pow), .Z(n34039) );
  XOR U34781 ( .A(g_input[657]), .B(creg[657]), .Z(n34040) );
  XOR U34782 ( .A(n34041), .B(n34042), .Z(n34032) );
  ANDN U34783 ( .A(n34043), .B(n26804), .Z(n34042) );
  XOR U34784 ( .A(n34044), .B(\modmult_1/zin[0][655] ), .Z(n26804) );
  IV U34785 ( .A(n34041), .Z(n34044) );
  XNOR U34786 ( .A(n34041), .B(n26803), .Z(n34043) );
  XOR U34787 ( .A(n34045), .B(n34046), .Z(n26803) );
  AND U34788 ( .A(\modmult_1/xin[1023] ), .B(n34047), .Z(n34046) );
  IV U34789 ( .A(n34045), .Z(n34047) );
  XOR U34790 ( .A(n34048), .B(g_input[656]), .Z(n34045) );
  NAND U34791 ( .A(n34049), .B(mul_pow), .Z(n34048) );
  XOR U34792 ( .A(g_input[656]), .B(creg[656]), .Z(n34049) );
  XOR U34793 ( .A(n34050), .B(n34051), .Z(n34041) );
  ANDN U34794 ( .A(n34052), .B(n26810), .Z(n34051) );
  XOR U34795 ( .A(n34053), .B(\modmult_1/zin[0][654] ), .Z(n26810) );
  IV U34796 ( .A(n34050), .Z(n34053) );
  XNOR U34797 ( .A(n34050), .B(n26809), .Z(n34052) );
  XOR U34798 ( .A(n34054), .B(n34055), .Z(n26809) );
  AND U34799 ( .A(\modmult_1/xin[1023] ), .B(n34056), .Z(n34055) );
  IV U34800 ( .A(n34054), .Z(n34056) );
  XOR U34801 ( .A(n34057), .B(g_input[655]), .Z(n34054) );
  NAND U34802 ( .A(n34058), .B(mul_pow), .Z(n34057) );
  XOR U34803 ( .A(g_input[655]), .B(creg[655]), .Z(n34058) );
  XOR U34804 ( .A(n34059), .B(n34060), .Z(n34050) );
  ANDN U34805 ( .A(n34061), .B(n26816), .Z(n34060) );
  XOR U34806 ( .A(n34062), .B(\modmult_1/zin[0][653] ), .Z(n26816) );
  IV U34807 ( .A(n34059), .Z(n34062) );
  XNOR U34808 ( .A(n34059), .B(n26815), .Z(n34061) );
  XOR U34809 ( .A(n34063), .B(n34064), .Z(n26815) );
  AND U34810 ( .A(\modmult_1/xin[1023] ), .B(n34065), .Z(n34064) );
  IV U34811 ( .A(n34063), .Z(n34065) );
  XOR U34812 ( .A(n34066), .B(g_input[654]), .Z(n34063) );
  NAND U34813 ( .A(n34067), .B(mul_pow), .Z(n34066) );
  XOR U34814 ( .A(g_input[654]), .B(creg[654]), .Z(n34067) );
  XOR U34815 ( .A(n34068), .B(n34069), .Z(n34059) );
  ANDN U34816 ( .A(n34070), .B(n26822), .Z(n34069) );
  XOR U34817 ( .A(n34071), .B(\modmult_1/zin[0][652] ), .Z(n26822) );
  IV U34818 ( .A(n34068), .Z(n34071) );
  XNOR U34819 ( .A(n34068), .B(n26821), .Z(n34070) );
  XOR U34820 ( .A(n34072), .B(n34073), .Z(n26821) );
  AND U34821 ( .A(\modmult_1/xin[1023] ), .B(n34074), .Z(n34073) );
  IV U34822 ( .A(n34072), .Z(n34074) );
  XOR U34823 ( .A(n34075), .B(g_input[653]), .Z(n34072) );
  NAND U34824 ( .A(n34076), .B(mul_pow), .Z(n34075) );
  XOR U34825 ( .A(g_input[653]), .B(creg[653]), .Z(n34076) );
  XOR U34826 ( .A(n34077), .B(n34078), .Z(n34068) );
  ANDN U34827 ( .A(n34079), .B(n26828), .Z(n34078) );
  XOR U34828 ( .A(n34080), .B(\modmult_1/zin[0][651] ), .Z(n26828) );
  IV U34829 ( .A(n34077), .Z(n34080) );
  XNOR U34830 ( .A(n34077), .B(n26827), .Z(n34079) );
  XOR U34831 ( .A(n34081), .B(n34082), .Z(n26827) );
  AND U34832 ( .A(\modmult_1/xin[1023] ), .B(n34083), .Z(n34082) );
  IV U34833 ( .A(n34081), .Z(n34083) );
  XOR U34834 ( .A(n34084), .B(g_input[652]), .Z(n34081) );
  NAND U34835 ( .A(n34085), .B(mul_pow), .Z(n34084) );
  XOR U34836 ( .A(g_input[652]), .B(creg[652]), .Z(n34085) );
  XOR U34837 ( .A(n34086), .B(n34087), .Z(n34077) );
  ANDN U34838 ( .A(n34088), .B(n26834), .Z(n34087) );
  XOR U34839 ( .A(n34089), .B(\modmult_1/zin[0][650] ), .Z(n26834) );
  IV U34840 ( .A(n34086), .Z(n34089) );
  XNOR U34841 ( .A(n34086), .B(n26833), .Z(n34088) );
  XOR U34842 ( .A(n34090), .B(n34091), .Z(n26833) );
  AND U34843 ( .A(\modmult_1/xin[1023] ), .B(n34092), .Z(n34091) );
  IV U34844 ( .A(n34090), .Z(n34092) );
  XOR U34845 ( .A(n34093), .B(g_input[651]), .Z(n34090) );
  NAND U34846 ( .A(n34094), .B(mul_pow), .Z(n34093) );
  XOR U34847 ( .A(g_input[651]), .B(creg[651]), .Z(n34094) );
  XOR U34848 ( .A(n34095), .B(n34096), .Z(n34086) );
  ANDN U34849 ( .A(n34097), .B(n26840), .Z(n34096) );
  XOR U34850 ( .A(n34098), .B(\modmult_1/zin[0][649] ), .Z(n26840) );
  IV U34851 ( .A(n34095), .Z(n34098) );
  XNOR U34852 ( .A(n34095), .B(n26839), .Z(n34097) );
  XOR U34853 ( .A(n34099), .B(n34100), .Z(n26839) );
  AND U34854 ( .A(\modmult_1/xin[1023] ), .B(n34101), .Z(n34100) );
  IV U34855 ( .A(n34099), .Z(n34101) );
  XOR U34856 ( .A(n34102), .B(g_input[650]), .Z(n34099) );
  NAND U34857 ( .A(n34103), .B(mul_pow), .Z(n34102) );
  XOR U34858 ( .A(g_input[650]), .B(creg[650]), .Z(n34103) );
  XOR U34859 ( .A(n34104), .B(n34105), .Z(n34095) );
  ANDN U34860 ( .A(n34106), .B(n26846), .Z(n34105) );
  XOR U34861 ( .A(n34107), .B(\modmult_1/zin[0][648] ), .Z(n26846) );
  IV U34862 ( .A(n34104), .Z(n34107) );
  XNOR U34863 ( .A(n34104), .B(n26845), .Z(n34106) );
  XOR U34864 ( .A(n34108), .B(n34109), .Z(n26845) );
  AND U34865 ( .A(\modmult_1/xin[1023] ), .B(n34110), .Z(n34109) );
  IV U34866 ( .A(n34108), .Z(n34110) );
  XOR U34867 ( .A(n34111), .B(g_input[649]), .Z(n34108) );
  NAND U34868 ( .A(n34112), .B(mul_pow), .Z(n34111) );
  XOR U34869 ( .A(g_input[649]), .B(creg[649]), .Z(n34112) );
  XOR U34870 ( .A(n34113), .B(n34114), .Z(n34104) );
  ANDN U34871 ( .A(n34115), .B(n26852), .Z(n34114) );
  XOR U34872 ( .A(n34116), .B(\modmult_1/zin[0][647] ), .Z(n26852) );
  IV U34873 ( .A(n34113), .Z(n34116) );
  XNOR U34874 ( .A(n34113), .B(n26851), .Z(n34115) );
  XOR U34875 ( .A(n34117), .B(n34118), .Z(n26851) );
  AND U34876 ( .A(\modmult_1/xin[1023] ), .B(n34119), .Z(n34118) );
  IV U34877 ( .A(n34117), .Z(n34119) );
  XOR U34878 ( .A(n34120), .B(g_input[648]), .Z(n34117) );
  NAND U34879 ( .A(n34121), .B(mul_pow), .Z(n34120) );
  XOR U34880 ( .A(g_input[648]), .B(creg[648]), .Z(n34121) );
  XOR U34881 ( .A(n34122), .B(n34123), .Z(n34113) );
  ANDN U34882 ( .A(n34124), .B(n26858), .Z(n34123) );
  XOR U34883 ( .A(n34125), .B(\modmult_1/zin[0][646] ), .Z(n26858) );
  IV U34884 ( .A(n34122), .Z(n34125) );
  XNOR U34885 ( .A(n34122), .B(n26857), .Z(n34124) );
  XOR U34886 ( .A(n34126), .B(n34127), .Z(n26857) );
  AND U34887 ( .A(\modmult_1/xin[1023] ), .B(n34128), .Z(n34127) );
  IV U34888 ( .A(n34126), .Z(n34128) );
  XOR U34889 ( .A(n34129), .B(g_input[647]), .Z(n34126) );
  NAND U34890 ( .A(n34130), .B(mul_pow), .Z(n34129) );
  XOR U34891 ( .A(g_input[647]), .B(creg[647]), .Z(n34130) );
  XOR U34892 ( .A(n34131), .B(n34132), .Z(n34122) );
  ANDN U34893 ( .A(n34133), .B(n26864), .Z(n34132) );
  XOR U34894 ( .A(n34134), .B(\modmult_1/zin[0][645] ), .Z(n26864) );
  IV U34895 ( .A(n34131), .Z(n34134) );
  XNOR U34896 ( .A(n34131), .B(n26863), .Z(n34133) );
  XOR U34897 ( .A(n34135), .B(n34136), .Z(n26863) );
  AND U34898 ( .A(\modmult_1/xin[1023] ), .B(n34137), .Z(n34136) );
  IV U34899 ( .A(n34135), .Z(n34137) );
  XOR U34900 ( .A(n34138), .B(g_input[646]), .Z(n34135) );
  NAND U34901 ( .A(n34139), .B(mul_pow), .Z(n34138) );
  XOR U34902 ( .A(g_input[646]), .B(creg[646]), .Z(n34139) );
  XOR U34903 ( .A(n34140), .B(n34141), .Z(n34131) );
  ANDN U34904 ( .A(n34142), .B(n26870), .Z(n34141) );
  XOR U34905 ( .A(n34143), .B(\modmult_1/zin[0][644] ), .Z(n26870) );
  IV U34906 ( .A(n34140), .Z(n34143) );
  XNOR U34907 ( .A(n34140), .B(n26869), .Z(n34142) );
  XOR U34908 ( .A(n34144), .B(n34145), .Z(n26869) );
  AND U34909 ( .A(\modmult_1/xin[1023] ), .B(n34146), .Z(n34145) );
  IV U34910 ( .A(n34144), .Z(n34146) );
  XOR U34911 ( .A(n34147), .B(g_input[645]), .Z(n34144) );
  NAND U34912 ( .A(n34148), .B(mul_pow), .Z(n34147) );
  XOR U34913 ( .A(g_input[645]), .B(creg[645]), .Z(n34148) );
  XOR U34914 ( .A(n34149), .B(n34150), .Z(n34140) );
  ANDN U34915 ( .A(n34151), .B(n26876), .Z(n34150) );
  XOR U34916 ( .A(n34152), .B(\modmult_1/zin[0][643] ), .Z(n26876) );
  IV U34917 ( .A(n34149), .Z(n34152) );
  XNOR U34918 ( .A(n34149), .B(n26875), .Z(n34151) );
  XOR U34919 ( .A(n34153), .B(n34154), .Z(n26875) );
  AND U34920 ( .A(\modmult_1/xin[1023] ), .B(n34155), .Z(n34154) );
  IV U34921 ( .A(n34153), .Z(n34155) );
  XOR U34922 ( .A(n34156), .B(g_input[644]), .Z(n34153) );
  NAND U34923 ( .A(n34157), .B(mul_pow), .Z(n34156) );
  XOR U34924 ( .A(g_input[644]), .B(creg[644]), .Z(n34157) );
  XOR U34925 ( .A(n34158), .B(n34159), .Z(n34149) );
  ANDN U34926 ( .A(n34160), .B(n26882), .Z(n34159) );
  XOR U34927 ( .A(n34161), .B(\modmult_1/zin[0][642] ), .Z(n26882) );
  IV U34928 ( .A(n34158), .Z(n34161) );
  XNOR U34929 ( .A(n34158), .B(n26881), .Z(n34160) );
  XOR U34930 ( .A(n34162), .B(n34163), .Z(n26881) );
  AND U34931 ( .A(\modmult_1/xin[1023] ), .B(n34164), .Z(n34163) );
  IV U34932 ( .A(n34162), .Z(n34164) );
  XOR U34933 ( .A(n34165), .B(g_input[643]), .Z(n34162) );
  NAND U34934 ( .A(n34166), .B(mul_pow), .Z(n34165) );
  XOR U34935 ( .A(g_input[643]), .B(creg[643]), .Z(n34166) );
  XOR U34936 ( .A(n34167), .B(n34168), .Z(n34158) );
  ANDN U34937 ( .A(n34169), .B(n26888), .Z(n34168) );
  XOR U34938 ( .A(n34170), .B(\modmult_1/zin[0][641] ), .Z(n26888) );
  IV U34939 ( .A(n34167), .Z(n34170) );
  XNOR U34940 ( .A(n34167), .B(n26887), .Z(n34169) );
  XOR U34941 ( .A(n34171), .B(n34172), .Z(n26887) );
  AND U34942 ( .A(\modmult_1/xin[1023] ), .B(n34173), .Z(n34172) );
  IV U34943 ( .A(n34171), .Z(n34173) );
  XOR U34944 ( .A(n34174), .B(g_input[642]), .Z(n34171) );
  NAND U34945 ( .A(n34175), .B(mul_pow), .Z(n34174) );
  XOR U34946 ( .A(g_input[642]), .B(creg[642]), .Z(n34175) );
  XOR U34947 ( .A(n34176), .B(n34177), .Z(n34167) );
  ANDN U34948 ( .A(n34178), .B(n26894), .Z(n34177) );
  XOR U34949 ( .A(n34179), .B(\modmult_1/zin[0][640] ), .Z(n26894) );
  IV U34950 ( .A(n34176), .Z(n34179) );
  XNOR U34951 ( .A(n34176), .B(n26893), .Z(n34178) );
  XOR U34952 ( .A(n34180), .B(n34181), .Z(n26893) );
  AND U34953 ( .A(\modmult_1/xin[1023] ), .B(n34182), .Z(n34181) );
  IV U34954 ( .A(n34180), .Z(n34182) );
  XOR U34955 ( .A(n34183), .B(g_input[641]), .Z(n34180) );
  NAND U34956 ( .A(n34184), .B(mul_pow), .Z(n34183) );
  XOR U34957 ( .A(g_input[641]), .B(creg[641]), .Z(n34184) );
  XOR U34958 ( .A(n34185), .B(n34186), .Z(n34176) );
  ANDN U34959 ( .A(n34187), .B(n26900), .Z(n34186) );
  XOR U34960 ( .A(n34188), .B(\modmult_1/zin[0][639] ), .Z(n26900) );
  IV U34961 ( .A(n34185), .Z(n34188) );
  XNOR U34962 ( .A(n34185), .B(n26899), .Z(n34187) );
  XOR U34963 ( .A(n34189), .B(n34190), .Z(n26899) );
  AND U34964 ( .A(\modmult_1/xin[1023] ), .B(n34191), .Z(n34190) );
  IV U34965 ( .A(n34189), .Z(n34191) );
  XOR U34966 ( .A(n34192), .B(g_input[640]), .Z(n34189) );
  NAND U34967 ( .A(n34193), .B(mul_pow), .Z(n34192) );
  XOR U34968 ( .A(g_input[640]), .B(creg[640]), .Z(n34193) );
  XOR U34969 ( .A(n34194), .B(n34195), .Z(n34185) );
  ANDN U34970 ( .A(n34196), .B(n26906), .Z(n34195) );
  XOR U34971 ( .A(n34197), .B(\modmult_1/zin[0][638] ), .Z(n26906) );
  IV U34972 ( .A(n34194), .Z(n34197) );
  XNOR U34973 ( .A(n34194), .B(n26905), .Z(n34196) );
  XOR U34974 ( .A(n34198), .B(n34199), .Z(n26905) );
  AND U34975 ( .A(\modmult_1/xin[1023] ), .B(n34200), .Z(n34199) );
  IV U34976 ( .A(n34198), .Z(n34200) );
  XOR U34977 ( .A(n34201), .B(g_input[639]), .Z(n34198) );
  NAND U34978 ( .A(n34202), .B(mul_pow), .Z(n34201) );
  XOR U34979 ( .A(g_input[639]), .B(creg[639]), .Z(n34202) );
  XOR U34980 ( .A(n34203), .B(n34204), .Z(n34194) );
  ANDN U34981 ( .A(n34205), .B(n26912), .Z(n34204) );
  XOR U34982 ( .A(n34206), .B(\modmult_1/zin[0][637] ), .Z(n26912) );
  IV U34983 ( .A(n34203), .Z(n34206) );
  XNOR U34984 ( .A(n34203), .B(n26911), .Z(n34205) );
  XOR U34985 ( .A(n34207), .B(n34208), .Z(n26911) );
  AND U34986 ( .A(\modmult_1/xin[1023] ), .B(n34209), .Z(n34208) );
  IV U34987 ( .A(n34207), .Z(n34209) );
  XOR U34988 ( .A(n34210), .B(g_input[638]), .Z(n34207) );
  NAND U34989 ( .A(n34211), .B(mul_pow), .Z(n34210) );
  XOR U34990 ( .A(g_input[638]), .B(creg[638]), .Z(n34211) );
  XOR U34991 ( .A(n34212), .B(n34213), .Z(n34203) );
  ANDN U34992 ( .A(n34214), .B(n26918), .Z(n34213) );
  XOR U34993 ( .A(n34215), .B(\modmult_1/zin[0][636] ), .Z(n26918) );
  IV U34994 ( .A(n34212), .Z(n34215) );
  XNOR U34995 ( .A(n34212), .B(n26917), .Z(n34214) );
  XOR U34996 ( .A(n34216), .B(n34217), .Z(n26917) );
  AND U34997 ( .A(\modmult_1/xin[1023] ), .B(n34218), .Z(n34217) );
  IV U34998 ( .A(n34216), .Z(n34218) );
  XOR U34999 ( .A(n34219), .B(g_input[637]), .Z(n34216) );
  NAND U35000 ( .A(n34220), .B(mul_pow), .Z(n34219) );
  XOR U35001 ( .A(g_input[637]), .B(creg[637]), .Z(n34220) );
  XOR U35002 ( .A(n34221), .B(n34222), .Z(n34212) );
  ANDN U35003 ( .A(n34223), .B(n26924), .Z(n34222) );
  XOR U35004 ( .A(n34224), .B(\modmult_1/zin[0][635] ), .Z(n26924) );
  IV U35005 ( .A(n34221), .Z(n34224) );
  XNOR U35006 ( .A(n34221), .B(n26923), .Z(n34223) );
  XOR U35007 ( .A(n34225), .B(n34226), .Z(n26923) );
  AND U35008 ( .A(\modmult_1/xin[1023] ), .B(n34227), .Z(n34226) );
  IV U35009 ( .A(n34225), .Z(n34227) );
  XOR U35010 ( .A(n34228), .B(g_input[636]), .Z(n34225) );
  NAND U35011 ( .A(n34229), .B(mul_pow), .Z(n34228) );
  XOR U35012 ( .A(g_input[636]), .B(creg[636]), .Z(n34229) );
  XOR U35013 ( .A(n34230), .B(n34231), .Z(n34221) );
  ANDN U35014 ( .A(n34232), .B(n26930), .Z(n34231) );
  XOR U35015 ( .A(n34233), .B(\modmult_1/zin[0][634] ), .Z(n26930) );
  IV U35016 ( .A(n34230), .Z(n34233) );
  XNOR U35017 ( .A(n34230), .B(n26929), .Z(n34232) );
  XOR U35018 ( .A(n34234), .B(n34235), .Z(n26929) );
  AND U35019 ( .A(\modmult_1/xin[1023] ), .B(n34236), .Z(n34235) );
  IV U35020 ( .A(n34234), .Z(n34236) );
  XOR U35021 ( .A(n34237), .B(g_input[635]), .Z(n34234) );
  NAND U35022 ( .A(n34238), .B(mul_pow), .Z(n34237) );
  XOR U35023 ( .A(g_input[635]), .B(creg[635]), .Z(n34238) );
  XOR U35024 ( .A(n34239), .B(n34240), .Z(n34230) );
  ANDN U35025 ( .A(n34241), .B(n26936), .Z(n34240) );
  XOR U35026 ( .A(n34242), .B(\modmult_1/zin[0][633] ), .Z(n26936) );
  IV U35027 ( .A(n34239), .Z(n34242) );
  XNOR U35028 ( .A(n34239), .B(n26935), .Z(n34241) );
  XOR U35029 ( .A(n34243), .B(n34244), .Z(n26935) );
  AND U35030 ( .A(\modmult_1/xin[1023] ), .B(n34245), .Z(n34244) );
  IV U35031 ( .A(n34243), .Z(n34245) );
  XOR U35032 ( .A(n34246), .B(g_input[634]), .Z(n34243) );
  NAND U35033 ( .A(n34247), .B(mul_pow), .Z(n34246) );
  XOR U35034 ( .A(g_input[634]), .B(creg[634]), .Z(n34247) );
  XOR U35035 ( .A(n34248), .B(n34249), .Z(n34239) );
  ANDN U35036 ( .A(n34250), .B(n26942), .Z(n34249) );
  XOR U35037 ( .A(n34251), .B(\modmult_1/zin[0][632] ), .Z(n26942) );
  IV U35038 ( .A(n34248), .Z(n34251) );
  XNOR U35039 ( .A(n34248), .B(n26941), .Z(n34250) );
  XOR U35040 ( .A(n34252), .B(n34253), .Z(n26941) );
  AND U35041 ( .A(\modmult_1/xin[1023] ), .B(n34254), .Z(n34253) );
  IV U35042 ( .A(n34252), .Z(n34254) );
  XOR U35043 ( .A(n34255), .B(g_input[633]), .Z(n34252) );
  NAND U35044 ( .A(n34256), .B(mul_pow), .Z(n34255) );
  XOR U35045 ( .A(g_input[633]), .B(creg[633]), .Z(n34256) );
  XOR U35046 ( .A(n34257), .B(n34258), .Z(n34248) );
  ANDN U35047 ( .A(n34259), .B(n26948), .Z(n34258) );
  XOR U35048 ( .A(n34260), .B(\modmult_1/zin[0][631] ), .Z(n26948) );
  IV U35049 ( .A(n34257), .Z(n34260) );
  XNOR U35050 ( .A(n34257), .B(n26947), .Z(n34259) );
  XOR U35051 ( .A(n34261), .B(n34262), .Z(n26947) );
  AND U35052 ( .A(\modmult_1/xin[1023] ), .B(n34263), .Z(n34262) );
  IV U35053 ( .A(n34261), .Z(n34263) );
  XOR U35054 ( .A(n34264), .B(g_input[632]), .Z(n34261) );
  NAND U35055 ( .A(n34265), .B(mul_pow), .Z(n34264) );
  XOR U35056 ( .A(g_input[632]), .B(creg[632]), .Z(n34265) );
  XOR U35057 ( .A(n34266), .B(n34267), .Z(n34257) );
  ANDN U35058 ( .A(n34268), .B(n26954), .Z(n34267) );
  XOR U35059 ( .A(n34269), .B(\modmult_1/zin[0][630] ), .Z(n26954) );
  IV U35060 ( .A(n34266), .Z(n34269) );
  XNOR U35061 ( .A(n34266), .B(n26953), .Z(n34268) );
  XOR U35062 ( .A(n34270), .B(n34271), .Z(n26953) );
  AND U35063 ( .A(\modmult_1/xin[1023] ), .B(n34272), .Z(n34271) );
  IV U35064 ( .A(n34270), .Z(n34272) );
  XOR U35065 ( .A(n34273), .B(g_input[631]), .Z(n34270) );
  NAND U35066 ( .A(n34274), .B(mul_pow), .Z(n34273) );
  XOR U35067 ( .A(g_input[631]), .B(creg[631]), .Z(n34274) );
  XOR U35068 ( .A(n34275), .B(n34276), .Z(n34266) );
  ANDN U35069 ( .A(n34277), .B(n26960), .Z(n34276) );
  XOR U35070 ( .A(n34278), .B(\modmult_1/zin[0][629] ), .Z(n26960) );
  IV U35071 ( .A(n34275), .Z(n34278) );
  XNOR U35072 ( .A(n34275), .B(n26959), .Z(n34277) );
  XOR U35073 ( .A(n34279), .B(n34280), .Z(n26959) );
  AND U35074 ( .A(\modmult_1/xin[1023] ), .B(n34281), .Z(n34280) );
  IV U35075 ( .A(n34279), .Z(n34281) );
  XOR U35076 ( .A(n34282), .B(g_input[630]), .Z(n34279) );
  NAND U35077 ( .A(n34283), .B(mul_pow), .Z(n34282) );
  XOR U35078 ( .A(g_input[630]), .B(creg[630]), .Z(n34283) );
  XOR U35079 ( .A(n34284), .B(n34285), .Z(n34275) );
  ANDN U35080 ( .A(n34286), .B(n26966), .Z(n34285) );
  XOR U35081 ( .A(n34287), .B(\modmult_1/zin[0][628] ), .Z(n26966) );
  IV U35082 ( .A(n34284), .Z(n34287) );
  XNOR U35083 ( .A(n34284), .B(n26965), .Z(n34286) );
  XOR U35084 ( .A(n34288), .B(n34289), .Z(n26965) );
  AND U35085 ( .A(\modmult_1/xin[1023] ), .B(n34290), .Z(n34289) );
  IV U35086 ( .A(n34288), .Z(n34290) );
  XOR U35087 ( .A(n34291), .B(g_input[629]), .Z(n34288) );
  NAND U35088 ( .A(n34292), .B(mul_pow), .Z(n34291) );
  XOR U35089 ( .A(g_input[629]), .B(creg[629]), .Z(n34292) );
  XOR U35090 ( .A(n34293), .B(n34294), .Z(n34284) );
  ANDN U35091 ( .A(n34295), .B(n26972), .Z(n34294) );
  XOR U35092 ( .A(n34296), .B(\modmult_1/zin[0][627] ), .Z(n26972) );
  IV U35093 ( .A(n34293), .Z(n34296) );
  XNOR U35094 ( .A(n34293), .B(n26971), .Z(n34295) );
  XOR U35095 ( .A(n34297), .B(n34298), .Z(n26971) );
  AND U35096 ( .A(\modmult_1/xin[1023] ), .B(n34299), .Z(n34298) );
  IV U35097 ( .A(n34297), .Z(n34299) );
  XOR U35098 ( .A(n34300), .B(g_input[628]), .Z(n34297) );
  NAND U35099 ( .A(n34301), .B(mul_pow), .Z(n34300) );
  XOR U35100 ( .A(g_input[628]), .B(creg[628]), .Z(n34301) );
  XOR U35101 ( .A(n34302), .B(n34303), .Z(n34293) );
  ANDN U35102 ( .A(n34304), .B(n26978), .Z(n34303) );
  XOR U35103 ( .A(n34305), .B(\modmult_1/zin[0][626] ), .Z(n26978) );
  IV U35104 ( .A(n34302), .Z(n34305) );
  XNOR U35105 ( .A(n34302), .B(n26977), .Z(n34304) );
  XOR U35106 ( .A(n34306), .B(n34307), .Z(n26977) );
  AND U35107 ( .A(\modmult_1/xin[1023] ), .B(n34308), .Z(n34307) );
  IV U35108 ( .A(n34306), .Z(n34308) );
  XOR U35109 ( .A(n34309), .B(g_input[627]), .Z(n34306) );
  NAND U35110 ( .A(n34310), .B(mul_pow), .Z(n34309) );
  XOR U35111 ( .A(g_input[627]), .B(creg[627]), .Z(n34310) );
  XOR U35112 ( .A(n34311), .B(n34312), .Z(n34302) );
  ANDN U35113 ( .A(n34313), .B(n26984), .Z(n34312) );
  XOR U35114 ( .A(n34314), .B(\modmult_1/zin[0][625] ), .Z(n26984) );
  IV U35115 ( .A(n34311), .Z(n34314) );
  XNOR U35116 ( .A(n34311), .B(n26983), .Z(n34313) );
  XOR U35117 ( .A(n34315), .B(n34316), .Z(n26983) );
  AND U35118 ( .A(\modmult_1/xin[1023] ), .B(n34317), .Z(n34316) );
  IV U35119 ( .A(n34315), .Z(n34317) );
  XOR U35120 ( .A(n34318), .B(g_input[626]), .Z(n34315) );
  NAND U35121 ( .A(n34319), .B(mul_pow), .Z(n34318) );
  XOR U35122 ( .A(g_input[626]), .B(creg[626]), .Z(n34319) );
  XOR U35123 ( .A(n34320), .B(n34321), .Z(n34311) );
  ANDN U35124 ( .A(n34322), .B(n26990), .Z(n34321) );
  XOR U35125 ( .A(n34323), .B(\modmult_1/zin[0][624] ), .Z(n26990) );
  IV U35126 ( .A(n34320), .Z(n34323) );
  XNOR U35127 ( .A(n34320), .B(n26989), .Z(n34322) );
  XOR U35128 ( .A(n34324), .B(n34325), .Z(n26989) );
  AND U35129 ( .A(\modmult_1/xin[1023] ), .B(n34326), .Z(n34325) );
  IV U35130 ( .A(n34324), .Z(n34326) );
  XOR U35131 ( .A(n34327), .B(g_input[625]), .Z(n34324) );
  NAND U35132 ( .A(n34328), .B(mul_pow), .Z(n34327) );
  XOR U35133 ( .A(g_input[625]), .B(creg[625]), .Z(n34328) );
  XOR U35134 ( .A(n34329), .B(n34330), .Z(n34320) );
  ANDN U35135 ( .A(n34331), .B(n26996), .Z(n34330) );
  XOR U35136 ( .A(n34332), .B(\modmult_1/zin[0][623] ), .Z(n26996) );
  IV U35137 ( .A(n34329), .Z(n34332) );
  XNOR U35138 ( .A(n34329), .B(n26995), .Z(n34331) );
  XOR U35139 ( .A(n34333), .B(n34334), .Z(n26995) );
  AND U35140 ( .A(\modmult_1/xin[1023] ), .B(n34335), .Z(n34334) );
  IV U35141 ( .A(n34333), .Z(n34335) );
  XOR U35142 ( .A(n34336), .B(g_input[624]), .Z(n34333) );
  NAND U35143 ( .A(n34337), .B(mul_pow), .Z(n34336) );
  XOR U35144 ( .A(g_input[624]), .B(creg[624]), .Z(n34337) );
  XOR U35145 ( .A(n34338), .B(n34339), .Z(n34329) );
  ANDN U35146 ( .A(n34340), .B(n27002), .Z(n34339) );
  XOR U35147 ( .A(n34341), .B(\modmult_1/zin[0][622] ), .Z(n27002) );
  IV U35148 ( .A(n34338), .Z(n34341) );
  XNOR U35149 ( .A(n34338), .B(n27001), .Z(n34340) );
  XOR U35150 ( .A(n34342), .B(n34343), .Z(n27001) );
  AND U35151 ( .A(\modmult_1/xin[1023] ), .B(n34344), .Z(n34343) );
  IV U35152 ( .A(n34342), .Z(n34344) );
  XOR U35153 ( .A(n34345), .B(g_input[623]), .Z(n34342) );
  NAND U35154 ( .A(n34346), .B(mul_pow), .Z(n34345) );
  XOR U35155 ( .A(g_input[623]), .B(creg[623]), .Z(n34346) );
  XOR U35156 ( .A(n34347), .B(n34348), .Z(n34338) );
  ANDN U35157 ( .A(n34349), .B(n27008), .Z(n34348) );
  XOR U35158 ( .A(n34350), .B(\modmult_1/zin[0][621] ), .Z(n27008) );
  IV U35159 ( .A(n34347), .Z(n34350) );
  XNOR U35160 ( .A(n34347), .B(n27007), .Z(n34349) );
  XOR U35161 ( .A(n34351), .B(n34352), .Z(n27007) );
  AND U35162 ( .A(\modmult_1/xin[1023] ), .B(n34353), .Z(n34352) );
  IV U35163 ( .A(n34351), .Z(n34353) );
  XOR U35164 ( .A(n34354), .B(g_input[622]), .Z(n34351) );
  NAND U35165 ( .A(n34355), .B(mul_pow), .Z(n34354) );
  XOR U35166 ( .A(g_input[622]), .B(creg[622]), .Z(n34355) );
  XOR U35167 ( .A(n34356), .B(n34357), .Z(n34347) );
  ANDN U35168 ( .A(n34358), .B(n27014), .Z(n34357) );
  XOR U35169 ( .A(n34359), .B(\modmult_1/zin[0][620] ), .Z(n27014) );
  IV U35170 ( .A(n34356), .Z(n34359) );
  XNOR U35171 ( .A(n34356), .B(n27013), .Z(n34358) );
  XOR U35172 ( .A(n34360), .B(n34361), .Z(n27013) );
  AND U35173 ( .A(\modmult_1/xin[1023] ), .B(n34362), .Z(n34361) );
  IV U35174 ( .A(n34360), .Z(n34362) );
  XOR U35175 ( .A(n34363), .B(g_input[621]), .Z(n34360) );
  NAND U35176 ( .A(n34364), .B(mul_pow), .Z(n34363) );
  XOR U35177 ( .A(g_input[621]), .B(creg[621]), .Z(n34364) );
  XOR U35178 ( .A(n34365), .B(n34366), .Z(n34356) );
  ANDN U35179 ( .A(n34367), .B(n27020), .Z(n34366) );
  XOR U35180 ( .A(n34368), .B(\modmult_1/zin[0][619] ), .Z(n27020) );
  IV U35181 ( .A(n34365), .Z(n34368) );
  XNOR U35182 ( .A(n34365), .B(n27019), .Z(n34367) );
  XOR U35183 ( .A(n34369), .B(n34370), .Z(n27019) );
  AND U35184 ( .A(\modmult_1/xin[1023] ), .B(n34371), .Z(n34370) );
  IV U35185 ( .A(n34369), .Z(n34371) );
  XOR U35186 ( .A(n34372), .B(g_input[620]), .Z(n34369) );
  NAND U35187 ( .A(n34373), .B(mul_pow), .Z(n34372) );
  XOR U35188 ( .A(g_input[620]), .B(creg[620]), .Z(n34373) );
  XOR U35189 ( .A(n34374), .B(n34375), .Z(n34365) );
  ANDN U35190 ( .A(n34376), .B(n27026), .Z(n34375) );
  XOR U35191 ( .A(n34377), .B(\modmult_1/zin[0][618] ), .Z(n27026) );
  IV U35192 ( .A(n34374), .Z(n34377) );
  XNOR U35193 ( .A(n34374), .B(n27025), .Z(n34376) );
  XOR U35194 ( .A(n34378), .B(n34379), .Z(n27025) );
  AND U35195 ( .A(\modmult_1/xin[1023] ), .B(n34380), .Z(n34379) );
  IV U35196 ( .A(n34378), .Z(n34380) );
  XOR U35197 ( .A(n34381), .B(g_input[619]), .Z(n34378) );
  NAND U35198 ( .A(n34382), .B(mul_pow), .Z(n34381) );
  XOR U35199 ( .A(g_input[619]), .B(creg[619]), .Z(n34382) );
  XOR U35200 ( .A(n34383), .B(n34384), .Z(n34374) );
  ANDN U35201 ( .A(n34385), .B(n27032), .Z(n34384) );
  XOR U35202 ( .A(n34386), .B(\modmult_1/zin[0][617] ), .Z(n27032) );
  IV U35203 ( .A(n34383), .Z(n34386) );
  XNOR U35204 ( .A(n34383), .B(n27031), .Z(n34385) );
  XOR U35205 ( .A(n34387), .B(n34388), .Z(n27031) );
  AND U35206 ( .A(\modmult_1/xin[1023] ), .B(n34389), .Z(n34388) );
  IV U35207 ( .A(n34387), .Z(n34389) );
  XOR U35208 ( .A(n34390), .B(g_input[618]), .Z(n34387) );
  NAND U35209 ( .A(n34391), .B(mul_pow), .Z(n34390) );
  XOR U35210 ( .A(g_input[618]), .B(creg[618]), .Z(n34391) );
  XOR U35211 ( .A(n34392), .B(n34393), .Z(n34383) );
  ANDN U35212 ( .A(n34394), .B(n27038), .Z(n34393) );
  XOR U35213 ( .A(n34395), .B(\modmult_1/zin[0][616] ), .Z(n27038) );
  IV U35214 ( .A(n34392), .Z(n34395) );
  XNOR U35215 ( .A(n34392), .B(n27037), .Z(n34394) );
  XOR U35216 ( .A(n34396), .B(n34397), .Z(n27037) );
  AND U35217 ( .A(\modmult_1/xin[1023] ), .B(n34398), .Z(n34397) );
  IV U35218 ( .A(n34396), .Z(n34398) );
  XOR U35219 ( .A(n34399), .B(g_input[617]), .Z(n34396) );
  NAND U35220 ( .A(n34400), .B(mul_pow), .Z(n34399) );
  XOR U35221 ( .A(g_input[617]), .B(creg[617]), .Z(n34400) );
  XOR U35222 ( .A(n34401), .B(n34402), .Z(n34392) );
  ANDN U35223 ( .A(n34403), .B(n27044), .Z(n34402) );
  XOR U35224 ( .A(n34404), .B(\modmult_1/zin[0][615] ), .Z(n27044) );
  IV U35225 ( .A(n34401), .Z(n34404) );
  XNOR U35226 ( .A(n34401), .B(n27043), .Z(n34403) );
  XOR U35227 ( .A(n34405), .B(n34406), .Z(n27043) );
  AND U35228 ( .A(\modmult_1/xin[1023] ), .B(n34407), .Z(n34406) );
  IV U35229 ( .A(n34405), .Z(n34407) );
  XOR U35230 ( .A(n34408), .B(g_input[616]), .Z(n34405) );
  NAND U35231 ( .A(n34409), .B(mul_pow), .Z(n34408) );
  XOR U35232 ( .A(g_input[616]), .B(creg[616]), .Z(n34409) );
  XOR U35233 ( .A(n34410), .B(n34411), .Z(n34401) );
  ANDN U35234 ( .A(n34412), .B(n27050), .Z(n34411) );
  XOR U35235 ( .A(n34413), .B(\modmult_1/zin[0][614] ), .Z(n27050) );
  IV U35236 ( .A(n34410), .Z(n34413) );
  XNOR U35237 ( .A(n34410), .B(n27049), .Z(n34412) );
  XOR U35238 ( .A(n34414), .B(n34415), .Z(n27049) );
  AND U35239 ( .A(\modmult_1/xin[1023] ), .B(n34416), .Z(n34415) );
  IV U35240 ( .A(n34414), .Z(n34416) );
  XOR U35241 ( .A(n34417), .B(g_input[615]), .Z(n34414) );
  NAND U35242 ( .A(n34418), .B(mul_pow), .Z(n34417) );
  XOR U35243 ( .A(g_input[615]), .B(creg[615]), .Z(n34418) );
  XOR U35244 ( .A(n34419), .B(n34420), .Z(n34410) );
  ANDN U35245 ( .A(n34421), .B(n27056), .Z(n34420) );
  XOR U35246 ( .A(n34422), .B(\modmult_1/zin[0][613] ), .Z(n27056) );
  IV U35247 ( .A(n34419), .Z(n34422) );
  XNOR U35248 ( .A(n34419), .B(n27055), .Z(n34421) );
  XOR U35249 ( .A(n34423), .B(n34424), .Z(n27055) );
  AND U35250 ( .A(\modmult_1/xin[1023] ), .B(n34425), .Z(n34424) );
  IV U35251 ( .A(n34423), .Z(n34425) );
  XOR U35252 ( .A(n34426), .B(g_input[614]), .Z(n34423) );
  NAND U35253 ( .A(n34427), .B(mul_pow), .Z(n34426) );
  XOR U35254 ( .A(g_input[614]), .B(creg[614]), .Z(n34427) );
  XOR U35255 ( .A(n34428), .B(n34429), .Z(n34419) );
  ANDN U35256 ( .A(n34430), .B(n27062), .Z(n34429) );
  XOR U35257 ( .A(n34431), .B(\modmult_1/zin[0][612] ), .Z(n27062) );
  IV U35258 ( .A(n34428), .Z(n34431) );
  XNOR U35259 ( .A(n34428), .B(n27061), .Z(n34430) );
  XOR U35260 ( .A(n34432), .B(n34433), .Z(n27061) );
  AND U35261 ( .A(\modmult_1/xin[1023] ), .B(n34434), .Z(n34433) );
  IV U35262 ( .A(n34432), .Z(n34434) );
  XOR U35263 ( .A(n34435), .B(g_input[613]), .Z(n34432) );
  NAND U35264 ( .A(n34436), .B(mul_pow), .Z(n34435) );
  XOR U35265 ( .A(g_input[613]), .B(creg[613]), .Z(n34436) );
  XOR U35266 ( .A(n34437), .B(n34438), .Z(n34428) );
  ANDN U35267 ( .A(n34439), .B(n27068), .Z(n34438) );
  XOR U35268 ( .A(n34440), .B(\modmult_1/zin[0][611] ), .Z(n27068) );
  IV U35269 ( .A(n34437), .Z(n34440) );
  XNOR U35270 ( .A(n34437), .B(n27067), .Z(n34439) );
  XOR U35271 ( .A(n34441), .B(n34442), .Z(n27067) );
  AND U35272 ( .A(\modmult_1/xin[1023] ), .B(n34443), .Z(n34442) );
  IV U35273 ( .A(n34441), .Z(n34443) );
  XOR U35274 ( .A(n34444), .B(g_input[612]), .Z(n34441) );
  NAND U35275 ( .A(n34445), .B(mul_pow), .Z(n34444) );
  XOR U35276 ( .A(g_input[612]), .B(creg[612]), .Z(n34445) );
  XOR U35277 ( .A(n34446), .B(n34447), .Z(n34437) );
  ANDN U35278 ( .A(n34448), .B(n27074), .Z(n34447) );
  XOR U35279 ( .A(n34449), .B(\modmult_1/zin[0][610] ), .Z(n27074) );
  IV U35280 ( .A(n34446), .Z(n34449) );
  XNOR U35281 ( .A(n34446), .B(n27073), .Z(n34448) );
  XOR U35282 ( .A(n34450), .B(n34451), .Z(n27073) );
  AND U35283 ( .A(\modmult_1/xin[1023] ), .B(n34452), .Z(n34451) );
  IV U35284 ( .A(n34450), .Z(n34452) );
  XOR U35285 ( .A(n34453), .B(g_input[611]), .Z(n34450) );
  NAND U35286 ( .A(n34454), .B(mul_pow), .Z(n34453) );
  XOR U35287 ( .A(g_input[611]), .B(creg[611]), .Z(n34454) );
  XOR U35288 ( .A(n34455), .B(n34456), .Z(n34446) );
  ANDN U35289 ( .A(n34457), .B(n27080), .Z(n34456) );
  XOR U35290 ( .A(n34458), .B(\modmult_1/zin[0][609] ), .Z(n27080) );
  IV U35291 ( .A(n34455), .Z(n34458) );
  XNOR U35292 ( .A(n34455), .B(n27079), .Z(n34457) );
  XOR U35293 ( .A(n34459), .B(n34460), .Z(n27079) );
  AND U35294 ( .A(\modmult_1/xin[1023] ), .B(n34461), .Z(n34460) );
  IV U35295 ( .A(n34459), .Z(n34461) );
  XOR U35296 ( .A(n34462), .B(g_input[610]), .Z(n34459) );
  NAND U35297 ( .A(n34463), .B(mul_pow), .Z(n34462) );
  XOR U35298 ( .A(g_input[610]), .B(creg[610]), .Z(n34463) );
  XOR U35299 ( .A(n34464), .B(n34465), .Z(n34455) );
  ANDN U35300 ( .A(n34466), .B(n27086), .Z(n34465) );
  XOR U35301 ( .A(n34467), .B(\modmult_1/zin[0][608] ), .Z(n27086) );
  IV U35302 ( .A(n34464), .Z(n34467) );
  XNOR U35303 ( .A(n34464), .B(n27085), .Z(n34466) );
  XOR U35304 ( .A(n34468), .B(n34469), .Z(n27085) );
  AND U35305 ( .A(\modmult_1/xin[1023] ), .B(n34470), .Z(n34469) );
  IV U35306 ( .A(n34468), .Z(n34470) );
  XOR U35307 ( .A(n34471), .B(g_input[609]), .Z(n34468) );
  NAND U35308 ( .A(n34472), .B(mul_pow), .Z(n34471) );
  XOR U35309 ( .A(g_input[609]), .B(creg[609]), .Z(n34472) );
  XOR U35310 ( .A(n34473), .B(n34474), .Z(n34464) );
  ANDN U35311 ( .A(n34475), .B(n27092), .Z(n34474) );
  XOR U35312 ( .A(n34476), .B(\modmult_1/zin[0][607] ), .Z(n27092) );
  IV U35313 ( .A(n34473), .Z(n34476) );
  XNOR U35314 ( .A(n34473), .B(n27091), .Z(n34475) );
  XOR U35315 ( .A(n34477), .B(n34478), .Z(n27091) );
  AND U35316 ( .A(\modmult_1/xin[1023] ), .B(n34479), .Z(n34478) );
  IV U35317 ( .A(n34477), .Z(n34479) );
  XOR U35318 ( .A(n34480), .B(g_input[608]), .Z(n34477) );
  NAND U35319 ( .A(n34481), .B(mul_pow), .Z(n34480) );
  XOR U35320 ( .A(g_input[608]), .B(creg[608]), .Z(n34481) );
  XOR U35321 ( .A(n34482), .B(n34483), .Z(n34473) );
  ANDN U35322 ( .A(n34484), .B(n27098), .Z(n34483) );
  XOR U35323 ( .A(n34485), .B(\modmult_1/zin[0][606] ), .Z(n27098) );
  IV U35324 ( .A(n34482), .Z(n34485) );
  XNOR U35325 ( .A(n34482), .B(n27097), .Z(n34484) );
  XOR U35326 ( .A(n34486), .B(n34487), .Z(n27097) );
  AND U35327 ( .A(\modmult_1/xin[1023] ), .B(n34488), .Z(n34487) );
  IV U35328 ( .A(n34486), .Z(n34488) );
  XOR U35329 ( .A(n34489), .B(g_input[607]), .Z(n34486) );
  NAND U35330 ( .A(n34490), .B(mul_pow), .Z(n34489) );
  XOR U35331 ( .A(g_input[607]), .B(creg[607]), .Z(n34490) );
  XOR U35332 ( .A(n34491), .B(n34492), .Z(n34482) );
  ANDN U35333 ( .A(n34493), .B(n27104), .Z(n34492) );
  XOR U35334 ( .A(n34494), .B(\modmult_1/zin[0][605] ), .Z(n27104) );
  IV U35335 ( .A(n34491), .Z(n34494) );
  XNOR U35336 ( .A(n34491), .B(n27103), .Z(n34493) );
  XOR U35337 ( .A(n34495), .B(n34496), .Z(n27103) );
  AND U35338 ( .A(\modmult_1/xin[1023] ), .B(n34497), .Z(n34496) );
  IV U35339 ( .A(n34495), .Z(n34497) );
  XOR U35340 ( .A(n34498), .B(g_input[606]), .Z(n34495) );
  NAND U35341 ( .A(n34499), .B(mul_pow), .Z(n34498) );
  XOR U35342 ( .A(g_input[606]), .B(creg[606]), .Z(n34499) );
  XOR U35343 ( .A(n34500), .B(n34501), .Z(n34491) );
  ANDN U35344 ( .A(n34502), .B(n27110), .Z(n34501) );
  XOR U35345 ( .A(n34503), .B(\modmult_1/zin[0][604] ), .Z(n27110) );
  IV U35346 ( .A(n34500), .Z(n34503) );
  XNOR U35347 ( .A(n34500), .B(n27109), .Z(n34502) );
  XOR U35348 ( .A(n34504), .B(n34505), .Z(n27109) );
  AND U35349 ( .A(\modmult_1/xin[1023] ), .B(n34506), .Z(n34505) );
  IV U35350 ( .A(n34504), .Z(n34506) );
  XOR U35351 ( .A(n34507), .B(g_input[605]), .Z(n34504) );
  NAND U35352 ( .A(n34508), .B(mul_pow), .Z(n34507) );
  XOR U35353 ( .A(g_input[605]), .B(creg[605]), .Z(n34508) );
  XOR U35354 ( .A(n34509), .B(n34510), .Z(n34500) );
  ANDN U35355 ( .A(n34511), .B(n27116), .Z(n34510) );
  XOR U35356 ( .A(n34512), .B(\modmult_1/zin[0][603] ), .Z(n27116) );
  IV U35357 ( .A(n34509), .Z(n34512) );
  XNOR U35358 ( .A(n34509), .B(n27115), .Z(n34511) );
  XOR U35359 ( .A(n34513), .B(n34514), .Z(n27115) );
  AND U35360 ( .A(\modmult_1/xin[1023] ), .B(n34515), .Z(n34514) );
  IV U35361 ( .A(n34513), .Z(n34515) );
  XOR U35362 ( .A(n34516), .B(g_input[604]), .Z(n34513) );
  NAND U35363 ( .A(n34517), .B(mul_pow), .Z(n34516) );
  XOR U35364 ( .A(g_input[604]), .B(creg[604]), .Z(n34517) );
  XOR U35365 ( .A(n34518), .B(n34519), .Z(n34509) );
  ANDN U35366 ( .A(n34520), .B(n27122), .Z(n34519) );
  XOR U35367 ( .A(n34521), .B(\modmult_1/zin[0][602] ), .Z(n27122) );
  IV U35368 ( .A(n34518), .Z(n34521) );
  XNOR U35369 ( .A(n34518), .B(n27121), .Z(n34520) );
  XOR U35370 ( .A(n34522), .B(n34523), .Z(n27121) );
  AND U35371 ( .A(\modmult_1/xin[1023] ), .B(n34524), .Z(n34523) );
  IV U35372 ( .A(n34522), .Z(n34524) );
  XOR U35373 ( .A(n34525), .B(g_input[603]), .Z(n34522) );
  NAND U35374 ( .A(n34526), .B(mul_pow), .Z(n34525) );
  XOR U35375 ( .A(g_input[603]), .B(creg[603]), .Z(n34526) );
  XOR U35376 ( .A(n34527), .B(n34528), .Z(n34518) );
  ANDN U35377 ( .A(n34529), .B(n27128), .Z(n34528) );
  XOR U35378 ( .A(n34530), .B(\modmult_1/zin[0][601] ), .Z(n27128) );
  IV U35379 ( .A(n34527), .Z(n34530) );
  XNOR U35380 ( .A(n34527), .B(n27127), .Z(n34529) );
  XOR U35381 ( .A(n34531), .B(n34532), .Z(n27127) );
  AND U35382 ( .A(\modmult_1/xin[1023] ), .B(n34533), .Z(n34532) );
  IV U35383 ( .A(n34531), .Z(n34533) );
  XOR U35384 ( .A(n34534), .B(g_input[602]), .Z(n34531) );
  NAND U35385 ( .A(n34535), .B(mul_pow), .Z(n34534) );
  XOR U35386 ( .A(g_input[602]), .B(creg[602]), .Z(n34535) );
  XOR U35387 ( .A(n34536), .B(n34537), .Z(n34527) );
  ANDN U35388 ( .A(n34538), .B(n27134), .Z(n34537) );
  XOR U35389 ( .A(n34539), .B(\modmult_1/zin[0][600] ), .Z(n27134) );
  IV U35390 ( .A(n34536), .Z(n34539) );
  XNOR U35391 ( .A(n34536), .B(n27133), .Z(n34538) );
  XOR U35392 ( .A(n34540), .B(n34541), .Z(n27133) );
  AND U35393 ( .A(\modmult_1/xin[1023] ), .B(n34542), .Z(n34541) );
  IV U35394 ( .A(n34540), .Z(n34542) );
  XOR U35395 ( .A(n34543), .B(g_input[601]), .Z(n34540) );
  NAND U35396 ( .A(n34544), .B(mul_pow), .Z(n34543) );
  XOR U35397 ( .A(g_input[601]), .B(creg[601]), .Z(n34544) );
  XOR U35398 ( .A(n34545), .B(n34546), .Z(n34536) );
  ANDN U35399 ( .A(n34547), .B(n27140), .Z(n34546) );
  XOR U35400 ( .A(n34548), .B(\modmult_1/zin[0][599] ), .Z(n27140) );
  IV U35401 ( .A(n34545), .Z(n34548) );
  XNOR U35402 ( .A(n34545), .B(n27139), .Z(n34547) );
  XOR U35403 ( .A(n34549), .B(n34550), .Z(n27139) );
  AND U35404 ( .A(\modmult_1/xin[1023] ), .B(n34551), .Z(n34550) );
  IV U35405 ( .A(n34549), .Z(n34551) );
  XOR U35406 ( .A(n34552), .B(g_input[600]), .Z(n34549) );
  NAND U35407 ( .A(n34553), .B(mul_pow), .Z(n34552) );
  XOR U35408 ( .A(g_input[600]), .B(creg[600]), .Z(n34553) );
  XOR U35409 ( .A(n34554), .B(n34555), .Z(n34545) );
  ANDN U35410 ( .A(n34556), .B(n27146), .Z(n34555) );
  XOR U35411 ( .A(n34557), .B(\modmult_1/zin[0][598] ), .Z(n27146) );
  IV U35412 ( .A(n34554), .Z(n34557) );
  XNOR U35413 ( .A(n34554), .B(n27145), .Z(n34556) );
  XOR U35414 ( .A(n34558), .B(n34559), .Z(n27145) );
  AND U35415 ( .A(\modmult_1/xin[1023] ), .B(n34560), .Z(n34559) );
  IV U35416 ( .A(n34558), .Z(n34560) );
  XOR U35417 ( .A(n34561), .B(g_input[599]), .Z(n34558) );
  NAND U35418 ( .A(n34562), .B(mul_pow), .Z(n34561) );
  XOR U35419 ( .A(g_input[599]), .B(creg[599]), .Z(n34562) );
  XOR U35420 ( .A(n34563), .B(n34564), .Z(n34554) );
  ANDN U35421 ( .A(n34565), .B(n27152), .Z(n34564) );
  XOR U35422 ( .A(n34566), .B(\modmult_1/zin[0][597] ), .Z(n27152) );
  IV U35423 ( .A(n34563), .Z(n34566) );
  XNOR U35424 ( .A(n34563), .B(n27151), .Z(n34565) );
  XOR U35425 ( .A(n34567), .B(n34568), .Z(n27151) );
  AND U35426 ( .A(\modmult_1/xin[1023] ), .B(n34569), .Z(n34568) );
  IV U35427 ( .A(n34567), .Z(n34569) );
  XOR U35428 ( .A(n34570), .B(g_input[598]), .Z(n34567) );
  NAND U35429 ( .A(n34571), .B(mul_pow), .Z(n34570) );
  XOR U35430 ( .A(g_input[598]), .B(creg[598]), .Z(n34571) );
  XOR U35431 ( .A(n34572), .B(n34573), .Z(n34563) );
  ANDN U35432 ( .A(n34574), .B(n27158), .Z(n34573) );
  XOR U35433 ( .A(n34575), .B(\modmult_1/zin[0][596] ), .Z(n27158) );
  IV U35434 ( .A(n34572), .Z(n34575) );
  XNOR U35435 ( .A(n34572), .B(n27157), .Z(n34574) );
  XOR U35436 ( .A(n34576), .B(n34577), .Z(n27157) );
  AND U35437 ( .A(\modmult_1/xin[1023] ), .B(n34578), .Z(n34577) );
  IV U35438 ( .A(n34576), .Z(n34578) );
  XOR U35439 ( .A(n34579), .B(g_input[597]), .Z(n34576) );
  NAND U35440 ( .A(n34580), .B(mul_pow), .Z(n34579) );
  XOR U35441 ( .A(g_input[597]), .B(creg[597]), .Z(n34580) );
  XOR U35442 ( .A(n34581), .B(n34582), .Z(n34572) );
  ANDN U35443 ( .A(n34583), .B(n27164), .Z(n34582) );
  XOR U35444 ( .A(n34584), .B(\modmult_1/zin[0][595] ), .Z(n27164) );
  IV U35445 ( .A(n34581), .Z(n34584) );
  XNOR U35446 ( .A(n34581), .B(n27163), .Z(n34583) );
  XOR U35447 ( .A(n34585), .B(n34586), .Z(n27163) );
  AND U35448 ( .A(\modmult_1/xin[1023] ), .B(n34587), .Z(n34586) );
  IV U35449 ( .A(n34585), .Z(n34587) );
  XOR U35450 ( .A(n34588), .B(g_input[596]), .Z(n34585) );
  NAND U35451 ( .A(n34589), .B(mul_pow), .Z(n34588) );
  XOR U35452 ( .A(g_input[596]), .B(creg[596]), .Z(n34589) );
  XOR U35453 ( .A(n34590), .B(n34591), .Z(n34581) );
  ANDN U35454 ( .A(n34592), .B(n27170), .Z(n34591) );
  XOR U35455 ( .A(n34593), .B(\modmult_1/zin[0][594] ), .Z(n27170) );
  IV U35456 ( .A(n34590), .Z(n34593) );
  XNOR U35457 ( .A(n34590), .B(n27169), .Z(n34592) );
  XOR U35458 ( .A(n34594), .B(n34595), .Z(n27169) );
  AND U35459 ( .A(\modmult_1/xin[1023] ), .B(n34596), .Z(n34595) );
  IV U35460 ( .A(n34594), .Z(n34596) );
  XOR U35461 ( .A(n34597), .B(g_input[595]), .Z(n34594) );
  NAND U35462 ( .A(n34598), .B(mul_pow), .Z(n34597) );
  XOR U35463 ( .A(g_input[595]), .B(creg[595]), .Z(n34598) );
  XOR U35464 ( .A(n34599), .B(n34600), .Z(n34590) );
  ANDN U35465 ( .A(n34601), .B(n27176), .Z(n34600) );
  XOR U35466 ( .A(n34602), .B(\modmult_1/zin[0][593] ), .Z(n27176) );
  IV U35467 ( .A(n34599), .Z(n34602) );
  XNOR U35468 ( .A(n34599), .B(n27175), .Z(n34601) );
  XOR U35469 ( .A(n34603), .B(n34604), .Z(n27175) );
  AND U35470 ( .A(\modmult_1/xin[1023] ), .B(n34605), .Z(n34604) );
  IV U35471 ( .A(n34603), .Z(n34605) );
  XOR U35472 ( .A(n34606), .B(g_input[594]), .Z(n34603) );
  NAND U35473 ( .A(n34607), .B(mul_pow), .Z(n34606) );
  XOR U35474 ( .A(g_input[594]), .B(creg[594]), .Z(n34607) );
  XOR U35475 ( .A(n34608), .B(n34609), .Z(n34599) );
  ANDN U35476 ( .A(n34610), .B(n27182), .Z(n34609) );
  XOR U35477 ( .A(n34611), .B(\modmult_1/zin[0][592] ), .Z(n27182) );
  IV U35478 ( .A(n34608), .Z(n34611) );
  XNOR U35479 ( .A(n34608), .B(n27181), .Z(n34610) );
  XOR U35480 ( .A(n34612), .B(n34613), .Z(n27181) );
  AND U35481 ( .A(\modmult_1/xin[1023] ), .B(n34614), .Z(n34613) );
  IV U35482 ( .A(n34612), .Z(n34614) );
  XOR U35483 ( .A(n34615), .B(g_input[593]), .Z(n34612) );
  NAND U35484 ( .A(n34616), .B(mul_pow), .Z(n34615) );
  XOR U35485 ( .A(g_input[593]), .B(creg[593]), .Z(n34616) );
  XOR U35486 ( .A(n34617), .B(n34618), .Z(n34608) );
  ANDN U35487 ( .A(n34619), .B(n27188), .Z(n34618) );
  XOR U35488 ( .A(n34620), .B(\modmult_1/zin[0][591] ), .Z(n27188) );
  IV U35489 ( .A(n34617), .Z(n34620) );
  XNOR U35490 ( .A(n34617), .B(n27187), .Z(n34619) );
  XOR U35491 ( .A(n34621), .B(n34622), .Z(n27187) );
  AND U35492 ( .A(\modmult_1/xin[1023] ), .B(n34623), .Z(n34622) );
  IV U35493 ( .A(n34621), .Z(n34623) );
  XOR U35494 ( .A(n34624), .B(g_input[592]), .Z(n34621) );
  NAND U35495 ( .A(n34625), .B(mul_pow), .Z(n34624) );
  XOR U35496 ( .A(g_input[592]), .B(creg[592]), .Z(n34625) );
  XOR U35497 ( .A(n34626), .B(n34627), .Z(n34617) );
  ANDN U35498 ( .A(n34628), .B(n27194), .Z(n34627) );
  XOR U35499 ( .A(n34629), .B(\modmult_1/zin[0][590] ), .Z(n27194) );
  IV U35500 ( .A(n34626), .Z(n34629) );
  XNOR U35501 ( .A(n34626), .B(n27193), .Z(n34628) );
  XOR U35502 ( .A(n34630), .B(n34631), .Z(n27193) );
  AND U35503 ( .A(\modmult_1/xin[1023] ), .B(n34632), .Z(n34631) );
  IV U35504 ( .A(n34630), .Z(n34632) );
  XOR U35505 ( .A(n34633), .B(g_input[591]), .Z(n34630) );
  NAND U35506 ( .A(n34634), .B(mul_pow), .Z(n34633) );
  XOR U35507 ( .A(g_input[591]), .B(creg[591]), .Z(n34634) );
  XOR U35508 ( .A(n34635), .B(n34636), .Z(n34626) );
  ANDN U35509 ( .A(n34637), .B(n27200), .Z(n34636) );
  XOR U35510 ( .A(n34638), .B(\modmult_1/zin[0][589] ), .Z(n27200) );
  IV U35511 ( .A(n34635), .Z(n34638) );
  XNOR U35512 ( .A(n34635), .B(n27199), .Z(n34637) );
  XOR U35513 ( .A(n34639), .B(n34640), .Z(n27199) );
  AND U35514 ( .A(\modmult_1/xin[1023] ), .B(n34641), .Z(n34640) );
  IV U35515 ( .A(n34639), .Z(n34641) );
  XOR U35516 ( .A(n34642), .B(g_input[590]), .Z(n34639) );
  NAND U35517 ( .A(n34643), .B(mul_pow), .Z(n34642) );
  XOR U35518 ( .A(g_input[590]), .B(creg[590]), .Z(n34643) );
  XOR U35519 ( .A(n34644), .B(n34645), .Z(n34635) );
  ANDN U35520 ( .A(n34646), .B(n27206), .Z(n34645) );
  XOR U35521 ( .A(n34647), .B(\modmult_1/zin[0][588] ), .Z(n27206) );
  IV U35522 ( .A(n34644), .Z(n34647) );
  XNOR U35523 ( .A(n34644), .B(n27205), .Z(n34646) );
  XOR U35524 ( .A(n34648), .B(n34649), .Z(n27205) );
  AND U35525 ( .A(\modmult_1/xin[1023] ), .B(n34650), .Z(n34649) );
  IV U35526 ( .A(n34648), .Z(n34650) );
  XOR U35527 ( .A(n34651), .B(g_input[589]), .Z(n34648) );
  NAND U35528 ( .A(n34652), .B(mul_pow), .Z(n34651) );
  XOR U35529 ( .A(g_input[589]), .B(creg[589]), .Z(n34652) );
  XOR U35530 ( .A(n34653), .B(n34654), .Z(n34644) );
  ANDN U35531 ( .A(n34655), .B(n27212), .Z(n34654) );
  XOR U35532 ( .A(n34656), .B(\modmult_1/zin[0][587] ), .Z(n27212) );
  IV U35533 ( .A(n34653), .Z(n34656) );
  XNOR U35534 ( .A(n34653), .B(n27211), .Z(n34655) );
  XOR U35535 ( .A(n34657), .B(n34658), .Z(n27211) );
  AND U35536 ( .A(\modmult_1/xin[1023] ), .B(n34659), .Z(n34658) );
  IV U35537 ( .A(n34657), .Z(n34659) );
  XOR U35538 ( .A(n34660), .B(g_input[588]), .Z(n34657) );
  NAND U35539 ( .A(n34661), .B(mul_pow), .Z(n34660) );
  XOR U35540 ( .A(g_input[588]), .B(creg[588]), .Z(n34661) );
  XOR U35541 ( .A(n34662), .B(n34663), .Z(n34653) );
  ANDN U35542 ( .A(n34664), .B(n27218), .Z(n34663) );
  XOR U35543 ( .A(n34665), .B(\modmult_1/zin[0][586] ), .Z(n27218) );
  IV U35544 ( .A(n34662), .Z(n34665) );
  XNOR U35545 ( .A(n34662), .B(n27217), .Z(n34664) );
  XOR U35546 ( .A(n34666), .B(n34667), .Z(n27217) );
  AND U35547 ( .A(\modmult_1/xin[1023] ), .B(n34668), .Z(n34667) );
  IV U35548 ( .A(n34666), .Z(n34668) );
  XOR U35549 ( .A(n34669), .B(g_input[587]), .Z(n34666) );
  NAND U35550 ( .A(n34670), .B(mul_pow), .Z(n34669) );
  XOR U35551 ( .A(g_input[587]), .B(creg[587]), .Z(n34670) );
  XOR U35552 ( .A(n34671), .B(n34672), .Z(n34662) );
  ANDN U35553 ( .A(n34673), .B(n27224), .Z(n34672) );
  XOR U35554 ( .A(n34674), .B(\modmult_1/zin[0][585] ), .Z(n27224) );
  IV U35555 ( .A(n34671), .Z(n34674) );
  XNOR U35556 ( .A(n34671), .B(n27223), .Z(n34673) );
  XOR U35557 ( .A(n34675), .B(n34676), .Z(n27223) );
  AND U35558 ( .A(\modmult_1/xin[1023] ), .B(n34677), .Z(n34676) );
  IV U35559 ( .A(n34675), .Z(n34677) );
  XOR U35560 ( .A(n34678), .B(g_input[586]), .Z(n34675) );
  NAND U35561 ( .A(n34679), .B(mul_pow), .Z(n34678) );
  XOR U35562 ( .A(g_input[586]), .B(creg[586]), .Z(n34679) );
  XOR U35563 ( .A(n34680), .B(n34681), .Z(n34671) );
  ANDN U35564 ( .A(n34682), .B(n27230), .Z(n34681) );
  XOR U35565 ( .A(n34683), .B(\modmult_1/zin[0][584] ), .Z(n27230) );
  IV U35566 ( .A(n34680), .Z(n34683) );
  XNOR U35567 ( .A(n34680), .B(n27229), .Z(n34682) );
  XOR U35568 ( .A(n34684), .B(n34685), .Z(n27229) );
  AND U35569 ( .A(\modmult_1/xin[1023] ), .B(n34686), .Z(n34685) );
  IV U35570 ( .A(n34684), .Z(n34686) );
  XOR U35571 ( .A(n34687), .B(g_input[585]), .Z(n34684) );
  NAND U35572 ( .A(n34688), .B(mul_pow), .Z(n34687) );
  XOR U35573 ( .A(g_input[585]), .B(creg[585]), .Z(n34688) );
  XOR U35574 ( .A(n34689), .B(n34690), .Z(n34680) );
  ANDN U35575 ( .A(n34691), .B(n27236), .Z(n34690) );
  XOR U35576 ( .A(n34692), .B(\modmult_1/zin[0][583] ), .Z(n27236) );
  IV U35577 ( .A(n34689), .Z(n34692) );
  XNOR U35578 ( .A(n34689), .B(n27235), .Z(n34691) );
  XOR U35579 ( .A(n34693), .B(n34694), .Z(n27235) );
  AND U35580 ( .A(\modmult_1/xin[1023] ), .B(n34695), .Z(n34694) );
  IV U35581 ( .A(n34693), .Z(n34695) );
  XOR U35582 ( .A(n34696), .B(g_input[584]), .Z(n34693) );
  NAND U35583 ( .A(n34697), .B(mul_pow), .Z(n34696) );
  XOR U35584 ( .A(g_input[584]), .B(creg[584]), .Z(n34697) );
  XOR U35585 ( .A(n34698), .B(n34699), .Z(n34689) );
  ANDN U35586 ( .A(n34700), .B(n27242), .Z(n34699) );
  XOR U35587 ( .A(n34701), .B(\modmult_1/zin[0][582] ), .Z(n27242) );
  IV U35588 ( .A(n34698), .Z(n34701) );
  XNOR U35589 ( .A(n34698), .B(n27241), .Z(n34700) );
  XOR U35590 ( .A(n34702), .B(n34703), .Z(n27241) );
  AND U35591 ( .A(\modmult_1/xin[1023] ), .B(n34704), .Z(n34703) );
  IV U35592 ( .A(n34702), .Z(n34704) );
  XOR U35593 ( .A(n34705), .B(g_input[583]), .Z(n34702) );
  NAND U35594 ( .A(n34706), .B(mul_pow), .Z(n34705) );
  XOR U35595 ( .A(g_input[583]), .B(creg[583]), .Z(n34706) );
  XOR U35596 ( .A(n34707), .B(n34708), .Z(n34698) );
  ANDN U35597 ( .A(n34709), .B(n27248), .Z(n34708) );
  XOR U35598 ( .A(n34710), .B(\modmult_1/zin[0][581] ), .Z(n27248) );
  IV U35599 ( .A(n34707), .Z(n34710) );
  XNOR U35600 ( .A(n34707), .B(n27247), .Z(n34709) );
  XOR U35601 ( .A(n34711), .B(n34712), .Z(n27247) );
  AND U35602 ( .A(\modmult_1/xin[1023] ), .B(n34713), .Z(n34712) );
  IV U35603 ( .A(n34711), .Z(n34713) );
  XOR U35604 ( .A(n34714), .B(g_input[582]), .Z(n34711) );
  NAND U35605 ( .A(n34715), .B(mul_pow), .Z(n34714) );
  XOR U35606 ( .A(g_input[582]), .B(creg[582]), .Z(n34715) );
  XOR U35607 ( .A(n34716), .B(n34717), .Z(n34707) );
  ANDN U35608 ( .A(n34718), .B(n27254), .Z(n34717) );
  XOR U35609 ( .A(n34719), .B(\modmult_1/zin[0][580] ), .Z(n27254) );
  IV U35610 ( .A(n34716), .Z(n34719) );
  XNOR U35611 ( .A(n34716), .B(n27253), .Z(n34718) );
  XOR U35612 ( .A(n34720), .B(n34721), .Z(n27253) );
  AND U35613 ( .A(\modmult_1/xin[1023] ), .B(n34722), .Z(n34721) );
  IV U35614 ( .A(n34720), .Z(n34722) );
  XOR U35615 ( .A(n34723), .B(g_input[581]), .Z(n34720) );
  NAND U35616 ( .A(n34724), .B(mul_pow), .Z(n34723) );
  XOR U35617 ( .A(g_input[581]), .B(creg[581]), .Z(n34724) );
  XOR U35618 ( .A(n34725), .B(n34726), .Z(n34716) );
  ANDN U35619 ( .A(n34727), .B(n27260), .Z(n34726) );
  XOR U35620 ( .A(n34728), .B(\modmult_1/zin[0][579] ), .Z(n27260) );
  IV U35621 ( .A(n34725), .Z(n34728) );
  XNOR U35622 ( .A(n34725), .B(n27259), .Z(n34727) );
  XOR U35623 ( .A(n34729), .B(n34730), .Z(n27259) );
  AND U35624 ( .A(\modmult_1/xin[1023] ), .B(n34731), .Z(n34730) );
  IV U35625 ( .A(n34729), .Z(n34731) );
  XOR U35626 ( .A(n34732), .B(g_input[580]), .Z(n34729) );
  NAND U35627 ( .A(n34733), .B(mul_pow), .Z(n34732) );
  XOR U35628 ( .A(g_input[580]), .B(creg[580]), .Z(n34733) );
  XOR U35629 ( .A(n34734), .B(n34735), .Z(n34725) );
  ANDN U35630 ( .A(n34736), .B(n27266), .Z(n34735) );
  XOR U35631 ( .A(n34737), .B(\modmult_1/zin[0][578] ), .Z(n27266) );
  IV U35632 ( .A(n34734), .Z(n34737) );
  XNOR U35633 ( .A(n34734), .B(n27265), .Z(n34736) );
  XOR U35634 ( .A(n34738), .B(n34739), .Z(n27265) );
  AND U35635 ( .A(\modmult_1/xin[1023] ), .B(n34740), .Z(n34739) );
  IV U35636 ( .A(n34738), .Z(n34740) );
  XOR U35637 ( .A(n34741), .B(g_input[579]), .Z(n34738) );
  NAND U35638 ( .A(n34742), .B(mul_pow), .Z(n34741) );
  XOR U35639 ( .A(g_input[579]), .B(creg[579]), .Z(n34742) );
  XOR U35640 ( .A(n34743), .B(n34744), .Z(n34734) );
  ANDN U35641 ( .A(n34745), .B(n27272), .Z(n34744) );
  XOR U35642 ( .A(n34746), .B(\modmult_1/zin[0][577] ), .Z(n27272) );
  IV U35643 ( .A(n34743), .Z(n34746) );
  XNOR U35644 ( .A(n34743), .B(n27271), .Z(n34745) );
  XOR U35645 ( .A(n34747), .B(n34748), .Z(n27271) );
  AND U35646 ( .A(\modmult_1/xin[1023] ), .B(n34749), .Z(n34748) );
  IV U35647 ( .A(n34747), .Z(n34749) );
  XOR U35648 ( .A(n34750), .B(g_input[578]), .Z(n34747) );
  NAND U35649 ( .A(n34751), .B(mul_pow), .Z(n34750) );
  XOR U35650 ( .A(g_input[578]), .B(creg[578]), .Z(n34751) );
  XOR U35651 ( .A(n34752), .B(n34753), .Z(n34743) );
  ANDN U35652 ( .A(n34754), .B(n27278), .Z(n34753) );
  XOR U35653 ( .A(n34755), .B(\modmult_1/zin[0][576] ), .Z(n27278) );
  IV U35654 ( .A(n34752), .Z(n34755) );
  XNOR U35655 ( .A(n34752), .B(n27277), .Z(n34754) );
  XOR U35656 ( .A(n34756), .B(n34757), .Z(n27277) );
  AND U35657 ( .A(\modmult_1/xin[1023] ), .B(n34758), .Z(n34757) );
  IV U35658 ( .A(n34756), .Z(n34758) );
  XOR U35659 ( .A(n34759), .B(g_input[577]), .Z(n34756) );
  NAND U35660 ( .A(n34760), .B(mul_pow), .Z(n34759) );
  XOR U35661 ( .A(g_input[577]), .B(creg[577]), .Z(n34760) );
  XOR U35662 ( .A(n34761), .B(n34762), .Z(n34752) );
  ANDN U35663 ( .A(n34763), .B(n27284), .Z(n34762) );
  XOR U35664 ( .A(n34764), .B(\modmult_1/zin[0][575] ), .Z(n27284) );
  IV U35665 ( .A(n34761), .Z(n34764) );
  XNOR U35666 ( .A(n34761), .B(n27283), .Z(n34763) );
  XOR U35667 ( .A(n34765), .B(n34766), .Z(n27283) );
  AND U35668 ( .A(\modmult_1/xin[1023] ), .B(n34767), .Z(n34766) );
  IV U35669 ( .A(n34765), .Z(n34767) );
  XOR U35670 ( .A(n34768), .B(g_input[576]), .Z(n34765) );
  NAND U35671 ( .A(n34769), .B(mul_pow), .Z(n34768) );
  XOR U35672 ( .A(g_input[576]), .B(creg[576]), .Z(n34769) );
  XOR U35673 ( .A(n34770), .B(n34771), .Z(n34761) );
  ANDN U35674 ( .A(n34772), .B(n27290), .Z(n34771) );
  XOR U35675 ( .A(n34773), .B(\modmult_1/zin[0][574] ), .Z(n27290) );
  IV U35676 ( .A(n34770), .Z(n34773) );
  XNOR U35677 ( .A(n34770), .B(n27289), .Z(n34772) );
  XOR U35678 ( .A(n34774), .B(n34775), .Z(n27289) );
  AND U35679 ( .A(\modmult_1/xin[1023] ), .B(n34776), .Z(n34775) );
  IV U35680 ( .A(n34774), .Z(n34776) );
  XOR U35681 ( .A(n34777), .B(g_input[575]), .Z(n34774) );
  NAND U35682 ( .A(n34778), .B(mul_pow), .Z(n34777) );
  XOR U35683 ( .A(g_input[575]), .B(creg[575]), .Z(n34778) );
  XOR U35684 ( .A(n34779), .B(n34780), .Z(n34770) );
  ANDN U35685 ( .A(n34781), .B(n27296), .Z(n34780) );
  XOR U35686 ( .A(n34782), .B(\modmult_1/zin[0][573] ), .Z(n27296) );
  IV U35687 ( .A(n34779), .Z(n34782) );
  XNOR U35688 ( .A(n34779), .B(n27295), .Z(n34781) );
  XOR U35689 ( .A(n34783), .B(n34784), .Z(n27295) );
  AND U35690 ( .A(\modmult_1/xin[1023] ), .B(n34785), .Z(n34784) );
  IV U35691 ( .A(n34783), .Z(n34785) );
  XOR U35692 ( .A(n34786), .B(g_input[574]), .Z(n34783) );
  NAND U35693 ( .A(n34787), .B(mul_pow), .Z(n34786) );
  XOR U35694 ( .A(g_input[574]), .B(creg[574]), .Z(n34787) );
  XOR U35695 ( .A(n34788), .B(n34789), .Z(n34779) );
  ANDN U35696 ( .A(n34790), .B(n27302), .Z(n34789) );
  XOR U35697 ( .A(n34791), .B(\modmult_1/zin[0][572] ), .Z(n27302) );
  IV U35698 ( .A(n34788), .Z(n34791) );
  XNOR U35699 ( .A(n34788), .B(n27301), .Z(n34790) );
  XOR U35700 ( .A(n34792), .B(n34793), .Z(n27301) );
  AND U35701 ( .A(\modmult_1/xin[1023] ), .B(n34794), .Z(n34793) );
  IV U35702 ( .A(n34792), .Z(n34794) );
  XOR U35703 ( .A(n34795), .B(g_input[573]), .Z(n34792) );
  NAND U35704 ( .A(n34796), .B(mul_pow), .Z(n34795) );
  XOR U35705 ( .A(g_input[573]), .B(creg[573]), .Z(n34796) );
  XOR U35706 ( .A(n34797), .B(n34798), .Z(n34788) );
  ANDN U35707 ( .A(n34799), .B(n27308), .Z(n34798) );
  XOR U35708 ( .A(n34800), .B(\modmult_1/zin[0][571] ), .Z(n27308) );
  IV U35709 ( .A(n34797), .Z(n34800) );
  XNOR U35710 ( .A(n34797), .B(n27307), .Z(n34799) );
  XOR U35711 ( .A(n34801), .B(n34802), .Z(n27307) );
  AND U35712 ( .A(\modmult_1/xin[1023] ), .B(n34803), .Z(n34802) );
  IV U35713 ( .A(n34801), .Z(n34803) );
  XOR U35714 ( .A(n34804), .B(g_input[572]), .Z(n34801) );
  NAND U35715 ( .A(n34805), .B(mul_pow), .Z(n34804) );
  XOR U35716 ( .A(g_input[572]), .B(creg[572]), .Z(n34805) );
  XOR U35717 ( .A(n34806), .B(n34807), .Z(n34797) );
  ANDN U35718 ( .A(n34808), .B(n27314), .Z(n34807) );
  XOR U35719 ( .A(n34809), .B(\modmult_1/zin[0][570] ), .Z(n27314) );
  IV U35720 ( .A(n34806), .Z(n34809) );
  XNOR U35721 ( .A(n34806), .B(n27313), .Z(n34808) );
  XOR U35722 ( .A(n34810), .B(n34811), .Z(n27313) );
  AND U35723 ( .A(\modmult_1/xin[1023] ), .B(n34812), .Z(n34811) );
  IV U35724 ( .A(n34810), .Z(n34812) );
  XOR U35725 ( .A(n34813), .B(g_input[571]), .Z(n34810) );
  NAND U35726 ( .A(n34814), .B(mul_pow), .Z(n34813) );
  XOR U35727 ( .A(g_input[571]), .B(creg[571]), .Z(n34814) );
  XOR U35728 ( .A(n34815), .B(n34816), .Z(n34806) );
  ANDN U35729 ( .A(n34817), .B(n27320), .Z(n34816) );
  XOR U35730 ( .A(n34818), .B(\modmult_1/zin[0][569] ), .Z(n27320) );
  IV U35731 ( .A(n34815), .Z(n34818) );
  XNOR U35732 ( .A(n34815), .B(n27319), .Z(n34817) );
  XOR U35733 ( .A(n34819), .B(n34820), .Z(n27319) );
  AND U35734 ( .A(\modmult_1/xin[1023] ), .B(n34821), .Z(n34820) );
  IV U35735 ( .A(n34819), .Z(n34821) );
  XOR U35736 ( .A(n34822), .B(g_input[570]), .Z(n34819) );
  NAND U35737 ( .A(n34823), .B(mul_pow), .Z(n34822) );
  XOR U35738 ( .A(g_input[570]), .B(creg[570]), .Z(n34823) );
  XOR U35739 ( .A(n34824), .B(n34825), .Z(n34815) );
  ANDN U35740 ( .A(n34826), .B(n27326), .Z(n34825) );
  XOR U35741 ( .A(n34827), .B(\modmult_1/zin[0][568] ), .Z(n27326) );
  IV U35742 ( .A(n34824), .Z(n34827) );
  XNOR U35743 ( .A(n34824), .B(n27325), .Z(n34826) );
  XOR U35744 ( .A(n34828), .B(n34829), .Z(n27325) );
  AND U35745 ( .A(\modmult_1/xin[1023] ), .B(n34830), .Z(n34829) );
  IV U35746 ( .A(n34828), .Z(n34830) );
  XOR U35747 ( .A(n34831), .B(g_input[569]), .Z(n34828) );
  NAND U35748 ( .A(n34832), .B(mul_pow), .Z(n34831) );
  XOR U35749 ( .A(g_input[569]), .B(creg[569]), .Z(n34832) );
  XOR U35750 ( .A(n34833), .B(n34834), .Z(n34824) );
  ANDN U35751 ( .A(n34835), .B(n27332), .Z(n34834) );
  XOR U35752 ( .A(n34836), .B(\modmult_1/zin[0][567] ), .Z(n27332) );
  IV U35753 ( .A(n34833), .Z(n34836) );
  XNOR U35754 ( .A(n34833), .B(n27331), .Z(n34835) );
  XOR U35755 ( .A(n34837), .B(n34838), .Z(n27331) );
  AND U35756 ( .A(\modmult_1/xin[1023] ), .B(n34839), .Z(n34838) );
  IV U35757 ( .A(n34837), .Z(n34839) );
  XOR U35758 ( .A(n34840), .B(g_input[568]), .Z(n34837) );
  NAND U35759 ( .A(n34841), .B(mul_pow), .Z(n34840) );
  XOR U35760 ( .A(g_input[568]), .B(creg[568]), .Z(n34841) );
  XOR U35761 ( .A(n34842), .B(n34843), .Z(n34833) );
  ANDN U35762 ( .A(n34844), .B(n27338), .Z(n34843) );
  XOR U35763 ( .A(n34845), .B(\modmult_1/zin[0][566] ), .Z(n27338) );
  IV U35764 ( .A(n34842), .Z(n34845) );
  XNOR U35765 ( .A(n34842), .B(n27337), .Z(n34844) );
  XOR U35766 ( .A(n34846), .B(n34847), .Z(n27337) );
  AND U35767 ( .A(\modmult_1/xin[1023] ), .B(n34848), .Z(n34847) );
  IV U35768 ( .A(n34846), .Z(n34848) );
  XOR U35769 ( .A(n34849), .B(g_input[567]), .Z(n34846) );
  NAND U35770 ( .A(n34850), .B(mul_pow), .Z(n34849) );
  XOR U35771 ( .A(g_input[567]), .B(creg[567]), .Z(n34850) );
  XOR U35772 ( .A(n34851), .B(n34852), .Z(n34842) );
  ANDN U35773 ( .A(n34853), .B(n27344), .Z(n34852) );
  XOR U35774 ( .A(n34854), .B(\modmult_1/zin[0][565] ), .Z(n27344) );
  IV U35775 ( .A(n34851), .Z(n34854) );
  XNOR U35776 ( .A(n34851), .B(n27343), .Z(n34853) );
  XOR U35777 ( .A(n34855), .B(n34856), .Z(n27343) );
  AND U35778 ( .A(\modmult_1/xin[1023] ), .B(n34857), .Z(n34856) );
  IV U35779 ( .A(n34855), .Z(n34857) );
  XOR U35780 ( .A(n34858), .B(g_input[566]), .Z(n34855) );
  NAND U35781 ( .A(n34859), .B(mul_pow), .Z(n34858) );
  XOR U35782 ( .A(g_input[566]), .B(creg[566]), .Z(n34859) );
  XOR U35783 ( .A(n34860), .B(n34861), .Z(n34851) );
  ANDN U35784 ( .A(n34862), .B(n27350), .Z(n34861) );
  XOR U35785 ( .A(n34863), .B(\modmult_1/zin[0][564] ), .Z(n27350) );
  IV U35786 ( .A(n34860), .Z(n34863) );
  XNOR U35787 ( .A(n34860), .B(n27349), .Z(n34862) );
  XOR U35788 ( .A(n34864), .B(n34865), .Z(n27349) );
  AND U35789 ( .A(\modmult_1/xin[1023] ), .B(n34866), .Z(n34865) );
  IV U35790 ( .A(n34864), .Z(n34866) );
  XOR U35791 ( .A(n34867), .B(g_input[565]), .Z(n34864) );
  NAND U35792 ( .A(n34868), .B(mul_pow), .Z(n34867) );
  XOR U35793 ( .A(g_input[565]), .B(creg[565]), .Z(n34868) );
  XOR U35794 ( .A(n34869), .B(n34870), .Z(n34860) );
  ANDN U35795 ( .A(n34871), .B(n27356), .Z(n34870) );
  XOR U35796 ( .A(n34872), .B(\modmult_1/zin[0][563] ), .Z(n27356) );
  IV U35797 ( .A(n34869), .Z(n34872) );
  XNOR U35798 ( .A(n34869), .B(n27355), .Z(n34871) );
  XOR U35799 ( .A(n34873), .B(n34874), .Z(n27355) );
  AND U35800 ( .A(\modmult_1/xin[1023] ), .B(n34875), .Z(n34874) );
  IV U35801 ( .A(n34873), .Z(n34875) );
  XOR U35802 ( .A(n34876), .B(g_input[564]), .Z(n34873) );
  NAND U35803 ( .A(n34877), .B(mul_pow), .Z(n34876) );
  XOR U35804 ( .A(g_input[564]), .B(creg[564]), .Z(n34877) );
  XOR U35805 ( .A(n34878), .B(n34879), .Z(n34869) );
  ANDN U35806 ( .A(n34880), .B(n27362), .Z(n34879) );
  XOR U35807 ( .A(n34881), .B(\modmult_1/zin[0][562] ), .Z(n27362) );
  IV U35808 ( .A(n34878), .Z(n34881) );
  XNOR U35809 ( .A(n34878), .B(n27361), .Z(n34880) );
  XOR U35810 ( .A(n34882), .B(n34883), .Z(n27361) );
  AND U35811 ( .A(\modmult_1/xin[1023] ), .B(n34884), .Z(n34883) );
  IV U35812 ( .A(n34882), .Z(n34884) );
  XOR U35813 ( .A(n34885), .B(g_input[563]), .Z(n34882) );
  NAND U35814 ( .A(n34886), .B(mul_pow), .Z(n34885) );
  XOR U35815 ( .A(g_input[563]), .B(creg[563]), .Z(n34886) );
  XOR U35816 ( .A(n34887), .B(n34888), .Z(n34878) );
  ANDN U35817 ( .A(n34889), .B(n27368), .Z(n34888) );
  XOR U35818 ( .A(n34890), .B(\modmult_1/zin[0][561] ), .Z(n27368) );
  IV U35819 ( .A(n34887), .Z(n34890) );
  XNOR U35820 ( .A(n34887), .B(n27367), .Z(n34889) );
  XOR U35821 ( .A(n34891), .B(n34892), .Z(n27367) );
  AND U35822 ( .A(\modmult_1/xin[1023] ), .B(n34893), .Z(n34892) );
  IV U35823 ( .A(n34891), .Z(n34893) );
  XOR U35824 ( .A(n34894), .B(g_input[562]), .Z(n34891) );
  NAND U35825 ( .A(n34895), .B(mul_pow), .Z(n34894) );
  XOR U35826 ( .A(g_input[562]), .B(creg[562]), .Z(n34895) );
  XOR U35827 ( .A(n34896), .B(n34897), .Z(n34887) );
  ANDN U35828 ( .A(n34898), .B(n27374), .Z(n34897) );
  XOR U35829 ( .A(n34899), .B(\modmult_1/zin[0][560] ), .Z(n27374) );
  IV U35830 ( .A(n34896), .Z(n34899) );
  XNOR U35831 ( .A(n34896), .B(n27373), .Z(n34898) );
  XOR U35832 ( .A(n34900), .B(n34901), .Z(n27373) );
  AND U35833 ( .A(\modmult_1/xin[1023] ), .B(n34902), .Z(n34901) );
  IV U35834 ( .A(n34900), .Z(n34902) );
  XOR U35835 ( .A(n34903), .B(g_input[561]), .Z(n34900) );
  NAND U35836 ( .A(n34904), .B(mul_pow), .Z(n34903) );
  XOR U35837 ( .A(g_input[561]), .B(creg[561]), .Z(n34904) );
  XOR U35838 ( .A(n34905), .B(n34906), .Z(n34896) );
  ANDN U35839 ( .A(n34907), .B(n27380), .Z(n34906) );
  XOR U35840 ( .A(n34908), .B(\modmult_1/zin[0][559] ), .Z(n27380) );
  IV U35841 ( .A(n34905), .Z(n34908) );
  XNOR U35842 ( .A(n34905), .B(n27379), .Z(n34907) );
  XOR U35843 ( .A(n34909), .B(n34910), .Z(n27379) );
  AND U35844 ( .A(\modmult_1/xin[1023] ), .B(n34911), .Z(n34910) );
  IV U35845 ( .A(n34909), .Z(n34911) );
  XOR U35846 ( .A(n34912), .B(g_input[560]), .Z(n34909) );
  NAND U35847 ( .A(n34913), .B(mul_pow), .Z(n34912) );
  XOR U35848 ( .A(g_input[560]), .B(creg[560]), .Z(n34913) );
  XOR U35849 ( .A(n34914), .B(n34915), .Z(n34905) );
  ANDN U35850 ( .A(n34916), .B(n27386), .Z(n34915) );
  XOR U35851 ( .A(n34917), .B(\modmult_1/zin[0][558] ), .Z(n27386) );
  IV U35852 ( .A(n34914), .Z(n34917) );
  XNOR U35853 ( .A(n34914), .B(n27385), .Z(n34916) );
  XOR U35854 ( .A(n34918), .B(n34919), .Z(n27385) );
  AND U35855 ( .A(\modmult_1/xin[1023] ), .B(n34920), .Z(n34919) );
  IV U35856 ( .A(n34918), .Z(n34920) );
  XOR U35857 ( .A(n34921), .B(g_input[559]), .Z(n34918) );
  NAND U35858 ( .A(n34922), .B(mul_pow), .Z(n34921) );
  XOR U35859 ( .A(g_input[559]), .B(creg[559]), .Z(n34922) );
  XOR U35860 ( .A(n34923), .B(n34924), .Z(n34914) );
  ANDN U35861 ( .A(n34925), .B(n27392), .Z(n34924) );
  XOR U35862 ( .A(n34926), .B(\modmult_1/zin[0][557] ), .Z(n27392) );
  IV U35863 ( .A(n34923), .Z(n34926) );
  XNOR U35864 ( .A(n34923), .B(n27391), .Z(n34925) );
  XOR U35865 ( .A(n34927), .B(n34928), .Z(n27391) );
  AND U35866 ( .A(\modmult_1/xin[1023] ), .B(n34929), .Z(n34928) );
  IV U35867 ( .A(n34927), .Z(n34929) );
  XOR U35868 ( .A(n34930), .B(g_input[558]), .Z(n34927) );
  NAND U35869 ( .A(n34931), .B(mul_pow), .Z(n34930) );
  XOR U35870 ( .A(g_input[558]), .B(creg[558]), .Z(n34931) );
  XOR U35871 ( .A(n34932), .B(n34933), .Z(n34923) );
  ANDN U35872 ( .A(n34934), .B(n27398), .Z(n34933) );
  XOR U35873 ( .A(n34935), .B(\modmult_1/zin[0][556] ), .Z(n27398) );
  IV U35874 ( .A(n34932), .Z(n34935) );
  XNOR U35875 ( .A(n34932), .B(n27397), .Z(n34934) );
  XOR U35876 ( .A(n34936), .B(n34937), .Z(n27397) );
  AND U35877 ( .A(\modmult_1/xin[1023] ), .B(n34938), .Z(n34937) );
  IV U35878 ( .A(n34936), .Z(n34938) );
  XOR U35879 ( .A(n34939), .B(g_input[557]), .Z(n34936) );
  NAND U35880 ( .A(n34940), .B(mul_pow), .Z(n34939) );
  XOR U35881 ( .A(g_input[557]), .B(creg[557]), .Z(n34940) );
  XOR U35882 ( .A(n34941), .B(n34942), .Z(n34932) );
  ANDN U35883 ( .A(n34943), .B(n27404), .Z(n34942) );
  XOR U35884 ( .A(n34944), .B(\modmult_1/zin[0][555] ), .Z(n27404) );
  IV U35885 ( .A(n34941), .Z(n34944) );
  XNOR U35886 ( .A(n34941), .B(n27403), .Z(n34943) );
  XOR U35887 ( .A(n34945), .B(n34946), .Z(n27403) );
  AND U35888 ( .A(\modmult_1/xin[1023] ), .B(n34947), .Z(n34946) );
  IV U35889 ( .A(n34945), .Z(n34947) );
  XOR U35890 ( .A(n34948), .B(g_input[556]), .Z(n34945) );
  NAND U35891 ( .A(n34949), .B(mul_pow), .Z(n34948) );
  XOR U35892 ( .A(g_input[556]), .B(creg[556]), .Z(n34949) );
  XOR U35893 ( .A(n34950), .B(n34951), .Z(n34941) );
  ANDN U35894 ( .A(n34952), .B(n27410), .Z(n34951) );
  XOR U35895 ( .A(n34953), .B(\modmult_1/zin[0][554] ), .Z(n27410) );
  IV U35896 ( .A(n34950), .Z(n34953) );
  XNOR U35897 ( .A(n34950), .B(n27409), .Z(n34952) );
  XOR U35898 ( .A(n34954), .B(n34955), .Z(n27409) );
  AND U35899 ( .A(\modmult_1/xin[1023] ), .B(n34956), .Z(n34955) );
  IV U35900 ( .A(n34954), .Z(n34956) );
  XOR U35901 ( .A(n34957), .B(g_input[555]), .Z(n34954) );
  NAND U35902 ( .A(n34958), .B(mul_pow), .Z(n34957) );
  XOR U35903 ( .A(g_input[555]), .B(creg[555]), .Z(n34958) );
  XOR U35904 ( .A(n34959), .B(n34960), .Z(n34950) );
  ANDN U35905 ( .A(n34961), .B(n27416), .Z(n34960) );
  XOR U35906 ( .A(n34962), .B(\modmult_1/zin[0][553] ), .Z(n27416) );
  IV U35907 ( .A(n34959), .Z(n34962) );
  XNOR U35908 ( .A(n34959), .B(n27415), .Z(n34961) );
  XOR U35909 ( .A(n34963), .B(n34964), .Z(n27415) );
  AND U35910 ( .A(\modmult_1/xin[1023] ), .B(n34965), .Z(n34964) );
  IV U35911 ( .A(n34963), .Z(n34965) );
  XOR U35912 ( .A(n34966), .B(g_input[554]), .Z(n34963) );
  NAND U35913 ( .A(n34967), .B(mul_pow), .Z(n34966) );
  XOR U35914 ( .A(g_input[554]), .B(creg[554]), .Z(n34967) );
  XOR U35915 ( .A(n34968), .B(n34969), .Z(n34959) );
  ANDN U35916 ( .A(n34970), .B(n27422), .Z(n34969) );
  XOR U35917 ( .A(n34971), .B(\modmult_1/zin[0][552] ), .Z(n27422) );
  IV U35918 ( .A(n34968), .Z(n34971) );
  XNOR U35919 ( .A(n34968), .B(n27421), .Z(n34970) );
  XOR U35920 ( .A(n34972), .B(n34973), .Z(n27421) );
  AND U35921 ( .A(\modmult_1/xin[1023] ), .B(n34974), .Z(n34973) );
  IV U35922 ( .A(n34972), .Z(n34974) );
  XOR U35923 ( .A(n34975), .B(g_input[553]), .Z(n34972) );
  NAND U35924 ( .A(n34976), .B(mul_pow), .Z(n34975) );
  XOR U35925 ( .A(g_input[553]), .B(creg[553]), .Z(n34976) );
  XOR U35926 ( .A(n34977), .B(n34978), .Z(n34968) );
  ANDN U35927 ( .A(n34979), .B(n27428), .Z(n34978) );
  XOR U35928 ( .A(n34980), .B(\modmult_1/zin[0][551] ), .Z(n27428) );
  IV U35929 ( .A(n34977), .Z(n34980) );
  XNOR U35930 ( .A(n34977), .B(n27427), .Z(n34979) );
  XOR U35931 ( .A(n34981), .B(n34982), .Z(n27427) );
  AND U35932 ( .A(\modmult_1/xin[1023] ), .B(n34983), .Z(n34982) );
  IV U35933 ( .A(n34981), .Z(n34983) );
  XOR U35934 ( .A(n34984), .B(g_input[552]), .Z(n34981) );
  NAND U35935 ( .A(n34985), .B(mul_pow), .Z(n34984) );
  XOR U35936 ( .A(g_input[552]), .B(creg[552]), .Z(n34985) );
  XOR U35937 ( .A(n34986), .B(n34987), .Z(n34977) );
  ANDN U35938 ( .A(n34988), .B(n27434), .Z(n34987) );
  XOR U35939 ( .A(n34989), .B(\modmult_1/zin[0][550] ), .Z(n27434) );
  IV U35940 ( .A(n34986), .Z(n34989) );
  XNOR U35941 ( .A(n34986), .B(n27433), .Z(n34988) );
  XOR U35942 ( .A(n34990), .B(n34991), .Z(n27433) );
  AND U35943 ( .A(\modmult_1/xin[1023] ), .B(n34992), .Z(n34991) );
  IV U35944 ( .A(n34990), .Z(n34992) );
  XOR U35945 ( .A(n34993), .B(g_input[551]), .Z(n34990) );
  NAND U35946 ( .A(n34994), .B(mul_pow), .Z(n34993) );
  XOR U35947 ( .A(g_input[551]), .B(creg[551]), .Z(n34994) );
  XOR U35948 ( .A(n34995), .B(n34996), .Z(n34986) );
  ANDN U35949 ( .A(n34997), .B(n27440), .Z(n34996) );
  XOR U35950 ( .A(n34998), .B(\modmult_1/zin[0][549] ), .Z(n27440) );
  IV U35951 ( .A(n34995), .Z(n34998) );
  XNOR U35952 ( .A(n34995), .B(n27439), .Z(n34997) );
  XOR U35953 ( .A(n34999), .B(n35000), .Z(n27439) );
  AND U35954 ( .A(\modmult_1/xin[1023] ), .B(n35001), .Z(n35000) );
  IV U35955 ( .A(n34999), .Z(n35001) );
  XOR U35956 ( .A(n35002), .B(g_input[550]), .Z(n34999) );
  NAND U35957 ( .A(n35003), .B(mul_pow), .Z(n35002) );
  XOR U35958 ( .A(g_input[550]), .B(creg[550]), .Z(n35003) );
  XOR U35959 ( .A(n35004), .B(n35005), .Z(n34995) );
  ANDN U35960 ( .A(n35006), .B(n27446), .Z(n35005) );
  XOR U35961 ( .A(n35007), .B(\modmult_1/zin[0][548] ), .Z(n27446) );
  IV U35962 ( .A(n35004), .Z(n35007) );
  XNOR U35963 ( .A(n35004), .B(n27445), .Z(n35006) );
  XOR U35964 ( .A(n35008), .B(n35009), .Z(n27445) );
  AND U35965 ( .A(\modmult_1/xin[1023] ), .B(n35010), .Z(n35009) );
  IV U35966 ( .A(n35008), .Z(n35010) );
  XOR U35967 ( .A(n35011), .B(g_input[549]), .Z(n35008) );
  NAND U35968 ( .A(n35012), .B(mul_pow), .Z(n35011) );
  XOR U35969 ( .A(g_input[549]), .B(creg[549]), .Z(n35012) );
  XOR U35970 ( .A(n35013), .B(n35014), .Z(n35004) );
  ANDN U35971 ( .A(n35015), .B(n27452), .Z(n35014) );
  XOR U35972 ( .A(n35016), .B(\modmult_1/zin[0][547] ), .Z(n27452) );
  IV U35973 ( .A(n35013), .Z(n35016) );
  XNOR U35974 ( .A(n35013), .B(n27451), .Z(n35015) );
  XOR U35975 ( .A(n35017), .B(n35018), .Z(n27451) );
  AND U35976 ( .A(\modmult_1/xin[1023] ), .B(n35019), .Z(n35018) );
  IV U35977 ( .A(n35017), .Z(n35019) );
  XOR U35978 ( .A(n35020), .B(g_input[548]), .Z(n35017) );
  NAND U35979 ( .A(n35021), .B(mul_pow), .Z(n35020) );
  XOR U35980 ( .A(g_input[548]), .B(creg[548]), .Z(n35021) );
  XOR U35981 ( .A(n35022), .B(n35023), .Z(n35013) );
  ANDN U35982 ( .A(n35024), .B(n27458), .Z(n35023) );
  XOR U35983 ( .A(n35025), .B(\modmult_1/zin[0][546] ), .Z(n27458) );
  IV U35984 ( .A(n35022), .Z(n35025) );
  XNOR U35985 ( .A(n35022), .B(n27457), .Z(n35024) );
  XOR U35986 ( .A(n35026), .B(n35027), .Z(n27457) );
  AND U35987 ( .A(\modmult_1/xin[1023] ), .B(n35028), .Z(n35027) );
  IV U35988 ( .A(n35026), .Z(n35028) );
  XOR U35989 ( .A(n35029), .B(g_input[547]), .Z(n35026) );
  NAND U35990 ( .A(n35030), .B(mul_pow), .Z(n35029) );
  XOR U35991 ( .A(g_input[547]), .B(creg[547]), .Z(n35030) );
  XOR U35992 ( .A(n35031), .B(n35032), .Z(n35022) );
  ANDN U35993 ( .A(n35033), .B(n27464), .Z(n35032) );
  XOR U35994 ( .A(n35034), .B(\modmult_1/zin[0][545] ), .Z(n27464) );
  IV U35995 ( .A(n35031), .Z(n35034) );
  XNOR U35996 ( .A(n35031), .B(n27463), .Z(n35033) );
  XOR U35997 ( .A(n35035), .B(n35036), .Z(n27463) );
  AND U35998 ( .A(\modmult_1/xin[1023] ), .B(n35037), .Z(n35036) );
  IV U35999 ( .A(n35035), .Z(n35037) );
  XOR U36000 ( .A(n35038), .B(g_input[546]), .Z(n35035) );
  NAND U36001 ( .A(n35039), .B(mul_pow), .Z(n35038) );
  XOR U36002 ( .A(g_input[546]), .B(creg[546]), .Z(n35039) );
  XOR U36003 ( .A(n35040), .B(n35041), .Z(n35031) );
  ANDN U36004 ( .A(n35042), .B(n27470), .Z(n35041) );
  XOR U36005 ( .A(n35043), .B(\modmult_1/zin[0][544] ), .Z(n27470) );
  IV U36006 ( .A(n35040), .Z(n35043) );
  XNOR U36007 ( .A(n35040), .B(n27469), .Z(n35042) );
  XOR U36008 ( .A(n35044), .B(n35045), .Z(n27469) );
  AND U36009 ( .A(\modmult_1/xin[1023] ), .B(n35046), .Z(n35045) );
  IV U36010 ( .A(n35044), .Z(n35046) );
  XOR U36011 ( .A(n35047), .B(g_input[545]), .Z(n35044) );
  NAND U36012 ( .A(n35048), .B(mul_pow), .Z(n35047) );
  XOR U36013 ( .A(g_input[545]), .B(creg[545]), .Z(n35048) );
  XOR U36014 ( .A(n35049), .B(n35050), .Z(n35040) );
  ANDN U36015 ( .A(n35051), .B(n27476), .Z(n35050) );
  XOR U36016 ( .A(n35052), .B(\modmult_1/zin[0][543] ), .Z(n27476) );
  IV U36017 ( .A(n35049), .Z(n35052) );
  XNOR U36018 ( .A(n35049), .B(n27475), .Z(n35051) );
  XOR U36019 ( .A(n35053), .B(n35054), .Z(n27475) );
  AND U36020 ( .A(\modmult_1/xin[1023] ), .B(n35055), .Z(n35054) );
  IV U36021 ( .A(n35053), .Z(n35055) );
  XOR U36022 ( .A(n35056), .B(g_input[544]), .Z(n35053) );
  NAND U36023 ( .A(n35057), .B(mul_pow), .Z(n35056) );
  XOR U36024 ( .A(g_input[544]), .B(creg[544]), .Z(n35057) );
  XOR U36025 ( .A(n35058), .B(n35059), .Z(n35049) );
  ANDN U36026 ( .A(n35060), .B(n27482), .Z(n35059) );
  XOR U36027 ( .A(n35061), .B(\modmult_1/zin[0][542] ), .Z(n27482) );
  IV U36028 ( .A(n35058), .Z(n35061) );
  XNOR U36029 ( .A(n35058), .B(n27481), .Z(n35060) );
  XOR U36030 ( .A(n35062), .B(n35063), .Z(n27481) );
  AND U36031 ( .A(\modmult_1/xin[1023] ), .B(n35064), .Z(n35063) );
  IV U36032 ( .A(n35062), .Z(n35064) );
  XOR U36033 ( .A(n35065), .B(g_input[543]), .Z(n35062) );
  NAND U36034 ( .A(n35066), .B(mul_pow), .Z(n35065) );
  XOR U36035 ( .A(g_input[543]), .B(creg[543]), .Z(n35066) );
  XOR U36036 ( .A(n35067), .B(n35068), .Z(n35058) );
  ANDN U36037 ( .A(n35069), .B(n27488), .Z(n35068) );
  XOR U36038 ( .A(n35070), .B(\modmult_1/zin[0][541] ), .Z(n27488) );
  IV U36039 ( .A(n35067), .Z(n35070) );
  XNOR U36040 ( .A(n35067), .B(n27487), .Z(n35069) );
  XOR U36041 ( .A(n35071), .B(n35072), .Z(n27487) );
  AND U36042 ( .A(\modmult_1/xin[1023] ), .B(n35073), .Z(n35072) );
  IV U36043 ( .A(n35071), .Z(n35073) );
  XOR U36044 ( .A(n35074), .B(g_input[542]), .Z(n35071) );
  NAND U36045 ( .A(n35075), .B(mul_pow), .Z(n35074) );
  XOR U36046 ( .A(g_input[542]), .B(creg[542]), .Z(n35075) );
  XOR U36047 ( .A(n35076), .B(n35077), .Z(n35067) );
  ANDN U36048 ( .A(n35078), .B(n27494), .Z(n35077) );
  XOR U36049 ( .A(n35079), .B(\modmult_1/zin[0][540] ), .Z(n27494) );
  IV U36050 ( .A(n35076), .Z(n35079) );
  XNOR U36051 ( .A(n35076), .B(n27493), .Z(n35078) );
  XOR U36052 ( .A(n35080), .B(n35081), .Z(n27493) );
  AND U36053 ( .A(\modmult_1/xin[1023] ), .B(n35082), .Z(n35081) );
  IV U36054 ( .A(n35080), .Z(n35082) );
  XOR U36055 ( .A(n35083), .B(g_input[541]), .Z(n35080) );
  NAND U36056 ( .A(n35084), .B(mul_pow), .Z(n35083) );
  XOR U36057 ( .A(g_input[541]), .B(creg[541]), .Z(n35084) );
  XOR U36058 ( .A(n35085), .B(n35086), .Z(n35076) );
  ANDN U36059 ( .A(n35087), .B(n27500), .Z(n35086) );
  XOR U36060 ( .A(n35088), .B(\modmult_1/zin[0][539] ), .Z(n27500) );
  IV U36061 ( .A(n35085), .Z(n35088) );
  XNOR U36062 ( .A(n35085), .B(n27499), .Z(n35087) );
  XOR U36063 ( .A(n35089), .B(n35090), .Z(n27499) );
  AND U36064 ( .A(\modmult_1/xin[1023] ), .B(n35091), .Z(n35090) );
  IV U36065 ( .A(n35089), .Z(n35091) );
  XOR U36066 ( .A(n35092), .B(g_input[540]), .Z(n35089) );
  NAND U36067 ( .A(n35093), .B(mul_pow), .Z(n35092) );
  XOR U36068 ( .A(g_input[540]), .B(creg[540]), .Z(n35093) );
  XOR U36069 ( .A(n35094), .B(n35095), .Z(n35085) );
  ANDN U36070 ( .A(n35096), .B(n27506), .Z(n35095) );
  XOR U36071 ( .A(n35097), .B(\modmult_1/zin[0][538] ), .Z(n27506) );
  IV U36072 ( .A(n35094), .Z(n35097) );
  XNOR U36073 ( .A(n35094), .B(n27505), .Z(n35096) );
  XOR U36074 ( .A(n35098), .B(n35099), .Z(n27505) );
  AND U36075 ( .A(\modmult_1/xin[1023] ), .B(n35100), .Z(n35099) );
  IV U36076 ( .A(n35098), .Z(n35100) );
  XOR U36077 ( .A(n35101), .B(g_input[539]), .Z(n35098) );
  NAND U36078 ( .A(n35102), .B(mul_pow), .Z(n35101) );
  XOR U36079 ( .A(g_input[539]), .B(creg[539]), .Z(n35102) );
  XOR U36080 ( .A(n35103), .B(n35104), .Z(n35094) );
  ANDN U36081 ( .A(n35105), .B(n27512), .Z(n35104) );
  XOR U36082 ( .A(n35106), .B(\modmult_1/zin[0][537] ), .Z(n27512) );
  IV U36083 ( .A(n35103), .Z(n35106) );
  XNOR U36084 ( .A(n35103), .B(n27511), .Z(n35105) );
  XOR U36085 ( .A(n35107), .B(n35108), .Z(n27511) );
  AND U36086 ( .A(\modmult_1/xin[1023] ), .B(n35109), .Z(n35108) );
  IV U36087 ( .A(n35107), .Z(n35109) );
  XOR U36088 ( .A(n35110), .B(g_input[538]), .Z(n35107) );
  NAND U36089 ( .A(n35111), .B(mul_pow), .Z(n35110) );
  XOR U36090 ( .A(g_input[538]), .B(creg[538]), .Z(n35111) );
  XOR U36091 ( .A(n35112), .B(n35113), .Z(n35103) );
  ANDN U36092 ( .A(n35114), .B(n27518), .Z(n35113) );
  XOR U36093 ( .A(n35115), .B(\modmult_1/zin[0][536] ), .Z(n27518) );
  IV U36094 ( .A(n35112), .Z(n35115) );
  XNOR U36095 ( .A(n35112), .B(n27517), .Z(n35114) );
  XOR U36096 ( .A(n35116), .B(n35117), .Z(n27517) );
  AND U36097 ( .A(\modmult_1/xin[1023] ), .B(n35118), .Z(n35117) );
  IV U36098 ( .A(n35116), .Z(n35118) );
  XOR U36099 ( .A(n35119), .B(g_input[537]), .Z(n35116) );
  NAND U36100 ( .A(n35120), .B(mul_pow), .Z(n35119) );
  XOR U36101 ( .A(g_input[537]), .B(creg[537]), .Z(n35120) );
  XOR U36102 ( .A(n35121), .B(n35122), .Z(n35112) );
  ANDN U36103 ( .A(n35123), .B(n27524), .Z(n35122) );
  XOR U36104 ( .A(n35124), .B(\modmult_1/zin[0][535] ), .Z(n27524) );
  IV U36105 ( .A(n35121), .Z(n35124) );
  XNOR U36106 ( .A(n35121), .B(n27523), .Z(n35123) );
  XOR U36107 ( .A(n35125), .B(n35126), .Z(n27523) );
  AND U36108 ( .A(\modmult_1/xin[1023] ), .B(n35127), .Z(n35126) );
  IV U36109 ( .A(n35125), .Z(n35127) );
  XOR U36110 ( .A(n35128), .B(g_input[536]), .Z(n35125) );
  NAND U36111 ( .A(n35129), .B(mul_pow), .Z(n35128) );
  XOR U36112 ( .A(g_input[536]), .B(creg[536]), .Z(n35129) );
  XOR U36113 ( .A(n35130), .B(n35131), .Z(n35121) );
  ANDN U36114 ( .A(n35132), .B(n27530), .Z(n35131) );
  XOR U36115 ( .A(n35133), .B(\modmult_1/zin[0][534] ), .Z(n27530) );
  IV U36116 ( .A(n35130), .Z(n35133) );
  XNOR U36117 ( .A(n35130), .B(n27529), .Z(n35132) );
  XOR U36118 ( .A(n35134), .B(n35135), .Z(n27529) );
  AND U36119 ( .A(\modmult_1/xin[1023] ), .B(n35136), .Z(n35135) );
  IV U36120 ( .A(n35134), .Z(n35136) );
  XOR U36121 ( .A(n35137), .B(g_input[535]), .Z(n35134) );
  NAND U36122 ( .A(n35138), .B(mul_pow), .Z(n35137) );
  XOR U36123 ( .A(g_input[535]), .B(creg[535]), .Z(n35138) );
  XOR U36124 ( .A(n35139), .B(n35140), .Z(n35130) );
  ANDN U36125 ( .A(n35141), .B(n27536), .Z(n35140) );
  XOR U36126 ( .A(n35142), .B(\modmult_1/zin[0][533] ), .Z(n27536) );
  IV U36127 ( .A(n35139), .Z(n35142) );
  XNOR U36128 ( .A(n35139), .B(n27535), .Z(n35141) );
  XOR U36129 ( .A(n35143), .B(n35144), .Z(n27535) );
  AND U36130 ( .A(\modmult_1/xin[1023] ), .B(n35145), .Z(n35144) );
  IV U36131 ( .A(n35143), .Z(n35145) );
  XOR U36132 ( .A(n35146), .B(g_input[534]), .Z(n35143) );
  NAND U36133 ( .A(n35147), .B(mul_pow), .Z(n35146) );
  XOR U36134 ( .A(g_input[534]), .B(creg[534]), .Z(n35147) );
  XOR U36135 ( .A(n35148), .B(n35149), .Z(n35139) );
  ANDN U36136 ( .A(n35150), .B(n27542), .Z(n35149) );
  XOR U36137 ( .A(n35151), .B(\modmult_1/zin[0][532] ), .Z(n27542) );
  IV U36138 ( .A(n35148), .Z(n35151) );
  XNOR U36139 ( .A(n35148), .B(n27541), .Z(n35150) );
  XOR U36140 ( .A(n35152), .B(n35153), .Z(n27541) );
  AND U36141 ( .A(\modmult_1/xin[1023] ), .B(n35154), .Z(n35153) );
  IV U36142 ( .A(n35152), .Z(n35154) );
  XOR U36143 ( .A(n35155), .B(g_input[533]), .Z(n35152) );
  NAND U36144 ( .A(n35156), .B(mul_pow), .Z(n35155) );
  XOR U36145 ( .A(g_input[533]), .B(creg[533]), .Z(n35156) );
  XOR U36146 ( .A(n35157), .B(n35158), .Z(n35148) );
  ANDN U36147 ( .A(n35159), .B(n27548), .Z(n35158) );
  XOR U36148 ( .A(n35160), .B(\modmult_1/zin[0][531] ), .Z(n27548) );
  IV U36149 ( .A(n35157), .Z(n35160) );
  XNOR U36150 ( .A(n35157), .B(n27547), .Z(n35159) );
  XOR U36151 ( .A(n35161), .B(n35162), .Z(n27547) );
  AND U36152 ( .A(\modmult_1/xin[1023] ), .B(n35163), .Z(n35162) );
  IV U36153 ( .A(n35161), .Z(n35163) );
  XOR U36154 ( .A(n35164), .B(g_input[532]), .Z(n35161) );
  NAND U36155 ( .A(n35165), .B(mul_pow), .Z(n35164) );
  XOR U36156 ( .A(g_input[532]), .B(creg[532]), .Z(n35165) );
  XOR U36157 ( .A(n35166), .B(n35167), .Z(n35157) );
  ANDN U36158 ( .A(n35168), .B(n27554), .Z(n35167) );
  XOR U36159 ( .A(n35169), .B(\modmult_1/zin[0][530] ), .Z(n27554) );
  IV U36160 ( .A(n35166), .Z(n35169) );
  XNOR U36161 ( .A(n35166), .B(n27553), .Z(n35168) );
  XOR U36162 ( .A(n35170), .B(n35171), .Z(n27553) );
  AND U36163 ( .A(\modmult_1/xin[1023] ), .B(n35172), .Z(n35171) );
  IV U36164 ( .A(n35170), .Z(n35172) );
  XOR U36165 ( .A(n35173), .B(g_input[531]), .Z(n35170) );
  NAND U36166 ( .A(n35174), .B(mul_pow), .Z(n35173) );
  XOR U36167 ( .A(g_input[531]), .B(creg[531]), .Z(n35174) );
  XOR U36168 ( .A(n35175), .B(n35176), .Z(n35166) );
  ANDN U36169 ( .A(n35177), .B(n27560), .Z(n35176) );
  XOR U36170 ( .A(n35178), .B(\modmult_1/zin[0][529] ), .Z(n27560) );
  IV U36171 ( .A(n35175), .Z(n35178) );
  XNOR U36172 ( .A(n35175), .B(n27559), .Z(n35177) );
  XOR U36173 ( .A(n35179), .B(n35180), .Z(n27559) );
  AND U36174 ( .A(\modmult_1/xin[1023] ), .B(n35181), .Z(n35180) );
  IV U36175 ( .A(n35179), .Z(n35181) );
  XOR U36176 ( .A(n35182), .B(g_input[530]), .Z(n35179) );
  NAND U36177 ( .A(n35183), .B(mul_pow), .Z(n35182) );
  XOR U36178 ( .A(g_input[530]), .B(creg[530]), .Z(n35183) );
  XOR U36179 ( .A(n35184), .B(n35185), .Z(n35175) );
  ANDN U36180 ( .A(n35186), .B(n27566), .Z(n35185) );
  XOR U36181 ( .A(n35187), .B(\modmult_1/zin[0][528] ), .Z(n27566) );
  IV U36182 ( .A(n35184), .Z(n35187) );
  XNOR U36183 ( .A(n35184), .B(n27565), .Z(n35186) );
  XOR U36184 ( .A(n35188), .B(n35189), .Z(n27565) );
  AND U36185 ( .A(\modmult_1/xin[1023] ), .B(n35190), .Z(n35189) );
  IV U36186 ( .A(n35188), .Z(n35190) );
  XOR U36187 ( .A(n35191), .B(g_input[529]), .Z(n35188) );
  NAND U36188 ( .A(n35192), .B(mul_pow), .Z(n35191) );
  XOR U36189 ( .A(g_input[529]), .B(creg[529]), .Z(n35192) );
  XOR U36190 ( .A(n35193), .B(n35194), .Z(n35184) );
  ANDN U36191 ( .A(n35195), .B(n27572), .Z(n35194) );
  XOR U36192 ( .A(n35196), .B(\modmult_1/zin[0][527] ), .Z(n27572) );
  IV U36193 ( .A(n35193), .Z(n35196) );
  XNOR U36194 ( .A(n35193), .B(n27571), .Z(n35195) );
  XOR U36195 ( .A(n35197), .B(n35198), .Z(n27571) );
  AND U36196 ( .A(\modmult_1/xin[1023] ), .B(n35199), .Z(n35198) );
  IV U36197 ( .A(n35197), .Z(n35199) );
  XOR U36198 ( .A(n35200), .B(g_input[528]), .Z(n35197) );
  NAND U36199 ( .A(n35201), .B(mul_pow), .Z(n35200) );
  XOR U36200 ( .A(g_input[528]), .B(creg[528]), .Z(n35201) );
  XOR U36201 ( .A(n35202), .B(n35203), .Z(n35193) );
  ANDN U36202 ( .A(n35204), .B(n27578), .Z(n35203) );
  XOR U36203 ( .A(n35205), .B(\modmult_1/zin[0][526] ), .Z(n27578) );
  IV U36204 ( .A(n35202), .Z(n35205) );
  XNOR U36205 ( .A(n35202), .B(n27577), .Z(n35204) );
  XOR U36206 ( .A(n35206), .B(n35207), .Z(n27577) );
  AND U36207 ( .A(\modmult_1/xin[1023] ), .B(n35208), .Z(n35207) );
  IV U36208 ( .A(n35206), .Z(n35208) );
  XOR U36209 ( .A(n35209), .B(g_input[527]), .Z(n35206) );
  NAND U36210 ( .A(n35210), .B(mul_pow), .Z(n35209) );
  XOR U36211 ( .A(g_input[527]), .B(creg[527]), .Z(n35210) );
  XOR U36212 ( .A(n35211), .B(n35212), .Z(n35202) );
  ANDN U36213 ( .A(n35213), .B(n27584), .Z(n35212) );
  XOR U36214 ( .A(n35214), .B(\modmult_1/zin[0][525] ), .Z(n27584) );
  IV U36215 ( .A(n35211), .Z(n35214) );
  XNOR U36216 ( .A(n35211), .B(n27583), .Z(n35213) );
  XOR U36217 ( .A(n35215), .B(n35216), .Z(n27583) );
  AND U36218 ( .A(\modmult_1/xin[1023] ), .B(n35217), .Z(n35216) );
  IV U36219 ( .A(n35215), .Z(n35217) );
  XOR U36220 ( .A(n35218), .B(g_input[526]), .Z(n35215) );
  NAND U36221 ( .A(n35219), .B(mul_pow), .Z(n35218) );
  XOR U36222 ( .A(g_input[526]), .B(creg[526]), .Z(n35219) );
  XOR U36223 ( .A(n35220), .B(n35221), .Z(n35211) );
  ANDN U36224 ( .A(n35222), .B(n27590), .Z(n35221) );
  XOR U36225 ( .A(n35223), .B(\modmult_1/zin[0][524] ), .Z(n27590) );
  IV U36226 ( .A(n35220), .Z(n35223) );
  XNOR U36227 ( .A(n35220), .B(n27589), .Z(n35222) );
  XOR U36228 ( .A(n35224), .B(n35225), .Z(n27589) );
  AND U36229 ( .A(\modmult_1/xin[1023] ), .B(n35226), .Z(n35225) );
  IV U36230 ( .A(n35224), .Z(n35226) );
  XOR U36231 ( .A(n35227), .B(g_input[525]), .Z(n35224) );
  NAND U36232 ( .A(n35228), .B(mul_pow), .Z(n35227) );
  XOR U36233 ( .A(g_input[525]), .B(creg[525]), .Z(n35228) );
  XOR U36234 ( .A(n35229), .B(n35230), .Z(n35220) );
  ANDN U36235 ( .A(n35231), .B(n27596), .Z(n35230) );
  XOR U36236 ( .A(n35232), .B(\modmult_1/zin[0][523] ), .Z(n27596) );
  IV U36237 ( .A(n35229), .Z(n35232) );
  XNOR U36238 ( .A(n35229), .B(n27595), .Z(n35231) );
  XOR U36239 ( .A(n35233), .B(n35234), .Z(n27595) );
  AND U36240 ( .A(\modmult_1/xin[1023] ), .B(n35235), .Z(n35234) );
  IV U36241 ( .A(n35233), .Z(n35235) );
  XOR U36242 ( .A(n35236), .B(g_input[524]), .Z(n35233) );
  NAND U36243 ( .A(n35237), .B(mul_pow), .Z(n35236) );
  XOR U36244 ( .A(g_input[524]), .B(creg[524]), .Z(n35237) );
  XOR U36245 ( .A(n35238), .B(n35239), .Z(n35229) );
  ANDN U36246 ( .A(n35240), .B(n27602), .Z(n35239) );
  XOR U36247 ( .A(n35241), .B(\modmult_1/zin[0][522] ), .Z(n27602) );
  IV U36248 ( .A(n35238), .Z(n35241) );
  XNOR U36249 ( .A(n35238), .B(n27601), .Z(n35240) );
  XOR U36250 ( .A(n35242), .B(n35243), .Z(n27601) );
  AND U36251 ( .A(\modmult_1/xin[1023] ), .B(n35244), .Z(n35243) );
  IV U36252 ( .A(n35242), .Z(n35244) );
  XOR U36253 ( .A(n35245), .B(g_input[523]), .Z(n35242) );
  NAND U36254 ( .A(n35246), .B(mul_pow), .Z(n35245) );
  XOR U36255 ( .A(g_input[523]), .B(creg[523]), .Z(n35246) );
  XOR U36256 ( .A(n35247), .B(n35248), .Z(n35238) );
  ANDN U36257 ( .A(n35249), .B(n27608), .Z(n35248) );
  XOR U36258 ( .A(n35250), .B(\modmult_1/zin[0][521] ), .Z(n27608) );
  IV U36259 ( .A(n35247), .Z(n35250) );
  XNOR U36260 ( .A(n35247), .B(n27607), .Z(n35249) );
  XOR U36261 ( .A(n35251), .B(n35252), .Z(n27607) );
  AND U36262 ( .A(\modmult_1/xin[1023] ), .B(n35253), .Z(n35252) );
  IV U36263 ( .A(n35251), .Z(n35253) );
  XOR U36264 ( .A(n35254), .B(g_input[522]), .Z(n35251) );
  NAND U36265 ( .A(n35255), .B(mul_pow), .Z(n35254) );
  XOR U36266 ( .A(g_input[522]), .B(creg[522]), .Z(n35255) );
  XOR U36267 ( .A(n35256), .B(n35257), .Z(n35247) );
  ANDN U36268 ( .A(n35258), .B(n27614), .Z(n35257) );
  XOR U36269 ( .A(n35259), .B(\modmult_1/zin[0][520] ), .Z(n27614) );
  IV U36270 ( .A(n35256), .Z(n35259) );
  XNOR U36271 ( .A(n35256), .B(n27613), .Z(n35258) );
  XOR U36272 ( .A(n35260), .B(n35261), .Z(n27613) );
  AND U36273 ( .A(\modmult_1/xin[1023] ), .B(n35262), .Z(n35261) );
  IV U36274 ( .A(n35260), .Z(n35262) );
  XOR U36275 ( .A(n35263), .B(g_input[521]), .Z(n35260) );
  NAND U36276 ( .A(n35264), .B(mul_pow), .Z(n35263) );
  XOR U36277 ( .A(g_input[521]), .B(creg[521]), .Z(n35264) );
  XOR U36278 ( .A(n35265), .B(n35266), .Z(n35256) );
  ANDN U36279 ( .A(n35267), .B(n27620), .Z(n35266) );
  XOR U36280 ( .A(n35268), .B(\modmult_1/zin[0][519] ), .Z(n27620) );
  IV U36281 ( .A(n35265), .Z(n35268) );
  XNOR U36282 ( .A(n35265), .B(n27619), .Z(n35267) );
  XOR U36283 ( .A(n35269), .B(n35270), .Z(n27619) );
  AND U36284 ( .A(\modmult_1/xin[1023] ), .B(n35271), .Z(n35270) );
  IV U36285 ( .A(n35269), .Z(n35271) );
  XOR U36286 ( .A(n35272), .B(g_input[520]), .Z(n35269) );
  NAND U36287 ( .A(n35273), .B(mul_pow), .Z(n35272) );
  XOR U36288 ( .A(g_input[520]), .B(creg[520]), .Z(n35273) );
  XOR U36289 ( .A(n35274), .B(n35275), .Z(n35265) );
  ANDN U36290 ( .A(n35276), .B(n27626), .Z(n35275) );
  XOR U36291 ( .A(n35277), .B(\modmult_1/zin[0][518] ), .Z(n27626) );
  IV U36292 ( .A(n35274), .Z(n35277) );
  XNOR U36293 ( .A(n35274), .B(n27625), .Z(n35276) );
  XOR U36294 ( .A(n35278), .B(n35279), .Z(n27625) );
  AND U36295 ( .A(\modmult_1/xin[1023] ), .B(n35280), .Z(n35279) );
  IV U36296 ( .A(n35278), .Z(n35280) );
  XOR U36297 ( .A(n35281), .B(g_input[519]), .Z(n35278) );
  NAND U36298 ( .A(n35282), .B(mul_pow), .Z(n35281) );
  XOR U36299 ( .A(g_input[519]), .B(creg[519]), .Z(n35282) );
  XOR U36300 ( .A(n35283), .B(n35284), .Z(n35274) );
  ANDN U36301 ( .A(n35285), .B(n27632), .Z(n35284) );
  XOR U36302 ( .A(n35286), .B(\modmult_1/zin[0][517] ), .Z(n27632) );
  IV U36303 ( .A(n35283), .Z(n35286) );
  XNOR U36304 ( .A(n35283), .B(n27631), .Z(n35285) );
  XOR U36305 ( .A(n35287), .B(n35288), .Z(n27631) );
  AND U36306 ( .A(\modmult_1/xin[1023] ), .B(n35289), .Z(n35288) );
  IV U36307 ( .A(n35287), .Z(n35289) );
  XOR U36308 ( .A(n35290), .B(g_input[518]), .Z(n35287) );
  NAND U36309 ( .A(n35291), .B(mul_pow), .Z(n35290) );
  XOR U36310 ( .A(g_input[518]), .B(creg[518]), .Z(n35291) );
  XOR U36311 ( .A(n35292), .B(n35293), .Z(n35283) );
  ANDN U36312 ( .A(n35294), .B(n27638), .Z(n35293) );
  XOR U36313 ( .A(n35295), .B(\modmult_1/zin[0][516] ), .Z(n27638) );
  IV U36314 ( .A(n35292), .Z(n35295) );
  XNOR U36315 ( .A(n35292), .B(n27637), .Z(n35294) );
  XOR U36316 ( .A(n35296), .B(n35297), .Z(n27637) );
  AND U36317 ( .A(\modmult_1/xin[1023] ), .B(n35298), .Z(n35297) );
  IV U36318 ( .A(n35296), .Z(n35298) );
  XOR U36319 ( .A(n35299), .B(g_input[517]), .Z(n35296) );
  NAND U36320 ( .A(n35300), .B(mul_pow), .Z(n35299) );
  XOR U36321 ( .A(g_input[517]), .B(creg[517]), .Z(n35300) );
  XOR U36322 ( .A(n35301), .B(n35302), .Z(n35292) );
  ANDN U36323 ( .A(n35303), .B(n27644), .Z(n35302) );
  XOR U36324 ( .A(n35304), .B(\modmult_1/zin[0][515] ), .Z(n27644) );
  IV U36325 ( .A(n35301), .Z(n35304) );
  XNOR U36326 ( .A(n35301), .B(n27643), .Z(n35303) );
  XOR U36327 ( .A(n35305), .B(n35306), .Z(n27643) );
  AND U36328 ( .A(\modmult_1/xin[1023] ), .B(n35307), .Z(n35306) );
  IV U36329 ( .A(n35305), .Z(n35307) );
  XOR U36330 ( .A(n35308), .B(g_input[516]), .Z(n35305) );
  NAND U36331 ( .A(n35309), .B(mul_pow), .Z(n35308) );
  XOR U36332 ( .A(g_input[516]), .B(creg[516]), .Z(n35309) );
  XOR U36333 ( .A(n35310), .B(n35311), .Z(n35301) );
  ANDN U36334 ( .A(n35312), .B(n27650), .Z(n35311) );
  XOR U36335 ( .A(n35313), .B(\modmult_1/zin[0][514] ), .Z(n27650) );
  IV U36336 ( .A(n35310), .Z(n35313) );
  XNOR U36337 ( .A(n35310), .B(n27649), .Z(n35312) );
  XOR U36338 ( .A(n35314), .B(n35315), .Z(n27649) );
  AND U36339 ( .A(\modmult_1/xin[1023] ), .B(n35316), .Z(n35315) );
  IV U36340 ( .A(n35314), .Z(n35316) );
  XOR U36341 ( .A(n35317), .B(g_input[515]), .Z(n35314) );
  NAND U36342 ( .A(n35318), .B(mul_pow), .Z(n35317) );
  XOR U36343 ( .A(g_input[515]), .B(creg[515]), .Z(n35318) );
  XOR U36344 ( .A(n35319), .B(n35320), .Z(n35310) );
  ANDN U36345 ( .A(n35321), .B(n27656), .Z(n35320) );
  XOR U36346 ( .A(n35322), .B(\modmult_1/zin[0][513] ), .Z(n27656) );
  IV U36347 ( .A(n35319), .Z(n35322) );
  XNOR U36348 ( .A(n35319), .B(n27655), .Z(n35321) );
  XOR U36349 ( .A(n35323), .B(n35324), .Z(n27655) );
  AND U36350 ( .A(\modmult_1/xin[1023] ), .B(n35325), .Z(n35324) );
  IV U36351 ( .A(n35323), .Z(n35325) );
  XOR U36352 ( .A(n35326), .B(g_input[514]), .Z(n35323) );
  NAND U36353 ( .A(n35327), .B(mul_pow), .Z(n35326) );
  XOR U36354 ( .A(g_input[514]), .B(creg[514]), .Z(n35327) );
  XOR U36355 ( .A(n35328), .B(n35329), .Z(n35319) );
  ANDN U36356 ( .A(n35330), .B(n27662), .Z(n35329) );
  XOR U36357 ( .A(n35331), .B(\modmult_1/zin[0][512] ), .Z(n27662) );
  IV U36358 ( .A(n35328), .Z(n35331) );
  XNOR U36359 ( .A(n35328), .B(n27661), .Z(n35330) );
  XOR U36360 ( .A(n35332), .B(n35333), .Z(n27661) );
  AND U36361 ( .A(\modmult_1/xin[1023] ), .B(n35334), .Z(n35333) );
  IV U36362 ( .A(n35332), .Z(n35334) );
  XOR U36363 ( .A(n35335), .B(g_input[513]), .Z(n35332) );
  NAND U36364 ( .A(n35336), .B(mul_pow), .Z(n35335) );
  XOR U36365 ( .A(g_input[513]), .B(creg[513]), .Z(n35336) );
  XOR U36366 ( .A(n35337), .B(n35338), .Z(n35328) );
  ANDN U36367 ( .A(n35339), .B(n27668), .Z(n35338) );
  XOR U36368 ( .A(n35340), .B(\modmult_1/zin[0][511] ), .Z(n27668) );
  IV U36369 ( .A(n35337), .Z(n35340) );
  XNOR U36370 ( .A(n35337), .B(n27667), .Z(n35339) );
  XOR U36371 ( .A(n35341), .B(n35342), .Z(n27667) );
  AND U36372 ( .A(\modmult_1/xin[1023] ), .B(n35343), .Z(n35342) );
  IV U36373 ( .A(n35341), .Z(n35343) );
  XOR U36374 ( .A(n35344), .B(g_input[512]), .Z(n35341) );
  NAND U36375 ( .A(n35345), .B(mul_pow), .Z(n35344) );
  XOR U36376 ( .A(g_input[512]), .B(creg[512]), .Z(n35345) );
  XOR U36377 ( .A(n35346), .B(n35347), .Z(n35337) );
  ANDN U36378 ( .A(n35348), .B(n27674), .Z(n35347) );
  XOR U36379 ( .A(n35349), .B(\modmult_1/zin[0][510] ), .Z(n27674) );
  IV U36380 ( .A(n35346), .Z(n35349) );
  XNOR U36381 ( .A(n35346), .B(n27673), .Z(n35348) );
  XOR U36382 ( .A(n35350), .B(n35351), .Z(n27673) );
  AND U36383 ( .A(\modmult_1/xin[1023] ), .B(n35352), .Z(n35351) );
  IV U36384 ( .A(n35350), .Z(n35352) );
  XOR U36385 ( .A(n35353), .B(g_input[511]), .Z(n35350) );
  NAND U36386 ( .A(n35354), .B(mul_pow), .Z(n35353) );
  XOR U36387 ( .A(g_input[511]), .B(creg[511]), .Z(n35354) );
  XOR U36388 ( .A(n35355), .B(n35356), .Z(n35346) );
  ANDN U36389 ( .A(n35357), .B(n27680), .Z(n35356) );
  XOR U36390 ( .A(n35358), .B(\modmult_1/zin[0][509] ), .Z(n27680) );
  IV U36391 ( .A(n35355), .Z(n35358) );
  XNOR U36392 ( .A(n35355), .B(n27679), .Z(n35357) );
  XOR U36393 ( .A(n35359), .B(n35360), .Z(n27679) );
  AND U36394 ( .A(\modmult_1/xin[1023] ), .B(n35361), .Z(n35360) );
  IV U36395 ( .A(n35359), .Z(n35361) );
  XOR U36396 ( .A(n35362), .B(g_input[510]), .Z(n35359) );
  NAND U36397 ( .A(n35363), .B(mul_pow), .Z(n35362) );
  XOR U36398 ( .A(g_input[510]), .B(creg[510]), .Z(n35363) );
  XOR U36399 ( .A(n35364), .B(n35365), .Z(n35355) );
  ANDN U36400 ( .A(n35366), .B(n27686), .Z(n35365) );
  XOR U36401 ( .A(n35367), .B(\modmult_1/zin[0][508] ), .Z(n27686) );
  IV U36402 ( .A(n35364), .Z(n35367) );
  XNOR U36403 ( .A(n35364), .B(n27685), .Z(n35366) );
  XOR U36404 ( .A(n35368), .B(n35369), .Z(n27685) );
  AND U36405 ( .A(\modmult_1/xin[1023] ), .B(n35370), .Z(n35369) );
  IV U36406 ( .A(n35368), .Z(n35370) );
  XOR U36407 ( .A(n35371), .B(g_input[509]), .Z(n35368) );
  NAND U36408 ( .A(n35372), .B(mul_pow), .Z(n35371) );
  XOR U36409 ( .A(g_input[509]), .B(creg[509]), .Z(n35372) );
  XOR U36410 ( .A(n35373), .B(n35374), .Z(n35364) );
  ANDN U36411 ( .A(n35375), .B(n27692), .Z(n35374) );
  XOR U36412 ( .A(n35376), .B(\modmult_1/zin[0][507] ), .Z(n27692) );
  IV U36413 ( .A(n35373), .Z(n35376) );
  XNOR U36414 ( .A(n35373), .B(n27691), .Z(n35375) );
  XOR U36415 ( .A(n35377), .B(n35378), .Z(n27691) );
  AND U36416 ( .A(\modmult_1/xin[1023] ), .B(n35379), .Z(n35378) );
  IV U36417 ( .A(n35377), .Z(n35379) );
  XOR U36418 ( .A(n35380), .B(g_input[508]), .Z(n35377) );
  NAND U36419 ( .A(n35381), .B(mul_pow), .Z(n35380) );
  XOR U36420 ( .A(g_input[508]), .B(creg[508]), .Z(n35381) );
  XOR U36421 ( .A(n35382), .B(n35383), .Z(n35373) );
  ANDN U36422 ( .A(n35384), .B(n27698), .Z(n35383) );
  XOR U36423 ( .A(n35385), .B(\modmult_1/zin[0][506] ), .Z(n27698) );
  IV U36424 ( .A(n35382), .Z(n35385) );
  XNOR U36425 ( .A(n35382), .B(n27697), .Z(n35384) );
  XOR U36426 ( .A(n35386), .B(n35387), .Z(n27697) );
  AND U36427 ( .A(\modmult_1/xin[1023] ), .B(n35388), .Z(n35387) );
  IV U36428 ( .A(n35386), .Z(n35388) );
  XOR U36429 ( .A(n35389), .B(g_input[507]), .Z(n35386) );
  NAND U36430 ( .A(n35390), .B(mul_pow), .Z(n35389) );
  XOR U36431 ( .A(g_input[507]), .B(creg[507]), .Z(n35390) );
  XOR U36432 ( .A(n35391), .B(n35392), .Z(n35382) );
  ANDN U36433 ( .A(n35393), .B(n27704), .Z(n35392) );
  XOR U36434 ( .A(n35394), .B(\modmult_1/zin[0][505] ), .Z(n27704) );
  IV U36435 ( .A(n35391), .Z(n35394) );
  XNOR U36436 ( .A(n35391), .B(n27703), .Z(n35393) );
  XOR U36437 ( .A(n35395), .B(n35396), .Z(n27703) );
  AND U36438 ( .A(\modmult_1/xin[1023] ), .B(n35397), .Z(n35396) );
  IV U36439 ( .A(n35395), .Z(n35397) );
  XOR U36440 ( .A(n35398), .B(g_input[506]), .Z(n35395) );
  NAND U36441 ( .A(n35399), .B(mul_pow), .Z(n35398) );
  XOR U36442 ( .A(g_input[506]), .B(creg[506]), .Z(n35399) );
  XOR U36443 ( .A(n35400), .B(n35401), .Z(n35391) );
  ANDN U36444 ( .A(n35402), .B(n27710), .Z(n35401) );
  XOR U36445 ( .A(n35403), .B(\modmult_1/zin[0][504] ), .Z(n27710) );
  IV U36446 ( .A(n35400), .Z(n35403) );
  XNOR U36447 ( .A(n35400), .B(n27709), .Z(n35402) );
  XOR U36448 ( .A(n35404), .B(n35405), .Z(n27709) );
  AND U36449 ( .A(\modmult_1/xin[1023] ), .B(n35406), .Z(n35405) );
  IV U36450 ( .A(n35404), .Z(n35406) );
  XOR U36451 ( .A(n35407), .B(g_input[505]), .Z(n35404) );
  NAND U36452 ( .A(n35408), .B(mul_pow), .Z(n35407) );
  XOR U36453 ( .A(g_input[505]), .B(creg[505]), .Z(n35408) );
  XOR U36454 ( .A(n35409), .B(n35410), .Z(n35400) );
  ANDN U36455 ( .A(n35411), .B(n27716), .Z(n35410) );
  XOR U36456 ( .A(n35412), .B(\modmult_1/zin[0][503] ), .Z(n27716) );
  IV U36457 ( .A(n35409), .Z(n35412) );
  XNOR U36458 ( .A(n35409), .B(n27715), .Z(n35411) );
  XOR U36459 ( .A(n35413), .B(n35414), .Z(n27715) );
  AND U36460 ( .A(\modmult_1/xin[1023] ), .B(n35415), .Z(n35414) );
  IV U36461 ( .A(n35413), .Z(n35415) );
  XOR U36462 ( .A(n35416), .B(g_input[504]), .Z(n35413) );
  NAND U36463 ( .A(n35417), .B(mul_pow), .Z(n35416) );
  XOR U36464 ( .A(g_input[504]), .B(creg[504]), .Z(n35417) );
  XOR U36465 ( .A(n35418), .B(n35419), .Z(n35409) );
  ANDN U36466 ( .A(n35420), .B(n27722), .Z(n35419) );
  XOR U36467 ( .A(n35421), .B(\modmult_1/zin[0][502] ), .Z(n27722) );
  IV U36468 ( .A(n35418), .Z(n35421) );
  XNOR U36469 ( .A(n35418), .B(n27721), .Z(n35420) );
  XOR U36470 ( .A(n35422), .B(n35423), .Z(n27721) );
  AND U36471 ( .A(\modmult_1/xin[1023] ), .B(n35424), .Z(n35423) );
  IV U36472 ( .A(n35422), .Z(n35424) );
  XOR U36473 ( .A(n35425), .B(g_input[503]), .Z(n35422) );
  NAND U36474 ( .A(n35426), .B(mul_pow), .Z(n35425) );
  XOR U36475 ( .A(g_input[503]), .B(creg[503]), .Z(n35426) );
  XOR U36476 ( .A(n35427), .B(n35428), .Z(n35418) );
  ANDN U36477 ( .A(n35429), .B(n27728), .Z(n35428) );
  XOR U36478 ( .A(n35430), .B(\modmult_1/zin[0][501] ), .Z(n27728) );
  IV U36479 ( .A(n35427), .Z(n35430) );
  XNOR U36480 ( .A(n35427), .B(n27727), .Z(n35429) );
  XOR U36481 ( .A(n35431), .B(n35432), .Z(n27727) );
  AND U36482 ( .A(\modmult_1/xin[1023] ), .B(n35433), .Z(n35432) );
  IV U36483 ( .A(n35431), .Z(n35433) );
  XOR U36484 ( .A(n35434), .B(g_input[502]), .Z(n35431) );
  NAND U36485 ( .A(n35435), .B(mul_pow), .Z(n35434) );
  XOR U36486 ( .A(g_input[502]), .B(creg[502]), .Z(n35435) );
  XOR U36487 ( .A(n35436), .B(n35437), .Z(n35427) );
  ANDN U36488 ( .A(n35438), .B(n27734), .Z(n35437) );
  XOR U36489 ( .A(n35439), .B(\modmult_1/zin[0][500] ), .Z(n27734) );
  IV U36490 ( .A(n35436), .Z(n35439) );
  XNOR U36491 ( .A(n35436), .B(n27733), .Z(n35438) );
  XOR U36492 ( .A(n35440), .B(n35441), .Z(n27733) );
  AND U36493 ( .A(\modmult_1/xin[1023] ), .B(n35442), .Z(n35441) );
  IV U36494 ( .A(n35440), .Z(n35442) );
  XOR U36495 ( .A(n35443), .B(g_input[501]), .Z(n35440) );
  NAND U36496 ( .A(n35444), .B(mul_pow), .Z(n35443) );
  XOR U36497 ( .A(g_input[501]), .B(creg[501]), .Z(n35444) );
  XOR U36498 ( .A(n35445), .B(n35446), .Z(n35436) );
  ANDN U36499 ( .A(n35447), .B(n27740), .Z(n35446) );
  XOR U36500 ( .A(n35448), .B(\modmult_1/zin[0][499] ), .Z(n27740) );
  IV U36501 ( .A(n35445), .Z(n35448) );
  XNOR U36502 ( .A(n35445), .B(n27739), .Z(n35447) );
  XOR U36503 ( .A(n35449), .B(n35450), .Z(n27739) );
  AND U36504 ( .A(\modmult_1/xin[1023] ), .B(n35451), .Z(n35450) );
  IV U36505 ( .A(n35449), .Z(n35451) );
  XOR U36506 ( .A(n35452), .B(g_input[500]), .Z(n35449) );
  NAND U36507 ( .A(n35453), .B(mul_pow), .Z(n35452) );
  XOR U36508 ( .A(g_input[500]), .B(creg[500]), .Z(n35453) );
  XOR U36509 ( .A(n35454), .B(n35455), .Z(n35445) );
  ANDN U36510 ( .A(n35456), .B(n27746), .Z(n35455) );
  XOR U36511 ( .A(n35457), .B(\modmult_1/zin[0][498] ), .Z(n27746) );
  IV U36512 ( .A(n35454), .Z(n35457) );
  XNOR U36513 ( .A(n35454), .B(n27745), .Z(n35456) );
  XOR U36514 ( .A(n35458), .B(n35459), .Z(n27745) );
  AND U36515 ( .A(\modmult_1/xin[1023] ), .B(n35460), .Z(n35459) );
  IV U36516 ( .A(n35458), .Z(n35460) );
  XOR U36517 ( .A(n35461), .B(g_input[499]), .Z(n35458) );
  NAND U36518 ( .A(n35462), .B(mul_pow), .Z(n35461) );
  XOR U36519 ( .A(g_input[499]), .B(creg[499]), .Z(n35462) );
  XOR U36520 ( .A(n35463), .B(n35464), .Z(n35454) );
  ANDN U36521 ( .A(n35465), .B(n27752), .Z(n35464) );
  XOR U36522 ( .A(n35466), .B(\modmult_1/zin[0][497] ), .Z(n27752) );
  IV U36523 ( .A(n35463), .Z(n35466) );
  XNOR U36524 ( .A(n35463), .B(n27751), .Z(n35465) );
  XOR U36525 ( .A(n35467), .B(n35468), .Z(n27751) );
  AND U36526 ( .A(\modmult_1/xin[1023] ), .B(n35469), .Z(n35468) );
  IV U36527 ( .A(n35467), .Z(n35469) );
  XOR U36528 ( .A(n35470), .B(g_input[498]), .Z(n35467) );
  NAND U36529 ( .A(n35471), .B(mul_pow), .Z(n35470) );
  XOR U36530 ( .A(g_input[498]), .B(creg[498]), .Z(n35471) );
  XOR U36531 ( .A(n35472), .B(n35473), .Z(n35463) );
  ANDN U36532 ( .A(n35474), .B(n27758), .Z(n35473) );
  XOR U36533 ( .A(n35475), .B(\modmult_1/zin[0][496] ), .Z(n27758) );
  IV U36534 ( .A(n35472), .Z(n35475) );
  XNOR U36535 ( .A(n35472), .B(n27757), .Z(n35474) );
  XOR U36536 ( .A(n35476), .B(n35477), .Z(n27757) );
  AND U36537 ( .A(\modmult_1/xin[1023] ), .B(n35478), .Z(n35477) );
  IV U36538 ( .A(n35476), .Z(n35478) );
  XOR U36539 ( .A(n35479), .B(g_input[497]), .Z(n35476) );
  NAND U36540 ( .A(n35480), .B(mul_pow), .Z(n35479) );
  XOR U36541 ( .A(g_input[497]), .B(creg[497]), .Z(n35480) );
  XOR U36542 ( .A(n35481), .B(n35482), .Z(n35472) );
  ANDN U36543 ( .A(n35483), .B(n27764), .Z(n35482) );
  XOR U36544 ( .A(n35484), .B(\modmult_1/zin[0][495] ), .Z(n27764) );
  IV U36545 ( .A(n35481), .Z(n35484) );
  XNOR U36546 ( .A(n35481), .B(n27763), .Z(n35483) );
  XOR U36547 ( .A(n35485), .B(n35486), .Z(n27763) );
  AND U36548 ( .A(\modmult_1/xin[1023] ), .B(n35487), .Z(n35486) );
  IV U36549 ( .A(n35485), .Z(n35487) );
  XOR U36550 ( .A(n35488), .B(g_input[496]), .Z(n35485) );
  NAND U36551 ( .A(n35489), .B(mul_pow), .Z(n35488) );
  XOR U36552 ( .A(g_input[496]), .B(creg[496]), .Z(n35489) );
  XOR U36553 ( .A(n35490), .B(n35491), .Z(n35481) );
  ANDN U36554 ( .A(n35492), .B(n27770), .Z(n35491) );
  XOR U36555 ( .A(n35493), .B(\modmult_1/zin[0][494] ), .Z(n27770) );
  IV U36556 ( .A(n35490), .Z(n35493) );
  XNOR U36557 ( .A(n35490), .B(n27769), .Z(n35492) );
  XOR U36558 ( .A(n35494), .B(n35495), .Z(n27769) );
  AND U36559 ( .A(\modmult_1/xin[1023] ), .B(n35496), .Z(n35495) );
  IV U36560 ( .A(n35494), .Z(n35496) );
  XOR U36561 ( .A(n35497), .B(g_input[495]), .Z(n35494) );
  NAND U36562 ( .A(n35498), .B(mul_pow), .Z(n35497) );
  XOR U36563 ( .A(g_input[495]), .B(creg[495]), .Z(n35498) );
  XOR U36564 ( .A(n35499), .B(n35500), .Z(n35490) );
  ANDN U36565 ( .A(n35501), .B(n27776), .Z(n35500) );
  XOR U36566 ( .A(n35502), .B(\modmult_1/zin[0][493] ), .Z(n27776) );
  IV U36567 ( .A(n35499), .Z(n35502) );
  XNOR U36568 ( .A(n35499), .B(n27775), .Z(n35501) );
  XOR U36569 ( .A(n35503), .B(n35504), .Z(n27775) );
  AND U36570 ( .A(\modmult_1/xin[1023] ), .B(n35505), .Z(n35504) );
  IV U36571 ( .A(n35503), .Z(n35505) );
  XOR U36572 ( .A(n35506), .B(g_input[494]), .Z(n35503) );
  NAND U36573 ( .A(n35507), .B(mul_pow), .Z(n35506) );
  XOR U36574 ( .A(g_input[494]), .B(creg[494]), .Z(n35507) );
  XOR U36575 ( .A(n35508), .B(n35509), .Z(n35499) );
  ANDN U36576 ( .A(n35510), .B(n27782), .Z(n35509) );
  XOR U36577 ( .A(n35511), .B(\modmult_1/zin[0][492] ), .Z(n27782) );
  IV U36578 ( .A(n35508), .Z(n35511) );
  XNOR U36579 ( .A(n35508), .B(n27781), .Z(n35510) );
  XOR U36580 ( .A(n35512), .B(n35513), .Z(n27781) );
  AND U36581 ( .A(\modmult_1/xin[1023] ), .B(n35514), .Z(n35513) );
  IV U36582 ( .A(n35512), .Z(n35514) );
  XOR U36583 ( .A(n35515), .B(g_input[493]), .Z(n35512) );
  NAND U36584 ( .A(n35516), .B(mul_pow), .Z(n35515) );
  XOR U36585 ( .A(g_input[493]), .B(creg[493]), .Z(n35516) );
  XOR U36586 ( .A(n35517), .B(n35518), .Z(n35508) );
  ANDN U36587 ( .A(n35519), .B(n27788), .Z(n35518) );
  XOR U36588 ( .A(n35520), .B(\modmult_1/zin[0][491] ), .Z(n27788) );
  IV U36589 ( .A(n35517), .Z(n35520) );
  XNOR U36590 ( .A(n35517), .B(n27787), .Z(n35519) );
  XOR U36591 ( .A(n35521), .B(n35522), .Z(n27787) );
  AND U36592 ( .A(\modmult_1/xin[1023] ), .B(n35523), .Z(n35522) );
  IV U36593 ( .A(n35521), .Z(n35523) );
  XOR U36594 ( .A(n35524), .B(g_input[492]), .Z(n35521) );
  NAND U36595 ( .A(n35525), .B(mul_pow), .Z(n35524) );
  XOR U36596 ( .A(g_input[492]), .B(creg[492]), .Z(n35525) );
  XOR U36597 ( .A(n35526), .B(n35527), .Z(n35517) );
  ANDN U36598 ( .A(n35528), .B(n27794), .Z(n35527) );
  XOR U36599 ( .A(n35529), .B(\modmult_1/zin[0][490] ), .Z(n27794) );
  IV U36600 ( .A(n35526), .Z(n35529) );
  XNOR U36601 ( .A(n35526), .B(n27793), .Z(n35528) );
  XOR U36602 ( .A(n35530), .B(n35531), .Z(n27793) );
  AND U36603 ( .A(\modmult_1/xin[1023] ), .B(n35532), .Z(n35531) );
  IV U36604 ( .A(n35530), .Z(n35532) );
  XOR U36605 ( .A(n35533), .B(g_input[491]), .Z(n35530) );
  NAND U36606 ( .A(n35534), .B(mul_pow), .Z(n35533) );
  XOR U36607 ( .A(g_input[491]), .B(creg[491]), .Z(n35534) );
  XOR U36608 ( .A(n35535), .B(n35536), .Z(n35526) );
  ANDN U36609 ( .A(n35537), .B(n27800), .Z(n35536) );
  XOR U36610 ( .A(n35538), .B(\modmult_1/zin[0][489] ), .Z(n27800) );
  IV U36611 ( .A(n35535), .Z(n35538) );
  XNOR U36612 ( .A(n35535), .B(n27799), .Z(n35537) );
  XOR U36613 ( .A(n35539), .B(n35540), .Z(n27799) );
  AND U36614 ( .A(\modmult_1/xin[1023] ), .B(n35541), .Z(n35540) );
  IV U36615 ( .A(n35539), .Z(n35541) );
  XOR U36616 ( .A(n35542), .B(g_input[490]), .Z(n35539) );
  NAND U36617 ( .A(n35543), .B(mul_pow), .Z(n35542) );
  XOR U36618 ( .A(g_input[490]), .B(creg[490]), .Z(n35543) );
  XOR U36619 ( .A(n35544), .B(n35545), .Z(n35535) );
  ANDN U36620 ( .A(n35546), .B(n27806), .Z(n35545) );
  XOR U36621 ( .A(n35547), .B(\modmult_1/zin[0][488] ), .Z(n27806) );
  IV U36622 ( .A(n35544), .Z(n35547) );
  XNOR U36623 ( .A(n35544), .B(n27805), .Z(n35546) );
  XOR U36624 ( .A(n35548), .B(n35549), .Z(n27805) );
  AND U36625 ( .A(\modmult_1/xin[1023] ), .B(n35550), .Z(n35549) );
  IV U36626 ( .A(n35548), .Z(n35550) );
  XOR U36627 ( .A(n35551), .B(g_input[489]), .Z(n35548) );
  NAND U36628 ( .A(n35552), .B(mul_pow), .Z(n35551) );
  XOR U36629 ( .A(g_input[489]), .B(creg[489]), .Z(n35552) );
  XOR U36630 ( .A(n35553), .B(n35554), .Z(n35544) );
  ANDN U36631 ( .A(n35555), .B(n27812), .Z(n35554) );
  XOR U36632 ( .A(n35556), .B(\modmult_1/zin[0][487] ), .Z(n27812) );
  IV U36633 ( .A(n35553), .Z(n35556) );
  XNOR U36634 ( .A(n35553), .B(n27811), .Z(n35555) );
  XOR U36635 ( .A(n35557), .B(n35558), .Z(n27811) );
  AND U36636 ( .A(\modmult_1/xin[1023] ), .B(n35559), .Z(n35558) );
  IV U36637 ( .A(n35557), .Z(n35559) );
  XOR U36638 ( .A(n35560), .B(g_input[488]), .Z(n35557) );
  NAND U36639 ( .A(n35561), .B(mul_pow), .Z(n35560) );
  XOR U36640 ( .A(g_input[488]), .B(creg[488]), .Z(n35561) );
  XOR U36641 ( .A(n35562), .B(n35563), .Z(n35553) );
  ANDN U36642 ( .A(n35564), .B(n27818), .Z(n35563) );
  XOR U36643 ( .A(n35565), .B(\modmult_1/zin[0][486] ), .Z(n27818) );
  IV U36644 ( .A(n35562), .Z(n35565) );
  XNOR U36645 ( .A(n35562), .B(n27817), .Z(n35564) );
  XOR U36646 ( .A(n35566), .B(n35567), .Z(n27817) );
  AND U36647 ( .A(\modmult_1/xin[1023] ), .B(n35568), .Z(n35567) );
  IV U36648 ( .A(n35566), .Z(n35568) );
  XOR U36649 ( .A(n35569), .B(g_input[487]), .Z(n35566) );
  NAND U36650 ( .A(n35570), .B(mul_pow), .Z(n35569) );
  XOR U36651 ( .A(g_input[487]), .B(creg[487]), .Z(n35570) );
  XOR U36652 ( .A(n35571), .B(n35572), .Z(n35562) );
  ANDN U36653 ( .A(n35573), .B(n27824), .Z(n35572) );
  XOR U36654 ( .A(n35574), .B(\modmult_1/zin[0][485] ), .Z(n27824) );
  IV U36655 ( .A(n35571), .Z(n35574) );
  XNOR U36656 ( .A(n35571), .B(n27823), .Z(n35573) );
  XOR U36657 ( .A(n35575), .B(n35576), .Z(n27823) );
  AND U36658 ( .A(\modmult_1/xin[1023] ), .B(n35577), .Z(n35576) );
  IV U36659 ( .A(n35575), .Z(n35577) );
  XOR U36660 ( .A(n35578), .B(g_input[486]), .Z(n35575) );
  NAND U36661 ( .A(n35579), .B(mul_pow), .Z(n35578) );
  XOR U36662 ( .A(g_input[486]), .B(creg[486]), .Z(n35579) );
  XOR U36663 ( .A(n35580), .B(n35581), .Z(n35571) );
  ANDN U36664 ( .A(n35582), .B(n27830), .Z(n35581) );
  XOR U36665 ( .A(n35583), .B(\modmult_1/zin[0][484] ), .Z(n27830) );
  IV U36666 ( .A(n35580), .Z(n35583) );
  XNOR U36667 ( .A(n35580), .B(n27829), .Z(n35582) );
  XOR U36668 ( .A(n35584), .B(n35585), .Z(n27829) );
  AND U36669 ( .A(\modmult_1/xin[1023] ), .B(n35586), .Z(n35585) );
  IV U36670 ( .A(n35584), .Z(n35586) );
  XOR U36671 ( .A(n35587), .B(g_input[485]), .Z(n35584) );
  NAND U36672 ( .A(n35588), .B(mul_pow), .Z(n35587) );
  XOR U36673 ( .A(g_input[485]), .B(creg[485]), .Z(n35588) );
  XOR U36674 ( .A(n35589), .B(n35590), .Z(n35580) );
  ANDN U36675 ( .A(n35591), .B(n27836), .Z(n35590) );
  XOR U36676 ( .A(n35592), .B(\modmult_1/zin[0][483] ), .Z(n27836) );
  IV U36677 ( .A(n35589), .Z(n35592) );
  XNOR U36678 ( .A(n35589), .B(n27835), .Z(n35591) );
  XOR U36679 ( .A(n35593), .B(n35594), .Z(n27835) );
  AND U36680 ( .A(\modmult_1/xin[1023] ), .B(n35595), .Z(n35594) );
  IV U36681 ( .A(n35593), .Z(n35595) );
  XOR U36682 ( .A(n35596), .B(g_input[484]), .Z(n35593) );
  NAND U36683 ( .A(n35597), .B(mul_pow), .Z(n35596) );
  XOR U36684 ( .A(g_input[484]), .B(creg[484]), .Z(n35597) );
  XOR U36685 ( .A(n35598), .B(n35599), .Z(n35589) );
  ANDN U36686 ( .A(n35600), .B(n27842), .Z(n35599) );
  XOR U36687 ( .A(n35601), .B(\modmult_1/zin[0][482] ), .Z(n27842) );
  IV U36688 ( .A(n35598), .Z(n35601) );
  XNOR U36689 ( .A(n35598), .B(n27841), .Z(n35600) );
  XOR U36690 ( .A(n35602), .B(n35603), .Z(n27841) );
  AND U36691 ( .A(\modmult_1/xin[1023] ), .B(n35604), .Z(n35603) );
  IV U36692 ( .A(n35602), .Z(n35604) );
  XOR U36693 ( .A(n35605), .B(g_input[483]), .Z(n35602) );
  NAND U36694 ( .A(n35606), .B(mul_pow), .Z(n35605) );
  XOR U36695 ( .A(g_input[483]), .B(creg[483]), .Z(n35606) );
  XOR U36696 ( .A(n35607), .B(n35608), .Z(n35598) );
  ANDN U36697 ( .A(n35609), .B(n27848), .Z(n35608) );
  XOR U36698 ( .A(n35610), .B(\modmult_1/zin[0][481] ), .Z(n27848) );
  IV U36699 ( .A(n35607), .Z(n35610) );
  XNOR U36700 ( .A(n35607), .B(n27847), .Z(n35609) );
  XOR U36701 ( .A(n35611), .B(n35612), .Z(n27847) );
  AND U36702 ( .A(\modmult_1/xin[1023] ), .B(n35613), .Z(n35612) );
  IV U36703 ( .A(n35611), .Z(n35613) );
  XOR U36704 ( .A(n35614), .B(g_input[482]), .Z(n35611) );
  NAND U36705 ( .A(n35615), .B(mul_pow), .Z(n35614) );
  XOR U36706 ( .A(g_input[482]), .B(creg[482]), .Z(n35615) );
  XOR U36707 ( .A(n35616), .B(n35617), .Z(n35607) );
  ANDN U36708 ( .A(n35618), .B(n27854), .Z(n35617) );
  XOR U36709 ( .A(n35619), .B(\modmult_1/zin[0][480] ), .Z(n27854) );
  IV U36710 ( .A(n35616), .Z(n35619) );
  XNOR U36711 ( .A(n35616), .B(n27853), .Z(n35618) );
  XOR U36712 ( .A(n35620), .B(n35621), .Z(n27853) );
  AND U36713 ( .A(\modmult_1/xin[1023] ), .B(n35622), .Z(n35621) );
  IV U36714 ( .A(n35620), .Z(n35622) );
  XOR U36715 ( .A(n35623), .B(g_input[481]), .Z(n35620) );
  NAND U36716 ( .A(n35624), .B(mul_pow), .Z(n35623) );
  XOR U36717 ( .A(g_input[481]), .B(creg[481]), .Z(n35624) );
  XOR U36718 ( .A(n35625), .B(n35626), .Z(n35616) );
  ANDN U36719 ( .A(n35627), .B(n27860), .Z(n35626) );
  XOR U36720 ( .A(n35628), .B(\modmult_1/zin[0][479] ), .Z(n27860) );
  IV U36721 ( .A(n35625), .Z(n35628) );
  XNOR U36722 ( .A(n35625), .B(n27859), .Z(n35627) );
  XOR U36723 ( .A(n35629), .B(n35630), .Z(n27859) );
  AND U36724 ( .A(\modmult_1/xin[1023] ), .B(n35631), .Z(n35630) );
  IV U36725 ( .A(n35629), .Z(n35631) );
  XOR U36726 ( .A(n35632), .B(g_input[480]), .Z(n35629) );
  NAND U36727 ( .A(n35633), .B(mul_pow), .Z(n35632) );
  XOR U36728 ( .A(g_input[480]), .B(creg[480]), .Z(n35633) );
  XOR U36729 ( .A(n35634), .B(n35635), .Z(n35625) );
  ANDN U36730 ( .A(n35636), .B(n27866), .Z(n35635) );
  XOR U36731 ( .A(n35637), .B(\modmult_1/zin[0][478] ), .Z(n27866) );
  IV U36732 ( .A(n35634), .Z(n35637) );
  XNOR U36733 ( .A(n35634), .B(n27865), .Z(n35636) );
  XOR U36734 ( .A(n35638), .B(n35639), .Z(n27865) );
  AND U36735 ( .A(\modmult_1/xin[1023] ), .B(n35640), .Z(n35639) );
  IV U36736 ( .A(n35638), .Z(n35640) );
  XOR U36737 ( .A(n35641), .B(g_input[479]), .Z(n35638) );
  NAND U36738 ( .A(n35642), .B(mul_pow), .Z(n35641) );
  XOR U36739 ( .A(g_input[479]), .B(creg[479]), .Z(n35642) );
  XOR U36740 ( .A(n35643), .B(n35644), .Z(n35634) );
  ANDN U36741 ( .A(n35645), .B(n27872), .Z(n35644) );
  XOR U36742 ( .A(n35646), .B(\modmult_1/zin[0][477] ), .Z(n27872) );
  IV U36743 ( .A(n35643), .Z(n35646) );
  XNOR U36744 ( .A(n35643), .B(n27871), .Z(n35645) );
  XOR U36745 ( .A(n35647), .B(n35648), .Z(n27871) );
  AND U36746 ( .A(\modmult_1/xin[1023] ), .B(n35649), .Z(n35648) );
  IV U36747 ( .A(n35647), .Z(n35649) );
  XOR U36748 ( .A(n35650), .B(g_input[478]), .Z(n35647) );
  NAND U36749 ( .A(n35651), .B(mul_pow), .Z(n35650) );
  XOR U36750 ( .A(g_input[478]), .B(creg[478]), .Z(n35651) );
  XOR U36751 ( .A(n35652), .B(n35653), .Z(n35643) );
  ANDN U36752 ( .A(n35654), .B(n27878), .Z(n35653) );
  XOR U36753 ( .A(n35655), .B(\modmult_1/zin[0][476] ), .Z(n27878) );
  IV U36754 ( .A(n35652), .Z(n35655) );
  XNOR U36755 ( .A(n35652), .B(n27877), .Z(n35654) );
  XOR U36756 ( .A(n35656), .B(n35657), .Z(n27877) );
  AND U36757 ( .A(\modmult_1/xin[1023] ), .B(n35658), .Z(n35657) );
  IV U36758 ( .A(n35656), .Z(n35658) );
  XOR U36759 ( .A(n35659), .B(g_input[477]), .Z(n35656) );
  NAND U36760 ( .A(n35660), .B(mul_pow), .Z(n35659) );
  XOR U36761 ( .A(g_input[477]), .B(creg[477]), .Z(n35660) );
  XOR U36762 ( .A(n35661), .B(n35662), .Z(n35652) );
  ANDN U36763 ( .A(n35663), .B(n27884), .Z(n35662) );
  XOR U36764 ( .A(n35664), .B(\modmult_1/zin[0][475] ), .Z(n27884) );
  IV U36765 ( .A(n35661), .Z(n35664) );
  XNOR U36766 ( .A(n35661), .B(n27883), .Z(n35663) );
  XOR U36767 ( .A(n35665), .B(n35666), .Z(n27883) );
  AND U36768 ( .A(\modmult_1/xin[1023] ), .B(n35667), .Z(n35666) );
  IV U36769 ( .A(n35665), .Z(n35667) );
  XOR U36770 ( .A(n35668), .B(g_input[476]), .Z(n35665) );
  NAND U36771 ( .A(n35669), .B(mul_pow), .Z(n35668) );
  XOR U36772 ( .A(g_input[476]), .B(creg[476]), .Z(n35669) );
  XOR U36773 ( .A(n35670), .B(n35671), .Z(n35661) );
  ANDN U36774 ( .A(n35672), .B(n27890), .Z(n35671) );
  XOR U36775 ( .A(n35673), .B(\modmult_1/zin[0][474] ), .Z(n27890) );
  IV U36776 ( .A(n35670), .Z(n35673) );
  XNOR U36777 ( .A(n35670), .B(n27889), .Z(n35672) );
  XOR U36778 ( .A(n35674), .B(n35675), .Z(n27889) );
  AND U36779 ( .A(\modmult_1/xin[1023] ), .B(n35676), .Z(n35675) );
  IV U36780 ( .A(n35674), .Z(n35676) );
  XOR U36781 ( .A(n35677), .B(g_input[475]), .Z(n35674) );
  NAND U36782 ( .A(n35678), .B(mul_pow), .Z(n35677) );
  XOR U36783 ( .A(g_input[475]), .B(creg[475]), .Z(n35678) );
  XOR U36784 ( .A(n35679), .B(n35680), .Z(n35670) );
  ANDN U36785 ( .A(n35681), .B(n27896), .Z(n35680) );
  XOR U36786 ( .A(n35682), .B(\modmult_1/zin[0][473] ), .Z(n27896) );
  IV U36787 ( .A(n35679), .Z(n35682) );
  XNOR U36788 ( .A(n35679), .B(n27895), .Z(n35681) );
  XOR U36789 ( .A(n35683), .B(n35684), .Z(n27895) );
  AND U36790 ( .A(\modmult_1/xin[1023] ), .B(n35685), .Z(n35684) );
  IV U36791 ( .A(n35683), .Z(n35685) );
  XOR U36792 ( .A(n35686), .B(g_input[474]), .Z(n35683) );
  NAND U36793 ( .A(n35687), .B(mul_pow), .Z(n35686) );
  XOR U36794 ( .A(g_input[474]), .B(creg[474]), .Z(n35687) );
  XOR U36795 ( .A(n35688), .B(n35689), .Z(n35679) );
  ANDN U36796 ( .A(n35690), .B(n27902), .Z(n35689) );
  XOR U36797 ( .A(n35691), .B(\modmult_1/zin[0][472] ), .Z(n27902) );
  IV U36798 ( .A(n35688), .Z(n35691) );
  XNOR U36799 ( .A(n35688), .B(n27901), .Z(n35690) );
  XOR U36800 ( .A(n35692), .B(n35693), .Z(n27901) );
  AND U36801 ( .A(\modmult_1/xin[1023] ), .B(n35694), .Z(n35693) );
  IV U36802 ( .A(n35692), .Z(n35694) );
  XOR U36803 ( .A(n35695), .B(g_input[473]), .Z(n35692) );
  NAND U36804 ( .A(n35696), .B(mul_pow), .Z(n35695) );
  XOR U36805 ( .A(g_input[473]), .B(creg[473]), .Z(n35696) );
  XOR U36806 ( .A(n35697), .B(n35698), .Z(n35688) );
  ANDN U36807 ( .A(n35699), .B(n27908), .Z(n35698) );
  XOR U36808 ( .A(n35700), .B(\modmult_1/zin[0][471] ), .Z(n27908) );
  IV U36809 ( .A(n35697), .Z(n35700) );
  XNOR U36810 ( .A(n35697), .B(n27907), .Z(n35699) );
  XOR U36811 ( .A(n35701), .B(n35702), .Z(n27907) );
  AND U36812 ( .A(\modmult_1/xin[1023] ), .B(n35703), .Z(n35702) );
  IV U36813 ( .A(n35701), .Z(n35703) );
  XOR U36814 ( .A(n35704), .B(g_input[472]), .Z(n35701) );
  NAND U36815 ( .A(n35705), .B(mul_pow), .Z(n35704) );
  XOR U36816 ( .A(g_input[472]), .B(creg[472]), .Z(n35705) );
  XOR U36817 ( .A(n35706), .B(n35707), .Z(n35697) );
  ANDN U36818 ( .A(n35708), .B(n27914), .Z(n35707) );
  XOR U36819 ( .A(n35709), .B(\modmult_1/zin[0][470] ), .Z(n27914) );
  IV U36820 ( .A(n35706), .Z(n35709) );
  XNOR U36821 ( .A(n35706), .B(n27913), .Z(n35708) );
  XOR U36822 ( .A(n35710), .B(n35711), .Z(n27913) );
  AND U36823 ( .A(\modmult_1/xin[1023] ), .B(n35712), .Z(n35711) );
  IV U36824 ( .A(n35710), .Z(n35712) );
  XOR U36825 ( .A(n35713), .B(g_input[471]), .Z(n35710) );
  NAND U36826 ( .A(n35714), .B(mul_pow), .Z(n35713) );
  XOR U36827 ( .A(g_input[471]), .B(creg[471]), .Z(n35714) );
  XOR U36828 ( .A(n35715), .B(n35716), .Z(n35706) );
  ANDN U36829 ( .A(n35717), .B(n27920), .Z(n35716) );
  XOR U36830 ( .A(n35718), .B(\modmult_1/zin[0][469] ), .Z(n27920) );
  IV U36831 ( .A(n35715), .Z(n35718) );
  XNOR U36832 ( .A(n35715), .B(n27919), .Z(n35717) );
  XOR U36833 ( .A(n35719), .B(n35720), .Z(n27919) );
  AND U36834 ( .A(\modmult_1/xin[1023] ), .B(n35721), .Z(n35720) );
  IV U36835 ( .A(n35719), .Z(n35721) );
  XOR U36836 ( .A(n35722), .B(g_input[470]), .Z(n35719) );
  NAND U36837 ( .A(n35723), .B(mul_pow), .Z(n35722) );
  XOR U36838 ( .A(g_input[470]), .B(creg[470]), .Z(n35723) );
  XOR U36839 ( .A(n35724), .B(n35725), .Z(n35715) );
  ANDN U36840 ( .A(n35726), .B(n27926), .Z(n35725) );
  XOR U36841 ( .A(n35727), .B(\modmult_1/zin[0][468] ), .Z(n27926) );
  IV U36842 ( .A(n35724), .Z(n35727) );
  XNOR U36843 ( .A(n35724), .B(n27925), .Z(n35726) );
  XOR U36844 ( .A(n35728), .B(n35729), .Z(n27925) );
  AND U36845 ( .A(\modmult_1/xin[1023] ), .B(n35730), .Z(n35729) );
  IV U36846 ( .A(n35728), .Z(n35730) );
  XOR U36847 ( .A(n35731), .B(g_input[469]), .Z(n35728) );
  NAND U36848 ( .A(n35732), .B(mul_pow), .Z(n35731) );
  XOR U36849 ( .A(g_input[469]), .B(creg[469]), .Z(n35732) );
  XOR U36850 ( .A(n35733), .B(n35734), .Z(n35724) );
  ANDN U36851 ( .A(n35735), .B(n27932), .Z(n35734) );
  XOR U36852 ( .A(n35736), .B(\modmult_1/zin[0][467] ), .Z(n27932) );
  IV U36853 ( .A(n35733), .Z(n35736) );
  XNOR U36854 ( .A(n35733), .B(n27931), .Z(n35735) );
  XOR U36855 ( .A(n35737), .B(n35738), .Z(n27931) );
  AND U36856 ( .A(\modmult_1/xin[1023] ), .B(n35739), .Z(n35738) );
  IV U36857 ( .A(n35737), .Z(n35739) );
  XOR U36858 ( .A(n35740), .B(g_input[468]), .Z(n35737) );
  NAND U36859 ( .A(n35741), .B(mul_pow), .Z(n35740) );
  XOR U36860 ( .A(g_input[468]), .B(creg[468]), .Z(n35741) );
  XOR U36861 ( .A(n35742), .B(n35743), .Z(n35733) );
  ANDN U36862 ( .A(n35744), .B(n27938), .Z(n35743) );
  XOR U36863 ( .A(n35745), .B(\modmult_1/zin[0][466] ), .Z(n27938) );
  IV U36864 ( .A(n35742), .Z(n35745) );
  XNOR U36865 ( .A(n35742), .B(n27937), .Z(n35744) );
  XOR U36866 ( .A(n35746), .B(n35747), .Z(n27937) );
  AND U36867 ( .A(\modmult_1/xin[1023] ), .B(n35748), .Z(n35747) );
  IV U36868 ( .A(n35746), .Z(n35748) );
  XOR U36869 ( .A(n35749), .B(g_input[467]), .Z(n35746) );
  NAND U36870 ( .A(n35750), .B(mul_pow), .Z(n35749) );
  XOR U36871 ( .A(g_input[467]), .B(creg[467]), .Z(n35750) );
  XOR U36872 ( .A(n35751), .B(n35752), .Z(n35742) );
  ANDN U36873 ( .A(n35753), .B(n27944), .Z(n35752) );
  XOR U36874 ( .A(n35754), .B(\modmult_1/zin[0][465] ), .Z(n27944) );
  IV U36875 ( .A(n35751), .Z(n35754) );
  XNOR U36876 ( .A(n35751), .B(n27943), .Z(n35753) );
  XOR U36877 ( .A(n35755), .B(n35756), .Z(n27943) );
  AND U36878 ( .A(\modmult_1/xin[1023] ), .B(n35757), .Z(n35756) );
  IV U36879 ( .A(n35755), .Z(n35757) );
  XOR U36880 ( .A(n35758), .B(g_input[466]), .Z(n35755) );
  NAND U36881 ( .A(n35759), .B(mul_pow), .Z(n35758) );
  XOR U36882 ( .A(g_input[466]), .B(creg[466]), .Z(n35759) );
  XOR U36883 ( .A(n35760), .B(n35761), .Z(n35751) );
  ANDN U36884 ( .A(n35762), .B(n27950), .Z(n35761) );
  XOR U36885 ( .A(n35763), .B(\modmult_1/zin[0][464] ), .Z(n27950) );
  IV U36886 ( .A(n35760), .Z(n35763) );
  XNOR U36887 ( .A(n35760), .B(n27949), .Z(n35762) );
  XOR U36888 ( .A(n35764), .B(n35765), .Z(n27949) );
  AND U36889 ( .A(\modmult_1/xin[1023] ), .B(n35766), .Z(n35765) );
  IV U36890 ( .A(n35764), .Z(n35766) );
  XOR U36891 ( .A(n35767), .B(g_input[465]), .Z(n35764) );
  NAND U36892 ( .A(n35768), .B(mul_pow), .Z(n35767) );
  XOR U36893 ( .A(g_input[465]), .B(creg[465]), .Z(n35768) );
  XOR U36894 ( .A(n35769), .B(n35770), .Z(n35760) );
  ANDN U36895 ( .A(n35771), .B(n27956), .Z(n35770) );
  XOR U36896 ( .A(n35772), .B(\modmult_1/zin[0][463] ), .Z(n27956) );
  IV U36897 ( .A(n35769), .Z(n35772) );
  XNOR U36898 ( .A(n35769), .B(n27955), .Z(n35771) );
  XOR U36899 ( .A(n35773), .B(n35774), .Z(n27955) );
  AND U36900 ( .A(\modmult_1/xin[1023] ), .B(n35775), .Z(n35774) );
  IV U36901 ( .A(n35773), .Z(n35775) );
  XOR U36902 ( .A(n35776), .B(g_input[464]), .Z(n35773) );
  NAND U36903 ( .A(n35777), .B(mul_pow), .Z(n35776) );
  XOR U36904 ( .A(g_input[464]), .B(creg[464]), .Z(n35777) );
  XOR U36905 ( .A(n35778), .B(n35779), .Z(n35769) );
  ANDN U36906 ( .A(n35780), .B(n27962), .Z(n35779) );
  XOR U36907 ( .A(n35781), .B(\modmult_1/zin[0][462] ), .Z(n27962) );
  IV U36908 ( .A(n35778), .Z(n35781) );
  XNOR U36909 ( .A(n35778), .B(n27961), .Z(n35780) );
  XOR U36910 ( .A(n35782), .B(n35783), .Z(n27961) );
  AND U36911 ( .A(\modmult_1/xin[1023] ), .B(n35784), .Z(n35783) );
  IV U36912 ( .A(n35782), .Z(n35784) );
  XOR U36913 ( .A(n35785), .B(g_input[463]), .Z(n35782) );
  NAND U36914 ( .A(n35786), .B(mul_pow), .Z(n35785) );
  XOR U36915 ( .A(g_input[463]), .B(creg[463]), .Z(n35786) );
  XOR U36916 ( .A(n35787), .B(n35788), .Z(n35778) );
  ANDN U36917 ( .A(n35789), .B(n27968), .Z(n35788) );
  XOR U36918 ( .A(n35790), .B(\modmult_1/zin[0][461] ), .Z(n27968) );
  IV U36919 ( .A(n35787), .Z(n35790) );
  XNOR U36920 ( .A(n35787), .B(n27967), .Z(n35789) );
  XOR U36921 ( .A(n35791), .B(n35792), .Z(n27967) );
  AND U36922 ( .A(\modmult_1/xin[1023] ), .B(n35793), .Z(n35792) );
  IV U36923 ( .A(n35791), .Z(n35793) );
  XOR U36924 ( .A(n35794), .B(g_input[462]), .Z(n35791) );
  NAND U36925 ( .A(n35795), .B(mul_pow), .Z(n35794) );
  XOR U36926 ( .A(g_input[462]), .B(creg[462]), .Z(n35795) );
  XOR U36927 ( .A(n35796), .B(n35797), .Z(n35787) );
  ANDN U36928 ( .A(n35798), .B(n27974), .Z(n35797) );
  XOR U36929 ( .A(n35799), .B(\modmult_1/zin[0][460] ), .Z(n27974) );
  IV U36930 ( .A(n35796), .Z(n35799) );
  XNOR U36931 ( .A(n35796), .B(n27973), .Z(n35798) );
  XOR U36932 ( .A(n35800), .B(n35801), .Z(n27973) );
  AND U36933 ( .A(\modmult_1/xin[1023] ), .B(n35802), .Z(n35801) );
  IV U36934 ( .A(n35800), .Z(n35802) );
  XOR U36935 ( .A(n35803), .B(g_input[461]), .Z(n35800) );
  NAND U36936 ( .A(n35804), .B(mul_pow), .Z(n35803) );
  XOR U36937 ( .A(g_input[461]), .B(creg[461]), .Z(n35804) );
  XOR U36938 ( .A(n35805), .B(n35806), .Z(n35796) );
  ANDN U36939 ( .A(n35807), .B(n27980), .Z(n35806) );
  XOR U36940 ( .A(n35808), .B(\modmult_1/zin[0][459] ), .Z(n27980) );
  IV U36941 ( .A(n35805), .Z(n35808) );
  XNOR U36942 ( .A(n35805), .B(n27979), .Z(n35807) );
  XOR U36943 ( .A(n35809), .B(n35810), .Z(n27979) );
  AND U36944 ( .A(\modmult_1/xin[1023] ), .B(n35811), .Z(n35810) );
  IV U36945 ( .A(n35809), .Z(n35811) );
  XOR U36946 ( .A(n35812), .B(g_input[460]), .Z(n35809) );
  NAND U36947 ( .A(n35813), .B(mul_pow), .Z(n35812) );
  XOR U36948 ( .A(g_input[460]), .B(creg[460]), .Z(n35813) );
  XOR U36949 ( .A(n35814), .B(n35815), .Z(n35805) );
  ANDN U36950 ( .A(n35816), .B(n27986), .Z(n35815) );
  XOR U36951 ( .A(n35817), .B(\modmult_1/zin[0][458] ), .Z(n27986) );
  IV U36952 ( .A(n35814), .Z(n35817) );
  XNOR U36953 ( .A(n35814), .B(n27985), .Z(n35816) );
  XOR U36954 ( .A(n35818), .B(n35819), .Z(n27985) );
  AND U36955 ( .A(\modmult_1/xin[1023] ), .B(n35820), .Z(n35819) );
  IV U36956 ( .A(n35818), .Z(n35820) );
  XOR U36957 ( .A(n35821), .B(g_input[459]), .Z(n35818) );
  NAND U36958 ( .A(n35822), .B(mul_pow), .Z(n35821) );
  XOR U36959 ( .A(g_input[459]), .B(creg[459]), .Z(n35822) );
  XOR U36960 ( .A(n35823), .B(n35824), .Z(n35814) );
  ANDN U36961 ( .A(n35825), .B(n27992), .Z(n35824) );
  XOR U36962 ( .A(n35826), .B(\modmult_1/zin[0][457] ), .Z(n27992) );
  IV U36963 ( .A(n35823), .Z(n35826) );
  XNOR U36964 ( .A(n35823), .B(n27991), .Z(n35825) );
  XOR U36965 ( .A(n35827), .B(n35828), .Z(n27991) );
  AND U36966 ( .A(\modmult_1/xin[1023] ), .B(n35829), .Z(n35828) );
  IV U36967 ( .A(n35827), .Z(n35829) );
  XOR U36968 ( .A(n35830), .B(g_input[458]), .Z(n35827) );
  NAND U36969 ( .A(n35831), .B(mul_pow), .Z(n35830) );
  XOR U36970 ( .A(g_input[458]), .B(creg[458]), .Z(n35831) );
  XOR U36971 ( .A(n35832), .B(n35833), .Z(n35823) );
  ANDN U36972 ( .A(n35834), .B(n27998), .Z(n35833) );
  XOR U36973 ( .A(n35835), .B(\modmult_1/zin[0][456] ), .Z(n27998) );
  IV U36974 ( .A(n35832), .Z(n35835) );
  XNOR U36975 ( .A(n35832), .B(n27997), .Z(n35834) );
  XOR U36976 ( .A(n35836), .B(n35837), .Z(n27997) );
  AND U36977 ( .A(\modmult_1/xin[1023] ), .B(n35838), .Z(n35837) );
  IV U36978 ( .A(n35836), .Z(n35838) );
  XOR U36979 ( .A(n35839), .B(g_input[457]), .Z(n35836) );
  NAND U36980 ( .A(n35840), .B(mul_pow), .Z(n35839) );
  XOR U36981 ( .A(g_input[457]), .B(creg[457]), .Z(n35840) );
  XOR U36982 ( .A(n35841), .B(n35842), .Z(n35832) );
  ANDN U36983 ( .A(n35843), .B(n28004), .Z(n35842) );
  XOR U36984 ( .A(n35844), .B(\modmult_1/zin[0][455] ), .Z(n28004) );
  IV U36985 ( .A(n35841), .Z(n35844) );
  XNOR U36986 ( .A(n35841), .B(n28003), .Z(n35843) );
  XOR U36987 ( .A(n35845), .B(n35846), .Z(n28003) );
  AND U36988 ( .A(\modmult_1/xin[1023] ), .B(n35847), .Z(n35846) );
  IV U36989 ( .A(n35845), .Z(n35847) );
  XOR U36990 ( .A(n35848), .B(g_input[456]), .Z(n35845) );
  NAND U36991 ( .A(n35849), .B(mul_pow), .Z(n35848) );
  XOR U36992 ( .A(g_input[456]), .B(creg[456]), .Z(n35849) );
  XOR U36993 ( .A(n35850), .B(n35851), .Z(n35841) );
  ANDN U36994 ( .A(n35852), .B(n28010), .Z(n35851) );
  XOR U36995 ( .A(n35853), .B(\modmult_1/zin[0][454] ), .Z(n28010) );
  IV U36996 ( .A(n35850), .Z(n35853) );
  XNOR U36997 ( .A(n35850), .B(n28009), .Z(n35852) );
  XOR U36998 ( .A(n35854), .B(n35855), .Z(n28009) );
  AND U36999 ( .A(\modmult_1/xin[1023] ), .B(n35856), .Z(n35855) );
  IV U37000 ( .A(n35854), .Z(n35856) );
  XOR U37001 ( .A(n35857), .B(g_input[455]), .Z(n35854) );
  NAND U37002 ( .A(n35858), .B(mul_pow), .Z(n35857) );
  XOR U37003 ( .A(g_input[455]), .B(creg[455]), .Z(n35858) );
  XOR U37004 ( .A(n35859), .B(n35860), .Z(n35850) );
  ANDN U37005 ( .A(n35861), .B(n28016), .Z(n35860) );
  XOR U37006 ( .A(n35862), .B(\modmult_1/zin[0][453] ), .Z(n28016) );
  IV U37007 ( .A(n35859), .Z(n35862) );
  XNOR U37008 ( .A(n35859), .B(n28015), .Z(n35861) );
  XOR U37009 ( .A(n35863), .B(n35864), .Z(n28015) );
  AND U37010 ( .A(\modmult_1/xin[1023] ), .B(n35865), .Z(n35864) );
  IV U37011 ( .A(n35863), .Z(n35865) );
  XOR U37012 ( .A(n35866), .B(g_input[454]), .Z(n35863) );
  NAND U37013 ( .A(n35867), .B(mul_pow), .Z(n35866) );
  XOR U37014 ( .A(g_input[454]), .B(creg[454]), .Z(n35867) );
  XOR U37015 ( .A(n35868), .B(n35869), .Z(n35859) );
  ANDN U37016 ( .A(n35870), .B(n28022), .Z(n35869) );
  XOR U37017 ( .A(n35871), .B(\modmult_1/zin[0][452] ), .Z(n28022) );
  IV U37018 ( .A(n35868), .Z(n35871) );
  XNOR U37019 ( .A(n35868), .B(n28021), .Z(n35870) );
  XOR U37020 ( .A(n35872), .B(n35873), .Z(n28021) );
  AND U37021 ( .A(\modmult_1/xin[1023] ), .B(n35874), .Z(n35873) );
  IV U37022 ( .A(n35872), .Z(n35874) );
  XOR U37023 ( .A(n35875), .B(g_input[453]), .Z(n35872) );
  NAND U37024 ( .A(n35876), .B(mul_pow), .Z(n35875) );
  XOR U37025 ( .A(g_input[453]), .B(creg[453]), .Z(n35876) );
  XOR U37026 ( .A(n35877), .B(n35878), .Z(n35868) );
  ANDN U37027 ( .A(n35879), .B(n28028), .Z(n35878) );
  XOR U37028 ( .A(n35880), .B(\modmult_1/zin[0][451] ), .Z(n28028) );
  IV U37029 ( .A(n35877), .Z(n35880) );
  XNOR U37030 ( .A(n35877), .B(n28027), .Z(n35879) );
  XOR U37031 ( .A(n35881), .B(n35882), .Z(n28027) );
  AND U37032 ( .A(\modmult_1/xin[1023] ), .B(n35883), .Z(n35882) );
  IV U37033 ( .A(n35881), .Z(n35883) );
  XOR U37034 ( .A(n35884), .B(g_input[452]), .Z(n35881) );
  NAND U37035 ( .A(n35885), .B(mul_pow), .Z(n35884) );
  XOR U37036 ( .A(g_input[452]), .B(creg[452]), .Z(n35885) );
  XOR U37037 ( .A(n35886), .B(n35887), .Z(n35877) );
  ANDN U37038 ( .A(n35888), .B(n28034), .Z(n35887) );
  XOR U37039 ( .A(n35889), .B(\modmult_1/zin[0][450] ), .Z(n28034) );
  IV U37040 ( .A(n35886), .Z(n35889) );
  XNOR U37041 ( .A(n35886), .B(n28033), .Z(n35888) );
  XOR U37042 ( .A(n35890), .B(n35891), .Z(n28033) );
  AND U37043 ( .A(\modmult_1/xin[1023] ), .B(n35892), .Z(n35891) );
  IV U37044 ( .A(n35890), .Z(n35892) );
  XOR U37045 ( .A(n35893), .B(g_input[451]), .Z(n35890) );
  NAND U37046 ( .A(n35894), .B(mul_pow), .Z(n35893) );
  XOR U37047 ( .A(g_input[451]), .B(creg[451]), .Z(n35894) );
  XOR U37048 ( .A(n35895), .B(n35896), .Z(n35886) );
  ANDN U37049 ( .A(n35897), .B(n28040), .Z(n35896) );
  XOR U37050 ( .A(n35898), .B(\modmult_1/zin[0][449] ), .Z(n28040) );
  IV U37051 ( .A(n35895), .Z(n35898) );
  XNOR U37052 ( .A(n35895), .B(n28039), .Z(n35897) );
  XOR U37053 ( .A(n35899), .B(n35900), .Z(n28039) );
  AND U37054 ( .A(\modmult_1/xin[1023] ), .B(n35901), .Z(n35900) );
  IV U37055 ( .A(n35899), .Z(n35901) );
  XOR U37056 ( .A(n35902), .B(g_input[450]), .Z(n35899) );
  NAND U37057 ( .A(n35903), .B(mul_pow), .Z(n35902) );
  XOR U37058 ( .A(g_input[450]), .B(creg[450]), .Z(n35903) );
  XOR U37059 ( .A(n35904), .B(n35905), .Z(n35895) );
  ANDN U37060 ( .A(n35906), .B(n28046), .Z(n35905) );
  XOR U37061 ( .A(n35907), .B(\modmult_1/zin[0][448] ), .Z(n28046) );
  IV U37062 ( .A(n35904), .Z(n35907) );
  XNOR U37063 ( .A(n35904), .B(n28045), .Z(n35906) );
  XOR U37064 ( .A(n35908), .B(n35909), .Z(n28045) );
  AND U37065 ( .A(\modmult_1/xin[1023] ), .B(n35910), .Z(n35909) );
  IV U37066 ( .A(n35908), .Z(n35910) );
  XOR U37067 ( .A(n35911), .B(g_input[449]), .Z(n35908) );
  NAND U37068 ( .A(n35912), .B(mul_pow), .Z(n35911) );
  XOR U37069 ( .A(g_input[449]), .B(creg[449]), .Z(n35912) );
  XOR U37070 ( .A(n35913), .B(n35914), .Z(n35904) );
  ANDN U37071 ( .A(n35915), .B(n28052), .Z(n35914) );
  XOR U37072 ( .A(n35916), .B(\modmult_1/zin[0][447] ), .Z(n28052) );
  IV U37073 ( .A(n35913), .Z(n35916) );
  XNOR U37074 ( .A(n35913), .B(n28051), .Z(n35915) );
  XOR U37075 ( .A(n35917), .B(n35918), .Z(n28051) );
  AND U37076 ( .A(\modmult_1/xin[1023] ), .B(n35919), .Z(n35918) );
  IV U37077 ( .A(n35917), .Z(n35919) );
  XOR U37078 ( .A(n35920), .B(g_input[448]), .Z(n35917) );
  NAND U37079 ( .A(n35921), .B(mul_pow), .Z(n35920) );
  XOR U37080 ( .A(g_input[448]), .B(creg[448]), .Z(n35921) );
  XOR U37081 ( .A(n35922), .B(n35923), .Z(n35913) );
  ANDN U37082 ( .A(n35924), .B(n28058), .Z(n35923) );
  XOR U37083 ( .A(n35925), .B(\modmult_1/zin[0][446] ), .Z(n28058) );
  IV U37084 ( .A(n35922), .Z(n35925) );
  XNOR U37085 ( .A(n35922), .B(n28057), .Z(n35924) );
  XOR U37086 ( .A(n35926), .B(n35927), .Z(n28057) );
  AND U37087 ( .A(\modmult_1/xin[1023] ), .B(n35928), .Z(n35927) );
  IV U37088 ( .A(n35926), .Z(n35928) );
  XOR U37089 ( .A(n35929), .B(g_input[447]), .Z(n35926) );
  NAND U37090 ( .A(n35930), .B(mul_pow), .Z(n35929) );
  XOR U37091 ( .A(g_input[447]), .B(creg[447]), .Z(n35930) );
  XOR U37092 ( .A(n35931), .B(n35932), .Z(n35922) );
  ANDN U37093 ( .A(n35933), .B(n28064), .Z(n35932) );
  XOR U37094 ( .A(n35934), .B(\modmult_1/zin[0][445] ), .Z(n28064) );
  IV U37095 ( .A(n35931), .Z(n35934) );
  XNOR U37096 ( .A(n35931), .B(n28063), .Z(n35933) );
  XOR U37097 ( .A(n35935), .B(n35936), .Z(n28063) );
  AND U37098 ( .A(\modmult_1/xin[1023] ), .B(n35937), .Z(n35936) );
  IV U37099 ( .A(n35935), .Z(n35937) );
  XOR U37100 ( .A(n35938), .B(g_input[446]), .Z(n35935) );
  NAND U37101 ( .A(n35939), .B(mul_pow), .Z(n35938) );
  XOR U37102 ( .A(g_input[446]), .B(creg[446]), .Z(n35939) );
  XOR U37103 ( .A(n35940), .B(n35941), .Z(n35931) );
  ANDN U37104 ( .A(n35942), .B(n28070), .Z(n35941) );
  XOR U37105 ( .A(n35943), .B(\modmult_1/zin[0][444] ), .Z(n28070) );
  IV U37106 ( .A(n35940), .Z(n35943) );
  XNOR U37107 ( .A(n35940), .B(n28069), .Z(n35942) );
  XOR U37108 ( .A(n35944), .B(n35945), .Z(n28069) );
  AND U37109 ( .A(\modmult_1/xin[1023] ), .B(n35946), .Z(n35945) );
  IV U37110 ( .A(n35944), .Z(n35946) );
  XOR U37111 ( .A(n35947), .B(g_input[445]), .Z(n35944) );
  NAND U37112 ( .A(n35948), .B(mul_pow), .Z(n35947) );
  XOR U37113 ( .A(g_input[445]), .B(creg[445]), .Z(n35948) );
  XOR U37114 ( .A(n35949), .B(n35950), .Z(n35940) );
  ANDN U37115 ( .A(n35951), .B(n28076), .Z(n35950) );
  XOR U37116 ( .A(n35952), .B(\modmult_1/zin[0][443] ), .Z(n28076) );
  IV U37117 ( .A(n35949), .Z(n35952) );
  XNOR U37118 ( .A(n35949), .B(n28075), .Z(n35951) );
  XOR U37119 ( .A(n35953), .B(n35954), .Z(n28075) );
  AND U37120 ( .A(\modmult_1/xin[1023] ), .B(n35955), .Z(n35954) );
  IV U37121 ( .A(n35953), .Z(n35955) );
  XOR U37122 ( .A(n35956), .B(g_input[444]), .Z(n35953) );
  NAND U37123 ( .A(n35957), .B(mul_pow), .Z(n35956) );
  XOR U37124 ( .A(g_input[444]), .B(creg[444]), .Z(n35957) );
  XOR U37125 ( .A(n35958), .B(n35959), .Z(n35949) );
  ANDN U37126 ( .A(n35960), .B(n28082), .Z(n35959) );
  XOR U37127 ( .A(n35961), .B(\modmult_1/zin[0][442] ), .Z(n28082) );
  IV U37128 ( .A(n35958), .Z(n35961) );
  XNOR U37129 ( .A(n35958), .B(n28081), .Z(n35960) );
  XOR U37130 ( .A(n35962), .B(n35963), .Z(n28081) );
  AND U37131 ( .A(\modmult_1/xin[1023] ), .B(n35964), .Z(n35963) );
  IV U37132 ( .A(n35962), .Z(n35964) );
  XOR U37133 ( .A(n35965), .B(g_input[443]), .Z(n35962) );
  NAND U37134 ( .A(n35966), .B(mul_pow), .Z(n35965) );
  XOR U37135 ( .A(g_input[443]), .B(creg[443]), .Z(n35966) );
  XOR U37136 ( .A(n35967), .B(n35968), .Z(n35958) );
  ANDN U37137 ( .A(n35969), .B(n28088), .Z(n35968) );
  XOR U37138 ( .A(n35970), .B(\modmult_1/zin[0][441] ), .Z(n28088) );
  IV U37139 ( .A(n35967), .Z(n35970) );
  XNOR U37140 ( .A(n35967), .B(n28087), .Z(n35969) );
  XOR U37141 ( .A(n35971), .B(n35972), .Z(n28087) );
  AND U37142 ( .A(\modmult_1/xin[1023] ), .B(n35973), .Z(n35972) );
  IV U37143 ( .A(n35971), .Z(n35973) );
  XOR U37144 ( .A(n35974), .B(g_input[442]), .Z(n35971) );
  NAND U37145 ( .A(n35975), .B(mul_pow), .Z(n35974) );
  XOR U37146 ( .A(g_input[442]), .B(creg[442]), .Z(n35975) );
  XOR U37147 ( .A(n35976), .B(n35977), .Z(n35967) );
  ANDN U37148 ( .A(n35978), .B(n28094), .Z(n35977) );
  XOR U37149 ( .A(n35979), .B(\modmult_1/zin[0][440] ), .Z(n28094) );
  IV U37150 ( .A(n35976), .Z(n35979) );
  XNOR U37151 ( .A(n35976), .B(n28093), .Z(n35978) );
  XOR U37152 ( .A(n35980), .B(n35981), .Z(n28093) );
  AND U37153 ( .A(\modmult_1/xin[1023] ), .B(n35982), .Z(n35981) );
  IV U37154 ( .A(n35980), .Z(n35982) );
  XOR U37155 ( .A(n35983), .B(g_input[441]), .Z(n35980) );
  NAND U37156 ( .A(n35984), .B(mul_pow), .Z(n35983) );
  XOR U37157 ( .A(g_input[441]), .B(creg[441]), .Z(n35984) );
  XOR U37158 ( .A(n35985), .B(n35986), .Z(n35976) );
  ANDN U37159 ( .A(n35987), .B(n28100), .Z(n35986) );
  XOR U37160 ( .A(n35988), .B(\modmult_1/zin[0][439] ), .Z(n28100) );
  IV U37161 ( .A(n35985), .Z(n35988) );
  XNOR U37162 ( .A(n35985), .B(n28099), .Z(n35987) );
  XOR U37163 ( .A(n35989), .B(n35990), .Z(n28099) );
  AND U37164 ( .A(\modmult_1/xin[1023] ), .B(n35991), .Z(n35990) );
  IV U37165 ( .A(n35989), .Z(n35991) );
  XOR U37166 ( .A(n35992), .B(g_input[440]), .Z(n35989) );
  NAND U37167 ( .A(n35993), .B(mul_pow), .Z(n35992) );
  XOR U37168 ( .A(g_input[440]), .B(creg[440]), .Z(n35993) );
  XOR U37169 ( .A(n35994), .B(n35995), .Z(n35985) );
  ANDN U37170 ( .A(n35996), .B(n28106), .Z(n35995) );
  XOR U37171 ( .A(n35997), .B(\modmult_1/zin[0][438] ), .Z(n28106) );
  IV U37172 ( .A(n35994), .Z(n35997) );
  XNOR U37173 ( .A(n35994), .B(n28105), .Z(n35996) );
  XOR U37174 ( .A(n35998), .B(n35999), .Z(n28105) );
  AND U37175 ( .A(\modmult_1/xin[1023] ), .B(n36000), .Z(n35999) );
  IV U37176 ( .A(n35998), .Z(n36000) );
  XOR U37177 ( .A(n36001), .B(g_input[439]), .Z(n35998) );
  NAND U37178 ( .A(n36002), .B(mul_pow), .Z(n36001) );
  XOR U37179 ( .A(g_input[439]), .B(creg[439]), .Z(n36002) );
  XOR U37180 ( .A(n36003), .B(n36004), .Z(n35994) );
  ANDN U37181 ( .A(n36005), .B(n28112), .Z(n36004) );
  XOR U37182 ( .A(n36006), .B(\modmult_1/zin[0][437] ), .Z(n28112) );
  IV U37183 ( .A(n36003), .Z(n36006) );
  XNOR U37184 ( .A(n36003), .B(n28111), .Z(n36005) );
  XOR U37185 ( .A(n36007), .B(n36008), .Z(n28111) );
  AND U37186 ( .A(\modmult_1/xin[1023] ), .B(n36009), .Z(n36008) );
  IV U37187 ( .A(n36007), .Z(n36009) );
  XOR U37188 ( .A(n36010), .B(g_input[438]), .Z(n36007) );
  NAND U37189 ( .A(n36011), .B(mul_pow), .Z(n36010) );
  XOR U37190 ( .A(g_input[438]), .B(creg[438]), .Z(n36011) );
  XOR U37191 ( .A(n36012), .B(n36013), .Z(n36003) );
  ANDN U37192 ( .A(n36014), .B(n28118), .Z(n36013) );
  XOR U37193 ( .A(n36015), .B(\modmult_1/zin[0][436] ), .Z(n28118) );
  IV U37194 ( .A(n36012), .Z(n36015) );
  XNOR U37195 ( .A(n36012), .B(n28117), .Z(n36014) );
  XOR U37196 ( .A(n36016), .B(n36017), .Z(n28117) );
  AND U37197 ( .A(\modmult_1/xin[1023] ), .B(n36018), .Z(n36017) );
  IV U37198 ( .A(n36016), .Z(n36018) );
  XOR U37199 ( .A(n36019), .B(g_input[437]), .Z(n36016) );
  NAND U37200 ( .A(n36020), .B(mul_pow), .Z(n36019) );
  XOR U37201 ( .A(g_input[437]), .B(creg[437]), .Z(n36020) );
  XOR U37202 ( .A(n36021), .B(n36022), .Z(n36012) );
  ANDN U37203 ( .A(n36023), .B(n28124), .Z(n36022) );
  XOR U37204 ( .A(n36024), .B(\modmult_1/zin[0][435] ), .Z(n28124) );
  IV U37205 ( .A(n36021), .Z(n36024) );
  XNOR U37206 ( .A(n36021), .B(n28123), .Z(n36023) );
  XOR U37207 ( .A(n36025), .B(n36026), .Z(n28123) );
  AND U37208 ( .A(\modmult_1/xin[1023] ), .B(n36027), .Z(n36026) );
  IV U37209 ( .A(n36025), .Z(n36027) );
  XOR U37210 ( .A(n36028), .B(g_input[436]), .Z(n36025) );
  NAND U37211 ( .A(n36029), .B(mul_pow), .Z(n36028) );
  XOR U37212 ( .A(g_input[436]), .B(creg[436]), .Z(n36029) );
  XOR U37213 ( .A(n36030), .B(n36031), .Z(n36021) );
  ANDN U37214 ( .A(n36032), .B(n28130), .Z(n36031) );
  XOR U37215 ( .A(n36033), .B(\modmult_1/zin[0][434] ), .Z(n28130) );
  IV U37216 ( .A(n36030), .Z(n36033) );
  XNOR U37217 ( .A(n36030), .B(n28129), .Z(n36032) );
  XOR U37218 ( .A(n36034), .B(n36035), .Z(n28129) );
  AND U37219 ( .A(\modmult_1/xin[1023] ), .B(n36036), .Z(n36035) );
  IV U37220 ( .A(n36034), .Z(n36036) );
  XOR U37221 ( .A(n36037), .B(g_input[435]), .Z(n36034) );
  NAND U37222 ( .A(n36038), .B(mul_pow), .Z(n36037) );
  XOR U37223 ( .A(g_input[435]), .B(creg[435]), .Z(n36038) );
  XOR U37224 ( .A(n36039), .B(n36040), .Z(n36030) );
  ANDN U37225 ( .A(n36041), .B(n28136), .Z(n36040) );
  XOR U37226 ( .A(n36042), .B(\modmult_1/zin[0][433] ), .Z(n28136) );
  IV U37227 ( .A(n36039), .Z(n36042) );
  XNOR U37228 ( .A(n36039), .B(n28135), .Z(n36041) );
  XOR U37229 ( .A(n36043), .B(n36044), .Z(n28135) );
  AND U37230 ( .A(\modmult_1/xin[1023] ), .B(n36045), .Z(n36044) );
  IV U37231 ( .A(n36043), .Z(n36045) );
  XOR U37232 ( .A(n36046), .B(g_input[434]), .Z(n36043) );
  NAND U37233 ( .A(n36047), .B(mul_pow), .Z(n36046) );
  XOR U37234 ( .A(g_input[434]), .B(creg[434]), .Z(n36047) );
  XOR U37235 ( .A(n36048), .B(n36049), .Z(n36039) );
  ANDN U37236 ( .A(n36050), .B(n28142), .Z(n36049) );
  XOR U37237 ( .A(n36051), .B(\modmult_1/zin[0][432] ), .Z(n28142) );
  IV U37238 ( .A(n36048), .Z(n36051) );
  XNOR U37239 ( .A(n36048), .B(n28141), .Z(n36050) );
  XOR U37240 ( .A(n36052), .B(n36053), .Z(n28141) );
  AND U37241 ( .A(\modmult_1/xin[1023] ), .B(n36054), .Z(n36053) );
  IV U37242 ( .A(n36052), .Z(n36054) );
  XOR U37243 ( .A(n36055), .B(g_input[433]), .Z(n36052) );
  NAND U37244 ( .A(n36056), .B(mul_pow), .Z(n36055) );
  XOR U37245 ( .A(g_input[433]), .B(creg[433]), .Z(n36056) );
  XOR U37246 ( .A(n36057), .B(n36058), .Z(n36048) );
  ANDN U37247 ( .A(n36059), .B(n28148), .Z(n36058) );
  XOR U37248 ( .A(n36060), .B(\modmult_1/zin[0][431] ), .Z(n28148) );
  IV U37249 ( .A(n36057), .Z(n36060) );
  XNOR U37250 ( .A(n36057), .B(n28147), .Z(n36059) );
  XOR U37251 ( .A(n36061), .B(n36062), .Z(n28147) );
  AND U37252 ( .A(\modmult_1/xin[1023] ), .B(n36063), .Z(n36062) );
  IV U37253 ( .A(n36061), .Z(n36063) );
  XOR U37254 ( .A(n36064), .B(g_input[432]), .Z(n36061) );
  NAND U37255 ( .A(n36065), .B(mul_pow), .Z(n36064) );
  XOR U37256 ( .A(g_input[432]), .B(creg[432]), .Z(n36065) );
  XOR U37257 ( .A(n36066), .B(n36067), .Z(n36057) );
  ANDN U37258 ( .A(n36068), .B(n28154), .Z(n36067) );
  XOR U37259 ( .A(n36069), .B(\modmult_1/zin[0][430] ), .Z(n28154) );
  IV U37260 ( .A(n36066), .Z(n36069) );
  XNOR U37261 ( .A(n36066), .B(n28153), .Z(n36068) );
  XOR U37262 ( .A(n36070), .B(n36071), .Z(n28153) );
  AND U37263 ( .A(\modmult_1/xin[1023] ), .B(n36072), .Z(n36071) );
  IV U37264 ( .A(n36070), .Z(n36072) );
  XOR U37265 ( .A(n36073), .B(g_input[431]), .Z(n36070) );
  NAND U37266 ( .A(n36074), .B(mul_pow), .Z(n36073) );
  XOR U37267 ( .A(g_input[431]), .B(creg[431]), .Z(n36074) );
  XOR U37268 ( .A(n36075), .B(n36076), .Z(n36066) );
  ANDN U37269 ( .A(n36077), .B(n28160), .Z(n36076) );
  XOR U37270 ( .A(n36078), .B(\modmult_1/zin[0][429] ), .Z(n28160) );
  IV U37271 ( .A(n36075), .Z(n36078) );
  XNOR U37272 ( .A(n36075), .B(n28159), .Z(n36077) );
  XOR U37273 ( .A(n36079), .B(n36080), .Z(n28159) );
  AND U37274 ( .A(\modmult_1/xin[1023] ), .B(n36081), .Z(n36080) );
  IV U37275 ( .A(n36079), .Z(n36081) );
  XOR U37276 ( .A(n36082), .B(g_input[430]), .Z(n36079) );
  NAND U37277 ( .A(n36083), .B(mul_pow), .Z(n36082) );
  XOR U37278 ( .A(g_input[430]), .B(creg[430]), .Z(n36083) );
  XOR U37279 ( .A(n36084), .B(n36085), .Z(n36075) );
  ANDN U37280 ( .A(n36086), .B(n28166), .Z(n36085) );
  XOR U37281 ( .A(n36087), .B(\modmult_1/zin[0][428] ), .Z(n28166) );
  IV U37282 ( .A(n36084), .Z(n36087) );
  XNOR U37283 ( .A(n36084), .B(n28165), .Z(n36086) );
  XOR U37284 ( .A(n36088), .B(n36089), .Z(n28165) );
  AND U37285 ( .A(\modmult_1/xin[1023] ), .B(n36090), .Z(n36089) );
  IV U37286 ( .A(n36088), .Z(n36090) );
  XOR U37287 ( .A(n36091), .B(g_input[429]), .Z(n36088) );
  NAND U37288 ( .A(n36092), .B(mul_pow), .Z(n36091) );
  XOR U37289 ( .A(g_input[429]), .B(creg[429]), .Z(n36092) );
  XOR U37290 ( .A(n36093), .B(n36094), .Z(n36084) );
  ANDN U37291 ( .A(n36095), .B(n28172), .Z(n36094) );
  XOR U37292 ( .A(n36096), .B(\modmult_1/zin[0][427] ), .Z(n28172) );
  IV U37293 ( .A(n36093), .Z(n36096) );
  XNOR U37294 ( .A(n36093), .B(n28171), .Z(n36095) );
  XOR U37295 ( .A(n36097), .B(n36098), .Z(n28171) );
  AND U37296 ( .A(\modmult_1/xin[1023] ), .B(n36099), .Z(n36098) );
  IV U37297 ( .A(n36097), .Z(n36099) );
  XOR U37298 ( .A(n36100), .B(g_input[428]), .Z(n36097) );
  NAND U37299 ( .A(n36101), .B(mul_pow), .Z(n36100) );
  XOR U37300 ( .A(g_input[428]), .B(creg[428]), .Z(n36101) );
  XOR U37301 ( .A(n36102), .B(n36103), .Z(n36093) );
  ANDN U37302 ( .A(n36104), .B(n28178), .Z(n36103) );
  XOR U37303 ( .A(n36105), .B(\modmult_1/zin[0][426] ), .Z(n28178) );
  IV U37304 ( .A(n36102), .Z(n36105) );
  XNOR U37305 ( .A(n36102), .B(n28177), .Z(n36104) );
  XOR U37306 ( .A(n36106), .B(n36107), .Z(n28177) );
  AND U37307 ( .A(\modmult_1/xin[1023] ), .B(n36108), .Z(n36107) );
  IV U37308 ( .A(n36106), .Z(n36108) );
  XOR U37309 ( .A(n36109), .B(g_input[427]), .Z(n36106) );
  NAND U37310 ( .A(n36110), .B(mul_pow), .Z(n36109) );
  XOR U37311 ( .A(g_input[427]), .B(creg[427]), .Z(n36110) );
  XOR U37312 ( .A(n36111), .B(n36112), .Z(n36102) );
  ANDN U37313 ( .A(n36113), .B(n28184), .Z(n36112) );
  XOR U37314 ( .A(n36114), .B(\modmult_1/zin[0][425] ), .Z(n28184) );
  IV U37315 ( .A(n36111), .Z(n36114) );
  XNOR U37316 ( .A(n36111), .B(n28183), .Z(n36113) );
  XOR U37317 ( .A(n36115), .B(n36116), .Z(n28183) );
  AND U37318 ( .A(\modmult_1/xin[1023] ), .B(n36117), .Z(n36116) );
  IV U37319 ( .A(n36115), .Z(n36117) );
  XOR U37320 ( .A(n36118), .B(g_input[426]), .Z(n36115) );
  NAND U37321 ( .A(n36119), .B(mul_pow), .Z(n36118) );
  XOR U37322 ( .A(g_input[426]), .B(creg[426]), .Z(n36119) );
  XOR U37323 ( .A(n36120), .B(n36121), .Z(n36111) );
  ANDN U37324 ( .A(n36122), .B(n28190), .Z(n36121) );
  XOR U37325 ( .A(n36123), .B(\modmult_1/zin[0][424] ), .Z(n28190) );
  IV U37326 ( .A(n36120), .Z(n36123) );
  XNOR U37327 ( .A(n36120), .B(n28189), .Z(n36122) );
  XOR U37328 ( .A(n36124), .B(n36125), .Z(n28189) );
  AND U37329 ( .A(\modmult_1/xin[1023] ), .B(n36126), .Z(n36125) );
  IV U37330 ( .A(n36124), .Z(n36126) );
  XOR U37331 ( .A(n36127), .B(g_input[425]), .Z(n36124) );
  NAND U37332 ( .A(n36128), .B(mul_pow), .Z(n36127) );
  XOR U37333 ( .A(g_input[425]), .B(creg[425]), .Z(n36128) );
  XOR U37334 ( .A(n36129), .B(n36130), .Z(n36120) );
  ANDN U37335 ( .A(n36131), .B(n28196), .Z(n36130) );
  XOR U37336 ( .A(n36132), .B(\modmult_1/zin[0][423] ), .Z(n28196) );
  IV U37337 ( .A(n36129), .Z(n36132) );
  XNOR U37338 ( .A(n36129), .B(n28195), .Z(n36131) );
  XOR U37339 ( .A(n36133), .B(n36134), .Z(n28195) );
  AND U37340 ( .A(\modmult_1/xin[1023] ), .B(n36135), .Z(n36134) );
  IV U37341 ( .A(n36133), .Z(n36135) );
  XOR U37342 ( .A(n36136), .B(g_input[424]), .Z(n36133) );
  NAND U37343 ( .A(n36137), .B(mul_pow), .Z(n36136) );
  XOR U37344 ( .A(g_input[424]), .B(creg[424]), .Z(n36137) );
  XOR U37345 ( .A(n36138), .B(n36139), .Z(n36129) );
  ANDN U37346 ( .A(n36140), .B(n28202), .Z(n36139) );
  XOR U37347 ( .A(n36141), .B(\modmult_1/zin[0][422] ), .Z(n28202) );
  IV U37348 ( .A(n36138), .Z(n36141) );
  XNOR U37349 ( .A(n36138), .B(n28201), .Z(n36140) );
  XOR U37350 ( .A(n36142), .B(n36143), .Z(n28201) );
  AND U37351 ( .A(\modmult_1/xin[1023] ), .B(n36144), .Z(n36143) );
  IV U37352 ( .A(n36142), .Z(n36144) );
  XOR U37353 ( .A(n36145), .B(g_input[423]), .Z(n36142) );
  NAND U37354 ( .A(n36146), .B(mul_pow), .Z(n36145) );
  XOR U37355 ( .A(g_input[423]), .B(creg[423]), .Z(n36146) );
  XOR U37356 ( .A(n36147), .B(n36148), .Z(n36138) );
  ANDN U37357 ( .A(n36149), .B(n28208), .Z(n36148) );
  XOR U37358 ( .A(n36150), .B(\modmult_1/zin[0][421] ), .Z(n28208) );
  IV U37359 ( .A(n36147), .Z(n36150) );
  XNOR U37360 ( .A(n36147), .B(n28207), .Z(n36149) );
  XOR U37361 ( .A(n36151), .B(n36152), .Z(n28207) );
  AND U37362 ( .A(\modmult_1/xin[1023] ), .B(n36153), .Z(n36152) );
  IV U37363 ( .A(n36151), .Z(n36153) );
  XOR U37364 ( .A(n36154), .B(g_input[422]), .Z(n36151) );
  NAND U37365 ( .A(n36155), .B(mul_pow), .Z(n36154) );
  XOR U37366 ( .A(g_input[422]), .B(creg[422]), .Z(n36155) );
  XOR U37367 ( .A(n36156), .B(n36157), .Z(n36147) );
  ANDN U37368 ( .A(n36158), .B(n28214), .Z(n36157) );
  XOR U37369 ( .A(n36159), .B(\modmult_1/zin[0][420] ), .Z(n28214) );
  IV U37370 ( .A(n36156), .Z(n36159) );
  XNOR U37371 ( .A(n36156), .B(n28213), .Z(n36158) );
  XOR U37372 ( .A(n36160), .B(n36161), .Z(n28213) );
  AND U37373 ( .A(\modmult_1/xin[1023] ), .B(n36162), .Z(n36161) );
  IV U37374 ( .A(n36160), .Z(n36162) );
  XOR U37375 ( .A(n36163), .B(g_input[421]), .Z(n36160) );
  NAND U37376 ( .A(n36164), .B(mul_pow), .Z(n36163) );
  XOR U37377 ( .A(g_input[421]), .B(creg[421]), .Z(n36164) );
  XOR U37378 ( .A(n36165), .B(n36166), .Z(n36156) );
  ANDN U37379 ( .A(n36167), .B(n28220), .Z(n36166) );
  XOR U37380 ( .A(n36168), .B(\modmult_1/zin[0][419] ), .Z(n28220) );
  IV U37381 ( .A(n36165), .Z(n36168) );
  XNOR U37382 ( .A(n36165), .B(n28219), .Z(n36167) );
  XOR U37383 ( .A(n36169), .B(n36170), .Z(n28219) );
  AND U37384 ( .A(\modmult_1/xin[1023] ), .B(n36171), .Z(n36170) );
  IV U37385 ( .A(n36169), .Z(n36171) );
  XOR U37386 ( .A(n36172), .B(g_input[420]), .Z(n36169) );
  NAND U37387 ( .A(n36173), .B(mul_pow), .Z(n36172) );
  XOR U37388 ( .A(g_input[420]), .B(creg[420]), .Z(n36173) );
  XOR U37389 ( .A(n36174), .B(n36175), .Z(n36165) );
  ANDN U37390 ( .A(n36176), .B(n28226), .Z(n36175) );
  XOR U37391 ( .A(n36177), .B(\modmult_1/zin[0][418] ), .Z(n28226) );
  IV U37392 ( .A(n36174), .Z(n36177) );
  XNOR U37393 ( .A(n36174), .B(n28225), .Z(n36176) );
  XOR U37394 ( .A(n36178), .B(n36179), .Z(n28225) );
  AND U37395 ( .A(\modmult_1/xin[1023] ), .B(n36180), .Z(n36179) );
  IV U37396 ( .A(n36178), .Z(n36180) );
  XOR U37397 ( .A(n36181), .B(g_input[419]), .Z(n36178) );
  NAND U37398 ( .A(n36182), .B(mul_pow), .Z(n36181) );
  XOR U37399 ( .A(g_input[419]), .B(creg[419]), .Z(n36182) );
  XOR U37400 ( .A(n36183), .B(n36184), .Z(n36174) );
  ANDN U37401 ( .A(n36185), .B(n28232), .Z(n36184) );
  XOR U37402 ( .A(n36186), .B(\modmult_1/zin[0][417] ), .Z(n28232) );
  IV U37403 ( .A(n36183), .Z(n36186) );
  XNOR U37404 ( .A(n36183), .B(n28231), .Z(n36185) );
  XOR U37405 ( .A(n36187), .B(n36188), .Z(n28231) );
  AND U37406 ( .A(\modmult_1/xin[1023] ), .B(n36189), .Z(n36188) );
  IV U37407 ( .A(n36187), .Z(n36189) );
  XOR U37408 ( .A(n36190), .B(g_input[418]), .Z(n36187) );
  NAND U37409 ( .A(n36191), .B(mul_pow), .Z(n36190) );
  XOR U37410 ( .A(g_input[418]), .B(creg[418]), .Z(n36191) );
  XOR U37411 ( .A(n36192), .B(n36193), .Z(n36183) );
  ANDN U37412 ( .A(n36194), .B(n28238), .Z(n36193) );
  XOR U37413 ( .A(n36195), .B(\modmult_1/zin[0][416] ), .Z(n28238) );
  IV U37414 ( .A(n36192), .Z(n36195) );
  XNOR U37415 ( .A(n36192), .B(n28237), .Z(n36194) );
  XOR U37416 ( .A(n36196), .B(n36197), .Z(n28237) );
  AND U37417 ( .A(\modmult_1/xin[1023] ), .B(n36198), .Z(n36197) );
  IV U37418 ( .A(n36196), .Z(n36198) );
  XOR U37419 ( .A(n36199), .B(g_input[417]), .Z(n36196) );
  NAND U37420 ( .A(n36200), .B(mul_pow), .Z(n36199) );
  XOR U37421 ( .A(g_input[417]), .B(creg[417]), .Z(n36200) );
  XOR U37422 ( .A(n36201), .B(n36202), .Z(n36192) );
  ANDN U37423 ( .A(n36203), .B(n28244), .Z(n36202) );
  XOR U37424 ( .A(n36204), .B(\modmult_1/zin[0][415] ), .Z(n28244) );
  IV U37425 ( .A(n36201), .Z(n36204) );
  XNOR U37426 ( .A(n36201), .B(n28243), .Z(n36203) );
  XOR U37427 ( .A(n36205), .B(n36206), .Z(n28243) );
  AND U37428 ( .A(\modmult_1/xin[1023] ), .B(n36207), .Z(n36206) );
  IV U37429 ( .A(n36205), .Z(n36207) );
  XOR U37430 ( .A(n36208), .B(g_input[416]), .Z(n36205) );
  NAND U37431 ( .A(n36209), .B(mul_pow), .Z(n36208) );
  XOR U37432 ( .A(g_input[416]), .B(creg[416]), .Z(n36209) );
  XOR U37433 ( .A(n36210), .B(n36211), .Z(n36201) );
  ANDN U37434 ( .A(n36212), .B(n28250), .Z(n36211) );
  XOR U37435 ( .A(n36213), .B(\modmult_1/zin[0][414] ), .Z(n28250) );
  IV U37436 ( .A(n36210), .Z(n36213) );
  XNOR U37437 ( .A(n36210), .B(n28249), .Z(n36212) );
  XOR U37438 ( .A(n36214), .B(n36215), .Z(n28249) );
  AND U37439 ( .A(\modmult_1/xin[1023] ), .B(n36216), .Z(n36215) );
  IV U37440 ( .A(n36214), .Z(n36216) );
  XOR U37441 ( .A(n36217), .B(g_input[415]), .Z(n36214) );
  NAND U37442 ( .A(n36218), .B(mul_pow), .Z(n36217) );
  XOR U37443 ( .A(g_input[415]), .B(creg[415]), .Z(n36218) );
  XOR U37444 ( .A(n36219), .B(n36220), .Z(n36210) );
  ANDN U37445 ( .A(n36221), .B(n28256), .Z(n36220) );
  XOR U37446 ( .A(n36222), .B(\modmult_1/zin[0][413] ), .Z(n28256) );
  IV U37447 ( .A(n36219), .Z(n36222) );
  XNOR U37448 ( .A(n36219), .B(n28255), .Z(n36221) );
  XOR U37449 ( .A(n36223), .B(n36224), .Z(n28255) );
  AND U37450 ( .A(\modmult_1/xin[1023] ), .B(n36225), .Z(n36224) );
  IV U37451 ( .A(n36223), .Z(n36225) );
  XOR U37452 ( .A(n36226), .B(g_input[414]), .Z(n36223) );
  NAND U37453 ( .A(n36227), .B(mul_pow), .Z(n36226) );
  XOR U37454 ( .A(g_input[414]), .B(creg[414]), .Z(n36227) );
  XOR U37455 ( .A(n36228), .B(n36229), .Z(n36219) );
  ANDN U37456 ( .A(n36230), .B(n28262), .Z(n36229) );
  XOR U37457 ( .A(n36231), .B(\modmult_1/zin[0][412] ), .Z(n28262) );
  IV U37458 ( .A(n36228), .Z(n36231) );
  XNOR U37459 ( .A(n36228), .B(n28261), .Z(n36230) );
  XOR U37460 ( .A(n36232), .B(n36233), .Z(n28261) );
  AND U37461 ( .A(\modmult_1/xin[1023] ), .B(n36234), .Z(n36233) );
  IV U37462 ( .A(n36232), .Z(n36234) );
  XOR U37463 ( .A(n36235), .B(g_input[413]), .Z(n36232) );
  NAND U37464 ( .A(n36236), .B(mul_pow), .Z(n36235) );
  XOR U37465 ( .A(g_input[413]), .B(creg[413]), .Z(n36236) );
  XOR U37466 ( .A(n36237), .B(n36238), .Z(n36228) );
  ANDN U37467 ( .A(n36239), .B(n28268), .Z(n36238) );
  XOR U37468 ( .A(n36240), .B(\modmult_1/zin[0][411] ), .Z(n28268) );
  IV U37469 ( .A(n36237), .Z(n36240) );
  XNOR U37470 ( .A(n36237), .B(n28267), .Z(n36239) );
  XOR U37471 ( .A(n36241), .B(n36242), .Z(n28267) );
  AND U37472 ( .A(\modmult_1/xin[1023] ), .B(n36243), .Z(n36242) );
  IV U37473 ( .A(n36241), .Z(n36243) );
  XOR U37474 ( .A(n36244), .B(g_input[412]), .Z(n36241) );
  NAND U37475 ( .A(n36245), .B(mul_pow), .Z(n36244) );
  XOR U37476 ( .A(g_input[412]), .B(creg[412]), .Z(n36245) );
  XOR U37477 ( .A(n36246), .B(n36247), .Z(n36237) );
  ANDN U37478 ( .A(n36248), .B(n28274), .Z(n36247) );
  XOR U37479 ( .A(n36249), .B(\modmult_1/zin[0][410] ), .Z(n28274) );
  IV U37480 ( .A(n36246), .Z(n36249) );
  XNOR U37481 ( .A(n36246), .B(n28273), .Z(n36248) );
  XOR U37482 ( .A(n36250), .B(n36251), .Z(n28273) );
  AND U37483 ( .A(\modmult_1/xin[1023] ), .B(n36252), .Z(n36251) );
  IV U37484 ( .A(n36250), .Z(n36252) );
  XOR U37485 ( .A(n36253), .B(g_input[411]), .Z(n36250) );
  NAND U37486 ( .A(n36254), .B(mul_pow), .Z(n36253) );
  XOR U37487 ( .A(g_input[411]), .B(creg[411]), .Z(n36254) );
  XOR U37488 ( .A(n36255), .B(n36256), .Z(n36246) );
  ANDN U37489 ( .A(n36257), .B(n28280), .Z(n36256) );
  XOR U37490 ( .A(n36258), .B(\modmult_1/zin[0][409] ), .Z(n28280) );
  IV U37491 ( .A(n36255), .Z(n36258) );
  XNOR U37492 ( .A(n36255), .B(n28279), .Z(n36257) );
  XOR U37493 ( .A(n36259), .B(n36260), .Z(n28279) );
  AND U37494 ( .A(\modmult_1/xin[1023] ), .B(n36261), .Z(n36260) );
  IV U37495 ( .A(n36259), .Z(n36261) );
  XOR U37496 ( .A(n36262), .B(g_input[410]), .Z(n36259) );
  NAND U37497 ( .A(n36263), .B(mul_pow), .Z(n36262) );
  XOR U37498 ( .A(g_input[410]), .B(creg[410]), .Z(n36263) );
  XOR U37499 ( .A(n36264), .B(n36265), .Z(n36255) );
  ANDN U37500 ( .A(n36266), .B(n28286), .Z(n36265) );
  XOR U37501 ( .A(n36267), .B(\modmult_1/zin[0][408] ), .Z(n28286) );
  IV U37502 ( .A(n36264), .Z(n36267) );
  XNOR U37503 ( .A(n36264), .B(n28285), .Z(n36266) );
  XOR U37504 ( .A(n36268), .B(n36269), .Z(n28285) );
  AND U37505 ( .A(\modmult_1/xin[1023] ), .B(n36270), .Z(n36269) );
  IV U37506 ( .A(n36268), .Z(n36270) );
  XOR U37507 ( .A(n36271), .B(g_input[409]), .Z(n36268) );
  NAND U37508 ( .A(n36272), .B(mul_pow), .Z(n36271) );
  XOR U37509 ( .A(g_input[409]), .B(creg[409]), .Z(n36272) );
  XOR U37510 ( .A(n36273), .B(n36274), .Z(n36264) );
  ANDN U37511 ( .A(n36275), .B(n28292), .Z(n36274) );
  XOR U37512 ( .A(n36276), .B(\modmult_1/zin[0][407] ), .Z(n28292) );
  IV U37513 ( .A(n36273), .Z(n36276) );
  XNOR U37514 ( .A(n36273), .B(n28291), .Z(n36275) );
  XOR U37515 ( .A(n36277), .B(n36278), .Z(n28291) );
  AND U37516 ( .A(\modmult_1/xin[1023] ), .B(n36279), .Z(n36278) );
  IV U37517 ( .A(n36277), .Z(n36279) );
  XOR U37518 ( .A(n36280), .B(g_input[408]), .Z(n36277) );
  NAND U37519 ( .A(n36281), .B(mul_pow), .Z(n36280) );
  XOR U37520 ( .A(g_input[408]), .B(creg[408]), .Z(n36281) );
  XOR U37521 ( .A(n36282), .B(n36283), .Z(n36273) );
  ANDN U37522 ( .A(n36284), .B(n28298), .Z(n36283) );
  XOR U37523 ( .A(n36285), .B(\modmult_1/zin[0][406] ), .Z(n28298) );
  IV U37524 ( .A(n36282), .Z(n36285) );
  XNOR U37525 ( .A(n36282), .B(n28297), .Z(n36284) );
  XOR U37526 ( .A(n36286), .B(n36287), .Z(n28297) );
  AND U37527 ( .A(\modmult_1/xin[1023] ), .B(n36288), .Z(n36287) );
  IV U37528 ( .A(n36286), .Z(n36288) );
  XOR U37529 ( .A(n36289), .B(g_input[407]), .Z(n36286) );
  NAND U37530 ( .A(n36290), .B(mul_pow), .Z(n36289) );
  XOR U37531 ( .A(g_input[407]), .B(creg[407]), .Z(n36290) );
  XOR U37532 ( .A(n36291), .B(n36292), .Z(n36282) );
  ANDN U37533 ( .A(n36293), .B(n28304), .Z(n36292) );
  XOR U37534 ( .A(n36294), .B(\modmult_1/zin[0][405] ), .Z(n28304) );
  IV U37535 ( .A(n36291), .Z(n36294) );
  XNOR U37536 ( .A(n36291), .B(n28303), .Z(n36293) );
  XOR U37537 ( .A(n36295), .B(n36296), .Z(n28303) );
  AND U37538 ( .A(\modmult_1/xin[1023] ), .B(n36297), .Z(n36296) );
  IV U37539 ( .A(n36295), .Z(n36297) );
  XOR U37540 ( .A(n36298), .B(g_input[406]), .Z(n36295) );
  NAND U37541 ( .A(n36299), .B(mul_pow), .Z(n36298) );
  XOR U37542 ( .A(g_input[406]), .B(creg[406]), .Z(n36299) );
  XOR U37543 ( .A(n36300), .B(n36301), .Z(n36291) );
  ANDN U37544 ( .A(n36302), .B(n28310), .Z(n36301) );
  XOR U37545 ( .A(n36303), .B(\modmult_1/zin[0][404] ), .Z(n28310) );
  IV U37546 ( .A(n36300), .Z(n36303) );
  XNOR U37547 ( .A(n36300), .B(n28309), .Z(n36302) );
  XOR U37548 ( .A(n36304), .B(n36305), .Z(n28309) );
  AND U37549 ( .A(\modmult_1/xin[1023] ), .B(n36306), .Z(n36305) );
  IV U37550 ( .A(n36304), .Z(n36306) );
  XOR U37551 ( .A(n36307), .B(g_input[405]), .Z(n36304) );
  NAND U37552 ( .A(n36308), .B(mul_pow), .Z(n36307) );
  XOR U37553 ( .A(g_input[405]), .B(creg[405]), .Z(n36308) );
  XOR U37554 ( .A(n36309), .B(n36310), .Z(n36300) );
  ANDN U37555 ( .A(n36311), .B(n28316), .Z(n36310) );
  XOR U37556 ( .A(n36312), .B(\modmult_1/zin[0][403] ), .Z(n28316) );
  IV U37557 ( .A(n36309), .Z(n36312) );
  XNOR U37558 ( .A(n36309), .B(n28315), .Z(n36311) );
  XOR U37559 ( .A(n36313), .B(n36314), .Z(n28315) );
  AND U37560 ( .A(\modmult_1/xin[1023] ), .B(n36315), .Z(n36314) );
  IV U37561 ( .A(n36313), .Z(n36315) );
  XOR U37562 ( .A(n36316), .B(g_input[404]), .Z(n36313) );
  NAND U37563 ( .A(n36317), .B(mul_pow), .Z(n36316) );
  XOR U37564 ( .A(g_input[404]), .B(creg[404]), .Z(n36317) );
  XOR U37565 ( .A(n36318), .B(n36319), .Z(n36309) );
  ANDN U37566 ( .A(n36320), .B(n28322), .Z(n36319) );
  XOR U37567 ( .A(n36321), .B(\modmult_1/zin[0][402] ), .Z(n28322) );
  IV U37568 ( .A(n36318), .Z(n36321) );
  XNOR U37569 ( .A(n36318), .B(n28321), .Z(n36320) );
  XOR U37570 ( .A(n36322), .B(n36323), .Z(n28321) );
  AND U37571 ( .A(\modmult_1/xin[1023] ), .B(n36324), .Z(n36323) );
  IV U37572 ( .A(n36322), .Z(n36324) );
  XOR U37573 ( .A(n36325), .B(g_input[403]), .Z(n36322) );
  NAND U37574 ( .A(n36326), .B(mul_pow), .Z(n36325) );
  XOR U37575 ( .A(g_input[403]), .B(creg[403]), .Z(n36326) );
  XOR U37576 ( .A(n36327), .B(n36328), .Z(n36318) );
  ANDN U37577 ( .A(n36329), .B(n28328), .Z(n36328) );
  XOR U37578 ( .A(n36330), .B(\modmult_1/zin[0][401] ), .Z(n28328) );
  IV U37579 ( .A(n36327), .Z(n36330) );
  XNOR U37580 ( .A(n36327), .B(n28327), .Z(n36329) );
  XOR U37581 ( .A(n36331), .B(n36332), .Z(n28327) );
  AND U37582 ( .A(\modmult_1/xin[1023] ), .B(n36333), .Z(n36332) );
  IV U37583 ( .A(n36331), .Z(n36333) );
  XOR U37584 ( .A(n36334), .B(g_input[402]), .Z(n36331) );
  NAND U37585 ( .A(n36335), .B(mul_pow), .Z(n36334) );
  XOR U37586 ( .A(g_input[402]), .B(creg[402]), .Z(n36335) );
  XOR U37587 ( .A(n36336), .B(n36337), .Z(n36327) );
  ANDN U37588 ( .A(n36338), .B(n28334), .Z(n36337) );
  XOR U37589 ( .A(n36339), .B(\modmult_1/zin[0][400] ), .Z(n28334) );
  IV U37590 ( .A(n36336), .Z(n36339) );
  XNOR U37591 ( .A(n36336), .B(n28333), .Z(n36338) );
  XOR U37592 ( .A(n36340), .B(n36341), .Z(n28333) );
  AND U37593 ( .A(\modmult_1/xin[1023] ), .B(n36342), .Z(n36341) );
  IV U37594 ( .A(n36340), .Z(n36342) );
  XOR U37595 ( .A(n36343), .B(g_input[401]), .Z(n36340) );
  NAND U37596 ( .A(n36344), .B(mul_pow), .Z(n36343) );
  XOR U37597 ( .A(g_input[401]), .B(creg[401]), .Z(n36344) );
  XOR U37598 ( .A(n36345), .B(n36346), .Z(n36336) );
  ANDN U37599 ( .A(n36347), .B(n28340), .Z(n36346) );
  XOR U37600 ( .A(n36348), .B(\modmult_1/zin[0][399] ), .Z(n28340) );
  IV U37601 ( .A(n36345), .Z(n36348) );
  XNOR U37602 ( .A(n36345), .B(n28339), .Z(n36347) );
  XOR U37603 ( .A(n36349), .B(n36350), .Z(n28339) );
  AND U37604 ( .A(\modmult_1/xin[1023] ), .B(n36351), .Z(n36350) );
  IV U37605 ( .A(n36349), .Z(n36351) );
  XOR U37606 ( .A(n36352), .B(g_input[400]), .Z(n36349) );
  NAND U37607 ( .A(n36353), .B(mul_pow), .Z(n36352) );
  XOR U37608 ( .A(g_input[400]), .B(creg[400]), .Z(n36353) );
  XOR U37609 ( .A(n36354), .B(n36355), .Z(n36345) );
  ANDN U37610 ( .A(n36356), .B(n28346), .Z(n36355) );
  XOR U37611 ( .A(n36357), .B(\modmult_1/zin[0][398] ), .Z(n28346) );
  IV U37612 ( .A(n36354), .Z(n36357) );
  XNOR U37613 ( .A(n36354), .B(n28345), .Z(n36356) );
  XOR U37614 ( .A(n36358), .B(n36359), .Z(n28345) );
  AND U37615 ( .A(\modmult_1/xin[1023] ), .B(n36360), .Z(n36359) );
  IV U37616 ( .A(n36358), .Z(n36360) );
  XOR U37617 ( .A(n36361), .B(g_input[399]), .Z(n36358) );
  NAND U37618 ( .A(n36362), .B(mul_pow), .Z(n36361) );
  XOR U37619 ( .A(g_input[399]), .B(creg[399]), .Z(n36362) );
  XOR U37620 ( .A(n36363), .B(n36364), .Z(n36354) );
  ANDN U37621 ( .A(n36365), .B(n28352), .Z(n36364) );
  XOR U37622 ( .A(n36366), .B(\modmult_1/zin[0][397] ), .Z(n28352) );
  IV U37623 ( .A(n36363), .Z(n36366) );
  XNOR U37624 ( .A(n36363), .B(n28351), .Z(n36365) );
  XOR U37625 ( .A(n36367), .B(n36368), .Z(n28351) );
  AND U37626 ( .A(\modmult_1/xin[1023] ), .B(n36369), .Z(n36368) );
  IV U37627 ( .A(n36367), .Z(n36369) );
  XOR U37628 ( .A(n36370), .B(g_input[398]), .Z(n36367) );
  NAND U37629 ( .A(n36371), .B(mul_pow), .Z(n36370) );
  XOR U37630 ( .A(g_input[398]), .B(creg[398]), .Z(n36371) );
  XOR U37631 ( .A(n36372), .B(n36373), .Z(n36363) );
  ANDN U37632 ( .A(n36374), .B(n28358), .Z(n36373) );
  XOR U37633 ( .A(n36375), .B(\modmult_1/zin[0][396] ), .Z(n28358) );
  IV U37634 ( .A(n36372), .Z(n36375) );
  XNOR U37635 ( .A(n36372), .B(n28357), .Z(n36374) );
  XOR U37636 ( .A(n36376), .B(n36377), .Z(n28357) );
  AND U37637 ( .A(\modmult_1/xin[1023] ), .B(n36378), .Z(n36377) );
  IV U37638 ( .A(n36376), .Z(n36378) );
  XOR U37639 ( .A(n36379), .B(g_input[397]), .Z(n36376) );
  NAND U37640 ( .A(n36380), .B(mul_pow), .Z(n36379) );
  XOR U37641 ( .A(g_input[397]), .B(creg[397]), .Z(n36380) );
  XOR U37642 ( .A(n36381), .B(n36382), .Z(n36372) );
  ANDN U37643 ( .A(n36383), .B(n28364), .Z(n36382) );
  XOR U37644 ( .A(n36384), .B(\modmult_1/zin[0][395] ), .Z(n28364) );
  IV U37645 ( .A(n36381), .Z(n36384) );
  XNOR U37646 ( .A(n36381), .B(n28363), .Z(n36383) );
  XOR U37647 ( .A(n36385), .B(n36386), .Z(n28363) );
  AND U37648 ( .A(\modmult_1/xin[1023] ), .B(n36387), .Z(n36386) );
  IV U37649 ( .A(n36385), .Z(n36387) );
  XOR U37650 ( .A(n36388), .B(g_input[396]), .Z(n36385) );
  NAND U37651 ( .A(n36389), .B(mul_pow), .Z(n36388) );
  XOR U37652 ( .A(g_input[396]), .B(creg[396]), .Z(n36389) );
  XOR U37653 ( .A(n36390), .B(n36391), .Z(n36381) );
  ANDN U37654 ( .A(n36392), .B(n28370), .Z(n36391) );
  XOR U37655 ( .A(n36393), .B(\modmult_1/zin[0][394] ), .Z(n28370) );
  IV U37656 ( .A(n36390), .Z(n36393) );
  XNOR U37657 ( .A(n36390), .B(n28369), .Z(n36392) );
  XOR U37658 ( .A(n36394), .B(n36395), .Z(n28369) );
  AND U37659 ( .A(\modmult_1/xin[1023] ), .B(n36396), .Z(n36395) );
  IV U37660 ( .A(n36394), .Z(n36396) );
  XOR U37661 ( .A(n36397), .B(g_input[395]), .Z(n36394) );
  NAND U37662 ( .A(n36398), .B(mul_pow), .Z(n36397) );
  XOR U37663 ( .A(g_input[395]), .B(creg[395]), .Z(n36398) );
  XOR U37664 ( .A(n36399), .B(n36400), .Z(n36390) );
  ANDN U37665 ( .A(n36401), .B(n28376), .Z(n36400) );
  XOR U37666 ( .A(n36402), .B(\modmult_1/zin[0][393] ), .Z(n28376) );
  IV U37667 ( .A(n36399), .Z(n36402) );
  XNOR U37668 ( .A(n36399), .B(n28375), .Z(n36401) );
  XOR U37669 ( .A(n36403), .B(n36404), .Z(n28375) );
  AND U37670 ( .A(\modmult_1/xin[1023] ), .B(n36405), .Z(n36404) );
  IV U37671 ( .A(n36403), .Z(n36405) );
  XOR U37672 ( .A(n36406), .B(g_input[394]), .Z(n36403) );
  NAND U37673 ( .A(n36407), .B(mul_pow), .Z(n36406) );
  XOR U37674 ( .A(g_input[394]), .B(creg[394]), .Z(n36407) );
  XOR U37675 ( .A(n36408), .B(n36409), .Z(n36399) );
  ANDN U37676 ( .A(n36410), .B(n28382), .Z(n36409) );
  XOR U37677 ( .A(n36411), .B(\modmult_1/zin[0][392] ), .Z(n28382) );
  IV U37678 ( .A(n36408), .Z(n36411) );
  XNOR U37679 ( .A(n36408), .B(n28381), .Z(n36410) );
  XOR U37680 ( .A(n36412), .B(n36413), .Z(n28381) );
  AND U37681 ( .A(\modmult_1/xin[1023] ), .B(n36414), .Z(n36413) );
  IV U37682 ( .A(n36412), .Z(n36414) );
  XOR U37683 ( .A(n36415), .B(g_input[393]), .Z(n36412) );
  NAND U37684 ( .A(n36416), .B(mul_pow), .Z(n36415) );
  XOR U37685 ( .A(g_input[393]), .B(creg[393]), .Z(n36416) );
  XOR U37686 ( .A(n36417), .B(n36418), .Z(n36408) );
  ANDN U37687 ( .A(n36419), .B(n28388), .Z(n36418) );
  XOR U37688 ( .A(n36420), .B(\modmult_1/zin[0][391] ), .Z(n28388) );
  IV U37689 ( .A(n36417), .Z(n36420) );
  XNOR U37690 ( .A(n36417), .B(n28387), .Z(n36419) );
  XOR U37691 ( .A(n36421), .B(n36422), .Z(n28387) );
  AND U37692 ( .A(\modmult_1/xin[1023] ), .B(n36423), .Z(n36422) );
  IV U37693 ( .A(n36421), .Z(n36423) );
  XOR U37694 ( .A(n36424), .B(g_input[392]), .Z(n36421) );
  NAND U37695 ( .A(n36425), .B(mul_pow), .Z(n36424) );
  XOR U37696 ( .A(g_input[392]), .B(creg[392]), .Z(n36425) );
  XOR U37697 ( .A(n36426), .B(n36427), .Z(n36417) );
  ANDN U37698 ( .A(n36428), .B(n28394), .Z(n36427) );
  XOR U37699 ( .A(n36429), .B(\modmult_1/zin[0][390] ), .Z(n28394) );
  IV U37700 ( .A(n36426), .Z(n36429) );
  XNOR U37701 ( .A(n36426), .B(n28393), .Z(n36428) );
  XOR U37702 ( .A(n36430), .B(n36431), .Z(n28393) );
  AND U37703 ( .A(\modmult_1/xin[1023] ), .B(n36432), .Z(n36431) );
  IV U37704 ( .A(n36430), .Z(n36432) );
  XOR U37705 ( .A(n36433), .B(g_input[391]), .Z(n36430) );
  NAND U37706 ( .A(n36434), .B(mul_pow), .Z(n36433) );
  XOR U37707 ( .A(g_input[391]), .B(creg[391]), .Z(n36434) );
  XOR U37708 ( .A(n36435), .B(n36436), .Z(n36426) );
  ANDN U37709 ( .A(n36437), .B(n28400), .Z(n36436) );
  XOR U37710 ( .A(n36438), .B(\modmult_1/zin[0][389] ), .Z(n28400) );
  IV U37711 ( .A(n36435), .Z(n36438) );
  XNOR U37712 ( .A(n36435), .B(n28399), .Z(n36437) );
  XOR U37713 ( .A(n36439), .B(n36440), .Z(n28399) );
  AND U37714 ( .A(\modmult_1/xin[1023] ), .B(n36441), .Z(n36440) );
  IV U37715 ( .A(n36439), .Z(n36441) );
  XOR U37716 ( .A(n36442), .B(g_input[390]), .Z(n36439) );
  NAND U37717 ( .A(n36443), .B(mul_pow), .Z(n36442) );
  XOR U37718 ( .A(g_input[390]), .B(creg[390]), .Z(n36443) );
  XOR U37719 ( .A(n36444), .B(n36445), .Z(n36435) );
  ANDN U37720 ( .A(n36446), .B(n28406), .Z(n36445) );
  XOR U37721 ( .A(n36447), .B(\modmult_1/zin[0][388] ), .Z(n28406) );
  IV U37722 ( .A(n36444), .Z(n36447) );
  XNOR U37723 ( .A(n36444), .B(n28405), .Z(n36446) );
  XOR U37724 ( .A(n36448), .B(n36449), .Z(n28405) );
  AND U37725 ( .A(\modmult_1/xin[1023] ), .B(n36450), .Z(n36449) );
  IV U37726 ( .A(n36448), .Z(n36450) );
  XOR U37727 ( .A(n36451), .B(g_input[389]), .Z(n36448) );
  NAND U37728 ( .A(n36452), .B(mul_pow), .Z(n36451) );
  XOR U37729 ( .A(g_input[389]), .B(creg[389]), .Z(n36452) );
  XOR U37730 ( .A(n36453), .B(n36454), .Z(n36444) );
  ANDN U37731 ( .A(n36455), .B(n28412), .Z(n36454) );
  XOR U37732 ( .A(n36456), .B(\modmult_1/zin[0][387] ), .Z(n28412) );
  IV U37733 ( .A(n36453), .Z(n36456) );
  XNOR U37734 ( .A(n36453), .B(n28411), .Z(n36455) );
  XOR U37735 ( .A(n36457), .B(n36458), .Z(n28411) );
  AND U37736 ( .A(\modmult_1/xin[1023] ), .B(n36459), .Z(n36458) );
  IV U37737 ( .A(n36457), .Z(n36459) );
  XOR U37738 ( .A(n36460), .B(g_input[388]), .Z(n36457) );
  NAND U37739 ( .A(n36461), .B(mul_pow), .Z(n36460) );
  XOR U37740 ( .A(g_input[388]), .B(creg[388]), .Z(n36461) );
  XOR U37741 ( .A(n36462), .B(n36463), .Z(n36453) );
  ANDN U37742 ( .A(n36464), .B(n28418), .Z(n36463) );
  XOR U37743 ( .A(n36465), .B(\modmult_1/zin[0][386] ), .Z(n28418) );
  IV U37744 ( .A(n36462), .Z(n36465) );
  XNOR U37745 ( .A(n36462), .B(n28417), .Z(n36464) );
  XOR U37746 ( .A(n36466), .B(n36467), .Z(n28417) );
  AND U37747 ( .A(\modmult_1/xin[1023] ), .B(n36468), .Z(n36467) );
  IV U37748 ( .A(n36466), .Z(n36468) );
  XOR U37749 ( .A(n36469), .B(g_input[387]), .Z(n36466) );
  NAND U37750 ( .A(n36470), .B(mul_pow), .Z(n36469) );
  XOR U37751 ( .A(g_input[387]), .B(creg[387]), .Z(n36470) );
  XOR U37752 ( .A(n36471), .B(n36472), .Z(n36462) );
  ANDN U37753 ( .A(n36473), .B(n28424), .Z(n36472) );
  XOR U37754 ( .A(n36474), .B(\modmult_1/zin[0][385] ), .Z(n28424) );
  IV U37755 ( .A(n36471), .Z(n36474) );
  XNOR U37756 ( .A(n36471), .B(n28423), .Z(n36473) );
  XOR U37757 ( .A(n36475), .B(n36476), .Z(n28423) );
  AND U37758 ( .A(\modmult_1/xin[1023] ), .B(n36477), .Z(n36476) );
  IV U37759 ( .A(n36475), .Z(n36477) );
  XOR U37760 ( .A(n36478), .B(g_input[386]), .Z(n36475) );
  NAND U37761 ( .A(n36479), .B(mul_pow), .Z(n36478) );
  XOR U37762 ( .A(g_input[386]), .B(creg[386]), .Z(n36479) );
  XOR U37763 ( .A(n36480), .B(n36481), .Z(n36471) );
  ANDN U37764 ( .A(n36482), .B(n28430), .Z(n36481) );
  XOR U37765 ( .A(n36483), .B(\modmult_1/zin[0][384] ), .Z(n28430) );
  IV U37766 ( .A(n36480), .Z(n36483) );
  XNOR U37767 ( .A(n36480), .B(n28429), .Z(n36482) );
  XOR U37768 ( .A(n36484), .B(n36485), .Z(n28429) );
  AND U37769 ( .A(\modmult_1/xin[1023] ), .B(n36486), .Z(n36485) );
  IV U37770 ( .A(n36484), .Z(n36486) );
  XOR U37771 ( .A(n36487), .B(g_input[385]), .Z(n36484) );
  NAND U37772 ( .A(n36488), .B(mul_pow), .Z(n36487) );
  XOR U37773 ( .A(g_input[385]), .B(creg[385]), .Z(n36488) );
  XOR U37774 ( .A(n36489), .B(n36490), .Z(n36480) );
  ANDN U37775 ( .A(n36491), .B(n28436), .Z(n36490) );
  XOR U37776 ( .A(n36492), .B(\modmult_1/zin[0][383] ), .Z(n28436) );
  IV U37777 ( .A(n36489), .Z(n36492) );
  XNOR U37778 ( .A(n36489), .B(n28435), .Z(n36491) );
  XOR U37779 ( .A(n36493), .B(n36494), .Z(n28435) );
  AND U37780 ( .A(\modmult_1/xin[1023] ), .B(n36495), .Z(n36494) );
  IV U37781 ( .A(n36493), .Z(n36495) );
  XOR U37782 ( .A(n36496), .B(g_input[384]), .Z(n36493) );
  NAND U37783 ( .A(n36497), .B(mul_pow), .Z(n36496) );
  XOR U37784 ( .A(g_input[384]), .B(creg[384]), .Z(n36497) );
  XOR U37785 ( .A(n36498), .B(n36499), .Z(n36489) );
  ANDN U37786 ( .A(n36500), .B(n28442), .Z(n36499) );
  XOR U37787 ( .A(n36501), .B(\modmult_1/zin[0][382] ), .Z(n28442) );
  IV U37788 ( .A(n36498), .Z(n36501) );
  XNOR U37789 ( .A(n36498), .B(n28441), .Z(n36500) );
  XOR U37790 ( .A(n36502), .B(n36503), .Z(n28441) );
  AND U37791 ( .A(\modmult_1/xin[1023] ), .B(n36504), .Z(n36503) );
  IV U37792 ( .A(n36502), .Z(n36504) );
  XOR U37793 ( .A(n36505), .B(g_input[383]), .Z(n36502) );
  NAND U37794 ( .A(n36506), .B(mul_pow), .Z(n36505) );
  XOR U37795 ( .A(g_input[383]), .B(creg[383]), .Z(n36506) );
  XOR U37796 ( .A(n36507), .B(n36508), .Z(n36498) );
  ANDN U37797 ( .A(n36509), .B(n28448), .Z(n36508) );
  XOR U37798 ( .A(n36510), .B(\modmult_1/zin[0][381] ), .Z(n28448) );
  IV U37799 ( .A(n36507), .Z(n36510) );
  XNOR U37800 ( .A(n36507), .B(n28447), .Z(n36509) );
  XOR U37801 ( .A(n36511), .B(n36512), .Z(n28447) );
  AND U37802 ( .A(\modmult_1/xin[1023] ), .B(n36513), .Z(n36512) );
  IV U37803 ( .A(n36511), .Z(n36513) );
  XOR U37804 ( .A(n36514), .B(g_input[382]), .Z(n36511) );
  NAND U37805 ( .A(n36515), .B(mul_pow), .Z(n36514) );
  XOR U37806 ( .A(g_input[382]), .B(creg[382]), .Z(n36515) );
  XOR U37807 ( .A(n36516), .B(n36517), .Z(n36507) );
  ANDN U37808 ( .A(n36518), .B(n28454), .Z(n36517) );
  XOR U37809 ( .A(n36519), .B(\modmult_1/zin[0][380] ), .Z(n28454) );
  IV U37810 ( .A(n36516), .Z(n36519) );
  XNOR U37811 ( .A(n36516), .B(n28453), .Z(n36518) );
  XOR U37812 ( .A(n36520), .B(n36521), .Z(n28453) );
  AND U37813 ( .A(\modmult_1/xin[1023] ), .B(n36522), .Z(n36521) );
  IV U37814 ( .A(n36520), .Z(n36522) );
  XOR U37815 ( .A(n36523), .B(g_input[381]), .Z(n36520) );
  NAND U37816 ( .A(n36524), .B(mul_pow), .Z(n36523) );
  XOR U37817 ( .A(g_input[381]), .B(creg[381]), .Z(n36524) );
  XOR U37818 ( .A(n36525), .B(n36526), .Z(n36516) );
  ANDN U37819 ( .A(n36527), .B(n28460), .Z(n36526) );
  XOR U37820 ( .A(n36528), .B(\modmult_1/zin[0][379] ), .Z(n28460) );
  IV U37821 ( .A(n36525), .Z(n36528) );
  XNOR U37822 ( .A(n36525), .B(n28459), .Z(n36527) );
  XOR U37823 ( .A(n36529), .B(n36530), .Z(n28459) );
  AND U37824 ( .A(\modmult_1/xin[1023] ), .B(n36531), .Z(n36530) );
  IV U37825 ( .A(n36529), .Z(n36531) );
  XOR U37826 ( .A(n36532), .B(g_input[380]), .Z(n36529) );
  NAND U37827 ( .A(n36533), .B(mul_pow), .Z(n36532) );
  XOR U37828 ( .A(g_input[380]), .B(creg[380]), .Z(n36533) );
  XOR U37829 ( .A(n36534), .B(n36535), .Z(n36525) );
  ANDN U37830 ( .A(n36536), .B(n28466), .Z(n36535) );
  XOR U37831 ( .A(n36537), .B(\modmult_1/zin[0][378] ), .Z(n28466) );
  IV U37832 ( .A(n36534), .Z(n36537) );
  XNOR U37833 ( .A(n36534), .B(n28465), .Z(n36536) );
  XOR U37834 ( .A(n36538), .B(n36539), .Z(n28465) );
  AND U37835 ( .A(\modmult_1/xin[1023] ), .B(n36540), .Z(n36539) );
  IV U37836 ( .A(n36538), .Z(n36540) );
  XOR U37837 ( .A(n36541), .B(g_input[379]), .Z(n36538) );
  NAND U37838 ( .A(n36542), .B(mul_pow), .Z(n36541) );
  XOR U37839 ( .A(g_input[379]), .B(creg[379]), .Z(n36542) );
  XOR U37840 ( .A(n36543), .B(n36544), .Z(n36534) );
  ANDN U37841 ( .A(n36545), .B(n28472), .Z(n36544) );
  XOR U37842 ( .A(n36546), .B(\modmult_1/zin[0][377] ), .Z(n28472) );
  IV U37843 ( .A(n36543), .Z(n36546) );
  XNOR U37844 ( .A(n36543), .B(n28471), .Z(n36545) );
  XOR U37845 ( .A(n36547), .B(n36548), .Z(n28471) );
  AND U37846 ( .A(\modmult_1/xin[1023] ), .B(n36549), .Z(n36548) );
  IV U37847 ( .A(n36547), .Z(n36549) );
  XOR U37848 ( .A(n36550), .B(g_input[378]), .Z(n36547) );
  NAND U37849 ( .A(n36551), .B(mul_pow), .Z(n36550) );
  XOR U37850 ( .A(g_input[378]), .B(creg[378]), .Z(n36551) );
  XOR U37851 ( .A(n36552), .B(n36553), .Z(n36543) );
  ANDN U37852 ( .A(n36554), .B(n28478), .Z(n36553) );
  XOR U37853 ( .A(n36555), .B(\modmult_1/zin[0][376] ), .Z(n28478) );
  IV U37854 ( .A(n36552), .Z(n36555) );
  XNOR U37855 ( .A(n36552), .B(n28477), .Z(n36554) );
  XOR U37856 ( .A(n36556), .B(n36557), .Z(n28477) );
  AND U37857 ( .A(\modmult_1/xin[1023] ), .B(n36558), .Z(n36557) );
  IV U37858 ( .A(n36556), .Z(n36558) );
  XOR U37859 ( .A(n36559), .B(g_input[377]), .Z(n36556) );
  NAND U37860 ( .A(n36560), .B(mul_pow), .Z(n36559) );
  XOR U37861 ( .A(g_input[377]), .B(creg[377]), .Z(n36560) );
  XOR U37862 ( .A(n36561), .B(n36562), .Z(n36552) );
  ANDN U37863 ( .A(n36563), .B(n28484), .Z(n36562) );
  XOR U37864 ( .A(n36564), .B(\modmult_1/zin[0][375] ), .Z(n28484) );
  IV U37865 ( .A(n36561), .Z(n36564) );
  XNOR U37866 ( .A(n36561), .B(n28483), .Z(n36563) );
  XOR U37867 ( .A(n36565), .B(n36566), .Z(n28483) );
  AND U37868 ( .A(\modmult_1/xin[1023] ), .B(n36567), .Z(n36566) );
  IV U37869 ( .A(n36565), .Z(n36567) );
  XOR U37870 ( .A(n36568), .B(g_input[376]), .Z(n36565) );
  NAND U37871 ( .A(n36569), .B(mul_pow), .Z(n36568) );
  XOR U37872 ( .A(g_input[376]), .B(creg[376]), .Z(n36569) );
  XOR U37873 ( .A(n36570), .B(n36571), .Z(n36561) );
  ANDN U37874 ( .A(n36572), .B(n28490), .Z(n36571) );
  XOR U37875 ( .A(n36573), .B(\modmult_1/zin[0][374] ), .Z(n28490) );
  IV U37876 ( .A(n36570), .Z(n36573) );
  XNOR U37877 ( .A(n36570), .B(n28489), .Z(n36572) );
  XOR U37878 ( .A(n36574), .B(n36575), .Z(n28489) );
  AND U37879 ( .A(\modmult_1/xin[1023] ), .B(n36576), .Z(n36575) );
  IV U37880 ( .A(n36574), .Z(n36576) );
  XOR U37881 ( .A(n36577), .B(g_input[375]), .Z(n36574) );
  NAND U37882 ( .A(n36578), .B(mul_pow), .Z(n36577) );
  XOR U37883 ( .A(g_input[375]), .B(creg[375]), .Z(n36578) );
  XOR U37884 ( .A(n36579), .B(n36580), .Z(n36570) );
  ANDN U37885 ( .A(n36581), .B(n28496), .Z(n36580) );
  XOR U37886 ( .A(n36582), .B(\modmult_1/zin[0][373] ), .Z(n28496) );
  IV U37887 ( .A(n36579), .Z(n36582) );
  XNOR U37888 ( .A(n36579), .B(n28495), .Z(n36581) );
  XOR U37889 ( .A(n36583), .B(n36584), .Z(n28495) );
  AND U37890 ( .A(\modmult_1/xin[1023] ), .B(n36585), .Z(n36584) );
  IV U37891 ( .A(n36583), .Z(n36585) );
  XOR U37892 ( .A(n36586), .B(g_input[374]), .Z(n36583) );
  NAND U37893 ( .A(n36587), .B(mul_pow), .Z(n36586) );
  XOR U37894 ( .A(g_input[374]), .B(creg[374]), .Z(n36587) );
  XOR U37895 ( .A(n36588), .B(n36589), .Z(n36579) );
  ANDN U37896 ( .A(n36590), .B(n28502), .Z(n36589) );
  XOR U37897 ( .A(n36591), .B(\modmult_1/zin[0][372] ), .Z(n28502) );
  IV U37898 ( .A(n36588), .Z(n36591) );
  XNOR U37899 ( .A(n36588), .B(n28501), .Z(n36590) );
  XOR U37900 ( .A(n36592), .B(n36593), .Z(n28501) );
  AND U37901 ( .A(\modmult_1/xin[1023] ), .B(n36594), .Z(n36593) );
  IV U37902 ( .A(n36592), .Z(n36594) );
  XOR U37903 ( .A(n36595), .B(g_input[373]), .Z(n36592) );
  NAND U37904 ( .A(n36596), .B(mul_pow), .Z(n36595) );
  XOR U37905 ( .A(g_input[373]), .B(creg[373]), .Z(n36596) );
  XOR U37906 ( .A(n36597), .B(n36598), .Z(n36588) );
  ANDN U37907 ( .A(n36599), .B(n28508), .Z(n36598) );
  XOR U37908 ( .A(n36600), .B(\modmult_1/zin[0][371] ), .Z(n28508) );
  IV U37909 ( .A(n36597), .Z(n36600) );
  XNOR U37910 ( .A(n36597), .B(n28507), .Z(n36599) );
  XOR U37911 ( .A(n36601), .B(n36602), .Z(n28507) );
  AND U37912 ( .A(\modmult_1/xin[1023] ), .B(n36603), .Z(n36602) );
  IV U37913 ( .A(n36601), .Z(n36603) );
  XOR U37914 ( .A(n36604), .B(g_input[372]), .Z(n36601) );
  NAND U37915 ( .A(n36605), .B(mul_pow), .Z(n36604) );
  XOR U37916 ( .A(g_input[372]), .B(creg[372]), .Z(n36605) );
  XOR U37917 ( .A(n36606), .B(n36607), .Z(n36597) );
  ANDN U37918 ( .A(n36608), .B(n28514), .Z(n36607) );
  XOR U37919 ( .A(n36609), .B(\modmult_1/zin[0][370] ), .Z(n28514) );
  IV U37920 ( .A(n36606), .Z(n36609) );
  XNOR U37921 ( .A(n36606), .B(n28513), .Z(n36608) );
  XOR U37922 ( .A(n36610), .B(n36611), .Z(n28513) );
  AND U37923 ( .A(\modmult_1/xin[1023] ), .B(n36612), .Z(n36611) );
  IV U37924 ( .A(n36610), .Z(n36612) );
  XOR U37925 ( .A(n36613), .B(g_input[371]), .Z(n36610) );
  NAND U37926 ( .A(n36614), .B(mul_pow), .Z(n36613) );
  XOR U37927 ( .A(g_input[371]), .B(creg[371]), .Z(n36614) );
  XOR U37928 ( .A(n36615), .B(n36616), .Z(n36606) );
  ANDN U37929 ( .A(n36617), .B(n28520), .Z(n36616) );
  XOR U37930 ( .A(n36618), .B(\modmult_1/zin[0][369] ), .Z(n28520) );
  IV U37931 ( .A(n36615), .Z(n36618) );
  XNOR U37932 ( .A(n36615), .B(n28519), .Z(n36617) );
  XOR U37933 ( .A(n36619), .B(n36620), .Z(n28519) );
  AND U37934 ( .A(\modmult_1/xin[1023] ), .B(n36621), .Z(n36620) );
  IV U37935 ( .A(n36619), .Z(n36621) );
  XOR U37936 ( .A(n36622), .B(g_input[370]), .Z(n36619) );
  NAND U37937 ( .A(n36623), .B(mul_pow), .Z(n36622) );
  XOR U37938 ( .A(g_input[370]), .B(creg[370]), .Z(n36623) );
  XOR U37939 ( .A(n36624), .B(n36625), .Z(n36615) );
  ANDN U37940 ( .A(n36626), .B(n28526), .Z(n36625) );
  XOR U37941 ( .A(n36627), .B(\modmult_1/zin[0][368] ), .Z(n28526) );
  IV U37942 ( .A(n36624), .Z(n36627) );
  XNOR U37943 ( .A(n36624), .B(n28525), .Z(n36626) );
  XOR U37944 ( .A(n36628), .B(n36629), .Z(n28525) );
  AND U37945 ( .A(\modmult_1/xin[1023] ), .B(n36630), .Z(n36629) );
  IV U37946 ( .A(n36628), .Z(n36630) );
  XOR U37947 ( .A(n36631), .B(g_input[369]), .Z(n36628) );
  NAND U37948 ( .A(n36632), .B(mul_pow), .Z(n36631) );
  XOR U37949 ( .A(g_input[369]), .B(creg[369]), .Z(n36632) );
  XOR U37950 ( .A(n36633), .B(n36634), .Z(n36624) );
  ANDN U37951 ( .A(n36635), .B(n28532), .Z(n36634) );
  XOR U37952 ( .A(n36636), .B(\modmult_1/zin[0][367] ), .Z(n28532) );
  IV U37953 ( .A(n36633), .Z(n36636) );
  XNOR U37954 ( .A(n36633), .B(n28531), .Z(n36635) );
  XOR U37955 ( .A(n36637), .B(n36638), .Z(n28531) );
  AND U37956 ( .A(\modmult_1/xin[1023] ), .B(n36639), .Z(n36638) );
  IV U37957 ( .A(n36637), .Z(n36639) );
  XOR U37958 ( .A(n36640), .B(g_input[368]), .Z(n36637) );
  NAND U37959 ( .A(n36641), .B(mul_pow), .Z(n36640) );
  XOR U37960 ( .A(g_input[368]), .B(creg[368]), .Z(n36641) );
  XOR U37961 ( .A(n36642), .B(n36643), .Z(n36633) );
  ANDN U37962 ( .A(n36644), .B(n28538), .Z(n36643) );
  XOR U37963 ( .A(n36645), .B(\modmult_1/zin[0][366] ), .Z(n28538) );
  IV U37964 ( .A(n36642), .Z(n36645) );
  XNOR U37965 ( .A(n36642), .B(n28537), .Z(n36644) );
  XOR U37966 ( .A(n36646), .B(n36647), .Z(n28537) );
  AND U37967 ( .A(\modmult_1/xin[1023] ), .B(n36648), .Z(n36647) );
  IV U37968 ( .A(n36646), .Z(n36648) );
  XOR U37969 ( .A(n36649), .B(g_input[367]), .Z(n36646) );
  NAND U37970 ( .A(n36650), .B(mul_pow), .Z(n36649) );
  XOR U37971 ( .A(g_input[367]), .B(creg[367]), .Z(n36650) );
  XOR U37972 ( .A(n36651), .B(n36652), .Z(n36642) );
  ANDN U37973 ( .A(n36653), .B(n28544), .Z(n36652) );
  XOR U37974 ( .A(n36654), .B(\modmult_1/zin[0][365] ), .Z(n28544) );
  IV U37975 ( .A(n36651), .Z(n36654) );
  XNOR U37976 ( .A(n36651), .B(n28543), .Z(n36653) );
  XOR U37977 ( .A(n36655), .B(n36656), .Z(n28543) );
  AND U37978 ( .A(\modmult_1/xin[1023] ), .B(n36657), .Z(n36656) );
  IV U37979 ( .A(n36655), .Z(n36657) );
  XOR U37980 ( .A(n36658), .B(g_input[366]), .Z(n36655) );
  NAND U37981 ( .A(n36659), .B(mul_pow), .Z(n36658) );
  XOR U37982 ( .A(g_input[366]), .B(creg[366]), .Z(n36659) );
  XOR U37983 ( .A(n36660), .B(n36661), .Z(n36651) );
  ANDN U37984 ( .A(n36662), .B(n28550), .Z(n36661) );
  XOR U37985 ( .A(n36663), .B(\modmult_1/zin[0][364] ), .Z(n28550) );
  IV U37986 ( .A(n36660), .Z(n36663) );
  XNOR U37987 ( .A(n36660), .B(n28549), .Z(n36662) );
  XOR U37988 ( .A(n36664), .B(n36665), .Z(n28549) );
  AND U37989 ( .A(\modmult_1/xin[1023] ), .B(n36666), .Z(n36665) );
  IV U37990 ( .A(n36664), .Z(n36666) );
  XOR U37991 ( .A(n36667), .B(g_input[365]), .Z(n36664) );
  NAND U37992 ( .A(n36668), .B(mul_pow), .Z(n36667) );
  XOR U37993 ( .A(g_input[365]), .B(creg[365]), .Z(n36668) );
  XOR U37994 ( .A(n36669), .B(n36670), .Z(n36660) );
  ANDN U37995 ( .A(n36671), .B(n28556), .Z(n36670) );
  XOR U37996 ( .A(n36672), .B(\modmult_1/zin[0][363] ), .Z(n28556) );
  IV U37997 ( .A(n36669), .Z(n36672) );
  XNOR U37998 ( .A(n36669), .B(n28555), .Z(n36671) );
  XOR U37999 ( .A(n36673), .B(n36674), .Z(n28555) );
  AND U38000 ( .A(\modmult_1/xin[1023] ), .B(n36675), .Z(n36674) );
  IV U38001 ( .A(n36673), .Z(n36675) );
  XOR U38002 ( .A(n36676), .B(g_input[364]), .Z(n36673) );
  NAND U38003 ( .A(n36677), .B(mul_pow), .Z(n36676) );
  XOR U38004 ( .A(g_input[364]), .B(creg[364]), .Z(n36677) );
  XOR U38005 ( .A(n36678), .B(n36679), .Z(n36669) );
  ANDN U38006 ( .A(n36680), .B(n28562), .Z(n36679) );
  XOR U38007 ( .A(n36681), .B(\modmult_1/zin[0][362] ), .Z(n28562) );
  IV U38008 ( .A(n36678), .Z(n36681) );
  XNOR U38009 ( .A(n36678), .B(n28561), .Z(n36680) );
  XOR U38010 ( .A(n36682), .B(n36683), .Z(n28561) );
  AND U38011 ( .A(\modmult_1/xin[1023] ), .B(n36684), .Z(n36683) );
  IV U38012 ( .A(n36682), .Z(n36684) );
  XOR U38013 ( .A(n36685), .B(g_input[363]), .Z(n36682) );
  NAND U38014 ( .A(n36686), .B(mul_pow), .Z(n36685) );
  XOR U38015 ( .A(g_input[363]), .B(creg[363]), .Z(n36686) );
  XOR U38016 ( .A(n36687), .B(n36688), .Z(n36678) );
  ANDN U38017 ( .A(n36689), .B(n28568), .Z(n36688) );
  XOR U38018 ( .A(n36690), .B(\modmult_1/zin[0][361] ), .Z(n28568) );
  IV U38019 ( .A(n36687), .Z(n36690) );
  XNOR U38020 ( .A(n36687), .B(n28567), .Z(n36689) );
  XOR U38021 ( .A(n36691), .B(n36692), .Z(n28567) );
  AND U38022 ( .A(\modmult_1/xin[1023] ), .B(n36693), .Z(n36692) );
  IV U38023 ( .A(n36691), .Z(n36693) );
  XOR U38024 ( .A(n36694), .B(g_input[362]), .Z(n36691) );
  NAND U38025 ( .A(n36695), .B(mul_pow), .Z(n36694) );
  XOR U38026 ( .A(g_input[362]), .B(creg[362]), .Z(n36695) );
  XOR U38027 ( .A(n36696), .B(n36697), .Z(n36687) );
  ANDN U38028 ( .A(n36698), .B(n28574), .Z(n36697) );
  XOR U38029 ( .A(n36699), .B(\modmult_1/zin[0][360] ), .Z(n28574) );
  IV U38030 ( .A(n36696), .Z(n36699) );
  XNOR U38031 ( .A(n36696), .B(n28573), .Z(n36698) );
  XOR U38032 ( .A(n36700), .B(n36701), .Z(n28573) );
  AND U38033 ( .A(\modmult_1/xin[1023] ), .B(n36702), .Z(n36701) );
  IV U38034 ( .A(n36700), .Z(n36702) );
  XOR U38035 ( .A(n36703), .B(g_input[361]), .Z(n36700) );
  NAND U38036 ( .A(n36704), .B(mul_pow), .Z(n36703) );
  XOR U38037 ( .A(g_input[361]), .B(creg[361]), .Z(n36704) );
  XOR U38038 ( .A(n36705), .B(n36706), .Z(n36696) );
  ANDN U38039 ( .A(n36707), .B(n28580), .Z(n36706) );
  XOR U38040 ( .A(n36708), .B(\modmult_1/zin[0][359] ), .Z(n28580) );
  IV U38041 ( .A(n36705), .Z(n36708) );
  XNOR U38042 ( .A(n36705), .B(n28579), .Z(n36707) );
  XOR U38043 ( .A(n36709), .B(n36710), .Z(n28579) );
  AND U38044 ( .A(\modmult_1/xin[1023] ), .B(n36711), .Z(n36710) );
  IV U38045 ( .A(n36709), .Z(n36711) );
  XOR U38046 ( .A(n36712), .B(g_input[360]), .Z(n36709) );
  NAND U38047 ( .A(n36713), .B(mul_pow), .Z(n36712) );
  XOR U38048 ( .A(g_input[360]), .B(creg[360]), .Z(n36713) );
  XOR U38049 ( .A(n36714), .B(n36715), .Z(n36705) );
  ANDN U38050 ( .A(n36716), .B(n28586), .Z(n36715) );
  XOR U38051 ( .A(n36717), .B(\modmult_1/zin[0][358] ), .Z(n28586) );
  IV U38052 ( .A(n36714), .Z(n36717) );
  XNOR U38053 ( .A(n36714), .B(n28585), .Z(n36716) );
  XOR U38054 ( .A(n36718), .B(n36719), .Z(n28585) );
  AND U38055 ( .A(\modmult_1/xin[1023] ), .B(n36720), .Z(n36719) );
  IV U38056 ( .A(n36718), .Z(n36720) );
  XOR U38057 ( .A(n36721), .B(g_input[359]), .Z(n36718) );
  NAND U38058 ( .A(n36722), .B(mul_pow), .Z(n36721) );
  XOR U38059 ( .A(g_input[359]), .B(creg[359]), .Z(n36722) );
  XOR U38060 ( .A(n36723), .B(n36724), .Z(n36714) );
  ANDN U38061 ( .A(n36725), .B(n28592), .Z(n36724) );
  XOR U38062 ( .A(n36726), .B(\modmult_1/zin[0][357] ), .Z(n28592) );
  IV U38063 ( .A(n36723), .Z(n36726) );
  XNOR U38064 ( .A(n36723), .B(n28591), .Z(n36725) );
  XOR U38065 ( .A(n36727), .B(n36728), .Z(n28591) );
  AND U38066 ( .A(\modmult_1/xin[1023] ), .B(n36729), .Z(n36728) );
  IV U38067 ( .A(n36727), .Z(n36729) );
  XOR U38068 ( .A(n36730), .B(g_input[358]), .Z(n36727) );
  NAND U38069 ( .A(n36731), .B(mul_pow), .Z(n36730) );
  XOR U38070 ( .A(g_input[358]), .B(creg[358]), .Z(n36731) );
  XOR U38071 ( .A(n36732), .B(n36733), .Z(n36723) );
  ANDN U38072 ( .A(n36734), .B(n28598), .Z(n36733) );
  XOR U38073 ( .A(n36735), .B(\modmult_1/zin[0][356] ), .Z(n28598) );
  IV U38074 ( .A(n36732), .Z(n36735) );
  XNOR U38075 ( .A(n36732), .B(n28597), .Z(n36734) );
  XOR U38076 ( .A(n36736), .B(n36737), .Z(n28597) );
  AND U38077 ( .A(\modmult_1/xin[1023] ), .B(n36738), .Z(n36737) );
  IV U38078 ( .A(n36736), .Z(n36738) );
  XOR U38079 ( .A(n36739), .B(g_input[357]), .Z(n36736) );
  NAND U38080 ( .A(n36740), .B(mul_pow), .Z(n36739) );
  XOR U38081 ( .A(g_input[357]), .B(creg[357]), .Z(n36740) );
  XOR U38082 ( .A(n36741), .B(n36742), .Z(n36732) );
  ANDN U38083 ( .A(n36743), .B(n28604), .Z(n36742) );
  XOR U38084 ( .A(n36744), .B(\modmult_1/zin[0][355] ), .Z(n28604) );
  IV U38085 ( .A(n36741), .Z(n36744) );
  XNOR U38086 ( .A(n36741), .B(n28603), .Z(n36743) );
  XOR U38087 ( .A(n36745), .B(n36746), .Z(n28603) );
  AND U38088 ( .A(\modmult_1/xin[1023] ), .B(n36747), .Z(n36746) );
  IV U38089 ( .A(n36745), .Z(n36747) );
  XOR U38090 ( .A(n36748), .B(g_input[356]), .Z(n36745) );
  NAND U38091 ( .A(n36749), .B(mul_pow), .Z(n36748) );
  XOR U38092 ( .A(g_input[356]), .B(creg[356]), .Z(n36749) );
  XOR U38093 ( .A(n36750), .B(n36751), .Z(n36741) );
  ANDN U38094 ( .A(n36752), .B(n28610), .Z(n36751) );
  XOR U38095 ( .A(n36753), .B(\modmult_1/zin[0][354] ), .Z(n28610) );
  IV U38096 ( .A(n36750), .Z(n36753) );
  XNOR U38097 ( .A(n36750), .B(n28609), .Z(n36752) );
  XOR U38098 ( .A(n36754), .B(n36755), .Z(n28609) );
  AND U38099 ( .A(\modmult_1/xin[1023] ), .B(n36756), .Z(n36755) );
  IV U38100 ( .A(n36754), .Z(n36756) );
  XOR U38101 ( .A(n36757), .B(g_input[355]), .Z(n36754) );
  NAND U38102 ( .A(n36758), .B(mul_pow), .Z(n36757) );
  XOR U38103 ( .A(g_input[355]), .B(creg[355]), .Z(n36758) );
  XOR U38104 ( .A(n36759), .B(n36760), .Z(n36750) );
  ANDN U38105 ( .A(n36761), .B(n28616), .Z(n36760) );
  XOR U38106 ( .A(n36762), .B(\modmult_1/zin[0][353] ), .Z(n28616) );
  IV U38107 ( .A(n36759), .Z(n36762) );
  XNOR U38108 ( .A(n36759), .B(n28615), .Z(n36761) );
  XOR U38109 ( .A(n36763), .B(n36764), .Z(n28615) );
  AND U38110 ( .A(\modmult_1/xin[1023] ), .B(n36765), .Z(n36764) );
  IV U38111 ( .A(n36763), .Z(n36765) );
  XOR U38112 ( .A(n36766), .B(g_input[354]), .Z(n36763) );
  NAND U38113 ( .A(n36767), .B(mul_pow), .Z(n36766) );
  XOR U38114 ( .A(g_input[354]), .B(creg[354]), .Z(n36767) );
  XOR U38115 ( .A(n36768), .B(n36769), .Z(n36759) );
  ANDN U38116 ( .A(n36770), .B(n28622), .Z(n36769) );
  XOR U38117 ( .A(n36771), .B(\modmult_1/zin[0][352] ), .Z(n28622) );
  IV U38118 ( .A(n36768), .Z(n36771) );
  XNOR U38119 ( .A(n36768), .B(n28621), .Z(n36770) );
  XOR U38120 ( .A(n36772), .B(n36773), .Z(n28621) );
  AND U38121 ( .A(\modmult_1/xin[1023] ), .B(n36774), .Z(n36773) );
  IV U38122 ( .A(n36772), .Z(n36774) );
  XOR U38123 ( .A(n36775), .B(g_input[353]), .Z(n36772) );
  NAND U38124 ( .A(n36776), .B(mul_pow), .Z(n36775) );
  XOR U38125 ( .A(g_input[353]), .B(creg[353]), .Z(n36776) );
  XOR U38126 ( .A(n36777), .B(n36778), .Z(n36768) );
  ANDN U38127 ( .A(n36779), .B(n28628), .Z(n36778) );
  XOR U38128 ( .A(n36780), .B(\modmult_1/zin[0][351] ), .Z(n28628) );
  IV U38129 ( .A(n36777), .Z(n36780) );
  XNOR U38130 ( .A(n36777), .B(n28627), .Z(n36779) );
  XOR U38131 ( .A(n36781), .B(n36782), .Z(n28627) );
  AND U38132 ( .A(\modmult_1/xin[1023] ), .B(n36783), .Z(n36782) );
  IV U38133 ( .A(n36781), .Z(n36783) );
  XOR U38134 ( .A(n36784), .B(g_input[352]), .Z(n36781) );
  NAND U38135 ( .A(n36785), .B(mul_pow), .Z(n36784) );
  XOR U38136 ( .A(g_input[352]), .B(creg[352]), .Z(n36785) );
  XOR U38137 ( .A(n36786), .B(n36787), .Z(n36777) );
  ANDN U38138 ( .A(n36788), .B(n28634), .Z(n36787) );
  XOR U38139 ( .A(n36789), .B(\modmult_1/zin[0][350] ), .Z(n28634) );
  IV U38140 ( .A(n36786), .Z(n36789) );
  XNOR U38141 ( .A(n36786), .B(n28633), .Z(n36788) );
  XOR U38142 ( .A(n36790), .B(n36791), .Z(n28633) );
  AND U38143 ( .A(\modmult_1/xin[1023] ), .B(n36792), .Z(n36791) );
  IV U38144 ( .A(n36790), .Z(n36792) );
  XOR U38145 ( .A(n36793), .B(g_input[351]), .Z(n36790) );
  NAND U38146 ( .A(n36794), .B(mul_pow), .Z(n36793) );
  XOR U38147 ( .A(g_input[351]), .B(creg[351]), .Z(n36794) );
  XOR U38148 ( .A(n36795), .B(n36796), .Z(n36786) );
  ANDN U38149 ( .A(n36797), .B(n28640), .Z(n36796) );
  XOR U38150 ( .A(n36798), .B(\modmult_1/zin[0][349] ), .Z(n28640) );
  IV U38151 ( .A(n36795), .Z(n36798) );
  XNOR U38152 ( .A(n36795), .B(n28639), .Z(n36797) );
  XOR U38153 ( .A(n36799), .B(n36800), .Z(n28639) );
  AND U38154 ( .A(\modmult_1/xin[1023] ), .B(n36801), .Z(n36800) );
  IV U38155 ( .A(n36799), .Z(n36801) );
  XOR U38156 ( .A(n36802), .B(g_input[350]), .Z(n36799) );
  NAND U38157 ( .A(n36803), .B(mul_pow), .Z(n36802) );
  XOR U38158 ( .A(g_input[350]), .B(creg[350]), .Z(n36803) );
  XOR U38159 ( .A(n36804), .B(n36805), .Z(n36795) );
  ANDN U38160 ( .A(n36806), .B(n28646), .Z(n36805) );
  XOR U38161 ( .A(n36807), .B(\modmult_1/zin[0][348] ), .Z(n28646) );
  IV U38162 ( .A(n36804), .Z(n36807) );
  XNOR U38163 ( .A(n36804), .B(n28645), .Z(n36806) );
  XOR U38164 ( .A(n36808), .B(n36809), .Z(n28645) );
  AND U38165 ( .A(\modmult_1/xin[1023] ), .B(n36810), .Z(n36809) );
  IV U38166 ( .A(n36808), .Z(n36810) );
  XOR U38167 ( .A(n36811), .B(g_input[349]), .Z(n36808) );
  NAND U38168 ( .A(n36812), .B(mul_pow), .Z(n36811) );
  XOR U38169 ( .A(g_input[349]), .B(creg[349]), .Z(n36812) );
  XOR U38170 ( .A(n36813), .B(n36814), .Z(n36804) );
  ANDN U38171 ( .A(n36815), .B(n28652), .Z(n36814) );
  XOR U38172 ( .A(n36816), .B(\modmult_1/zin[0][347] ), .Z(n28652) );
  IV U38173 ( .A(n36813), .Z(n36816) );
  XNOR U38174 ( .A(n36813), .B(n28651), .Z(n36815) );
  XOR U38175 ( .A(n36817), .B(n36818), .Z(n28651) );
  AND U38176 ( .A(\modmult_1/xin[1023] ), .B(n36819), .Z(n36818) );
  IV U38177 ( .A(n36817), .Z(n36819) );
  XOR U38178 ( .A(n36820), .B(g_input[348]), .Z(n36817) );
  NAND U38179 ( .A(n36821), .B(mul_pow), .Z(n36820) );
  XOR U38180 ( .A(g_input[348]), .B(creg[348]), .Z(n36821) );
  XOR U38181 ( .A(n36822), .B(n36823), .Z(n36813) );
  ANDN U38182 ( .A(n36824), .B(n28658), .Z(n36823) );
  XOR U38183 ( .A(n36825), .B(\modmult_1/zin[0][346] ), .Z(n28658) );
  IV U38184 ( .A(n36822), .Z(n36825) );
  XNOR U38185 ( .A(n36822), .B(n28657), .Z(n36824) );
  XOR U38186 ( .A(n36826), .B(n36827), .Z(n28657) );
  AND U38187 ( .A(\modmult_1/xin[1023] ), .B(n36828), .Z(n36827) );
  IV U38188 ( .A(n36826), .Z(n36828) );
  XOR U38189 ( .A(n36829), .B(g_input[347]), .Z(n36826) );
  NAND U38190 ( .A(n36830), .B(mul_pow), .Z(n36829) );
  XOR U38191 ( .A(g_input[347]), .B(creg[347]), .Z(n36830) );
  XOR U38192 ( .A(n36831), .B(n36832), .Z(n36822) );
  ANDN U38193 ( .A(n36833), .B(n28664), .Z(n36832) );
  XOR U38194 ( .A(n36834), .B(\modmult_1/zin[0][345] ), .Z(n28664) );
  IV U38195 ( .A(n36831), .Z(n36834) );
  XNOR U38196 ( .A(n36831), .B(n28663), .Z(n36833) );
  XOR U38197 ( .A(n36835), .B(n36836), .Z(n28663) );
  AND U38198 ( .A(\modmult_1/xin[1023] ), .B(n36837), .Z(n36836) );
  IV U38199 ( .A(n36835), .Z(n36837) );
  XOR U38200 ( .A(n36838), .B(g_input[346]), .Z(n36835) );
  NAND U38201 ( .A(n36839), .B(mul_pow), .Z(n36838) );
  XOR U38202 ( .A(g_input[346]), .B(creg[346]), .Z(n36839) );
  XOR U38203 ( .A(n36840), .B(n36841), .Z(n36831) );
  ANDN U38204 ( .A(n36842), .B(n28670), .Z(n36841) );
  XOR U38205 ( .A(n36843), .B(\modmult_1/zin[0][344] ), .Z(n28670) );
  IV U38206 ( .A(n36840), .Z(n36843) );
  XNOR U38207 ( .A(n36840), .B(n28669), .Z(n36842) );
  XOR U38208 ( .A(n36844), .B(n36845), .Z(n28669) );
  AND U38209 ( .A(\modmult_1/xin[1023] ), .B(n36846), .Z(n36845) );
  IV U38210 ( .A(n36844), .Z(n36846) );
  XOR U38211 ( .A(n36847), .B(g_input[345]), .Z(n36844) );
  NAND U38212 ( .A(n36848), .B(mul_pow), .Z(n36847) );
  XOR U38213 ( .A(g_input[345]), .B(creg[345]), .Z(n36848) );
  XOR U38214 ( .A(n36849), .B(n36850), .Z(n36840) );
  ANDN U38215 ( .A(n36851), .B(n28676), .Z(n36850) );
  XOR U38216 ( .A(n36852), .B(\modmult_1/zin[0][343] ), .Z(n28676) );
  IV U38217 ( .A(n36849), .Z(n36852) );
  XNOR U38218 ( .A(n36849), .B(n28675), .Z(n36851) );
  XOR U38219 ( .A(n36853), .B(n36854), .Z(n28675) );
  AND U38220 ( .A(\modmult_1/xin[1023] ), .B(n36855), .Z(n36854) );
  IV U38221 ( .A(n36853), .Z(n36855) );
  XOR U38222 ( .A(n36856), .B(g_input[344]), .Z(n36853) );
  NAND U38223 ( .A(n36857), .B(mul_pow), .Z(n36856) );
  XOR U38224 ( .A(g_input[344]), .B(creg[344]), .Z(n36857) );
  XOR U38225 ( .A(n36858), .B(n36859), .Z(n36849) );
  ANDN U38226 ( .A(n36860), .B(n28682), .Z(n36859) );
  XOR U38227 ( .A(n36861), .B(\modmult_1/zin[0][342] ), .Z(n28682) );
  IV U38228 ( .A(n36858), .Z(n36861) );
  XNOR U38229 ( .A(n36858), .B(n28681), .Z(n36860) );
  XOR U38230 ( .A(n36862), .B(n36863), .Z(n28681) );
  AND U38231 ( .A(\modmult_1/xin[1023] ), .B(n36864), .Z(n36863) );
  IV U38232 ( .A(n36862), .Z(n36864) );
  XOR U38233 ( .A(n36865), .B(g_input[343]), .Z(n36862) );
  NAND U38234 ( .A(n36866), .B(mul_pow), .Z(n36865) );
  XOR U38235 ( .A(g_input[343]), .B(creg[343]), .Z(n36866) );
  XOR U38236 ( .A(n36867), .B(n36868), .Z(n36858) );
  ANDN U38237 ( .A(n36869), .B(n28688), .Z(n36868) );
  XOR U38238 ( .A(n36870), .B(\modmult_1/zin[0][341] ), .Z(n28688) );
  IV U38239 ( .A(n36867), .Z(n36870) );
  XNOR U38240 ( .A(n36867), .B(n28687), .Z(n36869) );
  XOR U38241 ( .A(n36871), .B(n36872), .Z(n28687) );
  AND U38242 ( .A(\modmult_1/xin[1023] ), .B(n36873), .Z(n36872) );
  IV U38243 ( .A(n36871), .Z(n36873) );
  XOR U38244 ( .A(n36874), .B(g_input[342]), .Z(n36871) );
  NAND U38245 ( .A(n36875), .B(mul_pow), .Z(n36874) );
  XOR U38246 ( .A(g_input[342]), .B(creg[342]), .Z(n36875) );
  XOR U38247 ( .A(n36876), .B(n36877), .Z(n36867) );
  ANDN U38248 ( .A(n36878), .B(n28694), .Z(n36877) );
  XOR U38249 ( .A(n36879), .B(\modmult_1/zin[0][340] ), .Z(n28694) );
  IV U38250 ( .A(n36876), .Z(n36879) );
  XNOR U38251 ( .A(n36876), .B(n28693), .Z(n36878) );
  XOR U38252 ( .A(n36880), .B(n36881), .Z(n28693) );
  AND U38253 ( .A(\modmult_1/xin[1023] ), .B(n36882), .Z(n36881) );
  IV U38254 ( .A(n36880), .Z(n36882) );
  XOR U38255 ( .A(n36883), .B(g_input[341]), .Z(n36880) );
  NAND U38256 ( .A(n36884), .B(mul_pow), .Z(n36883) );
  XOR U38257 ( .A(g_input[341]), .B(creg[341]), .Z(n36884) );
  XOR U38258 ( .A(n36885), .B(n36886), .Z(n36876) );
  ANDN U38259 ( .A(n36887), .B(n28700), .Z(n36886) );
  XOR U38260 ( .A(n36888), .B(\modmult_1/zin[0][339] ), .Z(n28700) );
  IV U38261 ( .A(n36885), .Z(n36888) );
  XNOR U38262 ( .A(n36885), .B(n28699), .Z(n36887) );
  XOR U38263 ( .A(n36889), .B(n36890), .Z(n28699) );
  AND U38264 ( .A(\modmult_1/xin[1023] ), .B(n36891), .Z(n36890) );
  IV U38265 ( .A(n36889), .Z(n36891) );
  XOR U38266 ( .A(n36892), .B(g_input[340]), .Z(n36889) );
  NAND U38267 ( .A(n36893), .B(mul_pow), .Z(n36892) );
  XOR U38268 ( .A(g_input[340]), .B(creg[340]), .Z(n36893) );
  XOR U38269 ( .A(n36894), .B(n36895), .Z(n36885) );
  ANDN U38270 ( .A(n36896), .B(n28706), .Z(n36895) );
  XOR U38271 ( .A(n36897), .B(\modmult_1/zin[0][338] ), .Z(n28706) );
  IV U38272 ( .A(n36894), .Z(n36897) );
  XNOR U38273 ( .A(n36894), .B(n28705), .Z(n36896) );
  XOR U38274 ( .A(n36898), .B(n36899), .Z(n28705) );
  AND U38275 ( .A(\modmult_1/xin[1023] ), .B(n36900), .Z(n36899) );
  IV U38276 ( .A(n36898), .Z(n36900) );
  XOR U38277 ( .A(n36901), .B(g_input[339]), .Z(n36898) );
  NAND U38278 ( .A(n36902), .B(mul_pow), .Z(n36901) );
  XOR U38279 ( .A(g_input[339]), .B(creg[339]), .Z(n36902) );
  XOR U38280 ( .A(n36903), .B(n36904), .Z(n36894) );
  ANDN U38281 ( .A(n36905), .B(n28712), .Z(n36904) );
  XOR U38282 ( .A(n36906), .B(\modmult_1/zin[0][337] ), .Z(n28712) );
  IV U38283 ( .A(n36903), .Z(n36906) );
  XNOR U38284 ( .A(n36903), .B(n28711), .Z(n36905) );
  XOR U38285 ( .A(n36907), .B(n36908), .Z(n28711) );
  AND U38286 ( .A(\modmult_1/xin[1023] ), .B(n36909), .Z(n36908) );
  IV U38287 ( .A(n36907), .Z(n36909) );
  XOR U38288 ( .A(n36910), .B(g_input[338]), .Z(n36907) );
  NAND U38289 ( .A(n36911), .B(mul_pow), .Z(n36910) );
  XOR U38290 ( .A(g_input[338]), .B(creg[338]), .Z(n36911) );
  XOR U38291 ( .A(n36912), .B(n36913), .Z(n36903) );
  ANDN U38292 ( .A(n36914), .B(n28718), .Z(n36913) );
  XOR U38293 ( .A(n36915), .B(\modmult_1/zin[0][336] ), .Z(n28718) );
  IV U38294 ( .A(n36912), .Z(n36915) );
  XNOR U38295 ( .A(n36912), .B(n28717), .Z(n36914) );
  XOR U38296 ( .A(n36916), .B(n36917), .Z(n28717) );
  AND U38297 ( .A(\modmult_1/xin[1023] ), .B(n36918), .Z(n36917) );
  IV U38298 ( .A(n36916), .Z(n36918) );
  XOR U38299 ( .A(n36919), .B(g_input[337]), .Z(n36916) );
  NAND U38300 ( .A(n36920), .B(mul_pow), .Z(n36919) );
  XOR U38301 ( .A(g_input[337]), .B(creg[337]), .Z(n36920) );
  XOR U38302 ( .A(n36921), .B(n36922), .Z(n36912) );
  ANDN U38303 ( .A(n36923), .B(n28724), .Z(n36922) );
  XOR U38304 ( .A(n36924), .B(\modmult_1/zin[0][335] ), .Z(n28724) );
  IV U38305 ( .A(n36921), .Z(n36924) );
  XNOR U38306 ( .A(n36921), .B(n28723), .Z(n36923) );
  XOR U38307 ( .A(n36925), .B(n36926), .Z(n28723) );
  AND U38308 ( .A(\modmult_1/xin[1023] ), .B(n36927), .Z(n36926) );
  IV U38309 ( .A(n36925), .Z(n36927) );
  XOR U38310 ( .A(n36928), .B(g_input[336]), .Z(n36925) );
  NAND U38311 ( .A(n36929), .B(mul_pow), .Z(n36928) );
  XOR U38312 ( .A(g_input[336]), .B(creg[336]), .Z(n36929) );
  XOR U38313 ( .A(n36930), .B(n36931), .Z(n36921) );
  ANDN U38314 ( .A(n36932), .B(n28730), .Z(n36931) );
  XOR U38315 ( .A(n36933), .B(\modmult_1/zin[0][334] ), .Z(n28730) );
  IV U38316 ( .A(n36930), .Z(n36933) );
  XNOR U38317 ( .A(n36930), .B(n28729), .Z(n36932) );
  XOR U38318 ( .A(n36934), .B(n36935), .Z(n28729) );
  AND U38319 ( .A(\modmult_1/xin[1023] ), .B(n36936), .Z(n36935) );
  IV U38320 ( .A(n36934), .Z(n36936) );
  XOR U38321 ( .A(n36937), .B(g_input[335]), .Z(n36934) );
  NAND U38322 ( .A(n36938), .B(mul_pow), .Z(n36937) );
  XOR U38323 ( .A(g_input[335]), .B(creg[335]), .Z(n36938) );
  XOR U38324 ( .A(n36939), .B(n36940), .Z(n36930) );
  ANDN U38325 ( .A(n36941), .B(n28736), .Z(n36940) );
  XOR U38326 ( .A(n36942), .B(\modmult_1/zin[0][333] ), .Z(n28736) );
  IV U38327 ( .A(n36939), .Z(n36942) );
  XNOR U38328 ( .A(n36939), .B(n28735), .Z(n36941) );
  XOR U38329 ( .A(n36943), .B(n36944), .Z(n28735) );
  AND U38330 ( .A(\modmult_1/xin[1023] ), .B(n36945), .Z(n36944) );
  IV U38331 ( .A(n36943), .Z(n36945) );
  XOR U38332 ( .A(n36946), .B(g_input[334]), .Z(n36943) );
  NAND U38333 ( .A(n36947), .B(mul_pow), .Z(n36946) );
  XOR U38334 ( .A(g_input[334]), .B(creg[334]), .Z(n36947) );
  XOR U38335 ( .A(n36948), .B(n36949), .Z(n36939) );
  ANDN U38336 ( .A(n36950), .B(n28742), .Z(n36949) );
  XOR U38337 ( .A(n36951), .B(\modmult_1/zin[0][332] ), .Z(n28742) );
  IV U38338 ( .A(n36948), .Z(n36951) );
  XNOR U38339 ( .A(n36948), .B(n28741), .Z(n36950) );
  XOR U38340 ( .A(n36952), .B(n36953), .Z(n28741) );
  AND U38341 ( .A(\modmult_1/xin[1023] ), .B(n36954), .Z(n36953) );
  IV U38342 ( .A(n36952), .Z(n36954) );
  XOR U38343 ( .A(n36955), .B(g_input[333]), .Z(n36952) );
  NAND U38344 ( .A(n36956), .B(mul_pow), .Z(n36955) );
  XOR U38345 ( .A(g_input[333]), .B(creg[333]), .Z(n36956) );
  XOR U38346 ( .A(n36957), .B(n36958), .Z(n36948) );
  ANDN U38347 ( .A(n36959), .B(n28748), .Z(n36958) );
  XOR U38348 ( .A(n36960), .B(\modmult_1/zin[0][331] ), .Z(n28748) );
  IV U38349 ( .A(n36957), .Z(n36960) );
  XNOR U38350 ( .A(n36957), .B(n28747), .Z(n36959) );
  XOR U38351 ( .A(n36961), .B(n36962), .Z(n28747) );
  AND U38352 ( .A(\modmult_1/xin[1023] ), .B(n36963), .Z(n36962) );
  IV U38353 ( .A(n36961), .Z(n36963) );
  XOR U38354 ( .A(n36964), .B(g_input[332]), .Z(n36961) );
  NAND U38355 ( .A(n36965), .B(mul_pow), .Z(n36964) );
  XOR U38356 ( .A(g_input[332]), .B(creg[332]), .Z(n36965) );
  XOR U38357 ( .A(n36966), .B(n36967), .Z(n36957) );
  ANDN U38358 ( .A(n36968), .B(n28754), .Z(n36967) );
  XOR U38359 ( .A(n36969), .B(\modmult_1/zin[0][330] ), .Z(n28754) );
  IV U38360 ( .A(n36966), .Z(n36969) );
  XNOR U38361 ( .A(n36966), .B(n28753), .Z(n36968) );
  XOR U38362 ( .A(n36970), .B(n36971), .Z(n28753) );
  AND U38363 ( .A(\modmult_1/xin[1023] ), .B(n36972), .Z(n36971) );
  IV U38364 ( .A(n36970), .Z(n36972) );
  XOR U38365 ( .A(n36973), .B(g_input[331]), .Z(n36970) );
  NAND U38366 ( .A(n36974), .B(mul_pow), .Z(n36973) );
  XOR U38367 ( .A(g_input[331]), .B(creg[331]), .Z(n36974) );
  XOR U38368 ( .A(n36975), .B(n36976), .Z(n36966) );
  ANDN U38369 ( .A(n36977), .B(n28760), .Z(n36976) );
  XOR U38370 ( .A(n36978), .B(\modmult_1/zin[0][329] ), .Z(n28760) );
  IV U38371 ( .A(n36975), .Z(n36978) );
  XNOR U38372 ( .A(n36975), .B(n28759), .Z(n36977) );
  XOR U38373 ( .A(n36979), .B(n36980), .Z(n28759) );
  AND U38374 ( .A(\modmult_1/xin[1023] ), .B(n36981), .Z(n36980) );
  IV U38375 ( .A(n36979), .Z(n36981) );
  XOR U38376 ( .A(n36982), .B(g_input[330]), .Z(n36979) );
  NAND U38377 ( .A(n36983), .B(mul_pow), .Z(n36982) );
  XOR U38378 ( .A(g_input[330]), .B(creg[330]), .Z(n36983) );
  XOR U38379 ( .A(n36984), .B(n36985), .Z(n36975) );
  ANDN U38380 ( .A(n36986), .B(n28766), .Z(n36985) );
  XOR U38381 ( .A(n36987), .B(\modmult_1/zin[0][328] ), .Z(n28766) );
  IV U38382 ( .A(n36984), .Z(n36987) );
  XNOR U38383 ( .A(n36984), .B(n28765), .Z(n36986) );
  XOR U38384 ( .A(n36988), .B(n36989), .Z(n28765) );
  AND U38385 ( .A(\modmult_1/xin[1023] ), .B(n36990), .Z(n36989) );
  IV U38386 ( .A(n36988), .Z(n36990) );
  XOR U38387 ( .A(n36991), .B(g_input[329]), .Z(n36988) );
  NAND U38388 ( .A(n36992), .B(mul_pow), .Z(n36991) );
  XOR U38389 ( .A(g_input[329]), .B(creg[329]), .Z(n36992) );
  XOR U38390 ( .A(n36993), .B(n36994), .Z(n36984) );
  ANDN U38391 ( .A(n36995), .B(n28772), .Z(n36994) );
  XOR U38392 ( .A(n36996), .B(\modmult_1/zin[0][327] ), .Z(n28772) );
  IV U38393 ( .A(n36993), .Z(n36996) );
  XNOR U38394 ( .A(n36993), .B(n28771), .Z(n36995) );
  XOR U38395 ( .A(n36997), .B(n36998), .Z(n28771) );
  AND U38396 ( .A(\modmult_1/xin[1023] ), .B(n36999), .Z(n36998) );
  IV U38397 ( .A(n36997), .Z(n36999) );
  XOR U38398 ( .A(n37000), .B(g_input[328]), .Z(n36997) );
  NAND U38399 ( .A(n37001), .B(mul_pow), .Z(n37000) );
  XOR U38400 ( .A(g_input[328]), .B(creg[328]), .Z(n37001) );
  XOR U38401 ( .A(n37002), .B(n37003), .Z(n36993) );
  ANDN U38402 ( .A(n37004), .B(n28778), .Z(n37003) );
  XOR U38403 ( .A(n37005), .B(\modmult_1/zin[0][326] ), .Z(n28778) );
  IV U38404 ( .A(n37002), .Z(n37005) );
  XNOR U38405 ( .A(n37002), .B(n28777), .Z(n37004) );
  XOR U38406 ( .A(n37006), .B(n37007), .Z(n28777) );
  AND U38407 ( .A(\modmult_1/xin[1023] ), .B(n37008), .Z(n37007) );
  IV U38408 ( .A(n37006), .Z(n37008) );
  XOR U38409 ( .A(n37009), .B(g_input[327]), .Z(n37006) );
  NAND U38410 ( .A(n37010), .B(mul_pow), .Z(n37009) );
  XOR U38411 ( .A(g_input[327]), .B(creg[327]), .Z(n37010) );
  XOR U38412 ( .A(n37011), .B(n37012), .Z(n37002) );
  ANDN U38413 ( .A(n37013), .B(n28784), .Z(n37012) );
  XOR U38414 ( .A(n37014), .B(\modmult_1/zin[0][325] ), .Z(n28784) );
  IV U38415 ( .A(n37011), .Z(n37014) );
  XNOR U38416 ( .A(n37011), .B(n28783), .Z(n37013) );
  XOR U38417 ( .A(n37015), .B(n37016), .Z(n28783) );
  AND U38418 ( .A(\modmult_1/xin[1023] ), .B(n37017), .Z(n37016) );
  IV U38419 ( .A(n37015), .Z(n37017) );
  XOR U38420 ( .A(n37018), .B(g_input[326]), .Z(n37015) );
  NAND U38421 ( .A(n37019), .B(mul_pow), .Z(n37018) );
  XOR U38422 ( .A(g_input[326]), .B(creg[326]), .Z(n37019) );
  XOR U38423 ( .A(n37020), .B(n37021), .Z(n37011) );
  ANDN U38424 ( .A(n37022), .B(n28790), .Z(n37021) );
  XOR U38425 ( .A(n37023), .B(\modmult_1/zin[0][324] ), .Z(n28790) );
  IV U38426 ( .A(n37020), .Z(n37023) );
  XNOR U38427 ( .A(n37020), .B(n28789), .Z(n37022) );
  XOR U38428 ( .A(n37024), .B(n37025), .Z(n28789) );
  AND U38429 ( .A(\modmult_1/xin[1023] ), .B(n37026), .Z(n37025) );
  IV U38430 ( .A(n37024), .Z(n37026) );
  XOR U38431 ( .A(n37027), .B(g_input[325]), .Z(n37024) );
  NAND U38432 ( .A(n37028), .B(mul_pow), .Z(n37027) );
  XOR U38433 ( .A(g_input[325]), .B(creg[325]), .Z(n37028) );
  XOR U38434 ( .A(n37029), .B(n37030), .Z(n37020) );
  ANDN U38435 ( .A(n37031), .B(n28796), .Z(n37030) );
  XOR U38436 ( .A(n37032), .B(\modmult_1/zin[0][323] ), .Z(n28796) );
  IV U38437 ( .A(n37029), .Z(n37032) );
  XNOR U38438 ( .A(n37029), .B(n28795), .Z(n37031) );
  XOR U38439 ( .A(n37033), .B(n37034), .Z(n28795) );
  AND U38440 ( .A(\modmult_1/xin[1023] ), .B(n37035), .Z(n37034) );
  IV U38441 ( .A(n37033), .Z(n37035) );
  XOR U38442 ( .A(n37036), .B(g_input[324]), .Z(n37033) );
  NAND U38443 ( .A(n37037), .B(mul_pow), .Z(n37036) );
  XOR U38444 ( .A(g_input[324]), .B(creg[324]), .Z(n37037) );
  XOR U38445 ( .A(n37038), .B(n37039), .Z(n37029) );
  ANDN U38446 ( .A(n37040), .B(n28802), .Z(n37039) );
  XOR U38447 ( .A(n37041), .B(\modmult_1/zin[0][322] ), .Z(n28802) );
  IV U38448 ( .A(n37038), .Z(n37041) );
  XNOR U38449 ( .A(n37038), .B(n28801), .Z(n37040) );
  XOR U38450 ( .A(n37042), .B(n37043), .Z(n28801) );
  AND U38451 ( .A(\modmult_1/xin[1023] ), .B(n37044), .Z(n37043) );
  IV U38452 ( .A(n37042), .Z(n37044) );
  XOR U38453 ( .A(n37045), .B(g_input[323]), .Z(n37042) );
  NAND U38454 ( .A(n37046), .B(mul_pow), .Z(n37045) );
  XOR U38455 ( .A(g_input[323]), .B(creg[323]), .Z(n37046) );
  XOR U38456 ( .A(n37047), .B(n37048), .Z(n37038) );
  ANDN U38457 ( .A(n37049), .B(n28808), .Z(n37048) );
  XOR U38458 ( .A(n37050), .B(\modmult_1/zin[0][321] ), .Z(n28808) );
  IV U38459 ( .A(n37047), .Z(n37050) );
  XNOR U38460 ( .A(n37047), .B(n28807), .Z(n37049) );
  XOR U38461 ( .A(n37051), .B(n37052), .Z(n28807) );
  AND U38462 ( .A(\modmult_1/xin[1023] ), .B(n37053), .Z(n37052) );
  IV U38463 ( .A(n37051), .Z(n37053) );
  XOR U38464 ( .A(n37054), .B(g_input[322]), .Z(n37051) );
  NAND U38465 ( .A(n37055), .B(mul_pow), .Z(n37054) );
  XOR U38466 ( .A(g_input[322]), .B(creg[322]), .Z(n37055) );
  XOR U38467 ( .A(n37056), .B(n37057), .Z(n37047) );
  ANDN U38468 ( .A(n37058), .B(n28814), .Z(n37057) );
  XOR U38469 ( .A(n37059), .B(\modmult_1/zin[0][320] ), .Z(n28814) );
  IV U38470 ( .A(n37056), .Z(n37059) );
  XNOR U38471 ( .A(n37056), .B(n28813), .Z(n37058) );
  XOR U38472 ( .A(n37060), .B(n37061), .Z(n28813) );
  AND U38473 ( .A(\modmult_1/xin[1023] ), .B(n37062), .Z(n37061) );
  IV U38474 ( .A(n37060), .Z(n37062) );
  XOR U38475 ( .A(n37063), .B(g_input[321]), .Z(n37060) );
  NAND U38476 ( .A(n37064), .B(mul_pow), .Z(n37063) );
  XOR U38477 ( .A(g_input[321]), .B(creg[321]), .Z(n37064) );
  XOR U38478 ( .A(n37065), .B(n37066), .Z(n37056) );
  ANDN U38479 ( .A(n37067), .B(n28820), .Z(n37066) );
  XOR U38480 ( .A(n37068), .B(\modmult_1/zin[0][319] ), .Z(n28820) );
  IV U38481 ( .A(n37065), .Z(n37068) );
  XNOR U38482 ( .A(n37065), .B(n28819), .Z(n37067) );
  XOR U38483 ( .A(n37069), .B(n37070), .Z(n28819) );
  AND U38484 ( .A(\modmult_1/xin[1023] ), .B(n37071), .Z(n37070) );
  IV U38485 ( .A(n37069), .Z(n37071) );
  XOR U38486 ( .A(n37072), .B(g_input[320]), .Z(n37069) );
  NAND U38487 ( .A(n37073), .B(mul_pow), .Z(n37072) );
  XOR U38488 ( .A(g_input[320]), .B(creg[320]), .Z(n37073) );
  XOR U38489 ( .A(n37074), .B(n37075), .Z(n37065) );
  ANDN U38490 ( .A(n37076), .B(n28826), .Z(n37075) );
  XOR U38491 ( .A(n37077), .B(\modmult_1/zin[0][318] ), .Z(n28826) );
  IV U38492 ( .A(n37074), .Z(n37077) );
  XNOR U38493 ( .A(n37074), .B(n28825), .Z(n37076) );
  XOR U38494 ( .A(n37078), .B(n37079), .Z(n28825) );
  AND U38495 ( .A(\modmult_1/xin[1023] ), .B(n37080), .Z(n37079) );
  IV U38496 ( .A(n37078), .Z(n37080) );
  XOR U38497 ( .A(n37081), .B(g_input[319]), .Z(n37078) );
  NAND U38498 ( .A(n37082), .B(mul_pow), .Z(n37081) );
  XOR U38499 ( .A(g_input[319]), .B(creg[319]), .Z(n37082) );
  XOR U38500 ( .A(n37083), .B(n37084), .Z(n37074) );
  ANDN U38501 ( .A(n37085), .B(n28832), .Z(n37084) );
  XOR U38502 ( .A(n37086), .B(\modmult_1/zin[0][317] ), .Z(n28832) );
  IV U38503 ( .A(n37083), .Z(n37086) );
  XNOR U38504 ( .A(n37083), .B(n28831), .Z(n37085) );
  XOR U38505 ( .A(n37087), .B(n37088), .Z(n28831) );
  AND U38506 ( .A(\modmult_1/xin[1023] ), .B(n37089), .Z(n37088) );
  IV U38507 ( .A(n37087), .Z(n37089) );
  XOR U38508 ( .A(n37090), .B(g_input[318]), .Z(n37087) );
  NAND U38509 ( .A(n37091), .B(mul_pow), .Z(n37090) );
  XOR U38510 ( .A(g_input[318]), .B(creg[318]), .Z(n37091) );
  XOR U38511 ( .A(n37092), .B(n37093), .Z(n37083) );
  ANDN U38512 ( .A(n37094), .B(n28838), .Z(n37093) );
  XOR U38513 ( .A(n37095), .B(\modmult_1/zin[0][316] ), .Z(n28838) );
  IV U38514 ( .A(n37092), .Z(n37095) );
  XNOR U38515 ( .A(n37092), .B(n28837), .Z(n37094) );
  XOR U38516 ( .A(n37096), .B(n37097), .Z(n28837) );
  AND U38517 ( .A(\modmult_1/xin[1023] ), .B(n37098), .Z(n37097) );
  IV U38518 ( .A(n37096), .Z(n37098) );
  XOR U38519 ( .A(n37099), .B(g_input[317]), .Z(n37096) );
  NAND U38520 ( .A(n37100), .B(mul_pow), .Z(n37099) );
  XOR U38521 ( .A(g_input[317]), .B(creg[317]), .Z(n37100) );
  XOR U38522 ( .A(n37101), .B(n37102), .Z(n37092) );
  ANDN U38523 ( .A(n37103), .B(n28844), .Z(n37102) );
  XOR U38524 ( .A(n37104), .B(\modmult_1/zin[0][315] ), .Z(n28844) );
  IV U38525 ( .A(n37101), .Z(n37104) );
  XNOR U38526 ( .A(n37101), .B(n28843), .Z(n37103) );
  XOR U38527 ( .A(n37105), .B(n37106), .Z(n28843) );
  AND U38528 ( .A(\modmult_1/xin[1023] ), .B(n37107), .Z(n37106) );
  IV U38529 ( .A(n37105), .Z(n37107) );
  XOR U38530 ( .A(n37108), .B(g_input[316]), .Z(n37105) );
  NAND U38531 ( .A(n37109), .B(mul_pow), .Z(n37108) );
  XOR U38532 ( .A(g_input[316]), .B(creg[316]), .Z(n37109) );
  XOR U38533 ( .A(n37110), .B(n37111), .Z(n37101) );
  ANDN U38534 ( .A(n37112), .B(n28850), .Z(n37111) );
  XOR U38535 ( .A(n37113), .B(\modmult_1/zin[0][314] ), .Z(n28850) );
  IV U38536 ( .A(n37110), .Z(n37113) );
  XNOR U38537 ( .A(n37110), .B(n28849), .Z(n37112) );
  XOR U38538 ( .A(n37114), .B(n37115), .Z(n28849) );
  AND U38539 ( .A(\modmult_1/xin[1023] ), .B(n37116), .Z(n37115) );
  IV U38540 ( .A(n37114), .Z(n37116) );
  XOR U38541 ( .A(n37117), .B(g_input[315]), .Z(n37114) );
  NAND U38542 ( .A(n37118), .B(mul_pow), .Z(n37117) );
  XOR U38543 ( .A(g_input[315]), .B(creg[315]), .Z(n37118) );
  XOR U38544 ( .A(n37119), .B(n37120), .Z(n37110) );
  ANDN U38545 ( .A(n37121), .B(n28856), .Z(n37120) );
  XOR U38546 ( .A(n37122), .B(\modmult_1/zin[0][313] ), .Z(n28856) );
  IV U38547 ( .A(n37119), .Z(n37122) );
  XNOR U38548 ( .A(n37119), .B(n28855), .Z(n37121) );
  XOR U38549 ( .A(n37123), .B(n37124), .Z(n28855) );
  AND U38550 ( .A(\modmult_1/xin[1023] ), .B(n37125), .Z(n37124) );
  IV U38551 ( .A(n37123), .Z(n37125) );
  XOR U38552 ( .A(n37126), .B(g_input[314]), .Z(n37123) );
  NAND U38553 ( .A(n37127), .B(mul_pow), .Z(n37126) );
  XOR U38554 ( .A(g_input[314]), .B(creg[314]), .Z(n37127) );
  XOR U38555 ( .A(n37128), .B(n37129), .Z(n37119) );
  ANDN U38556 ( .A(n37130), .B(n28862), .Z(n37129) );
  XOR U38557 ( .A(n37131), .B(\modmult_1/zin[0][312] ), .Z(n28862) );
  IV U38558 ( .A(n37128), .Z(n37131) );
  XNOR U38559 ( .A(n37128), .B(n28861), .Z(n37130) );
  XOR U38560 ( .A(n37132), .B(n37133), .Z(n28861) );
  AND U38561 ( .A(\modmult_1/xin[1023] ), .B(n37134), .Z(n37133) );
  IV U38562 ( .A(n37132), .Z(n37134) );
  XOR U38563 ( .A(n37135), .B(g_input[313]), .Z(n37132) );
  NAND U38564 ( .A(n37136), .B(mul_pow), .Z(n37135) );
  XOR U38565 ( .A(g_input[313]), .B(creg[313]), .Z(n37136) );
  XOR U38566 ( .A(n37137), .B(n37138), .Z(n37128) );
  ANDN U38567 ( .A(n37139), .B(n28868), .Z(n37138) );
  XOR U38568 ( .A(n37140), .B(\modmult_1/zin[0][311] ), .Z(n28868) );
  IV U38569 ( .A(n37137), .Z(n37140) );
  XNOR U38570 ( .A(n37137), .B(n28867), .Z(n37139) );
  XOR U38571 ( .A(n37141), .B(n37142), .Z(n28867) );
  AND U38572 ( .A(\modmult_1/xin[1023] ), .B(n37143), .Z(n37142) );
  IV U38573 ( .A(n37141), .Z(n37143) );
  XOR U38574 ( .A(n37144), .B(g_input[312]), .Z(n37141) );
  NAND U38575 ( .A(n37145), .B(mul_pow), .Z(n37144) );
  XOR U38576 ( .A(g_input[312]), .B(creg[312]), .Z(n37145) );
  XOR U38577 ( .A(n37146), .B(n37147), .Z(n37137) );
  ANDN U38578 ( .A(n37148), .B(n28874), .Z(n37147) );
  XOR U38579 ( .A(n37149), .B(\modmult_1/zin[0][310] ), .Z(n28874) );
  IV U38580 ( .A(n37146), .Z(n37149) );
  XNOR U38581 ( .A(n37146), .B(n28873), .Z(n37148) );
  XOR U38582 ( .A(n37150), .B(n37151), .Z(n28873) );
  AND U38583 ( .A(\modmult_1/xin[1023] ), .B(n37152), .Z(n37151) );
  IV U38584 ( .A(n37150), .Z(n37152) );
  XOR U38585 ( .A(n37153), .B(g_input[311]), .Z(n37150) );
  NAND U38586 ( .A(n37154), .B(mul_pow), .Z(n37153) );
  XOR U38587 ( .A(g_input[311]), .B(creg[311]), .Z(n37154) );
  XOR U38588 ( .A(n37155), .B(n37156), .Z(n37146) );
  ANDN U38589 ( .A(n37157), .B(n28880), .Z(n37156) );
  XOR U38590 ( .A(n37158), .B(\modmult_1/zin[0][309] ), .Z(n28880) );
  IV U38591 ( .A(n37155), .Z(n37158) );
  XNOR U38592 ( .A(n37155), .B(n28879), .Z(n37157) );
  XOR U38593 ( .A(n37159), .B(n37160), .Z(n28879) );
  AND U38594 ( .A(\modmult_1/xin[1023] ), .B(n37161), .Z(n37160) );
  IV U38595 ( .A(n37159), .Z(n37161) );
  XOR U38596 ( .A(n37162), .B(g_input[310]), .Z(n37159) );
  NAND U38597 ( .A(n37163), .B(mul_pow), .Z(n37162) );
  XOR U38598 ( .A(g_input[310]), .B(creg[310]), .Z(n37163) );
  XOR U38599 ( .A(n37164), .B(n37165), .Z(n37155) );
  ANDN U38600 ( .A(n37166), .B(n28886), .Z(n37165) );
  XOR U38601 ( .A(n37167), .B(\modmult_1/zin[0][308] ), .Z(n28886) );
  IV U38602 ( .A(n37164), .Z(n37167) );
  XNOR U38603 ( .A(n37164), .B(n28885), .Z(n37166) );
  XOR U38604 ( .A(n37168), .B(n37169), .Z(n28885) );
  AND U38605 ( .A(\modmult_1/xin[1023] ), .B(n37170), .Z(n37169) );
  IV U38606 ( .A(n37168), .Z(n37170) );
  XOR U38607 ( .A(n37171), .B(g_input[309]), .Z(n37168) );
  NAND U38608 ( .A(n37172), .B(mul_pow), .Z(n37171) );
  XOR U38609 ( .A(g_input[309]), .B(creg[309]), .Z(n37172) );
  XOR U38610 ( .A(n37173), .B(n37174), .Z(n37164) );
  ANDN U38611 ( .A(n37175), .B(n28892), .Z(n37174) );
  XOR U38612 ( .A(n37176), .B(\modmult_1/zin[0][307] ), .Z(n28892) );
  IV U38613 ( .A(n37173), .Z(n37176) );
  XNOR U38614 ( .A(n37173), .B(n28891), .Z(n37175) );
  XOR U38615 ( .A(n37177), .B(n37178), .Z(n28891) );
  AND U38616 ( .A(\modmult_1/xin[1023] ), .B(n37179), .Z(n37178) );
  IV U38617 ( .A(n37177), .Z(n37179) );
  XOR U38618 ( .A(n37180), .B(g_input[308]), .Z(n37177) );
  NAND U38619 ( .A(n37181), .B(mul_pow), .Z(n37180) );
  XOR U38620 ( .A(g_input[308]), .B(creg[308]), .Z(n37181) );
  XOR U38621 ( .A(n37182), .B(n37183), .Z(n37173) );
  ANDN U38622 ( .A(n37184), .B(n28898), .Z(n37183) );
  XOR U38623 ( .A(n37185), .B(\modmult_1/zin[0][306] ), .Z(n28898) );
  IV U38624 ( .A(n37182), .Z(n37185) );
  XNOR U38625 ( .A(n37182), .B(n28897), .Z(n37184) );
  XOR U38626 ( .A(n37186), .B(n37187), .Z(n28897) );
  AND U38627 ( .A(\modmult_1/xin[1023] ), .B(n37188), .Z(n37187) );
  IV U38628 ( .A(n37186), .Z(n37188) );
  XOR U38629 ( .A(n37189), .B(g_input[307]), .Z(n37186) );
  NAND U38630 ( .A(n37190), .B(mul_pow), .Z(n37189) );
  XOR U38631 ( .A(g_input[307]), .B(creg[307]), .Z(n37190) );
  XOR U38632 ( .A(n37191), .B(n37192), .Z(n37182) );
  ANDN U38633 ( .A(n37193), .B(n28904), .Z(n37192) );
  XOR U38634 ( .A(n37194), .B(\modmult_1/zin[0][305] ), .Z(n28904) );
  IV U38635 ( .A(n37191), .Z(n37194) );
  XNOR U38636 ( .A(n37191), .B(n28903), .Z(n37193) );
  XOR U38637 ( .A(n37195), .B(n37196), .Z(n28903) );
  AND U38638 ( .A(\modmult_1/xin[1023] ), .B(n37197), .Z(n37196) );
  IV U38639 ( .A(n37195), .Z(n37197) );
  XOR U38640 ( .A(n37198), .B(g_input[306]), .Z(n37195) );
  NAND U38641 ( .A(n37199), .B(mul_pow), .Z(n37198) );
  XOR U38642 ( .A(g_input[306]), .B(creg[306]), .Z(n37199) );
  XOR U38643 ( .A(n37200), .B(n37201), .Z(n37191) );
  ANDN U38644 ( .A(n37202), .B(n28910), .Z(n37201) );
  XOR U38645 ( .A(n37203), .B(\modmult_1/zin[0][304] ), .Z(n28910) );
  IV U38646 ( .A(n37200), .Z(n37203) );
  XNOR U38647 ( .A(n37200), .B(n28909), .Z(n37202) );
  XOR U38648 ( .A(n37204), .B(n37205), .Z(n28909) );
  AND U38649 ( .A(\modmult_1/xin[1023] ), .B(n37206), .Z(n37205) );
  IV U38650 ( .A(n37204), .Z(n37206) );
  XOR U38651 ( .A(n37207), .B(g_input[305]), .Z(n37204) );
  NAND U38652 ( .A(n37208), .B(mul_pow), .Z(n37207) );
  XOR U38653 ( .A(g_input[305]), .B(creg[305]), .Z(n37208) );
  XOR U38654 ( .A(n37209), .B(n37210), .Z(n37200) );
  ANDN U38655 ( .A(n37211), .B(n28916), .Z(n37210) );
  XOR U38656 ( .A(n37212), .B(\modmult_1/zin[0][303] ), .Z(n28916) );
  IV U38657 ( .A(n37209), .Z(n37212) );
  XNOR U38658 ( .A(n37209), .B(n28915), .Z(n37211) );
  XOR U38659 ( .A(n37213), .B(n37214), .Z(n28915) );
  AND U38660 ( .A(\modmult_1/xin[1023] ), .B(n37215), .Z(n37214) );
  IV U38661 ( .A(n37213), .Z(n37215) );
  XOR U38662 ( .A(n37216), .B(g_input[304]), .Z(n37213) );
  NAND U38663 ( .A(n37217), .B(mul_pow), .Z(n37216) );
  XOR U38664 ( .A(g_input[304]), .B(creg[304]), .Z(n37217) );
  XOR U38665 ( .A(n37218), .B(n37219), .Z(n37209) );
  ANDN U38666 ( .A(n37220), .B(n28922), .Z(n37219) );
  XOR U38667 ( .A(n37221), .B(\modmult_1/zin[0][302] ), .Z(n28922) );
  IV U38668 ( .A(n37218), .Z(n37221) );
  XNOR U38669 ( .A(n37218), .B(n28921), .Z(n37220) );
  XOR U38670 ( .A(n37222), .B(n37223), .Z(n28921) );
  AND U38671 ( .A(\modmult_1/xin[1023] ), .B(n37224), .Z(n37223) );
  IV U38672 ( .A(n37222), .Z(n37224) );
  XOR U38673 ( .A(n37225), .B(g_input[303]), .Z(n37222) );
  NAND U38674 ( .A(n37226), .B(mul_pow), .Z(n37225) );
  XOR U38675 ( .A(g_input[303]), .B(creg[303]), .Z(n37226) );
  XOR U38676 ( .A(n37227), .B(n37228), .Z(n37218) );
  ANDN U38677 ( .A(n37229), .B(n28928), .Z(n37228) );
  XOR U38678 ( .A(n37230), .B(\modmult_1/zin[0][301] ), .Z(n28928) );
  IV U38679 ( .A(n37227), .Z(n37230) );
  XNOR U38680 ( .A(n37227), .B(n28927), .Z(n37229) );
  XOR U38681 ( .A(n37231), .B(n37232), .Z(n28927) );
  AND U38682 ( .A(\modmult_1/xin[1023] ), .B(n37233), .Z(n37232) );
  IV U38683 ( .A(n37231), .Z(n37233) );
  XOR U38684 ( .A(n37234), .B(g_input[302]), .Z(n37231) );
  NAND U38685 ( .A(n37235), .B(mul_pow), .Z(n37234) );
  XOR U38686 ( .A(g_input[302]), .B(creg[302]), .Z(n37235) );
  XOR U38687 ( .A(n37236), .B(n37237), .Z(n37227) );
  ANDN U38688 ( .A(n37238), .B(n28934), .Z(n37237) );
  XOR U38689 ( .A(n37239), .B(\modmult_1/zin[0][300] ), .Z(n28934) );
  IV U38690 ( .A(n37236), .Z(n37239) );
  XNOR U38691 ( .A(n37236), .B(n28933), .Z(n37238) );
  XOR U38692 ( .A(n37240), .B(n37241), .Z(n28933) );
  AND U38693 ( .A(\modmult_1/xin[1023] ), .B(n37242), .Z(n37241) );
  IV U38694 ( .A(n37240), .Z(n37242) );
  XOR U38695 ( .A(n37243), .B(g_input[301]), .Z(n37240) );
  NAND U38696 ( .A(n37244), .B(mul_pow), .Z(n37243) );
  XOR U38697 ( .A(g_input[301]), .B(creg[301]), .Z(n37244) );
  XOR U38698 ( .A(n37245), .B(n37246), .Z(n37236) );
  ANDN U38699 ( .A(n37247), .B(n28940), .Z(n37246) );
  XOR U38700 ( .A(n37248), .B(\modmult_1/zin[0][299] ), .Z(n28940) );
  IV U38701 ( .A(n37245), .Z(n37248) );
  XNOR U38702 ( .A(n37245), .B(n28939), .Z(n37247) );
  XOR U38703 ( .A(n37249), .B(n37250), .Z(n28939) );
  AND U38704 ( .A(\modmult_1/xin[1023] ), .B(n37251), .Z(n37250) );
  IV U38705 ( .A(n37249), .Z(n37251) );
  XOR U38706 ( .A(n37252), .B(g_input[300]), .Z(n37249) );
  NAND U38707 ( .A(n37253), .B(mul_pow), .Z(n37252) );
  XOR U38708 ( .A(g_input[300]), .B(creg[300]), .Z(n37253) );
  XOR U38709 ( .A(n37254), .B(n37255), .Z(n37245) );
  ANDN U38710 ( .A(n37256), .B(n28946), .Z(n37255) );
  XOR U38711 ( .A(n37257), .B(\modmult_1/zin[0][298] ), .Z(n28946) );
  IV U38712 ( .A(n37254), .Z(n37257) );
  XNOR U38713 ( .A(n37254), .B(n28945), .Z(n37256) );
  XOR U38714 ( .A(n37258), .B(n37259), .Z(n28945) );
  AND U38715 ( .A(\modmult_1/xin[1023] ), .B(n37260), .Z(n37259) );
  IV U38716 ( .A(n37258), .Z(n37260) );
  XOR U38717 ( .A(n37261), .B(g_input[299]), .Z(n37258) );
  NAND U38718 ( .A(n37262), .B(mul_pow), .Z(n37261) );
  XOR U38719 ( .A(g_input[299]), .B(creg[299]), .Z(n37262) );
  XOR U38720 ( .A(n37263), .B(n37264), .Z(n37254) );
  ANDN U38721 ( .A(n37265), .B(n28952), .Z(n37264) );
  XOR U38722 ( .A(n37266), .B(\modmult_1/zin[0][297] ), .Z(n28952) );
  IV U38723 ( .A(n37263), .Z(n37266) );
  XNOR U38724 ( .A(n37263), .B(n28951), .Z(n37265) );
  XOR U38725 ( .A(n37267), .B(n37268), .Z(n28951) );
  AND U38726 ( .A(\modmult_1/xin[1023] ), .B(n37269), .Z(n37268) );
  IV U38727 ( .A(n37267), .Z(n37269) );
  XOR U38728 ( .A(n37270), .B(g_input[298]), .Z(n37267) );
  NAND U38729 ( .A(n37271), .B(mul_pow), .Z(n37270) );
  XOR U38730 ( .A(g_input[298]), .B(creg[298]), .Z(n37271) );
  XOR U38731 ( .A(n37272), .B(n37273), .Z(n37263) );
  ANDN U38732 ( .A(n37274), .B(n28958), .Z(n37273) );
  XOR U38733 ( .A(n37275), .B(\modmult_1/zin[0][296] ), .Z(n28958) );
  IV U38734 ( .A(n37272), .Z(n37275) );
  XNOR U38735 ( .A(n37272), .B(n28957), .Z(n37274) );
  XOR U38736 ( .A(n37276), .B(n37277), .Z(n28957) );
  AND U38737 ( .A(\modmult_1/xin[1023] ), .B(n37278), .Z(n37277) );
  IV U38738 ( .A(n37276), .Z(n37278) );
  XOR U38739 ( .A(n37279), .B(g_input[297]), .Z(n37276) );
  NAND U38740 ( .A(n37280), .B(mul_pow), .Z(n37279) );
  XOR U38741 ( .A(g_input[297]), .B(creg[297]), .Z(n37280) );
  XOR U38742 ( .A(n37281), .B(n37282), .Z(n37272) );
  ANDN U38743 ( .A(n37283), .B(n28964), .Z(n37282) );
  XOR U38744 ( .A(n37284), .B(\modmult_1/zin[0][295] ), .Z(n28964) );
  IV U38745 ( .A(n37281), .Z(n37284) );
  XNOR U38746 ( .A(n37281), .B(n28963), .Z(n37283) );
  XOR U38747 ( .A(n37285), .B(n37286), .Z(n28963) );
  AND U38748 ( .A(\modmult_1/xin[1023] ), .B(n37287), .Z(n37286) );
  IV U38749 ( .A(n37285), .Z(n37287) );
  XOR U38750 ( .A(n37288), .B(g_input[296]), .Z(n37285) );
  NAND U38751 ( .A(n37289), .B(mul_pow), .Z(n37288) );
  XOR U38752 ( .A(g_input[296]), .B(creg[296]), .Z(n37289) );
  XOR U38753 ( .A(n37290), .B(n37291), .Z(n37281) );
  ANDN U38754 ( .A(n37292), .B(n28970), .Z(n37291) );
  XOR U38755 ( .A(n37293), .B(\modmult_1/zin[0][294] ), .Z(n28970) );
  IV U38756 ( .A(n37290), .Z(n37293) );
  XNOR U38757 ( .A(n37290), .B(n28969), .Z(n37292) );
  XOR U38758 ( .A(n37294), .B(n37295), .Z(n28969) );
  AND U38759 ( .A(\modmult_1/xin[1023] ), .B(n37296), .Z(n37295) );
  IV U38760 ( .A(n37294), .Z(n37296) );
  XOR U38761 ( .A(n37297), .B(g_input[295]), .Z(n37294) );
  NAND U38762 ( .A(n37298), .B(mul_pow), .Z(n37297) );
  XOR U38763 ( .A(g_input[295]), .B(creg[295]), .Z(n37298) );
  XOR U38764 ( .A(n37299), .B(n37300), .Z(n37290) );
  ANDN U38765 ( .A(n37301), .B(n28976), .Z(n37300) );
  XOR U38766 ( .A(n37302), .B(\modmult_1/zin[0][293] ), .Z(n28976) );
  IV U38767 ( .A(n37299), .Z(n37302) );
  XNOR U38768 ( .A(n37299), .B(n28975), .Z(n37301) );
  XOR U38769 ( .A(n37303), .B(n37304), .Z(n28975) );
  AND U38770 ( .A(\modmult_1/xin[1023] ), .B(n37305), .Z(n37304) );
  IV U38771 ( .A(n37303), .Z(n37305) );
  XOR U38772 ( .A(n37306), .B(g_input[294]), .Z(n37303) );
  NAND U38773 ( .A(n37307), .B(mul_pow), .Z(n37306) );
  XOR U38774 ( .A(g_input[294]), .B(creg[294]), .Z(n37307) );
  XOR U38775 ( .A(n37308), .B(n37309), .Z(n37299) );
  ANDN U38776 ( .A(n37310), .B(n28982), .Z(n37309) );
  XOR U38777 ( .A(n37311), .B(\modmult_1/zin[0][292] ), .Z(n28982) );
  IV U38778 ( .A(n37308), .Z(n37311) );
  XNOR U38779 ( .A(n37308), .B(n28981), .Z(n37310) );
  XOR U38780 ( .A(n37312), .B(n37313), .Z(n28981) );
  AND U38781 ( .A(\modmult_1/xin[1023] ), .B(n37314), .Z(n37313) );
  IV U38782 ( .A(n37312), .Z(n37314) );
  XOR U38783 ( .A(n37315), .B(g_input[293]), .Z(n37312) );
  NAND U38784 ( .A(n37316), .B(mul_pow), .Z(n37315) );
  XOR U38785 ( .A(g_input[293]), .B(creg[293]), .Z(n37316) );
  XOR U38786 ( .A(n37317), .B(n37318), .Z(n37308) );
  ANDN U38787 ( .A(n37319), .B(n28988), .Z(n37318) );
  XOR U38788 ( .A(n37320), .B(\modmult_1/zin[0][291] ), .Z(n28988) );
  IV U38789 ( .A(n37317), .Z(n37320) );
  XNOR U38790 ( .A(n37317), .B(n28987), .Z(n37319) );
  XOR U38791 ( .A(n37321), .B(n37322), .Z(n28987) );
  AND U38792 ( .A(\modmult_1/xin[1023] ), .B(n37323), .Z(n37322) );
  IV U38793 ( .A(n37321), .Z(n37323) );
  XOR U38794 ( .A(n37324), .B(g_input[292]), .Z(n37321) );
  NAND U38795 ( .A(n37325), .B(mul_pow), .Z(n37324) );
  XOR U38796 ( .A(g_input[292]), .B(creg[292]), .Z(n37325) );
  XOR U38797 ( .A(n37326), .B(n37327), .Z(n37317) );
  ANDN U38798 ( .A(n37328), .B(n28994), .Z(n37327) );
  XOR U38799 ( .A(n37329), .B(\modmult_1/zin[0][290] ), .Z(n28994) );
  IV U38800 ( .A(n37326), .Z(n37329) );
  XNOR U38801 ( .A(n37326), .B(n28993), .Z(n37328) );
  XOR U38802 ( .A(n37330), .B(n37331), .Z(n28993) );
  AND U38803 ( .A(\modmult_1/xin[1023] ), .B(n37332), .Z(n37331) );
  IV U38804 ( .A(n37330), .Z(n37332) );
  XOR U38805 ( .A(n37333), .B(g_input[291]), .Z(n37330) );
  NAND U38806 ( .A(n37334), .B(mul_pow), .Z(n37333) );
  XOR U38807 ( .A(g_input[291]), .B(creg[291]), .Z(n37334) );
  XOR U38808 ( .A(n37335), .B(n37336), .Z(n37326) );
  ANDN U38809 ( .A(n37337), .B(n29000), .Z(n37336) );
  XOR U38810 ( .A(n37338), .B(\modmult_1/zin[0][289] ), .Z(n29000) );
  IV U38811 ( .A(n37335), .Z(n37338) );
  XNOR U38812 ( .A(n37335), .B(n28999), .Z(n37337) );
  XOR U38813 ( .A(n37339), .B(n37340), .Z(n28999) );
  AND U38814 ( .A(\modmult_1/xin[1023] ), .B(n37341), .Z(n37340) );
  IV U38815 ( .A(n37339), .Z(n37341) );
  XOR U38816 ( .A(n37342), .B(g_input[290]), .Z(n37339) );
  NAND U38817 ( .A(n37343), .B(mul_pow), .Z(n37342) );
  XOR U38818 ( .A(g_input[290]), .B(creg[290]), .Z(n37343) );
  XOR U38819 ( .A(n37344), .B(n37345), .Z(n37335) );
  ANDN U38820 ( .A(n37346), .B(n29006), .Z(n37345) );
  XOR U38821 ( .A(n37347), .B(\modmult_1/zin[0][288] ), .Z(n29006) );
  IV U38822 ( .A(n37344), .Z(n37347) );
  XNOR U38823 ( .A(n37344), .B(n29005), .Z(n37346) );
  XOR U38824 ( .A(n37348), .B(n37349), .Z(n29005) );
  AND U38825 ( .A(\modmult_1/xin[1023] ), .B(n37350), .Z(n37349) );
  IV U38826 ( .A(n37348), .Z(n37350) );
  XOR U38827 ( .A(n37351), .B(g_input[289]), .Z(n37348) );
  NAND U38828 ( .A(n37352), .B(mul_pow), .Z(n37351) );
  XOR U38829 ( .A(g_input[289]), .B(creg[289]), .Z(n37352) );
  XOR U38830 ( .A(n37353), .B(n37354), .Z(n37344) );
  ANDN U38831 ( .A(n37355), .B(n29012), .Z(n37354) );
  XOR U38832 ( .A(n37356), .B(\modmult_1/zin[0][287] ), .Z(n29012) );
  IV U38833 ( .A(n37353), .Z(n37356) );
  XNOR U38834 ( .A(n37353), .B(n29011), .Z(n37355) );
  XOR U38835 ( .A(n37357), .B(n37358), .Z(n29011) );
  AND U38836 ( .A(\modmult_1/xin[1023] ), .B(n37359), .Z(n37358) );
  IV U38837 ( .A(n37357), .Z(n37359) );
  XOR U38838 ( .A(n37360), .B(g_input[288]), .Z(n37357) );
  NAND U38839 ( .A(n37361), .B(mul_pow), .Z(n37360) );
  XOR U38840 ( .A(g_input[288]), .B(creg[288]), .Z(n37361) );
  XOR U38841 ( .A(n37362), .B(n37363), .Z(n37353) );
  ANDN U38842 ( .A(n37364), .B(n29018), .Z(n37363) );
  XOR U38843 ( .A(n37365), .B(\modmult_1/zin[0][286] ), .Z(n29018) );
  IV U38844 ( .A(n37362), .Z(n37365) );
  XNOR U38845 ( .A(n37362), .B(n29017), .Z(n37364) );
  XOR U38846 ( .A(n37366), .B(n37367), .Z(n29017) );
  AND U38847 ( .A(\modmult_1/xin[1023] ), .B(n37368), .Z(n37367) );
  IV U38848 ( .A(n37366), .Z(n37368) );
  XOR U38849 ( .A(n37369), .B(g_input[287]), .Z(n37366) );
  NAND U38850 ( .A(n37370), .B(mul_pow), .Z(n37369) );
  XOR U38851 ( .A(g_input[287]), .B(creg[287]), .Z(n37370) );
  XOR U38852 ( .A(n37371), .B(n37372), .Z(n37362) );
  ANDN U38853 ( .A(n37373), .B(n29024), .Z(n37372) );
  XOR U38854 ( .A(n37374), .B(\modmult_1/zin[0][285] ), .Z(n29024) );
  IV U38855 ( .A(n37371), .Z(n37374) );
  XNOR U38856 ( .A(n37371), .B(n29023), .Z(n37373) );
  XOR U38857 ( .A(n37375), .B(n37376), .Z(n29023) );
  AND U38858 ( .A(\modmult_1/xin[1023] ), .B(n37377), .Z(n37376) );
  IV U38859 ( .A(n37375), .Z(n37377) );
  XOR U38860 ( .A(n37378), .B(g_input[286]), .Z(n37375) );
  NAND U38861 ( .A(n37379), .B(mul_pow), .Z(n37378) );
  XOR U38862 ( .A(g_input[286]), .B(creg[286]), .Z(n37379) );
  XOR U38863 ( .A(n37380), .B(n37381), .Z(n37371) );
  ANDN U38864 ( .A(n37382), .B(n29030), .Z(n37381) );
  XOR U38865 ( .A(n37383), .B(\modmult_1/zin[0][284] ), .Z(n29030) );
  IV U38866 ( .A(n37380), .Z(n37383) );
  XNOR U38867 ( .A(n37380), .B(n29029), .Z(n37382) );
  XOR U38868 ( .A(n37384), .B(n37385), .Z(n29029) );
  AND U38869 ( .A(\modmult_1/xin[1023] ), .B(n37386), .Z(n37385) );
  IV U38870 ( .A(n37384), .Z(n37386) );
  XOR U38871 ( .A(n37387), .B(g_input[285]), .Z(n37384) );
  NAND U38872 ( .A(n37388), .B(mul_pow), .Z(n37387) );
  XOR U38873 ( .A(g_input[285]), .B(creg[285]), .Z(n37388) );
  XOR U38874 ( .A(n37389), .B(n37390), .Z(n37380) );
  ANDN U38875 ( .A(n37391), .B(n29036), .Z(n37390) );
  XOR U38876 ( .A(n37392), .B(\modmult_1/zin[0][283] ), .Z(n29036) );
  IV U38877 ( .A(n37389), .Z(n37392) );
  XNOR U38878 ( .A(n37389), .B(n29035), .Z(n37391) );
  XOR U38879 ( .A(n37393), .B(n37394), .Z(n29035) );
  AND U38880 ( .A(\modmult_1/xin[1023] ), .B(n37395), .Z(n37394) );
  IV U38881 ( .A(n37393), .Z(n37395) );
  XOR U38882 ( .A(n37396), .B(g_input[284]), .Z(n37393) );
  NAND U38883 ( .A(n37397), .B(mul_pow), .Z(n37396) );
  XOR U38884 ( .A(g_input[284]), .B(creg[284]), .Z(n37397) );
  XOR U38885 ( .A(n37398), .B(n37399), .Z(n37389) );
  ANDN U38886 ( .A(n37400), .B(n29042), .Z(n37399) );
  XOR U38887 ( .A(n37401), .B(\modmult_1/zin[0][282] ), .Z(n29042) );
  IV U38888 ( .A(n37398), .Z(n37401) );
  XNOR U38889 ( .A(n37398), .B(n29041), .Z(n37400) );
  XOR U38890 ( .A(n37402), .B(n37403), .Z(n29041) );
  AND U38891 ( .A(\modmult_1/xin[1023] ), .B(n37404), .Z(n37403) );
  IV U38892 ( .A(n37402), .Z(n37404) );
  XOR U38893 ( .A(n37405), .B(g_input[283]), .Z(n37402) );
  NAND U38894 ( .A(n37406), .B(mul_pow), .Z(n37405) );
  XOR U38895 ( .A(g_input[283]), .B(creg[283]), .Z(n37406) );
  XOR U38896 ( .A(n37407), .B(n37408), .Z(n37398) );
  ANDN U38897 ( .A(n37409), .B(n29048), .Z(n37408) );
  XOR U38898 ( .A(n37410), .B(\modmult_1/zin[0][281] ), .Z(n29048) );
  IV U38899 ( .A(n37407), .Z(n37410) );
  XNOR U38900 ( .A(n37407), .B(n29047), .Z(n37409) );
  XOR U38901 ( .A(n37411), .B(n37412), .Z(n29047) );
  AND U38902 ( .A(\modmult_1/xin[1023] ), .B(n37413), .Z(n37412) );
  IV U38903 ( .A(n37411), .Z(n37413) );
  XOR U38904 ( .A(n37414), .B(g_input[282]), .Z(n37411) );
  NAND U38905 ( .A(n37415), .B(mul_pow), .Z(n37414) );
  XOR U38906 ( .A(g_input[282]), .B(creg[282]), .Z(n37415) );
  XOR U38907 ( .A(n37416), .B(n37417), .Z(n37407) );
  ANDN U38908 ( .A(n37418), .B(n29054), .Z(n37417) );
  XOR U38909 ( .A(n37419), .B(\modmult_1/zin[0][280] ), .Z(n29054) );
  IV U38910 ( .A(n37416), .Z(n37419) );
  XNOR U38911 ( .A(n37416), .B(n29053), .Z(n37418) );
  XOR U38912 ( .A(n37420), .B(n37421), .Z(n29053) );
  AND U38913 ( .A(\modmult_1/xin[1023] ), .B(n37422), .Z(n37421) );
  IV U38914 ( .A(n37420), .Z(n37422) );
  XOR U38915 ( .A(n37423), .B(g_input[281]), .Z(n37420) );
  NAND U38916 ( .A(n37424), .B(mul_pow), .Z(n37423) );
  XOR U38917 ( .A(g_input[281]), .B(creg[281]), .Z(n37424) );
  XOR U38918 ( .A(n37425), .B(n37426), .Z(n37416) );
  ANDN U38919 ( .A(n37427), .B(n29060), .Z(n37426) );
  XOR U38920 ( .A(n37428), .B(\modmult_1/zin[0][279] ), .Z(n29060) );
  IV U38921 ( .A(n37425), .Z(n37428) );
  XNOR U38922 ( .A(n37425), .B(n29059), .Z(n37427) );
  XOR U38923 ( .A(n37429), .B(n37430), .Z(n29059) );
  AND U38924 ( .A(\modmult_1/xin[1023] ), .B(n37431), .Z(n37430) );
  IV U38925 ( .A(n37429), .Z(n37431) );
  XOR U38926 ( .A(n37432), .B(g_input[280]), .Z(n37429) );
  NAND U38927 ( .A(n37433), .B(mul_pow), .Z(n37432) );
  XOR U38928 ( .A(g_input[280]), .B(creg[280]), .Z(n37433) );
  XOR U38929 ( .A(n37434), .B(n37435), .Z(n37425) );
  ANDN U38930 ( .A(n37436), .B(n29066), .Z(n37435) );
  XOR U38931 ( .A(n37437), .B(\modmult_1/zin[0][278] ), .Z(n29066) );
  IV U38932 ( .A(n37434), .Z(n37437) );
  XNOR U38933 ( .A(n37434), .B(n29065), .Z(n37436) );
  XOR U38934 ( .A(n37438), .B(n37439), .Z(n29065) );
  AND U38935 ( .A(\modmult_1/xin[1023] ), .B(n37440), .Z(n37439) );
  IV U38936 ( .A(n37438), .Z(n37440) );
  XOR U38937 ( .A(n37441), .B(g_input[279]), .Z(n37438) );
  NAND U38938 ( .A(n37442), .B(mul_pow), .Z(n37441) );
  XOR U38939 ( .A(g_input[279]), .B(creg[279]), .Z(n37442) );
  XOR U38940 ( .A(n37443), .B(n37444), .Z(n37434) );
  ANDN U38941 ( .A(n37445), .B(n29072), .Z(n37444) );
  XOR U38942 ( .A(n37446), .B(\modmult_1/zin[0][277] ), .Z(n29072) );
  IV U38943 ( .A(n37443), .Z(n37446) );
  XNOR U38944 ( .A(n37443), .B(n29071), .Z(n37445) );
  XOR U38945 ( .A(n37447), .B(n37448), .Z(n29071) );
  AND U38946 ( .A(\modmult_1/xin[1023] ), .B(n37449), .Z(n37448) );
  IV U38947 ( .A(n37447), .Z(n37449) );
  XOR U38948 ( .A(n37450), .B(g_input[278]), .Z(n37447) );
  NAND U38949 ( .A(n37451), .B(mul_pow), .Z(n37450) );
  XOR U38950 ( .A(g_input[278]), .B(creg[278]), .Z(n37451) );
  XOR U38951 ( .A(n37452), .B(n37453), .Z(n37443) );
  ANDN U38952 ( .A(n37454), .B(n29078), .Z(n37453) );
  XOR U38953 ( .A(n37455), .B(\modmult_1/zin[0][276] ), .Z(n29078) );
  IV U38954 ( .A(n37452), .Z(n37455) );
  XNOR U38955 ( .A(n37452), .B(n29077), .Z(n37454) );
  XOR U38956 ( .A(n37456), .B(n37457), .Z(n29077) );
  AND U38957 ( .A(\modmult_1/xin[1023] ), .B(n37458), .Z(n37457) );
  IV U38958 ( .A(n37456), .Z(n37458) );
  XOR U38959 ( .A(n37459), .B(g_input[277]), .Z(n37456) );
  NAND U38960 ( .A(n37460), .B(mul_pow), .Z(n37459) );
  XOR U38961 ( .A(g_input[277]), .B(creg[277]), .Z(n37460) );
  XOR U38962 ( .A(n37461), .B(n37462), .Z(n37452) );
  ANDN U38963 ( .A(n37463), .B(n29084), .Z(n37462) );
  XOR U38964 ( .A(n37464), .B(\modmult_1/zin[0][275] ), .Z(n29084) );
  IV U38965 ( .A(n37461), .Z(n37464) );
  XNOR U38966 ( .A(n37461), .B(n29083), .Z(n37463) );
  XOR U38967 ( .A(n37465), .B(n37466), .Z(n29083) );
  AND U38968 ( .A(\modmult_1/xin[1023] ), .B(n37467), .Z(n37466) );
  IV U38969 ( .A(n37465), .Z(n37467) );
  XOR U38970 ( .A(n37468), .B(g_input[276]), .Z(n37465) );
  NAND U38971 ( .A(n37469), .B(mul_pow), .Z(n37468) );
  XOR U38972 ( .A(g_input[276]), .B(creg[276]), .Z(n37469) );
  XOR U38973 ( .A(n37470), .B(n37471), .Z(n37461) );
  ANDN U38974 ( .A(n37472), .B(n29090), .Z(n37471) );
  XOR U38975 ( .A(n37473), .B(\modmult_1/zin[0][274] ), .Z(n29090) );
  IV U38976 ( .A(n37470), .Z(n37473) );
  XNOR U38977 ( .A(n37470), .B(n29089), .Z(n37472) );
  XOR U38978 ( .A(n37474), .B(n37475), .Z(n29089) );
  AND U38979 ( .A(\modmult_1/xin[1023] ), .B(n37476), .Z(n37475) );
  IV U38980 ( .A(n37474), .Z(n37476) );
  XOR U38981 ( .A(n37477), .B(g_input[275]), .Z(n37474) );
  NAND U38982 ( .A(n37478), .B(mul_pow), .Z(n37477) );
  XOR U38983 ( .A(g_input[275]), .B(creg[275]), .Z(n37478) );
  XOR U38984 ( .A(n37479), .B(n37480), .Z(n37470) );
  ANDN U38985 ( .A(n37481), .B(n29096), .Z(n37480) );
  XOR U38986 ( .A(n37482), .B(\modmult_1/zin[0][273] ), .Z(n29096) );
  IV U38987 ( .A(n37479), .Z(n37482) );
  XNOR U38988 ( .A(n37479), .B(n29095), .Z(n37481) );
  XOR U38989 ( .A(n37483), .B(n37484), .Z(n29095) );
  AND U38990 ( .A(\modmult_1/xin[1023] ), .B(n37485), .Z(n37484) );
  IV U38991 ( .A(n37483), .Z(n37485) );
  XOR U38992 ( .A(n37486), .B(g_input[274]), .Z(n37483) );
  NAND U38993 ( .A(n37487), .B(mul_pow), .Z(n37486) );
  XOR U38994 ( .A(g_input[274]), .B(creg[274]), .Z(n37487) );
  XOR U38995 ( .A(n37488), .B(n37489), .Z(n37479) );
  ANDN U38996 ( .A(n37490), .B(n29102), .Z(n37489) );
  XOR U38997 ( .A(n37491), .B(\modmult_1/zin[0][272] ), .Z(n29102) );
  IV U38998 ( .A(n37488), .Z(n37491) );
  XNOR U38999 ( .A(n37488), .B(n29101), .Z(n37490) );
  XOR U39000 ( .A(n37492), .B(n37493), .Z(n29101) );
  AND U39001 ( .A(\modmult_1/xin[1023] ), .B(n37494), .Z(n37493) );
  IV U39002 ( .A(n37492), .Z(n37494) );
  XOR U39003 ( .A(n37495), .B(g_input[273]), .Z(n37492) );
  NAND U39004 ( .A(n37496), .B(mul_pow), .Z(n37495) );
  XOR U39005 ( .A(g_input[273]), .B(creg[273]), .Z(n37496) );
  XOR U39006 ( .A(n37497), .B(n37498), .Z(n37488) );
  ANDN U39007 ( .A(n37499), .B(n29108), .Z(n37498) );
  XOR U39008 ( .A(n37500), .B(\modmult_1/zin[0][271] ), .Z(n29108) );
  IV U39009 ( .A(n37497), .Z(n37500) );
  XNOR U39010 ( .A(n37497), .B(n29107), .Z(n37499) );
  XOR U39011 ( .A(n37501), .B(n37502), .Z(n29107) );
  AND U39012 ( .A(\modmult_1/xin[1023] ), .B(n37503), .Z(n37502) );
  IV U39013 ( .A(n37501), .Z(n37503) );
  XOR U39014 ( .A(n37504), .B(g_input[272]), .Z(n37501) );
  NAND U39015 ( .A(n37505), .B(mul_pow), .Z(n37504) );
  XOR U39016 ( .A(g_input[272]), .B(creg[272]), .Z(n37505) );
  XOR U39017 ( .A(n37506), .B(n37507), .Z(n37497) );
  ANDN U39018 ( .A(n37508), .B(n29114), .Z(n37507) );
  XOR U39019 ( .A(n37509), .B(\modmult_1/zin[0][270] ), .Z(n29114) );
  IV U39020 ( .A(n37506), .Z(n37509) );
  XNOR U39021 ( .A(n37506), .B(n29113), .Z(n37508) );
  XOR U39022 ( .A(n37510), .B(n37511), .Z(n29113) );
  AND U39023 ( .A(\modmult_1/xin[1023] ), .B(n37512), .Z(n37511) );
  IV U39024 ( .A(n37510), .Z(n37512) );
  XOR U39025 ( .A(n37513), .B(g_input[271]), .Z(n37510) );
  NAND U39026 ( .A(n37514), .B(mul_pow), .Z(n37513) );
  XOR U39027 ( .A(g_input[271]), .B(creg[271]), .Z(n37514) );
  XOR U39028 ( .A(n37515), .B(n37516), .Z(n37506) );
  ANDN U39029 ( .A(n37517), .B(n29120), .Z(n37516) );
  XOR U39030 ( .A(n37518), .B(\modmult_1/zin[0][269] ), .Z(n29120) );
  IV U39031 ( .A(n37515), .Z(n37518) );
  XNOR U39032 ( .A(n37515), .B(n29119), .Z(n37517) );
  XOR U39033 ( .A(n37519), .B(n37520), .Z(n29119) );
  AND U39034 ( .A(\modmult_1/xin[1023] ), .B(n37521), .Z(n37520) );
  IV U39035 ( .A(n37519), .Z(n37521) );
  XOR U39036 ( .A(n37522), .B(g_input[270]), .Z(n37519) );
  NAND U39037 ( .A(n37523), .B(mul_pow), .Z(n37522) );
  XOR U39038 ( .A(g_input[270]), .B(creg[270]), .Z(n37523) );
  XOR U39039 ( .A(n37524), .B(n37525), .Z(n37515) );
  ANDN U39040 ( .A(n37526), .B(n29126), .Z(n37525) );
  XOR U39041 ( .A(n37527), .B(\modmult_1/zin[0][268] ), .Z(n29126) );
  IV U39042 ( .A(n37524), .Z(n37527) );
  XNOR U39043 ( .A(n37524), .B(n29125), .Z(n37526) );
  XOR U39044 ( .A(n37528), .B(n37529), .Z(n29125) );
  AND U39045 ( .A(\modmult_1/xin[1023] ), .B(n37530), .Z(n37529) );
  IV U39046 ( .A(n37528), .Z(n37530) );
  XOR U39047 ( .A(n37531), .B(g_input[269]), .Z(n37528) );
  NAND U39048 ( .A(n37532), .B(mul_pow), .Z(n37531) );
  XOR U39049 ( .A(g_input[269]), .B(creg[269]), .Z(n37532) );
  XOR U39050 ( .A(n37533), .B(n37534), .Z(n37524) );
  ANDN U39051 ( .A(n37535), .B(n29132), .Z(n37534) );
  XOR U39052 ( .A(n37536), .B(\modmult_1/zin[0][267] ), .Z(n29132) );
  IV U39053 ( .A(n37533), .Z(n37536) );
  XNOR U39054 ( .A(n37533), .B(n29131), .Z(n37535) );
  XOR U39055 ( .A(n37537), .B(n37538), .Z(n29131) );
  AND U39056 ( .A(\modmult_1/xin[1023] ), .B(n37539), .Z(n37538) );
  IV U39057 ( .A(n37537), .Z(n37539) );
  XOR U39058 ( .A(n37540), .B(g_input[268]), .Z(n37537) );
  NAND U39059 ( .A(n37541), .B(mul_pow), .Z(n37540) );
  XOR U39060 ( .A(g_input[268]), .B(creg[268]), .Z(n37541) );
  XOR U39061 ( .A(n37542), .B(n37543), .Z(n37533) );
  ANDN U39062 ( .A(n37544), .B(n29138), .Z(n37543) );
  XOR U39063 ( .A(n37545), .B(\modmult_1/zin[0][266] ), .Z(n29138) );
  IV U39064 ( .A(n37542), .Z(n37545) );
  XNOR U39065 ( .A(n37542), .B(n29137), .Z(n37544) );
  XOR U39066 ( .A(n37546), .B(n37547), .Z(n29137) );
  AND U39067 ( .A(\modmult_1/xin[1023] ), .B(n37548), .Z(n37547) );
  IV U39068 ( .A(n37546), .Z(n37548) );
  XOR U39069 ( .A(n37549), .B(g_input[267]), .Z(n37546) );
  NAND U39070 ( .A(n37550), .B(mul_pow), .Z(n37549) );
  XOR U39071 ( .A(g_input[267]), .B(creg[267]), .Z(n37550) );
  XOR U39072 ( .A(n37551), .B(n37552), .Z(n37542) );
  ANDN U39073 ( .A(n37553), .B(n29144), .Z(n37552) );
  XOR U39074 ( .A(n37554), .B(\modmult_1/zin[0][265] ), .Z(n29144) );
  IV U39075 ( .A(n37551), .Z(n37554) );
  XNOR U39076 ( .A(n37551), .B(n29143), .Z(n37553) );
  XOR U39077 ( .A(n37555), .B(n37556), .Z(n29143) );
  AND U39078 ( .A(\modmult_1/xin[1023] ), .B(n37557), .Z(n37556) );
  IV U39079 ( .A(n37555), .Z(n37557) );
  XOR U39080 ( .A(n37558), .B(g_input[266]), .Z(n37555) );
  NAND U39081 ( .A(n37559), .B(mul_pow), .Z(n37558) );
  XOR U39082 ( .A(g_input[266]), .B(creg[266]), .Z(n37559) );
  XOR U39083 ( .A(n37560), .B(n37561), .Z(n37551) );
  ANDN U39084 ( .A(n37562), .B(n29150), .Z(n37561) );
  XOR U39085 ( .A(n37563), .B(\modmult_1/zin[0][264] ), .Z(n29150) );
  IV U39086 ( .A(n37560), .Z(n37563) );
  XNOR U39087 ( .A(n37560), .B(n29149), .Z(n37562) );
  XOR U39088 ( .A(n37564), .B(n37565), .Z(n29149) );
  AND U39089 ( .A(\modmult_1/xin[1023] ), .B(n37566), .Z(n37565) );
  IV U39090 ( .A(n37564), .Z(n37566) );
  XOR U39091 ( .A(n37567), .B(g_input[265]), .Z(n37564) );
  NAND U39092 ( .A(n37568), .B(mul_pow), .Z(n37567) );
  XOR U39093 ( .A(g_input[265]), .B(creg[265]), .Z(n37568) );
  XOR U39094 ( .A(n37569), .B(n37570), .Z(n37560) );
  ANDN U39095 ( .A(n37571), .B(n29156), .Z(n37570) );
  XOR U39096 ( .A(n37572), .B(\modmult_1/zin[0][263] ), .Z(n29156) );
  IV U39097 ( .A(n37569), .Z(n37572) );
  XNOR U39098 ( .A(n37569), .B(n29155), .Z(n37571) );
  XOR U39099 ( .A(n37573), .B(n37574), .Z(n29155) );
  AND U39100 ( .A(\modmult_1/xin[1023] ), .B(n37575), .Z(n37574) );
  IV U39101 ( .A(n37573), .Z(n37575) );
  XOR U39102 ( .A(n37576), .B(g_input[264]), .Z(n37573) );
  NAND U39103 ( .A(n37577), .B(mul_pow), .Z(n37576) );
  XOR U39104 ( .A(g_input[264]), .B(creg[264]), .Z(n37577) );
  XOR U39105 ( .A(n37578), .B(n37579), .Z(n37569) );
  ANDN U39106 ( .A(n37580), .B(n29162), .Z(n37579) );
  XOR U39107 ( .A(n37581), .B(\modmult_1/zin[0][262] ), .Z(n29162) );
  IV U39108 ( .A(n37578), .Z(n37581) );
  XNOR U39109 ( .A(n37578), .B(n29161), .Z(n37580) );
  XOR U39110 ( .A(n37582), .B(n37583), .Z(n29161) );
  AND U39111 ( .A(\modmult_1/xin[1023] ), .B(n37584), .Z(n37583) );
  IV U39112 ( .A(n37582), .Z(n37584) );
  XOR U39113 ( .A(n37585), .B(g_input[263]), .Z(n37582) );
  NAND U39114 ( .A(n37586), .B(mul_pow), .Z(n37585) );
  XOR U39115 ( .A(g_input[263]), .B(creg[263]), .Z(n37586) );
  XOR U39116 ( .A(n37587), .B(n37588), .Z(n37578) );
  ANDN U39117 ( .A(n37589), .B(n29168), .Z(n37588) );
  XOR U39118 ( .A(n37590), .B(\modmult_1/zin[0][261] ), .Z(n29168) );
  IV U39119 ( .A(n37587), .Z(n37590) );
  XNOR U39120 ( .A(n37587), .B(n29167), .Z(n37589) );
  XOR U39121 ( .A(n37591), .B(n37592), .Z(n29167) );
  AND U39122 ( .A(\modmult_1/xin[1023] ), .B(n37593), .Z(n37592) );
  IV U39123 ( .A(n37591), .Z(n37593) );
  XOR U39124 ( .A(n37594), .B(g_input[262]), .Z(n37591) );
  NAND U39125 ( .A(n37595), .B(mul_pow), .Z(n37594) );
  XOR U39126 ( .A(g_input[262]), .B(creg[262]), .Z(n37595) );
  XOR U39127 ( .A(n37596), .B(n37597), .Z(n37587) );
  ANDN U39128 ( .A(n37598), .B(n29174), .Z(n37597) );
  XOR U39129 ( .A(n37599), .B(\modmult_1/zin[0][260] ), .Z(n29174) );
  IV U39130 ( .A(n37596), .Z(n37599) );
  XNOR U39131 ( .A(n37596), .B(n29173), .Z(n37598) );
  XOR U39132 ( .A(n37600), .B(n37601), .Z(n29173) );
  AND U39133 ( .A(\modmult_1/xin[1023] ), .B(n37602), .Z(n37601) );
  IV U39134 ( .A(n37600), .Z(n37602) );
  XOR U39135 ( .A(n37603), .B(g_input[261]), .Z(n37600) );
  NAND U39136 ( .A(n37604), .B(mul_pow), .Z(n37603) );
  XOR U39137 ( .A(g_input[261]), .B(creg[261]), .Z(n37604) );
  XOR U39138 ( .A(n37605), .B(n37606), .Z(n37596) );
  ANDN U39139 ( .A(n37607), .B(n29180), .Z(n37606) );
  XOR U39140 ( .A(n37608), .B(\modmult_1/zin[0][259] ), .Z(n29180) );
  IV U39141 ( .A(n37605), .Z(n37608) );
  XNOR U39142 ( .A(n37605), .B(n29179), .Z(n37607) );
  XOR U39143 ( .A(n37609), .B(n37610), .Z(n29179) );
  AND U39144 ( .A(\modmult_1/xin[1023] ), .B(n37611), .Z(n37610) );
  IV U39145 ( .A(n37609), .Z(n37611) );
  XOR U39146 ( .A(n37612), .B(g_input[260]), .Z(n37609) );
  NAND U39147 ( .A(n37613), .B(mul_pow), .Z(n37612) );
  XOR U39148 ( .A(g_input[260]), .B(creg[260]), .Z(n37613) );
  XOR U39149 ( .A(n37614), .B(n37615), .Z(n37605) );
  ANDN U39150 ( .A(n37616), .B(n29186), .Z(n37615) );
  XOR U39151 ( .A(n37617), .B(\modmult_1/zin[0][258] ), .Z(n29186) );
  IV U39152 ( .A(n37614), .Z(n37617) );
  XNOR U39153 ( .A(n37614), .B(n29185), .Z(n37616) );
  XOR U39154 ( .A(n37618), .B(n37619), .Z(n29185) );
  AND U39155 ( .A(\modmult_1/xin[1023] ), .B(n37620), .Z(n37619) );
  IV U39156 ( .A(n37618), .Z(n37620) );
  XOR U39157 ( .A(n37621), .B(g_input[259]), .Z(n37618) );
  NAND U39158 ( .A(n37622), .B(mul_pow), .Z(n37621) );
  XOR U39159 ( .A(g_input[259]), .B(creg[259]), .Z(n37622) );
  XOR U39160 ( .A(n37623), .B(n37624), .Z(n37614) );
  ANDN U39161 ( .A(n37625), .B(n29192), .Z(n37624) );
  XOR U39162 ( .A(n37626), .B(\modmult_1/zin[0][257] ), .Z(n29192) );
  IV U39163 ( .A(n37623), .Z(n37626) );
  XNOR U39164 ( .A(n37623), .B(n29191), .Z(n37625) );
  XOR U39165 ( .A(n37627), .B(n37628), .Z(n29191) );
  AND U39166 ( .A(\modmult_1/xin[1023] ), .B(n37629), .Z(n37628) );
  IV U39167 ( .A(n37627), .Z(n37629) );
  XOR U39168 ( .A(n37630), .B(g_input[258]), .Z(n37627) );
  NAND U39169 ( .A(n37631), .B(mul_pow), .Z(n37630) );
  XOR U39170 ( .A(g_input[258]), .B(creg[258]), .Z(n37631) );
  XOR U39171 ( .A(n37632), .B(n37633), .Z(n37623) );
  ANDN U39172 ( .A(n37634), .B(n29198), .Z(n37633) );
  XOR U39173 ( .A(n37635), .B(\modmult_1/zin[0][256] ), .Z(n29198) );
  IV U39174 ( .A(n37632), .Z(n37635) );
  XNOR U39175 ( .A(n37632), .B(n29197), .Z(n37634) );
  XOR U39176 ( .A(n37636), .B(n37637), .Z(n29197) );
  AND U39177 ( .A(\modmult_1/xin[1023] ), .B(n37638), .Z(n37637) );
  IV U39178 ( .A(n37636), .Z(n37638) );
  XOR U39179 ( .A(n37639), .B(g_input[257]), .Z(n37636) );
  NAND U39180 ( .A(n37640), .B(mul_pow), .Z(n37639) );
  XOR U39181 ( .A(g_input[257]), .B(creg[257]), .Z(n37640) );
  XOR U39182 ( .A(n37641), .B(n37642), .Z(n37632) );
  ANDN U39183 ( .A(n37643), .B(n29204), .Z(n37642) );
  XOR U39184 ( .A(n37644), .B(\modmult_1/zin[0][255] ), .Z(n29204) );
  IV U39185 ( .A(n37641), .Z(n37644) );
  XNOR U39186 ( .A(n37641), .B(n29203), .Z(n37643) );
  XOR U39187 ( .A(n37645), .B(n37646), .Z(n29203) );
  AND U39188 ( .A(\modmult_1/xin[1023] ), .B(n37647), .Z(n37646) );
  IV U39189 ( .A(n37645), .Z(n37647) );
  XOR U39190 ( .A(n37648), .B(g_input[256]), .Z(n37645) );
  NAND U39191 ( .A(n37649), .B(mul_pow), .Z(n37648) );
  XOR U39192 ( .A(g_input[256]), .B(creg[256]), .Z(n37649) );
  XOR U39193 ( .A(n37650), .B(n37651), .Z(n37641) );
  ANDN U39194 ( .A(n37652), .B(n29210), .Z(n37651) );
  XOR U39195 ( .A(n37653), .B(\modmult_1/zin[0][254] ), .Z(n29210) );
  IV U39196 ( .A(n37650), .Z(n37653) );
  XNOR U39197 ( .A(n37650), .B(n29209), .Z(n37652) );
  XOR U39198 ( .A(n37654), .B(n37655), .Z(n29209) );
  AND U39199 ( .A(\modmult_1/xin[1023] ), .B(n37656), .Z(n37655) );
  IV U39200 ( .A(n37654), .Z(n37656) );
  XOR U39201 ( .A(n37657), .B(g_input[255]), .Z(n37654) );
  NAND U39202 ( .A(n37658), .B(mul_pow), .Z(n37657) );
  XOR U39203 ( .A(g_input[255]), .B(creg[255]), .Z(n37658) );
  XOR U39204 ( .A(n37659), .B(n37660), .Z(n37650) );
  ANDN U39205 ( .A(n37661), .B(n29216), .Z(n37660) );
  XOR U39206 ( .A(n37662), .B(\modmult_1/zin[0][253] ), .Z(n29216) );
  IV U39207 ( .A(n37659), .Z(n37662) );
  XNOR U39208 ( .A(n37659), .B(n29215), .Z(n37661) );
  XOR U39209 ( .A(n37663), .B(n37664), .Z(n29215) );
  AND U39210 ( .A(\modmult_1/xin[1023] ), .B(n37665), .Z(n37664) );
  IV U39211 ( .A(n37663), .Z(n37665) );
  XOR U39212 ( .A(n37666), .B(g_input[254]), .Z(n37663) );
  NAND U39213 ( .A(n37667), .B(mul_pow), .Z(n37666) );
  XOR U39214 ( .A(g_input[254]), .B(creg[254]), .Z(n37667) );
  XOR U39215 ( .A(n37668), .B(n37669), .Z(n37659) );
  ANDN U39216 ( .A(n37670), .B(n29222), .Z(n37669) );
  XOR U39217 ( .A(n37671), .B(\modmult_1/zin[0][252] ), .Z(n29222) );
  IV U39218 ( .A(n37668), .Z(n37671) );
  XNOR U39219 ( .A(n37668), .B(n29221), .Z(n37670) );
  XOR U39220 ( .A(n37672), .B(n37673), .Z(n29221) );
  AND U39221 ( .A(\modmult_1/xin[1023] ), .B(n37674), .Z(n37673) );
  IV U39222 ( .A(n37672), .Z(n37674) );
  XOR U39223 ( .A(n37675), .B(g_input[253]), .Z(n37672) );
  NAND U39224 ( .A(n37676), .B(mul_pow), .Z(n37675) );
  XOR U39225 ( .A(g_input[253]), .B(creg[253]), .Z(n37676) );
  XOR U39226 ( .A(n37677), .B(n37678), .Z(n37668) );
  ANDN U39227 ( .A(n37679), .B(n29228), .Z(n37678) );
  XOR U39228 ( .A(n37680), .B(\modmult_1/zin[0][251] ), .Z(n29228) );
  IV U39229 ( .A(n37677), .Z(n37680) );
  XNOR U39230 ( .A(n37677), .B(n29227), .Z(n37679) );
  XOR U39231 ( .A(n37681), .B(n37682), .Z(n29227) );
  AND U39232 ( .A(\modmult_1/xin[1023] ), .B(n37683), .Z(n37682) );
  IV U39233 ( .A(n37681), .Z(n37683) );
  XOR U39234 ( .A(n37684), .B(g_input[252]), .Z(n37681) );
  NAND U39235 ( .A(n37685), .B(mul_pow), .Z(n37684) );
  XOR U39236 ( .A(g_input[252]), .B(creg[252]), .Z(n37685) );
  XOR U39237 ( .A(n37686), .B(n37687), .Z(n37677) );
  ANDN U39238 ( .A(n37688), .B(n29234), .Z(n37687) );
  XOR U39239 ( .A(n37689), .B(\modmult_1/zin[0][250] ), .Z(n29234) );
  IV U39240 ( .A(n37686), .Z(n37689) );
  XNOR U39241 ( .A(n37686), .B(n29233), .Z(n37688) );
  XOR U39242 ( .A(n37690), .B(n37691), .Z(n29233) );
  AND U39243 ( .A(\modmult_1/xin[1023] ), .B(n37692), .Z(n37691) );
  IV U39244 ( .A(n37690), .Z(n37692) );
  XOR U39245 ( .A(n37693), .B(g_input[251]), .Z(n37690) );
  NAND U39246 ( .A(n37694), .B(mul_pow), .Z(n37693) );
  XOR U39247 ( .A(g_input[251]), .B(creg[251]), .Z(n37694) );
  XOR U39248 ( .A(n37695), .B(n37696), .Z(n37686) );
  ANDN U39249 ( .A(n37697), .B(n29240), .Z(n37696) );
  XOR U39250 ( .A(n37698), .B(\modmult_1/zin[0][249] ), .Z(n29240) );
  IV U39251 ( .A(n37695), .Z(n37698) );
  XNOR U39252 ( .A(n37695), .B(n29239), .Z(n37697) );
  XOR U39253 ( .A(n37699), .B(n37700), .Z(n29239) );
  AND U39254 ( .A(\modmult_1/xin[1023] ), .B(n37701), .Z(n37700) );
  IV U39255 ( .A(n37699), .Z(n37701) );
  XOR U39256 ( .A(n37702), .B(g_input[250]), .Z(n37699) );
  NAND U39257 ( .A(n37703), .B(mul_pow), .Z(n37702) );
  XOR U39258 ( .A(g_input[250]), .B(creg[250]), .Z(n37703) );
  XOR U39259 ( .A(n37704), .B(n37705), .Z(n37695) );
  ANDN U39260 ( .A(n37706), .B(n29246), .Z(n37705) );
  XOR U39261 ( .A(n37707), .B(\modmult_1/zin[0][248] ), .Z(n29246) );
  IV U39262 ( .A(n37704), .Z(n37707) );
  XNOR U39263 ( .A(n37704), .B(n29245), .Z(n37706) );
  XOR U39264 ( .A(n37708), .B(n37709), .Z(n29245) );
  AND U39265 ( .A(\modmult_1/xin[1023] ), .B(n37710), .Z(n37709) );
  IV U39266 ( .A(n37708), .Z(n37710) );
  XOR U39267 ( .A(n37711), .B(g_input[249]), .Z(n37708) );
  NAND U39268 ( .A(n37712), .B(mul_pow), .Z(n37711) );
  XOR U39269 ( .A(g_input[249]), .B(creg[249]), .Z(n37712) );
  XOR U39270 ( .A(n37713), .B(n37714), .Z(n37704) );
  ANDN U39271 ( .A(n37715), .B(n29252), .Z(n37714) );
  XOR U39272 ( .A(n37716), .B(\modmult_1/zin[0][247] ), .Z(n29252) );
  IV U39273 ( .A(n37713), .Z(n37716) );
  XNOR U39274 ( .A(n37713), .B(n29251), .Z(n37715) );
  XOR U39275 ( .A(n37717), .B(n37718), .Z(n29251) );
  AND U39276 ( .A(\modmult_1/xin[1023] ), .B(n37719), .Z(n37718) );
  IV U39277 ( .A(n37717), .Z(n37719) );
  XOR U39278 ( .A(n37720), .B(g_input[248]), .Z(n37717) );
  NAND U39279 ( .A(n37721), .B(mul_pow), .Z(n37720) );
  XOR U39280 ( .A(g_input[248]), .B(creg[248]), .Z(n37721) );
  XOR U39281 ( .A(n37722), .B(n37723), .Z(n37713) );
  ANDN U39282 ( .A(n37724), .B(n29258), .Z(n37723) );
  XOR U39283 ( .A(n37725), .B(\modmult_1/zin[0][246] ), .Z(n29258) );
  IV U39284 ( .A(n37722), .Z(n37725) );
  XNOR U39285 ( .A(n37722), .B(n29257), .Z(n37724) );
  XOR U39286 ( .A(n37726), .B(n37727), .Z(n29257) );
  AND U39287 ( .A(\modmult_1/xin[1023] ), .B(n37728), .Z(n37727) );
  IV U39288 ( .A(n37726), .Z(n37728) );
  XOR U39289 ( .A(n37729), .B(g_input[247]), .Z(n37726) );
  NAND U39290 ( .A(n37730), .B(mul_pow), .Z(n37729) );
  XOR U39291 ( .A(g_input[247]), .B(creg[247]), .Z(n37730) );
  XOR U39292 ( .A(n37731), .B(n37732), .Z(n37722) );
  ANDN U39293 ( .A(n37733), .B(n29264), .Z(n37732) );
  XOR U39294 ( .A(n37734), .B(\modmult_1/zin[0][245] ), .Z(n29264) );
  IV U39295 ( .A(n37731), .Z(n37734) );
  XNOR U39296 ( .A(n37731), .B(n29263), .Z(n37733) );
  XOR U39297 ( .A(n37735), .B(n37736), .Z(n29263) );
  AND U39298 ( .A(\modmult_1/xin[1023] ), .B(n37737), .Z(n37736) );
  IV U39299 ( .A(n37735), .Z(n37737) );
  XOR U39300 ( .A(n37738), .B(g_input[246]), .Z(n37735) );
  NAND U39301 ( .A(n37739), .B(mul_pow), .Z(n37738) );
  XOR U39302 ( .A(g_input[246]), .B(creg[246]), .Z(n37739) );
  XOR U39303 ( .A(n37740), .B(n37741), .Z(n37731) );
  ANDN U39304 ( .A(n37742), .B(n29270), .Z(n37741) );
  XOR U39305 ( .A(n37743), .B(\modmult_1/zin[0][244] ), .Z(n29270) );
  IV U39306 ( .A(n37740), .Z(n37743) );
  XNOR U39307 ( .A(n37740), .B(n29269), .Z(n37742) );
  XOR U39308 ( .A(n37744), .B(n37745), .Z(n29269) );
  AND U39309 ( .A(\modmult_1/xin[1023] ), .B(n37746), .Z(n37745) );
  IV U39310 ( .A(n37744), .Z(n37746) );
  XOR U39311 ( .A(n37747), .B(g_input[245]), .Z(n37744) );
  NAND U39312 ( .A(n37748), .B(mul_pow), .Z(n37747) );
  XOR U39313 ( .A(g_input[245]), .B(creg[245]), .Z(n37748) );
  XOR U39314 ( .A(n37749), .B(n37750), .Z(n37740) );
  ANDN U39315 ( .A(n37751), .B(n29276), .Z(n37750) );
  XOR U39316 ( .A(n37752), .B(\modmult_1/zin[0][243] ), .Z(n29276) );
  IV U39317 ( .A(n37749), .Z(n37752) );
  XNOR U39318 ( .A(n37749), .B(n29275), .Z(n37751) );
  XOR U39319 ( .A(n37753), .B(n37754), .Z(n29275) );
  AND U39320 ( .A(\modmult_1/xin[1023] ), .B(n37755), .Z(n37754) );
  IV U39321 ( .A(n37753), .Z(n37755) );
  XOR U39322 ( .A(n37756), .B(g_input[244]), .Z(n37753) );
  NAND U39323 ( .A(n37757), .B(mul_pow), .Z(n37756) );
  XOR U39324 ( .A(g_input[244]), .B(creg[244]), .Z(n37757) );
  XOR U39325 ( .A(n37758), .B(n37759), .Z(n37749) );
  ANDN U39326 ( .A(n37760), .B(n29282), .Z(n37759) );
  XOR U39327 ( .A(n37761), .B(\modmult_1/zin[0][242] ), .Z(n29282) );
  IV U39328 ( .A(n37758), .Z(n37761) );
  XNOR U39329 ( .A(n37758), .B(n29281), .Z(n37760) );
  XOR U39330 ( .A(n37762), .B(n37763), .Z(n29281) );
  AND U39331 ( .A(\modmult_1/xin[1023] ), .B(n37764), .Z(n37763) );
  IV U39332 ( .A(n37762), .Z(n37764) );
  XOR U39333 ( .A(n37765), .B(g_input[243]), .Z(n37762) );
  NAND U39334 ( .A(n37766), .B(mul_pow), .Z(n37765) );
  XOR U39335 ( .A(g_input[243]), .B(creg[243]), .Z(n37766) );
  XOR U39336 ( .A(n37767), .B(n37768), .Z(n37758) );
  ANDN U39337 ( .A(n37769), .B(n29288), .Z(n37768) );
  XOR U39338 ( .A(n37770), .B(\modmult_1/zin[0][241] ), .Z(n29288) );
  IV U39339 ( .A(n37767), .Z(n37770) );
  XNOR U39340 ( .A(n37767), .B(n29287), .Z(n37769) );
  XOR U39341 ( .A(n37771), .B(n37772), .Z(n29287) );
  AND U39342 ( .A(\modmult_1/xin[1023] ), .B(n37773), .Z(n37772) );
  IV U39343 ( .A(n37771), .Z(n37773) );
  XOR U39344 ( .A(n37774), .B(g_input[242]), .Z(n37771) );
  NAND U39345 ( .A(n37775), .B(mul_pow), .Z(n37774) );
  XOR U39346 ( .A(g_input[242]), .B(creg[242]), .Z(n37775) );
  XOR U39347 ( .A(n37776), .B(n37777), .Z(n37767) );
  ANDN U39348 ( .A(n37778), .B(n29294), .Z(n37777) );
  XOR U39349 ( .A(n37779), .B(\modmult_1/zin[0][240] ), .Z(n29294) );
  IV U39350 ( .A(n37776), .Z(n37779) );
  XNOR U39351 ( .A(n37776), .B(n29293), .Z(n37778) );
  XOR U39352 ( .A(n37780), .B(n37781), .Z(n29293) );
  AND U39353 ( .A(\modmult_1/xin[1023] ), .B(n37782), .Z(n37781) );
  IV U39354 ( .A(n37780), .Z(n37782) );
  XOR U39355 ( .A(n37783), .B(g_input[241]), .Z(n37780) );
  NAND U39356 ( .A(n37784), .B(mul_pow), .Z(n37783) );
  XOR U39357 ( .A(g_input[241]), .B(creg[241]), .Z(n37784) );
  XOR U39358 ( .A(n37785), .B(n37786), .Z(n37776) );
  ANDN U39359 ( .A(n37787), .B(n29300), .Z(n37786) );
  XOR U39360 ( .A(n37788), .B(\modmult_1/zin[0][239] ), .Z(n29300) );
  IV U39361 ( .A(n37785), .Z(n37788) );
  XNOR U39362 ( .A(n37785), .B(n29299), .Z(n37787) );
  XOR U39363 ( .A(n37789), .B(n37790), .Z(n29299) );
  AND U39364 ( .A(\modmult_1/xin[1023] ), .B(n37791), .Z(n37790) );
  IV U39365 ( .A(n37789), .Z(n37791) );
  XOR U39366 ( .A(n37792), .B(g_input[240]), .Z(n37789) );
  NAND U39367 ( .A(n37793), .B(mul_pow), .Z(n37792) );
  XOR U39368 ( .A(g_input[240]), .B(creg[240]), .Z(n37793) );
  XOR U39369 ( .A(n37794), .B(n37795), .Z(n37785) );
  ANDN U39370 ( .A(n37796), .B(n29306), .Z(n37795) );
  XOR U39371 ( .A(n37797), .B(\modmult_1/zin[0][238] ), .Z(n29306) );
  IV U39372 ( .A(n37794), .Z(n37797) );
  XNOR U39373 ( .A(n37794), .B(n29305), .Z(n37796) );
  XOR U39374 ( .A(n37798), .B(n37799), .Z(n29305) );
  AND U39375 ( .A(\modmult_1/xin[1023] ), .B(n37800), .Z(n37799) );
  IV U39376 ( .A(n37798), .Z(n37800) );
  XOR U39377 ( .A(n37801), .B(g_input[239]), .Z(n37798) );
  NAND U39378 ( .A(n37802), .B(mul_pow), .Z(n37801) );
  XOR U39379 ( .A(g_input[239]), .B(creg[239]), .Z(n37802) );
  XOR U39380 ( .A(n37803), .B(n37804), .Z(n37794) );
  ANDN U39381 ( .A(n37805), .B(n29312), .Z(n37804) );
  XOR U39382 ( .A(n37806), .B(\modmult_1/zin[0][237] ), .Z(n29312) );
  IV U39383 ( .A(n37803), .Z(n37806) );
  XNOR U39384 ( .A(n37803), .B(n29311), .Z(n37805) );
  XOR U39385 ( .A(n37807), .B(n37808), .Z(n29311) );
  AND U39386 ( .A(\modmult_1/xin[1023] ), .B(n37809), .Z(n37808) );
  IV U39387 ( .A(n37807), .Z(n37809) );
  XOR U39388 ( .A(n37810), .B(g_input[238]), .Z(n37807) );
  NAND U39389 ( .A(n37811), .B(mul_pow), .Z(n37810) );
  XOR U39390 ( .A(g_input[238]), .B(creg[238]), .Z(n37811) );
  XOR U39391 ( .A(n37812), .B(n37813), .Z(n37803) );
  ANDN U39392 ( .A(n37814), .B(n29318), .Z(n37813) );
  XOR U39393 ( .A(n37815), .B(\modmult_1/zin[0][236] ), .Z(n29318) );
  IV U39394 ( .A(n37812), .Z(n37815) );
  XNOR U39395 ( .A(n37812), .B(n29317), .Z(n37814) );
  XOR U39396 ( .A(n37816), .B(n37817), .Z(n29317) );
  AND U39397 ( .A(\modmult_1/xin[1023] ), .B(n37818), .Z(n37817) );
  IV U39398 ( .A(n37816), .Z(n37818) );
  XOR U39399 ( .A(n37819), .B(g_input[237]), .Z(n37816) );
  NAND U39400 ( .A(n37820), .B(mul_pow), .Z(n37819) );
  XOR U39401 ( .A(g_input[237]), .B(creg[237]), .Z(n37820) );
  XOR U39402 ( .A(n37821), .B(n37822), .Z(n37812) );
  ANDN U39403 ( .A(n37823), .B(n29324), .Z(n37822) );
  XOR U39404 ( .A(n37824), .B(\modmult_1/zin[0][235] ), .Z(n29324) );
  IV U39405 ( .A(n37821), .Z(n37824) );
  XNOR U39406 ( .A(n37821), .B(n29323), .Z(n37823) );
  XOR U39407 ( .A(n37825), .B(n37826), .Z(n29323) );
  AND U39408 ( .A(\modmult_1/xin[1023] ), .B(n37827), .Z(n37826) );
  IV U39409 ( .A(n37825), .Z(n37827) );
  XOR U39410 ( .A(n37828), .B(g_input[236]), .Z(n37825) );
  NAND U39411 ( .A(n37829), .B(mul_pow), .Z(n37828) );
  XOR U39412 ( .A(g_input[236]), .B(creg[236]), .Z(n37829) );
  XOR U39413 ( .A(n37830), .B(n37831), .Z(n37821) );
  ANDN U39414 ( .A(n37832), .B(n29330), .Z(n37831) );
  XOR U39415 ( .A(n37833), .B(\modmult_1/zin[0][234] ), .Z(n29330) );
  IV U39416 ( .A(n37830), .Z(n37833) );
  XNOR U39417 ( .A(n37830), .B(n29329), .Z(n37832) );
  XOR U39418 ( .A(n37834), .B(n37835), .Z(n29329) );
  AND U39419 ( .A(\modmult_1/xin[1023] ), .B(n37836), .Z(n37835) );
  IV U39420 ( .A(n37834), .Z(n37836) );
  XOR U39421 ( .A(n37837), .B(g_input[235]), .Z(n37834) );
  NAND U39422 ( .A(n37838), .B(mul_pow), .Z(n37837) );
  XOR U39423 ( .A(g_input[235]), .B(creg[235]), .Z(n37838) );
  XOR U39424 ( .A(n37839), .B(n37840), .Z(n37830) );
  ANDN U39425 ( .A(n37841), .B(n29336), .Z(n37840) );
  XOR U39426 ( .A(n37842), .B(\modmult_1/zin[0][233] ), .Z(n29336) );
  IV U39427 ( .A(n37839), .Z(n37842) );
  XNOR U39428 ( .A(n37839), .B(n29335), .Z(n37841) );
  XOR U39429 ( .A(n37843), .B(n37844), .Z(n29335) );
  AND U39430 ( .A(\modmult_1/xin[1023] ), .B(n37845), .Z(n37844) );
  IV U39431 ( .A(n37843), .Z(n37845) );
  XOR U39432 ( .A(n37846), .B(g_input[234]), .Z(n37843) );
  NAND U39433 ( .A(n37847), .B(mul_pow), .Z(n37846) );
  XOR U39434 ( .A(g_input[234]), .B(creg[234]), .Z(n37847) );
  XOR U39435 ( .A(n37848), .B(n37849), .Z(n37839) );
  ANDN U39436 ( .A(n37850), .B(n29342), .Z(n37849) );
  XOR U39437 ( .A(n37851), .B(\modmult_1/zin[0][232] ), .Z(n29342) );
  IV U39438 ( .A(n37848), .Z(n37851) );
  XNOR U39439 ( .A(n37848), .B(n29341), .Z(n37850) );
  XOR U39440 ( .A(n37852), .B(n37853), .Z(n29341) );
  AND U39441 ( .A(\modmult_1/xin[1023] ), .B(n37854), .Z(n37853) );
  IV U39442 ( .A(n37852), .Z(n37854) );
  XOR U39443 ( .A(n37855), .B(g_input[233]), .Z(n37852) );
  NAND U39444 ( .A(n37856), .B(mul_pow), .Z(n37855) );
  XOR U39445 ( .A(g_input[233]), .B(creg[233]), .Z(n37856) );
  XOR U39446 ( .A(n37857), .B(n37858), .Z(n37848) );
  ANDN U39447 ( .A(n37859), .B(n29348), .Z(n37858) );
  XOR U39448 ( .A(n37860), .B(\modmult_1/zin[0][231] ), .Z(n29348) );
  IV U39449 ( .A(n37857), .Z(n37860) );
  XNOR U39450 ( .A(n37857), .B(n29347), .Z(n37859) );
  XOR U39451 ( .A(n37861), .B(n37862), .Z(n29347) );
  AND U39452 ( .A(\modmult_1/xin[1023] ), .B(n37863), .Z(n37862) );
  IV U39453 ( .A(n37861), .Z(n37863) );
  XOR U39454 ( .A(n37864), .B(g_input[232]), .Z(n37861) );
  NAND U39455 ( .A(n37865), .B(mul_pow), .Z(n37864) );
  XOR U39456 ( .A(g_input[232]), .B(creg[232]), .Z(n37865) );
  XOR U39457 ( .A(n37866), .B(n37867), .Z(n37857) );
  ANDN U39458 ( .A(n37868), .B(n29354), .Z(n37867) );
  XOR U39459 ( .A(n37869), .B(\modmult_1/zin[0][230] ), .Z(n29354) );
  IV U39460 ( .A(n37866), .Z(n37869) );
  XNOR U39461 ( .A(n37866), .B(n29353), .Z(n37868) );
  XOR U39462 ( .A(n37870), .B(n37871), .Z(n29353) );
  AND U39463 ( .A(\modmult_1/xin[1023] ), .B(n37872), .Z(n37871) );
  IV U39464 ( .A(n37870), .Z(n37872) );
  XOR U39465 ( .A(n37873), .B(g_input[231]), .Z(n37870) );
  NAND U39466 ( .A(n37874), .B(mul_pow), .Z(n37873) );
  XOR U39467 ( .A(g_input[231]), .B(creg[231]), .Z(n37874) );
  XOR U39468 ( .A(n37875), .B(n37876), .Z(n37866) );
  ANDN U39469 ( .A(n37877), .B(n29360), .Z(n37876) );
  XOR U39470 ( .A(n37878), .B(\modmult_1/zin[0][229] ), .Z(n29360) );
  IV U39471 ( .A(n37875), .Z(n37878) );
  XNOR U39472 ( .A(n37875), .B(n29359), .Z(n37877) );
  XOR U39473 ( .A(n37879), .B(n37880), .Z(n29359) );
  AND U39474 ( .A(\modmult_1/xin[1023] ), .B(n37881), .Z(n37880) );
  IV U39475 ( .A(n37879), .Z(n37881) );
  XOR U39476 ( .A(n37882), .B(g_input[230]), .Z(n37879) );
  NAND U39477 ( .A(n37883), .B(mul_pow), .Z(n37882) );
  XOR U39478 ( .A(g_input[230]), .B(creg[230]), .Z(n37883) );
  XOR U39479 ( .A(n37884), .B(n37885), .Z(n37875) );
  ANDN U39480 ( .A(n37886), .B(n29366), .Z(n37885) );
  XOR U39481 ( .A(n37887), .B(\modmult_1/zin[0][228] ), .Z(n29366) );
  IV U39482 ( .A(n37884), .Z(n37887) );
  XNOR U39483 ( .A(n37884), .B(n29365), .Z(n37886) );
  XOR U39484 ( .A(n37888), .B(n37889), .Z(n29365) );
  AND U39485 ( .A(\modmult_1/xin[1023] ), .B(n37890), .Z(n37889) );
  IV U39486 ( .A(n37888), .Z(n37890) );
  XOR U39487 ( .A(n37891), .B(g_input[229]), .Z(n37888) );
  NAND U39488 ( .A(n37892), .B(mul_pow), .Z(n37891) );
  XOR U39489 ( .A(g_input[229]), .B(creg[229]), .Z(n37892) );
  XOR U39490 ( .A(n37893), .B(n37894), .Z(n37884) );
  ANDN U39491 ( .A(n37895), .B(n29372), .Z(n37894) );
  XOR U39492 ( .A(n37896), .B(\modmult_1/zin[0][227] ), .Z(n29372) );
  IV U39493 ( .A(n37893), .Z(n37896) );
  XNOR U39494 ( .A(n37893), .B(n29371), .Z(n37895) );
  XOR U39495 ( .A(n37897), .B(n37898), .Z(n29371) );
  AND U39496 ( .A(\modmult_1/xin[1023] ), .B(n37899), .Z(n37898) );
  IV U39497 ( .A(n37897), .Z(n37899) );
  XOR U39498 ( .A(n37900), .B(g_input[228]), .Z(n37897) );
  NAND U39499 ( .A(n37901), .B(mul_pow), .Z(n37900) );
  XOR U39500 ( .A(g_input[228]), .B(creg[228]), .Z(n37901) );
  XOR U39501 ( .A(n37902), .B(n37903), .Z(n37893) );
  ANDN U39502 ( .A(n37904), .B(n29378), .Z(n37903) );
  XOR U39503 ( .A(n37905), .B(\modmult_1/zin[0][226] ), .Z(n29378) );
  IV U39504 ( .A(n37902), .Z(n37905) );
  XNOR U39505 ( .A(n37902), .B(n29377), .Z(n37904) );
  XOR U39506 ( .A(n37906), .B(n37907), .Z(n29377) );
  AND U39507 ( .A(\modmult_1/xin[1023] ), .B(n37908), .Z(n37907) );
  IV U39508 ( .A(n37906), .Z(n37908) );
  XOR U39509 ( .A(n37909), .B(g_input[227]), .Z(n37906) );
  NAND U39510 ( .A(n37910), .B(mul_pow), .Z(n37909) );
  XOR U39511 ( .A(g_input[227]), .B(creg[227]), .Z(n37910) );
  XOR U39512 ( .A(n37911), .B(n37912), .Z(n37902) );
  ANDN U39513 ( .A(n37913), .B(n29384), .Z(n37912) );
  XOR U39514 ( .A(n37914), .B(\modmult_1/zin[0][225] ), .Z(n29384) );
  IV U39515 ( .A(n37911), .Z(n37914) );
  XNOR U39516 ( .A(n37911), .B(n29383), .Z(n37913) );
  XOR U39517 ( .A(n37915), .B(n37916), .Z(n29383) );
  AND U39518 ( .A(\modmult_1/xin[1023] ), .B(n37917), .Z(n37916) );
  IV U39519 ( .A(n37915), .Z(n37917) );
  XOR U39520 ( .A(n37918), .B(g_input[226]), .Z(n37915) );
  NAND U39521 ( .A(n37919), .B(mul_pow), .Z(n37918) );
  XOR U39522 ( .A(g_input[226]), .B(creg[226]), .Z(n37919) );
  XOR U39523 ( .A(n37920), .B(n37921), .Z(n37911) );
  ANDN U39524 ( .A(n37922), .B(n29390), .Z(n37921) );
  XOR U39525 ( .A(n37923), .B(\modmult_1/zin[0][224] ), .Z(n29390) );
  IV U39526 ( .A(n37920), .Z(n37923) );
  XNOR U39527 ( .A(n37920), .B(n29389), .Z(n37922) );
  XOR U39528 ( .A(n37924), .B(n37925), .Z(n29389) );
  AND U39529 ( .A(\modmult_1/xin[1023] ), .B(n37926), .Z(n37925) );
  IV U39530 ( .A(n37924), .Z(n37926) );
  XOR U39531 ( .A(n37927), .B(g_input[225]), .Z(n37924) );
  NAND U39532 ( .A(n37928), .B(mul_pow), .Z(n37927) );
  XOR U39533 ( .A(g_input[225]), .B(creg[225]), .Z(n37928) );
  XOR U39534 ( .A(n37929), .B(n37930), .Z(n37920) );
  ANDN U39535 ( .A(n37931), .B(n29396), .Z(n37930) );
  XOR U39536 ( .A(n37932), .B(\modmult_1/zin[0][223] ), .Z(n29396) );
  IV U39537 ( .A(n37929), .Z(n37932) );
  XNOR U39538 ( .A(n37929), .B(n29395), .Z(n37931) );
  XOR U39539 ( .A(n37933), .B(n37934), .Z(n29395) );
  AND U39540 ( .A(\modmult_1/xin[1023] ), .B(n37935), .Z(n37934) );
  IV U39541 ( .A(n37933), .Z(n37935) );
  XOR U39542 ( .A(n37936), .B(g_input[224]), .Z(n37933) );
  NAND U39543 ( .A(n37937), .B(mul_pow), .Z(n37936) );
  XOR U39544 ( .A(g_input[224]), .B(creg[224]), .Z(n37937) );
  XOR U39545 ( .A(n37938), .B(n37939), .Z(n37929) );
  ANDN U39546 ( .A(n37940), .B(n29402), .Z(n37939) );
  XOR U39547 ( .A(n37941), .B(\modmult_1/zin[0][222] ), .Z(n29402) );
  IV U39548 ( .A(n37938), .Z(n37941) );
  XNOR U39549 ( .A(n37938), .B(n29401), .Z(n37940) );
  XOR U39550 ( .A(n37942), .B(n37943), .Z(n29401) );
  AND U39551 ( .A(\modmult_1/xin[1023] ), .B(n37944), .Z(n37943) );
  IV U39552 ( .A(n37942), .Z(n37944) );
  XOR U39553 ( .A(n37945), .B(g_input[223]), .Z(n37942) );
  NAND U39554 ( .A(n37946), .B(mul_pow), .Z(n37945) );
  XOR U39555 ( .A(g_input[223]), .B(creg[223]), .Z(n37946) );
  XOR U39556 ( .A(n37947), .B(n37948), .Z(n37938) );
  ANDN U39557 ( .A(n37949), .B(n29408), .Z(n37948) );
  XOR U39558 ( .A(n37950), .B(\modmult_1/zin[0][221] ), .Z(n29408) );
  IV U39559 ( .A(n37947), .Z(n37950) );
  XNOR U39560 ( .A(n37947), .B(n29407), .Z(n37949) );
  XOR U39561 ( .A(n37951), .B(n37952), .Z(n29407) );
  AND U39562 ( .A(\modmult_1/xin[1023] ), .B(n37953), .Z(n37952) );
  IV U39563 ( .A(n37951), .Z(n37953) );
  XOR U39564 ( .A(n37954), .B(g_input[222]), .Z(n37951) );
  NAND U39565 ( .A(n37955), .B(mul_pow), .Z(n37954) );
  XOR U39566 ( .A(g_input[222]), .B(creg[222]), .Z(n37955) );
  XOR U39567 ( .A(n37956), .B(n37957), .Z(n37947) );
  ANDN U39568 ( .A(n37958), .B(n29414), .Z(n37957) );
  XOR U39569 ( .A(n37959), .B(\modmult_1/zin[0][220] ), .Z(n29414) );
  IV U39570 ( .A(n37956), .Z(n37959) );
  XNOR U39571 ( .A(n37956), .B(n29413), .Z(n37958) );
  XOR U39572 ( .A(n37960), .B(n37961), .Z(n29413) );
  AND U39573 ( .A(\modmult_1/xin[1023] ), .B(n37962), .Z(n37961) );
  IV U39574 ( .A(n37960), .Z(n37962) );
  XOR U39575 ( .A(n37963), .B(g_input[221]), .Z(n37960) );
  NAND U39576 ( .A(n37964), .B(mul_pow), .Z(n37963) );
  XOR U39577 ( .A(g_input[221]), .B(creg[221]), .Z(n37964) );
  XOR U39578 ( .A(n37965), .B(n37966), .Z(n37956) );
  ANDN U39579 ( .A(n37967), .B(n29420), .Z(n37966) );
  XOR U39580 ( .A(n37968), .B(\modmult_1/zin[0][219] ), .Z(n29420) );
  IV U39581 ( .A(n37965), .Z(n37968) );
  XNOR U39582 ( .A(n37965), .B(n29419), .Z(n37967) );
  XOR U39583 ( .A(n37969), .B(n37970), .Z(n29419) );
  AND U39584 ( .A(\modmult_1/xin[1023] ), .B(n37971), .Z(n37970) );
  IV U39585 ( .A(n37969), .Z(n37971) );
  XOR U39586 ( .A(n37972), .B(g_input[220]), .Z(n37969) );
  NAND U39587 ( .A(n37973), .B(mul_pow), .Z(n37972) );
  XOR U39588 ( .A(g_input[220]), .B(creg[220]), .Z(n37973) );
  XOR U39589 ( .A(n37974), .B(n37975), .Z(n37965) );
  ANDN U39590 ( .A(n37976), .B(n29426), .Z(n37975) );
  XOR U39591 ( .A(n37977), .B(\modmult_1/zin[0][218] ), .Z(n29426) );
  IV U39592 ( .A(n37974), .Z(n37977) );
  XNOR U39593 ( .A(n37974), .B(n29425), .Z(n37976) );
  XOR U39594 ( .A(n37978), .B(n37979), .Z(n29425) );
  AND U39595 ( .A(\modmult_1/xin[1023] ), .B(n37980), .Z(n37979) );
  IV U39596 ( .A(n37978), .Z(n37980) );
  XOR U39597 ( .A(n37981), .B(g_input[219]), .Z(n37978) );
  NAND U39598 ( .A(n37982), .B(mul_pow), .Z(n37981) );
  XOR U39599 ( .A(g_input[219]), .B(creg[219]), .Z(n37982) );
  XOR U39600 ( .A(n37983), .B(n37984), .Z(n37974) );
  ANDN U39601 ( .A(n37985), .B(n29432), .Z(n37984) );
  XOR U39602 ( .A(n37986), .B(\modmult_1/zin[0][217] ), .Z(n29432) );
  IV U39603 ( .A(n37983), .Z(n37986) );
  XNOR U39604 ( .A(n37983), .B(n29431), .Z(n37985) );
  XOR U39605 ( .A(n37987), .B(n37988), .Z(n29431) );
  AND U39606 ( .A(\modmult_1/xin[1023] ), .B(n37989), .Z(n37988) );
  IV U39607 ( .A(n37987), .Z(n37989) );
  XOR U39608 ( .A(n37990), .B(g_input[218]), .Z(n37987) );
  NAND U39609 ( .A(n37991), .B(mul_pow), .Z(n37990) );
  XOR U39610 ( .A(g_input[218]), .B(creg[218]), .Z(n37991) );
  XOR U39611 ( .A(n37992), .B(n37993), .Z(n37983) );
  ANDN U39612 ( .A(n37994), .B(n29438), .Z(n37993) );
  XOR U39613 ( .A(n37995), .B(\modmult_1/zin[0][216] ), .Z(n29438) );
  IV U39614 ( .A(n37992), .Z(n37995) );
  XNOR U39615 ( .A(n37992), .B(n29437), .Z(n37994) );
  XOR U39616 ( .A(n37996), .B(n37997), .Z(n29437) );
  AND U39617 ( .A(\modmult_1/xin[1023] ), .B(n37998), .Z(n37997) );
  IV U39618 ( .A(n37996), .Z(n37998) );
  XOR U39619 ( .A(n37999), .B(g_input[217]), .Z(n37996) );
  NAND U39620 ( .A(n38000), .B(mul_pow), .Z(n37999) );
  XOR U39621 ( .A(g_input[217]), .B(creg[217]), .Z(n38000) );
  XOR U39622 ( .A(n38001), .B(n38002), .Z(n37992) );
  ANDN U39623 ( .A(n38003), .B(n29444), .Z(n38002) );
  XOR U39624 ( .A(n38004), .B(\modmult_1/zin[0][215] ), .Z(n29444) );
  IV U39625 ( .A(n38001), .Z(n38004) );
  XNOR U39626 ( .A(n38001), .B(n29443), .Z(n38003) );
  XOR U39627 ( .A(n38005), .B(n38006), .Z(n29443) );
  AND U39628 ( .A(\modmult_1/xin[1023] ), .B(n38007), .Z(n38006) );
  IV U39629 ( .A(n38005), .Z(n38007) );
  XOR U39630 ( .A(n38008), .B(g_input[216]), .Z(n38005) );
  NAND U39631 ( .A(n38009), .B(mul_pow), .Z(n38008) );
  XOR U39632 ( .A(g_input[216]), .B(creg[216]), .Z(n38009) );
  XOR U39633 ( .A(n38010), .B(n38011), .Z(n38001) );
  ANDN U39634 ( .A(n38012), .B(n29450), .Z(n38011) );
  XOR U39635 ( .A(n38013), .B(\modmult_1/zin[0][214] ), .Z(n29450) );
  IV U39636 ( .A(n38010), .Z(n38013) );
  XNOR U39637 ( .A(n38010), .B(n29449), .Z(n38012) );
  XOR U39638 ( .A(n38014), .B(n38015), .Z(n29449) );
  AND U39639 ( .A(\modmult_1/xin[1023] ), .B(n38016), .Z(n38015) );
  IV U39640 ( .A(n38014), .Z(n38016) );
  XOR U39641 ( .A(n38017), .B(g_input[215]), .Z(n38014) );
  NAND U39642 ( .A(n38018), .B(mul_pow), .Z(n38017) );
  XOR U39643 ( .A(g_input[215]), .B(creg[215]), .Z(n38018) );
  XOR U39644 ( .A(n38019), .B(n38020), .Z(n38010) );
  ANDN U39645 ( .A(n38021), .B(n29456), .Z(n38020) );
  XOR U39646 ( .A(n38022), .B(\modmult_1/zin[0][213] ), .Z(n29456) );
  IV U39647 ( .A(n38019), .Z(n38022) );
  XNOR U39648 ( .A(n38019), .B(n29455), .Z(n38021) );
  XOR U39649 ( .A(n38023), .B(n38024), .Z(n29455) );
  AND U39650 ( .A(\modmult_1/xin[1023] ), .B(n38025), .Z(n38024) );
  IV U39651 ( .A(n38023), .Z(n38025) );
  XOR U39652 ( .A(n38026), .B(g_input[214]), .Z(n38023) );
  NAND U39653 ( .A(n38027), .B(mul_pow), .Z(n38026) );
  XOR U39654 ( .A(g_input[214]), .B(creg[214]), .Z(n38027) );
  XOR U39655 ( .A(n38028), .B(n38029), .Z(n38019) );
  ANDN U39656 ( .A(n38030), .B(n29462), .Z(n38029) );
  XOR U39657 ( .A(n38031), .B(\modmult_1/zin[0][212] ), .Z(n29462) );
  IV U39658 ( .A(n38028), .Z(n38031) );
  XNOR U39659 ( .A(n38028), .B(n29461), .Z(n38030) );
  XOR U39660 ( .A(n38032), .B(n38033), .Z(n29461) );
  AND U39661 ( .A(\modmult_1/xin[1023] ), .B(n38034), .Z(n38033) );
  IV U39662 ( .A(n38032), .Z(n38034) );
  XOR U39663 ( .A(n38035), .B(g_input[213]), .Z(n38032) );
  NAND U39664 ( .A(n38036), .B(mul_pow), .Z(n38035) );
  XOR U39665 ( .A(g_input[213]), .B(creg[213]), .Z(n38036) );
  XOR U39666 ( .A(n38037), .B(n38038), .Z(n38028) );
  ANDN U39667 ( .A(n38039), .B(n29468), .Z(n38038) );
  XOR U39668 ( .A(n38040), .B(\modmult_1/zin[0][211] ), .Z(n29468) );
  IV U39669 ( .A(n38037), .Z(n38040) );
  XNOR U39670 ( .A(n38037), .B(n29467), .Z(n38039) );
  XOR U39671 ( .A(n38041), .B(n38042), .Z(n29467) );
  AND U39672 ( .A(\modmult_1/xin[1023] ), .B(n38043), .Z(n38042) );
  IV U39673 ( .A(n38041), .Z(n38043) );
  XOR U39674 ( .A(n38044), .B(g_input[212]), .Z(n38041) );
  NAND U39675 ( .A(n38045), .B(mul_pow), .Z(n38044) );
  XOR U39676 ( .A(g_input[212]), .B(creg[212]), .Z(n38045) );
  XOR U39677 ( .A(n38046), .B(n38047), .Z(n38037) );
  ANDN U39678 ( .A(n38048), .B(n29474), .Z(n38047) );
  XOR U39679 ( .A(n38049), .B(\modmult_1/zin[0][210] ), .Z(n29474) );
  IV U39680 ( .A(n38046), .Z(n38049) );
  XNOR U39681 ( .A(n38046), .B(n29473), .Z(n38048) );
  XOR U39682 ( .A(n38050), .B(n38051), .Z(n29473) );
  AND U39683 ( .A(\modmult_1/xin[1023] ), .B(n38052), .Z(n38051) );
  IV U39684 ( .A(n38050), .Z(n38052) );
  XOR U39685 ( .A(n38053), .B(g_input[211]), .Z(n38050) );
  NAND U39686 ( .A(n38054), .B(mul_pow), .Z(n38053) );
  XOR U39687 ( .A(g_input[211]), .B(creg[211]), .Z(n38054) );
  XOR U39688 ( .A(n38055), .B(n38056), .Z(n38046) );
  ANDN U39689 ( .A(n38057), .B(n29480), .Z(n38056) );
  XOR U39690 ( .A(n38058), .B(\modmult_1/zin[0][209] ), .Z(n29480) );
  IV U39691 ( .A(n38055), .Z(n38058) );
  XNOR U39692 ( .A(n38055), .B(n29479), .Z(n38057) );
  XOR U39693 ( .A(n38059), .B(n38060), .Z(n29479) );
  AND U39694 ( .A(\modmult_1/xin[1023] ), .B(n38061), .Z(n38060) );
  IV U39695 ( .A(n38059), .Z(n38061) );
  XOR U39696 ( .A(n38062), .B(g_input[210]), .Z(n38059) );
  NAND U39697 ( .A(n38063), .B(mul_pow), .Z(n38062) );
  XOR U39698 ( .A(g_input[210]), .B(creg[210]), .Z(n38063) );
  XOR U39699 ( .A(n38064), .B(n38065), .Z(n38055) );
  ANDN U39700 ( .A(n38066), .B(n29486), .Z(n38065) );
  XOR U39701 ( .A(n38067), .B(\modmult_1/zin[0][208] ), .Z(n29486) );
  IV U39702 ( .A(n38064), .Z(n38067) );
  XNOR U39703 ( .A(n38064), .B(n29485), .Z(n38066) );
  XOR U39704 ( .A(n38068), .B(n38069), .Z(n29485) );
  AND U39705 ( .A(\modmult_1/xin[1023] ), .B(n38070), .Z(n38069) );
  IV U39706 ( .A(n38068), .Z(n38070) );
  XOR U39707 ( .A(n38071), .B(g_input[209]), .Z(n38068) );
  NAND U39708 ( .A(n38072), .B(mul_pow), .Z(n38071) );
  XOR U39709 ( .A(g_input[209]), .B(creg[209]), .Z(n38072) );
  XOR U39710 ( .A(n38073), .B(n38074), .Z(n38064) );
  ANDN U39711 ( .A(n38075), .B(n29492), .Z(n38074) );
  XOR U39712 ( .A(n38076), .B(\modmult_1/zin[0][207] ), .Z(n29492) );
  IV U39713 ( .A(n38073), .Z(n38076) );
  XNOR U39714 ( .A(n38073), .B(n29491), .Z(n38075) );
  XOR U39715 ( .A(n38077), .B(n38078), .Z(n29491) );
  AND U39716 ( .A(\modmult_1/xin[1023] ), .B(n38079), .Z(n38078) );
  IV U39717 ( .A(n38077), .Z(n38079) );
  XOR U39718 ( .A(n38080), .B(g_input[208]), .Z(n38077) );
  NAND U39719 ( .A(n38081), .B(mul_pow), .Z(n38080) );
  XOR U39720 ( .A(g_input[208]), .B(creg[208]), .Z(n38081) );
  XOR U39721 ( .A(n38082), .B(n38083), .Z(n38073) );
  ANDN U39722 ( .A(n38084), .B(n29498), .Z(n38083) );
  XOR U39723 ( .A(n38085), .B(\modmult_1/zin[0][206] ), .Z(n29498) );
  IV U39724 ( .A(n38082), .Z(n38085) );
  XNOR U39725 ( .A(n38082), .B(n29497), .Z(n38084) );
  XOR U39726 ( .A(n38086), .B(n38087), .Z(n29497) );
  AND U39727 ( .A(\modmult_1/xin[1023] ), .B(n38088), .Z(n38087) );
  IV U39728 ( .A(n38086), .Z(n38088) );
  XOR U39729 ( .A(n38089), .B(g_input[207]), .Z(n38086) );
  NAND U39730 ( .A(n38090), .B(mul_pow), .Z(n38089) );
  XOR U39731 ( .A(g_input[207]), .B(creg[207]), .Z(n38090) );
  XOR U39732 ( .A(n38091), .B(n38092), .Z(n38082) );
  ANDN U39733 ( .A(n38093), .B(n29504), .Z(n38092) );
  XOR U39734 ( .A(n38094), .B(\modmult_1/zin[0][205] ), .Z(n29504) );
  IV U39735 ( .A(n38091), .Z(n38094) );
  XNOR U39736 ( .A(n38091), .B(n29503), .Z(n38093) );
  XOR U39737 ( .A(n38095), .B(n38096), .Z(n29503) );
  AND U39738 ( .A(\modmult_1/xin[1023] ), .B(n38097), .Z(n38096) );
  IV U39739 ( .A(n38095), .Z(n38097) );
  XOR U39740 ( .A(n38098), .B(g_input[206]), .Z(n38095) );
  NAND U39741 ( .A(n38099), .B(mul_pow), .Z(n38098) );
  XOR U39742 ( .A(g_input[206]), .B(creg[206]), .Z(n38099) );
  XOR U39743 ( .A(n38100), .B(n38101), .Z(n38091) );
  ANDN U39744 ( .A(n38102), .B(n29510), .Z(n38101) );
  XOR U39745 ( .A(n38103), .B(\modmult_1/zin[0][204] ), .Z(n29510) );
  IV U39746 ( .A(n38100), .Z(n38103) );
  XNOR U39747 ( .A(n38100), .B(n29509), .Z(n38102) );
  XOR U39748 ( .A(n38104), .B(n38105), .Z(n29509) );
  AND U39749 ( .A(\modmult_1/xin[1023] ), .B(n38106), .Z(n38105) );
  IV U39750 ( .A(n38104), .Z(n38106) );
  XOR U39751 ( .A(n38107), .B(g_input[205]), .Z(n38104) );
  NAND U39752 ( .A(n38108), .B(mul_pow), .Z(n38107) );
  XOR U39753 ( .A(g_input[205]), .B(creg[205]), .Z(n38108) );
  XOR U39754 ( .A(n38109), .B(n38110), .Z(n38100) );
  ANDN U39755 ( .A(n38111), .B(n29516), .Z(n38110) );
  XOR U39756 ( .A(n38112), .B(\modmult_1/zin[0][203] ), .Z(n29516) );
  IV U39757 ( .A(n38109), .Z(n38112) );
  XNOR U39758 ( .A(n38109), .B(n29515), .Z(n38111) );
  XOR U39759 ( .A(n38113), .B(n38114), .Z(n29515) );
  AND U39760 ( .A(\modmult_1/xin[1023] ), .B(n38115), .Z(n38114) );
  IV U39761 ( .A(n38113), .Z(n38115) );
  XOR U39762 ( .A(n38116), .B(g_input[204]), .Z(n38113) );
  NAND U39763 ( .A(n38117), .B(mul_pow), .Z(n38116) );
  XOR U39764 ( .A(g_input[204]), .B(creg[204]), .Z(n38117) );
  XOR U39765 ( .A(n38118), .B(n38119), .Z(n38109) );
  ANDN U39766 ( .A(n38120), .B(n29522), .Z(n38119) );
  XOR U39767 ( .A(n38121), .B(\modmult_1/zin[0][202] ), .Z(n29522) );
  IV U39768 ( .A(n38118), .Z(n38121) );
  XNOR U39769 ( .A(n38118), .B(n29521), .Z(n38120) );
  XOR U39770 ( .A(n38122), .B(n38123), .Z(n29521) );
  AND U39771 ( .A(\modmult_1/xin[1023] ), .B(n38124), .Z(n38123) );
  IV U39772 ( .A(n38122), .Z(n38124) );
  XOR U39773 ( .A(n38125), .B(g_input[203]), .Z(n38122) );
  NAND U39774 ( .A(n38126), .B(mul_pow), .Z(n38125) );
  XOR U39775 ( .A(g_input[203]), .B(creg[203]), .Z(n38126) );
  XOR U39776 ( .A(n38127), .B(n38128), .Z(n38118) );
  ANDN U39777 ( .A(n38129), .B(n29528), .Z(n38128) );
  XOR U39778 ( .A(n38130), .B(\modmult_1/zin[0][201] ), .Z(n29528) );
  IV U39779 ( .A(n38127), .Z(n38130) );
  XNOR U39780 ( .A(n38127), .B(n29527), .Z(n38129) );
  XOR U39781 ( .A(n38131), .B(n38132), .Z(n29527) );
  AND U39782 ( .A(\modmult_1/xin[1023] ), .B(n38133), .Z(n38132) );
  IV U39783 ( .A(n38131), .Z(n38133) );
  XOR U39784 ( .A(n38134), .B(g_input[202]), .Z(n38131) );
  NAND U39785 ( .A(n38135), .B(mul_pow), .Z(n38134) );
  XOR U39786 ( .A(g_input[202]), .B(creg[202]), .Z(n38135) );
  XOR U39787 ( .A(n38136), .B(n38137), .Z(n38127) );
  ANDN U39788 ( .A(n38138), .B(n29534), .Z(n38137) );
  XOR U39789 ( .A(n38139), .B(\modmult_1/zin[0][200] ), .Z(n29534) );
  IV U39790 ( .A(n38136), .Z(n38139) );
  XNOR U39791 ( .A(n38136), .B(n29533), .Z(n38138) );
  XOR U39792 ( .A(n38140), .B(n38141), .Z(n29533) );
  AND U39793 ( .A(\modmult_1/xin[1023] ), .B(n38142), .Z(n38141) );
  IV U39794 ( .A(n38140), .Z(n38142) );
  XOR U39795 ( .A(n38143), .B(g_input[201]), .Z(n38140) );
  NAND U39796 ( .A(n38144), .B(mul_pow), .Z(n38143) );
  XOR U39797 ( .A(g_input[201]), .B(creg[201]), .Z(n38144) );
  XOR U39798 ( .A(n38145), .B(n38146), .Z(n38136) );
  ANDN U39799 ( .A(n38147), .B(n29540), .Z(n38146) );
  XOR U39800 ( .A(n38148), .B(\modmult_1/zin[0][199] ), .Z(n29540) );
  IV U39801 ( .A(n38145), .Z(n38148) );
  XNOR U39802 ( .A(n38145), .B(n29539), .Z(n38147) );
  XOR U39803 ( .A(n38149), .B(n38150), .Z(n29539) );
  AND U39804 ( .A(\modmult_1/xin[1023] ), .B(n38151), .Z(n38150) );
  IV U39805 ( .A(n38149), .Z(n38151) );
  XOR U39806 ( .A(n38152), .B(g_input[200]), .Z(n38149) );
  NAND U39807 ( .A(n38153), .B(mul_pow), .Z(n38152) );
  XOR U39808 ( .A(g_input[200]), .B(creg[200]), .Z(n38153) );
  XOR U39809 ( .A(n38154), .B(n38155), .Z(n38145) );
  ANDN U39810 ( .A(n38156), .B(n29546), .Z(n38155) );
  XOR U39811 ( .A(n38157), .B(\modmult_1/zin[0][198] ), .Z(n29546) );
  IV U39812 ( .A(n38154), .Z(n38157) );
  XNOR U39813 ( .A(n38154), .B(n29545), .Z(n38156) );
  XOR U39814 ( .A(n38158), .B(n38159), .Z(n29545) );
  AND U39815 ( .A(\modmult_1/xin[1023] ), .B(n38160), .Z(n38159) );
  IV U39816 ( .A(n38158), .Z(n38160) );
  XOR U39817 ( .A(n38161), .B(g_input[199]), .Z(n38158) );
  NAND U39818 ( .A(n38162), .B(mul_pow), .Z(n38161) );
  XOR U39819 ( .A(g_input[199]), .B(creg[199]), .Z(n38162) );
  XOR U39820 ( .A(n38163), .B(n38164), .Z(n38154) );
  ANDN U39821 ( .A(n38165), .B(n29552), .Z(n38164) );
  XOR U39822 ( .A(n38166), .B(\modmult_1/zin[0][197] ), .Z(n29552) );
  IV U39823 ( .A(n38163), .Z(n38166) );
  XNOR U39824 ( .A(n38163), .B(n29551), .Z(n38165) );
  XOR U39825 ( .A(n38167), .B(n38168), .Z(n29551) );
  AND U39826 ( .A(\modmult_1/xin[1023] ), .B(n38169), .Z(n38168) );
  IV U39827 ( .A(n38167), .Z(n38169) );
  XOR U39828 ( .A(n38170), .B(g_input[198]), .Z(n38167) );
  NAND U39829 ( .A(n38171), .B(mul_pow), .Z(n38170) );
  XOR U39830 ( .A(g_input[198]), .B(creg[198]), .Z(n38171) );
  XOR U39831 ( .A(n38172), .B(n38173), .Z(n38163) );
  ANDN U39832 ( .A(n38174), .B(n29558), .Z(n38173) );
  XOR U39833 ( .A(n38175), .B(\modmult_1/zin[0][196] ), .Z(n29558) );
  IV U39834 ( .A(n38172), .Z(n38175) );
  XNOR U39835 ( .A(n38172), .B(n29557), .Z(n38174) );
  XOR U39836 ( .A(n38176), .B(n38177), .Z(n29557) );
  AND U39837 ( .A(\modmult_1/xin[1023] ), .B(n38178), .Z(n38177) );
  IV U39838 ( .A(n38176), .Z(n38178) );
  XOR U39839 ( .A(n38179), .B(g_input[197]), .Z(n38176) );
  NAND U39840 ( .A(n38180), .B(mul_pow), .Z(n38179) );
  XOR U39841 ( .A(g_input[197]), .B(creg[197]), .Z(n38180) );
  XOR U39842 ( .A(n38181), .B(n38182), .Z(n38172) );
  ANDN U39843 ( .A(n38183), .B(n29564), .Z(n38182) );
  XOR U39844 ( .A(n38184), .B(\modmult_1/zin[0][195] ), .Z(n29564) );
  IV U39845 ( .A(n38181), .Z(n38184) );
  XNOR U39846 ( .A(n38181), .B(n29563), .Z(n38183) );
  XOR U39847 ( .A(n38185), .B(n38186), .Z(n29563) );
  AND U39848 ( .A(\modmult_1/xin[1023] ), .B(n38187), .Z(n38186) );
  IV U39849 ( .A(n38185), .Z(n38187) );
  XOR U39850 ( .A(n38188), .B(g_input[196]), .Z(n38185) );
  NAND U39851 ( .A(n38189), .B(mul_pow), .Z(n38188) );
  XOR U39852 ( .A(g_input[196]), .B(creg[196]), .Z(n38189) );
  XOR U39853 ( .A(n38190), .B(n38191), .Z(n38181) );
  ANDN U39854 ( .A(n38192), .B(n29570), .Z(n38191) );
  XOR U39855 ( .A(n38193), .B(\modmult_1/zin[0][194] ), .Z(n29570) );
  IV U39856 ( .A(n38190), .Z(n38193) );
  XNOR U39857 ( .A(n38190), .B(n29569), .Z(n38192) );
  XOR U39858 ( .A(n38194), .B(n38195), .Z(n29569) );
  AND U39859 ( .A(\modmult_1/xin[1023] ), .B(n38196), .Z(n38195) );
  IV U39860 ( .A(n38194), .Z(n38196) );
  XOR U39861 ( .A(n38197), .B(g_input[195]), .Z(n38194) );
  NAND U39862 ( .A(n38198), .B(mul_pow), .Z(n38197) );
  XOR U39863 ( .A(g_input[195]), .B(creg[195]), .Z(n38198) );
  XOR U39864 ( .A(n38199), .B(n38200), .Z(n38190) );
  ANDN U39865 ( .A(n38201), .B(n29576), .Z(n38200) );
  XOR U39866 ( .A(n38202), .B(\modmult_1/zin[0][193] ), .Z(n29576) );
  IV U39867 ( .A(n38199), .Z(n38202) );
  XNOR U39868 ( .A(n38199), .B(n29575), .Z(n38201) );
  XOR U39869 ( .A(n38203), .B(n38204), .Z(n29575) );
  AND U39870 ( .A(\modmult_1/xin[1023] ), .B(n38205), .Z(n38204) );
  IV U39871 ( .A(n38203), .Z(n38205) );
  XOR U39872 ( .A(n38206), .B(g_input[194]), .Z(n38203) );
  NAND U39873 ( .A(n38207), .B(mul_pow), .Z(n38206) );
  XOR U39874 ( .A(g_input[194]), .B(creg[194]), .Z(n38207) );
  XOR U39875 ( .A(n38208), .B(n38209), .Z(n38199) );
  ANDN U39876 ( .A(n38210), .B(n29582), .Z(n38209) );
  XOR U39877 ( .A(n38211), .B(\modmult_1/zin[0][192] ), .Z(n29582) );
  IV U39878 ( .A(n38208), .Z(n38211) );
  XNOR U39879 ( .A(n38208), .B(n29581), .Z(n38210) );
  XOR U39880 ( .A(n38212), .B(n38213), .Z(n29581) );
  AND U39881 ( .A(\modmult_1/xin[1023] ), .B(n38214), .Z(n38213) );
  IV U39882 ( .A(n38212), .Z(n38214) );
  XOR U39883 ( .A(n38215), .B(g_input[193]), .Z(n38212) );
  NAND U39884 ( .A(n38216), .B(mul_pow), .Z(n38215) );
  XOR U39885 ( .A(g_input[193]), .B(creg[193]), .Z(n38216) );
  XOR U39886 ( .A(n38217), .B(n38218), .Z(n38208) );
  ANDN U39887 ( .A(n38219), .B(n29588), .Z(n38218) );
  XOR U39888 ( .A(n38220), .B(\modmult_1/zin[0][191] ), .Z(n29588) );
  IV U39889 ( .A(n38217), .Z(n38220) );
  XNOR U39890 ( .A(n38217), .B(n29587), .Z(n38219) );
  XOR U39891 ( .A(n38221), .B(n38222), .Z(n29587) );
  AND U39892 ( .A(\modmult_1/xin[1023] ), .B(n38223), .Z(n38222) );
  IV U39893 ( .A(n38221), .Z(n38223) );
  XOR U39894 ( .A(n38224), .B(g_input[192]), .Z(n38221) );
  NAND U39895 ( .A(n38225), .B(mul_pow), .Z(n38224) );
  XOR U39896 ( .A(g_input[192]), .B(creg[192]), .Z(n38225) );
  XOR U39897 ( .A(n38226), .B(n38227), .Z(n38217) );
  ANDN U39898 ( .A(n38228), .B(n29594), .Z(n38227) );
  XOR U39899 ( .A(n38229), .B(\modmult_1/zin[0][190] ), .Z(n29594) );
  IV U39900 ( .A(n38226), .Z(n38229) );
  XNOR U39901 ( .A(n38226), .B(n29593), .Z(n38228) );
  XOR U39902 ( .A(n38230), .B(n38231), .Z(n29593) );
  AND U39903 ( .A(\modmult_1/xin[1023] ), .B(n38232), .Z(n38231) );
  IV U39904 ( .A(n38230), .Z(n38232) );
  XOR U39905 ( .A(n38233), .B(g_input[191]), .Z(n38230) );
  NAND U39906 ( .A(n38234), .B(mul_pow), .Z(n38233) );
  XOR U39907 ( .A(g_input[191]), .B(creg[191]), .Z(n38234) );
  XOR U39908 ( .A(n38235), .B(n38236), .Z(n38226) );
  ANDN U39909 ( .A(n38237), .B(n29600), .Z(n38236) );
  XOR U39910 ( .A(n38238), .B(\modmult_1/zin[0][189] ), .Z(n29600) );
  IV U39911 ( .A(n38235), .Z(n38238) );
  XNOR U39912 ( .A(n38235), .B(n29599), .Z(n38237) );
  XOR U39913 ( .A(n38239), .B(n38240), .Z(n29599) );
  AND U39914 ( .A(\modmult_1/xin[1023] ), .B(n38241), .Z(n38240) );
  IV U39915 ( .A(n38239), .Z(n38241) );
  XOR U39916 ( .A(n38242), .B(g_input[190]), .Z(n38239) );
  NAND U39917 ( .A(n38243), .B(mul_pow), .Z(n38242) );
  XOR U39918 ( .A(g_input[190]), .B(creg[190]), .Z(n38243) );
  XOR U39919 ( .A(n38244), .B(n38245), .Z(n38235) );
  ANDN U39920 ( .A(n38246), .B(n29606), .Z(n38245) );
  XOR U39921 ( .A(n38247), .B(\modmult_1/zin[0][188] ), .Z(n29606) );
  IV U39922 ( .A(n38244), .Z(n38247) );
  XNOR U39923 ( .A(n38244), .B(n29605), .Z(n38246) );
  XOR U39924 ( .A(n38248), .B(n38249), .Z(n29605) );
  AND U39925 ( .A(\modmult_1/xin[1023] ), .B(n38250), .Z(n38249) );
  IV U39926 ( .A(n38248), .Z(n38250) );
  XOR U39927 ( .A(n38251), .B(g_input[189]), .Z(n38248) );
  NAND U39928 ( .A(n38252), .B(mul_pow), .Z(n38251) );
  XOR U39929 ( .A(g_input[189]), .B(creg[189]), .Z(n38252) );
  XOR U39930 ( .A(n38253), .B(n38254), .Z(n38244) );
  ANDN U39931 ( .A(n38255), .B(n29612), .Z(n38254) );
  XOR U39932 ( .A(n38256), .B(\modmult_1/zin[0][187] ), .Z(n29612) );
  IV U39933 ( .A(n38253), .Z(n38256) );
  XNOR U39934 ( .A(n38253), .B(n29611), .Z(n38255) );
  XOR U39935 ( .A(n38257), .B(n38258), .Z(n29611) );
  AND U39936 ( .A(\modmult_1/xin[1023] ), .B(n38259), .Z(n38258) );
  IV U39937 ( .A(n38257), .Z(n38259) );
  XOR U39938 ( .A(n38260), .B(g_input[188]), .Z(n38257) );
  NAND U39939 ( .A(n38261), .B(mul_pow), .Z(n38260) );
  XOR U39940 ( .A(g_input[188]), .B(creg[188]), .Z(n38261) );
  XOR U39941 ( .A(n38262), .B(n38263), .Z(n38253) );
  ANDN U39942 ( .A(n38264), .B(n29618), .Z(n38263) );
  XOR U39943 ( .A(n38265), .B(\modmult_1/zin[0][186] ), .Z(n29618) );
  IV U39944 ( .A(n38262), .Z(n38265) );
  XNOR U39945 ( .A(n38262), .B(n29617), .Z(n38264) );
  XOR U39946 ( .A(n38266), .B(n38267), .Z(n29617) );
  AND U39947 ( .A(\modmult_1/xin[1023] ), .B(n38268), .Z(n38267) );
  IV U39948 ( .A(n38266), .Z(n38268) );
  XOR U39949 ( .A(n38269), .B(g_input[187]), .Z(n38266) );
  NAND U39950 ( .A(n38270), .B(mul_pow), .Z(n38269) );
  XOR U39951 ( .A(g_input[187]), .B(creg[187]), .Z(n38270) );
  XOR U39952 ( .A(n38271), .B(n38272), .Z(n38262) );
  ANDN U39953 ( .A(n38273), .B(n29624), .Z(n38272) );
  XOR U39954 ( .A(n38274), .B(\modmult_1/zin[0][185] ), .Z(n29624) );
  IV U39955 ( .A(n38271), .Z(n38274) );
  XNOR U39956 ( .A(n38271), .B(n29623), .Z(n38273) );
  XOR U39957 ( .A(n38275), .B(n38276), .Z(n29623) );
  AND U39958 ( .A(\modmult_1/xin[1023] ), .B(n38277), .Z(n38276) );
  IV U39959 ( .A(n38275), .Z(n38277) );
  XOR U39960 ( .A(n38278), .B(g_input[186]), .Z(n38275) );
  NAND U39961 ( .A(n38279), .B(mul_pow), .Z(n38278) );
  XOR U39962 ( .A(g_input[186]), .B(creg[186]), .Z(n38279) );
  XOR U39963 ( .A(n38280), .B(n38281), .Z(n38271) );
  ANDN U39964 ( .A(n38282), .B(n29630), .Z(n38281) );
  XOR U39965 ( .A(n38283), .B(\modmult_1/zin[0][184] ), .Z(n29630) );
  IV U39966 ( .A(n38280), .Z(n38283) );
  XNOR U39967 ( .A(n38280), .B(n29629), .Z(n38282) );
  XOR U39968 ( .A(n38284), .B(n38285), .Z(n29629) );
  AND U39969 ( .A(\modmult_1/xin[1023] ), .B(n38286), .Z(n38285) );
  IV U39970 ( .A(n38284), .Z(n38286) );
  XOR U39971 ( .A(n38287), .B(g_input[185]), .Z(n38284) );
  NAND U39972 ( .A(n38288), .B(mul_pow), .Z(n38287) );
  XOR U39973 ( .A(g_input[185]), .B(creg[185]), .Z(n38288) );
  XOR U39974 ( .A(n38289), .B(n38290), .Z(n38280) );
  ANDN U39975 ( .A(n38291), .B(n29636), .Z(n38290) );
  XOR U39976 ( .A(n38292), .B(\modmult_1/zin[0][183] ), .Z(n29636) );
  IV U39977 ( .A(n38289), .Z(n38292) );
  XNOR U39978 ( .A(n38289), .B(n29635), .Z(n38291) );
  XOR U39979 ( .A(n38293), .B(n38294), .Z(n29635) );
  AND U39980 ( .A(\modmult_1/xin[1023] ), .B(n38295), .Z(n38294) );
  IV U39981 ( .A(n38293), .Z(n38295) );
  XOR U39982 ( .A(n38296), .B(g_input[184]), .Z(n38293) );
  NAND U39983 ( .A(n38297), .B(mul_pow), .Z(n38296) );
  XOR U39984 ( .A(g_input[184]), .B(creg[184]), .Z(n38297) );
  XOR U39985 ( .A(n38298), .B(n38299), .Z(n38289) );
  ANDN U39986 ( .A(n38300), .B(n29642), .Z(n38299) );
  XOR U39987 ( .A(n38301), .B(\modmult_1/zin[0][182] ), .Z(n29642) );
  IV U39988 ( .A(n38298), .Z(n38301) );
  XNOR U39989 ( .A(n38298), .B(n29641), .Z(n38300) );
  XOR U39990 ( .A(n38302), .B(n38303), .Z(n29641) );
  AND U39991 ( .A(\modmult_1/xin[1023] ), .B(n38304), .Z(n38303) );
  IV U39992 ( .A(n38302), .Z(n38304) );
  XOR U39993 ( .A(n38305), .B(g_input[183]), .Z(n38302) );
  NAND U39994 ( .A(n38306), .B(mul_pow), .Z(n38305) );
  XOR U39995 ( .A(g_input[183]), .B(creg[183]), .Z(n38306) );
  XOR U39996 ( .A(n38307), .B(n38308), .Z(n38298) );
  ANDN U39997 ( .A(n38309), .B(n29648), .Z(n38308) );
  XOR U39998 ( .A(n38310), .B(\modmult_1/zin[0][181] ), .Z(n29648) );
  IV U39999 ( .A(n38307), .Z(n38310) );
  XNOR U40000 ( .A(n38307), .B(n29647), .Z(n38309) );
  XOR U40001 ( .A(n38311), .B(n38312), .Z(n29647) );
  AND U40002 ( .A(\modmult_1/xin[1023] ), .B(n38313), .Z(n38312) );
  IV U40003 ( .A(n38311), .Z(n38313) );
  XOR U40004 ( .A(n38314), .B(g_input[182]), .Z(n38311) );
  NAND U40005 ( .A(n38315), .B(mul_pow), .Z(n38314) );
  XOR U40006 ( .A(g_input[182]), .B(creg[182]), .Z(n38315) );
  XOR U40007 ( .A(n38316), .B(n38317), .Z(n38307) );
  ANDN U40008 ( .A(n38318), .B(n29654), .Z(n38317) );
  XOR U40009 ( .A(n38319), .B(\modmult_1/zin[0][180] ), .Z(n29654) );
  IV U40010 ( .A(n38316), .Z(n38319) );
  XNOR U40011 ( .A(n38316), .B(n29653), .Z(n38318) );
  XOR U40012 ( .A(n38320), .B(n38321), .Z(n29653) );
  AND U40013 ( .A(\modmult_1/xin[1023] ), .B(n38322), .Z(n38321) );
  IV U40014 ( .A(n38320), .Z(n38322) );
  XOR U40015 ( .A(n38323), .B(g_input[181]), .Z(n38320) );
  NAND U40016 ( .A(n38324), .B(mul_pow), .Z(n38323) );
  XOR U40017 ( .A(g_input[181]), .B(creg[181]), .Z(n38324) );
  XOR U40018 ( .A(n38325), .B(n38326), .Z(n38316) );
  ANDN U40019 ( .A(n38327), .B(n29660), .Z(n38326) );
  XOR U40020 ( .A(n38328), .B(\modmult_1/zin[0][179] ), .Z(n29660) );
  IV U40021 ( .A(n38325), .Z(n38328) );
  XNOR U40022 ( .A(n38325), .B(n29659), .Z(n38327) );
  XOR U40023 ( .A(n38329), .B(n38330), .Z(n29659) );
  AND U40024 ( .A(\modmult_1/xin[1023] ), .B(n38331), .Z(n38330) );
  IV U40025 ( .A(n38329), .Z(n38331) );
  XOR U40026 ( .A(n38332), .B(g_input[180]), .Z(n38329) );
  NAND U40027 ( .A(n38333), .B(mul_pow), .Z(n38332) );
  XOR U40028 ( .A(g_input[180]), .B(creg[180]), .Z(n38333) );
  XOR U40029 ( .A(n38334), .B(n38335), .Z(n38325) );
  ANDN U40030 ( .A(n38336), .B(n29666), .Z(n38335) );
  XOR U40031 ( .A(n38337), .B(\modmult_1/zin[0][178] ), .Z(n29666) );
  IV U40032 ( .A(n38334), .Z(n38337) );
  XNOR U40033 ( .A(n38334), .B(n29665), .Z(n38336) );
  XOR U40034 ( .A(n38338), .B(n38339), .Z(n29665) );
  AND U40035 ( .A(\modmult_1/xin[1023] ), .B(n38340), .Z(n38339) );
  IV U40036 ( .A(n38338), .Z(n38340) );
  XOR U40037 ( .A(n38341), .B(g_input[179]), .Z(n38338) );
  NAND U40038 ( .A(n38342), .B(mul_pow), .Z(n38341) );
  XOR U40039 ( .A(g_input[179]), .B(creg[179]), .Z(n38342) );
  XOR U40040 ( .A(n38343), .B(n38344), .Z(n38334) );
  ANDN U40041 ( .A(n38345), .B(n29672), .Z(n38344) );
  XOR U40042 ( .A(n38346), .B(\modmult_1/zin[0][177] ), .Z(n29672) );
  IV U40043 ( .A(n38343), .Z(n38346) );
  XNOR U40044 ( .A(n38343), .B(n29671), .Z(n38345) );
  XOR U40045 ( .A(n38347), .B(n38348), .Z(n29671) );
  AND U40046 ( .A(\modmult_1/xin[1023] ), .B(n38349), .Z(n38348) );
  IV U40047 ( .A(n38347), .Z(n38349) );
  XOR U40048 ( .A(n38350), .B(g_input[178]), .Z(n38347) );
  NAND U40049 ( .A(n38351), .B(mul_pow), .Z(n38350) );
  XOR U40050 ( .A(g_input[178]), .B(creg[178]), .Z(n38351) );
  XOR U40051 ( .A(n38352), .B(n38353), .Z(n38343) );
  ANDN U40052 ( .A(n38354), .B(n29678), .Z(n38353) );
  XOR U40053 ( .A(n38355), .B(\modmult_1/zin[0][176] ), .Z(n29678) );
  IV U40054 ( .A(n38352), .Z(n38355) );
  XNOR U40055 ( .A(n38352), .B(n29677), .Z(n38354) );
  XOR U40056 ( .A(n38356), .B(n38357), .Z(n29677) );
  AND U40057 ( .A(\modmult_1/xin[1023] ), .B(n38358), .Z(n38357) );
  IV U40058 ( .A(n38356), .Z(n38358) );
  XOR U40059 ( .A(n38359), .B(g_input[177]), .Z(n38356) );
  NAND U40060 ( .A(n38360), .B(mul_pow), .Z(n38359) );
  XOR U40061 ( .A(g_input[177]), .B(creg[177]), .Z(n38360) );
  XOR U40062 ( .A(n38361), .B(n38362), .Z(n38352) );
  ANDN U40063 ( .A(n38363), .B(n29684), .Z(n38362) );
  XOR U40064 ( .A(n38364), .B(\modmult_1/zin[0][175] ), .Z(n29684) );
  IV U40065 ( .A(n38361), .Z(n38364) );
  XNOR U40066 ( .A(n38361), .B(n29683), .Z(n38363) );
  XOR U40067 ( .A(n38365), .B(n38366), .Z(n29683) );
  AND U40068 ( .A(\modmult_1/xin[1023] ), .B(n38367), .Z(n38366) );
  IV U40069 ( .A(n38365), .Z(n38367) );
  XOR U40070 ( .A(n38368), .B(g_input[176]), .Z(n38365) );
  NAND U40071 ( .A(n38369), .B(mul_pow), .Z(n38368) );
  XOR U40072 ( .A(g_input[176]), .B(creg[176]), .Z(n38369) );
  XOR U40073 ( .A(n38370), .B(n38371), .Z(n38361) );
  ANDN U40074 ( .A(n38372), .B(n29690), .Z(n38371) );
  XOR U40075 ( .A(n38373), .B(\modmult_1/zin[0][174] ), .Z(n29690) );
  IV U40076 ( .A(n38370), .Z(n38373) );
  XNOR U40077 ( .A(n38370), .B(n29689), .Z(n38372) );
  XOR U40078 ( .A(n38374), .B(n38375), .Z(n29689) );
  AND U40079 ( .A(\modmult_1/xin[1023] ), .B(n38376), .Z(n38375) );
  IV U40080 ( .A(n38374), .Z(n38376) );
  XOR U40081 ( .A(n38377), .B(g_input[175]), .Z(n38374) );
  NAND U40082 ( .A(n38378), .B(mul_pow), .Z(n38377) );
  XOR U40083 ( .A(g_input[175]), .B(creg[175]), .Z(n38378) );
  XOR U40084 ( .A(n38379), .B(n38380), .Z(n38370) );
  ANDN U40085 ( .A(n38381), .B(n29696), .Z(n38380) );
  XOR U40086 ( .A(n38382), .B(\modmult_1/zin[0][173] ), .Z(n29696) );
  IV U40087 ( .A(n38379), .Z(n38382) );
  XNOR U40088 ( .A(n38379), .B(n29695), .Z(n38381) );
  XOR U40089 ( .A(n38383), .B(n38384), .Z(n29695) );
  AND U40090 ( .A(\modmult_1/xin[1023] ), .B(n38385), .Z(n38384) );
  IV U40091 ( .A(n38383), .Z(n38385) );
  XOR U40092 ( .A(n38386), .B(g_input[174]), .Z(n38383) );
  NAND U40093 ( .A(n38387), .B(mul_pow), .Z(n38386) );
  XOR U40094 ( .A(g_input[174]), .B(creg[174]), .Z(n38387) );
  XOR U40095 ( .A(n38388), .B(n38389), .Z(n38379) );
  ANDN U40096 ( .A(n38390), .B(n29702), .Z(n38389) );
  XOR U40097 ( .A(n38391), .B(\modmult_1/zin[0][172] ), .Z(n29702) );
  IV U40098 ( .A(n38388), .Z(n38391) );
  XNOR U40099 ( .A(n38388), .B(n29701), .Z(n38390) );
  XOR U40100 ( .A(n38392), .B(n38393), .Z(n29701) );
  AND U40101 ( .A(\modmult_1/xin[1023] ), .B(n38394), .Z(n38393) );
  IV U40102 ( .A(n38392), .Z(n38394) );
  XOR U40103 ( .A(n38395), .B(g_input[173]), .Z(n38392) );
  NAND U40104 ( .A(n38396), .B(mul_pow), .Z(n38395) );
  XOR U40105 ( .A(g_input[173]), .B(creg[173]), .Z(n38396) );
  XOR U40106 ( .A(n38397), .B(n38398), .Z(n38388) );
  ANDN U40107 ( .A(n38399), .B(n29708), .Z(n38398) );
  XOR U40108 ( .A(n38400), .B(\modmult_1/zin[0][171] ), .Z(n29708) );
  IV U40109 ( .A(n38397), .Z(n38400) );
  XNOR U40110 ( .A(n38397), .B(n29707), .Z(n38399) );
  XOR U40111 ( .A(n38401), .B(n38402), .Z(n29707) );
  AND U40112 ( .A(\modmult_1/xin[1023] ), .B(n38403), .Z(n38402) );
  IV U40113 ( .A(n38401), .Z(n38403) );
  XOR U40114 ( .A(n38404), .B(g_input[172]), .Z(n38401) );
  NAND U40115 ( .A(n38405), .B(mul_pow), .Z(n38404) );
  XOR U40116 ( .A(g_input[172]), .B(creg[172]), .Z(n38405) );
  XOR U40117 ( .A(n38406), .B(n38407), .Z(n38397) );
  ANDN U40118 ( .A(n38408), .B(n29714), .Z(n38407) );
  XOR U40119 ( .A(n38409), .B(\modmult_1/zin[0][170] ), .Z(n29714) );
  IV U40120 ( .A(n38406), .Z(n38409) );
  XNOR U40121 ( .A(n38406), .B(n29713), .Z(n38408) );
  XOR U40122 ( .A(n38410), .B(n38411), .Z(n29713) );
  AND U40123 ( .A(\modmult_1/xin[1023] ), .B(n38412), .Z(n38411) );
  IV U40124 ( .A(n38410), .Z(n38412) );
  XOR U40125 ( .A(n38413), .B(g_input[171]), .Z(n38410) );
  NAND U40126 ( .A(n38414), .B(mul_pow), .Z(n38413) );
  XOR U40127 ( .A(g_input[171]), .B(creg[171]), .Z(n38414) );
  XOR U40128 ( .A(n38415), .B(n38416), .Z(n38406) );
  ANDN U40129 ( .A(n38417), .B(n29720), .Z(n38416) );
  XOR U40130 ( .A(n38418), .B(\modmult_1/zin[0][169] ), .Z(n29720) );
  IV U40131 ( .A(n38415), .Z(n38418) );
  XNOR U40132 ( .A(n38415), .B(n29719), .Z(n38417) );
  XOR U40133 ( .A(n38419), .B(n38420), .Z(n29719) );
  AND U40134 ( .A(\modmult_1/xin[1023] ), .B(n38421), .Z(n38420) );
  IV U40135 ( .A(n38419), .Z(n38421) );
  XOR U40136 ( .A(n38422), .B(g_input[170]), .Z(n38419) );
  NAND U40137 ( .A(n38423), .B(mul_pow), .Z(n38422) );
  XOR U40138 ( .A(g_input[170]), .B(creg[170]), .Z(n38423) );
  XOR U40139 ( .A(n38424), .B(n38425), .Z(n38415) );
  ANDN U40140 ( .A(n38426), .B(n29726), .Z(n38425) );
  XOR U40141 ( .A(n38427), .B(\modmult_1/zin[0][168] ), .Z(n29726) );
  IV U40142 ( .A(n38424), .Z(n38427) );
  XNOR U40143 ( .A(n38424), .B(n29725), .Z(n38426) );
  XOR U40144 ( .A(n38428), .B(n38429), .Z(n29725) );
  AND U40145 ( .A(\modmult_1/xin[1023] ), .B(n38430), .Z(n38429) );
  IV U40146 ( .A(n38428), .Z(n38430) );
  XOR U40147 ( .A(n38431), .B(g_input[169]), .Z(n38428) );
  NAND U40148 ( .A(n38432), .B(mul_pow), .Z(n38431) );
  XOR U40149 ( .A(g_input[169]), .B(creg[169]), .Z(n38432) );
  XOR U40150 ( .A(n38433), .B(n38434), .Z(n38424) );
  ANDN U40151 ( .A(n38435), .B(n29732), .Z(n38434) );
  XOR U40152 ( .A(n38436), .B(\modmult_1/zin[0][167] ), .Z(n29732) );
  IV U40153 ( .A(n38433), .Z(n38436) );
  XNOR U40154 ( .A(n38433), .B(n29731), .Z(n38435) );
  XOR U40155 ( .A(n38437), .B(n38438), .Z(n29731) );
  AND U40156 ( .A(\modmult_1/xin[1023] ), .B(n38439), .Z(n38438) );
  IV U40157 ( .A(n38437), .Z(n38439) );
  XOR U40158 ( .A(n38440), .B(g_input[168]), .Z(n38437) );
  NAND U40159 ( .A(n38441), .B(mul_pow), .Z(n38440) );
  XOR U40160 ( .A(g_input[168]), .B(creg[168]), .Z(n38441) );
  XOR U40161 ( .A(n38442), .B(n38443), .Z(n38433) );
  ANDN U40162 ( .A(n38444), .B(n29738), .Z(n38443) );
  XOR U40163 ( .A(n38445), .B(\modmult_1/zin[0][166] ), .Z(n29738) );
  IV U40164 ( .A(n38442), .Z(n38445) );
  XNOR U40165 ( .A(n38442), .B(n29737), .Z(n38444) );
  XOR U40166 ( .A(n38446), .B(n38447), .Z(n29737) );
  AND U40167 ( .A(\modmult_1/xin[1023] ), .B(n38448), .Z(n38447) );
  IV U40168 ( .A(n38446), .Z(n38448) );
  XOR U40169 ( .A(n38449), .B(g_input[167]), .Z(n38446) );
  NAND U40170 ( .A(n38450), .B(mul_pow), .Z(n38449) );
  XOR U40171 ( .A(g_input[167]), .B(creg[167]), .Z(n38450) );
  XOR U40172 ( .A(n38451), .B(n38452), .Z(n38442) );
  ANDN U40173 ( .A(n38453), .B(n29744), .Z(n38452) );
  XOR U40174 ( .A(n38454), .B(\modmult_1/zin[0][165] ), .Z(n29744) );
  IV U40175 ( .A(n38451), .Z(n38454) );
  XNOR U40176 ( .A(n38451), .B(n29743), .Z(n38453) );
  XOR U40177 ( .A(n38455), .B(n38456), .Z(n29743) );
  AND U40178 ( .A(\modmult_1/xin[1023] ), .B(n38457), .Z(n38456) );
  IV U40179 ( .A(n38455), .Z(n38457) );
  XOR U40180 ( .A(n38458), .B(g_input[166]), .Z(n38455) );
  NAND U40181 ( .A(n38459), .B(mul_pow), .Z(n38458) );
  XOR U40182 ( .A(g_input[166]), .B(creg[166]), .Z(n38459) );
  XOR U40183 ( .A(n38460), .B(n38461), .Z(n38451) );
  ANDN U40184 ( .A(n38462), .B(n29750), .Z(n38461) );
  XOR U40185 ( .A(n38463), .B(\modmult_1/zin[0][164] ), .Z(n29750) );
  IV U40186 ( .A(n38460), .Z(n38463) );
  XNOR U40187 ( .A(n38460), .B(n29749), .Z(n38462) );
  XOR U40188 ( .A(n38464), .B(n38465), .Z(n29749) );
  AND U40189 ( .A(\modmult_1/xin[1023] ), .B(n38466), .Z(n38465) );
  IV U40190 ( .A(n38464), .Z(n38466) );
  XOR U40191 ( .A(n38467), .B(g_input[165]), .Z(n38464) );
  NAND U40192 ( .A(n38468), .B(mul_pow), .Z(n38467) );
  XOR U40193 ( .A(g_input[165]), .B(creg[165]), .Z(n38468) );
  XOR U40194 ( .A(n38469), .B(n38470), .Z(n38460) );
  ANDN U40195 ( .A(n38471), .B(n29756), .Z(n38470) );
  XOR U40196 ( .A(n38472), .B(\modmult_1/zin[0][163] ), .Z(n29756) );
  IV U40197 ( .A(n38469), .Z(n38472) );
  XNOR U40198 ( .A(n38469), .B(n29755), .Z(n38471) );
  XOR U40199 ( .A(n38473), .B(n38474), .Z(n29755) );
  AND U40200 ( .A(\modmult_1/xin[1023] ), .B(n38475), .Z(n38474) );
  IV U40201 ( .A(n38473), .Z(n38475) );
  XOR U40202 ( .A(n38476), .B(g_input[164]), .Z(n38473) );
  NAND U40203 ( .A(n38477), .B(mul_pow), .Z(n38476) );
  XOR U40204 ( .A(g_input[164]), .B(creg[164]), .Z(n38477) );
  XOR U40205 ( .A(n38478), .B(n38479), .Z(n38469) );
  ANDN U40206 ( .A(n38480), .B(n29762), .Z(n38479) );
  XOR U40207 ( .A(n38481), .B(\modmult_1/zin[0][162] ), .Z(n29762) );
  IV U40208 ( .A(n38478), .Z(n38481) );
  XNOR U40209 ( .A(n38478), .B(n29761), .Z(n38480) );
  XOR U40210 ( .A(n38482), .B(n38483), .Z(n29761) );
  AND U40211 ( .A(\modmult_1/xin[1023] ), .B(n38484), .Z(n38483) );
  IV U40212 ( .A(n38482), .Z(n38484) );
  XOR U40213 ( .A(n38485), .B(g_input[163]), .Z(n38482) );
  NAND U40214 ( .A(n38486), .B(mul_pow), .Z(n38485) );
  XOR U40215 ( .A(g_input[163]), .B(creg[163]), .Z(n38486) );
  XOR U40216 ( .A(n38487), .B(n38488), .Z(n38478) );
  ANDN U40217 ( .A(n38489), .B(n29768), .Z(n38488) );
  XOR U40218 ( .A(n38490), .B(\modmult_1/zin[0][161] ), .Z(n29768) );
  IV U40219 ( .A(n38487), .Z(n38490) );
  XNOR U40220 ( .A(n38487), .B(n29767), .Z(n38489) );
  XOR U40221 ( .A(n38491), .B(n38492), .Z(n29767) );
  AND U40222 ( .A(\modmult_1/xin[1023] ), .B(n38493), .Z(n38492) );
  IV U40223 ( .A(n38491), .Z(n38493) );
  XOR U40224 ( .A(n38494), .B(g_input[162]), .Z(n38491) );
  NAND U40225 ( .A(n38495), .B(mul_pow), .Z(n38494) );
  XOR U40226 ( .A(g_input[162]), .B(creg[162]), .Z(n38495) );
  XOR U40227 ( .A(n38496), .B(n38497), .Z(n38487) );
  ANDN U40228 ( .A(n38498), .B(n29774), .Z(n38497) );
  XOR U40229 ( .A(n38499), .B(\modmult_1/zin[0][160] ), .Z(n29774) );
  IV U40230 ( .A(n38496), .Z(n38499) );
  XNOR U40231 ( .A(n38496), .B(n29773), .Z(n38498) );
  XOR U40232 ( .A(n38500), .B(n38501), .Z(n29773) );
  AND U40233 ( .A(\modmult_1/xin[1023] ), .B(n38502), .Z(n38501) );
  IV U40234 ( .A(n38500), .Z(n38502) );
  XOR U40235 ( .A(n38503), .B(g_input[161]), .Z(n38500) );
  NAND U40236 ( .A(n38504), .B(mul_pow), .Z(n38503) );
  XOR U40237 ( .A(g_input[161]), .B(creg[161]), .Z(n38504) );
  XOR U40238 ( .A(n38505), .B(n38506), .Z(n38496) );
  ANDN U40239 ( .A(n38507), .B(n29780), .Z(n38506) );
  XOR U40240 ( .A(n38508), .B(\modmult_1/zin[0][159] ), .Z(n29780) );
  IV U40241 ( .A(n38505), .Z(n38508) );
  XNOR U40242 ( .A(n38505), .B(n29779), .Z(n38507) );
  XOR U40243 ( .A(n38509), .B(n38510), .Z(n29779) );
  AND U40244 ( .A(\modmult_1/xin[1023] ), .B(n38511), .Z(n38510) );
  IV U40245 ( .A(n38509), .Z(n38511) );
  XOR U40246 ( .A(n38512), .B(g_input[160]), .Z(n38509) );
  NAND U40247 ( .A(n38513), .B(mul_pow), .Z(n38512) );
  XOR U40248 ( .A(g_input[160]), .B(creg[160]), .Z(n38513) );
  XOR U40249 ( .A(n38514), .B(n38515), .Z(n38505) );
  ANDN U40250 ( .A(n38516), .B(n29786), .Z(n38515) );
  XOR U40251 ( .A(n38517), .B(\modmult_1/zin[0][158] ), .Z(n29786) );
  IV U40252 ( .A(n38514), .Z(n38517) );
  XNOR U40253 ( .A(n38514), .B(n29785), .Z(n38516) );
  XOR U40254 ( .A(n38518), .B(n38519), .Z(n29785) );
  AND U40255 ( .A(\modmult_1/xin[1023] ), .B(n38520), .Z(n38519) );
  IV U40256 ( .A(n38518), .Z(n38520) );
  XOR U40257 ( .A(n38521), .B(g_input[159]), .Z(n38518) );
  NAND U40258 ( .A(n38522), .B(mul_pow), .Z(n38521) );
  XOR U40259 ( .A(g_input[159]), .B(creg[159]), .Z(n38522) );
  XOR U40260 ( .A(n38523), .B(n38524), .Z(n38514) );
  ANDN U40261 ( .A(n38525), .B(n29792), .Z(n38524) );
  XOR U40262 ( .A(n38526), .B(\modmult_1/zin[0][157] ), .Z(n29792) );
  IV U40263 ( .A(n38523), .Z(n38526) );
  XNOR U40264 ( .A(n38523), .B(n29791), .Z(n38525) );
  XOR U40265 ( .A(n38527), .B(n38528), .Z(n29791) );
  AND U40266 ( .A(\modmult_1/xin[1023] ), .B(n38529), .Z(n38528) );
  IV U40267 ( .A(n38527), .Z(n38529) );
  XOR U40268 ( .A(n38530), .B(g_input[158]), .Z(n38527) );
  NAND U40269 ( .A(n38531), .B(mul_pow), .Z(n38530) );
  XOR U40270 ( .A(g_input[158]), .B(creg[158]), .Z(n38531) );
  XOR U40271 ( .A(n38532), .B(n38533), .Z(n38523) );
  ANDN U40272 ( .A(n38534), .B(n29798), .Z(n38533) );
  XOR U40273 ( .A(n38535), .B(\modmult_1/zin[0][156] ), .Z(n29798) );
  IV U40274 ( .A(n38532), .Z(n38535) );
  XNOR U40275 ( .A(n38532), .B(n29797), .Z(n38534) );
  XOR U40276 ( .A(n38536), .B(n38537), .Z(n29797) );
  AND U40277 ( .A(\modmult_1/xin[1023] ), .B(n38538), .Z(n38537) );
  IV U40278 ( .A(n38536), .Z(n38538) );
  XOR U40279 ( .A(n38539), .B(g_input[157]), .Z(n38536) );
  NAND U40280 ( .A(n38540), .B(mul_pow), .Z(n38539) );
  XOR U40281 ( .A(g_input[157]), .B(creg[157]), .Z(n38540) );
  XOR U40282 ( .A(n38541), .B(n38542), .Z(n38532) );
  ANDN U40283 ( .A(n38543), .B(n29804), .Z(n38542) );
  XOR U40284 ( .A(n38544), .B(\modmult_1/zin[0][155] ), .Z(n29804) );
  IV U40285 ( .A(n38541), .Z(n38544) );
  XNOR U40286 ( .A(n38541), .B(n29803), .Z(n38543) );
  XOR U40287 ( .A(n38545), .B(n38546), .Z(n29803) );
  AND U40288 ( .A(\modmult_1/xin[1023] ), .B(n38547), .Z(n38546) );
  IV U40289 ( .A(n38545), .Z(n38547) );
  XOR U40290 ( .A(n38548), .B(g_input[156]), .Z(n38545) );
  NAND U40291 ( .A(n38549), .B(mul_pow), .Z(n38548) );
  XOR U40292 ( .A(g_input[156]), .B(creg[156]), .Z(n38549) );
  XOR U40293 ( .A(n38550), .B(n38551), .Z(n38541) );
  ANDN U40294 ( .A(n38552), .B(n29810), .Z(n38551) );
  XOR U40295 ( .A(n38553), .B(\modmult_1/zin[0][154] ), .Z(n29810) );
  IV U40296 ( .A(n38550), .Z(n38553) );
  XNOR U40297 ( .A(n38550), .B(n29809), .Z(n38552) );
  XOR U40298 ( .A(n38554), .B(n38555), .Z(n29809) );
  AND U40299 ( .A(\modmult_1/xin[1023] ), .B(n38556), .Z(n38555) );
  IV U40300 ( .A(n38554), .Z(n38556) );
  XOR U40301 ( .A(n38557), .B(g_input[155]), .Z(n38554) );
  NAND U40302 ( .A(n38558), .B(mul_pow), .Z(n38557) );
  XOR U40303 ( .A(g_input[155]), .B(creg[155]), .Z(n38558) );
  XOR U40304 ( .A(n38559), .B(n38560), .Z(n38550) );
  ANDN U40305 ( .A(n38561), .B(n29816), .Z(n38560) );
  XOR U40306 ( .A(n38562), .B(\modmult_1/zin[0][153] ), .Z(n29816) );
  IV U40307 ( .A(n38559), .Z(n38562) );
  XNOR U40308 ( .A(n38559), .B(n29815), .Z(n38561) );
  XOR U40309 ( .A(n38563), .B(n38564), .Z(n29815) );
  AND U40310 ( .A(\modmult_1/xin[1023] ), .B(n38565), .Z(n38564) );
  IV U40311 ( .A(n38563), .Z(n38565) );
  XOR U40312 ( .A(n38566), .B(g_input[154]), .Z(n38563) );
  NAND U40313 ( .A(n38567), .B(mul_pow), .Z(n38566) );
  XOR U40314 ( .A(g_input[154]), .B(creg[154]), .Z(n38567) );
  XOR U40315 ( .A(n38568), .B(n38569), .Z(n38559) );
  ANDN U40316 ( .A(n38570), .B(n29822), .Z(n38569) );
  XOR U40317 ( .A(n38571), .B(\modmult_1/zin[0][152] ), .Z(n29822) );
  IV U40318 ( .A(n38568), .Z(n38571) );
  XNOR U40319 ( .A(n38568), .B(n29821), .Z(n38570) );
  XOR U40320 ( .A(n38572), .B(n38573), .Z(n29821) );
  AND U40321 ( .A(\modmult_1/xin[1023] ), .B(n38574), .Z(n38573) );
  IV U40322 ( .A(n38572), .Z(n38574) );
  XOR U40323 ( .A(n38575), .B(g_input[153]), .Z(n38572) );
  NAND U40324 ( .A(n38576), .B(mul_pow), .Z(n38575) );
  XOR U40325 ( .A(g_input[153]), .B(creg[153]), .Z(n38576) );
  XOR U40326 ( .A(n38577), .B(n38578), .Z(n38568) );
  ANDN U40327 ( .A(n38579), .B(n29828), .Z(n38578) );
  XOR U40328 ( .A(n38580), .B(\modmult_1/zin[0][151] ), .Z(n29828) );
  IV U40329 ( .A(n38577), .Z(n38580) );
  XNOR U40330 ( .A(n38577), .B(n29827), .Z(n38579) );
  XOR U40331 ( .A(n38581), .B(n38582), .Z(n29827) );
  AND U40332 ( .A(\modmult_1/xin[1023] ), .B(n38583), .Z(n38582) );
  IV U40333 ( .A(n38581), .Z(n38583) );
  XOR U40334 ( .A(n38584), .B(g_input[152]), .Z(n38581) );
  NAND U40335 ( .A(n38585), .B(mul_pow), .Z(n38584) );
  XOR U40336 ( .A(g_input[152]), .B(creg[152]), .Z(n38585) );
  XOR U40337 ( .A(n38586), .B(n38587), .Z(n38577) );
  ANDN U40338 ( .A(n38588), .B(n29834), .Z(n38587) );
  XOR U40339 ( .A(n38589), .B(\modmult_1/zin[0][150] ), .Z(n29834) );
  IV U40340 ( .A(n38586), .Z(n38589) );
  XNOR U40341 ( .A(n38586), .B(n29833), .Z(n38588) );
  XOR U40342 ( .A(n38590), .B(n38591), .Z(n29833) );
  AND U40343 ( .A(\modmult_1/xin[1023] ), .B(n38592), .Z(n38591) );
  IV U40344 ( .A(n38590), .Z(n38592) );
  XOR U40345 ( .A(n38593), .B(g_input[151]), .Z(n38590) );
  NAND U40346 ( .A(n38594), .B(mul_pow), .Z(n38593) );
  XOR U40347 ( .A(g_input[151]), .B(creg[151]), .Z(n38594) );
  XOR U40348 ( .A(n38595), .B(n38596), .Z(n38586) );
  ANDN U40349 ( .A(n38597), .B(n29840), .Z(n38596) );
  XOR U40350 ( .A(n38598), .B(\modmult_1/zin[0][149] ), .Z(n29840) );
  IV U40351 ( .A(n38595), .Z(n38598) );
  XNOR U40352 ( .A(n38595), .B(n29839), .Z(n38597) );
  XOR U40353 ( .A(n38599), .B(n38600), .Z(n29839) );
  AND U40354 ( .A(\modmult_1/xin[1023] ), .B(n38601), .Z(n38600) );
  IV U40355 ( .A(n38599), .Z(n38601) );
  XOR U40356 ( .A(n38602), .B(g_input[150]), .Z(n38599) );
  NAND U40357 ( .A(n38603), .B(mul_pow), .Z(n38602) );
  XOR U40358 ( .A(g_input[150]), .B(creg[150]), .Z(n38603) );
  XOR U40359 ( .A(n38604), .B(n38605), .Z(n38595) );
  ANDN U40360 ( .A(n38606), .B(n29846), .Z(n38605) );
  XOR U40361 ( .A(n38607), .B(\modmult_1/zin[0][148] ), .Z(n29846) );
  IV U40362 ( .A(n38604), .Z(n38607) );
  XNOR U40363 ( .A(n38604), .B(n29845), .Z(n38606) );
  XOR U40364 ( .A(n38608), .B(n38609), .Z(n29845) );
  AND U40365 ( .A(\modmult_1/xin[1023] ), .B(n38610), .Z(n38609) );
  IV U40366 ( .A(n38608), .Z(n38610) );
  XOR U40367 ( .A(n38611), .B(g_input[149]), .Z(n38608) );
  NAND U40368 ( .A(n38612), .B(mul_pow), .Z(n38611) );
  XOR U40369 ( .A(g_input[149]), .B(creg[149]), .Z(n38612) );
  XOR U40370 ( .A(n38613), .B(n38614), .Z(n38604) );
  ANDN U40371 ( .A(n38615), .B(n29852), .Z(n38614) );
  XOR U40372 ( .A(n38616), .B(\modmult_1/zin[0][147] ), .Z(n29852) );
  IV U40373 ( .A(n38613), .Z(n38616) );
  XNOR U40374 ( .A(n38613), .B(n29851), .Z(n38615) );
  XOR U40375 ( .A(n38617), .B(n38618), .Z(n29851) );
  AND U40376 ( .A(\modmult_1/xin[1023] ), .B(n38619), .Z(n38618) );
  IV U40377 ( .A(n38617), .Z(n38619) );
  XOR U40378 ( .A(n38620), .B(g_input[148]), .Z(n38617) );
  NAND U40379 ( .A(n38621), .B(mul_pow), .Z(n38620) );
  XOR U40380 ( .A(g_input[148]), .B(creg[148]), .Z(n38621) );
  XOR U40381 ( .A(n38622), .B(n38623), .Z(n38613) );
  ANDN U40382 ( .A(n38624), .B(n29858), .Z(n38623) );
  XOR U40383 ( .A(n38625), .B(\modmult_1/zin[0][146] ), .Z(n29858) );
  IV U40384 ( .A(n38622), .Z(n38625) );
  XNOR U40385 ( .A(n38622), .B(n29857), .Z(n38624) );
  XOR U40386 ( .A(n38626), .B(n38627), .Z(n29857) );
  AND U40387 ( .A(\modmult_1/xin[1023] ), .B(n38628), .Z(n38627) );
  IV U40388 ( .A(n38626), .Z(n38628) );
  XOR U40389 ( .A(n38629), .B(g_input[147]), .Z(n38626) );
  NAND U40390 ( .A(n38630), .B(mul_pow), .Z(n38629) );
  XOR U40391 ( .A(g_input[147]), .B(creg[147]), .Z(n38630) );
  XOR U40392 ( .A(n38631), .B(n38632), .Z(n38622) );
  ANDN U40393 ( .A(n38633), .B(n29864), .Z(n38632) );
  XOR U40394 ( .A(n38634), .B(\modmult_1/zin[0][145] ), .Z(n29864) );
  IV U40395 ( .A(n38631), .Z(n38634) );
  XNOR U40396 ( .A(n38631), .B(n29863), .Z(n38633) );
  XOR U40397 ( .A(n38635), .B(n38636), .Z(n29863) );
  AND U40398 ( .A(\modmult_1/xin[1023] ), .B(n38637), .Z(n38636) );
  IV U40399 ( .A(n38635), .Z(n38637) );
  XOR U40400 ( .A(n38638), .B(g_input[146]), .Z(n38635) );
  NAND U40401 ( .A(n38639), .B(mul_pow), .Z(n38638) );
  XOR U40402 ( .A(g_input[146]), .B(creg[146]), .Z(n38639) );
  XOR U40403 ( .A(n38640), .B(n38641), .Z(n38631) );
  ANDN U40404 ( .A(n38642), .B(n29870), .Z(n38641) );
  XOR U40405 ( .A(n38643), .B(\modmult_1/zin[0][144] ), .Z(n29870) );
  IV U40406 ( .A(n38640), .Z(n38643) );
  XNOR U40407 ( .A(n38640), .B(n29869), .Z(n38642) );
  XOR U40408 ( .A(n38644), .B(n38645), .Z(n29869) );
  AND U40409 ( .A(\modmult_1/xin[1023] ), .B(n38646), .Z(n38645) );
  IV U40410 ( .A(n38644), .Z(n38646) );
  XOR U40411 ( .A(n38647), .B(g_input[145]), .Z(n38644) );
  NAND U40412 ( .A(n38648), .B(mul_pow), .Z(n38647) );
  XOR U40413 ( .A(g_input[145]), .B(creg[145]), .Z(n38648) );
  XOR U40414 ( .A(n38649), .B(n38650), .Z(n38640) );
  ANDN U40415 ( .A(n38651), .B(n29876), .Z(n38650) );
  XOR U40416 ( .A(n38652), .B(\modmult_1/zin[0][143] ), .Z(n29876) );
  IV U40417 ( .A(n38649), .Z(n38652) );
  XNOR U40418 ( .A(n38649), .B(n29875), .Z(n38651) );
  XOR U40419 ( .A(n38653), .B(n38654), .Z(n29875) );
  AND U40420 ( .A(\modmult_1/xin[1023] ), .B(n38655), .Z(n38654) );
  IV U40421 ( .A(n38653), .Z(n38655) );
  XOR U40422 ( .A(n38656), .B(g_input[144]), .Z(n38653) );
  NAND U40423 ( .A(n38657), .B(mul_pow), .Z(n38656) );
  XOR U40424 ( .A(g_input[144]), .B(creg[144]), .Z(n38657) );
  XOR U40425 ( .A(n38658), .B(n38659), .Z(n38649) );
  ANDN U40426 ( .A(n38660), .B(n29882), .Z(n38659) );
  XOR U40427 ( .A(n38661), .B(\modmult_1/zin[0][142] ), .Z(n29882) );
  IV U40428 ( .A(n38658), .Z(n38661) );
  XNOR U40429 ( .A(n38658), .B(n29881), .Z(n38660) );
  XOR U40430 ( .A(n38662), .B(n38663), .Z(n29881) );
  AND U40431 ( .A(\modmult_1/xin[1023] ), .B(n38664), .Z(n38663) );
  IV U40432 ( .A(n38662), .Z(n38664) );
  XOR U40433 ( .A(n38665), .B(g_input[143]), .Z(n38662) );
  NAND U40434 ( .A(n38666), .B(mul_pow), .Z(n38665) );
  XOR U40435 ( .A(g_input[143]), .B(creg[143]), .Z(n38666) );
  XOR U40436 ( .A(n38667), .B(n38668), .Z(n38658) );
  ANDN U40437 ( .A(n38669), .B(n29888), .Z(n38668) );
  XOR U40438 ( .A(n38670), .B(\modmult_1/zin[0][141] ), .Z(n29888) );
  IV U40439 ( .A(n38667), .Z(n38670) );
  XNOR U40440 ( .A(n38667), .B(n29887), .Z(n38669) );
  XOR U40441 ( .A(n38671), .B(n38672), .Z(n29887) );
  AND U40442 ( .A(\modmult_1/xin[1023] ), .B(n38673), .Z(n38672) );
  IV U40443 ( .A(n38671), .Z(n38673) );
  XOR U40444 ( .A(n38674), .B(g_input[142]), .Z(n38671) );
  NAND U40445 ( .A(n38675), .B(mul_pow), .Z(n38674) );
  XOR U40446 ( .A(g_input[142]), .B(creg[142]), .Z(n38675) );
  XOR U40447 ( .A(n38676), .B(n38677), .Z(n38667) );
  ANDN U40448 ( .A(n38678), .B(n29894), .Z(n38677) );
  XOR U40449 ( .A(n38679), .B(\modmult_1/zin[0][140] ), .Z(n29894) );
  IV U40450 ( .A(n38676), .Z(n38679) );
  XNOR U40451 ( .A(n38676), .B(n29893), .Z(n38678) );
  XOR U40452 ( .A(n38680), .B(n38681), .Z(n29893) );
  AND U40453 ( .A(\modmult_1/xin[1023] ), .B(n38682), .Z(n38681) );
  IV U40454 ( .A(n38680), .Z(n38682) );
  XOR U40455 ( .A(n38683), .B(g_input[141]), .Z(n38680) );
  NAND U40456 ( .A(n38684), .B(mul_pow), .Z(n38683) );
  XOR U40457 ( .A(g_input[141]), .B(creg[141]), .Z(n38684) );
  XOR U40458 ( .A(n38685), .B(n38686), .Z(n38676) );
  ANDN U40459 ( .A(n38687), .B(n29900), .Z(n38686) );
  XOR U40460 ( .A(n38688), .B(\modmult_1/zin[0][139] ), .Z(n29900) );
  IV U40461 ( .A(n38685), .Z(n38688) );
  XNOR U40462 ( .A(n38685), .B(n29899), .Z(n38687) );
  XOR U40463 ( .A(n38689), .B(n38690), .Z(n29899) );
  AND U40464 ( .A(\modmult_1/xin[1023] ), .B(n38691), .Z(n38690) );
  IV U40465 ( .A(n38689), .Z(n38691) );
  XOR U40466 ( .A(n38692), .B(g_input[140]), .Z(n38689) );
  NAND U40467 ( .A(n38693), .B(mul_pow), .Z(n38692) );
  XOR U40468 ( .A(g_input[140]), .B(creg[140]), .Z(n38693) );
  XOR U40469 ( .A(n38694), .B(n38695), .Z(n38685) );
  ANDN U40470 ( .A(n38696), .B(n29906), .Z(n38695) );
  XOR U40471 ( .A(n38697), .B(\modmult_1/zin[0][138] ), .Z(n29906) );
  IV U40472 ( .A(n38694), .Z(n38697) );
  XNOR U40473 ( .A(n38694), .B(n29905), .Z(n38696) );
  XOR U40474 ( .A(n38698), .B(n38699), .Z(n29905) );
  AND U40475 ( .A(\modmult_1/xin[1023] ), .B(n38700), .Z(n38699) );
  IV U40476 ( .A(n38698), .Z(n38700) );
  XOR U40477 ( .A(n38701), .B(g_input[139]), .Z(n38698) );
  NAND U40478 ( .A(n38702), .B(mul_pow), .Z(n38701) );
  XOR U40479 ( .A(g_input[139]), .B(creg[139]), .Z(n38702) );
  XOR U40480 ( .A(n38703), .B(n38704), .Z(n38694) );
  ANDN U40481 ( .A(n38705), .B(n29912), .Z(n38704) );
  XOR U40482 ( .A(n38706), .B(\modmult_1/zin[0][137] ), .Z(n29912) );
  IV U40483 ( .A(n38703), .Z(n38706) );
  XNOR U40484 ( .A(n38703), .B(n29911), .Z(n38705) );
  XOR U40485 ( .A(n38707), .B(n38708), .Z(n29911) );
  AND U40486 ( .A(\modmult_1/xin[1023] ), .B(n38709), .Z(n38708) );
  IV U40487 ( .A(n38707), .Z(n38709) );
  XOR U40488 ( .A(n38710), .B(g_input[138]), .Z(n38707) );
  NAND U40489 ( .A(n38711), .B(mul_pow), .Z(n38710) );
  XOR U40490 ( .A(g_input[138]), .B(creg[138]), .Z(n38711) );
  XOR U40491 ( .A(n38712), .B(n38713), .Z(n38703) );
  ANDN U40492 ( .A(n38714), .B(n29918), .Z(n38713) );
  XOR U40493 ( .A(n38715), .B(\modmult_1/zin[0][136] ), .Z(n29918) );
  IV U40494 ( .A(n38712), .Z(n38715) );
  XNOR U40495 ( .A(n38712), .B(n29917), .Z(n38714) );
  XOR U40496 ( .A(n38716), .B(n38717), .Z(n29917) );
  AND U40497 ( .A(\modmult_1/xin[1023] ), .B(n38718), .Z(n38717) );
  IV U40498 ( .A(n38716), .Z(n38718) );
  XOR U40499 ( .A(n38719), .B(g_input[137]), .Z(n38716) );
  NAND U40500 ( .A(n38720), .B(mul_pow), .Z(n38719) );
  XOR U40501 ( .A(g_input[137]), .B(creg[137]), .Z(n38720) );
  XOR U40502 ( .A(n38721), .B(n38722), .Z(n38712) );
  ANDN U40503 ( .A(n38723), .B(n29924), .Z(n38722) );
  XOR U40504 ( .A(n38724), .B(\modmult_1/zin[0][135] ), .Z(n29924) );
  IV U40505 ( .A(n38721), .Z(n38724) );
  XNOR U40506 ( .A(n38721), .B(n29923), .Z(n38723) );
  XOR U40507 ( .A(n38725), .B(n38726), .Z(n29923) );
  AND U40508 ( .A(\modmult_1/xin[1023] ), .B(n38727), .Z(n38726) );
  IV U40509 ( .A(n38725), .Z(n38727) );
  XOR U40510 ( .A(n38728), .B(g_input[136]), .Z(n38725) );
  NAND U40511 ( .A(n38729), .B(mul_pow), .Z(n38728) );
  XOR U40512 ( .A(g_input[136]), .B(creg[136]), .Z(n38729) );
  XOR U40513 ( .A(n38730), .B(n38731), .Z(n38721) );
  ANDN U40514 ( .A(n38732), .B(n29930), .Z(n38731) );
  XOR U40515 ( .A(n38733), .B(\modmult_1/zin[0][134] ), .Z(n29930) );
  IV U40516 ( .A(n38730), .Z(n38733) );
  XNOR U40517 ( .A(n38730), .B(n29929), .Z(n38732) );
  XOR U40518 ( .A(n38734), .B(n38735), .Z(n29929) );
  AND U40519 ( .A(\modmult_1/xin[1023] ), .B(n38736), .Z(n38735) );
  IV U40520 ( .A(n38734), .Z(n38736) );
  XOR U40521 ( .A(n38737), .B(g_input[135]), .Z(n38734) );
  NAND U40522 ( .A(n38738), .B(mul_pow), .Z(n38737) );
  XOR U40523 ( .A(g_input[135]), .B(creg[135]), .Z(n38738) );
  XOR U40524 ( .A(n38739), .B(n38740), .Z(n38730) );
  ANDN U40525 ( .A(n38741), .B(n29936), .Z(n38740) );
  XOR U40526 ( .A(n38742), .B(\modmult_1/zin[0][133] ), .Z(n29936) );
  IV U40527 ( .A(n38739), .Z(n38742) );
  XNOR U40528 ( .A(n38739), .B(n29935), .Z(n38741) );
  XOR U40529 ( .A(n38743), .B(n38744), .Z(n29935) );
  AND U40530 ( .A(\modmult_1/xin[1023] ), .B(n38745), .Z(n38744) );
  IV U40531 ( .A(n38743), .Z(n38745) );
  XOR U40532 ( .A(n38746), .B(g_input[134]), .Z(n38743) );
  NAND U40533 ( .A(n38747), .B(mul_pow), .Z(n38746) );
  XOR U40534 ( .A(g_input[134]), .B(creg[134]), .Z(n38747) );
  XOR U40535 ( .A(n38748), .B(n38749), .Z(n38739) );
  ANDN U40536 ( .A(n38750), .B(n29942), .Z(n38749) );
  XOR U40537 ( .A(n38751), .B(\modmult_1/zin[0][132] ), .Z(n29942) );
  IV U40538 ( .A(n38748), .Z(n38751) );
  XNOR U40539 ( .A(n38748), .B(n29941), .Z(n38750) );
  XOR U40540 ( .A(n38752), .B(n38753), .Z(n29941) );
  AND U40541 ( .A(\modmult_1/xin[1023] ), .B(n38754), .Z(n38753) );
  IV U40542 ( .A(n38752), .Z(n38754) );
  XOR U40543 ( .A(n38755), .B(g_input[133]), .Z(n38752) );
  NAND U40544 ( .A(n38756), .B(mul_pow), .Z(n38755) );
  XOR U40545 ( .A(g_input[133]), .B(creg[133]), .Z(n38756) );
  XOR U40546 ( .A(n38757), .B(n38758), .Z(n38748) );
  ANDN U40547 ( .A(n38759), .B(n29948), .Z(n38758) );
  XOR U40548 ( .A(n38760), .B(\modmult_1/zin[0][131] ), .Z(n29948) );
  IV U40549 ( .A(n38757), .Z(n38760) );
  XNOR U40550 ( .A(n38757), .B(n29947), .Z(n38759) );
  XOR U40551 ( .A(n38761), .B(n38762), .Z(n29947) );
  AND U40552 ( .A(\modmult_1/xin[1023] ), .B(n38763), .Z(n38762) );
  IV U40553 ( .A(n38761), .Z(n38763) );
  XOR U40554 ( .A(n38764), .B(g_input[132]), .Z(n38761) );
  NAND U40555 ( .A(n38765), .B(mul_pow), .Z(n38764) );
  XOR U40556 ( .A(g_input[132]), .B(creg[132]), .Z(n38765) );
  XOR U40557 ( .A(n38766), .B(n38767), .Z(n38757) );
  ANDN U40558 ( .A(n38768), .B(n29954), .Z(n38767) );
  XOR U40559 ( .A(n38769), .B(\modmult_1/zin[0][130] ), .Z(n29954) );
  IV U40560 ( .A(n38766), .Z(n38769) );
  XNOR U40561 ( .A(n38766), .B(n29953), .Z(n38768) );
  XOR U40562 ( .A(n38770), .B(n38771), .Z(n29953) );
  AND U40563 ( .A(\modmult_1/xin[1023] ), .B(n38772), .Z(n38771) );
  IV U40564 ( .A(n38770), .Z(n38772) );
  XOR U40565 ( .A(n38773), .B(g_input[131]), .Z(n38770) );
  NAND U40566 ( .A(n38774), .B(mul_pow), .Z(n38773) );
  XOR U40567 ( .A(g_input[131]), .B(creg[131]), .Z(n38774) );
  XOR U40568 ( .A(n38775), .B(n38776), .Z(n38766) );
  ANDN U40569 ( .A(n38777), .B(n29960), .Z(n38776) );
  XOR U40570 ( .A(n38778), .B(\modmult_1/zin[0][129] ), .Z(n29960) );
  IV U40571 ( .A(n38775), .Z(n38778) );
  XNOR U40572 ( .A(n38775), .B(n29959), .Z(n38777) );
  XOR U40573 ( .A(n38779), .B(n38780), .Z(n29959) );
  AND U40574 ( .A(\modmult_1/xin[1023] ), .B(n38781), .Z(n38780) );
  IV U40575 ( .A(n38779), .Z(n38781) );
  XOR U40576 ( .A(n38782), .B(g_input[130]), .Z(n38779) );
  NAND U40577 ( .A(n38783), .B(mul_pow), .Z(n38782) );
  XOR U40578 ( .A(g_input[130]), .B(creg[130]), .Z(n38783) );
  XOR U40579 ( .A(n38784), .B(n38785), .Z(n38775) );
  ANDN U40580 ( .A(n38786), .B(n29966), .Z(n38785) );
  XOR U40581 ( .A(n38787), .B(\modmult_1/zin[0][128] ), .Z(n29966) );
  IV U40582 ( .A(n38784), .Z(n38787) );
  XNOR U40583 ( .A(n38784), .B(n29965), .Z(n38786) );
  XOR U40584 ( .A(n38788), .B(n38789), .Z(n29965) );
  AND U40585 ( .A(\modmult_1/xin[1023] ), .B(n38790), .Z(n38789) );
  IV U40586 ( .A(n38788), .Z(n38790) );
  XOR U40587 ( .A(n38791), .B(g_input[129]), .Z(n38788) );
  NAND U40588 ( .A(n38792), .B(mul_pow), .Z(n38791) );
  XOR U40589 ( .A(g_input[129]), .B(creg[129]), .Z(n38792) );
  XOR U40590 ( .A(n38793), .B(n38794), .Z(n38784) );
  ANDN U40591 ( .A(n38795), .B(n29972), .Z(n38794) );
  XOR U40592 ( .A(n38796), .B(\modmult_1/zin[0][127] ), .Z(n29972) );
  IV U40593 ( .A(n38793), .Z(n38796) );
  XNOR U40594 ( .A(n38793), .B(n29971), .Z(n38795) );
  XOR U40595 ( .A(n38797), .B(n38798), .Z(n29971) );
  AND U40596 ( .A(\modmult_1/xin[1023] ), .B(n38799), .Z(n38798) );
  IV U40597 ( .A(n38797), .Z(n38799) );
  XOR U40598 ( .A(n38800), .B(g_input[128]), .Z(n38797) );
  NAND U40599 ( .A(n38801), .B(mul_pow), .Z(n38800) );
  XOR U40600 ( .A(g_input[128]), .B(creg[128]), .Z(n38801) );
  XOR U40601 ( .A(n38802), .B(n38803), .Z(n38793) );
  ANDN U40602 ( .A(n38804), .B(n29978), .Z(n38803) );
  XOR U40603 ( .A(n38805), .B(\modmult_1/zin[0][126] ), .Z(n29978) );
  IV U40604 ( .A(n38802), .Z(n38805) );
  XNOR U40605 ( .A(n38802), .B(n29977), .Z(n38804) );
  XOR U40606 ( .A(n38806), .B(n38807), .Z(n29977) );
  AND U40607 ( .A(\modmult_1/xin[1023] ), .B(n38808), .Z(n38807) );
  IV U40608 ( .A(n38806), .Z(n38808) );
  XOR U40609 ( .A(n38809), .B(g_input[127]), .Z(n38806) );
  NAND U40610 ( .A(n38810), .B(mul_pow), .Z(n38809) );
  XOR U40611 ( .A(g_input[127]), .B(creg[127]), .Z(n38810) );
  XOR U40612 ( .A(n38811), .B(n38812), .Z(n38802) );
  ANDN U40613 ( .A(n38813), .B(n29984), .Z(n38812) );
  XOR U40614 ( .A(n38814), .B(\modmult_1/zin[0][125] ), .Z(n29984) );
  IV U40615 ( .A(n38811), .Z(n38814) );
  XNOR U40616 ( .A(n38811), .B(n29983), .Z(n38813) );
  XOR U40617 ( .A(n38815), .B(n38816), .Z(n29983) );
  AND U40618 ( .A(\modmult_1/xin[1023] ), .B(n38817), .Z(n38816) );
  IV U40619 ( .A(n38815), .Z(n38817) );
  XOR U40620 ( .A(n38818), .B(g_input[126]), .Z(n38815) );
  NAND U40621 ( .A(n38819), .B(mul_pow), .Z(n38818) );
  XOR U40622 ( .A(g_input[126]), .B(creg[126]), .Z(n38819) );
  XOR U40623 ( .A(n38820), .B(n38821), .Z(n38811) );
  ANDN U40624 ( .A(n38822), .B(n29990), .Z(n38821) );
  XOR U40625 ( .A(n38823), .B(\modmult_1/zin[0][124] ), .Z(n29990) );
  IV U40626 ( .A(n38820), .Z(n38823) );
  XNOR U40627 ( .A(n38820), .B(n29989), .Z(n38822) );
  XOR U40628 ( .A(n38824), .B(n38825), .Z(n29989) );
  AND U40629 ( .A(\modmult_1/xin[1023] ), .B(n38826), .Z(n38825) );
  IV U40630 ( .A(n38824), .Z(n38826) );
  XOR U40631 ( .A(n38827), .B(g_input[125]), .Z(n38824) );
  NAND U40632 ( .A(n38828), .B(mul_pow), .Z(n38827) );
  XOR U40633 ( .A(g_input[125]), .B(creg[125]), .Z(n38828) );
  XOR U40634 ( .A(n38829), .B(n38830), .Z(n38820) );
  ANDN U40635 ( .A(n38831), .B(n29996), .Z(n38830) );
  XOR U40636 ( .A(n38832), .B(\modmult_1/zin[0][123] ), .Z(n29996) );
  IV U40637 ( .A(n38829), .Z(n38832) );
  XNOR U40638 ( .A(n38829), .B(n29995), .Z(n38831) );
  XOR U40639 ( .A(n38833), .B(n38834), .Z(n29995) );
  AND U40640 ( .A(\modmult_1/xin[1023] ), .B(n38835), .Z(n38834) );
  IV U40641 ( .A(n38833), .Z(n38835) );
  XOR U40642 ( .A(n38836), .B(g_input[124]), .Z(n38833) );
  NAND U40643 ( .A(n38837), .B(mul_pow), .Z(n38836) );
  XOR U40644 ( .A(g_input[124]), .B(creg[124]), .Z(n38837) );
  XOR U40645 ( .A(n38838), .B(n38839), .Z(n38829) );
  ANDN U40646 ( .A(n38840), .B(n30002), .Z(n38839) );
  XOR U40647 ( .A(n38841), .B(\modmult_1/zin[0][122] ), .Z(n30002) );
  IV U40648 ( .A(n38838), .Z(n38841) );
  XNOR U40649 ( .A(n38838), .B(n30001), .Z(n38840) );
  XOR U40650 ( .A(n38842), .B(n38843), .Z(n30001) );
  AND U40651 ( .A(\modmult_1/xin[1023] ), .B(n38844), .Z(n38843) );
  IV U40652 ( .A(n38842), .Z(n38844) );
  XOR U40653 ( .A(n38845), .B(g_input[123]), .Z(n38842) );
  NAND U40654 ( .A(n38846), .B(mul_pow), .Z(n38845) );
  XOR U40655 ( .A(g_input[123]), .B(creg[123]), .Z(n38846) );
  XOR U40656 ( .A(n38847), .B(n38848), .Z(n38838) );
  ANDN U40657 ( .A(n38849), .B(n30008), .Z(n38848) );
  XOR U40658 ( .A(n38850), .B(\modmult_1/zin[0][121] ), .Z(n30008) );
  IV U40659 ( .A(n38847), .Z(n38850) );
  XNOR U40660 ( .A(n38847), .B(n30007), .Z(n38849) );
  XOR U40661 ( .A(n38851), .B(n38852), .Z(n30007) );
  AND U40662 ( .A(\modmult_1/xin[1023] ), .B(n38853), .Z(n38852) );
  IV U40663 ( .A(n38851), .Z(n38853) );
  XOR U40664 ( .A(n38854), .B(g_input[122]), .Z(n38851) );
  NAND U40665 ( .A(n38855), .B(mul_pow), .Z(n38854) );
  XOR U40666 ( .A(g_input[122]), .B(creg[122]), .Z(n38855) );
  XOR U40667 ( .A(n38856), .B(n38857), .Z(n38847) );
  ANDN U40668 ( .A(n38858), .B(n30014), .Z(n38857) );
  XOR U40669 ( .A(n38859), .B(\modmult_1/zin[0][120] ), .Z(n30014) );
  IV U40670 ( .A(n38856), .Z(n38859) );
  XNOR U40671 ( .A(n38856), .B(n30013), .Z(n38858) );
  XOR U40672 ( .A(n38860), .B(n38861), .Z(n30013) );
  AND U40673 ( .A(\modmult_1/xin[1023] ), .B(n38862), .Z(n38861) );
  IV U40674 ( .A(n38860), .Z(n38862) );
  XOR U40675 ( .A(n38863), .B(g_input[121]), .Z(n38860) );
  NAND U40676 ( .A(n38864), .B(mul_pow), .Z(n38863) );
  XOR U40677 ( .A(g_input[121]), .B(creg[121]), .Z(n38864) );
  XOR U40678 ( .A(n38865), .B(n38866), .Z(n38856) );
  ANDN U40679 ( .A(n38867), .B(n30020), .Z(n38866) );
  XOR U40680 ( .A(n38868), .B(\modmult_1/zin[0][119] ), .Z(n30020) );
  IV U40681 ( .A(n38865), .Z(n38868) );
  XNOR U40682 ( .A(n38865), .B(n30019), .Z(n38867) );
  XOR U40683 ( .A(n38869), .B(n38870), .Z(n30019) );
  AND U40684 ( .A(\modmult_1/xin[1023] ), .B(n38871), .Z(n38870) );
  IV U40685 ( .A(n38869), .Z(n38871) );
  XOR U40686 ( .A(n38872), .B(g_input[120]), .Z(n38869) );
  NAND U40687 ( .A(n38873), .B(mul_pow), .Z(n38872) );
  XOR U40688 ( .A(g_input[120]), .B(creg[120]), .Z(n38873) );
  XOR U40689 ( .A(n38874), .B(n38875), .Z(n38865) );
  ANDN U40690 ( .A(n38876), .B(n30026), .Z(n38875) );
  XOR U40691 ( .A(n38877), .B(\modmult_1/zin[0][118] ), .Z(n30026) );
  IV U40692 ( .A(n38874), .Z(n38877) );
  XNOR U40693 ( .A(n38874), .B(n30025), .Z(n38876) );
  XOR U40694 ( .A(n38878), .B(n38879), .Z(n30025) );
  AND U40695 ( .A(\modmult_1/xin[1023] ), .B(n38880), .Z(n38879) );
  IV U40696 ( .A(n38878), .Z(n38880) );
  XOR U40697 ( .A(n38881), .B(g_input[119]), .Z(n38878) );
  NAND U40698 ( .A(n38882), .B(mul_pow), .Z(n38881) );
  XOR U40699 ( .A(g_input[119]), .B(creg[119]), .Z(n38882) );
  XOR U40700 ( .A(n38883), .B(n38884), .Z(n38874) );
  ANDN U40701 ( .A(n38885), .B(n30032), .Z(n38884) );
  XOR U40702 ( .A(n38886), .B(\modmult_1/zin[0][117] ), .Z(n30032) );
  IV U40703 ( .A(n38883), .Z(n38886) );
  XNOR U40704 ( .A(n38883), .B(n30031), .Z(n38885) );
  XOR U40705 ( .A(n38887), .B(n38888), .Z(n30031) );
  AND U40706 ( .A(\modmult_1/xin[1023] ), .B(n38889), .Z(n38888) );
  IV U40707 ( .A(n38887), .Z(n38889) );
  XOR U40708 ( .A(n38890), .B(g_input[118]), .Z(n38887) );
  NAND U40709 ( .A(n38891), .B(mul_pow), .Z(n38890) );
  XOR U40710 ( .A(g_input[118]), .B(creg[118]), .Z(n38891) );
  XOR U40711 ( .A(n38892), .B(n38893), .Z(n38883) );
  ANDN U40712 ( .A(n38894), .B(n30038), .Z(n38893) );
  XOR U40713 ( .A(n38895), .B(\modmult_1/zin[0][116] ), .Z(n30038) );
  IV U40714 ( .A(n38892), .Z(n38895) );
  XNOR U40715 ( .A(n38892), .B(n30037), .Z(n38894) );
  XOR U40716 ( .A(n38896), .B(n38897), .Z(n30037) );
  AND U40717 ( .A(\modmult_1/xin[1023] ), .B(n38898), .Z(n38897) );
  IV U40718 ( .A(n38896), .Z(n38898) );
  XOR U40719 ( .A(n38899), .B(g_input[117]), .Z(n38896) );
  NAND U40720 ( .A(n38900), .B(mul_pow), .Z(n38899) );
  XOR U40721 ( .A(g_input[117]), .B(creg[117]), .Z(n38900) );
  XOR U40722 ( .A(n38901), .B(n38902), .Z(n38892) );
  ANDN U40723 ( .A(n38903), .B(n30044), .Z(n38902) );
  XOR U40724 ( .A(n38904), .B(\modmult_1/zin[0][115] ), .Z(n30044) );
  IV U40725 ( .A(n38901), .Z(n38904) );
  XNOR U40726 ( .A(n38901), .B(n30043), .Z(n38903) );
  XOR U40727 ( .A(n38905), .B(n38906), .Z(n30043) );
  AND U40728 ( .A(\modmult_1/xin[1023] ), .B(n38907), .Z(n38906) );
  IV U40729 ( .A(n38905), .Z(n38907) );
  XOR U40730 ( .A(n38908), .B(g_input[116]), .Z(n38905) );
  NAND U40731 ( .A(n38909), .B(mul_pow), .Z(n38908) );
  XOR U40732 ( .A(g_input[116]), .B(creg[116]), .Z(n38909) );
  XOR U40733 ( .A(n38910), .B(n38911), .Z(n38901) );
  ANDN U40734 ( .A(n38912), .B(n30050), .Z(n38911) );
  XOR U40735 ( .A(n38913), .B(\modmult_1/zin[0][114] ), .Z(n30050) );
  IV U40736 ( .A(n38910), .Z(n38913) );
  XNOR U40737 ( .A(n38910), .B(n30049), .Z(n38912) );
  XOR U40738 ( .A(n38914), .B(n38915), .Z(n30049) );
  AND U40739 ( .A(\modmult_1/xin[1023] ), .B(n38916), .Z(n38915) );
  IV U40740 ( .A(n38914), .Z(n38916) );
  XOR U40741 ( .A(n38917), .B(g_input[115]), .Z(n38914) );
  NAND U40742 ( .A(n38918), .B(mul_pow), .Z(n38917) );
  XOR U40743 ( .A(g_input[115]), .B(creg[115]), .Z(n38918) );
  XOR U40744 ( .A(n38919), .B(n38920), .Z(n38910) );
  ANDN U40745 ( .A(n38921), .B(n30056), .Z(n38920) );
  XOR U40746 ( .A(n38922), .B(\modmult_1/zin[0][113] ), .Z(n30056) );
  IV U40747 ( .A(n38919), .Z(n38922) );
  XNOR U40748 ( .A(n38919), .B(n30055), .Z(n38921) );
  XOR U40749 ( .A(n38923), .B(n38924), .Z(n30055) );
  AND U40750 ( .A(\modmult_1/xin[1023] ), .B(n38925), .Z(n38924) );
  IV U40751 ( .A(n38923), .Z(n38925) );
  XOR U40752 ( .A(n38926), .B(g_input[114]), .Z(n38923) );
  NAND U40753 ( .A(n38927), .B(mul_pow), .Z(n38926) );
  XOR U40754 ( .A(g_input[114]), .B(creg[114]), .Z(n38927) );
  XOR U40755 ( .A(n38928), .B(n38929), .Z(n38919) );
  ANDN U40756 ( .A(n38930), .B(n30062), .Z(n38929) );
  XOR U40757 ( .A(n38931), .B(\modmult_1/zin[0][112] ), .Z(n30062) );
  IV U40758 ( .A(n38928), .Z(n38931) );
  XNOR U40759 ( .A(n38928), .B(n30061), .Z(n38930) );
  XOR U40760 ( .A(n38932), .B(n38933), .Z(n30061) );
  AND U40761 ( .A(\modmult_1/xin[1023] ), .B(n38934), .Z(n38933) );
  IV U40762 ( .A(n38932), .Z(n38934) );
  XOR U40763 ( .A(n38935), .B(g_input[113]), .Z(n38932) );
  NAND U40764 ( .A(n38936), .B(mul_pow), .Z(n38935) );
  XOR U40765 ( .A(g_input[113]), .B(creg[113]), .Z(n38936) );
  XOR U40766 ( .A(n38937), .B(n38938), .Z(n38928) );
  ANDN U40767 ( .A(n38939), .B(n30068), .Z(n38938) );
  XOR U40768 ( .A(n38940), .B(\modmult_1/zin[0][111] ), .Z(n30068) );
  IV U40769 ( .A(n38937), .Z(n38940) );
  XNOR U40770 ( .A(n38937), .B(n30067), .Z(n38939) );
  XOR U40771 ( .A(n38941), .B(n38942), .Z(n30067) );
  AND U40772 ( .A(\modmult_1/xin[1023] ), .B(n38943), .Z(n38942) );
  IV U40773 ( .A(n38941), .Z(n38943) );
  XOR U40774 ( .A(n38944), .B(g_input[112]), .Z(n38941) );
  NAND U40775 ( .A(n38945), .B(mul_pow), .Z(n38944) );
  XOR U40776 ( .A(g_input[112]), .B(creg[112]), .Z(n38945) );
  XOR U40777 ( .A(n38946), .B(n38947), .Z(n38937) );
  ANDN U40778 ( .A(n38948), .B(n30074), .Z(n38947) );
  XOR U40779 ( .A(n38949), .B(\modmult_1/zin[0][110] ), .Z(n30074) );
  IV U40780 ( .A(n38946), .Z(n38949) );
  XNOR U40781 ( .A(n38946), .B(n30073), .Z(n38948) );
  XOR U40782 ( .A(n38950), .B(n38951), .Z(n30073) );
  AND U40783 ( .A(\modmult_1/xin[1023] ), .B(n38952), .Z(n38951) );
  IV U40784 ( .A(n38950), .Z(n38952) );
  XOR U40785 ( .A(n38953), .B(g_input[111]), .Z(n38950) );
  NAND U40786 ( .A(n38954), .B(mul_pow), .Z(n38953) );
  XOR U40787 ( .A(g_input[111]), .B(creg[111]), .Z(n38954) );
  XOR U40788 ( .A(n38955), .B(n38956), .Z(n38946) );
  ANDN U40789 ( .A(n38957), .B(n30080), .Z(n38956) );
  XOR U40790 ( .A(n38958), .B(\modmult_1/zin[0][109] ), .Z(n30080) );
  IV U40791 ( .A(n38955), .Z(n38958) );
  XNOR U40792 ( .A(n38955), .B(n30079), .Z(n38957) );
  XOR U40793 ( .A(n38959), .B(n38960), .Z(n30079) );
  AND U40794 ( .A(\modmult_1/xin[1023] ), .B(n38961), .Z(n38960) );
  IV U40795 ( .A(n38959), .Z(n38961) );
  XOR U40796 ( .A(n38962), .B(g_input[110]), .Z(n38959) );
  NAND U40797 ( .A(n38963), .B(mul_pow), .Z(n38962) );
  XOR U40798 ( .A(g_input[110]), .B(creg[110]), .Z(n38963) );
  XOR U40799 ( .A(n38964), .B(n38965), .Z(n38955) );
  ANDN U40800 ( .A(n38966), .B(n30086), .Z(n38965) );
  XOR U40801 ( .A(n38967), .B(\modmult_1/zin[0][108] ), .Z(n30086) );
  IV U40802 ( .A(n38964), .Z(n38967) );
  XNOR U40803 ( .A(n38964), .B(n30085), .Z(n38966) );
  XOR U40804 ( .A(n38968), .B(n38969), .Z(n30085) );
  AND U40805 ( .A(\modmult_1/xin[1023] ), .B(n38970), .Z(n38969) );
  IV U40806 ( .A(n38968), .Z(n38970) );
  XOR U40807 ( .A(n38971), .B(g_input[109]), .Z(n38968) );
  NAND U40808 ( .A(n38972), .B(mul_pow), .Z(n38971) );
  XOR U40809 ( .A(g_input[109]), .B(creg[109]), .Z(n38972) );
  XOR U40810 ( .A(n38973), .B(n38974), .Z(n38964) );
  ANDN U40811 ( .A(n38975), .B(n30092), .Z(n38974) );
  XOR U40812 ( .A(n38976), .B(\modmult_1/zin[0][107] ), .Z(n30092) );
  IV U40813 ( .A(n38973), .Z(n38976) );
  XNOR U40814 ( .A(n38973), .B(n30091), .Z(n38975) );
  XOR U40815 ( .A(n38977), .B(n38978), .Z(n30091) );
  AND U40816 ( .A(\modmult_1/xin[1023] ), .B(n38979), .Z(n38978) );
  IV U40817 ( .A(n38977), .Z(n38979) );
  XOR U40818 ( .A(n38980), .B(g_input[108]), .Z(n38977) );
  NAND U40819 ( .A(n38981), .B(mul_pow), .Z(n38980) );
  XOR U40820 ( .A(g_input[108]), .B(creg[108]), .Z(n38981) );
  XOR U40821 ( .A(n38982), .B(n38983), .Z(n38973) );
  ANDN U40822 ( .A(n38984), .B(n30098), .Z(n38983) );
  XOR U40823 ( .A(n38985), .B(\modmult_1/zin[0][106] ), .Z(n30098) );
  IV U40824 ( .A(n38982), .Z(n38985) );
  XNOR U40825 ( .A(n38982), .B(n30097), .Z(n38984) );
  XOR U40826 ( .A(n38986), .B(n38987), .Z(n30097) );
  AND U40827 ( .A(\modmult_1/xin[1023] ), .B(n38988), .Z(n38987) );
  IV U40828 ( .A(n38986), .Z(n38988) );
  XOR U40829 ( .A(n38989), .B(g_input[107]), .Z(n38986) );
  NAND U40830 ( .A(n38990), .B(mul_pow), .Z(n38989) );
  XOR U40831 ( .A(g_input[107]), .B(creg[107]), .Z(n38990) );
  XOR U40832 ( .A(n38991), .B(n38992), .Z(n38982) );
  ANDN U40833 ( .A(n38993), .B(n30104), .Z(n38992) );
  XOR U40834 ( .A(n38994), .B(\modmult_1/zin[0][105] ), .Z(n30104) );
  IV U40835 ( .A(n38991), .Z(n38994) );
  XNOR U40836 ( .A(n38991), .B(n30103), .Z(n38993) );
  XOR U40837 ( .A(n38995), .B(n38996), .Z(n30103) );
  AND U40838 ( .A(\modmult_1/xin[1023] ), .B(n38997), .Z(n38996) );
  IV U40839 ( .A(n38995), .Z(n38997) );
  XOR U40840 ( .A(n38998), .B(g_input[106]), .Z(n38995) );
  NAND U40841 ( .A(n38999), .B(mul_pow), .Z(n38998) );
  XOR U40842 ( .A(g_input[106]), .B(creg[106]), .Z(n38999) );
  XOR U40843 ( .A(n39000), .B(n39001), .Z(n38991) );
  ANDN U40844 ( .A(n39002), .B(n30110), .Z(n39001) );
  XOR U40845 ( .A(n39003), .B(\modmult_1/zin[0][104] ), .Z(n30110) );
  IV U40846 ( .A(n39000), .Z(n39003) );
  XNOR U40847 ( .A(n39000), .B(n30109), .Z(n39002) );
  XOR U40848 ( .A(n39004), .B(n39005), .Z(n30109) );
  AND U40849 ( .A(\modmult_1/xin[1023] ), .B(n39006), .Z(n39005) );
  IV U40850 ( .A(n39004), .Z(n39006) );
  XOR U40851 ( .A(n39007), .B(g_input[105]), .Z(n39004) );
  NAND U40852 ( .A(n39008), .B(mul_pow), .Z(n39007) );
  XOR U40853 ( .A(g_input[105]), .B(creg[105]), .Z(n39008) );
  XOR U40854 ( .A(n39009), .B(n39010), .Z(n39000) );
  ANDN U40855 ( .A(n39011), .B(n30116), .Z(n39010) );
  XOR U40856 ( .A(n39012), .B(\modmult_1/zin[0][103] ), .Z(n30116) );
  IV U40857 ( .A(n39009), .Z(n39012) );
  XNOR U40858 ( .A(n39009), .B(n30115), .Z(n39011) );
  XOR U40859 ( .A(n39013), .B(n39014), .Z(n30115) );
  AND U40860 ( .A(\modmult_1/xin[1023] ), .B(n39015), .Z(n39014) );
  IV U40861 ( .A(n39013), .Z(n39015) );
  XOR U40862 ( .A(n39016), .B(g_input[104]), .Z(n39013) );
  NAND U40863 ( .A(n39017), .B(mul_pow), .Z(n39016) );
  XOR U40864 ( .A(g_input[104]), .B(creg[104]), .Z(n39017) );
  XOR U40865 ( .A(n39018), .B(n39019), .Z(n39009) );
  ANDN U40866 ( .A(n39020), .B(n30122), .Z(n39019) );
  XOR U40867 ( .A(n39021), .B(\modmult_1/zin[0][102] ), .Z(n30122) );
  IV U40868 ( .A(n39018), .Z(n39021) );
  XNOR U40869 ( .A(n39018), .B(n30121), .Z(n39020) );
  XOR U40870 ( .A(n39022), .B(n39023), .Z(n30121) );
  AND U40871 ( .A(\modmult_1/xin[1023] ), .B(n39024), .Z(n39023) );
  IV U40872 ( .A(n39022), .Z(n39024) );
  XOR U40873 ( .A(n39025), .B(g_input[103]), .Z(n39022) );
  NAND U40874 ( .A(n39026), .B(mul_pow), .Z(n39025) );
  XOR U40875 ( .A(g_input[103]), .B(creg[103]), .Z(n39026) );
  XOR U40876 ( .A(n39027), .B(n39028), .Z(n39018) );
  ANDN U40877 ( .A(n39029), .B(n30128), .Z(n39028) );
  XOR U40878 ( .A(n39030), .B(\modmult_1/zin[0][101] ), .Z(n30128) );
  IV U40879 ( .A(n39027), .Z(n39030) );
  XNOR U40880 ( .A(n39027), .B(n30127), .Z(n39029) );
  XOR U40881 ( .A(n39031), .B(n39032), .Z(n30127) );
  AND U40882 ( .A(\modmult_1/xin[1023] ), .B(n39033), .Z(n39032) );
  IV U40883 ( .A(n39031), .Z(n39033) );
  XOR U40884 ( .A(n39034), .B(g_input[102]), .Z(n39031) );
  NAND U40885 ( .A(n39035), .B(mul_pow), .Z(n39034) );
  XOR U40886 ( .A(g_input[102]), .B(creg[102]), .Z(n39035) );
  XOR U40887 ( .A(n39036), .B(n39037), .Z(n39027) );
  ANDN U40888 ( .A(n39038), .B(n30134), .Z(n39037) );
  XOR U40889 ( .A(n39039), .B(\modmult_1/zin[0][100] ), .Z(n30134) );
  IV U40890 ( .A(n39036), .Z(n39039) );
  XNOR U40891 ( .A(n39036), .B(n30133), .Z(n39038) );
  XOR U40892 ( .A(n39040), .B(n39041), .Z(n30133) );
  AND U40893 ( .A(\modmult_1/xin[1023] ), .B(n39042), .Z(n39041) );
  IV U40894 ( .A(n39040), .Z(n39042) );
  XOR U40895 ( .A(n39043), .B(g_input[101]), .Z(n39040) );
  NAND U40896 ( .A(n39044), .B(mul_pow), .Z(n39043) );
  XOR U40897 ( .A(g_input[101]), .B(creg[101]), .Z(n39044) );
  XOR U40898 ( .A(n39045), .B(n39046), .Z(n39036) );
  ANDN U40899 ( .A(n39047), .B(n30140), .Z(n39046) );
  XOR U40900 ( .A(n39048), .B(\modmult_1/zin[0][99] ), .Z(n30140) );
  IV U40901 ( .A(n39045), .Z(n39048) );
  XNOR U40902 ( .A(n39045), .B(n30139), .Z(n39047) );
  XOR U40903 ( .A(n39049), .B(n39050), .Z(n30139) );
  AND U40904 ( .A(\modmult_1/xin[1023] ), .B(n39051), .Z(n39050) );
  IV U40905 ( .A(n39049), .Z(n39051) );
  XOR U40906 ( .A(n39052), .B(g_input[100]), .Z(n39049) );
  NAND U40907 ( .A(n39053), .B(mul_pow), .Z(n39052) );
  XOR U40908 ( .A(g_input[100]), .B(creg[100]), .Z(n39053) );
  XOR U40909 ( .A(n39054), .B(n39055), .Z(n39045) );
  ANDN U40910 ( .A(n39056), .B(n30146), .Z(n39055) );
  XOR U40911 ( .A(n39057), .B(\modmult_1/zin[0][98] ), .Z(n30146) );
  IV U40912 ( .A(n39054), .Z(n39057) );
  XNOR U40913 ( .A(n39054), .B(n30145), .Z(n39056) );
  XOR U40914 ( .A(n39058), .B(n39059), .Z(n30145) );
  AND U40915 ( .A(\modmult_1/xin[1023] ), .B(n39060), .Z(n39059) );
  IV U40916 ( .A(n39058), .Z(n39060) );
  XOR U40917 ( .A(n39061), .B(g_input[99]), .Z(n39058) );
  NAND U40918 ( .A(n39062), .B(mul_pow), .Z(n39061) );
  XOR U40919 ( .A(g_input[99]), .B(creg[99]), .Z(n39062) );
  XOR U40920 ( .A(n39063), .B(n39064), .Z(n39054) );
  ANDN U40921 ( .A(n39065), .B(n30152), .Z(n39064) );
  XOR U40922 ( .A(n39066), .B(\modmult_1/zin[0][97] ), .Z(n30152) );
  IV U40923 ( .A(n39063), .Z(n39066) );
  XNOR U40924 ( .A(n39063), .B(n30151), .Z(n39065) );
  XOR U40925 ( .A(n39067), .B(n39068), .Z(n30151) );
  AND U40926 ( .A(\modmult_1/xin[1023] ), .B(n39069), .Z(n39068) );
  IV U40927 ( .A(n39067), .Z(n39069) );
  XOR U40928 ( .A(n39070), .B(g_input[98]), .Z(n39067) );
  NAND U40929 ( .A(n39071), .B(mul_pow), .Z(n39070) );
  XOR U40930 ( .A(g_input[98]), .B(creg[98]), .Z(n39071) );
  XOR U40931 ( .A(n39072), .B(n39073), .Z(n39063) );
  ANDN U40932 ( .A(n39074), .B(n30158), .Z(n39073) );
  XOR U40933 ( .A(n39075), .B(\modmult_1/zin[0][96] ), .Z(n30158) );
  IV U40934 ( .A(n39072), .Z(n39075) );
  XNOR U40935 ( .A(n39072), .B(n30157), .Z(n39074) );
  XOR U40936 ( .A(n39076), .B(n39077), .Z(n30157) );
  AND U40937 ( .A(\modmult_1/xin[1023] ), .B(n39078), .Z(n39077) );
  IV U40938 ( .A(n39076), .Z(n39078) );
  XOR U40939 ( .A(n39079), .B(g_input[97]), .Z(n39076) );
  NAND U40940 ( .A(n39080), .B(mul_pow), .Z(n39079) );
  XOR U40941 ( .A(g_input[97]), .B(creg[97]), .Z(n39080) );
  XOR U40942 ( .A(n39081), .B(n39082), .Z(n39072) );
  ANDN U40943 ( .A(n39083), .B(n30164), .Z(n39082) );
  XOR U40944 ( .A(n39084), .B(\modmult_1/zin[0][95] ), .Z(n30164) );
  IV U40945 ( .A(n39081), .Z(n39084) );
  XNOR U40946 ( .A(n39081), .B(n30163), .Z(n39083) );
  XOR U40947 ( .A(n39085), .B(n39086), .Z(n30163) );
  AND U40948 ( .A(\modmult_1/xin[1023] ), .B(n39087), .Z(n39086) );
  IV U40949 ( .A(n39085), .Z(n39087) );
  XOR U40950 ( .A(n39088), .B(g_input[96]), .Z(n39085) );
  NAND U40951 ( .A(n39089), .B(mul_pow), .Z(n39088) );
  XOR U40952 ( .A(g_input[96]), .B(creg[96]), .Z(n39089) );
  XOR U40953 ( .A(n39090), .B(n39091), .Z(n39081) );
  ANDN U40954 ( .A(n39092), .B(n30170), .Z(n39091) );
  XOR U40955 ( .A(n39093), .B(\modmult_1/zin[0][94] ), .Z(n30170) );
  IV U40956 ( .A(n39090), .Z(n39093) );
  XNOR U40957 ( .A(n39090), .B(n30169), .Z(n39092) );
  XOR U40958 ( .A(n39094), .B(n39095), .Z(n30169) );
  AND U40959 ( .A(\modmult_1/xin[1023] ), .B(n39096), .Z(n39095) );
  IV U40960 ( .A(n39094), .Z(n39096) );
  XOR U40961 ( .A(n39097), .B(g_input[95]), .Z(n39094) );
  NAND U40962 ( .A(n39098), .B(mul_pow), .Z(n39097) );
  XOR U40963 ( .A(g_input[95]), .B(creg[95]), .Z(n39098) );
  XOR U40964 ( .A(n39099), .B(n39100), .Z(n39090) );
  ANDN U40965 ( .A(n39101), .B(n30176), .Z(n39100) );
  XOR U40966 ( .A(n39102), .B(\modmult_1/zin[0][93] ), .Z(n30176) );
  IV U40967 ( .A(n39099), .Z(n39102) );
  XNOR U40968 ( .A(n39099), .B(n30175), .Z(n39101) );
  XOR U40969 ( .A(n39103), .B(n39104), .Z(n30175) );
  AND U40970 ( .A(\modmult_1/xin[1023] ), .B(n39105), .Z(n39104) );
  IV U40971 ( .A(n39103), .Z(n39105) );
  XOR U40972 ( .A(n39106), .B(g_input[94]), .Z(n39103) );
  NAND U40973 ( .A(n39107), .B(mul_pow), .Z(n39106) );
  XOR U40974 ( .A(g_input[94]), .B(creg[94]), .Z(n39107) );
  XOR U40975 ( .A(n39108), .B(n39109), .Z(n39099) );
  ANDN U40976 ( .A(n39110), .B(n30182), .Z(n39109) );
  XOR U40977 ( .A(n39111), .B(\modmult_1/zin[0][92] ), .Z(n30182) );
  IV U40978 ( .A(n39108), .Z(n39111) );
  XNOR U40979 ( .A(n39108), .B(n30181), .Z(n39110) );
  XOR U40980 ( .A(n39112), .B(n39113), .Z(n30181) );
  AND U40981 ( .A(\modmult_1/xin[1023] ), .B(n39114), .Z(n39113) );
  IV U40982 ( .A(n39112), .Z(n39114) );
  XOR U40983 ( .A(n39115), .B(g_input[93]), .Z(n39112) );
  NAND U40984 ( .A(n39116), .B(mul_pow), .Z(n39115) );
  XOR U40985 ( .A(g_input[93]), .B(creg[93]), .Z(n39116) );
  XOR U40986 ( .A(n39117), .B(n39118), .Z(n39108) );
  ANDN U40987 ( .A(n39119), .B(n30188), .Z(n39118) );
  XOR U40988 ( .A(n39120), .B(\modmult_1/zin[0][91] ), .Z(n30188) );
  IV U40989 ( .A(n39117), .Z(n39120) );
  XNOR U40990 ( .A(n39117), .B(n30187), .Z(n39119) );
  XOR U40991 ( .A(n39121), .B(n39122), .Z(n30187) );
  AND U40992 ( .A(\modmult_1/xin[1023] ), .B(n39123), .Z(n39122) );
  IV U40993 ( .A(n39121), .Z(n39123) );
  XOR U40994 ( .A(n39124), .B(g_input[92]), .Z(n39121) );
  NAND U40995 ( .A(n39125), .B(mul_pow), .Z(n39124) );
  XOR U40996 ( .A(g_input[92]), .B(creg[92]), .Z(n39125) );
  XOR U40997 ( .A(n39126), .B(n39127), .Z(n39117) );
  ANDN U40998 ( .A(n39128), .B(n30194), .Z(n39127) );
  XOR U40999 ( .A(n39129), .B(\modmult_1/zin[0][90] ), .Z(n30194) );
  IV U41000 ( .A(n39126), .Z(n39129) );
  XNOR U41001 ( .A(n39126), .B(n30193), .Z(n39128) );
  XOR U41002 ( .A(n39130), .B(n39131), .Z(n30193) );
  AND U41003 ( .A(\modmult_1/xin[1023] ), .B(n39132), .Z(n39131) );
  IV U41004 ( .A(n39130), .Z(n39132) );
  XOR U41005 ( .A(n39133), .B(g_input[91]), .Z(n39130) );
  NAND U41006 ( .A(n39134), .B(mul_pow), .Z(n39133) );
  XOR U41007 ( .A(g_input[91]), .B(creg[91]), .Z(n39134) );
  XOR U41008 ( .A(n39135), .B(n39136), .Z(n39126) );
  ANDN U41009 ( .A(n39137), .B(n30200), .Z(n39136) );
  XOR U41010 ( .A(n39138), .B(\modmult_1/zin[0][89] ), .Z(n30200) );
  IV U41011 ( .A(n39135), .Z(n39138) );
  XNOR U41012 ( .A(n39135), .B(n30199), .Z(n39137) );
  XOR U41013 ( .A(n39139), .B(n39140), .Z(n30199) );
  AND U41014 ( .A(\modmult_1/xin[1023] ), .B(n39141), .Z(n39140) );
  IV U41015 ( .A(n39139), .Z(n39141) );
  XOR U41016 ( .A(n39142), .B(g_input[90]), .Z(n39139) );
  NAND U41017 ( .A(n39143), .B(mul_pow), .Z(n39142) );
  XOR U41018 ( .A(g_input[90]), .B(creg[90]), .Z(n39143) );
  XOR U41019 ( .A(n39144), .B(n39145), .Z(n39135) );
  ANDN U41020 ( .A(n39146), .B(n30206), .Z(n39145) );
  XOR U41021 ( .A(n39147), .B(\modmult_1/zin[0][88] ), .Z(n30206) );
  IV U41022 ( .A(n39144), .Z(n39147) );
  XNOR U41023 ( .A(n39144), .B(n30205), .Z(n39146) );
  XOR U41024 ( .A(n39148), .B(n39149), .Z(n30205) );
  AND U41025 ( .A(\modmult_1/xin[1023] ), .B(n39150), .Z(n39149) );
  IV U41026 ( .A(n39148), .Z(n39150) );
  XOR U41027 ( .A(n39151), .B(g_input[89]), .Z(n39148) );
  NAND U41028 ( .A(n39152), .B(mul_pow), .Z(n39151) );
  XOR U41029 ( .A(g_input[89]), .B(creg[89]), .Z(n39152) );
  XOR U41030 ( .A(n39153), .B(n39154), .Z(n39144) );
  ANDN U41031 ( .A(n39155), .B(n30212), .Z(n39154) );
  XOR U41032 ( .A(n39156), .B(\modmult_1/zin[0][87] ), .Z(n30212) );
  IV U41033 ( .A(n39153), .Z(n39156) );
  XNOR U41034 ( .A(n39153), .B(n30211), .Z(n39155) );
  XOR U41035 ( .A(n39157), .B(n39158), .Z(n30211) );
  AND U41036 ( .A(\modmult_1/xin[1023] ), .B(n39159), .Z(n39158) );
  IV U41037 ( .A(n39157), .Z(n39159) );
  XOR U41038 ( .A(n39160), .B(g_input[88]), .Z(n39157) );
  NAND U41039 ( .A(n39161), .B(mul_pow), .Z(n39160) );
  XOR U41040 ( .A(g_input[88]), .B(creg[88]), .Z(n39161) );
  XOR U41041 ( .A(n39162), .B(n39163), .Z(n39153) );
  ANDN U41042 ( .A(n39164), .B(n30218), .Z(n39163) );
  XOR U41043 ( .A(n39165), .B(\modmult_1/zin[0][86] ), .Z(n30218) );
  IV U41044 ( .A(n39162), .Z(n39165) );
  XNOR U41045 ( .A(n39162), .B(n30217), .Z(n39164) );
  XOR U41046 ( .A(n39166), .B(n39167), .Z(n30217) );
  AND U41047 ( .A(\modmult_1/xin[1023] ), .B(n39168), .Z(n39167) );
  IV U41048 ( .A(n39166), .Z(n39168) );
  XOR U41049 ( .A(n39169), .B(g_input[87]), .Z(n39166) );
  NAND U41050 ( .A(n39170), .B(mul_pow), .Z(n39169) );
  XOR U41051 ( .A(g_input[87]), .B(creg[87]), .Z(n39170) );
  XOR U41052 ( .A(n39171), .B(n39172), .Z(n39162) );
  ANDN U41053 ( .A(n39173), .B(n30224), .Z(n39172) );
  XOR U41054 ( .A(n39174), .B(\modmult_1/zin[0][85] ), .Z(n30224) );
  IV U41055 ( .A(n39171), .Z(n39174) );
  XNOR U41056 ( .A(n39171), .B(n30223), .Z(n39173) );
  XOR U41057 ( .A(n39175), .B(n39176), .Z(n30223) );
  AND U41058 ( .A(\modmult_1/xin[1023] ), .B(n39177), .Z(n39176) );
  IV U41059 ( .A(n39175), .Z(n39177) );
  XOR U41060 ( .A(n39178), .B(g_input[86]), .Z(n39175) );
  NAND U41061 ( .A(n39179), .B(mul_pow), .Z(n39178) );
  XOR U41062 ( .A(g_input[86]), .B(creg[86]), .Z(n39179) );
  XOR U41063 ( .A(n39180), .B(n39181), .Z(n39171) );
  ANDN U41064 ( .A(n39182), .B(n30230), .Z(n39181) );
  XOR U41065 ( .A(n39183), .B(\modmult_1/zin[0][84] ), .Z(n30230) );
  IV U41066 ( .A(n39180), .Z(n39183) );
  XNOR U41067 ( .A(n39180), .B(n30229), .Z(n39182) );
  XOR U41068 ( .A(n39184), .B(n39185), .Z(n30229) );
  AND U41069 ( .A(\modmult_1/xin[1023] ), .B(n39186), .Z(n39185) );
  IV U41070 ( .A(n39184), .Z(n39186) );
  XOR U41071 ( .A(n39187), .B(g_input[85]), .Z(n39184) );
  NAND U41072 ( .A(n39188), .B(mul_pow), .Z(n39187) );
  XOR U41073 ( .A(g_input[85]), .B(creg[85]), .Z(n39188) );
  XOR U41074 ( .A(n39189), .B(n39190), .Z(n39180) );
  ANDN U41075 ( .A(n39191), .B(n30236), .Z(n39190) );
  XOR U41076 ( .A(n39192), .B(\modmult_1/zin[0][83] ), .Z(n30236) );
  IV U41077 ( .A(n39189), .Z(n39192) );
  XNOR U41078 ( .A(n39189), .B(n30235), .Z(n39191) );
  XOR U41079 ( .A(n39193), .B(n39194), .Z(n30235) );
  AND U41080 ( .A(\modmult_1/xin[1023] ), .B(n39195), .Z(n39194) );
  IV U41081 ( .A(n39193), .Z(n39195) );
  XOR U41082 ( .A(n39196), .B(g_input[84]), .Z(n39193) );
  NAND U41083 ( .A(n39197), .B(mul_pow), .Z(n39196) );
  XOR U41084 ( .A(g_input[84]), .B(creg[84]), .Z(n39197) );
  XOR U41085 ( .A(n39198), .B(n39199), .Z(n39189) );
  ANDN U41086 ( .A(n39200), .B(n30242), .Z(n39199) );
  XOR U41087 ( .A(n39201), .B(\modmult_1/zin[0][82] ), .Z(n30242) );
  IV U41088 ( .A(n39198), .Z(n39201) );
  XNOR U41089 ( .A(n39198), .B(n30241), .Z(n39200) );
  XOR U41090 ( .A(n39202), .B(n39203), .Z(n30241) );
  AND U41091 ( .A(\modmult_1/xin[1023] ), .B(n39204), .Z(n39203) );
  IV U41092 ( .A(n39202), .Z(n39204) );
  XOR U41093 ( .A(n39205), .B(g_input[83]), .Z(n39202) );
  NAND U41094 ( .A(n39206), .B(mul_pow), .Z(n39205) );
  XOR U41095 ( .A(g_input[83]), .B(creg[83]), .Z(n39206) );
  XOR U41096 ( .A(n39207), .B(n39208), .Z(n39198) );
  ANDN U41097 ( .A(n39209), .B(n30248), .Z(n39208) );
  XOR U41098 ( .A(n39210), .B(\modmult_1/zin[0][81] ), .Z(n30248) );
  IV U41099 ( .A(n39207), .Z(n39210) );
  XNOR U41100 ( .A(n39207), .B(n30247), .Z(n39209) );
  XOR U41101 ( .A(n39211), .B(n39212), .Z(n30247) );
  AND U41102 ( .A(\modmult_1/xin[1023] ), .B(n39213), .Z(n39212) );
  IV U41103 ( .A(n39211), .Z(n39213) );
  XOR U41104 ( .A(n39214), .B(g_input[82]), .Z(n39211) );
  NAND U41105 ( .A(n39215), .B(mul_pow), .Z(n39214) );
  XOR U41106 ( .A(g_input[82]), .B(creg[82]), .Z(n39215) );
  XOR U41107 ( .A(n39216), .B(n39217), .Z(n39207) );
  ANDN U41108 ( .A(n39218), .B(n30254), .Z(n39217) );
  XOR U41109 ( .A(n39219), .B(\modmult_1/zin[0][80] ), .Z(n30254) );
  IV U41110 ( .A(n39216), .Z(n39219) );
  XNOR U41111 ( .A(n39216), .B(n30253), .Z(n39218) );
  XOR U41112 ( .A(n39220), .B(n39221), .Z(n30253) );
  AND U41113 ( .A(\modmult_1/xin[1023] ), .B(n39222), .Z(n39221) );
  IV U41114 ( .A(n39220), .Z(n39222) );
  XOR U41115 ( .A(n39223), .B(g_input[81]), .Z(n39220) );
  NAND U41116 ( .A(n39224), .B(mul_pow), .Z(n39223) );
  XOR U41117 ( .A(g_input[81]), .B(creg[81]), .Z(n39224) );
  XOR U41118 ( .A(n39225), .B(n39226), .Z(n39216) );
  ANDN U41119 ( .A(n39227), .B(n30260), .Z(n39226) );
  XOR U41120 ( .A(n39228), .B(\modmult_1/zin[0][79] ), .Z(n30260) );
  IV U41121 ( .A(n39225), .Z(n39228) );
  XNOR U41122 ( .A(n39225), .B(n30259), .Z(n39227) );
  XOR U41123 ( .A(n39229), .B(n39230), .Z(n30259) );
  AND U41124 ( .A(\modmult_1/xin[1023] ), .B(n39231), .Z(n39230) );
  IV U41125 ( .A(n39229), .Z(n39231) );
  XOR U41126 ( .A(n39232), .B(g_input[80]), .Z(n39229) );
  NAND U41127 ( .A(n39233), .B(mul_pow), .Z(n39232) );
  XOR U41128 ( .A(g_input[80]), .B(creg[80]), .Z(n39233) );
  XOR U41129 ( .A(n39234), .B(n39235), .Z(n39225) );
  ANDN U41130 ( .A(n39236), .B(n30266), .Z(n39235) );
  XOR U41131 ( .A(n39237), .B(\modmult_1/zin[0][78] ), .Z(n30266) );
  IV U41132 ( .A(n39234), .Z(n39237) );
  XNOR U41133 ( .A(n39234), .B(n30265), .Z(n39236) );
  XOR U41134 ( .A(n39238), .B(n39239), .Z(n30265) );
  AND U41135 ( .A(\modmult_1/xin[1023] ), .B(n39240), .Z(n39239) );
  IV U41136 ( .A(n39238), .Z(n39240) );
  XOR U41137 ( .A(n39241), .B(g_input[79]), .Z(n39238) );
  NAND U41138 ( .A(n39242), .B(mul_pow), .Z(n39241) );
  XOR U41139 ( .A(g_input[79]), .B(creg[79]), .Z(n39242) );
  XOR U41140 ( .A(n39243), .B(n39244), .Z(n39234) );
  ANDN U41141 ( .A(n39245), .B(n30272), .Z(n39244) );
  XOR U41142 ( .A(n39246), .B(\modmult_1/zin[0][77] ), .Z(n30272) );
  IV U41143 ( .A(n39243), .Z(n39246) );
  XNOR U41144 ( .A(n39243), .B(n30271), .Z(n39245) );
  XOR U41145 ( .A(n39247), .B(n39248), .Z(n30271) );
  AND U41146 ( .A(\modmult_1/xin[1023] ), .B(n39249), .Z(n39248) );
  IV U41147 ( .A(n39247), .Z(n39249) );
  XOR U41148 ( .A(n39250), .B(g_input[78]), .Z(n39247) );
  NAND U41149 ( .A(n39251), .B(mul_pow), .Z(n39250) );
  XOR U41150 ( .A(g_input[78]), .B(creg[78]), .Z(n39251) );
  XOR U41151 ( .A(n39252), .B(n39253), .Z(n39243) );
  ANDN U41152 ( .A(n39254), .B(n30278), .Z(n39253) );
  XOR U41153 ( .A(n39255), .B(\modmult_1/zin[0][76] ), .Z(n30278) );
  IV U41154 ( .A(n39252), .Z(n39255) );
  XNOR U41155 ( .A(n39252), .B(n30277), .Z(n39254) );
  XOR U41156 ( .A(n39256), .B(n39257), .Z(n30277) );
  AND U41157 ( .A(\modmult_1/xin[1023] ), .B(n39258), .Z(n39257) );
  IV U41158 ( .A(n39256), .Z(n39258) );
  XOR U41159 ( .A(n39259), .B(g_input[77]), .Z(n39256) );
  NAND U41160 ( .A(n39260), .B(mul_pow), .Z(n39259) );
  XOR U41161 ( .A(g_input[77]), .B(creg[77]), .Z(n39260) );
  XOR U41162 ( .A(n39261), .B(n39262), .Z(n39252) );
  ANDN U41163 ( .A(n39263), .B(n30284), .Z(n39262) );
  XOR U41164 ( .A(n39264), .B(\modmult_1/zin[0][75] ), .Z(n30284) );
  IV U41165 ( .A(n39261), .Z(n39264) );
  XNOR U41166 ( .A(n39261), .B(n30283), .Z(n39263) );
  XOR U41167 ( .A(n39265), .B(n39266), .Z(n30283) );
  AND U41168 ( .A(\modmult_1/xin[1023] ), .B(n39267), .Z(n39266) );
  IV U41169 ( .A(n39265), .Z(n39267) );
  XOR U41170 ( .A(n39268), .B(g_input[76]), .Z(n39265) );
  NAND U41171 ( .A(n39269), .B(mul_pow), .Z(n39268) );
  XOR U41172 ( .A(g_input[76]), .B(creg[76]), .Z(n39269) );
  XOR U41173 ( .A(n39270), .B(n39271), .Z(n39261) );
  ANDN U41174 ( .A(n39272), .B(n30290), .Z(n39271) );
  XOR U41175 ( .A(n39273), .B(\modmult_1/zin[0][74] ), .Z(n30290) );
  IV U41176 ( .A(n39270), .Z(n39273) );
  XNOR U41177 ( .A(n39270), .B(n30289), .Z(n39272) );
  XOR U41178 ( .A(n39274), .B(n39275), .Z(n30289) );
  AND U41179 ( .A(\modmult_1/xin[1023] ), .B(n39276), .Z(n39275) );
  IV U41180 ( .A(n39274), .Z(n39276) );
  XOR U41181 ( .A(n39277), .B(g_input[75]), .Z(n39274) );
  NAND U41182 ( .A(n39278), .B(mul_pow), .Z(n39277) );
  XOR U41183 ( .A(g_input[75]), .B(creg[75]), .Z(n39278) );
  XOR U41184 ( .A(n39279), .B(n39280), .Z(n39270) );
  ANDN U41185 ( .A(n39281), .B(n30296), .Z(n39280) );
  XOR U41186 ( .A(n39282), .B(\modmult_1/zin[0][73] ), .Z(n30296) );
  IV U41187 ( .A(n39279), .Z(n39282) );
  XNOR U41188 ( .A(n39279), .B(n30295), .Z(n39281) );
  XOR U41189 ( .A(n39283), .B(n39284), .Z(n30295) );
  AND U41190 ( .A(\modmult_1/xin[1023] ), .B(n39285), .Z(n39284) );
  IV U41191 ( .A(n39283), .Z(n39285) );
  XOR U41192 ( .A(n39286), .B(g_input[74]), .Z(n39283) );
  NAND U41193 ( .A(n39287), .B(mul_pow), .Z(n39286) );
  XOR U41194 ( .A(g_input[74]), .B(creg[74]), .Z(n39287) );
  XOR U41195 ( .A(n39288), .B(n39289), .Z(n39279) );
  ANDN U41196 ( .A(n39290), .B(n30302), .Z(n39289) );
  XOR U41197 ( .A(n39291), .B(\modmult_1/zin[0][72] ), .Z(n30302) );
  IV U41198 ( .A(n39288), .Z(n39291) );
  XNOR U41199 ( .A(n39288), .B(n30301), .Z(n39290) );
  XOR U41200 ( .A(n39292), .B(n39293), .Z(n30301) );
  AND U41201 ( .A(\modmult_1/xin[1023] ), .B(n39294), .Z(n39293) );
  IV U41202 ( .A(n39292), .Z(n39294) );
  XOR U41203 ( .A(n39295), .B(g_input[73]), .Z(n39292) );
  NAND U41204 ( .A(n39296), .B(mul_pow), .Z(n39295) );
  XOR U41205 ( .A(g_input[73]), .B(creg[73]), .Z(n39296) );
  XOR U41206 ( .A(n39297), .B(n39298), .Z(n39288) );
  ANDN U41207 ( .A(n39299), .B(n30308), .Z(n39298) );
  XOR U41208 ( .A(n39300), .B(\modmult_1/zin[0][71] ), .Z(n30308) );
  IV U41209 ( .A(n39297), .Z(n39300) );
  XNOR U41210 ( .A(n39297), .B(n30307), .Z(n39299) );
  XOR U41211 ( .A(n39301), .B(n39302), .Z(n30307) );
  AND U41212 ( .A(\modmult_1/xin[1023] ), .B(n39303), .Z(n39302) );
  IV U41213 ( .A(n39301), .Z(n39303) );
  XOR U41214 ( .A(n39304), .B(g_input[72]), .Z(n39301) );
  NAND U41215 ( .A(n39305), .B(mul_pow), .Z(n39304) );
  XOR U41216 ( .A(g_input[72]), .B(creg[72]), .Z(n39305) );
  XOR U41217 ( .A(n39306), .B(n39307), .Z(n39297) );
  ANDN U41218 ( .A(n39308), .B(n30314), .Z(n39307) );
  XOR U41219 ( .A(n39309), .B(\modmult_1/zin[0][70] ), .Z(n30314) );
  IV U41220 ( .A(n39306), .Z(n39309) );
  XNOR U41221 ( .A(n39306), .B(n30313), .Z(n39308) );
  XOR U41222 ( .A(n39310), .B(n39311), .Z(n30313) );
  AND U41223 ( .A(\modmult_1/xin[1023] ), .B(n39312), .Z(n39311) );
  IV U41224 ( .A(n39310), .Z(n39312) );
  XOR U41225 ( .A(n39313), .B(g_input[71]), .Z(n39310) );
  NAND U41226 ( .A(n39314), .B(mul_pow), .Z(n39313) );
  XOR U41227 ( .A(g_input[71]), .B(creg[71]), .Z(n39314) );
  XOR U41228 ( .A(n39315), .B(n39316), .Z(n39306) );
  ANDN U41229 ( .A(n39317), .B(n30320), .Z(n39316) );
  XOR U41230 ( .A(n39318), .B(\modmult_1/zin[0][69] ), .Z(n30320) );
  IV U41231 ( .A(n39315), .Z(n39318) );
  XNOR U41232 ( .A(n39315), .B(n30319), .Z(n39317) );
  XOR U41233 ( .A(n39319), .B(n39320), .Z(n30319) );
  AND U41234 ( .A(\modmult_1/xin[1023] ), .B(n39321), .Z(n39320) );
  IV U41235 ( .A(n39319), .Z(n39321) );
  XOR U41236 ( .A(n39322), .B(g_input[70]), .Z(n39319) );
  NAND U41237 ( .A(n39323), .B(mul_pow), .Z(n39322) );
  XOR U41238 ( .A(g_input[70]), .B(creg[70]), .Z(n39323) );
  XOR U41239 ( .A(n39324), .B(n39325), .Z(n39315) );
  ANDN U41240 ( .A(n39326), .B(n30326), .Z(n39325) );
  XOR U41241 ( .A(n39327), .B(\modmult_1/zin[0][68] ), .Z(n30326) );
  IV U41242 ( .A(n39324), .Z(n39327) );
  XNOR U41243 ( .A(n39324), .B(n30325), .Z(n39326) );
  XOR U41244 ( .A(n39328), .B(n39329), .Z(n30325) );
  AND U41245 ( .A(\modmult_1/xin[1023] ), .B(n39330), .Z(n39329) );
  IV U41246 ( .A(n39328), .Z(n39330) );
  XOR U41247 ( .A(n39331), .B(g_input[69]), .Z(n39328) );
  NAND U41248 ( .A(n39332), .B(mul_pow), .Z(n39331) );
  XOR U41249 ( .A(g_input[69]), .B(creg[69]), .Z(n39332) );
  XOR U41250 ( .A(n39333), .B(n39334), .Z(n39324) );
  ANDN U41251 ( .A(n39335), .B(n30332), .Z(n39334) );
  XOR U41252 ( .A(n39336), .B(\modmult_1/zin[0][67] ), .Z(n30332) );
  IV U41253 ( .A(n39333), .Z(n39336) );
  XNOR U41254 ( .A(n39333), .B(n30331), .Z(n39335) );
  XOR U41255 ( .A(n39337), .B(n39338), .Z(n30331) );
  AND U41256 ( .A(\modmult_1/xin[1023] ), .B(n39339), .Z(n39338) );
  IV U41257 ( .A(n39337), .Z(n39339) );
  XOR U41258 ( .A(n39340), .B(g_input[68]), .Z(n39337) );
  NAND U41259 ( .A(n39341), .B(mul_pow), .Z(n39340) );
  XOR U41260 ( .A(g_input[68]), .B(creg[68]), .Z(n39341) );
  XOR U41261 ( .A(n39342), .B(n39343), .Z(n39333) );
  ANDN U41262 ( .A(n39344), .B(n30338), .Z(n39343) );
  XOR U41263 ( .A(n39345), .B(\modmult_1/zin[0][66] ), .Z(n30338) );
  IV U41264 ( .A(n39342), .Z(n39345) );
  XNOR U41265 ( .A(n39342), .B(n30337), .Z(n39344) );
  XOR U41266 ( .A(n39346), .B(n39347), .Z(n30337) );
  AND U41267 ( .A(\modmult_1/xin[1023] ), .B(n39348), .Z(n39347) );
  IV U41268 ( .A(n39346), .Z(n39348) );
  XOR U41269 ( .A(n39349), .B(g_input[67]), .Z(n39346) );
  NAND U41270 ( .A(n39350), .B(mul_pow), .Z(n39349) );
  XOR U41271 ( .A(g_input[67]), .B(creg[67]), .Z(n39350) );
  XOR U41272 ( .A(n39351), .B(n39352), .Z(n39342) );
  ANDN U41273 ( .A(n39353), .B(n30344), .Z(n39352) );
  XOR U41274 ( .A(n39354), .B(\modmult_1/zin[0][65] ), .Z(n30344) );
  IV U41275 ( .A(n39351), .Z(n39354) );
  XNOR U41276 ( .A(n39351), .B(n30343), .Z(n39353) );
  XOR U41277 ( .A(n39355), .B(n39356), .Z(n30343) );
  AND U41278 ( .A(\modmult_1/xin[1023] ), .B(n39357), .Z(n39356) );
  IV U41279 ( .A(n39355), .Z(n39357) );
  XOR U41280 ( .A(n39358), .B(g_input[66]), .Z(n39355) );
  NAND U41281 ( .A(n39359), .B(mul_pow), .Z(n39358) );
  XOR U41282 ( .A(g_input[66]), .B(creg[66]), .Z(n39359) );
  XOR U41283 ( .A(n39360), .B(n39361), .Z(n39351) );
  ANDN U41284 ( .A(n39362), .B(n30350), .Z(n39361) );
  XOR U41285 ( .A(n39363), .B(\modmult_1/zin[0][64] ), .Z(n30350) );
  IV U41286 ( .A(n39360), .Z(n39363) );
  XNOR U41287 ( .A(n39360), .B(n30349), .Z(n39362) );
  XOR U41288 ( .A(n39364), .B(n39365), .Z(n30349) );
  AND U41289 ( .A(\modmult_1/xin[1023] ), .B(n39366), .Z(n39365) );
  IV U41290 ( .A(n39364), .Z(n39366) );
  XOR U41291 ( .A(n39367), .B(g_input[65]), .Z(n39364) );
  NAND U41292 ( .A(n39368), .B(mul_pow), .Z(n39367) );
  XOR U41293 ( .A(g_input[65]), .B(creg[65]), .Z(n39368) );
  XOR U41294 ( .A(n39369), .B(n39370), .Z(n39360) );
  ANDN U41295 ( .A(n39371), .B(n30356), .Z(n39370) );
  XOR U41296 ( .A(n39372), .B(\modmult_1/zin[0][63] ), .Z(n30356) );
  IV U41297 ( .A(n39369), .Z(n39372) );
  XNOR U41298 ( .A(n39369), .B(n30355), .Z(n39371) );
  XOR U41299 ( .A(n39373), .B(n39374), .Z(n30355) );
  AND U41300 ( .A(\modmult_1/xin[1023] ), .B(n39375), .Z(n39374) );
  IV U41301 ( .A(n39373), .Z(n39375) );
  XOR U41302 ( .A(n39376), .B(g_input[64]), .Z(n39373) );
  NAND U41303 ( .A(n39377), .B(mul_pow), .Z(n39376) );
  XOR U41304 ( .A(g_input[64]), .B(creg[64]), .Z(n39377) );
  XOR U41305 ( .A(n39378), .B(n39379), .Z(n39369) );
  ANDN U41306 ( .A(n39380), .B(n30362), .Z(n39379) );
  XOR U41307 ( .A(n39381), .B(\modmult_1/zin[0][62] ), .Z(n30362) );
  IV U41308 ( .A(n39378), .Z(n39381) );
  XNOR U41309 ( .A(n39378), .B(n30361), .Z(n39380) );
  XOR U41310 ( .A(n39382), .B(n39383), .Z(n30361) );
  AND U41311 ( .A(\modmult_1/xin[1023] ), .B(n39384), .Z(n39383) );
  IV U41312 ( .A(n39382), .Z(n39384) );
  XOR U41313 ( .A(n39385), .B(g_input[63]), .Z(n39382) );
  NAND U41314 ( .A(n39386), .B(mul_pow), .Z(n39385) );
  XOR U41315 ( .A(g_input[63]), .B(creg[63]), .Z(n39386) );
  XOR U41316 ( .A(n39387), .B(n39388), .Z(n39378) );
  ANDN U41317 ( .A(n39389), .B(n30368), .Z(n39388) );
  XOR U41318 ( .A(n39390), .B(\modmult_1/zin[0][61] ), .Z(n30368) );
  IV U41319 ( .A(n39387), .Z(n39390) );
  XNOR U41320 ( .A(n39387), .B(n30367), .Z(n39389) );
  XOR U41321 ( .A(n39391), .B(n39392), .Z(n30367) );
  AND U41322 ( .A(\modmult_1/xin[1023] ), .B(n39393), .Z(n39392) );
  IV U41323 ( .A(n39391), .Z(n39393) );
  XOR U41324 ( .A(n39394), .B(g_input[62]), .Z(n39391) );
  NAND U41325 ( .A(n39395), .B(mul_pow), .Z(n39394) );
  XOR U41326 ( .A(g_input[62]), .B(creg[62]), .Z(n39395) );
  XOR U41327 ( .A(n39396), .B(n39397), .Z(n39387) );
  ANDN U41328 ( .A(n39398), .B(n30374), .Z(n39397) );
  XOR U41329 ( .A(n39399), .B(\modmult_1/zin[0][60] ), .Z(n30374) );
  IV U41330 ( .A(n39396), .Z(n39399) );
  XNOR U41331 ( .A(n39396), .B(n30373), .Z(n39398) );
  XOR U41332 ( .A(n39400), .B(n39401), .Z(n30373) );
  AND U41333 ( .A(\modmult_1/xin[1023] ), .B(n39402), .Z(n39401) );
  IV U41334 ( .A(n39400), .Z(n39402) );
  XOR U41335 ( .A(n39403), .B(g_input[61]), .Z(n39400) );
  NAND U41336 ( .A(n39404), .B(mul_pow), .Z(n39403) );
  XOR U41337 ( .A(g_input[61]), .B(creg[61]), .Z(n39404) );
  XOR U41338 ( .A(n39405), .B(n39406), .Z(n39396) );
  ANDN U41339 ( .A(n39407), .B(n30380), .Z(n39406) );
  XOR U41340 ( .A(n39408), .B(\modmult_1/zin[0][59] ), .Z(n30380) );
  IV U41341 ( .A(n39405), .Z(n39408) );
  XNOR U41342 ( .A(n39405), .B(n30379), .Z(n39407) );
  XOR U41343 ( .A(n39409), .B(n39410), .Z(n30379) );
  AND U41344 ( .A(\modmult_1/xin[1023] ), .B(n39411), .Z(n39410) );
  IV U41345 ( .A(n39409), .Z(n39411) );
  XOR U41346 ( .A(n39412), .B(g_input[60]), .Z(n39409) );
  NAND U41347 ( .A(n39413), .B(mul_pow), .Z(n39412) );
  XOR U41348 ( .A(g_input[60]), .B(creg[60]), .Z(n39413) );
  XOR U41349 ( .A(n39414), .B(n39415), .Z(n39405) );
  ANDN U41350 ( .A(n39416), .B(n30386), .Z(n39415) );
  XOR U41351 ( .A(n39417), .B(\modmult_1/zin[0][58] ), .Z(n30386) );
  IV U41352 ( .A(n39414), .Z(n39417) );
  XNOR U41353 ( .A(n39414), .B(n30385), .Z(n39416) );
  XOR U41354 ( .A(n39418), .B(n39419), .Z(n30385) );
  AND U41355 ( .A(\modmult_1/xin[1023] ), .B(n39420), .Z(n39419) );
  IV U41356 ( .A(n39418), .Z(n39420) );
  XOR U41357 ( .A(n39421), .B(g_input[59]), .Z(n39418) );
  NAND U41358 ( .A(n39422), .B(mul_pow), .Z(n39421) );
  XOR U41359 ( .A(g_input[59]), .B(creg[59]), .Z(n39422) );
  XOR U41360 ( .A(n39423), .B(n39424), .Z(n39414) );
  ANDN U41361 ( .A(n39425), .B(n30392), .Z(n39424) );
  XOR U41362 ( .A(n39426), .B(\modmult_1/zin[0][57] ), .Z(n30392) );
  IV U41363 ( .A(n39423), .Z(n39426) );
  XNOR U41364 ( .A(n39423), .B(n30391), .Z(n39425) );
  XOR U41365 ( .A(n39427), .B(n39428), .Z(n30391) );
  AND U41366 ( .A(\modmult_1/xin[1023] ), .B(n39429), .Z(n39428) );
  IV U41367 ( .A(n39427), .Z(n39429) );
  XOR U41368 ( .A(n39430), .B(g_input[58]), .Z(n39427) );
  NAND U41369 ( .A(n39431), .B(mul_pow), .Z(n39430) );
  XOR U41370 ( .A(g_input[58]), .B(creg[58]), .Z(n39431) );
  XOR U41371 ( .A(n39432), .B(n39433), .Z(n39423) );
  ANDN U41372 ( .A(n39434), .B(n30398), .Z(n39433) );
  XOR U41373 ( .A(n39435), .B(\modmult_1/zin[0][56] ), .Z(n30398) );
  IV U41374 ( .A(n39432), .Z(n39435) );
  XNOR U41375 ( .A(n39432), .B(n30397), .Z(n39434) );
  XOR U41376 ( .A(n39436), .B(n39437), .Z(n30397) );
  AND U41377 ( .A(\modmult_1/xin[1023] ), .B(n39438), .Z(n39437) );
  IV U41378 ( .A(n39436), .Z(n39438) );
  XOR U41379 ( .A(n39439), .B(g_input[57]), .Z(n39436) );
  NAND U41380 ( .A(n39440), .B(mul_pow), .Z(n39439) );
  XOR U41381 ( .A(g_input[57]), .B(creg[57]), .Z(n39440) );
  XOR U41382 ( .A(n39441), .B(n39442), .Z(n39432) );
  ANDN U41383 ( .A(n39443), .B(n30404), .Z(n39442) );
  XOR U41384 ( .A(n39444), .B(\modmult_1/zin[0][55] ), .Z(n30404) );
  IV U41385 ( .A(n39441), .Z(n39444) );
  XNOR U41386 ( .A(n39441), .B(n30403), .Z(n39443) );
  XOR U41387 ( .A(n39445), .B(n39446), .Z(n30403) );
  AND U41388 ( .A(\modmult_1/xin[1023] ), .B(n39447), .Z(n39446) );
  IV U41389 ( .A(n39445), .Z(n39447) );
  XOR U41390 ( .A(n39448), .B(g_input[56]), .Z(n39445) );
  NAND U41391 ( .A(n39449), .B(mul_pow), .Z(n39448) );
  XOR U41392 ( .A(g_input[56]), .B(creg[56]), .Z(n39449) );
  XOR U41393 ( .A(n39450), .B(n39451), .Z(n39441) );
  ANDN U41394 ( .A(n39452), .B(n30410), .Z(n39451) );
  XOR U41395 ( .A(n39453), .B(\modmult_1/zin[0][54] ), .Z(n30410) );
  IV U41396 ( .A(n39450), .Z(n39453) );
  XNOR U41397 ( .A(n39450), .B(n30409), .Z(n39452) );
  XOR U41398 ( .A(n39454), .B(n39455), .Z(n30409) );
  AND U41399 ( .A(\modmult_1/xin[1023] ), .B(n39456), .Z(n39455) );
  IV U41400 ( .A(n39454), .Z(n39456) );
  XOR U41401 ( .A(n39457), .B(g_input[55]), .Z(n39454) );
  NAND U41402 ( .A(n39458), .B(mul_pow), .Z(n39457) );
  XOR U41403 ( .A(g_input[55]), .B(creg[55]), .Z(n39458) );
  XOR U41404 ( .A(n39459), .B(n39460), .Z(n39450) );
  ANDN U41405 ( .A(n39461), .B(n30416), .Z(n39460) );
  XOR U41406 ( .A(n39462), .B(\modmult_1/zin[0][53] ), .Z(n30416) );
  IV U41407 ( .A(n39459), .Z(n39462) );
  XNOR U41408 ( .A(n39459), .B(n30415), .Z(n39461) );
  XOR U41409 ( .A(n39463), .B(n39464), .Z(n30415) );
  AND U41410 ( .A(\modmult_1/xin[1023] ), .B(n39465), .Z(n39464) );
  IV U41411 ( .A(n39463), .Z(n39465) );
  XOR U41412 ( .A(n39466), .B(g_input[54]), .Z(n39463) );
  NAND U41413 ( .A(n39467), .B(mul_pow), .Z(n39466) );
  XOR U41414 ( .A(g_input[54]), .B(creg[54]), .Z(n39467) );
  XOR U41415 ( .A(n39468), .B(n39469), .Z(n39459) );
  ANDN U41416 ( .A(n39470), .B(n30422), .Z(n39469) );
  XOR U41417 ( .A(n39471), .B(\modmult_1/zin[0][52] ), .Z(n30422) );
  IV U41418 ( .A(n39468), .Z(n39471) );
  XNOR U41419 ( .A(n39468), .B(n30421), .Z(n39470) );
  XOR U41420 ( .A(n39472), .B(n39473), .Z(n30421) );
  AND U41421 ( .A(\modmult_1/xin[1023] ), .B(n39474), .Z(n39473) );
  IV U41422 ( .A(n39472), .Z(n39474) );
  XOR U41423 ( .A(n39475), .B(g_input[53]), .Z(n39472) );
  NAND U41424 ( .A(n39476), .B(mul_pow), .Z(n39475) );
  XOR U41425 ( .A(g_input[53]), .B(creg[53]), .Z(n39476) );
  XOR U41426 ( .A(n39477), .B(n39478), .Z(n39468) );
  ANDN U41427 ( .A(n39479), .B(n30428), .Z(n39478) );
  XOR U41428 ( .A(n39480), .B(\modmult_1/zin[0][51] ), .Z(n30428) );
  IV U41429 ( .A(n39477), .Z(n39480) );
  XNOR U41430 ( .A(n39477), .B(n30427), .Z(n39479) );
  XOR U41431 ( .A(n39481), .B(n39482), .Z(n30427) );
  AND U41432 ( .A(\modmult_1/xin[1023] ), .B(n39483), .Z(n39482) );
  IV U41433 ( .A(n39481), .Z(n39483) );
  XOR U41434 ( .A(n39484), .B(g_input[52]), .Z(n39481) );
  NAND U41435 ( .A(n39485), .B(mul_pow), .Z(n39484) );
  XOR U41436 ( .A(g_input[52]), .B(creg[52]), .Z(n39485) );
  XOR U41437 ( .A(n39486), .B(n39487), .Z(n39477) );
  ANDN U41438 ( .A(n39488), .B(n30434), .Z(n39487) );
  XOR U41439 ( .A(n39489), .B(\modmult_1/zin[0][50] ), .Z(n30434) );
  IV U41440 ( .A(n39486), .Z(n39489) );
  XNOR U41441 ( .A(n39486), .B(n30433), .Z(n39488) );
  XOR U41442 ( .A(n39490), .B(n39491), .Z(n30433) );
  AND U41443 ( .A(\modmult_1/xin[1023] ), .B(n39492), .Z(n39491) );
  IV U41444 ( .A(n39490), .Z(n39492) );
  XOR U41445 ( .A(n39493), .B(g_input[51]), .Z(n39490) );
  NAND U41446 ( .A(n39494), .B(mul_pow), .Z(n39493) );
  XOR U41447 ( .A(g_input[51]), .B(creg[51]), .Z(n39494) );
  XOR U41448 ( .A(n39495), .B(n39496), .Z(n39486) );
  ANDN U41449 ( .A(n39497), .B(n30440), .Z(n39496) );
  XOR U41450 ( .A(n39498), .B(\modmult_1/zin[0][49] ), .Z(n30440) );
  IV U41451 ( .A(n39495), .Z(n39498) );
  XNOR U41452 ( .A(n39495), .B(n30439), .Z(n39497) );
  XOR U41453 ( .A(n39499), .B(n39500), .Z(n30439) );
  AND U41454 ( .A(\modmult_1/xin[1023] ), .B(n39501), .Z(n39500) );
  IV U41455 ( .A(n39499), .Z(n39501) );
  XOR U41456 ( .A(n39502), .B(g_input[50]), .Z(n39499) );
  NAND U41457 ( .A(n39503), .B(mul_pow), .Z(n39502) );
  XOR U41458 ( .A(g_input[50]), .B(creg[50]), .Z(n39503) );
  XOR U41459 ( .A(n39504), .B(n39505), .Z(n39495) );
  ANDN U41460 ( .A(n39506), .B(n30446), .Z(n39505) );
  XOR U41461 ( .A(n39507), .B(\modmult_1/zin[0][48] ), .Z(n30446) );
  IV U41462 ( .A(n39504), .Z(n39507) );
  XNOR U41463 ( .A(n39504), .B(n30445), .Z(n39506) );
  XOR U41464 ( .A(n39508), .B(n39509), .Z(n30445) );
  AND U41465 ( .A(\modmult_1/xin[1023] ), .B(n39510), .Z(n39509) );
  IV U41466 ( .A(n39508), .Z(n39510) );
  XOR U41467 ( .A(n39511), .B(g_input[49]), .Z(n39508) );
  NAND U41468 ( .A(n39512), .B(mul_pow), .Z(n39511) );
  XOR U41469 ( .A(g_input[49]), .B(creg[49]), .Z(n39512) );
  XOR U41470 ( .A(n39513), .B(n39514), .Z(n39504) );
  ANDN U41471 ( .A(n39515), .B(n30452), .Z(n39514) );
  XOR U41472 ( .A(n39516), .B(\modmult_1/zin[0][47] ), .Z(n30452) );
  IV U41473 ( .A(n39513), .Z(n39516) );
  XNOR U41474 ( .A(n39513), .B(n30451), .Z(n39515) );
  XOR U41475 ( .A(n39517), .B(n39518), .Z(n30451) );
  AND U41476 ( .A(\modmult_1/xin[1023] ), .B(n39519), .Z(n39518) );
  IV U41477 ( .A(n39517), .Z(n39519) );
  XOR U41478 ( .A(n39520), .B(g_input[48]), .Z(n39517) );
  NAND U41479 ( .A(n39521), .B(mul_pow), .Z(n39520) );
  XOR U41480 ( .A(g_input[48]), .B(creg[48]), .Z(n39521) );
  XOR U41481 ( .A(n39522), .B(n39523), .Z(n39513) );
  ANDN U41482 ( .A(n39524), .B(n30458), .Z(n39523) );
  XOR U41483 ( .A(n39525), .B(\modmult_1/zin[0][46] ), .Z(n30458) );
  IV U41484 ( .A(n39522), .Z(n39525) );
  XNOR U41485 ( .A(n39522), .B(n30457), .Z(n39524) );
  XOR U41486 ( .A(n39526), .B(n39527), .Z(n30457) );
  AND U41487 ( .A(\modmult_1/xin[1023] ), .B(n39528), .Z(n39527) );
  IV U41488 ( .A(n39526), .Z(n39528) );
  XOR U41489 ( .A(n39529), .B(g_input[47]), .Z(n39526) );
  NAND U41490 ( .A(n39530), .B(mul_pow), .Z(n39529) );
  XOR U41491 ( .A(g_input[47]), .B(creg[47]), .Z(n39530) );
  XOR U41492 ( .A(n39531), .B(n39532), .Z(n39522) );
  ANDN U41493 ( .A(n39533), .B(n30464), .Z(n39532) );
  XOR U41494 ( .A(n39534), .B(\modmult_1/zin[0][45] ), .Z(n30464) );
  IV U41495 ( .A(n39531), .Z(n39534) );
  XNOR U41496 ( .A(n39531), .B(n30463), .Z(n39533) );
  XOR U41497 ( .A(n39535), .B(n39536), .Z(n30463) );
  AND U41498 ( .A(\modmult_1/xin[1023] ), .B(n39537), .Z(n39536) );
  IV U41499 ( .A(n39535), .Z(n39537) );
  XOR U41500 ( .A(n39538), .B(g_input[46]), .Z(n39535) );
  NAND U41501 ( .A(n39539), .B(mul_pow), .Z(n39538) );
  XOR U41502 ( .A(g_input[46]), .B(creg[46]), .Z(n39539) );
  XOR U41503 ( .A(n39540), .B(n39541), .Z(n39531) );
  ANDN U41504 ( .A(n39542), .B(n30470), .Z(n39541) );
  XOR U41505 ( .A(n39543), .B(\modmult_1/zin[0][44] ), .Z(n30470) );
  IV U41506 ( .A(n39540), .Z(n39543) );
  XNOR U41507 ( .A(n39540), .B(n30469), .Z(n39542) );
  XOR U41508 ( .A(n39544), .B(n39545), .Z(n30469) );
  AND U41509 ( .A(\modmult_1/xin[1023] ), .B(n39546), .Z(n39545) );
  IV U41510 ( .A(n39544), .Z(n39546) );
  XOR U41511 ( .A(n39547), .B(g_input[45]), .Z(n39544) );
  NAND U41512 ( .A(n39548), .B(mul_pow), .Z(n39547) );
  XOR U41513 ( .A(g_input[45]), .B(creg[45]), .Z(n39548) );
  XOR U41514 ( .A(n39549), .B(n39550), .Z(n39540) );
  ANDN U41515 ( .A(n39551), .B(n30476), .Z(n39550) );
  XOR U41516 ( .A(n39552), .B(\modmult_1/zin[0][43] ), .Z(n30476) );
  IV U41517 ( .A(n39549), .Z(n39552) );
  XNOR U41518 ( .A(n39549), .B(n30475), .Z(n39551) );
  XOR U41519 ( .A(n39553), .B(n39554), .Z(n30475) );
  AND U41520 ( .A(\modmult_1/xin[1023] ), .B(n39555), .Z(n39554) );
  IV U41521 ( .A(n39553), .Z(n39555) );
  XOR U41522 ( .A(n39556), .B(g_input[44]), .Z(n39553) );
  NAND U41523 ( .A(n39557), .B(mul_pow), .Z(n39556) );
  XOR U41524 ( .A(g_input[44]), .B(creg[44]), .Z(n39557) );
  XOR U41525 ( .A(n39558), .B(n39559), .Z(n39549) );
  ANDN U41526 ( .A(n39560), .B(n30482), .Z(n39559) );
  XOR U41527 ( .A(n39561), .B(\modmult_1/zin[0][42] ), .Z(n30482) );
  IV U41528 ( .A(n39558), .Z(n39561) );
  XNOR U41529 ( .A(n39558), .B(n30481), .Z(n39560) );
  XOR U41530 ( .A(n39562), .B(n39563), .Z(n30481) );
  AND U41531 ( .A(\modmult_1/xin[1023] ), .B(n39564), .Z(n39563) );
  IV U41532 ( .A(n39562), .Z(n39564) );
  XOR U41533 ( .A(n39565), .B(g_input[43]), .Z(n39562) );
  NAND U41534 ( .A(n39566), .B(mul_pow), .Z(n39565) );
  XOR U41535 ( .A(g_input[43]), .B(creg[43]), .Z(n39566) );
  XOR U41536 ( .A(n39567), .B(n39568), .Z(n39558) );
  ANDN U41537 ( .A(n39569), .B(n30488), .Z(n39568) );
  XOR U41538 ( .A(n39570), .B(\modmult_1/zin[0][41] ), .Z(n30488) );
  IV U41539 ( .A(n39567), .Z(n39570) );
  XNOR U41540 ( .A(n39567), .B(n30487), .Z(n39569) );
  XOR U41541 ( .A(n39571), .B(n39572), .Z(n30487) );
  AND U41542 ( .A(\modmult_1/xin[1023] ), .B(n39573), .Z(n39572) );
  IV U41543 ( .A(n39571), .Z(n39573) );
  XOR U41544 ( .A(n39574), .B(g_input[42]), .Z(n39571) );
  NAND U41545 ( .A(n39575), .B(mul_pow), .Z(n39574) );
  XOR U41546 ( .A(g_input[42]), .B(creg[42]), .Z(n39575) );
  XOR U41547 ( .A(n39576), .B(n39577), .Z(n39567) );
  ANDN U41548 ( .A(n39578), .B(n30494), .Z(n39577) );
  XOR U41549 ( .A(n39579), .B(\modmult_1/zin[0][40] ), .Z(n30494) );
  IV U41550 ( .A(n39576), .Z(n39579) );
  XNOR U41551 ( .A(n39576), .B(n30493), .Z(n39578) );
  XOR U41552 ( .A(n39580), .B(n39581), .Z(n30493) );
  AND U41553 ( .A(\modmult_1/xin[1023] ), .B(n39582), .Z(n39581) );
  IV U41554 ( .A(n39580), .Z(n39582) );
  XOR U41555 ( .A(n39583), .B(g_input[41]), .Z(n39580) );
  NAND U41556 ( .A(n39584), .B(mul_pow), .Z(n39583) );
  XOR U41557 ( .A(g_input[41]), .B(creg[41]), .Z(n39584) );
  XOR U41558 ( .A(n39585), .B(n39586), .Z(n39576) );
  ANDN U41559 ( .A(n39587), .B(n30500), .Z(n39586) );
  XOR U41560 ( .A(n39588), .B(\modmult_1/zin[0][39] ), .Z(n30500) );
  IV U41561 ( .A(n39585), .Z(n39588) );
  XNOR U41562 ( .A(n39585), .B(n30499), .Z(n39587) );
  XOR U41563 ( .A(n39589), .B(n39590), .Z(n30499) );
  AND U41564 ( .A(\modmult_1/xin[1023] ), .B(n39591), .Z(n39590) );
  IV U41565 ( .A(n39589), .Z(n39591) );
  XOR U41566 ( .A(n39592), .B(g_input[40]), .Z(n39589) );
  NAND U41567 ( .A(n39593), .B(mul_pow), .Z(n39592) );
  XOR U41568 ( .A(g_input[40]), .B(creg[40]), .Z(n39593) );
  XOR U41569 ( .A(n39594), .B(n39595), .Z(n39585) );
  ANDN U41570 ( .A(n39596), .B(n30506), .Z(n39595) );
  XOR U41571 ( .A(n39597), .B(\modmult_1/zin[0][38] ), .Z(n30506) );
  IV U41572 ( .A(n39594), .Z(n39597) );
  XNOR U41573 ( .A(n39594), .B(n30505), .Z(n39596) );
  XOR U41574 ( .A(n39598), .B(n39599), .Z(n30505) );
  AND U41575 ( .A(\modmult_1/xin[1023] ), .B(n39600), .Z(n39599) );
  IV U41576 ( .A(n39598), .Z(n39600) );
  XOR U41577 ( .A(n39601), .B(g_input[39]), .Z(n39598) );
  NAND U41578 ( .A(n39602), .B(mul_pow), .Z(n39601) );
  XOR U41579 ( .A(g_input[39]), .B(creg[39]), .Z(n39602) );
  XOR U41580 ( .A(n39603), .B(n39604), .Z(n39594) );
  ANDN U41581 ( .A(n39605), .B(n30512), .Z(n39604) );
  XOR U41582 ( .A(n39606), .B(\modmult_1/zin[0][37] ), .Z(n30512) );
  IV U41583 ( .A(n39603), .Z(n39606) );
  XNOR U41584 ( .A(n39603), .B(n30511), .Z(n39605) );
  XOR U41585 ( .A(n39607), .B(n39608), .Z(n30511) );
  AND U41586 ( .A(\modmult_1/xin[1023] ), .B(n39609), .Z(n39608) );
  IV U41587 ( .A(n39607), .Z(n39609) );
  XOR U41588 ( .A(n39610), .B(g_input[38]), .Z(n39607) );
  NAND U41589 ( .A(n39611), .B(mul_pow), .Z(n39610) );
  XOR U41590 ( .A(g_input[38]), .B(creg[38]), .Z(n39611) );
  XOR U41591 ( .A(n39612), .B(n39613), .Z(n39603) );
  ANDN U41592 ( .A(n39614), .B(n30518), .Z(n39613) );
  XOR U41593 ( .A(n39615), .B(\modmult_1/zin[0][36] ), .Z(n30518) );
  IV U41594 ( .A(n39612), .Z(n39615) );
  XNOR U41595 ( .A(n39612), .B(n30517), .Z(n39614) );
  XOR U41596 ( .A(n39616), .B(n39617), .Z(n30517) );
  AND U41597 ( .A(\modmult_1/xin[1023] ), .B(n39618), .Z(n39617) );
  IV U41598 ( .A(n39616), .Z(n39618) );
  XOR U41599 ( .A(n39619), .B(g_input[37]), .Z(n39616) );
  NAND U41600 ( .A(n39620), .B(mul_pow), .Z(n39619) );
  XOR U41601 ( .A(g_input[37]), .B(creg[37]), .Z(n39620) );
  XOR U41602 ( .A(n39621), .B(n39622), .Z(n39612) );
  ANDN U41603 ( .A(n39623), .B(n30524), .Z(n39622) );
  XOR U41604 ( .A(n39624), .B(\modmult_1/zin[0][35] ), .Z(n30524) );
  IV U41605 ( .A(n39621), .Z(n39624) );
  XNOR U41606 ( .A(n39621), .B(n30523), .Z(n39623) );
  XOR U41607 ( .A(n39625), .B(n39626), .Z(n30523) );
  AND U41608 ( .A(\modmult_1/xin[1023] ), .B(n39627), .Z(n39626) );
  IV U41609 ( .A(n39625), .Z(n39627) );
  XOR U41610 ( .A(n39628), .B(g_input[36]), .Z(n39625) );
  NAND U41611 ( .A(n39629), .B(mul_pow), .Z(n39628) );
  XOR U41612 ( .A(g_input[36]), .B(creg[36]), .Z(n39629) );
  XOR U41613 ( .A(n39630), .B(n39631), .Z(n39621) );
  ANDN U41614 ( .A(n39632), .B(n30530), .Z(n39631) );
  XOR U41615 ( .A(n39633), .B(\modmult_1/zin[0][34] ), .Z(n30530) );
  IV U41616 ( .A(n39630), .Z(n39633) );
  XNOR U41617 ( .A(n39630), .B(n30529), .Z(n39632) );
  XOR U41618 ( .A(n39634), .B(n39635), .Z(n30529) );
  AND U41619 ( .A(\modmult_1/xin[1023] ), .B(n39636), .Z(n39635) );
  IV U41620 ( .A(n39634), .Z(n39636) );
  XOR U41621 ( .A(n39637), .B(g_input[35]), .Z(n39634) );
  NAND U41622 ( .A(n39638), .B(mul_pow), .Z(n39637) );
  XOR U41623 ( .A(g_input[35]), .B(creg[35]), .Z(n39638) );
  XOR U41624 ( .A(n39639), .B(n39640), .Z(n39630) );
  ANDN U41625 ( .A(n39641), .B(n30536), .Z(n39640) );
  XOR U41626 ( .A(n39642), .B(\modmult_1/zin[0][33] ), .Z(n30536) );
  IV U41627 ( .A(n39639), .Z(n39642) );
  XNOR U41628 ( .A(n39639), .B(n30535), .Z(n39641) );
  XOR U41629 ( .A(n39643), .B(n39644), .Z(n30535) );
  AND U41630 ( .A(\modmult_1/xin[1023] ), .B(n39645), .Z(n39644) );
  IV U41631 ( .A(n39643), .Z(n39645) );
  XOR U41632 ( .A(n39646), .B(g_input[34]), .Z(n39643) );
  NAND U41633 ( .A(n39647), .B(mul_pow), .Z(n39646) );
  XOR U41634 ( .A(g_input[34]), .B(creg[34]), .Z(n39647) );
  XOR U41635 ( .A(n39648), .B(n39649), .Z(n39639) );
  ANDN U41636 ( .A(n39650), .B(n30542), .Z(n39649) );
  XOR U41637 ( .A(n39651), .B(\modmult_1/zin[0][32] ), .Z(n30542) );
  IV U41638 ( .A(n39648), .Z(n39651) );
  XNOR U41639 ( .A(n39648), .B(n30541), .Z(n39650) );
  XOR U41640 ( .A(n39652), .B(n39653), .Z(n30541) );
  AND U41641 ( .A(\modmult_1/xin[1023] ), .B(n39654), .Z(n39653) );
  IV U41642 ( .A(n39652), .Z(n39654) );
  XOR U41643 ( .A(n39655), .B(g_input[33]), .Z(n39652) );
  NAND U41644 ( .A(n39656), .B(mul_pow), .Z(n39655) );
  XOR U41645 ( .A(g_input[33]), .B(creg[33]), .Z(n39656) );
  XOR U41646 ( .A(n39657), .B(n39658), .Z(n39648) );
  ANDN U41647 ( .A(n39659), .B(n30548), .Z(n39658) );
  XOR U41648 ( .A(n39660), .B(\modmult_1/zin[0][31] ), .Z(n30548) );
  IV U41649 ( .A(n39657), .Z(n39660) );
  XNOR U41650 ( .A(n39657), .B(n30547), .Z(n39659) );
  XOR U41651 ( .A(n39661), .B(n39662), .Z(n30547) );
  AND U41652 ( .A(\modmult_1/xin[1023] ), .B(n39663), .Z(n39662) );
  IV U41653 ( .A(n39661), .Z(n39663) );
  XOR U41654 ( .A(n39664), .B(g_input[32]), .Z(n39661) );
  NAND U41655 ( .A(n39665), .B(mul_pow), .Z(n39664) );
  XOR U41656 ( .A(g_input[32]), .B(creg[32]), .Z(n39665) );
  XOR U41657 ( .A(n39666), .B(n39667), .Z(n39657) );
  ANDN U41658 ( .A(n39668), .B(n30554), .Z(n39667) );
  XOR U41659 ( .A(n39669), .B(\modmult_1/zin[0][30] ), .Z(n30554) );
  IV U41660 ( .A(n39666), .Z(n39669) );
  XNOR U41661 ( .A(n39666), .B(n30553), .Z(n39668) );
  XOR U41662 ( .A(n39670), .B(n39671), .Z(n30553) );
  AND U41663 ( .A(\modmult_1/xin[1023] ), .B(n39672), .Z(n39671) );
  IV U41664 ( .A(n39670), .Z(n39672) );
  XOR U41665 ( .A(n39673), .B(g_input[31]), .Z(n39670) );
  NAND U41666 ( .A(n39674), .B(mul_pow), .Z(n39673) );
  XOR U41667 ( .A(g_input[31]), .B(creg[31]), .Z(n39674) );
  XOR U41668 ( .A(n39675), .B(n39676), .Z(n39666) );
  ANDN U41669 ( .A(n39677), .B(n30560), .Z(n39676) );
  XOR U41670 ( .A(n39678), .B(\modmult_1/zin[0][29] ), .Z(n30560) );
  IV U41671 ( .A(n39675), .Z(n39678) );
  XNOR U41672 ( .A(n39675), .B(n30559), .Z(n39677) );
  XOR U41673 ( .A(n39679), .B(n39680), .Z(n30559) );
  AND U41674 ( .A(\modmult_1/xin[1023] ), .B(n39681), .Z(n39680) );
  IV U41675 ( .A(n39679), .Z(n39681) );
  XOR U41676 ( .A(n39682), .B(g_input[30]), .Z(n39679) );
  NAND U41677 ( .A(n39683), .B(mul_pow), .Z(n39682) );
  XOR U41678 ( .A(g_input[30]), .B(creg[30]), .Z(n39683) );
  XOR U41679 ( .A(n39684), .B(n39685), .Z(n39675) );
  ANDN U41680 ( .A(n39686), .B(n30566), .Z(n39685) );
  XOR U41681 ( .A(n39687), .B(\modmult_1/zin[0][28] ), .Z(n30566) );
  IV U41682 ( .A(n39684), .Z(n39687) );
  XNOR U41683 ( .A(n39684), .B(n30565), .Z(n39686) );
  XOR U41684 ( .A(n39688), .B(n39689), .Z(n30565) );
  AND U41685 ( .A(\modmult_1/xin[1023] ), .B(n39690), .Z(n39689) );
  IV U41686 ( .A(n39688), .Z(n39690) );
  XOR U41687 ( .A(n39691), .B(g_input[29]), .Z(n39688) );
  NAND U41688 ( .A(n39692), .B(mul_pow), .Z(n39691) );
  XOR U41689 ( .A(g_input[29]), .B(creg[29]), .Z(n39692) );
  XOR U41690 ( .A(n39693), .B(n39694), .Z(n39684) );
  ANDN U41691 ( .A(n39695), .B(n30572), .Z(n39694) );
  XOR U41692 ( .A(n39696), .B(\modmult_1/zin[0][27] ), .Z(n30572) );
  IV U41693 ( .A(n39693), .Z(n39696) );
  XNOR U41694 ( .A(n39693), .B(n30571), .Z(n39695) );
  XOR U41695 ( .A(n39697), .B(n39698), .Z(n30571) );
  AND U41696 ( .A(\modmult_1/xin[1023] ), .B(n39699), .Z(n39698) );
  IV U41697 ( .A(n39697), .Z(n39699) );
  XOR U41698 ( .A(n39700), .B(g_input[28]), .Z(n39697) );
  NAND U41699 ( .A(n39701), .B(mul_pow), .Z(n39700) );
  XOR U41700 ( .A(g_input[28]), .B(creg[28]), .Z(n39701) );
  XOR U41701 ( .A(n39702), .B(n39703), .Z(n39693) );
  ANDN U41702 ( .A(n39704), .B(n30578), .Z(n39703) );
  XOR U41703 ( .A(n39705), .B(\modmult_1/zin[0][26] ), .Z(n30578) );
  IV U41704 ( .A(n39702), .Z(n39705) );
  XNOR U41705 ( .A(n39702), .B(n30577), .Z(n39704) );
  XOR U41706 ( .A(n39706), .B(n39707), .Z(n30577) );
  AND U41707 ( .A(\modmult_1/xin[1023] ), .B(n39708), .Z(n39707) );
  IV U41708 ( .A(n39706), .Z(n39708) );
  XOR U41709 ( .A(n39709), .B(g_input[27]), .Z(n39706) );
  NAND U41710 ( .A(n39710), .B(mul_pow), .Z(n39709) );
  XOR U41711 ( .A(g_input[27]), .B(creg[27]), .Z(n39710) );
  XOR U41712 ( .A(n39711), .B(n39712), .Z(n39702) );
  ANDN U41713 ( .A(n39713), .B(n30584), .Z(n39712) );
  XOR U41714 ( .A(n39714), .B(\modmult_1/zin[0][25] ), .Z(n30584) );
  IV U41715 ( .A(n39711), .Z(n39714) );
  XNOR U41716 ( .A(n39711), .B(n30583), .Z(n39713) );
  XOR U41717 ( .A(n39715), .B(n39716), .Z(n30583) );
  AND U41718 ( .A(\modmult_1/xin[1023] ), .B(n39717), .Z(n39716) );
  IV U41719 ( .A(n39715), .Z(n39717) );
  XOR U41720 ( .A(n39718), .B(g_input[26]), .Z(n39715) );
  NAND U41721 ( .A(n39719), .B(mul_pow), .Z(n39718) );
  XOR U41722 ( .A(g_input[26]), .B(creg[26]), .Z(n39719) );
  XOR U41723 ( .A(n39720), .B(n39721), .Z(n39711) );
  ANDN U41724 ( .A(n39722), .B(n30590), .Z(n39721) );
  XOR U41725 ( .A(n39723), .B(\modmult_1/zin[0][24] ), .Z(n30590) );
  IV U41726 ( .A(n39720), .Z(n39723) );
  XNOR U41727 ( .A(n39720), .B(n30589), .Z(n39722) );
  XOR U41728 ( .A(n39724), .B(n39725), .Z(n30589) );
  AND U41729 ( .A(\modmult_1/xin[1023] ), .B(n39726), .Z(n39725) );
  IV U41730 ( .A(n39724), .Z(n39726) );
  XOR U41731 ( .A(n39727), .B(g_input[25]), .Z(n39724) );
  NAND U41732 ( .A(n39728), .B(mul_pow), .Z(n39727) );
  XOR U41733 ( .A(g_input[25]), .B(creg[25]), .Z(n39728) );
  XOR U41734 ( .A(n39729), .B(n39730), .Z(n39720) );
  ANDN U41735 ( .A(n39731), .B(n30596), .Z(n39730) );
  XOR U41736 ( .A(n39732), .B(\modmult_1/zin[0][23] ), .Z(n30596) );
  IV U41737 ( .A(n39729), .Z(n39732) );
  XNOR U41738 ( .A(n39729), .B(n30595), .Z(n39731) );
  XOR U41739 ( .A(n39733), .B(n39734), .Z(n30595) );
  AND U41740 ( .A(\modmult_1/xin[1023] ), .B(n39735), .Z(n39734) );
  IV U41741 ( .A(n39733), .Z(n39735) );
  XOR U41742 ( .A(n39736), .B(g_input[24]), .Z(n39733) );
  NAND U41743 ( .A(n39737), .B(mul_pow), .Z(n39736) );
  XOR U41744 ( .A(g_input[24]), .B(creg[24]), .Z(n39737) );
  XOR U41745 ( .A(n39738), .B(n39739), .Z(n39729) );
  ANDN U41746 ( .A(n39740), .B(n30602), .Z(n39739) );
  XOR U41747 ( .A(n39741), .B(\modmult_1/zin[0][22] ), .Z(n30602) );
  IV U41748 ( .A(n39738), .Z(n39741) );
  XNOR U41749 ( .A(n39738), .B(n30601), .Z(n39740) );
  XOR U41750 ( .A(n39742), .B(n39743), .Z(n30601) );
  AND U41751 ( .A(\modmult_1/xin[1023] ), .B(n39744), .Z(n39743) );
  IV U41752 ( .A(n39742), .Z(n39744) );
  XOR U41753 ( .A(n39745), .B(g_input[23]), .Z(n39742) );
  NAND U41754 ( .A(n39746), .B(mul_pow), .Z(n39745) );
  XOR U41755 ( .A(g_input[23]), .B(creg[23]), .Z(n39746) );
  XOR U41756 ( .A(n39747), .B(n39748), .Z(n39738) );
  ANDN U41757 ( .A(n39749), .B(n30608), .Z(n39748) );
  XOR U41758 ( .A(n39750), .B(\modmult_1/zin[0][21] ), .Z(n30608) );
  IV U41759 ( .A(n39747), .Z(n39750) );
  XNOR U41760 ( .A(n39747), .B(n30607), .Z(n39749) );
  XOR U41761 ( .A(n39751), .B(n39752), .Z(n30607) );
  AND U41762 ( .A(\modmult_1/xin[1023] ), .B(n39753), .Z(n39752) );
  IV U41763 ( .A(n39751), .Z(n39753) );
  XOR U41764 ( .A(n39754), .B(g_input[22]), .Z(n39751) );
  NAND U41765 ( .A(n39755), .B(mul_pow), .Z(n39754) );
  XOR U41766 ( .A(g_input[22]), .B(creg[22]), .Z(n39755) );
  XOR U41767 ( .A(n39756), .B(n39757), .Z(n39747) );
  ANDN U41768 ( .A(n39758), .B(n30614), .Z(n39757) );
  XOR U41769 ( .A(n39759), .B(\modmult_1/zin[0][20] ), .Z(n30614) );
  IV U41770 ( .A(n39756), .Z(n39759) );
  XNOR U41771 ( .A(n39756), .B(n30613), .Z(n39758) );
  XOR U41772 ( .A(n39760), .B(n39761), .Z(n30613) );
  AND U41773 ( .A(\modmult_1/xin[1023] ), .B(n39762), .Z(n39761) );
  IV U41774 ( .A(n39760), .Z(n39762) );
  XOR U41775 ( .A(n39763), .B(g_input[21]), .Z(n39760) );
  NAND U41776 ( .A(n39764), .B(mul_pow), .Z(n39763) );
  XOR U41777 ( .A(g_input[21]), .B(creg[21]), .Z(n39764) );
  XOR U41778 ( .A(n39765), .B(n39766), .Z(n39756) );
  ANDN U41779 ( .A(n39767), .B(n30620), .Z(n39766) );
  XOR U41780 ( .A(n39768), .B(\modmult_1/zin[0][19] ), .Z(n30620) );
  IV U41781 ( .A(n39765), .Z(n39768) );
  XNOR U41782 ( .A(n39765), .B(n30619), .Z(n39767) );
  XOR U41783 ( .A(n39769), .B(n39770), .Z(n30619) );
  AND U41784 ( .A(\modmult_1/xin[1023] ), .B(n39771), .Z(n39770) );
  IV U41785 ( .A(n39769), .Z(n39771) );
  XOR U41786 ( .A(n39772), .B(g_input[20]), .Z(n39769) );
  NAND U41787 ( .A(n39773), .B(mul_pow), .Z(n39772) );
  XOR U41788 ( .A(g_input[20]), .B(creg[20]), .Z(n39773) );
  XOR U41789 ( .A(n39774), .B(n39775), .Z(n39765) );
  ANDN U41790 ( .A(n39776), .B(n30626), .Z(n39775) );
  XOR U41791 ( .A(n39777), .B(\modmult_1/zin[0][18] ), .Z(n30626) );
  IV U41792 ( .A(n39774), .Z(n39777) );
  XNOR U41793 ( .A(n39774), .B(n30625), .Z(n39776) );
  XOR U41794 ( .A(n39778), .B(n39779), .Z(n30625) );
  AND U41795 ( .A(\modmult_1/xin[1023] ), .B(n39780), .Z(n39779) );
  IV U41796 ( .A(n39778), .Z(n39780) );
  XOR U41797 ( .A(n39781), .B(g_input[19]), .Z(n39778) );
  NAND U41798 ( .A(n39782), .B(mul_pow), .Z(n39781) );
  XOR U41799 ( .A(g_input[19]), .B(creg[19]), .Z(n39782) );
  XOR U41800 ( .A(n39783), .B(n39784), .Z(n39774) );
  ANDN U41801 ( .A(n39785), .B(n30632), .Z(n39784) );
  XOR U41802 ( .A(n39786), .B(\modmult_1/zin[0][17] ), .Z(n30632) );
  IV U41803 ( .A(n39783), .Z(n39786) );
  XNOR U41804 ( .A(n39783), .B(n30631), .Z(n39785) );
  XOR U41805 ( .A(n39787), .B(n39788), .Z(n30631) );
  AND U41806 ( .A(\modmult_1/xin[1023] ), .B(n39789), .Z(n39788) );
  IV U41807 ( .A(n39787), .Z(n39789) );
  XOR U41808 ( .A(n39790), .B(g_input[18]), .Z(n39787) );
  NAND U41809 ( .A(n39791), .B(mul_pow), .Z(n39790) );
  XOR U41810 ( .A(g_input[18]), .B(creg[18]), .Z(n39791) );
  XOR U41811 ( .A(n39792), .B(n39793), .Z(n39783) );
  ANDN U41812 ( .A(n39794), .B(n30638), .Z(n39793) );
  XOR U41813 ( .A(n39795), .B(\modmult_1/zin[0][16] ), .Z(n30638) );
  IV U41814 ( .A(n39792), .Z(n39795) );
  XNOR U41815 ( .A(n39792), .B(n30637), .Z(n39794) );
  XOR U41816 ( .A(n39796), .B(n39797), .Z(n30637) );
  AND U41817 ( .A(\modmult_1/xin[1023] ), .B(n39798), .Z(n39797) );
  IV U41818 ( .A(n39796), .Z(n39798) );
  XOR U41819 ( .A(n39799), .B(g_input[17]), .Z(n39796) );
  NAND U41820 ( .A(n39800), .B(mul_pow), .Z(n39799) );
  XOR U41821 ( .A(g_input[17]), .B(creg[17]), .Z(n39800) );
  XOR U41822 ( .A(n39801), .B(n39802), .Z(n39792) );
  ANDN U41823 ( .A(n39803), .B(n30644), .Z(n39802) );
  XOR U41824 ( .A(n39804), .B(\modmult_1/zin[0][15] ), .Z(n30644) );
  IV U41825 ( .A(n39801), .Z(n39804) );
  XNOR U41826 ( .A(n39801), .B(n30643), .Z(n39803) );
  XOR U41827 ( .A(n39805), .B(n39806), .Z(n30643) );
  AND U41828 ( .A(\modmult_1/xin[1023] ), .B(n39807), .Z(n39806) );
  IV U41829 ( .A(n39805), .Z(n39807) );
  XOR U41830 ( .A(n39808), .B(g_input[16]), .Z(n39805) );
  NAND U41831 ( .A(n39809), .B(mul_pow), .Z(n39808) );
  XOR U41832 ( .A(g_input[16]), .B(creg[16]), .Z(n39809) );
  XOR U41833 ( .A(n39810), .B(n39811), .Z(n39801) );
  ANDN U41834 ( .A(n39812), .B(n30650), .Z(n39811) );
  XOR U41835 ( .A(n39813), .B(\modmult_1/zin[0][14] ), .Z(n30650) );
  IV U41836 ( .A(n39810), .Z(n39813) );
  XNOR U41837 ( .A(n39810), .B(n30649), .Z(n39812) );
  XOR U41838 ( .A(n39814), .B(n39815), .Z(n30649) );
  AND U41839 ( .A(\modmult_1/xin[1023] ), .B(n39816), .Z(n39815) );
  IV U41840 ( .A(n39814), .Z(n39816) );
  XOR U41841 ( .A(n39817), .B(g_input[15]), .Z(n39814) );
  NAND U41842 ( .A(n39818), .B(mul_pow), .Z(n39817) );
  XOR U41843 ( .A(g_input[15]), .B(creg[15]), .Z(n39818) );
  XOR U41844 ( .A(n39819), .B(n39820), .Z(n39810) );
  ANDN U41845 ( .A(n39821), .B(n30656), .Z(n39820) );
  XOR U41846 ( .A(n39822), .B(\modmult_1/zin[0][13] ), .Z(n30656) );
  IV U41847 ( .A(n39819), .Z(n39822) );
  XNOR U41848 ( .A(n39819), .B(n30655), .Z(n39821) );
  XOR U41849 ( .A(n39823), .B(n39824), .Z(n30655) );
  AND U41850 ( .A(\modmult_1/xin[1023] ), .B(n39825), .Z(n39824) );
  IV U41851 ( .A(n39823), .Z(n39825) );
  XOR U41852 ( .A(n39826), .B(g_input[14]), .Z(n39823) );
  NAND U41853 ( .A(n39827), .B(mul_pow), .Z(n39826) );
  XOR U41854 ( .A(g_input[14]), .B(creg[14]), .Z(n39827) );
  XOR U41855 ( .A(n39828), .B(n39829), .Z(n39819) );
  ANDN U41856 ( .A(n39830), .B(n30662), .Z(n39829) );
  XOR U41857 ( .A(n39831), .B(\modmult_1/zin[0][12] ), .Z(n30662) );
  IV U41858 ( .A(n39828), .Z(n39831) );
  XNOR U41859 ( .A(n39828), .B(n30661), .Z(n39830) );
  XOR U41860 ( .A(n39832), .B(n39833), .Z(n30661) );
  AND U41861 ( .A(\modmult_1/xin[1023] ), .B(n39834), .Z(n39833) );
  IV U41862 ( .A(n39832), .Z(n39834) );
  XOR U41863 ( .A(n39835), .B(g_input[13]), .Z(n39832) );
  NAND U41864 ( .A(n39836), .B(mul_pow), .Z(n39835) );
  XOR U41865 ( .A(g_input[13]), .B(creg[13]), .Z(n39836) );
  XOR U41866 ( .A(n39837), .B(n39838), .Z(n39828) );
  ANDN U41867 ( .A(n39839), .B(n30668), .Z(n39838) );
  XOR U41868 ( .A(n39840), .B(\modmult_1/zin[0][11] ), .Z(n30668) );
  IV U41869 ( .A(n39837), .Z(n39840) );
  XNOR U41870 ( .A(n39837), .B(n30667), .Z(n39839) );
  XOR U41871 ( .A(n39841), .B(n39842), .Z(n30667) );
  AND U41872 ( .A(\modmult_1/xin[1023] ), .B(n39843), .Z(n39842) );
  IV U41873 ( .A(n39841), .Z(n39843) );
  XOR U41874 ( .A(n39844), .B(g_input[12]), .Z(n39841) );
  NAND U41875 ( .A(n39845), .B(mul_pow), .Z(n39844) );
  XOR U41876 ( .A(g_input[12]), .B(creg[12]), .Z(n39845) );
  XOR U41877 ( .A(n39846), .B(n39847), .Z(n39837) );
  ANDN U41878 ( .A(n39848), .B(n30674), .Z(n39847) );
  XOR U41879 ( .A(n39849), .B(\modmult_1/zin[0][10] ), .Z(n30674) );
  IV U41880 ( .A(n39846), .Z(n39849) );
  XNOR U41881 ( .A(n39846), .B(n30673), .Z(n39848) );
  XOR U41882 ( .A(n39850), .B(n39851), .Z(n30673) );
  AND U41883 ( .A(\modmult_1/xin[1023] ), .B(n39852), .Z(n39851) );
  IV U41884 ( .A(n39850), .Z(n39852) );
  XOR U41885 ( .A(n39853), .B(g_input[11]), .Z(n39850) );
  NAND U41886 ( .A(n39854), .B(mul_pow), .Z(n39853) );
  XOR U41887 ( .A(g_input[11]), .B(creg[11]), .Z(n39854) );
  XOR U41888 ( .A(n39855), .B(n39856), .Z(n39846) );
  ANDN U41889 ( .A(n39857), .B(n30680), .Z(n39856) );
  XOR U41890 ( .A(n39858), .B(\modmult_1/zin[0][9] ), .Z(n30680) );
  IV U41891 ( .A(n39855), .Z(n39858) );
  XNOR U41892 ( .A(n39855), .B(n30679), .Z(n39857) );
  XOR U41893 ( .A(n39859), .B(n39860), .Z(n30679) );
  AND U41894 ( .A(\modmult_1/xin[1023] ), .B(n39861), .Z(n39860) );
  IV U41895 ( .A(n39859), .Z(n39861) );
  XOR U41896 ( .A(n39862), .B(g_input[10]), .Z(n39859) );
  NAND U41897 ( .A(n39863), .B(mul_pow), .Z(n39862) );
  XOR U41898 ( .A(g_input[10]), .B(creg[10]), .Z(n39863) );
  XOR U41899 ( .A(n39864), .B(n39865), .Z(n39855) );
  ANDN U41900 ( .A(n39866), .B(n30686), .Z(n39865) );
  XOR U41901 ( .A(n39867), .B(\modmult_1/zin[0][8] ), .Z(n30686) );
  IV U41902 ( .A(n39864), .Z(n39867) );
  XNOR U41903 ( .A(n39864), .B(n30685), .Z(n39866) );
  XOR U41904 ( .A(n39868), .B(n39869), .Z(n30685) );
  AND U41905 ( .A(\modmult_1/xin[1023] ), .B(n39870), .Z(n39869) );
  IV U41906 ( .A(n39868), .Z(n39870) );
  XOR U41907 ( .A(n39871), .B(g_input[9]), .Z(n39868) );
  NAND U41908 ( .A(n39872), .B(mul_pow), .Z(n39871) );
  XOR U41909 ( .A(g_input[9]), .B(creg[9]), .Z(n39872) );
  XOR U41910 ( .A(n39873), .B(n39874), .Z(n39864) );
  ANDN U41911 ( .A(n39875), .B(n30692), .Z(n39874) );
  XOR U41912 ( .A(n39876), .B(\modmult_1/zin[0][7] ), .Z(n30692) );
  IV U41913 ( .A(n39873), .Z(n39876) );
  XNOR U41914 ( .A(n39873), .B(n30691), .Z(n39875) );
  XOR U41915 ( .A(n39877), .B(n39878), .Z(n30691) );
  AND U41916 ( .A(\modmult_1/xin[1023] ), .B(n39879), .Z(n39878) );
  IV U41917 ( .A(n39877), .Z(n39879) );
  XOR U41918 ( .A(n39880), .B(g_input[8]), .Z(n39877) );
  NAND U41919 ( .A(n39881), .B(mul_pow), .Z(n39880) );
  XOR U41920 ( .A(g_input[8]), .B(creg[8]), .Z(n39881) );
  XOR U41921 ( .A(n39882), .B(n39883), .Z(n39873) );
  ANDN U41922 ( .A(n39884), .B(n30698), .Z(n39883) );
  XOR U41923 ( .A(n39885), .B(\modmult_1/zin[0][6] ), .Z(n30698) );
  IV U41924 ( .A(n39882), .Z(n39885) );
  XNOR U41925 ( .A(n39882), .B(n30697), .Z(n39884) );
  XOR U41926 ( .A(n39886), .B(n39887), .Z(n30697) );
  AND U41927 ( .A(\modmult_1/xin[1023] ), .B(n39888), .Z(n39887) );
  IV U41928 ( .A(n39886), .Z(n39888) );
  XOR U41929 ( .A(n39889), .B(g_input[7]), .Z(n39886) );
  NAND U41930 ( .A(n39890), .B(mul_pow), .Z(n39889) );
  XOR U41931 ( .A(g_input[7]), .B(creg[7]), .Z(n39890) );
  XOR U41932 ( .A(n39891), .B(n39892), .Z(n39882) );
  ANDN U41933 ( .A(n39893), .B(n30704), .Z(n39892) );
  XOR U41934 ( .A(n39894), .B(\modmult_1/zin[0][5] ), .Z(n30704) );
  IV U41935 ( .A(n39891), .Z(n39894) );
  XNOR U41936 ( .A(n39891), .B(n30703), .Z(n39893) );
  XOR U41937 ( .A(n39895), .B(n39896), .Z(n30703) );
  AND U41938 ( .A(\modmult_1/xin[1023] ), .B(n39897), .Z(n39896) );
  IV U41939 ( .A(n39895), .Z(n39897) );
  XOR U41940 ( .A(n39898), .B(g_input[6]), .Z(n39895) );
  NAND U41941 ( .A(n39899), .B(mul_pow), .Z(n39898) );
  XOR U41942 ( .A(g_input[6]), .B(creg[6]), .Z(n39899) );
  XOR U41943 ( .A(n39900), .B(n39901), .Z(n39891) );
  ANDN U41944 ( .A(n39902), .B(n30710), .Z(n39901) );
  XOR U41945 ( .A(n39903), .B(\modmult_1/zin[0][4] ), .Z(n30710) );
  IV U41946 ( .A(n39900), .Z(n39903) );
  XNOR U41947 ( .A(n39900), .B(n30709), .Z(n39902) );
  XOR U41948 ( .A(n39904), .B(n39905), .Z(n30709) );
  AND U41949 ( .A(\modmult_1/xin[1023] ), .B(n39906), .Z(n39905) );
  IV U41950 ( .A(n39904), .Z(n39906) );
  XOR U41951 ( .A(n39907), .B(g_input[5]), .Z(n39904) );
  NAND U41952 ( .A(n39908), .B(mul_pow), .Z(n39907) );
  XOR U41953 ( .A(g_input[5]), .B(creg[5]), .Z(n39908) );
  XOR U41954 ( .A(n39909), .B(n39910), .Z(n39900) );
  ANDN U41955 ( .A(n39911), .B(n30716), .Z(n39910) );
  XOR U41956 ( .A(n39912), .B(\modmult_1/zin[0][3] ), .Z(n30716) );
  IV U41957 ( .A(n39909), .Z(n39912) );
  XNOR U41958 ( .A(n39909), .B(n30715), .Z(n39911) );
  XOR U41959 ( .A(n39913), .B(n39914), .Z(n30715) );
  AND U41960 ( .A(\modmult_1/xin[1023] ), .B(n39915), .Z(n39914) );
  IV U41961 ( .A(n39913), .Z(n39915) );
  XOR U41962 ( .A(n39916), .B(g_input[4]), .Z(n39913) );
  NAND U41963 ( .A(n39917), .B(mul_pow), .Z(n39916) );
  XOR U41964 ( .A(g_input[4]), .B(creg[4]), .Z(n39917) );
  XNOR U41965 ( .A(n39918), .B(n39919), .Z(n39909) );
  ANDN U41966 ( .A(n39920), .B(n30722), .Z(n39919) );
  XOR U41967 ( .A(n39918), .B(\modmult_1/zin[0][2] ), .Z(n30722) );
  XOR U41968 ( .A(n39918), .B(n30721), .Z(n39920) );
  XOR U41969 ( .A(n39921), .B(n39922), .Z(n30721) );
  AND U41970 ( .A(\modmult_1/xin[1023] ), .B(n39923), .Z(n39922) );
  IV U41971 ( .A(n39921), .Z(n39923) );
  XOR U41972 ( .A(n39924), .B(g_input[3]), .Z(n39921) );
  NAND U41973 ( .A(n39925), .B(mul_pow), .Z(n39924) );
  XOR U41974 ( .A(g_input[3]), .B(creg[3]), .Z(n39925) );
  XOR U41975 ( .A(n39926), .B(n39927), .Z(n39918) );
  NAND U41976 ( .A(n39928), .B(n30728), .Z(n39926) );
  XNOR U41977 ( .A(n39929), .B(\modmult_1/zin[0][1] ), .Z(n30728) );
  IV U41978 ( .A(n39927), .Z(n39929) );
  XNOR U41979 ( .A(n39927), .B(n30727), .Z(n39928) );
  XOR U41980 ( .A(n39930), .B(n39931), .Z(n30727) );
  AND U41981 ( .A(\modmult_1/xin[1023] ), .B(n39932), .Z(n39931) );
  IV U41982 ( .A(n39930), .Z(n39932) );
  XOR U41983 ( .A(n39933), .B(g_input[2]), .Z(n39930) );
  NAND U41984 ( .A(n39934), .B(mul_pow), .Z(n39933) );
  XOR U41985 ( .A(g_input[2]), .B(creg[2]), .Z(n39934) );
  ANDN U41986 ( .A(\modmult_1/zin[0][0] ), .B(n30734), .Z(n39927) );
  XOR U41987 ( .A(n39935), .B(n39936), .Z(n30734) );
  AND U41988 ( .A(\modmult_1/xin[1023] ), .B(n39937), .Z(n39936) );
  IV U41989 ( .A(n39935), .Z(n39937) );
  XOR U41990 ( .A(n39938), .B(g_input[1]), .Z(n39935) );
  NAND U41991 ( .A(n39939), .B(mul_pow), .Z(n39938) );
  XOR U41992 ( .A(g_input[1]), .B(creg[1]), .Z(n39939) );
  XOR U41993 ( .A(n39940), .B(n39941), .Z(n24588) );
  AND U41994 ( .A(n39940), .B(\modmult_1/xin[1023] ), .Z(n39941) );
  XNOR U41995 ( .A(n39942), .B(g_input[0]), .Z(n39940) );
  NAND U41996 ( .A(n39943), .B(mul_pow), .Z(n39942) );
  XOR U41997 ( .A(g_input[0]), .B(creg[0]), .Z(n39943) );
  XOR U41998 ( .A(ein[8]), .B(n39944), .Z(ereg_next[9]) );
  AND U41999 ( .A(mul_pow), .B(n39945), .Z(n39944) );
  XOR U42000 ( .A(ein[9]), .B(ein[8]), .Z(n39945) );
  XOR U42001 ( .A(ein[98]), .B(n39946), .Z(ereg_next[99]) );
  AND U42002 ( .A(mul_pow), .B(n39947), .Z(n39946) );
  XOR U42003 ( .A(ein[99]), .B(ein[98]), .Z(n39947) );
  XOR U42004 ( .A(ein[998]), .B(n39948), .Z(ereg_next[999]) );
  AND U42005 ( .A(mul_pow), .B(n39949), .Z(n39948) );
  XOR U42006 ( .A(ein[999]), .B(ein[998]), .Z(n39949) );
  XOR U42007 ( .A(ein[997]), .B(n39950), .Z(ereg_next[998]) );
  AND U42008 ( .A(mul_pow), .B(n39951), .Z(n39950) );
  XOR U42009 ( .A(ein[998]), .B(ein[997]), .Z(n39951) );
  XOR U42010 ( .A(ein[996]), .B(n39952), .Z(ereg_next[997]) );
  AND U42011 ( .A(mul_pow), .B(n39953), .Z(n39952) );
  XOR U42012 ( .A(ein[997]), .B(ein[996]), .Z(n39953) );
  XOR U42013 ( .A(ein[995]), .B(n39954), .Z(ereg_next[996]) );
  AND U42014 ( .A(mul_pow), .B(n39955), .Z(n39954) );
  XOR U42015 ( .A(ein[996]), .B(ein[995]), .Z(n39955) );
  XOR U42016 ( .A(ein[994]), .B(n39956), .Z(ereg_next[995]) );
  AND U42017 ( .A(mul_pow), .B(n39957), .Z(n39956) );
  XOR U42018 ( .A(ein[995]), .B(ein[994]), .Z(n39957) );
  XOR U42019 ( .A(ein[993]), .B(n39958), .Z(ereg_next[994]) );
  AND U42020 ( .A(mul_pow), .B(n39959), .Z(n39958) );
  XOR U42021 ( .A(ein[994]), .B(ein[993]), .Z(n39959) );
  XOR U42022 ( .A(ein[992]), .B(n39960), .Z(ereg_next[993]) );
  AND U42023 ( .A(mul_pow), .B(n39961), .Z(n39960) );
  XOR U42024 ( .A(ein[993]), .B(ein[992]), .Z(n39961) );
  XOR U42025 ( .A(ein[991]), .B(n39962), .Z(ereg_next[992]) );
  AND U42026 ( .A(mul_pow), .B(n39963), .Z(n39962) );
  XOR U42027 ( .A(ein[992]), .B(ein[991]), .Z(n39963) );
  XOR U42028 ( .A(ein[990]), .B(n39964), .Z(ereg_next[991]) );
  AND U42029 ( .A(mul_pow), .B(n39965), .Z(n39964) );
  XOR U42030 ( .A(ein[991]), .B(ein[990]), .Z(n39965) );
  XOR U42031 ( .A(ein[989]), .B(n39966), .Z(ereg_next[990]) );
  AND U42032 ( .A(mul_pow), .B(n39967), .Z(n39966) );
  XOR U42033 ( .A(ein[990]), .B(ein[989]), .Z(n39967) );
  XOR U42034 ( .A(ein[97]), .B(n39968), .Z(ereg_next[98]) );
  AND U42035 ( .A(mul_pow), .B(n39969), .Z(n39968) );
  XOR U42036 ( .A(ein[98]), .B(ein[97]), .Z(n39969) );
  XOR U42037 ( .A(ein[988]), .B(n39970), .Z(ereg_next[989]) );
  AND U42038 ( .A(mul_pow), .B(n39971), .Z(n39970) );
  XOR U42039 ( .A(ein[989]), .B(ein[988]), .Z(n39971) );
  XOR U42040 ( .A(ein[987]), .B(n39972), .Z(ereg_next[988]) );
  AND U42041 ( .A(mul_pow), .B(n39973), .Z(n39972) );
  XOR U42042 ( .A(ein[988]), .B(ein[987]), .Z(n39973) );
  XOR U42043 ( .A(ein[986]), .B(n39974), .Z(ereg_next[987]) );
  AND U42044 ( .A(mul_pow), .B(n39975), .Z(n39974) );
  XOR U42045 ( .A(ein[987]), .B(ein[986]), .Z(n39975) );
  XOR U42046 ( .A(ein[985]), .B(n39976), .Z(ereg_next[986]) );
  AND U42047 ( .A(mul_pow), .B(n39977), .Z(n39976) );
  XOR U42048 ( .A(ein[986]), .B(ein[985]), .Z(n39977) );
  XOR U42049 ( .A(ein[984]), .B(n39978), .Z(ereg_next[985]) );
  AND U42050 ( .A(mul_pow), .B(n39979), .Z(n39978) );
  XOR U42051 ( .A(ein[985]), .B(ein[984]), .Z(n39979) );
  XOR U42052 ( .A(ein[983]), .B(n39980), .Z(ereg_next[984]) );
  AND U42053 ( .A(mul_pow), .B(n39981), .Z(n39980) );
  XOR U42054 ( .A(ein[984]), .B(ein[983]), .Z(n39981) );
  XOR U42055 ( .A(ein[982]), .B(n39982), .Z(ereg_next[983]) );
  AND U42056 ( .A(mul_pow), .B(n39983), .Z(n39982) );
  XOR U42057 ( .A(ein[983]), .B(ein[982]), .Z(n39983) );
  XOR U42058 ( .A(ein[981]), .B(n39984), .Z(ereg_next[982]) );
  AND U42059 ( .A(mul_pow), .B(n39985), .Z(n39984) );
  XOR U42060 ( .A(ein[982]), .B(ein[981]), .Z(n39985) );
  XOR U42061 ( .A(ein[980]), .B(n39986), .Z(ereg_next[981]) );
  AND U42062 ( .A(mul_pow), .B(n39987), .Z(n39986) );
  XOR U42063 ( .A(ein[981]), .B(ein[980]), .Z(n39987) );
  XOR U42064 ( .A(ein[979]), .B(n39988), .Z(ereg_next[980]) );
  AND U42065 ( .A(mul_pow), .B(n39989), .Z(n39988) );
  XOR U42066 ( .A(ein[980]), .B(ein[979]), .Z(n39989) );
  XOR U42067 ( .A(ein[96]), .B(n39990), .Z(ereg_next[97]) );
  AND U42068 ( .A(mul_pow), .B(n39991), .Z(n39990) );
  XOR U42069 ( .A(ein[97]), .B(ein[96]), .Z(n39991) );
  XOR U42070 ( .A(ein[978]), .B(n39992), .Z(ereg_next[979]) );
  AND U42071 ( .A(mul_pow), .B(n39993), .Z(n39992) );
  XOR U42072 ( .A(ein[979]), .B(ein[978]), .Z(n39993) );
  XOR U42073 ( .A(ein[977]), .B(n39994), .Z(ereg_next[978]) );
  AND U42074 ( .A(mul_pow), .B(n39995), .Z(n39994) );
  XOR U42075 ( .A(ein[978]), .B(ein[977]), .Z(n39995) );
  XOR U42076 ( .A(ein[976]), .B(n39996), .Z(ereg_next[977]) );
  AND U42077 ( .A(mul_pow), .B(n39997), .Z(n39996) );
  XOR U42078 ( .A(ein[977]), .B(ein[976]), .Z(n39997) );
  XOR U42079 ( .A(ein[975]), .B(n39998), .Z(ereg_next[976]) );
  AND U42080 ( .A(mul_pow), .B(n39999), .Z(n39998) );
  XOR U42081 ( .A(ein[976]), .B(ein[975]), .Z(n39999) );
  XOR U42082 ( .A(ein[974]), .B(n40000), .Z(ereg_next[975]) );
  AND U42083 ( .A(mul_pow), .B(n40001), .Z(n40000) );
  XOR U42084 ( .A(ein[975]), .B(ein[974]), .Z(n40001) );
  XOR U42085 ( .A(ein[973]), .B(n40002), .Z(ereg_next[974]) );
  AND U42086 ( .A(mul_pow), .B(n40003), .Z(n40002) );
  XOR U42087 ( .A(ein[974]), .B(ein[973]), .Z(n40003) );
  XOR U42088 ( .A(ein[972]), .B(n40004), .Z(ereg_next[973]) );
  AND U42089 ( .A(mul_pow), .B(n40005), .Z(n40004) );
  XOR U42090 ( .A(ein[973]), .B(ein[972]), .Z(n40005) );
  XOR U42091 ( .A(ein[971]), .B(n40006), .Z(ereg_next[972]) );
  AND U42092 ( .A(mul_pow), .B(n40007), .Z(n40006) );
  XOR U42093 ( .A(ein[972]), .B(ein[971]), .Z(n40007) );
  XOR U42094 ( .A(ein[970]), .B(n40008), .Z(ereg_next[971]) );
  AND U42095 ( .A(mul_pow), .B(n40009), .Z(n40008) );
  XOR U42096 ( .A(ein[971]), .B(ein[970]), .Z(n40009) );
  XOR U42097 ( .A(ein[969]), .B(n40010), .Z(ereg_next[970]) );
  AND U42098 ( .A(mul_pow), .B(n40011), .Z(n40010) );
  XOR U42099 ( .A(ein[970]), .B(ein[969]), .Z(n40011) );
  XOR U42100 ( .A(ein[95]), .B(n40012), .Z(ereg_next[96]) );
  AND U42101 ( .A(mul_pow), .B(n40013), .Z(n40012) );
  XOR U42102 ( .A(ein[96]), .B(ein[95]), .Z(n40013) );
  XOR U42103 ( .A(ein[968]), .B(n40014), .Z(ereg_next[969]) );
  AND U42104 ( .A(mul_pow), .B(n40015), .Z(n40014) );
  XOR U42105 ( .A(ein[969]), .B(ein[968]), .Z(n40015) );
  XOR U42106 ( .A(ein[967]), .B(n40016), .Z(ereg_next[968]) );
  AND U42107 ( .A(mul_pow), .B(n40017), .Z(n40016) );
  XOR U42108 ( .A(ein[968]), .B(ein[967]), .Z(n40017) );
  XOR U42109 ( .A(ein[966]), .B(n40018), .Z(ereg_next[967]) );
  AND U42110 ( .A(mul_pow), .B(n40019), .Z(n40018) );
  XOR U42111 ( .A(ein[967]), .B(ein[966]), .Z(n40019) );
  XOR U42112 ( .A(ein[965]), .B(n40020), .Z(ereg_next[966]) );
  AND U42113 ( .A(mul_pow), .B(n40021), .Z(n40020) );
  XOR U42114 ( .A(ein[966]), .B(ein[965]), .Z(n40021) );
  XOR U42115 ( .A(ein[964]), .B(n40022), .Z(ereg_next[965]) );
  AND U42116 ( .A(mul_pow), .B(n40023), .Z(n40022) );
  XOR U42117 ( .A(ein[965]), .B(ein[964]), .Z(n40023) );
  XOR U42118 ( .A(ein[963]), .B(n40024), .Z(ereg_next[964]) );
  AND U42119 ( .A(mul_pow), .B(n40025), .Z(n40024) );
  XOR U42120 ( .A(ein[964]), .B(ein[963]), .Z(n40025) );
  XOR U42121 ( .A(ein[962]), .B(n40026), .Z(ereg_next[963]) );
  AND U42122 ( .A(mul_pow), .B(n40027), .Z(n40026) );
  XOR U42123 ( .A(ein[963]), .B(ein[962]), .Z(n40027) );
  XOR U42124 ( .A(ein[961]), .B(n40028), .Z(ereg_next[962]) );
  AND U42125 ( .A(mul_pow), .B(n40029), .Z(n40028) );
  XOR U42126 ( .A(ein[962]), .B(ein[961]), .Z(n40029) );
  XOR U42127 ( .A(ein[960]), .B(n40030), .Z(ereg_next[961]) );
  AND U42128 ( .A(mul_pow), .B(n40031), .Z(n40030) );
  XOR U42129 ( .A(ein[961]), .B(ein[960]), .Z(n40031) );
  XOR U42130 ( .A(ein[959]), .B(n40032), .Z(ereg_next[960]) );
  AND U42131 ( .A(mul_pow), .B(n40033), .Z(n40032) );
  XOR U42132 ( .A(ein[960]), .B(ein[959]), .Z(n40033) );
  XOR U42133 ( .A(ein[94]), .B(n40034), .Z(ereg_next[95]) );
  AND U42134 ( .A(mul_pow), .B(n40035), .Z(n40034) );
  XOR U42135 ( .A(ein[95]), .B(ein[94]), .Z(n40035) );
  XOR U42136 ( .A(ein[958]), .B(n40036), .Z(ereg_next[959]) );
  AND U42137 ( .A(mul_pow), .B(n40037), .Z(n40036) );
  XOR U42138 ( .A(ein[959]), .B(ein[958]), .Z(n40037) );
  XOR U42139 ( .A(ein[957]), .B(n40038), .Z(ereg_next[958]) );
  AND U42140 ( .A(mul_pow), .B(n40039), .Z(n40038) );
  XOR U42141 ( .A(ein[958]), .B(ein[957]), .Z(n40039) );
  XOR U42142 ( .A(ein[956]), .B(n40040), .Z(ereg_next[957]) );
  AND U42143 ( .A(mul_pow), .B(n40041), .Z(n40040) );
  XOR U42144 ( .A(ein[957]), .B(ein[956]), .Z(n40041) );
  XOR U42145 ( .A(ein[955]), .B(n40042), .Z(ereg_next[956]) );
  AND U42146 ( .A(mul_pow), .B(n40043), .Z(n40042) );
  XOR U42147 ( .A(ein[956]), .B(ein[955]), .Z(n40043) );
  XOR U42148 ( .A(ein[954]), .B(n40044), .Z(ereg_next[955]) );
  AND U42149 ( .A(mul_pow), .B(n40045), .Z(n40044) );
  XOR U42150 ( .A(ein[955]), .B(ein[954]), .Z(n40045) );
  XOR U42151 ( .A(ein[953]), .B(n40046), .Z(ereg_next[954]) );
  AND U42152 ( .A(mul_pow), .B(n40047), .Z(n40046) );
  XOR U42153 ( .A(ein[954]), .B(ein[953]), .Z(n40047) );
  XOR U42154 ( .A(ein[952]), .B(n40048), .Z(ereg_next[953]) );
  AND U42155 ( .A(mul_pow), .B(n40049), .Z(n40048) );
  XOR U42156 ( .A(ein[953]), .B(ein[952]), .Z(n40049) );
  XOR U42157 ( .A(ein[951]), .B(n40050), .Z(ereg_next[952]) );
  AND U42158 ( .A(mul_pow), .B(n40051), .Z(n40050) );
  XOR U42159 ( .A(ein[952]), .B(ein[951]), .Z(n40051) );
  XOR U42160 ( .A(ein[950]), .B(n40052), .Z(ereg_next[951]) );
  AND U42161 ( .A(mul_pow), .B(n40053), .Z(n40052) );
  XOR U42162 ( .A(ein[951]), .B(ein[950]), .Z(n40053) );
  XOR U42163 ( .A(ein[949]), .B(n40054), .Z(ereg_next[950]) );
  AND U42164 ( .A(mul_pow), .B(n40055), .Z(n40054) );
  XOR U42165 ( .A(ein[950]), .B(ein[949]), .Z(n40055) );
  XOR U42166 ( .A(ein[93]), .B(n40056), .Z(ereg_next[94]) );
  AND U42167 ( .A(mul_pow), .B(n40057), .Z(n40056) );
  XOR U42168 ( .A(ein[94]), .B(ein[93]), .Z(n40057) );
  XOR U42169 ( .A(ein[948]), .B(n40058), .Z(ereg_next[949]) );
  AND U42170 ( .A(mul_pow), .B(n40059), .Z(n40058) );
  XOR U42171 ( .A(ein[949]), .B(ein[948]), .Z(n40059) );
  XOR U42172 ( .A(ein[947]), .B(n40060), .Z(ereg_next[948]) );
  AND U42173 ( .A(mul_pow), .B(n40061), .Z(n40060) );
  XOR U42174 ( .A(ein[948]), .B(ein[947]), .Z(n40061) );
  XOR U42175 ( .A(ein[946]), .B(n40062), .Z(ereg_next[947]) );
  AND U42176 ( .A(mul_pow), .B(n40063), .Z(n40062) );
  XOR U42177 ( .A(ein[947]), .B(ein[946]), .Z(n40063) );
  XOR U42178 ( .A(ein[945]), .B(n40064), .Z(ereg_next[946]) );
  AND U42179 ( .A(mul_pow), .B(n40065), .Z(n40064) );
  XOR U42180 ( .A(ein[946]), .B(ein[945]), .Z(n40065) );
  XOR U42181 ( .A(ein[944]), .B(n40066), .Z(ereg_next[945]) );
  AND U42182 ( .A(mul_pow), .B(n40067), .Z(n40066) );
  XOR U42183 ( .A(ein[945]), .B(ein[944]), .Z(n40067) );
  XOR U42184 ( .A(ein[943]), .B(n40068), .Z(ereg_next[944]) );
  AND U42185 ( .A(mul_pow), .B(n40069), .Z(n40068) );
  XOR U42186 ( .A(ein[944]), .B(ein[943]), .Z(n40069) );
  XOR U42187 ( .A(ein[942]), .B(n40070), .Z(ereg_next[943]) );
  AND U42188 ( .A(mul_pow), .B(n40071), .Z(n40070) );
  XOR U42189 ( .A(ein[943]), .B(ein[942]), .Z(n40071) );
  XOR U42190 ( .A(ein[941]), .B(n40072), .Z(ereg_next[942]) );
  AND U42191 ( .A(mul_pow), .B(n40073), .Z(n40072) );
  XOR U42192 ( .A(ein[942]), .B(ein[941]), .Z(n40073) );
  XOR U42193 ( .A(ein[940]), .B(n40074), .Z(ereg_next[941]) );
  AND U42194 ( .A(mul_pow), .B(n40075), .Z(n40074) );
  XOR U42195 ( .A(ein[941]), .B(ein[940]), .Z(n40075) );
  XOR U42196 ( .A(ein[939]), .B(n40076), .Z(ereg_next[940]) );
  AND U42197 ( .A(mul_pow), .B(n40077), .Z(n40076) );
  XOR U42198 ( .A(ein[940]), .B(ein[939]), .Z(n40077) );
  XOR U42199 ( .A(ein[92]), .B(n40078), .Z(ereg_next[93]) );
  AND U42200 ( .A(mul_pow), .B(n40079), .Z(n40078) );
  XOR U42201 ( .A(ein[93]), .B(ein[92]), .Z(n40079) );
  XOR U42202 ( .A(ein[938]), .B(n40080), .Z(ereg_next[939]) );
  AND U42203 ( .A(mul_pow), .B(n40081), .Z(n40080) );
  XOR U42204 ( .A(ein[939]), .B(ein[938]), .Z(n40081) );
  XOR U42205 ( .A(ein[937]), .B(n40082), .Z(ereg_next[938]) );
  AND U42206 ( .A(mul_pow), .B(n40083), .Z(n40082) );
  XOR U42207 ( .A(ein[938]), .B(ein[937]), .Z(n40083) );
  XOR U42208 ( .A(ein[936]), .B(n40084), .Z(ereg_next[937]) );
  AND U42209 ( .A(mul_pow), .B(n40085), .Z(n40084) );
  XOR U42210 ( .A(ein[937]), .B(ein[936]), .Z(n40085) );
  XOR U42211 ( .A(ein[935]), .B(n40086), .Z(ereg_next[936]) );
  AND U42212 ( .A(mul_pow), .B(n40087), .Z(n40086) );
  XOR U42213 ( .A(ein[936]), .B(ein[935]), .Z(n40087) );
  XOR U42214 ( .A(ein[934]), .B(n40088), .Z(ereg_next[935]) );
  AND U42215 ( .A(mul_pow), .B(n40089), .Z(n40088) );
  XOR U42216 ( .A(ein[935]), .B(ein[934]), .Z(n40089) );
  XOR U42217 ( .A(ein[933]), .B(n40090), .Z(ereg_next[934]) );
  AND U42218 ( .A(mul_pow), .B(n40091), .Z(n40090) );
  XOR U42219 ( .A(ein[934]), .B(ein[933]), .Z(n40091) );
  XOR U42220 ( .A(ein[932]), .B(n40092), .Z(ereg_next[933]) );
  AND U42221 ( .A(mul_pow), .B(n40093), .Z(n40092) );
  XOR U42222 ( .A(ein[933]), .B(ein[932]), .Z(n40093) );
  XOR U42223 ( .A(ein[931]), .B(n40094), .Z(ereg_next[932]) );
  AND U42224 ( .A(mul_pow), .B(n40095), .Z(n40094) );
  XOR U42225 ( .A(ein[932]), .B(ein[931]), .Z(n40095) );
  XOR U42226 ( .A(ein[930]), .B(n40096), .Z(ereg_next[931]) );
  AND U42227 ( .A(mul_pow), .B(n40097), .Z(n40096) );
  XOR U42228 ( .A(ein[931]), .B(ein[930]), .Z(n40097) );
  XOR U42229 ( .A(ein[929]), .B(n40098), .Z(ereg_next[930]) );
  AND U42230 ( .A(mul_pow), .B(n40099), .Z(n40098) );
  XOR U42231 ( .A(ein[930]), .B(ein[929]), .Z(n40099) );
  XOR U42232 ( .A(ein[91]), .B(n40100), .Z(ereg_next[92]) );
  AND U42233 ( .A(mul_pow), .B(n40101), .Z(n40100) );
  XOR U42234 ( .A(ein[92]), .B(ein[91]), .Z(n40101) );
  XOR U42235 ( .A(ein[928]), .B(n40102), .Z(ereg_next[929]) );
  AND U42236 ( .A(mul_pow), .B(n40103), .Z(n40102) );
  XOR U42237 ( .A(ein[929]), .B(ein[928]), .Z(n40103) );
  XOR U42238 ( .A(ein[927]), .B(n40104), .Z(ereg_next[928]) );
  AND U42239 ( .A(mul_pow), .B(n40105), .Z(n40104) );
  XOR U42240 ( .A(ein[928]), .B(ein[927]), .Z(n40105) );
  XOR U42241 ( .A(ein[926]), .B(n40106), .Z(ereg_next[927]) );
  AND U42242 ( .A(mul_pow), .B(n40107), .Z(n40106) );
  XOR U42243 ( .A(ein[927]), .B(ein[926]), .Z(n40107) );
  XOR U42244 ( .A(ein[925]), .B(n40108), .Z(ereg_next[926]) );
  AND U42245 ( .A(mul_pow), .B(n40109), .Z(n40108) );
  XOR U42246 ( .A(ein[926]), .B(ein[925]), .Z(n40109) );
  XOR U42247 ( .A(ein[924]), .B(n40110), .Z(ereg_next[925]) );
  AND U42248 ( .A(mul_pow), .B(n40111), .Z(n40110) );
  XOR U42249 ( .A(ein[925]), .B(ein[924]), .Z(n40111) );
  XOR U42250 ( .A(ein[923]), .B(n40112), .Z(ereg_next[924]) );
  AND U42251 ( .A(mul_pow), .B(n40113), .Z(n40112) );
  XOR U42252 ( .A(ein[924]), .B(ein[923]), .Z(n40113) );
  XOR U42253 ( .A(ein[922]), .B(n40114), .Z(ereg_next[923]) );
  AND U42254 ( .A(mul_pow), .B(n40115), .Z(n40114) );
  XOR U42255 ( .A(ein[923]), .B(ein[922]), .Z(n40115) );
  XOR U42256 ( .A(ein[921]), .B(n40116), .Z(ereg_next[922]) );
  AND U42257 ( .A(mul_pow), .B(n40117), .Z(n40116) );
  XOR U42258 ( .A(ein[922]), .B(ein[921]), .Z(n40117) );
  XOR U42259 ( .A(ein[920]), .B(n40118), .Z(ereg_next[921]) );
  AND U42260 ( .A(mul_pow), .B(n40119), .Z(n40118) );
  XOR U42261 ( .A(ein[921]), .B(ein[920]), .Z(n40119) );
  XOR U42262 ( .A(ein[919]), .B(n40120), .Z(ereg_next[920]) );
  AND U42263 ( .A(mul_pow), .B(n40121), .Z(n40120) );
  XOR U42264 ( .A(ein[920]), .B(ein[919]), .Z(n40121) );
  XOR U42265 ( .A(ein[90]), .B(n40122), .Z(ereg_next[91]) );
  AND U42266 ( .A(mul_pow), .B(n40123), .Z(n40122) );
  XOR U42267 ( .A(ein[91]), .B(ein[90]), .Z(n40123) );
  XOR U42268 ( .A(ein[918]), .B(n40124), .Z(ereg_next[919]) );
  AND U42269 ( .A(mul_pow), .B(n40125), .Z(n40124) );
  XOR U42270 ( .A(ein[919]), .B(ein[918]), .Z(n40125) );
  XOR U42271 ( .A(ein[917]), .B(n40126), .Z(ereg_next[918]) );
  AND U42272 ( .A(mul_pow), .B(n40127), .Z(n40126) );
  XOR U42273 ( .A(ein[918]), .B(ein[917]), .Z(n40127) );
  XOR U42274 ( .A(ein[916]), .B(n40128), .Z(ereg_next[917]) );
  AND U42275 ( .A(mul_pow), .B(n40129), .Z(n40128) );
  XOR U42276 ( .A(ein[917]), .B(ein[916]), .Z(n40129) );
  XOR U42277 ( .A(ein[915]), .B(n40130), .Z(ereg_next[916]) );
  AND U42278 ( .A(mul_pow), .B(n40131), .Z(n40130) );
  XOR U42279 ( .A(ein[916]), .B(ein[915]), .Z(n40131) );
  XOR U42280 ( .A(ein[914]), .B(n40132), .Z(ereg_next[915]) );
  AND U42281 ( .A(mul_pow), .B(n40133), .Z(n40132) );
  XOR U42282 ( .A(ein[915]), .B(ein[914]), .Z(n40133) );
  XOR U42283 ( .A(ein[913]), .B(n40134), .Z(ereg_next[914]) );
  AND U42284 ( .A(mul_pow), .B(n40135), .Z(n40134) );
  XOR U42285 ( .A(ein[914]), .B(ein[913]), .Z(n40135) );
  XOR U42286 ( .A(ein[912]), .B(n40136), .Z(ereg_next[913]) );
  AND U42287 ( .A(mul_pow), .B(n40137), .Z(n40136) );
  XOR U42288 ( .A(ein[913]), .B(ein[912]), .Z(n40137) );
  XOR U42289 ( .A(ein[911]), .B(n40138), .Z(ereg_next[912]) );
  AND U42290 ( .A(mul_pow), .B(n40139), .Z(n40138) );
  XOR U42291 ( .A(ein[912]), .B(ein[911]), .Z(n40139) );
  XOR U42292 ( .A(ein[910]), .B(n40140), .Z(ereg_next[911]) );
  AND U42293 ( .A(mul_pow), .B(n40141), .Z(n40140) );
  XOR U42294 ( .A(ein[911]), .B(ein[910]), .Z(n40141) );
  XOR U42295 ( .A(ein[909]), .B(n40142), .Z(ereg_next[910]) );
  AND U42296 ( .A(mul_pow), .B(n40143), .Z(n40142) );
  XOR U42297 ( .A(ein[910]), .B(ein[909]), .Z(n40143) );
  XOR U42298 ( .A(ein[89]), .B(n40144), .Z(ereg_next[90]) );
  AND U42299 ( .A(mul_pow), .B(n40145), .Z(n40144) );
  XOR U42300 ( .A(ein[90]), .B(ein[89]), .Z(n40145) );
  XOR U42301 ( .A(ein[908]), .B(n40146), .Z(ereg_next[909]) );
  AND U42302 ( .A(mul_pow), .B(n40147), .Z(n40146) );
  XOR U42303 ( .A(ein[909]), .B(ein[908]), .Z(n40147) );
  XOR U42304 ( .A(ein[907]), .B(n40148), .Z(ereg_next[908]) );
  AND U42305 ( .A(mul_pow), .B(n40149), .Z(n40148) );
  XOR U42306 ( .A(ein[908]), .B(ein[907]), .Z(n40149) );
  XOR U42307 ( .A(ein[906]), .B(n40150), .Z(ereg_next[907]) );
  AND U42308 ( .A(mul_pow), .B(n40151), .Z(n40150) );
  XOR U42309 ( .A(ein[907]), .B(ein[906]), .Z(n40151) );
  XOR U42310 ( .A(ein[905]), .B(n40152), .Z(ereg_next[906]) );
  AND U42311 ( .A(mul_pow), .B(n40153), .Z(n40152) );
  XOR U42312 ( .A(ein[906]), .B(ein[905]), .Z(n40153) );
  XOR U42313 ( .A(ein[904]), .B(n40154), .Z(ereg_next[905]) );
  AND U42314 ( .A(mul_pow), .B(n40155), .Z(n40154) );
  XOR U42315 ( .A(ein[905]), .B(ein[904]), .Z(n40155) );
  XOR U42316 ( .A(ein[903]), .B(n40156), .Z(ereg_next[904]) );
  AND U42317 ( .A(mul_pow), .B(n40157), .Z(n40156) );
  XOR U42318 ( .A(ein[904]), .B(ein[903]), .Z(n40157) );
  XOR U42319 ( .A(ein[902]), .B(n40158), .Z(ereg_next[903]) );
  AND U42320 ( .A(mul_pow), .B(n40159), .Z(n40158) );
  XOR U42321 ( .A(ein[903]), .B(ein[902]), .Z(n40159) );
  XOR U42322 ( .A(ein[901]), .B(n40160), .Z(ereg_next[902]) );
  AND U42323 ( .A(mul_pow), .B(n40161), .Z(n40160) );
  XOR U42324 ( .A(ein[902]), .B(ein[901]), .Z(n40161) );
  XOR U42325 ( .A(ein[900]), .B(n40162), .Z(ereg_next[901]) );
  AND U42326 ( .A(mul_pow), .B(n40163), .Z(n40162) );
  XOR U42327 ( .A(ein[901]), .B(ein[900]), .Z(n40163) );
  XOR U42328 ( .A(ein[899]), .B(n40164), .Z(ereg_next[900]) );
  AND U42329 ( .A(mul_pow), .B(n40165), .Z(n40164) );
  XOR U42330 ( .A(ein[900]), .B(ein[899]), .Z(n40165) );
  XOR U42331 ( .A(ein[7]), .B(n40166), .Z(ereg_next[8]) );
  AND U42332 ( .A(mul_pow), .B(n40167), .Z(n40166) );
  XOR U42333 ( .A(ein[8]), .B(ein[7]), .Z(n40167) );
  XOR U42334 ( .A(ein[88]), .B(n40168), .Z(ereg_next[89]) );
  AND U42335 ( .A(mul_pow), .B(n40169), .Z(n40168) );
  XOR U42336 ( .A(ein[89]), .B(ein[88]), .Z(n40169) );
  XOR U42337 ( .A(ein[898]), .B(n40170), .Z(ereg_next[899]) );
  AND U42338 ( .A(mul_pow), .B(n40171), .Z(n40170) );
  XOR U42339 ( .A(ein[899]), .B(ein[898]), .Z(n40171) );
  XOR U42340 ( .A(ein[897]), .B(n40172), .Z(ereg_next[898]) );
  AND U42341 ( .A(mul_pow), .B(n40173), .Z(n40172) );
  XOR U42342 ( .A(ein[898]), .B(ein[897]), .Z(n40173) );
  XOR U42343 ( .A(ein[896]), .B(n40174), .Z(ereg_next[897]) );
  AND U42344 ( .A(mul_pow), .B(n40175), .Z(n40174) );
  XOR U42345 ( .A(ein[897]), .B(ein[896]), .Z(n40175) );
  XOR U42346 ( .A(ein[895]), .B(n40176), .Z(ereg_next[896]) );
  AND U42347 ( .A(mul_pow), .B(n40177), .Z(n40176) );
  XOR U42348 ( .A(ein[896]), .B(ein[895]), .Z(n40177) );
  XOR U42349 ( .A(ein[894]), .B(n40178), .Z(ereg_next[895]) );
  AND U42350 ( .A(mul_pow), .B(n40179), .Z(n40178) );
  XOR U42351 ( .A(ein[895]), .B(ein[894]), .Z(n40179) );
  XOR U42352 ( .A(ein[893]), .B(n40180), .Z(ereg_next[894]) );
  AND U42353 ( .A(mul_pow), .B(n40181), .Z(n40180) );
  XOR U42354 ( .A(ein[894]), .B(ein[893]), .Z(n40181) );
  XOR U42355 ( .A(ein[892]), .B(n40182), .Z(ereg_next[893]) );
  AND U42356 ( .A(mul_pow), .B(n40183), .Z(n40182) );
  XOR U42357 ( .A(ein[893]), .B(ein[892]), .Z(n40183) );
  XOR U42358 ( .A(ein[891]), .B(n40184), .Z(ereg_next[892]) );
  AND U42359 ( .A(mul_pow), .B(n40185), .Z(n40184) );
  XOR U42360 ( .A(ein[892]), .B(ein[891]), .Z(n40185) );
  XOR U42361 ( .A(ein[890]), .B(n40186), .Z(ereg_next[891]) );
  AND U42362 ( .A(mul_pow), .B(n40187), .Z(n40186) );
  XOR U42363 ( .A(ein[891]), .B(ein[890]), .Z(n40187) );
  XOR U42364 ( .A(ein[889]), .B(n40188), .Z(ereg_next[890]) );
  AND U42365 ( .A(mul_pow), .B(n40189), .Z(n40188) );
  XOR U42366 ( .A(ein[890]), .B(ein[889]), .Z(n40189) );
  XOR U42367 ( .A(ein[87]), .B(n40190), .Z(ereg_next[88]) );
  AND U42368 ( .A(mul_pow), .B(n40191), .Z(n40190) );
  XOR U42369 ( .A(ein[88]), .B(ein[87]), .Z(n40191) );
  XOR U42370 ( .A(ein[888]), .B(n40192), .Z(ereg_next[889]) );
  AND U42371 ( .A(mul_pow), .B(n40193), .Z(n40192) );
  XOR U42372 ( .A(ein[889]), .B(ein[888]), .Z(n40193) );
  XOR U42373 ( .A(ein[887]), .B(n40194), .Z(ereg_next[888]) );
  AND U42374 ( .A(mul_pow), .B(n40195), .Z(n40194) );
  XOR U42375 ( .A(ein[888]), .B(ein[887]), .Z(n40195) );
  XOR U42376 ( .A(ein[886]), .B(n40196), .Z(ereg_next[887]) );
  AND U42377 ( .A(mul_pow), .B(n40197), .Z(n40196) );
  XOR U42378 ( .A(ein[887]), .B(ein[886]), .Z(n40197) );
  XOR U42379 ( .A(ein[885]), .B(n40198), .Z(ereg_next[886]) );
  AND U42380 ( .A(mul_pow), .B(n40199), .Z(n40198) );
  XOR U42381 ( .A(ein[886]), .B(ein[885]), .Z(n40199) );
  XOR U42382 ( .A(ein[884]), .B(n40200), .Z(ereg_next[885]) );
  AND U42383 ( .A(mul_pow), .B(n40201), .Z(n40200) );
  XOR U42384 ( .A(ein[885]), .B(ein[884]), .Z(n40201) );
  XOR U42385 ( .A(ein[883]), .B(n40202), .Z(ereg_next[884]) );
  AND U42386 ( .A(mul_pow), .B(n40203), .Z(n40202) );
  XOR U42387 ( .A(ein[884]), .B(ein[883]), .Z(n40203) );
  XOR U42388 ( .A(ein[882]), .B(n40204), .Z(ereg_next[883]) );
  AND U42389 ( .A(mul_pow), .B(n40205), .Z(n40204) );
  XOR U42390 ( .A(ein[883]), .B(ein[882]), .Z(n40205) );
  XOR U42391 ( .A(ein[881]), .B(n40206), .Z(ereg_next[882]) );
  AND U42392 ( .A(mul_pow), .B(n40207), .Z(n40206) );
  XOR U42393 ( .A(ein[882]), .B(ein[881]), .Z(n40207) );
  XOR U42394 ( .A(ein[880]), .B(n40208), .Z(ereg_next[881]) );
  AND U42395 ( .A(mul_pow), .B(n40209), .Z(n40208) );
  XOR U42396 ( .A(ein[881]), .B(ein[880]), .Z(n40209) );
  XOR U42397 ( .A(ein[879]), .B(n40210), .Z(ereg_next[880]) );
  AND U42398 ( .A(mul_pow), .B(n40211), .Z(n40210) );
  XOR U42399 ( .A(ein[880]), .B(ein[879]), .Z(n40211) );
  XOR U42400 ( .A(ein[86]), .B(n40212), .Z(ereg_next[87]) );
  AND U42401 ( .A(mul_pow), .B(n40213), .Z(n40212) );
  XOR U42402 ( .A(ein[87]), .B(ein[86]), .Z(n40213) );
  XOR U42403 ( .A(ein[878]), .B(n40214), .Z(ereg_next[879]) );
  AND U42404 ( .A(mul_pow), .B(n40215), .Z(n40214) );
  XOR U42405 ( .A(ein[879]), .B(ein[878]), .Z(n40215) );
  XOR U42406 ( .A(ein[877]), .B(n40216), .Z(ereg_next[878]) );
  AND U42407 ( .A(mul_pow), .B(n40217), .Z(n40216) );
  XOR U42408 ( .A(ein[878]), .B(ein[877]), .Z(n40217) );
  XOR U42409 ( .A(ein[876]), .B(n40218), .Z(ereg_next[877]) );
  AND U42410 ( .A(mul_pow), .B(n40219), .Z(n40218) );
  XOR U42411 ( .A(ein[877]), .B(ein[876]), .Z(n40219) );
  XOR U42412 ( .A(ein[875]), .B(n40220), .Z(ereg_next[876]) );
  AND U42413 ( .A(mul_pow), .B(n40221), .Z(n40220) );
  XOR U42414 ( .A(ein[876]), .B(ein[875]), .Z(n40221) );
  XOR U42415 ( .A(ein[874]), .B(n40222), .Z(ereg_next[875]) );
  AND U42416 ( .A(mul_pow), .B(n40223), .Z(n40222) );
  XOR U42417 ( .A(ein[875]), .B(ein[874]), .Z(n40223) );
  XOR U42418 ( .A(ein[873]), .B(n40224), .Z(ereg_next[874]) );
  AND U42419 ( .A(mul_pow), .B(n40225), .Z(n40224) );
  XOR U42420 ( .A(ein[874]), .B(ein[873]), .Z(n40225) );
  XOR U42421 ( .A(ein[872]), .B(n40226), .Z(ereg_next[873]) );
  AND U42422 ( .A(mul_pow), .B(n40227), .Z(n40226) );
  XOR U42423 ( .A(ein[873]), .B(ein[872]), .Z(n40227) );
  XOR U42424 ( .A(ein[871]), .B(n40228), .Z(ereg_next[872]) );
  AND U42425 ( .A(mul_pow), .B(n40229), .Z(n40228) );
  XOR U42426 ( .A(ein[872]), .B(ein[871]), .Z(n40229) );
  XOR U42427 ( .A(ein[870]), .B(n40230), .Z(ereg_next[871]) );
  AND U42428 ( .A(mul_pow), .B(n40231), .Z(n40230) );
  XOR U42429 ( .A(ein[871]), .B(ein[870]), .Z(n40231) );
  XOR U42430 ( .A(ein[869]), .B(n40232), .Z(ereg_next[870]) );
  AND U42431 ( .A(mul_pow), .B(n40233), .Z(n40232) );
  XOR U42432 ( .A(ein[870]), .B(ein[869]), .Z(n40233) );
  XOR U42433 ( .A(ein[85]), .B(n40234), .Z(ereg_next[86]) );
  AND U42434 ( .A(mul_pow), .B(n40235), .Z(n40234) );
  XOR U42435 ( .A(ein[86]), .B(ein[85]), .Z(n40235) );
  XOR U42436 ( .A(ein[868]), .B(n40236), .Z(ereg_next[869]) );
  AND U42437 ( .A(mul_pow), .B(n40237), .Z(n40236) );
  XOR U42438 ( .A(ein[869]), .B(ein[868]), .Z(n40237) );
  XOR U42439 ( .A(ein[867]), .B(n40238), .Z(ereg_next[868]) );
  AND U42440 ( .A(mul_pow), .B(n40239), .Z(n40238) );
  XOR U42441 ( .A(ein[868]), .B(ein[867]), .Z(n40239) );
  XOR U42442 ( .A(ein[866]), .B(n40240), .Z(ereg_next[867]) );
  AND U42443 ( .A(mul_pow), .B(n40241), .Z(n40240) );
  XOR U42444 ( .A(ein[867]), .B(ein[866]), .Z(n40241) );
  XOR U42445 ( .A(ein[865]), .B(n40242), .Z(ereg_next[866]) );
  AND U42446 ( .A(mul_pow), .B(n40243), .Z(n40242) );
  XOR U42447 ( .A(ein[866]), .B(ein[865]), .Z(n40243) );
  XOR U42448 ( .A(ein[864]), .B(n40244), .Z(ereg_next[865]) );
  AND U42449 ( .A(mul_pow), .B(n40245), .Z(n40244) );
  XOR U42450 ( .A(ein[865]), .B(ein[864]), .Z(n40245) );
  XOR U42451 ( .A(ein[863]), .B(n40246), .Z(ereg_next[864]) );
  AND U42452 ( .A(mul_pow), .B(n40247), .Z(n40246) );
  XOR U42453 ( .A(ein[864]), .B(ein[863]), .Z(n40247) );
  XOR U42454 ( .A(ein[862]), .B(n40248), .Z(ereg_next[863]) );
  AND U42455 ( .A(mul_pow), .B(n40249), .Z(n40248) );
  XOR U42456 ( .A(ein[863]), .B(ein[862]), .Z(n40249) );
  XOR U42457 ( .A(ein[861]), .B(n40250), .Z(ereg_next[862]) );
  AND U42458 ( .A(mul_pow), .B(n40251), .Z(n40250) );
  XOR U42459 ( .A(ein[862]), .B(ein[861]), .Z(n40251) );
  XOR U42460 ( .A(ein[860]), .B(n40252), .Z(ereg_next[861]) );
  AND U42461 ( .A(mul_pow), .B(n40253), .Z(n40252) );
  XOR U42462 ( .A(ein[861]), .B(ein[860]), .Z(n40253) );
  XOR U42463 ( .A(ein[859]), .B(n40254), .Z(ereg_next[860]) );
  AND U42464 ( .A(mul_pow), .B(n40255), .Z(n40254) );
  XOR U42465 ( .A(ein[860]), .B(ein[859]), .Z(n40255) );
  XOR U42466 ( .A(ein[84]), .B(n40256), .Z(ereg_next[85]) );
  AND U42467 ( .A(mul_pow), .B(n40257), .Z(n40256) );
  XOR U42468 ( .A(ein[85]), .B(ein[84]), .Z(n40257) );
  XOR U42469 ( .A(ein[858]), .B(n40258), .Z(ereg_next[859]) );
  AND U42470 ( .A(mul_pow), .B(n40259), .Z(n40258) );
  XOR U42471 ( .A(ein[859]), .B(ein[858]), .Z(n40259) );
  XOR U42472 ( .A(ein[857]), .B(n40260), .Z(ereg_next[858]) );
  AND U42473 ( .A(mul_pow), .B(n40261), .Z(n40260) );
  XOR U42474 ( .A(ein[858]), .B(ein[857]), .Z(n40261) );
  XOR U42475 ( .A(ein[856]), .B(n40262), .Z(ereg_next[857]) );
  AND U42476 ( .A(mul_pow), .B(n40263), .Z(n40262) );
  XOR U42477 ( .A(ein[857]), .B(ein[856]), .Z(n40263) );
  XOR U42478 ( .A(ein[855]), .B(n40264), .Z(ereg_next[856]) );
  AND U42479 ( .A(mul_pow), .B(n40265), .Z(n40264) );
  XOR U42480 ( .A(ein[856]), .B(ein[855]), .Z(n40265) );
  XOR U42481 ( .A(ein[854]), .B(n40266), .Z(ereg_next[855]) );
  AND U42482 ( .A(mul_pow), .B(n40267), .Z(n40266) );
  XOR U42483 ( .A(ein[855]), .B(ein[854]), .Z(n40267) );
  XOR U42484 ( .A(ein[853]), .B(n40268), .Z(ereg_next[854]) );
  AND U42485 ( .A(mul_pow), .B(n40269), .Z(n40268) );
  XOR U42486 ( .A(ein[854]), .B(ein[853]), .Z(n40269) );
  XOR U42487 ( .A(ein[852]), .B(n40270), .Z(ereg_next[853]) );
  AND U42488 ( .A(mul_pow), .B(n40271), .Z(n40270) );
  XOR U42489 ( .A(ein[853]), .B(ein[852]), .Z(n40271) );
  XOR U42490 ( .A(ein[851]), .B(n40272), .Z(ereg_next[852]) );
  AND U42491 ( .A(mul_pow), .B(n40273), .Z(n40272) );
  XOR U42492 ( .A(ein[852]), .B(ein[851]), .Z(n40273) );
  XOR U42493 ( .A(ein[850]), .B(n40274), .Z(ereg_next[851]) );
  AND U42494 ( .A(mul_pow), .B(n40275), .Z(n40274) );
  XOR U42495 ( .A(ein[851]), .B(ein[850]), .Z(n40275) );
  XOR U42496 ( .A(ein[849]), .B(n40276), .Z(ereg_next[850]) );
  AND U42497 ( .A(mul_pow), .B(n40277), .Z(n40276) );
  XOR U42498 ( .A(ein[850]), .B(ein[849]), .Z(n40277) );
  XOR U42499 ( .A(ein[83]), .B(n40278), .Z(ereg_next[84]) );
  AND U42500 ( .A(mul_pow), .B(n40279), .Z(n40278) );
  XOR U42501 ( .A(ein[84]), .B(ein[83]), .Z(n40279) );
  XOR U42502 ( .A(ein[848]), .B(n40280), .Z(ereg_next[849]) );
  AND U42503 ( .A(mul_pow), .B(n40281), .Z(n40280) );
  XOR U42504 ( .A(ein[849]), .B(ein[848]), .Z(n40281) );
  XOR U42505 ( .A(ein[847]), .B(n40282), .Z(ereg_next[848]) );
  AND U42506 ( .A(mul_pow), .B(n40283), .Z(n40282) );
  XOR U42507 ( .A(ein[848]), .B(ein[847]), .Z(n40283) );
  XOR U42508 ( .A(ein[846]), .B(n40284), .Z(ereg_next[847]) );
  AND U42509 ( .A(mul_pow), .B(n40285), .Z(n40284) );
  XOR U42510 ( .A(ein[847]), .B(ein[846]), .Z(n40285) );
  XOR U42511 ( .A(ein[845]), .B(n40286), .Z(ereg_next[846]) );
  AND U42512 ( .A(mul_pow), .B(n40287), .Z(n40286) );
  XOR U42513 ( .A(ein[846]), .B(ein[845]), .Z(n40287) );
  XOR U42514 ( .A(ein[844]), .B(n40288), .Z(ereg_next[845]) );
  AND U42515 ( .A(mul_pow), .B(n40289), .Z(n40288) );
  XOR U42516 ( .A(ein[845]), .B(ein[844]), .Z(n40289) );
  XOR U42517 ( .A(ein[843]), .B(n40290), .Z(ereg_next[844]) );
  AND U42518 ( .A(mul_pow), .B(n40291), .Z(n40290) );
  XOR U42519 ( .A(ein[844]), .B(ein[843]), .Z(n40291) );
  XOR U42520 ( .A(ein[842]), .B(n40292), .Z(ereg_next[843]) );
  AND U42521 ( .A(mul_pow), .B(n40293), .Z(n40292) );
  XOR U42522 ( .A(ein[843]), .B(ein[842]), .Z(n40293) );
  XOR U42523 ( .A(ein[841]), .B(n40294), .Z(ereg_next[842]) );
  AND U42524 ( .A(mul_pow), .B(n40295), .Z(n40294) );
  XOR U42525 ( .A(ein[842]), .B(ein[841]), .Z(n40295) );
  XOR U42526 ( .A(ein[840]), .B(n40296), .Z(ereg_next[841]) );
  AND U42527 ( .A(mul_pow), .B(n40297), .Z(n40296) );
  XOR U42528 ( .A(ein[841]), .B(ein[840]), .Z(n40297) );
  XOR U42529 ( .A(ein[839]), .B(n40298), .Z(ereg_next[840]) );
  AND U42530 ( .A(mul_pow), .B(n40299), .Z(n40298) );
  XOR U42531 ( .A(ein[840]), .B(ein[839]), .Z(n40299) );
  XOR U42532 ( .A(ein[82]), .B(n40300), .Z(ereg_next[83]) );
  AND U42533 ( .A(mul_pow), .B(n40301), .Z(n40300) );
  XOR U42534 ( .A(ein[83]), .B(ein[82]), .Z(n40301) );
  XOR U42535 ( .A(ein[838]), .B(n40302), .Z(ereg_next[839]) );
  AND U42536 ( .A(mul_pow), .B(n40303), .Z(n40302) );
  XOR U42537 ( .A(ein[839]), .B(ein[838]), .Z(n40303) );
  XOR U42538 ( .A(ein[837]), .B(n40304), .Z(ereg_next[838]) );
  AND U42539 ( .A(mul_pow), .B(n40305), .Z(n40304) );
  XOR U42540 ( .A(ein[838]), .B(ein[837]), .Z(n40305) );
  XOR U42541 ( .A(ein[836]), .B(n40306), .Z(ereg_next[837]) );
  AND U42542 ( .A(mul_pow), .B(n40307), .Z(n40306) );
  XOR U42543 ( .A(ein[837]), .B(ein[836]), .Z(n40307) );
  XOR U42544 ( .A(ein[835]), .B(n40308), .Z(ereg_next[836]) );
  AND U42545 ( .A(mul_pow), .B(n40309), .Z(n40308) );
  XOR U42546 ( .A(ein[836]), .B(ein[835]), .Z(n40309) );
  XOR U42547 ( .A(ein[834]), .B(n40310), .Z(ereg_next[835]) );
  AND U42548 ( .A(mul_pow), .B(n40311), .Z(n40310) );
  XOR U42549 ( .A(ein[835]), .B(ein[834]), .Z(n40311) );
  XOR U42550 ( .A(ein[833]), .B(n40312), .Z(ereg_next[834]) );
  AND U42551 ( .A(mul_pow), .B(n40313), .Z(n40312) );
  XOR U42552 ( .A(ein[834]), .B(ein[833]), .Z(n40313) );
  XOR U42553 ( .A(ein[832]), .B(n40314), .Z(ereg_next[833]) );
  AND U42554 ( .A(mul_pow), .B(n40315), .Z(n40314) );
  XOR U42555 ( .A(ein[833]), .B(ein[832]), .Z(n40315) );
  XOR U42556 ( .A(ein[831]), .B(n40316), .Z(ereg_next[832]) );
  AND U42557 ( .A(mul_pow), .B(n40317), .Z(n40316) );
  XOR U42558 ( .A(ein[832]), .B(ein[831]), .Z(n40317) );
  XOR U42559 ( .A(ein[830]), .B(n40318), .Z(ereg_next[831]) );
  AND U42560 ( .A(mul_pow), .B(n40319), .Z(n40318) );
  XOR U42561 ( .A(ein[831]), .B(ein[830]), .Z(n40319) );
  XOR U42562 ( .A(ein[829]), .B(n40320), .Z(ereg_next[830]) );
  AND U42563 ( .A(mul_pow), .B(n40321), .Z(n40320) );
  XOR U42564 ( .A(ein[830]), .B(ein[829]), .Z(n40321) );
  XOR U42565 ( .A(ein[81]), .B(n40322), .Z(ereg_next[82]) );
  AND U42566 ( .A(mul_pow), .B(n40323), .Z(n40322) );
  XOR U42567 ( .A(ein[82]), .B(ein[81]), .Z(n40323) );
  XOR U42568 ( .A(ein[828]), .B(n40324), .Z(ereg_next[829]) );
  AND U42569 ( .A(mul_pow), .B(n40325), .Z(n40324) );
  XOR U42570 ( .A(ein[829]), .B(ein[828]), .Z(n40325) );
  XOR U42571 ( .A(ein[827]), .B(n40326), .Z(ereg_next[828]) );
  AND U42572 ( .A(mul_pow), .B(n40327), .Z(n40326) );
  XOR U42573 ( .A(ein[828]), .B(ein[827]), .Z(n40327) );
  XOR U42574 ( .A(ein[826]), .B(n40328), .Z(ereg_next[827]) );
  AND U42575 ( .A(mul_pow), .B(n40329), .Z(n40328) );
  XOR U42576 ( .A(ein[827]), .B(ein[826]), .Z(n40329) );
  XOR U42577 ( .A(ein[825]), .B(n40330), .Z(ereg_next[826]) );
  AND U42578 ( .A(mul_pow), .B(n40331), .Z(n40330) );
  XOR U42579 ( .A(ein[826]), .B(ein[825]), .Z(n40331) );
  XOR U42580 ( .A(ein[824]), .B(n40332), .Z(ereg_next[825]) );
  AND U42581 ( .A(mul_pow), .B(n40333), .Z(n40332) );
  XOR U42582 ( .A(ein[825]), .B(ein[824]), .Z(n40333) );
  XOR U42583 ( .A(ein[823]), .B(n40334), .Z(ereg_next[824]) );
  AND U42584 ( .A(mul_pow), .B(n40335), .Z(n40334) );
  XOR U42585 ( .A(ein[824]), .B(ein[823]), .Z(n40335) );
  XOR U42586 ( .A(ein[822]), .B(n40336), .Z(ereg_next[823]) );
  AND U42587 ( .A(mul_pow), .B(n40337), .Z(n40336) );
  XOR U42588 ( .A(ein[823]), .B(ein[822]), .Z(n40337) );
  XOR U42589 ( .A(ein[821]), .B(n40338), .Z(ereg_next[822]) );
  AND U42590 ( .A(mul_pow), .B(n40339), .Z(n40338) );
  XOR U42591 ( .A(ein[822]), .B(ein[821]), .Z(n40339) );
  XOR U42592 ( .A(ein[820]), .B(n40340), .Z(ereg_next[821]) );
  AND U42593 ( .A(mul_pow), .B(n40341), .Z(n40340) );
  XOR U42594 ( .A(ein[821]), .B(ein[820]), .Z(n40341) );
  XOR U42595 ( .A(ein[819]), .B(n40342), .Z(ereg_next[820]) );
  AND U42596 ( .A(mul_pow), .B(n40343), .Z(n40342) );
  XOR U42597 ( .A(ein[820]), .B(ein[819]), .Z(n40343) );
  XOR U42598 ( .A(ein[80]), .B(n40344), .Z(ereg_next[81]) );
  AND U42599 ( .A(mul_pow), .B(n40345), .Z(n40344) );
  XOR U42600 ( .A(ein[81]), .B(ein[80]), .Z(n40345) );
  XOR U42601 ( .A(ein[818]), .B(n40346), .Z(ereg_next[819]) );
  AND U42602 ( .A(mul_pow), .B(n40347), .Z(n40346) );
  XOR U42603 ( .A(ein[819]), .B(ein[818]), .Z(n40347) );
  XOR U42604 ( .A(ein[817]), .B(n40348), .Z(ereg_next[818]) );
  AND U42605 ( .A(mul_pow), .B(n40349), .Z(n40348) );
  XOR U42606 ( .A(ein[818]), .B(ein[817]), .Z(n40349) );
  XOR U42607 ( .A(ein[816]), .B(n40350), .Z(ereg_next[817]) );
  AND U42608 ( .A(mul_pow), .B(n40351), .Z(n40350) );
  XOR U42609 ( .A(ein[817]), .B(ein[816]), .Z(n40351) );
  XOR U42610 ( .A(ein[815]), .B(n40352), .Z(ereg_next[816]) );
  AND U42611 ( .A(mul_pow), .B(n40353), .Z(n40352) );
  XOR U42612 ( .A(ein[816]), .B(ein[815]), .Z(n40353) );
  XOR U42613 ( .A(ein[814]), .B(n40354), .Z(ereg_next[815]) );
  AND U42614 ( .A(mul_pow), .B(n40355), .Z(n40354) );
  XOR U42615 ( .A(ein[815]), .B(ein[814]), .Z(n40355) );
  XOR U42616 ( .A(ein[813]), .B(n40356), .Z(ereg_next[814]) );
  AND U42617 ( .A(mul_pow), .B(n40357), .Z(n40356) );
  XOR U42618 ( .A(ein[814]), .B(ein[813]), .Z(n40357) );
  XOR U42619 ( .A(ein[812]), .B(n40358), .Z(ereg_next[813]) );
  AND U42620 ( .A(mul_pow), .B(n40359), .Z(n40358) );
  XOR U42621 ( .A(ein[813]), .B(ein[812]), .Z(n40359) );
  XOR U42622 ( .A(ein[811]), .B(n40360), .Z(ereg_next[812]) );
  AND U42623 ( .A(mul_pow), .B(n40361), .Z(n40360) );
  XOR U42624 ( .A(ein[812]), .B(ein[811]), .Z(n40361) );
  XOR U42625 ( .A(ein[810]), .B(n40362), .Z(ereg_next[811]) );
  AND U42626 ( .A(mul_pow), .B(n40363), .Z(n40362) );
  XOR U42627 ( .A(ein[811]), .B(ein[810]), .Z(n40363) );
  XOR U42628 ( .A(ein[809]), .B(n40364), .Z(ereg_next[810]) );
  AND U42629 ( .A(mul_pow), .B(n40365), .Z(n40364) );
  XOR U42630 ( .A(ein[810]), .B(ein[809]), .Z(n40365) );
  XOR U42631 ( .A(ein[79]), .B(n40366), .Z(ereg_next[80]) );
  AND U42632 ( .A(mul_pow), .B(n40367), .Z(n40366) );
  XOR U42633 ( .A(ein[80]), .B(ein[79]), .Z(n40367) );
  XOR U42634 ( .A(ein[808]), .B(n40368), .Z(ereg_next[809]) );
  AND U42635 ( .A(mul_pow), .B(n40369), .Z(n40368) );
  XOR U42636 ( .A(ein[809]), .B(ein[808]), .Z(n40369) );
  XOR U42637 ( .A(ein[807]), .B(n40370), .Z(ereg_next[808]) );
  AND U42638 ( .A(mul_pow), .B(n40371), .Z(n40370) );
  XOR U42639 ( .A(ein[808]), .B(ein[807]), .Z(n40371) );
  XOR U42640 ( .A(ein[806]), .B(n40372), .Z(ereg_next[807]) );
  AND U42641 ( .A(mul_pow), .B(n40373), .Z(n40372) );
  XOR U42642 ( .A(ein[807]), .B(ein[806]), .Z(n40373) );
  XOR U42643 ( .A(ein[805]), .B(n40374), .Z(ereg_next[806]) );
  AND U42644 ( .A(mul_pow), .B(n40375), .Z(n40374) );
  XOR U42645 ( .A(ein[806]), .B(ein[805]), .Z(n40375) );
  XOR U42646 ( .A(ein[804]), .B(n40376), .Z(ereg_next[805]) );
  AND U42647 ( .A(mul_pow), .B(n40377), .Z(n40376) );
  XOR U42648 ( .A(ein[805]), .B(ein[804]), .Z(n40377) );
  XOR U42649 ( .A(ein[803]), .B(n40378), .Z(ereg_next[804]) );
  AND U42650 ( .A(mul_pow), .B(n40379), .Z(n40378) );
  XOR U42651 ( .A(ein[804]), .B(ein[803]), .Z(n40379) );
  XOR U42652 ( .A(ein[802]), .B(n40380), .Z(ereg_next[803]) );
  AND U42653 ( .A(mul_pow), .B(n40381), .Z(n40380) );
  XOR U42654 ( .A(ein[803]), .B(ein[802]), .Z(n40381) );
  XOR U42655 ( .A(ein[801]), .B(n40382), .Z(ereg_next[802]) );
  AND U42656 ( .A(mul_pow), .B(n40383), .Z(n40382) );
  XOR U42657 ( .A(ein[802]), .B(ein[801]), .Z(n40383) );
  XOR U42658 ( .A(ein[800]), .B(n40384), .Z(ereg_next[801]) );
  AND U42659 ( .A(mul_pow), .B(n40385), .Z(n40384) );
  XOR U42660 ( .A(ein[801]), .B(ein[800]), .Z(n40385) );
  XOR U42661 ( .A(ein[799]), .B(n40386), .Z(ereg_next[800]) );
  AND U42662 ( .A(mul_pow), .B(n40387), .Z(n40386) );
  XOR U42663 ( .A(ein[800]), .B(ein[799]), .Z(n40387) );
  XOR U42664 ( .A(ein[6]), .B(n40388), .Z(ereg_next[7]) );
  AND U42665 ( .A(mul_pow), .B(n40389), .Z(n40388) );
  XOR U42666 ( .A(ein[7]), .B(ein[6]), .Z(n40389) );
  XOR U42667 ( .A(ein[78]), .B(n40390), .Z(ereg_next[79]) );
  AND U42668 ( .A(mul_pow), .B(n40391), .Z(n40390) );
  XOR U42669 ( .A(ein[79]), .B(ein[78]), .Z(n40391) );
  XOR U42670 ( .A(ein[798]), .B(n40392), .Z(ereg_next[799]) );
  AND U42671 ( .A(mul_pow), .B(n40393), .Z(n40392) );
  XOR U42672 ( .A(ein[799]), .B(ein[798]), .Z(n40393) );
  XOR U42673 ( .A(ein[797]), .B(n40394), .Z(ereg_next[798]) );
  AND U42674 ( .A(mul_pow), .B(n40395), .Z(n40394) );
  XOR U42675 ( .A(ein[798]), .B(ein[797]), .Z(n40395) );
  XOR U42676 ( .A(ein[796]), .B(n40396), .Z(ereg_next[797]) );
  AND U42677 ( .A(mul_pow), .B(n40397), .Z(n40396) );
  XOR U42678 ( .A(ein[797]), .B(ein[796]), .Z(n40397) );
  XOR U42679 ( .A(ein[795]), .B(n40398), .Z(ereg_next[796]) );
  AND U42680 ( .A(mul_pow), .B(n40399), .Z(n40398) );
  XOR U42681 ( .A(ein[796]), .B(ein[795]), .Z(n40399) );
  XOR U42682 ( .A(ein[794]), .B(n40400), .Z(ereg_next[795]) );
  AND U42683 ( .A(mul_pow), .B(n40401), .Z(n40400) );
  XOR U42684 ( .A(ein[795]), .B(ein[794]), .Z(n40401) );
  XOR U42685 ( .A(ein[793]), .B(n40402), .Z(ereg_next[794]) );
  AND U42686 ( .A(mul_pow), .B(n40403), .Z(n40402) );
  XOR U42687 ( .A(ein[794]), .B(ein[793]), .Z(n40403) );
  XOR U42688 ( .A(ein[792]), .B(n40404), .Z(ereg_next[793]) );
  AND U42689 ( .A(mul_pow), .B(n40405), .Z(n40404) );
  XOR U42690 ( .A(ein[793]), .B(ein[792]), .Z(n40405) );
  XOR U42691 ( .A(ein[791]), .B(n40406), .Z(ereg_next[792]) );
  AND U42692 ( .A(mul_pow), .B(n40407), .Z(n40406) );
  XOR U42693 ( .A(ein[792]), .B(ein[791]), .Z(n40407) );
  XOR U42694 ( .A(ein[790]), .B(n40408), .Z(ereg_next[791]) );
  AND U42695 ( .A(mul_pow), .B(n40409), .Z(n40408) );
  XOR U42696 ( .A(ein[791]), .B(ein[790]), .Z(n40409) );
  XOR U42697 ( .A(ein[789]), .B(n40410), .Z(ereg_next[790]) );
  AND U42698 ( .A(mul_pow), .B(n40411), .Z(n40410) );
  XOR U42699 ( .A(ein[790]), .B(ein[789]), .Z(n40411) );
  XOR U42700 ( .A(ein[77]), .B(n40412), .Z(ereg_next[78]) );
  AND U42701 ( .A(mul_pow), .B(n40413), .Z(n40412) );
  XOR U42702 ( .A(ein[78]), .B(ein[77]), .Z(n40413) );
  XOR U42703 ( .A(ein[788]), .B(n40414), .Z(ereg_next[789]) );
  AND U42704 ( .A(mul_pow), .B(n40415), .Z(n40414) );
  XOR U42705 ( .A(ein[789]), .B(ein[788]), .Z(n40415) );
  XOR U42706 ( .A(ein[787]), .B(n40416), .Z(ereg_next[788]) );
  AND U42707 ( .A(mul_pow), .B(n40417), .Z(n40416) );
  XOR U42708 ( .A(ein[788]), .B(ein[787]), .Z(n40417) );
  XOR U42709 ( .A(ein[786]), .B(n40418), .Z(ereg_next[787]) );
  AND U42710 ( .A(mul_pow), .B(n40419), .Z(n40418) );
  XOR U42711 ( .A(ein[787]), .B(ein[786]), .Z(n40419) );
  XOR U42712 ( .A(ein[785]), .B(n40420), .Z(ereg_next[786]) );
  AND U42713 ( .A(mul_pow), .B(n40421), .Z(n40420) );
  XOR U42714 ( .A(ein[786]), .B(ein[785]), .Z(n40421) );
  XOR U42715 ( .A(ein[784]), .B(n40422), .Z(ereg_next[785]) );
  AND U42716 ( .A(mul_pow), .B(n40423), .Z(n40422) );
  XOR U42717 ( .A(ein[785]), .B(ein[784]), .Z(n40423) );
  XOR U42718 ( .A(ein[783]), .B(n40424), .Z(ereg_next[784]) );
  AND U42719 ( .A(mul_pow), .B(n40425), .Z(n40424) );
  XOR U42720 ( .A(ein[784]), .B(ein[783]), .Z(n40425) );
  XOR U42721 ( .A(ein[782]), .B(n40426), .Z(ereg_next[783]) );
  AND U42722 ( .A(mul_pow), .B(n40427), .Z(n40426) );
  XOR U42723 ( .A(ein[783]), .B(ein[782]), .Z(n40427) );
  XOR U42724 ( .A(ein[781]), .B(n40428), .Z(ereg_next[782]) );
  AND U42725 ( .A(mul_pow), .B(n40429), .Z(n40428) );
  XOR U42726 ( .A(ein[782]), .B(ein[781]), .Z(n40429) );
  XOR U42727 ( .A(ein[780]), .B(n40430), .Z(ereg_next[781]) );
  AND U42728 ( .A(mul_pow), .B(n40431), .Z(n40430) );
  XOR U42729 ( .A(ein[781]), .B(ein[780]), .Z(n40431) );
  XOR U42730 ( .A(ein[779]), .B(n40432), .Z(ereg_next[780]) );
  AND U42731 ( .A(mul_pow), .B(n40433), .Z(n40432) );
  XOR U42732 ( .A(ein[780]), .B(ein[779]), .Z(n40433) );
  XOR U42733 ( .A(ein[76]), .B(n40434), .Z(ereg_next[77]) );
  AND U42734 ( .A(mul_pow), .B(n40435), .Z(n40434) );
  XOR U42735 ( .A(ein[77]), .B(ein[76]), .Z(n40435) );
  XOR U42736 ( .A(ein[778]), .B(n40436), .Z(ereg_next[779]) );
  AND U42737 ( .A(mul_pow), .B(n40437), .Z(n40436) );
  XOR U42738 ( .A(ein[779]), .B(ein[778]), .Z(n40437) );
  XOR U42739 ( .A(ein[777]), .B(n40438), .Z(ereg_next[778]) );
  AND U42740 ( .A(mul_pow), .B(n40439), .Z(n40438) );
  XOR U42741 ( .A(ein[778]), .B(ein[777]), .Z(n40439) );
  XOR U42742 ( .A(ein[776]), .B(n40440), .Z(ereg_next[777]) );
  AND U42743 ( .A(mul_pow), .B(n40441), .Z(n40440) );
  XOR U42744 ( .A(ein[777]), .B(ein[776]), .Z(n40441) );
  XOR U42745 ( .A(ein[775]), .B(n40442), .Z(ereg_next[776]) );
  AND U42746 ( .A(mul_pow), .B(n40443), .Z(n40442) );
  XOR U42747 ( .A(ein[776]), .B(ein[775]), .Z(n40443) );
  XOR U42748 ( .A(ein[774]), .B(n40444), .Z(ereg_next[775]) );
  AND U42749 ( .A(mul_pow), .B(n40445), .Z(n40444) );
  XOR U42750 ( .A(ein[775]), .B(ein[774]), .Z(n40445) );
  XOR U42751 ( .A(ein[773]), .B(n40446), .Z(ereg_next[774]) );
  AND U42752 ( .A(mul_pow), .B(n40447), .Z(n40446) );
  XOR U42753 ( .A(ein[774]), .B(ein[773]), .Z(n40447) );
  XOR U42754 ( .A(ein[772]), .B(n40448), .Z(ereg_next[773]) );
  AND U42755 ( .A(mul_pow), .B(n40449), .Z(n40448) );
  XOR U42756 ( .A(ein[773]), .B(ein[772]), .Z(n40449) );
  XOR U42757 ( .A(ein[771]), .B(n40450), .Z(ereg_next[772]) );
  AND U42758 ( .A(mul_pow), .B(n40451), .Z(n40450) );
  XOR U42759 ( .A(ein[772]), .B(ein[771]), .Z(n40451) );
  XOR U42760 ( .A(ein[770]), .B(n40452), .Z(ereg_next[771]) );
  AND U42761 ( .A(mul_pow), .B(n40453), .Z(n40452) );
  XOR U42762 ( .A(ein[771]), .B(ein[770]), .Z(n40453) );
  XOR U42763 ( .A(ein[769]), .B(n40454), .Z(ereg_next[770]) );
  AND U42764 ( .A(mul_pow), .B(n40455), .Z(n40454) );
  XOR U42765 ( .A(ein[770]), .B(ein[769]), .Z(n40455) );
  XOR U42766 ( .A(ein[75]), .B(n40456), .Z(ereg_next[76]) );
  AND U42767 ( .A(mul_pow), .B(n40457), .Z(n40456) );
  XOR U42768 ( .A(ein[76]), .B(ein[75]), .Z(n40457) );
  XOR U42769 ( .A(ein[768]), .B(n40458), .Z(ereg_next[769]) );
  AND U42770 ( .A(mul_pow), .B(n40459), .Z(n40458) );
  XOR U42771 ( .A(ein[769]), .B(ein[768]), .Z(n40459) );
  XOR U42772 ( .A(ein[767]), .B(n40460), .Z(ereg_next[768]) );
  AND U42773 ( .A(mul_pow), .B(n40461), .Z(n40460) );
  XOR U42774 ( .A(ein[768]), .B(ein[767]), .Z(n40461) );
  XOR U42775 ( .A(ein[766]), .B(n40462), .Z(ereg_next[767]) );
  AND U42776 ( .A(mul_pow), .B(n40463), .Z(n40462) );
  XOR U42777 ( .A(ein[767]), .B(ein[766]), .Z(n40463) );
  XOR U42778 ( .A(ein[765]), .B(n40464), .Z(ereg_next[766]) );
  AND U42779 ( .A(mul_pow), .B(n40465), .Z(n40464) );
  XOR U42780 ( .A(ein[766]), .B(ein[765]), .Z(n40465) );
  XOR U42781 ( .A(ein[764]), .B(n40466), .Z(ereg_next[765]) );
  AND U42782 ( .A(mul_pow), .B(n40467), .Z(n40466) );
  XOR U42783 ( .A(ein[765]), .B(ein[764]), .Z(n40467) );
  XOR U42784 ( .A(ein[763]), .B(n40468), .Z(ereg_next[764]) );
  AND U42785 ( .A(mul_pow), .B(n40469), .Z(n40468) );
  XOR U42786 ( .A(ein[764]), .B(ein[763]), .Z(n40469) );
  XOR U42787 ( .A(ein[762]), .B(n40470), .Z(ereg_next[763]) );
  AND U42788 ( .A(mul_pow), .B(n40471), .Z(n40470) );
  XOR U42789 ( .A(ein[763]), .B(ein[762]), .Z(n40471) );
  XOR U42790 ( .A(ein[761]), .B(n40472), .Z(ereg_next[762]) );
  AND U42791 ( .A(mul_pow), .B(n40473), .Z(n40472) );
  XOR U42792 ( .A(ein[762]), .B(ein[761]), .Z(n40473) );
  XOR U42793 ( .A(ein[760]), .B(n40474), .Z(ereg_next[761]) );
  AND U42794 ( .A(mul_pow), .B(n40475), .Z(n40474) );
  XOR U42795 ( .A(ein[761]), .B(ein[760]), .Z(n40475) );
  XOR U42796 ( .A(ein[759]), .B(n40476), .Z(ereg_next[760]) );
  AND U42797 ( .A(mul_pow), .B(n40477), .Z(n40476) );
  XOR U42798 ( .A(ein[760]), .B(ein[759]), .Z(n40477) );
  XOR U42799 ( .A(ein[74]), .B(n40478), .Z(ereg_next[75]) );
  AND U42800 ( .A(mul_pow), .B(n40479), .Z(n40478) );
  XOR U42801 ( .A(ein[75]), .B(ein[74]), .Z(n40479) );
  XOR U42802 ( .A(ein[758]), .B(n40480), .Z(ereg_next[759]) );
  AND U42803 ( .A(mul_pow), .B(n40481), .Z(n40480) );
  XOR U42804 ( .A(ein[759]), .B(ein[758]), .Z(n40481) );
  XOR U42805 ( .A(ein[757]), .B(n40482), .Z(ereg_next[758]) );
  AND U42806 ( .A(mul_pow), .B(n40483), .Z(n40482) );
  XOR U42807 ( .A(ein[758]), .B(ein[757]), .Z(n40483) );
  XOR U42808 ( .A(ein[756]), .B(n40484), .Z(ereg_next[757]) );
  AND U42809 ( .A(mul_pow), .B(n40485), .Z(n40484) );
  XOR U42810 ( .A(ein[757]), .B(ein[756]), .Z(n40485) );
  XOR U42811 ( .A(ein[755]), .B(n40486), .Z(ereg_next[756]) );
  AND U42812 ( .A(mul_pow), .B(n40487), .Z(n40486) );
  XOR U42813 ( .A(ein[756]), .B(ein[755]), .Z(n40487) );
  XOR U42814 ( .A(ein[754]), .B(n40488), .Z(ereg_next[755]) );
  AND U42815 ( .A(mul_pow), .B(n40489), .Z(n40488) );
  XOR U42816 ( .A(ein[755]), .B(ein[754]), .Z(n40489) );
  XOR U42817 ( .A(ein[753]), .B(n40490), .Z(ereg_next[754]) );
  AND U42818 ( .A(mul_pow), .B(n40491), .Z(n40490) );
  XOR U42819 ( .A(ein[754]), .B(ein[753]), .Z(n40491) );
  XOR U42820 ( .A(ein[752]), .B(n40492), .Z(ereg_next[753]) );
  AND U42821 ( .A(mul_pow), .B(n40493), .Z(n40492) );
  XOR U42822 ( .A(ein[753]), .B(ein[752]), .Z(n40493) );
  XOR U42823 ( .A(ein[751]), .B(n40494), .Z(ereg_next[752]) );
  AND U42824 ( .A(mul_pow), .B(n40495), .Z(n40494) );
  XOR U42825 ( .A(ein[752]), .B(ein[751]), .Z(n40495) );
  XOR U42826 ( .A(ein[750]), .B(n40496), .Z(ereg_next[751]) );
  AND U42827 ( .A(mul_pow), .B(n40497), .Z(n40496) );
  XOR U42828 ( .A(ein[751]), .B(ein[750]), .Z(n40497) );
  XOR U42829 ( .A(ein[749]), .B(n40498), .Z(ereg_next[750]) );
  AND U42830 ( .A(mul_pow), .B(n40499), .Z(n40498) );
  XOR U42831 ( .A(ein[750]), .B(ein[749]), .Z(n40499) );
  XOR U42832 ( .A(ein[73]), .B(n40500), .Z(ereg_next[74]) );
  AND U42833 ( .A(mul_pow), .B(n40501), .Z(n40500) );
  XOR U42834 ( .A(ein[74]), .B(ein[73]), .Z(n40501) );
  XOR U42835 ( .A(ein[748]), .B(n40502), .Z(ereg_next[749]) );
  AND U42836 ( .A(mul_pow), .B(n40503), .Z(n40502) );
  XOR U42837 ( .A(ein[749]), .B(ein[748]), .Z(n40503) );
  XOR U42838 ( .A(ein[747]), .B(n40504), .Z(ereg_next[748]) );
  AND U42839 ( .A(mul_pow), .B(n40505), .Z(n40504) );
  XOR U42840 ( .A(ein[748]), .B(ein[747]), .Z(n40505) );
  XOR U42841 ( .A(ein[746]), .B(n40506), .Z(ereg_next[747]) );
  AND U42842 ( .A(mul_pow), .B(n40507), .Z(n40506) );
  XOR U42843 ( .A(ein[747]), .B(ein[746]), .Z(n40507) );
  XOR U42844 ( .A(ein[745]), .B(n40508), .Z(ereg_next[746]) );
  AND U42845 ( .A(mul_pow), .B(n40509), .Z(n40508) );
  XOR U42846 ( .A(ein[746]), .B(ein[745]), .Z(n40509) );
  XOR U42847 ( .A(ein[744]), .B(n40510), .Z(ereg_next[745]) );
  AND U42848 ( .A(mul_pow), .B(n40511), .Z(n40510) );
  XOR U42849 ( .A(ein[745]), .B(ein[744]), .Z(n40511) );
  XOR U42850 ( .A(ein[743]), .B(n40512), .Z(ereg_next[744]) );
  AND U42851 ( .A(mul_pow), .B(n40513), .Z(n40512) );
  XOR U42852 ( .A(ein[744]), .B(ein[743]), .Z(n40513) );
  XOR U42853 ( .A(ein[742]), .B(n40514), .Z(ereg_next[743]) );
  AND U42854 ( .A(mul_pow), .B(n40515), .Z(n40514) );
  XOR U42855 ( .A(ein[743]), .B(ein[742]), .Z(n40515) );
  XOR U42856 ( .A(ein[741]), .B(n40516), .Z(ereg_next[742]) );
  AND U42857 ( .A(mul_pow), .B(n40517), .Z(n40516) );
  XOR U42858 ( .A(ein[742]), .B(ein[741]), .Z(n40517) );
  XOR U42859 ( .A(ein[740]), .B(n40518), .Z(ereg_next[741]) );
  AND U42860 ( .A(mul_pow), .B(n40519), .Z(n40518) );
  XOR U42861 ( .A(ein[741]), .B(ein[740]), .Z(n40519) );
  XOR U42862 ( .A(ein[739]), .B(n40520), .Z(ereg_next[740]) );
  AND U42863 ( .A(mul_pow), .B(n40521), .Z(n40520) );
  XOR U42864 ( .A(ein[740]), .B(ein[739]), .Z(n40521) );
  XOR U42865 ( .A(ein[72]), .B(n40522), .Z(ereg_next[73]) );
  AND U42866 ( .A(mul_pow), .B(n40523), .Z(n40522) );
  XOR U42867 ( .A(ein[73]), .B(ein[72]), .Z(n40523) );
  XOR U42868 ( .A(ein[738]), .B(n40524), .Z(ereg_next[739]) );
  AND U42869 ( .A(mul_pow), .B(n40525), .Z(n40524) );
  XOR U42870 ( .A(ein[739]), .B(ein[738]), .Z(n40525) );
  XOR U42871 ( .A(ein[737]), .B(n40526), .Z(ereg_next[738]) );
  AND U42872 ( .A(mul_pow), .B(n40527), .Z(n40526) );
  XOR U42873 ( .A(ein[738]), .B(ein[737]), .Z(n40527) );
  XOR U42874 ( .A(ein[736]), .B(n40528), .Z(ereg_next[737]) );
  AND U42875 ( .A(mul_pow), .B(n40529), .Z(n40528) );
  XOR U42876 ( .A(ein[737]), .B(ein[736]), .Z(n40529) );
  XOR U42877 ( .A(ein[735]), .B(n40530), .Z(ereg_next[736]) );
  AND U42878 ( .A(mul_pow), .B(n40531), .Z(n40530) );
  XOR U42879 ( .A(ein[736]), .B(ein[735]), .Z(n40531) );
  XOR U42880 ( .A(ein[734]), .B(n40532), .Z(ereg_next[735]) );
  AND U42881 ( .A(mul_pow), .B(n40533), .Z(n40532) );
  XOR U42882 ( .A(ein[735]), .B(ein[734]), .Z(n40533) );
  XOR U42883 ( .A(ein[733]), .B(n40534), .Z(ereg_next[734]) );
  AND U42884 ( .A(mul_pow), .B(n40535), .Z(n40534) );
  XOR U42885 ( .A(ein[734]), .B(ein[733]), .Z(n40535) );
  XOR U42886 ( .A(ein[732]), .B(n40536), .Z(ereg_next[733]) );
  AND U42887 ( .A(mul_pow), .B(n40537), .Z(n40536) );
  XOR U42888 ( .A(ein[733]), .B(ein[732]), .Z(n40537) );
  XOR U42889 ( .A(ein[731]), .B(n40538), .Z(ereg_next[732]) );
  AND U42890 ( .A(mul_pow), .B(n40539), .Z(n40538) );
  XOR U42891 ( .A(ein[732]), .B(ein[731]), .Z(n40539) );
  XOR U42892 ( .A(ein[730]), .B(n40540), .Z(ereg_next[731]) );
  AND U42893 ( .A(mul_pow), .B(n40541), .Z(n40540) );
  XOR U42894 ( .A(ein[731]), .B(ein[730]), .Z(n40541) );
  XOR U42895 ( .A(ein[729]), .B(n40542), .Z(ereg_next[730]) );
  AND U42896 ( .A(mul_pow), .B(n40543), .Z(n40542) );
  XOR U42897 ( .A(ein[730]), .B(ein[729]), .Z(n40543) );
  XOR U42898 ( .A(ein[71]), .B(n40544), .Z(ereg_next[72]) );
  AND U42899 ( .A(mul_pow), .B(n40545), .Z(n40544) );
  XOR U42900 ( .A(ein[72]), .B(ein[71]), .Z(n40545) );
  XOR U42901 ( .A(ein[728]), .B(n40546), .Z(ereg_next[729]) );
  AND U42902 ( .A(mul_pow), .B(n40547), .Z(n40546) );
  XOR U42903 ( .A(ein[729]), .B(ein[728]), .Z(n40547) );
  XOR U42904 ( .A(ein[727]), .B(n40548), .Z(ereg_next[728]) );
  AND U42905 ( .A(mul_pow), .B(n40549), .Z(n40548) );
  XOR U42906 ( .A(ein[728]), .B(ein[727]), .Z(n40549) );
  XOR U42907 ( .A(ein[726]), .B(n40550), .Z(ereg_next[727]) );
  AND U42908 ( .A(mul_pow), .B(n40551), .Z(n40550) );
  XOR U42909 ( .A(ein[727]), .B(ein[726]), .Z(n40551) );
  XOR U42910 ( .A(ein[725]), .B(n40552), .Z(ereg_next[726]) );
  AND U42911 ( .A(mul_pow), .B(n40553), .Z(n40552) );
  XOR U42912 ( .A(ein[726]), .B(ein[725]), .Z(n40553) );
  XOR U42913 ( .A(ein[724]), .B(n40554), .Z(ereg_next[725]) );
  AND U42914 ( .A(mul_pow), .B(n40555), .Z(n40554) );
  XOR U42915 ( .A(ein[725]), .B(ein[724]), .Z(n40555) );
  XOR U42916 ( .A(ein[723]), .B(n40556), .Z(ereg_next[724]) );
  AND U42917 ( .A(mul_pow), .B(n40557), .Z(n40556) );
  XOR U42918 ( .A(ein[724]), .B(ein[723]), .Z(n40557) );
  XOR U42919 ( .A(ein[722]), .B(n40558), .Z(ereg_next[723]) );
  AND U42920 ( .A(mul_pow), .B(n40559), .Z(n40558) );
  XOR U42921 ( .A(ein[723]), .B(ein[722]), .Z(n40559) );
  XOR U42922 ( .A(ein[721]), .B(n40560), .Z(ereg_next[722]) );
  AND U42923 ( .A(mul_pow), .B(n40561), .Z(n40560) );
  XOR U42924 ( .A(ein[722]), .B(ein[721]), .Z(n40561) );
  XOR U42925 ( .A(ein[720]), .B(n40562), .Z(ereg_next[721]) );
  AND U42926 ( .A(mul_pow), .B(n40563), .Z(n40562) );
  XOR U42927 ( .A(ein[721]), .B(ein[720]), .Z(n40563) );
  XOR U42928 ( .A(ein[719]), .B(n40564), .Z(ereg_next[720]) );
  AND U42929 ( .A(mul_pow), .B(n40565), .Z(n40564) );
  XOR U42930 ( .A(ein[720]), .B(ein[719]), .Z(n40565) );
  XOR U42931 ( .A(ein[70]), .B(n40566), .Z(ereg_next[71]) );
  AND U42932 ( .A(mul_pow), .B(n40567), .Z(n40566) );
  XOR U42933 ( .A(ein[71]), .B(ein[70]), .Z(n40567) );
  XOR U42934 ( .A(ein[718]), .B(n40568), .Z(ereg_next[719]) );
  AND U42935 ( .A(mul_pow), .B(n40569), .Z(n40568) );
  XOR U42936 ( .A(ein[719]), .B(ein[718]), .Z(n40569) );
  XOR U42937 ( .A(ein[717]), .B(n40570), .Z(ereg_next[718]) );
  AND U42938 ( .A(mul_pow), .B(n40571), .Z(n40570) );
  XOR U42939 ( .A(ein[718]), .B(ein[717]), .Z(n40571) );
  XOR U42940 ( .A(ein[716]), .B(n40572), .Z(ereg_next[717]) );
  AND U42941 ( .A(mul_pow), .B(n40573), .Z(n40572) );
  XOR U42942 ( .A(ein[717]), .B(ein[716]), .Z(n40573) );
  XOR U42943 ( .A(ein[715]), .B(n40574), .Z(ereg_next[716]) );
  AND U42944 ( .A(mul_pow), .B(n40575), .Z(n40574) );
  XOR U42945 ( .A(ein[716]), .B(ein[715]), .Z(n40575) );
  XOR U42946 ( .A(ein[714]), .B(n40576), .Z(ereg_next[715]) );
  AND U42947 ( .A(mul_pow), .B(n40577), .Z(n40576) );
  XOR U42948 ( .A(ein[715]), .B(ein[714]), .Z(n40577) );
  XOR U42949 ( .A(ein[713]), .B(n40578), .Z(ereg_next[714]) );
  AND U42950 ( .A(mul_pow), .B(n40579), .Z(n40578) );
  XOR U42951 ( .A(ein[714]), .B(ein[713]), .Z(n40579) );
  XOR U42952 ( .A(ein[712]), .B(n40580), .Z(ereg_next[713]) );
  AND U42953 ( .A(mul_pow), .B(n40581), .Z(n40580) );
  XOR U42954 ( .A(ein[713]), .B(ein[712]), .Z(n40581) );
  XOR U42955 ( .A(ein[711]), .B(n40582), .Z(ereg_next[712]) );
  AND U42956 ( .A(mul_pow), .B(n40583), .Z(n40582) );
  XOR U42957 ( .A(ein[712]), .B(ein[711]), .Z(n40583) );
  XOR U42958 ( .A(ein[710]), .B(n40584), .Z(ereg_next[711]) );
  AND U42959 ( .A(mul_pow), .B(n40585), .Z(n40584) );
  XOR U42960 ( .A(ein[711]), .B(ein[710]), .Z(n40585) );
  XOR U42961 ( .A(ein[709]), .B(n40586), .Z(ereg_next[710]) );
  AND U42962 ( .A(mul_pow), .B(n40587), .Z(n40586) );
  XOR U42963 ( .A(ein[710]), .B(ein[709]), .Z(n40587) );
  XOR U42964 ( .A(ein[69]), .B(n40588), .Z(ereg_next[70]) );
  AND U42965 ( .A(mul_pow), .B(n40589), .Z(n40588) );
  XOR U42966 ( .A(ein[70]), .B(ein[69]), .Z(n40589) );
  XOR U42967 ( .A(ein[708]), .B(n40590), .Z(ereg_next[709]) );
  AND U42968 ( .A(mul_pow), .B(n40591), .Z(n40590) );
  XOR U42969 ( .A(ein[709]), .B(ein[708]), .Z(n40591) );
  XOR U42970 ( .A(ein[707]), .B(n40592), .Z(ereg_next[708]) );
  AND U42971 ( .A(mul_pow), .B(n40593), .Z(n40592) );
  XOR U42972 ( .A(ein[708]), .B(ein[707]), .Z(n40593) );
  XOR U42973 ( .A(ein[706]), .B(n40594), .Z(ereg_next[707]) );
  AND U42974 ( .A(mul_pow), .B(n40595), .Z(n40594) );
  XOR U42975 ( .A(ein[707]), .B(ein[706]), .Z(n40595) );
  XOR U42976 ( .A(ein[705]), .B(n40596), .Z(ereg_next[706]) );
  AND U42977 ( .A(mul_pow), .B(n40597), .Z(n40596) );
  XOR U42978 ( .A(ein[706]), .B(ein[705]), .Z(n40597) );
  XOR U42979 ( .A(ein[704]), .B(n40598), .Z(ereg_next[705]) );
  AND U42980 ( .A(mul_pow), .B(n40599), .Z(n40598) );
  XOR U42981 ( .A(ein[705]), .B(ein[704]), .Z(n40599) );
  XOR U42982 ( .A(ein[703]), .B(n40600), .Z(ereg_next[704]) );
  AND U42983 ( .A(mul_pow), .B(n40601), .Z(n40600) );
  XOR U42984 ( .A(ein[704]), .B(ein[703]), .Z(n40601) );
  XOR U42985 ( .A(ein[702]), .B(n40602), .Z(ereg_next[703]) );
  AND U42986 ( .A(mul_pow), .B(n40603), .Z(n40602) );
  XOR U42987 ( .A(ein[703]), .B(ein[702]), .Z(n40603) );
  XOR U42988 ( .A(ein[701]), .B(n40604), .Z(ereg_next[702]) );
  AND U42989 ( .A(mul_pow), .B(n40605), .Z(n40604) );
  XOR U42990 ( .A(ein[702]), .B(ein[701]), .Z(n40605) );
  XOR U42991 ( .A(ein[700]), .B(n40606), .Z(ereg_next[701]) );
  AND U42992 ( .A(mul_pow), .B(n40607), .Z(n40606) );
  XOR U42993 ( .A(ein[701]), .B(ein[700]), .Z(n40607) );
  XOR U42994 ( .A(ein[699]), .B(n40608), .Z(ereg_next[700]) );
  AND U42995 ( .A(mul_pow), .B(n40609), .Z(n40608) );
  XOR U42996 ( .A(ein[700]), .B(ein[699]), .Z(n40609) );
  XOR U42997 ( .A(ein[5]), .B(n40610), .Z(ereg_next[6]) );
  AND U42998 ( .A(mul_pow), .B(n40611), .Z(n40610) );
  XOR U42999 ( .A(ein[6]), .B(ein[5]), .Z(n40611) );
  XOR U43000 ( .A(ein[68]), .B(n40612), .Z(ereg_next[69]) );
  AND U43001 ( .A(mul_pow), .B(n40613), .Z(n40612) );
  XOR U43002 ( .A(ein[69]), .B(ein[68]), .Z(n40613) );
  XOR U43003 ( .A(ein[698]), .B(n40614), .Z(ereg_next[699]) );
  AND U43004 ( .A(mul_pow), .B(n40615), .Z(n40614) );
  XOR U43005 ( .A(ein[699]), .B(ein[698]), .Z(n40615) );
  XOR U43006 ( .A(ein[697]), .B(n40616), .Z(ereg_next[698]) );
  AND U43007 ( .A(mul_pow), .B(n40617), .Z(n40616) );
  XOR U43008 ( .A(ein[698]), .B(ein[697]), .Z(n40617) );
  XOR U43009 ( .A(ein[696]), .B(n40618), .Z(ereg_next[697]) );
  AND U43010 ( .A(mul_pow), .B(n40619), .Z(n40618) );
  XOR U43011 ( .A(ein[697]), .B(ein[696]), .Z(n40619) );
  XOR U43012 ( .A(ein[695]), .B(n40620), .Z(ereg_next[696]) );
  AND U43013 ( .A(mul_pow), .B(n40621), .Z(n40620) );
  XOR U43014 ( .A(ein[696]), .B(ein[695]), .Z(n40621) );
  XOR U43015 ( .A(ein[694]), .B(n40622), .Z(ereg_next[695]) );
  AND U43016 ( .A(mul_pow), .B(n40623), .Z(n40622) );
  XOR U43017 ( .A(ein[695]), .B(ein[694]), .Z(n40623) );
  XOR U43018 ( .A(ein[693]), .B(n40624), .Z(ereg_next[694]) );
  AND U43019 ( .A(mul_pow), .B(n40625), .Z(n40624) );
  XOR U43020 ( .A(ein[694]), .B(ein[693]), .Z(n40625) );
  XOR U43021 ( .A(ein[692]), .B(n40626), .Z(ereg_next[693]) );
  AND U43022 ( .A(mul_pow), .B(n40627), .Z(n40626) );
  XOR U43023 ( .A(ein[693]), .B(ein[692]), .Z(n40627) );
  XOR U43024 ( .A(ein[691]), .B(n40628), .Z(ereg_next[692]) );
  AND U43025 ( .A(mul_pow), .B(n40629), .Z(n40628) );
  XOR U43026 ( .A(ein[692]), .B(ein[691]), .Z(n40629) );
  XOR U43027 ( .A(ein[690]), .B(n40630), .Z(ereg_next[691]) );
  AND U43028 ( .A(mul_pow), .B(n40631), .Z(n40630) );
  XOR U43029 ( .A(ein[691]), .B(ein[690]), .Z(n40631) );
  XOR U43030 ( .A(ein[689]), .B(n40632), .Z(ereg_next[690]) );
  AND U43031 ( .A(mul_pow), .B(n40633), .Z(n40632) );
  XOR U43032 ( .A(ein[690]), .B(ein[689]), .Z(n40633) );
  XOR U43033 ( .A(ein[67]), .B(n40634), .Z(ereg_next[68]) );
  AND U43034 ( .A(mul_pow), .B(n40635), .Z(n40634) );
  XOR U43035 ( .A(ein[68]), .B(ein[67]), .Z(n40635) );
  XOR U43036 ( .A(ein[688]), .B(n40636), .Z(ereg_next[689]) );
  AND U43037 ( .A(mul_pow), .B(n40637), .Z(n40636) );
  XOR U43038 ( .A(ein[689]), .B(ein[688]), .Z(n40637) );
  XOR U43039 ( .A(ein[687]), .B(n40638), .Z(ereg_next[688]) );
  AND U43040 ( .A(mul_pow), .B(n40639), .Z(n40638) );
  XOR U43041 ( .A(ein[688]), .B(ein[687]), .Z(n40639) );
  XOR U43042 ( .A(ein[686]), .B(n40640), .Z(ereg_next[687]) );
  AND U43043 ( .A(mul_pow), .B(n40641), .Z(n40640) );
  XOR U43044 ( .A(ein[687]), .B(ein[686]), .Z(n40641) );
  XOR U43045 ( .A(ein[685]), .B(n40642), .Z(ereg_next[686]) );
  AND U43046 ( .A(mul_pow), .B(n40643), .Z(n40642) );
  XOR U43047 ( .A(ein[686]), .B(ein[685]), .Z(n40643) );
  XOR U43048 ( .A(ein[684]), .B(n40644), .Z(ereg_next[685]) );
  AND U43049 ( .A(mul_pow), .B(n40645), .Z(n40644) );
  XOR U43050 ( .A(ein[685]), .B(ein[684]), .Z(n40645) );
  XOR U43051 ( .A(ein[683]), .B(n40646), .Z(ereg_next[684]) );
  AND U43052 ( .A(mul_pow), .B(n40647), .Z(n40646) );
  XOR U43053 ( .A(ein[684]), .B(ein[683]), .Z(n40647) );
  XOR U43054 ( .A(ein[682]), .B(n40648), .Z(ereg_next[683]) );
  AND U43055 ( .A(mul_pow), .B(n40649), .Z(n40648) );
  XOR U43056 ( .A(ein[683]), .B(ein[682]), .Z(n40649) );
  XOR U43057 ( .A(ein[681]), .B(n40650), .Z(ereg_next[682]) );
  AND U43058 ( .A(mul_pow), .B(n40651), .Z(n40650) );
  XOR U43059 ( .A(ein[682]), .B(ein[681]), .Z(n40651) );
  XOR U43060 ( .A(ein[680]), .B(n40652), .Z(ereg_next[681]) );
  AND U43061 ( .A(mul_pow), .B(n40653), .Z(n40652) );
  XOR U43062 ( .A(ein[681]), .B(ein[680]), .Z(n40653) );
  XOR U43063 ( .A(ein[679]), .B(n40654), .Z(ereg_next[680]) );
  AND U43064 ( .A(mul_pow), .B(n40655), .Z(n40654) );
  XOR U43065 ( .A(ein[680]), .B(ein[679]), .Z(n40655) );
  XOR U43066 ( .A(ein[66]), .B(n40656), .Z(ereg_next[67]) );
  AND U43067 ( .A(mul_pow), .B(n40657), .Z(n40656) );
  XOR U43068 ( .A(ein[67]), .B(ein[66]), .Z(n40657) );
  XOR U43069 ( .A(ein[678]), .B(n40658), .Z(ereg_next[679]) );
  AND U43070 ( .A(mul_pow), .B(n40659), .Z(n40658) );
  XOR U43071 ( .A(ein[679]), .B(ein[678]), .Z(n40659) );
  XOR U43072 ( .A(ein[677]), .B(n40660), .Z(ereg_next[678]) );
  AND U43073 ( .A(mul_pow), .B(n40661), .Z(n40660) );
  XOR U43074 ( .A(ein[678]), .B(ein[677]), .Z(n40661) );
  XOR U43075 ( .A(ein[676]), .B(n40662), .Z(ereg_next[677]) );
  AND U43076 ( .A(mul_pow), .B(n40663), .Z(n40662) );
  XOR U43077 ( .A(ein[677]), .B(ein[676]), .Z(n40663) );
  XOR U43078 ( .A(ein[675]), .B(n40664), .Z(ereg_next[676]) );
  AND U43079 ( .A(mul_pow), .B(n40665), .Z(n40664) );
  XOR U43080 ( .A(ein[676]), .B(ein[675]), .Z(n40665) );
  XOR U43081 ( .A(ein[674]), .B(n40666), .Z(ereg_next[675]) );
  AND U43082 ( .A(mul_pow), .B(n40667), .Z(n40666) );
  XOR U43083 ( .A(ein[675]), .B(ein[674]), .Z(n40667) );
  XOR U43084 ( .A(ein[673]), .B(n40668), .Z(ereg_next[674]) );
  AND U43085 ( .A(mul_pow), .B(n40669), .Z(n40668) );
  XOR U43086 ( .A(ein[674]), .B(ein[673]), .Z(n40669) );
  XOR U43087 ( .A(ein[672]), .B(n40670), .Z(ereg_next[673]) );
  AND U43088 ( .A(mul_pow), .B(n40671), .Z(n40670) );
  XOR U43089 ( .A(ein[673]), .B(ein[672]), .Z(n40671) );
  XOR U43090 ( .A(ein[671]), .B(n40672), .Z(ereg_next[672]) );
  AND U43091 ( .A(mul_pow), .B(n40673), .Z(n40672) );
  XOR U43092 ( .A(ein[672]), .B(ein[671]), .Z(n40673) );
  XOR U43093 ( .A(ein[670]), .B(n40674), .Z(ereg_next[671]) );
  AND U43094 ( .A(mul_pow), .B(n40675), .Z(n40674) );
  XOR U43095 ( .A(ein[671]), .B(ein[670]), .Z(n40675) );
  XOR U43096 ( .A(ein[669]), .B(n40676), .Z(ereg_next[670]) );
  AND U43097 ( .A(mul_pow), .B(n40677), .Z(n40676) );
  XOR U43098 ( .A(ein[670]), .B(ein[669]), .Z(n40677) );
  XOR U43099 ( .A(ein[65]), .B(n40678), .Z(ereg_next[66]) );
  AND U43100 ( .A(mul_pow), .B(n40679), .Z(n40678) );
  XOR U43101 ( .A(ein[66]), .B(ein[65]), .Z(n40679) );
  XOR U43102 ( .A(ein[668]), .B(n40680), .Z(ereg_next[669]) );
  AND U43103 ( .A(mul_pow), .B(n40681), .Z(n40680) );
  XOR U43104 ( .A(ein[669]), .B(ein[668]), .Z(n40681) );
  XOR U43105 ( .A(ein[667]), .B(n40682), .Z(ereg_next[668]) );
  AND U43106 ( .A(mul_pow), .B(n40683), .Z(n40682) );
  XOR U43107 ( .A(ein[668]), .B(ein[667]), .Z(n40683) );
  XOR U43108 ( .A(ein[666]), .B(n40684), .Z(ereg_next[667]) );
  AND U43109 ( .A(mul_pow), .B(n40685), .Z(n40684) );
  XOR U43110 ( .A(ein[667]), .B(ein[666]), .Z(n40685) );
  XOR U43111 ( .A(ein[665]), .B(n40686), .Z(ereg_next[666]) );
  AND U43112 ( .A(mul_pow), .B(n40687), .Z(n40686) );
  XOR U43113 ( .A(ein[666]), .B(ein[665]), .Z(n40687) );
  XOR U43114 ( .A(ein[664]), .B(n40688), .Z(ereg_next[665]) );
  AND U43115 ( .A(mul_pow), .B(n40689), .Z(n40688) );
  XOR U43116 ( .A(ein[665]), .B(ein[664]), .Z(n40689) );
  XOR U43117 ( .A(ein[663]), .B(n40690), .Z(ereg_next[664]) );
  AND U43118 ( .A(mul_pow), .B(n40691), .Z(n40690) );
  XOR U43119 ( .A(ein[664]), .B(ein[663]), .Z(n40691) );
  XOR U43120 ( .A(ein[662]), .B(n40692), .Z(ereg_next[663]) );
  AND U43121 ( .A(mul_pow), .B(n40693), .Z(n40692) );
  XOR U43122 ( .A(ein[663]), .B(ein[662]), .Z(n40693) );
  XOR U43123 ( .A(ein[661]), .B(n40694), .Z(ereg_next[662]) );
  AND U43124 ( .A(mul_pow), .B(n40695), .Z(n40694) );
  XOR U43125 ( .A(ein[662]), .B(ein[661]), .Z(n40695) );
  XOR U43126 ( .A(ein[660]), .B(n40696), .Z(ereg_next[661]) );
  AND U43127 ( .A(mul_pow), .B(n40697), .Z(n40696) );
  XOR U43128 ( .A(ein[661]), .B(ein[660]), .Z(n40697) );
  XOR U43129 ( .A(ein[659]), .B(n40698), .Z(ereg_next[660]) );
  AND U43130 ( .A(mul_pow), .B(n40699), .Z(n40698) );
  XOR U43131 ( .A(ein[660]), .B(ein[659]), .Z(n40699) );
  XOR U43132 ( .A(ein[64]), .B(n40700), .Z(ereg_next[65]) );
  AND U43133 ( .A(mul_pow), .B(n40701), .Z(n40700) );
  XOR U43134 ( .A(ein[65]), .B(ein[64]), .Z(n40701) );
  XOR U43135 ( .A(ein[658]), .B(n40702), .Z(ereg_next[659]) );
  AND U43136 ( .A(mul_pow), .B(n40703), .Z(n40702) );
  XOR U43137 ( .A(ein[659]), .B(ein[658]), .Z(n40703) );
  XOR U43138 ( .A(ein[657]), .B(n40704), .Z(ereg_next[658]) );
  AND U43139 ( .A(mul_pow), .B(n40705), .Z(n40704) );
  XOR U43140 ( .A(ein[658]), .B(ein[657]), .Z(n40705) );
  XOR U43141 ( .A(ein[656]), .B(n40706), .Z(ereg_next[657]) );
  AND U43142 ( .A(mul_pow), .B(n40707), .Z(n40706) );
  XOR U43143 ( .A(ein[657]), .B(ein[656]), .Z(n40707) );
  XOR U43144 ( .A(ein[655]), .B(n40708), .Z(ereg_next[656]) );
  AND U43145 ( .A(mul_pow), .B(n40709), .Z(n40708) );
  XOR U43146 ( .A(ein[656]), .B(ein[655]), .Z(n40709) );
  XOR U43147 ( .A(ein[654]), .B(n40710), .Z(ereg_next[655]) );
  AND U43148 ( .A(mul_pow), .B(n40711), .Z(n40710) );
  XOR U43149 ( .A(ein[655]), .B(ein[654]), .Z(n40711) );
  XOR U43150 ( .A(ein[653]), .B(n40712), .Z(ereg_next[654]) );
  AND U43151 ( .A(mul_pow), .B(n40713), .Z(n40712) );
  XOR U43152 ( .A(ein[654]), .B(ein[653]), .Z(n40713) );
  XOR U43153 ( .A(ein[652]), .B(n40714), .Z(ereg_next[653]) );
  AND U43154 ( .A(mul_pow), .B(n40715), .Z(n40714) );
  XOR U43155 ( .A(ein[653]), .B(ein[652]), .Z(n40715) );
  XOR U43156 ( .A(ein[651]), .B(n40716), .Z(ereg_next[652]) );
  AND U43157 ( .A(mul_pow), .B(n40717), .Z(n40716) );
  XOR U43158 ( .A(ein[652]), .B(ein[651]), .Z(n40717) );
  XOR U43159 ( .A(ein[650]), .B(n40718), .Z(ereg_next[651]) );
  AND U43160 ( .A(mul_pow), .B(n40719), .Z(n40718) );
  XOR U43161 ( .A(ein[651]), .B(ein[650]), .Z(n40719) );
  XOR U43162 ( .A(ein[649]), .B(n40720), .Z(ereg_next[650]) );
  AND U43163 ( .A(mul_pow), .B(n40721), .Z(n40720) );
  XOR U43164 ( .A(ein[650]), .B(ein[649]), .Z(n40721) );
  XOR U43165 ( .A(ein[63]), .B(n40722), .Z(ereg_next[64]) );
  AND U43166 ( .A(mul_pow), .B(n40723), .Z(n40722) );
  XOR U43167 ( .A(ein[64]), .B(ein[63]), .Z(n40723) );
  XOR U43168 ( .A(ein[648]), .B(n40724), .Z(ereg_next[649]) );
  AND U43169 ( .A(mul_pow), .B(n40725), .Z(n40724) );
  XOR U43170 ( .A(ein[649]), .B(ein[648]), .Z(n40725) );
  XOR U43171 ( .A(ein[647]), .B(n40726), .Z(ereg_next[648]) );
  AND U43172 ( .A(mul_pow), .B(n40727), .Z(n40726) );
  XOR U43173 ( .A(ein[648]), .B(ein[647]), .Z(n40727) );
  XOR U43174 ( .A(ein[646]), .B(n40728), .Z(ereg_next[647]) );
  AND U43175 ( .A(mul_pow), .B(n40729), .Z(n40728) );
  XOR U43176 ( .A(ein[647]), .B(ein[646]), .Z(n40729) );
  XOR U43177 ( .A(ein[645]), .B(n40730), .Z(ereg_next[646]) );
  AND U43178 ( .A(mul_pow), .B(n40731), .Z(n40730) );
  XOR U43179 ( .A(ein[646]), .B(ein[645]), .Z(n40731) );
  XOR U43180 ( .A(ein[644]), .B(n40732), .Z(ereg_next[645]) );
  AND U43181 ( .A(mul_pow), .B(n40733), .Z(n40732) );
  XOR U43182 ( .A(ein[645]), .B(ein[644]), .Z(n40733) );
  XOR U43183 ( .A(ein[643]), .B(n40734), .Z(ereg_next[644]) );
  AND U43184 ( .A(mul_pow), .B(n40735), .Z(n40734) );
  XOR U43185 ( .A(ein[644]), .B(ein[643]), .Z(n40735) );
  XOR U43186 ( .A(ein[642]), .B(n40736), .Z(ereg_next[643]) );
  AND U43187 ( .A(mul_pow), .B(n40737), .Z(n40736) );
  XOR U43188 ( .A(ein[643]), .B(ein[642]), .Z(n40737) );
  XOR U43189 ( .A(ein[641]), .B(n40738), .Z(ereg_next[642]) );
  AND U43190 ( .A(mul_pow), .B(n40739), .Z(n40738) );
  XOR U43191 ( .A(ein[642]), .B(ein[641]), .Z(n40739) );
  XOR U43192 ( .A(ein[640]), .B(n40740), .Z(ereg_next[641]) );
  AND U43193 ( .A(mul_pow), .B(n40741), .Z(n40740) );
  XOR U43194 ( .A(ein[641]), .B(ein[640]), .Z(n40741) );
  XOR U43195 ( .A(ein[639]), .B(n40742), .Z(ereg_next[640]) );
  AND U43196 ( .A(mul_pow), .B(n40743), .Z(n40742) );
  XOR U43197 ( .A(ein[640]), .B(ein[639]), .Z(n40743) );
  XOR U43198 ( .A(ein[62]), .B(n40744), .Z(ereg_next[63]) );
  AND U43199 ( .A(mul_pow), .B(n40745), .Z(n40744) );
  XOR U43200 ( .A(ein[63]), .B(ein[62]), .Z(n40745) );
  XOR U43201 ( .A(ein[638]), .B(n40746), .Z(ereg_next[639]) );
  AND U43202 ( .A(mul_pow), .B(n40747), .Z(n40746) );
  XOR U43203 ( .A(ein[639]), .B(ein[638]), .Z(n40747) );
  XOR U43204 ( .A(ein[637]), .B(n40748), .Z(ereg_next[638]) );
  AND U43205 ( .A(mul_pow), .B(n40749), .Z(n40748) );
  XOR U43206 ( .A(ein[638]), .B(ein[637]), .Z(n40749) );
  XOR U43207 ( .A(ein[636]), .B(n40750), .Z(ereg_next[637]) );
  AND U43208 ( .A(mul_pow), .B(n40751), .Z(n40750) );
  XOR U43209 ( .A(ein[637]), .B(ein[636]), .Z(n40751) );
  XOR U43210 ( .A(ein[635]), .B(n40752), .Z(ereg_next[636]) );
  AND U43211 ( .A(mul_pow), .B(n40753), .Z(n40752) );
  XOR U43212 ( .A(ein[636]), .B(ein[635]), .Z(n40753) );
  XOR U43213 ( .A(ein[634]), .B(n40754), .Z(ereg_next[635]) );
  AND U43214 ( .A(mul_pow), .B(n40755), .Z(n40754) );
  XOR U43215 ( .A(ein[635]), .B(ein[634]), .Z(n40755) );
  XOR U43216 ( .A(ein[633]), .B(n40756), .Z(ereg_next[634]) );
  AND U43217 ( .A(mul_pow), .B(n40757), .Z(n40756) );
  XOR U43218 ( .A(ein[634]), .B(ein[633]), .Z(n40757) );
  XOR U43219 ( .A(ein[632]), .B(n40758), .Z(ereg_next[633]) );
  AND U43220 ( .A(mul_pow), .B(n40759), .Z(n40758) );
  XOR U43221 ( .A(ein[633]), .B(ein[632]), .Z(n40759) );
  XOR U43222 ( .A(ein[631]), .B(n40760), .Z(ereg_next[632]) );
  AND U43223 ( .A(mul_pow), .B(n40761), .Z(n40760) );
  XOR U43224 ( .A(ein[632]), .B(ein[631]), .Z(n40761) );
  XOR U43225 ( .A(ein[630]), .B(n40762), .Z(ereg_next[631]) );
  AND U43226 ( .A(mul_pow), .B(n40763), .Z(n40762) );
  XOR U43227 ( .A(ein[631]), .B(ein[630]), .Z(n40763) );
  XOR U43228 ( .A(ein[629]), .B(n40764), .Z(ereg_next[630]) );
  AND U43229 ( .A(mul_pow), .B(n40765), .Z(n40764) );
  XOR U43230 ( .A(ein[630]), .B(ein[629]), .Z(n40765) );
  XOR U43231 ( .A(ein[61]), .B(n40766), .Z(ereg_next[62]) );
  AND U43232 ( .A(mul_pow), .B(n40767), .Z(n40766) );
  XOR U43233 ( .A(ein[62]), .B(ein[61]), .Z(n40767) );
  XOR U43234 ( .A(ein[628]), .B(n40768), .Z(ereg_next[629]) );
  AND U43235 ( .A(mul_pow), .B(n40769), .Z(n40768) );
  XOR U43236 ( .A(ein[629]), .B(ein[628]), .Z(n40769) );
  XOR U43237 ( .A(ein[627]), .B(n40770), .Z(ereg_next[628]) );
  AND U43238 ( .A(mul_pow), .B(n40771), .Z(n40770) );
  XOR U43239 ( .A(ein[628]), .B(ein[627]), .Z(n40771) );
  XOR U43240 ( .A(ein[626]), .B(n40772), .Z(ereg_next[627]) );
  AND U43241 ( .A(mul_pow), .B(n40773), .Z(n40772) );
  XOR U43242 ( .A(ein[627]), .B(ein[626]), .Z(n40773) );
  XOR U43243 ( .A(ein[625]), .B(n40774), .Z(ereg_next[626]) );
  AND U43244 ( .A(mul_pow), .B(n40775), .Z(n40774) );
  XOR U43245 ( .A(ein[626]), .B(ein[625]), .Z(n40775) );
  XOR U43246 ( .A(ein[624]), .B(n40776), .Z(ereg_next[625]) );
  AND U43247 ( .A(mul_pow), .B(n40777), .Z(n40776) );
  XOR U43248 ( .A(ein[625]), .B(ein[624]), .Z(n40777) );
  XOR U43249 ( .A(ein[623]), .B(n40778), .Z(ereg_next[624]) );
  AND U43250 ( .A(mul_pow), .B(n40779), .Z(n40778) );
  XOR U43251 ( .A(ein[624]), .B(ein[623]), .Z(n40779) );
  XOR U43252 ( .A(ein[622]), .B(n40780), .Z(ereg_next[623]) );
  AND U43253 ( .A(mul_pow), .B(n40781), .Z(n40780) );
  XOR U43254 ( .A(ein[623]), .B(ein[622]), .Z(n40781) );
  XOR U43255 ( .A(ein[621]), .B(n40782), .Z(ereg_next[622]) );
  AND U43256 ( .A(mul_pow), .B(n40783), .Z(n40782) );
  XOR U43257 ( .A(ein[622]), .B(ein[621]), .Z(n40783) );
  XOR U43258 ( .A(ein[620]), .B(n40784), .Z(ereg_next[621]) );
  AND U43259 ( .A(mul_pow), .B(n40785), .Z(n40784) );
  XOR U43260 ( .A(ein[621]), .B(ein[620]), .Z(n40785) );
  XOR U43261 ( .A(ein[619]), .B(n40786), .Z(ereg_next[620]) );
  AND U43262 ( .A(mul_pow), .B(n40787), .Z(n40786) );
  XOR U43263 ( .A(ein[620]), .B(ein[619]), .Z(n40787) );
  XOR U43264 ( .A(ein[60]), .B(n40788), .Z(ereg_next[61]) );
  AND U43265 ( .A(mul_pow), .B(n40789), .Z(n40788) );
  XOR U43266 ( .A(ein[61]), .B(ein[60]), .Z(n40789) );
  XOR U43267 ( .A(ein[618]), .B(n40790), .Z(ereg_next[619]) );
  AND U43268 ( .A(mul_pow), .B(n40791), .Z(n40790) );
  XOR U43269 ( .A(ein[619]), .B(ein[618]), .Z(n40791) );
  XOR U43270 ( .A(ein[617]), .B(n40792), .Z(ereg_next[618]) );
  AND U43271 ( .A(mul_pow), .B(n40793), .Z(n40792) );
  XOR U43272 ( .A(ein[618]), .B(ein[617]), .Z(n40793) );
  XOR U43273 ( .A(ein[616]), .B(n40794), .Z(ereg_next[617]) );
  AND U43274 ( .A(mul_pow), .B(n40795), .Z(n40794) );
  XOR U43275 ( .A(ein[617]), .B(ein[616]), .Z(n40795) );
  XOR U43276 ( .A(ein[615]), .B(n40796), .Z(ereg_next[616]) );
  AND U43277 ( .A(mul_pow), .B(n40797), .Z(n40796) );
  XOR U43278 ( .A(ein[616]), .B(ein[615]), .Z(n40797) );
  XOR U43279 ( .A(ein[614]), .B(n40798), .Z(ereg_next[615]) );
  AND U43280 ( .A(mul_pow), .B(n40799), .Z(n40798) );
  XOR U43281 ( .A(ein[615]), .B(ein[614]), .Z(n40799) );
  XOR U43282 ( .A(ein[613]), .B(n40800), .Z(ereg_next[614]) );
  AND U43283 ( .A(mul_pow), .B(n40801), .Z(n40800) );
  XOR U43284 ( .A(ein[614]), .B(ein[613]), .Z(n40801) );
  XOR U43285 ( .A(ein[612]), .B(n40802), .Z(ereg_next[613]) );
  AND U43286 ( .A(mul_pow), .B(n40803), .Z(n40802) );
  XOR U43287 ( .A(ein[613]), .B(ein[612]), .Z(n40803) );
  XOR U43288 ( .A(ein[611]), .B(n40804), .Z(ereg_next[612]) );
  AND U43289 ( .A(mul_pow), .B(n40805), .Z(n40804) );
  XOR U43290 ( .A(ein[612]), .B(ein[611]), .Z(n40805) );
  XOR U43291 ( .A(ein[610]), .B(n40806), .Z(ereg_next[611]) );
  AND U43292 ( .A(mul_pow), .B(n40807), .Z(n40806) );
  XOR U43293 ( .A(ein[611]), .B(ein[610]), .Z(n40807) );
  XOR U43294 ( .A(ein[609]), .B(n40808), .Z(ereg_next[610]) );
  AND U43295 ( .A(mul_pow), .B(n40809), .Z(n40808) );
  XOR U43296 ( .A(ein[610]), .B(ein[609]), .Z(n40809) );
  XOR U43297 ( .A(ein[59]), .B(n40810), .Z(ereg_next[60]) );
  AND U43298 ( .A(mul_pow), .B(n40811), .Z(n40810) );
  XOR U43299 ( .A(ein[60]), .B(ein[59]), .Z(n40811) );
  XOR U43300 ( .A(ein[608]), .B(n40812), .Z(ereg_next[609]) );
  AND U43301 ( .A(mul_pow), .B(n40813), .Z(n40812) );
  XOR U43302 ( .A(ein[609]), .B(ein[608]), .Z(n40813) );
  XOR U43303 ( .A(ein[607]), .B(n40814), .Z(ereg_next[608]) );
  AND U43304 ( .A(mul_pow), .B(n40815), .Z(n40814) );
  XOR U43305 ( .A(ein[608]), .B(ein[607]), .Z(n40815) );
  XOR U43306 ( .A(ein[606]), .B(n40816), .Z(ereg_next[607]) );
  AND U43307 ( .A(mul_pow), .B(n40817), .Z(n40816) );
  XOR U43308 ( .A(ein[607]), .B(ein[606]), .Z(n40817) );
  XOR U43309 ( .A(ein[605]), .B(n40818), .Z(ereg_next[606]) );
  AND U43310 ( .A(mul_pow), .B(n40819), .Z(n40818) );
  XOR U43311 ( .A(ein[606]), .B(ein[605]), .Z(n40819) );
  XOR U43312 ( .A(ein[604]), .B(n40820), .Z(ereg_next[605]) );
  AND U43313 ( .A(mul_pow), .B(n40821), .Z(n40820) );
  XOR U43314 ( .A(ein[605]), .B(ein[604]), .Z(n40821) );
  XOR U43315 ( .A(ein[603]), .B(n40822), .Z(ereg_next[604]) );
  AND U43316 ( .A(mul_pow), .B(n40823), .Z(n40822) );
  XOR U43317 ( .A(ein[604]), .B(ein[603]), .Z(n40823) );
  XOR U43318 ( .A(ein[602]), .B(n40824), .Z(ereg_next[603]) );
  AND U43319 ( .A(mul_pow), .B(n40825), .Z(n40824) );
  XOR U43320 ( .A(ein[603]), .B(ein[602]), .Z(n40825) );
  XOR U43321 ( .A(ein[601]), .B(n40826), .Z(ereg_next[602]) );
  AND U43322 ( .A(mul_pow), .B(n40827), .Z(n40826) );
  XOR U43323 ( .A(ein[602]), .B(ein[601]), .Z(n40827) );
  XOR U43324 ( .A(ein[600]), .B(n40828), .Z(ereg_next[601]) );
  AND U43325 ( .A(mul_pow), .B(n40829), .Z(n40828) );
  XOR U43326 ( .A(ein[601]), .B(ein[600]), .Z(n40829) );
  XOR U43327 ( .A(ein[599]), .B(n40830), .Z(ereg_next[600]) );
  AND U43328 ( .A(mul_pow), .B(n40831), .Z(n40830) );
  XOR U43329 ( .A(ein[600]), .B(ein[599]), .Z(n40831) );
  XOR U43330 ( .A(ein[4]), .B(n40832), .Z(ereg_next[5]) );
  AND U43331 ( .A(mul_pow), .B(n40833), .Z(n40832) );
  XOR U43332 ( .A(ein[5]), .B(ein[4]), .Z(n40833) );
  XOR U43333 ( .A(ein[58]), .B(n40834), .Z(ereg_next[59]) );
  AND U43334 ( .A(mul_pow), .B(n40835), .Z(n40834) );
  XOR U43335 ( .A(ein[59]), .B(ein[58]), .Z(n40835) );
  XOR U43336 ( .A(ein[598]), .B(n40836), .Z(ereg_next[599]) );
  AND U43337 ( .A(mul_pow), .B(n40837), .Z(n40836) );
  XOR U43338 ( .A(ein[599]), .B(ein[598]), .Z(n40837) );
  XOR U43339 ( .A(ein[597]), .B(n40838), .Z(ereg_next[598]) );
  AND U43340 ( .A(mul_pow), .B(n40839), .Z(n40838) );
  XOR U43341 ( .A(ein[598]), .B(ein[597]), .Z(n40839) );
  XOR U43342 ( .A(ein[596]), .B(n40840), .Z(ereg_next[597]) );
  AND U43343 ( .A(mul_pow), .B(n40841), .Z(n40840) );
  XOR U43344 ( .A(ein[597]), .B(ein[596]), .Z(n40841) );
  XOR U43345 ( .A(ein[595]), .B(n40842), .Z(ereg_next[596]) );
  AND U43346 ( .A(mul_pow), .B(n40843), .Z(n40842) );
  XOR U43347 ( .A(ein[596]), .B(ein[595]), .Z(n40843) );
  XOR U43348 ( .A(ein[594]), .B(n40844), .Z(ereg_next[595]) );
  AND U43349 ( .A(mul_pow), .B(n40845), .Z(n40844) );
  XOR U43350 ( .A(ein[595]), .B(ein[594]), .Z(n40845) );
  XOR U43351 ( .A(ein[593]), .B(n40846), .Z(ereg_next[594]) );
  AND U43352 ( .A(mul_pow), .B(n40847), .Z(n40846) );
  XOR U43353 ( .A(ein[594]), .B(ein[593]), .Z(n40847) );
  XOR U43354 ( .A(ein[592]), .B(n40848), .Z(ereg_next[593]) );
  AND U43355 ( .A(mul_pow), .B(n40849), .Z(n40848) );
  XOR U43356 ( .A(ein[593]), .B(ein[592]), .Z(n40849) );
  XOR U43357 ( .A(ein[591]), .B(n40850), .Z(ereg_next[592]) );
  AND U43358 ( .A(mul_pow), .B(n40851), .Z(n40850) );
  XOR U43359 ( .A(ein[592]), .B(ein[591]), .Z(n40851) );
  XOR U43360 ( .A(ein[590]), .B(n40852), .Z(ereg_next[591]) );
  AND U43361 ( .A(mul_pow), .B(n40853), .Z(n40852) );
  XOR U43362 ( .A(ein[591]), .B(ein[590]), .Z(n40853) );
  XOR U43363 ( .A(ein[589]), .B(n40854), .Z(ereg_next[590]) );
  AND U43364 ( .A(mul_pow), .B(n40855), .Z(n40854) );
  XOR U43365 ( .A(ein[590]), .B(ein[589]), .Z(n40855) );
  XOR U43366 ( .A(ein[57]), .B(n40856), .Z(ereg_next[58]) );
  AND U43367 ( .A(mul_pow), .B(n40857), .Z(n40856) );
  XOR U43368 ( .A(ein[58]), .B(ein[57]), .Z(n40857) );
  XOR U43369 ( .A(ein[588]), .B(n40858), .Z(ereg_next[589]) );
  AND U43370 ( .A(mul_pow), .B(n40859), .Z(n40858) );
  XOR U43371 ( .A(ein[589]), .B(ein[588]), .Z(n40859) );
  XOR U43372 ( .A(ein[587]), .B(n40860), .Z(ereg_next[588]) );
  AND U43373 ( .A(mul_pow), .B(n40861), .Z(n40860) );
  XOR U43374 ( .A(ein[588]), .B(ein[587]), .Z(n40861) );
  XOR U43375 ( .A(ein[586]), .B(n40862), .Z(ereg_next[587]) );
  AND U43376 ( .A(mul_pow), .B(n40863), .Z(n40862) );
  XOR U43377 ( .A(ein[587]), .B(ein[586]), .Z(n40863) );
  XOR U43378 ( .A(ein[585]), .B(n40864), .Z(ereg_next[586]) );
  AND U43379 ( .A(mul_pow), .B(n40865), .Z(n40864) );
  XOR U43380 ( .A(ein[586]), .B(ein[585]), .Z(n40865) );
  XOR U43381 ( .A(ein[584]), .B(n40866), .Z(ereg_next[585]) );
  AND U43382 ( .A(mul_pow), .B(n40867), .Z(n40866) );
  XOR U43383 ( .A(ein[585]), .B(ein[584]), .Z(n40867) );
  XOR U43384 ( .A(ein[583]), .B(n40868), .Z(ereg_next[584]) );
  AND U43385 ( .A(mul_pow), .B(n40869), .Z(n40868) );
  XOR U43386 ( .A(ein[584]), .B(ein[583]), .Z(n40869) );
  XOR U43387 ( .A(ein[582]), .B(n40870), .Z(ereg_next[583]) );
  AND U43388 ( .A(mul_pow), .B(n40871), .Z(n40870) );
  XOR U43389 ( .A(ein[583]), .B(ein[582]), .Z(n40871) );
  XOR U43390 ( .A(ein[581]), .B(n40872), .Z(ereg_next[582]) );
  AND U43391 ( .A(mul_pow), .B(n40873), .Z(n40872) );
  XOR U43392 ( .A(ein[582]), .B(ein[581]), .Z(n40873) );
  XOR U43393 ( .A(ein[580]), .B(n40874), .Z(ereg_next[581]) );
  AND U43394 ( .A(mul_pow), .B(n40875), .Z(n40874) );
  XOR U43395 ( .A(ein[581]), .B(ein[580]), .Z(n40875) );
  XOR U43396 ( .A(ein[579]), .B(n40876), .Z(ereg_next[580]) );
  AND U43397 ( .A(mul_pow), .B(n40877), .Z(n40876) );
  XOR U43398 ( .A(ein[580]), .B(ein[579]), .Z(n40877) );
  XOR U43399 ( .A(ein[56]), .B(n40878), .Z(ereg_next[57]) );
  AND U43400 ( .A(mul_pow), .B(n40879), .Z(n40878) );
  XOR U43401 ( .A(ein[57]), .B(ein[56]), .Z(n40879) );
  XOR U43402 ( .A(ein[578]), .B(n40880), .Z(ereg_next[579]) );
  AND U43403 ( .A(mul_pow), .B(n40881), .Z(n40880) );
  XOR U43404 ( .A(ein[579]), .B(ein[578]), .Z(n40881) );
  XOR U43405 ( .A(ein[577]), .B(n40882), .Z(ereg_next[578]) );
  AND U43406 ( .A(mul_pow), .B(n40883), .Z(n40882) );
  XOR U43407 ( .A(ein[578]), .B(ein[577]), .Z(n40883) );
  XOR U43408 ( .A(ein[576]), .B(n40884), .Z(ereg_next[577]) );
  AND U43409 ( .A(mul_pow), .B(n40885), .Z(n40884) );
  XOR U43410 ( .A(ein[577]), .B(ein[576]), .Z(n40885) );
  XOR U43411 ( .A(ein[575]), .B(n40886), .Z(ereg_next[576]) );
  AND U43412 ( .A(mul_pow), .B(n40887), .Z(n40886) );
  XOR U43413 ( .A(ein[576]), .B(ein[575]), .Z(n40887) );
  XOR U43414 ( .A(ein[574]), .B(n40888), .Z(ereg_next[575]) );
  AND U43415 ( .A(mul_pow), .B(n40889), .Z(n40888) );
  XOR U43416 ( .A(ein[575]), .B(ein[574]), .Z(n40889) );
  XOR U43417 ( .A(ein[573]), .B(n40890), .Z(ereg_next[574]) );
  AND U43418 ( .A(mul_pow), .B(n40891), .Z(n40890) );
  XOR U43419 ( .A(ein[574]), .B(ein[573]), .Z(n40891) );
  XOR U43420 ( .A(ein[572]), .B(n40892), .Z(ereg_next[573]) );
  AND U43421 ( .A(mul_pow), .B(n40893), .Z(n40892) );
  XOR U43422 ( .A(ein[573]), .B(ein[572]), .Z(n40893) );
  XOR U43423 ( .A(ein[571]), .B(n40894), .Z(ereg_next[572]) );
  AND U43424 ( .A(mul_pow), .B(n40895), .Z(n40894) );
  XOR U43425 ( .A(ein[572]), .B(ein[571]), .Z(n40895) );
  XOR U43426 ( .A(ein[570]), .B(n40896), .Z(ereg_next[571]) );
  AND U43427 ( .A(mul_pow), .B(n40897), .Z(n40896) );
  XOR U43428 ( .A(ein[571]), .B(ein[570]), .Z(n40897) );
  XOR U43429 ( .A(ein[569]), .B(n40898), .Z(ereg_next[570]) );
  AND U43430 ( .A(mul_pow), .B(n40899), .Z(n40898) );
  XOR U43431 ( .A(ein[570]), .B(ein[569]), .Z(n40899) );
  XOR U43432 ( .A(ein[55]), .B(n40900), .Z(ereg_next[56]) );
  AND U43433 ( .A(mul_pow), .B(n40901), .Z(n40900) );
  XOR U43434 ( .A(ein[56]), .B(ein[55]), .Z(n40901) );
  XOR U43435 ( .A(ein[568]), .B(n40902), .Z(ereg_next[569]) );
  AND U43436 ( .A(mul_pow), .B(n40903), .Z(n40902) );
  XOR U43437 ( .A(ein[569]), .B(ein[568]), .Z(n40903) );
  XOR U43438 ( .A(ein[567]), .B(n40904), .Z(ereg_next[568]) );
  AND U43439 ( .A(mul_pow), .B(n40905), .Z(n40904) );
  XOR U43440 ( .A(ein[568]), .B(ein[567]), .Z(n40905) );
  XOR U43441 ( .A(ein[566]), .B(n40906), .Z(ereg_next[567]) );
  AND U43442 ( .A(mul_pow), .B(n40907), .Z(n40906) );
  XOR U43443 ( .A(ein[567]), .B(ein[566]), .Z(n40907) );
  XOR U43444 ( .A(ein[565]), .B(n40908), .Z(ereg_next[566]) );
  AND U43445 ( .A(mul_pow), .B(n40909), .Z(n40908) );
  XOR U43446 ( .A(ein[566]), .B(ein[565]), .Z(n40909) );
  XOR U43447 ( .A(ein[564]), .B(n40910), .Z(ereg_next[565]) );
  AND U43448 ( .A(mul_pow), .B(n40911), .Z(n40910) );
  XOR U43449 ( .A(ein[565]), .B(ein[564]), .Z(n40911) );
  XOR U43450 ( .A(ein[563]), .B(n40912), .Z(ereg_next[564]) );
  AND U43451 ( .A(mul_pow), .B(n40913), .Z(n40912) );
  XOR U43452 ( .A(ein[564]), .B(ein[563]), .Z(n40913) );
  XOR U43453 ( .A(ein[562]), .B(n40914), .Z(ereg_next[563]) );
  AND U43454 ( .A(mul_pow), .B(n40915), .Z(n40914) );
  XOR U43455 ( .A(ein[563]), .B(ein[562]), .Z(n40915) );
  XOR U43456 ( .A(ein[561]), .B(n40916), .Z(ereg_next[562]) );
  AND U43457 ( .A(mul_pow), .B(n40917), .Z(n40916) );
  XOR U43458 ( .A(ein[562]), .B(ein[561]), .Z(n40917) );
  XOR U43459 ( .A(ein[560]), .B(n40918), .Z(ereg_next[561]) );
  AND U43460 ( .A(mul_pow), .B(n40919), .Z(n40918) );
  XOR U43461 ( .A(ein[561]), .B(ein[560]), .Z(n40919) );
  XOR U43462 ( .A(ein[559]), .B(n40920), .Z(ereg_next[560]) );
  AND U43463 ( .A(mul_pow), .B(n40921), .Z(n40920) );
  XOR U43464 ( .A(ein[560]), .B(ein[559]), .Z(n40921) );
  XOR U43465 ( .A(ein[54]), .B(n40922), .Z(ereg_next[55]) );
  AND U43466 ( .A(mul_pow), .B(n40923), .Z(n40922) );
  XOR U43467 ( .A(ein[55]), .B(ein[54]), .Z(n40923) );
  XOR U43468 ( .A(ein[558]), .B(n40924), .Z(ereg_next[559]) );
  AND U43469 ( .A(mul_pow), .B(n40925), .Z(n40924) );
  XOR U43470 ( .A(ein[559]), .B(ein[558]), .Z(n40925) );
  XOR U43471 ( .A(ein[557]), .B(n40926), .Z(ereg_next[558]) );
  AND U43472 ( .A(mul_pow), .B(n40927), .Z(n40926) );
  XOR U43473 ( .A(ein[558]), .B(ein[557]), .Z(n40927) );
  XOR U43474 ( .A(ein[556]), .B(n40928), .Z(ereg_next[557]) );
  AND U43475 ( .A(mul_pow), .B(n40929), .Z(n40928) );
  XOR U43476 ( .A(ein[557]), .B(ein[556]), .Z(n40929) );
  XOR U43477 ( .A(ein[555]), .B(n40930), .Z(ereg_next[556]) );
  AND U43478 ( .A(mul_pow), .B(n40931), .Z(n40930) );
  XOR U43479 ( .A(ein[556]), .B(ein[555]), .Z(n40931) );
  XOR U43480 ( .A(ein[554]), .B(n40932), .Z(ereg_next[555]) );
  AND U43481 ( .A(mul_pow), .B(n40933), .Z(n40932) );
  XOR U43482 ( .A(ein[555]), .B(ein[554]), .Z(n40933) );
  XOR U43483 ( .A(ein[553]), .B(n40934), .Z(ereg_next[554]) );
  AND U43484 ( .A(mul_pow), .B(n40935), .Z(n40934) );
  XOR U43485 ( .A(ein[554]), .B(ein[553]), .Z(n40935) );
  XOR U43486 ( .A(ein[552]), .B(n40936), .Z(ereg_next[553]) );
  AND U43487 ( .A(mul_pow), .B(n40937), .Z(n40936) );
  XOR U43488 ( .A(ein[553]), .B(ein[552]), .Z(n40937) );
  XOR U43489 ( .A(ein[551]), .B(n40938), .Z(ereg_next[552]) );
  AND U43490 ( .A(mul_pow), .B(n40939), .Z(n40938) );
  XOR U43491 ( .A(ein[552]), .B(ein[551]), .Z(n40939) );
  XOR U43492 ( .A(ein[550]), .B(n40940), .Z(ereg_next[551]) );
  AND U43493 ( .A(mul_pow), .B(n40941), .Z(n40940) );
  XOR U43494 ( .A(ein[551]), .B(ein[550]), .Z(n40941) );
  XOR U43495 ( .A(ein[549]), .B(n40942), .Z(ereg_next[550]) );
  AND U43496 ( .A(mul_pow), .B(n40943), .Z(n40942) );
  XOR U43497 ( .A(ein[550]), .B(ein[549]), .Z(n40943) );
  XOR U43498 ( .A(ein[53]), .B(n40944), .Z(ereg_next[54]) );
  AND U43499 ( .A(mul_pow), .B(n40945), .Z(n40944) );
  XOR U43500 ( .A(ein[54]), .B(ein[53]), .Z(n40945) );
  XOR U43501 ( .A(ein[548]), .B(n40946), .Z(ereg_next[549]) );
  AND U43502 ( .A(mul_pow), .B(n40947), .Z(n40946) );
  XOR U43503 ( .A(ein[549]), .B(ein[548]), .Z(n40947) );
  XOR U43504 ( .A(ein[547]), .B(n40948), .Z(ereg_next[548]) );
  AND U43505 ( .A(mul_pow), .B(n40949), .Z(n40948) );
  XOR U43506 ( .A(ein[548]), .B(ein[547]), .Z(n40949) );
  XOR U43507 ( .A(ein[546]), .B(n40950), .Z(ereg_next[547]) );
  AND U43508 ( .A(mul_pow), .B(n40951), .Z(n40950) );
  XOR U43509 ( .A(ein[547]), .B(ein[546]), .Z(n40951) );
  XOR U43510 ( .A(ein[545]), .B(n40952), .Z(ereg_next[546]) );
  AND U43511 ( .A(mul_pow), .B(n40953), .Z(n40952) );
  XOR U43512 ( .A(ein[546]), .B(ein[545]), .Z(n40953) );
  XOR U43513 ( .A(ein[544]), .B(n40954), .Z(ereg_next[545]) );
  AND U43514 ( .A(mul_pow), .B(n40955), .Z(n40954) );
  XOR U43515 ( .A(ein[545]), .B(ein[544]), .Z(n40955) );
  XOR U43516 ( .A(ein[543]), .B(n40956), .Z(ereg_next[544]) );
  AND U43517 ( .A(mul_pow), .B(n40957), .Z(n40956) );
  XOR U43518 ( .A(ein[544]), .B(ein[543]), .Z(n40957) );
  XOR U43519 ( .A(ein[542]), .B(n40958), .Z(ereg_next[543]) );
  AND U43520 ( .A(mul_pow), .B(n40959), .Z(n40958) );
  XOR U43521 ( .A(ein[543]), .B(ein[542]), .Z(n40959) );
  XOR U43522 ( .A(ein[541]), .B(n40960), .Z(ereg_next[542]) );
  AND U43523 ( .A(mul_pow), .B(n40961), .Z(n40960) );
  XOR U43524 ( .A(ein[542]), .B(ein[541]), .Z(n40961) );
  XOR U43525 ( .A(ein[540]), .B(n40962), .Z(ereg_next[541]) );
  AND U43526 ( .A(mul_pow), .B(n40963), .Z(n40962) );
  XOR U43527 ( .A(ein[541]), .B(ein[540]), .Z(n40963) );
  XOR U43528 ( .A(ein[539]), .B(n40964), .Z(ereg_next[540]) );
  AND U43529 ( .A(mul_pow), .B(n40965), .Z(n40964) );
  XOR U43530 ( .A(ein[540]), .B(ein[539]), .Z(n40965) );
  XOR U43531 ( .A(ein[52]), .B(n40966), .Z(ereg_next[53]) );
  AND U43532 ( .A(mul_pow), .B(n40967), .Z(n40966) );
  XOR U43533 ( .A(ein[53]), .B(ein[52]), .Z(n40967) );
  XOR U43534 ( .A(ein[538]), .B(n40968), .Z(ereg_next[539]) );
  AND U43535 ( .A(mul_pow), .B(n40969), .Z(n40968) );
  XOR U43536 ( .A(ein[539]), .B(ein[538]), .Z(n40969) );
  XOR U43537 ( .A(ein[537]), .B(n40970), .Z(ereg_next[538]) );
  AND U43538 ( .A(mul_pow), .B(n40971), .Z(n40970) );
  XOR U43539 ( .A(ein[538]), .B(ein[537]), .Z(n40971) );
  XOR U43540 ( .A(ein[536]), .B(n40972), .Z(ereg_next[537]) );
  AND U43541 ( .A(mul_pow), .B(n40973), .Z(n40972) );
  XOR U43542 ( .A(ein[537]), .B(ein[536]), .Z(n40973) );
  XOR U43543 ( .A(ein[535]), .B(n40974), .Z(ereg_next[536]) );
  AND U43544 ( .A(mul_pow), .B(n40975), .Z(n40974) );
  XOR U43545 ( .A(ein[536]), .B(ein[535]), .Z(n40975) );
  XOR U43546 ( .A(ein[534]), .B(n40976), .Z(ereg_next[535]) );
  AND U43547 ( .A(mul_pow), .B(n40977), .Z(n40976) );
  XOR U43548 ( .A(ein[535]), .B(ein[534]), .Z(n40977) );
  XOR U43549 ( .A(ein[533]), .B(n40978), .Z(ereg_next[534]) );
  AND U43550 ( .A(mul_pow), .B(n40979), .Z(n40978) );
  XOR U43551 ( .A(ein[534]), .B(ein[533]), .Z(n40979) );
  XOR U43552 ( .A(ein[532]), .B(n40980), .Z(ereg_next[533]) );
  AND U43553 ( .A(mul_pow), .B(n40981), .Z(n40980) );
  XOR U43554 ( .A(ein[533]), .B(ein[532]), .Z(n40981) );
  XOR U43555 ( .A(ein[531]), .B(n40982), .Z(ereg_next[532]) );
  AND U43556 ( .A(mul_pow), .B(n40983), .Z(n40982) );
  XOR U43557 ( .A(ein[532]), .B(ein[531]), .Z(n40983) );
  XOR U43558 ( .A(ein[530]), .B(n40984), .Z(ereg_next[531]) );
  AND U43559 ( .A(mul_pow), .B(n40985), .Z(n40984) );
  XOR U43560 ( .A(ein[531]), .B(ein[530]), .Z(n40985) );
  XOR U43561 ( .A(ein[529]), .B(n40986), .Z(ereg_next[530]) );
  AND U43562 ( .A(mul_pow), .B(n40987), .Z(n40986) );
  XOR U43563 ( .A(ein[530]), .B(ein[529]), .Z(n40987) );
  XOR U43564 ( .A(ein[51]), .B(n40988), .Z(ereg_next[52]) );
  AND U43565 ( .A(mul_pow), .B(n40989), .Z(n40988) );
  XOR U43566 ( .A(ein[52]), .B(ein[51]), .Z(n40989) );
  XOR U43567 ( .A(ein[528]), .B(n40990), .Z(ereg_next[529]) );
  AND U43568 ( .A(mul_pow), .B(n40991), .Z(n40990) );
  XOR U43569 ( .A(ein[529]), .B(ein[528]), .Z(n40991) );
  XOR U43570 ( .A(ein[527]), .B(n40992), .Z(ereg_next[528]) );
  AND U43571 ( .A(mul_pow), .B(n40993), .Z(n40992) );
  XOR U43572 ( .A(ein[528]), .B(ein[527]), .Z(n40993) );
  XOR U43573 ( .A(ein[526]), .B(n40994), .Z(ereg_next[527]) );
  AND U43574 ( .A(mul_pow), .B(n40995), .Z(n40994) );
  XOR U43575 ( .A(ein[527]), .B(ein[526]), .Z(n40995) );
  XOR U43576 ( .A(ein[525]), .B(n40996), .Z(ereg_next[526]) );
  AND U43577 ( .A(mul_pow), .B(n40997), .Z(n40996) );
  XOR U43578 ( .A(ein[526]), .B(ein[525]), .Z(n40997) );
  XOR U43579 ( .A(ein[524]), .B(n40998), .Z(ereg_next[525]) );
  AND U43580 ( .A(mul_pow), .B(n40999), .Z(n40998) );
  XOR U43581 ( .A(ein[525]), .B(ein[524]), .Z(n40999) );
  XOR U43582 ( .A(ein[523]), .B(n41000), .Z(ereg_next[524]) );
  AND U43583 ( .A(mul_pow), .B(n41001), .Z(n41000) );
  XOR U43584 ( .A(ein[524]), .B(ein[523]), .Z(n41001) );
  XOR U43585 ( .A(ein[522]), .B(n41002), .Z(ereg_next[523]) );
  AND U43586 ( .A(mul_pow), .B(n41003), .Z(n41002) );
  XOR U43587 ( .A(ein[523]), .B(ein[522]), .Z(n41003) );
  XOR U43588 ( .A(ein[521]), .B(n41004), .Z(ereg_next[522]) );
  AND U43589 ( .A(mul_pow), .B(n41005), .Z(n41004) );
  XOR U43590 ( .A(ein[522]), .B(ein[521]), .Z(n41005) );
  XOR U43591 ( .A(ein[520]), .B(n41006), .Z(ereg_next[521]) );
  AND U43592 ( .A(mul_pow), .B(n41007), .Z(n41006) );
  XOR U43593 ( .A(ein[521]), .B(ein[520]), .Z(n41007) );
  XOR U43594 ( .A(ein[519]), .B(n41008), .Z(ereg_next[520]) );
  AND U43595 ( .A(mul_pow), .B(n41009), .Z(n41008) );
  XOR U43596 ( .A(ein[520]), .B(ein[519]), .Z(n41009) );
  XOR U43597 ( .A(ein[50]), .B(n41010), .Z(ereg_next[51]) );
  AND U43598 ( .A(mul_pow), .B(n41011), .Z(n41010) );
  XOR U43599 ( .A(ein[51]), .B(ein[50]), .Z(n41011) );
  XOR U43600 ( .A(ein[518]), .B(n41012), .Z(ereg_next[519]) );
  AND U43601 ( .A(mul_pow), .B(n41013), .Z(n41012) );
  XOR U43602 ( .A(ein[519]), .B(ein[518]), .Z(n41013) );
  XOR U43603 ( .A(ein[517]), .B(n41014), .Z(ereg_next[518]) );
  AND U43604 ( .A(mul_pow), .B(n41015), .Z(n41014) );
  XOR U43605 ( .A(ein[518]), .B(ein[517]), .Z(n41015) );
  XOR U43606 ( .A(ein[516]), .B(n41016), .Z(ereg_next[517]) );
  AND U43607 ( .A(mul_pow), .B(n41017), .Z(n41016) );
  XOR U43608 ( .A(ein[517]), .B(ein[516]), .Z(n41017) );
  XOR U43609 ( .A(ein[515]), .B(n41018), .Z(ereg_next[516]) );
  AND U43610 ( .A(mul_pow), .B(n41019), .Z(n41018) );
  XOR U43611 ( .A(ein[516]), .B(ein[515]), .Z(n41019) );
  XOR U43612 ( .A(ein[514]), .B(n41020), .Z(ereg_next[515]) );
  AND U43613 ( .A(mul_pow), .B(n41021), .Z(n41020) );
  XOR U43614 ( .A(ein[515]), .B(ein[514]), .Z(n41021) );
  XOR U43615 ( .A(ein[513]), .B(n41022), .Z(ereg_next[514]) );
  AND U43616 ( .A(mul_pow), .B(n41023), .Z(n41022) );
  XOR U43617 ( .A(ein[514]), .B(ein[513]), .Z(n41023) );
  XOR U43618 ( .A(ein[512]), .B(n41024), .Z(ereg_next[513]) );
  AND U43619 ( .A(mul_pow), .B(n41025), .Z(n41024) );
  XOR U43620 ( .A(ein[513]), .B(ein[512]), .Z(n41025) );
  XOR U43621 ( .A(ein[511]), .B(n41026), .Z(ereg_next[512]) );
  AND U43622 ( .A(mul_pow), .B(n41027), .Z(n41026) );
  XOR U43623 ( .A(ein[512]), .B(ein[511]), .Z(n41027) );
  XOR U43624 ( .A(ein[510]), .B(n41028), .Z(ereg_next[511]) );
  AND U43625 ( .A(mul_pow), .B(n41029), .Z(n41028) );
  XOR U43626 ( .A(ein[511]), .B(ein[510]), .Z(n41029) );
  XOR U43627 ( .A(ein[509]), .B(n41030), .Z(ereg_next[510]) );
  AND U43628 ( .A(mul_pow), .B(n41031), .Z(n41030) );
  XOR U43629 ( .A(ein[510]), .B(ein[509]), .Z(n41031) );
  XOR U43630 ( .A(ein[49]), .B(n41032), .Z(ereg_next[50]) );
  AND U43631 ( .A(mul_pow), .B(n41033), .Z(n41032) );
  XOR U43632 ( .A(ein[50]), .B(ein[49]), .Z(n41033) );
  XOR U43633 ( .A(ein[508]), .B(n41034), .Z(ereg_next[509]) );
  AND U43634 ( .A(mul_pow), .B(n41035), .Z(n41034) );
  XOR U43635 ( .A(ein[509]), .B(ein[508]), .Z(n41035) );
  XOR U43636 ( .A(ein[507]), .B(n41036), .Z(ereg_next[508]) );
  AND U43637 ( .A(mul_pow), .B(n41037), .Z(n41036) );
  XOR U43638 ( .A(ein[508]), .B(ein[507]), .Z(n41037) );
  XOR U43639 ( .A(ein[506]), .B(n41038), .Z(ereg_next[507]) );
  AND U43640 ( .A(mul_pow), .B(n41039), .Z(n41038) );
  XOR U43641 ( .A(ein[507]), .B(ein[506]), .Z(n41039) );
  XOR U43642 ( .A(ein[505]), .B(n41040), .Z(ereg_next[506]) );
  AND U43643 ( .A(mul_pow), .B(n41041), .Z(n41040) );
  XOR U43644 ( .A(ein[506]), .B(ein[505]), .Z(n41041) );
  XOR U43645 ( .A(ein[504]), .B(n41042), .Z(ereg_next[505]) );
  AND U43646 ( .A(mul_pow), .B(n41043), .Z(n41042) );
  XOR U43647 ( .A(ein[505]), .B(ein[504]), .Z(n41043) );
  XOR U43648 ( .A(ein[503]), .B(n41044), .Z(ereg_next[504]) );
  AND U43649 ( .A(mul_pow), .B(n41045), .Z(n41044) );
  XOR U43650 ( .A(ein[504]), .B(ein[503]), .Z(n41045) );
  XOR U43651 ( .A(ein[502]), .B(n41046), .Z(ereg_next[503]) );
  AND U43652 ( .A(mul_pow), .B(n41047), .Z(n41046) );
  XOR U43653 ( .A(ein[503]), .B(ein[502]), .Z(n41047) );
  XOR U43654 ( .A(ein[501]), .B(n41048), .Z(ereg_next[502]) );
  AND U43655 ( .A(mul_pow), .B(n41049), .Z(n41048) );
  XOR U43656 ( .A(ein[502]), .B(ein[501]), .Z(n41049) );
  XOR U43657 ( .A(ein[500]), .B(n41050), .Z(ereg_next[501]) );
  AND U43658 ( .A(mul_pow), .B(n41051), .Z(n41050) );
  XOR U43659 ( .A(ein[501]), .B(ein[500]), .Z(n41051) );
  XOR U43660 ( .A(ein[499]), .B(n41052), .Z(ereg_next[500]) );
  AND U43661 ( .A(mul_pow), .B(n41053), .Z(n41052) );
  XOR U43662 ( .A(ein[500]), .B(ein[499]), .Z(n41053) );
  XOR U43663 ( .A(ein[3]), .B(n41054), .Z(ereg_next[4]) );
  AND U43664 ( .A(mul_pow), .B(n41055), .Z(n41054) );
  XOR U43665 ( .A(ein[4]), .B(ein[3]), .Z(n41055) );
  XOR U43666 ( .A(ein[48]), .B(n41056), .Z(ereg_next[49]) );
  AND U43667 ( .A(mul_pow), .B(n41057), .Z(n41056) );
  XOR U43668 ( .A(ein[49]), .B(ein[48]), .Z(n41057) );
  XOR U43669 ( .A(ein[498]), .B(n41058), .Z(ereg_next[499]) );
  AND U43670 ( .A(mul_pow), .B(n41059), .Z(n41058) );
  XOR U43671 ( .A(ein[499]), .B(ein[498]), .Z(n41059) );
  XOR U43672 ( .A(ein[497]), .B(n41060), .Z(ereg_next[498]) );
  AND U43673 ( .A(mul_pow), .B(n41061), .Z(n41060) );
  XOR U43674 ( .A(ein[498]), .B(ein[497]), .Z(n41061) );
  XOR U43675 ( .A(ein[496]), .B(n41062), .Z(ereg_next[497]) );
  AND U43676 ( .A(mul_pow), .B(n41063), .Z(n41062) );
  XOR U43677 ( .A(ein[497]), .B(ein[496]), .Z(n41063) );
  XOR U43678 ( .A(ein[495]), .B(n41064), .Z(ereg_next[496]) );
  AND U43679 ( .A(mul_pow), .B(n41065), .Z(n41064) );
  XOR U43680 ( .A(ein[496]), .B(ein[495]), .Z(n41065) );
  XOR U43681 ( .A(ein[494]), .B(n41066), .Z(ereg_next[495]) );
  AND U43682 ( .A(mul_pow), .B(n41067), .Z(n41066) );
  XOR U43683 ( .A(ein[495]), .B(ein[494]), .Z(n41067) );
  XOR U43684 ( .A(ein[493]), .B(n41068), .Z(ereg_next[494]) );
  AND U43685 ( .A(mul_pow), .B(n41069), .Z(n41068) );
  XOR U43686 ( .A(ein[494]), .B(ein[493]), .Z(n41069) );
  XOR U43687 ( .A(ein[492]), .B(n41070), .Z(ereg_next[493]) );
  AND U43688 ( .A(mul_pow), .B(n41071), .Z(n41070) );
  XOR U43689 ( .A(ein[493]), .B(ein[492]), .Z(n41071) );
  XOR U43690 ( .A(ein[491]), .B(n41072), .Z(ereg_next[492]) );
  AND U43691 ( .A(mul_pow), .B(n41073), .Z(n41072) );
  XOR U43692 ( .A(ein[492]), .B(ein[491]), .Z(n41073) );
  XOR U43693 ( .A(ein[490]), .B(n41074), .Z(ereg_next[491]) );
  AND U43694 ( .A(mul_pow), .B(n41075), .Z(n41074) );
  XOR U43695 ( .A(ein[491]), .B(ein[490]), .Z(n41075) );
  XOR U43696 ( .A(ein[489]), .B(n41076), .Z(ereg_next[490]) );
  AND U43697 ( .A(mul_pow), .B(n41077), .Z(n41076) );
  XOR U43698 ( .A(ein[490]), .B(ein[489]), .Z(n41077) );
  XOR U43699 ( .A(ein[47]), .B(n41078), .Z(ereg_next[48]) );
  AND U43700 ( .A(mul_pow), .B(n41079), .Z(n41078) );
  XOR U43701 ( .A(ein[48]), .B(ein[47]), .Z(n41079) );
  XOR U43702 ( .A(ein[488]), .B(n41080), .Z(ereg_next[489]) );
  AND U43703 ( .A(mul_pow), .B(n41081), .Z(n41080) );
  XOR U43704 ( .A(ein[489]), .B(ein[488]), .Z(n41081) );
  XOR U43705 ( .A(ein[487]), .B(n41082), .Z(ereg_next[488]) );
  AND U43706 ( .A(mul_pow), .B(n41083), .Z(n41082) );
  XOR U43707 ( .A(ein[488]), .B(ein[487]), .Z(n41083) );
  XOR U43708 ( .A(ein[486]), .B(n41084), .Z(ereg_next[487]) );
  AND U43709 ( .A(mul_pow), .B(n41085), .Z(n41084) );
  XOR U43710 ( .A(ein[487]), .B(ein[486]), .Z(n41085) );
  XOR U43711 ( .A(ein[485]), .B(n41086), .Z(ereg_next[486]) );
  AND U43712 ( .A(mul_pow), .B(n41087), .Z(n41086) );
  XOR U43713 ( .A(ein[486]), .B(ein[485]), .Z(n41087) );
  XOR U43714 ( .A(ein[484]), .B(n41088), .Z(ereg_next[485]) );
  AND U43715 ( .A(mul_pow), .B(n41089), .Z(n41088) );
  XOR U43716 ( .A(ein[485]), .B(ein[484]), .Z(n41089) );
  XOR U43717 ( .A(ein[483]), .B(n41090), .Z(ereg_next[484]) );
  AND U43718 ( .A(mul_pow), .B(n41091), .Z(n41090) );
  XOR U43719 ( .A(ein[484]), .B(ein[483]), .Z(n41091) );
  XOR U43720 ( .A(ein[482]), .B(n41092), .Z(ereg_next[483]) );
  AND U43721 ( .A(mul_pow), .B(n41093), .Z(n41092) );
  XOR U43722 ( .A(ein[483]), .B(ein[482]), .Z(n41093) );
  XOR U43723 ( .A(ein[481]), .B(n41094), .Z(ereg_next[482]) );
  AND U43724 ( .A(mul_pow), .B(n41095), .Z(n41094) );
  XOR U43725 ( .A(ein[482]), .B(ein[481]), .Z(n41095) );
  XOR U43726 ( .A(ein[480]), .B(n41096), .Z(ereg_next[481]) );
  AND U43727 ( .A(mul_pow), .B(n41097), .Z(n41096) );
  XOR U43728 ( .A(ein[481]), .B(ein[480]), .Z(n41097) );
  XOR U43729 ( .A(ein[479]), .B(n41098), .Z(ereg_next[480]) );
  AND U43730 ( .A(mul_pow), .B(n41099), .Z(n41098) );
  XOR U43731 ( .A(ein[480]), .B(ein[479]), .Z(n41099) );
  XOR U43732 ( .A(ein[46]), .B(n41100), .Z(ereg_next[47]) );
  AND U43733 ( .A(mul_pow), .B(n41101), .Z(n41100) );
  XOR U43734 ( .A(ein[47]), .B(ein[46]), .Z(n41101) );
  XOR U43735 ( .A(ein[478]), .B(n41102), .Z(ereg_next[479]) );
  AND U43736 ( .A(mul_pow), .B(n41103), .Z(n41102) );
  XOR U43737 ( .A(ein[479]), .B(ein[478]), .Z(n41103) );
  XOR U43738 ( .A(ein[477]), .B(n41104), .Z(ereg_next[478]) );
  AND U43739 ( .A(mul_pow), .B(n41105), .Z(n41104) );
  XOR U43740 ( .A(ein[478]), .B(ein[477]), .Z(n41105) );
  XOR U43741 ( .A(ein[476]), .B(n41106), .Z(ereg_next[477]) );
  AND U43742 ( .A(mul_pow), .B(n41107), .Z(n41106) );
  XOR U43743 ( .A(ein[477]), .B(ein[476]), .Z(n41107) );
  XOR U43744 ( .A(ein[475]), .B(n41108), .Z(ereg_next[476]) );
  AND U43745 ( .A(mul_pow), .B(n41109), .Z(n41108) );
  XOR U43746 ( .A(ein[476]), .B(ein[475]), .Z(n41109) );
  XOR U43747 ( .A(ein[474]), .B(n41110), .Z(ereg_next[475]) );
  AND U43748 ( .A(mul_pow), .B(n41111), .Z(n41110) );
  XOR U43749 ( .A(ein[475]), .B(ein[474]), .Z(n41111) );
  XOR U43750 ( .A(ein[473]), .B(n41112), .Z(ereg_next[474]) );
  AND U43751 ( .A(mul_pow), .B(n41113), .Z(n41112) );
  XOR U43752 ( .A(ein[474]), .B(ein[473]), .Z(n41113) );
  XOR U43753 ( .A(ein[472]), .B(n41114), .Z(ereg_next[473]) );
  AND U43754 ( .A(mul_pow), .B(n41115), .Z(n41114) );
  XOR U43755 ( .A(ein[473]), .B(ein[472]), .Z(n41115) );
  XOR U43756 ( .A(ein[471]), .B(n41116), .Z(ereg_next[472]) );
  AND U43757 ( .A(mul_pow), .B(n41117), .Z(n41116) );
  XOR U43758 ( .A(ein[472]), .B(ein[471]), .Z(n41117) );
  XOR U43759 ( .A(ein[470]), .B(n41118), .Z(ereg_next[471]) );
  AND U43760 ( .A(mul_pow), .B(n41119), .Z(n41118) );
  XOR U43761 ( .A(ein[471]), .B(ein[470]), .Z(n41119) );
  XOR U43762 ( .A(ein[469]), .B(n41120), .Z(ereg_next[470]) );
  AND U43763 ( .A(mul_pow), .B(n41121), .Z(n41120) );
  XOR U43764 ( .A(ein[470]), .B(ein[469]), .Z(n41121) );
  XOR U43765 ( .A(ein[45]), .B(n41122), .Z(ereg_next[46]) );
  AND U43766 ( .A(mul_pow), .B(n41123), .Z(n41122) );
  XOR U43767 ( .A(ein[46]), .B(ein[45]), .Z(n41123) );
  XOR U43768 ( .A(ein[468]), .B(n41124), .Z(ereg_next[469]) );
  AND U43769 ( .A(mul_pow), .B(n41125), .Z(n41124) );
  XOR U43770 ( .A(ein[469]), .B(ein[468]), .Z(n41125) );
  XOR U43771 ( .A(ein[467]), .B(n41126), .Z(ereg_next[468]) );
  AND U43772 ( .A(mul_pow), .B(n41127), .Z(n41126) );
  XOR U43773 ( .A(ein[468]), .B(ein[467]), .Z(n41127) );
  XOR U43774 ( .A(ein[466]), .B(n41128), .Z(ereg_next[467]) );
  AND U43775 ( .A(mul_pow), .B(n41129), .Z(n41128) );
  XOR U43776 ( .A(ein[467]), .B(ein[466]), .Z(n41129) );
  XOR U43777 ( .A(ein[465]), .B(n41130), .Z(ereg_next[466]) );
  AND U43778 ( .A(mul_pow), .B(n41131), .Z(n41130) );
  XOR U43779 ( .A(ein[466]), .B(ein[465]), .Z(n41131) );
  XOR U43780 ( .A(ein[464]), .B(n41132), .Z(ereg_next[465]) );
  AND U43781 ( .A(mul_pow), .B(n41133), .Z(n41132) );
  XOR U43782 ( .A(ein[465]), .B(ein[464]), .Z(n41133) );
  XOR U43783 ( .A(ein[463]), .B(n41134), .Z(ereg_next[464]) );
  AND U43784 ( .A(mul_pow), .B(n41135), .Z(n41134) );
  XOR U43785 ( .A(ein[464]), .B(ein[463]), .Z(n41135) );
  XOR U43786 ( .A(ein[462]), .B(n41136), .Z(ereg_next[463]) );
  AND U43787 ( .A(mul_pow), .B(n41137), .Z(n41136) );
  XOR U43788 ( .A(ein[463]), .B(ein[462]), .Z(n41137) );
  XOR U43789 ( .A(ein[461]), .B(n41138), .Z(ereg_next[462]) );
  AND U43790 ( .A(mul_pow), .B(n41139), .Z(n41138) );
  XOR U43791 ( .A(ein[462]), .B(ein[461]), .Z(n41139) );
  XOR U43792 ( .A(ein[460]), .B(n41140), .Z(ereg_next[461]) );
  AND U43793 ( .A(mul_pow), .B(n41141), .Z(n41140) );
  XOR U43794 ( .A(ein[461]), .B(ein[460]), .Z(n41141) );
  XOR U43795 ( .A(ein[459]), .B(n41142), .Z(ereg_next[460]) );
  AND U43796 ( .A(mul_pow), .B(n41143), .Z(n41142) );
  XOR U43797 ( .A(ein[460]), .B(ein[459]), .Z(n41143) );
  XOR U43798 ( .A(ein[44]), .B(n41144), .Z(ereg_next[45]) );
  AND U43799 ( .A(mul_pow), .B(n41145), .Z(n41144) );
  XOR U43800 ( .A(ein[45]), .B(ein[44]), .Z(n41145) );
  XOR U43801 ( .A(ein[458]), .B(n41146), .Z(ereg_next[459]) );
  AND U43802 ( .A(mul_pow), .B(n41147), .Z(n41146) );
  XOR U43803 ( .A(ein[459]), .B(ein[458]), .Z(n41147) );
  XOR U43804 ( .A(ein[457]), .B(n41148), .Z(ereg_next[458]) );
  AND U43805 ( .A(mul_pow), .B(n41149), .Z(n41148) );
  XOR U43806 ( .A(ein[458]), .B(ein[457]), .Z(n41149) );
  XOR U43807 ( .A(ein[456]), .B(n41150), .Z(ereg_next[457]) );
  AND U43808 ( .A(mul_pow), .B(n41151), .Z(n41150) );
  XOR U43809 ( .A(ein[457]), .B(ein[456]), .Z(n41151) );
  XOR U43810 ( .A(ein[455]), .B(n41152), .Z(ereg_next[456]) );
  AND U43811 ( .A(mul_pow), .B(n41153), .Z(n41152) );
  XOR U43812 ( .A(ein[456]), .B(ein[455]), .Z(n41153) );
  XOR U43813 ( .A(ein[454]), .B(n41154), .Z(ereg_next[455]) );
  AND U43814 ( .A(mul_pow), .B(n41155), .Z(n41154) );
  XOR U43815 ( .A(ein[455]), .B(ein[454]), .Z(n41155) );
  XOR U43816 ( .A(ein[453]), .B(n41156), .Z(ereg_next[454]) );
  AND U43817 ( .A(mul_pow), .B(n41157), .Z(n41156) );
  XOR U43818 ( .A(ein[454]), .B(ein[453]), .Z(n41157) );
  XOR U43819 ( .A(ein[452]), .B(n41158), .Z(ereg_next[453]) );
  AND U43820 ( .A(mul_pow), .B(n41159), .Z(n41158) );
  XOR U43821 ( .A(ein[453]), .B(ein[452]), .Z(n41159) );
  XOR U43822 ( .A(ein[451]), .B(n41160), .Z(ereg_next[452]) );
  AND U43823 ( .A(mul_pow), .B(n41161), .Z(n41160) );
  XOR U43824 ( .A(ein[452]), .B(ein[451]), .Z(n41161) );
  XOR U43825 ( .A(ein[450]), .B(n41162), .Z(ereg_next[451]) );
  AND U43826 ( .A(mul_pow), .B(n41163), .Z(n41162) );
  XOR U43827 ( .A(ein[451]), .B(ein[450]), .Z(n41163) );
  XOR U43828 ( .A(ein[449]), .B(n41164), .Z(ereg_next[450]) );
  AND U43829 ( .A(mul_pow), .B(n41165), .Z(n41164) );
  XOR U43830 ( .A(ein[450]), .B(ein[449]), .Z(n41165) );
  XOR U43831 ( .A(ein[43]), .B(n41166), .Z(ereg_next[44]) );
  AND U43832 ( .A(mul_pow), .B(n41167), .Z(n41166) );
  XOR U43833 ( .A(ein[44]), .B(ein[43]), .Z(n41167) );
  XOR U43834 ( .A(ein[448]), .B(n41168), .Z(ereg_next[449]) );
  AND U43835 ( .A(mul_pow), .B(n41169), .Z(n41168) );
  XOR U43836 ( .A(ein[449]), .B(ein[448]), .Z(n41169) );
  XOR U43837 ( .A(ein[447]), .B(n41170), .Z(ereg_next[448]) );
  AND U43838 ( .A(mul_pow), .B(n41171), .Z(n41170) );
  XOR U43839 ( .A(ein[448]), .B(ein[447]), .Z(n41171) );
  XOR U43840 ( .A(ein[446]), .B(n41172), .Z(ereg_next[447]) );
  AND U43841 ( .A(mul_pow), .B(n41173), .Z(n41172) );
  XOR U43842 ( .A(ein[447]), .B(ein[446]), .Z(n41173) );
  XOR U43843 ( .A(ein[445]), .B(n41174), .Z(ereg_next[446]) );
  AND U43844 ( .A(mul_pow), .B(n41175), .Z(n41174) );
  XOR U43845 ( .A(ein[446]), .B(ein[445]), .Z(n41175) );
  XOR U43846 ( .A(ein[444]), .B(n41176), .Z(ereg_next[445]) );
  AND U43847 ( .A(mul_pow), .B(n41177), .Z(n41176) );
  XOR U43848 ( .A(ein[445]), .B(ein[444]), .Z(n41177) );
  XOR U43849 ( .A(ein[443]), .B(n41178), .Z(ereg_next[444]) );
  AND U43850 ( .A(mul_pow), .B(n41179), .Z(n41178) );
  XOR U43851 ( .A(ein[444]), .B(ein[443]), .Z(n41179) );
  XOR U43852 ( .A(ein[442]), .B(n41180), .Z(ereg_next[443]) );
  AND U43853 ( .A(mul_pow), .B(n41181), .Z(n41180) );
  XOR U43854 ( .A(ein[443]), .B(ein[442]), .Z(n41181) );
  XOR U43855 ( .A(ein[441]), .B(n41182), .Z(ereg_next[442]) );
  AND U43856 ( .A(mul_pow), .B(n41183), .Z(n41182) );
  XOR U43857 ( .A(ein[442]), .B(ein[441]), .Z(n41183) );
  XOR U43858 ( .A(ein[440]), .B(n41184), .Z(ereg_next[441]) );
  AND U43859 ( .A(mul_pow), .B(n41185), .Z(n41184) );
  XOR U43860 ( .A(ein[441]), .B(ein[440]), .Z(n41185) );
  XOR U43861 ( .A(ein[439]), .B(n41186), .Z(ereg_next[440]) );
  AND U43862 ( .A(mul_pow), .B(n41187), .Z(n41186) );
  XOR U43863 ( .A(ein[440]), .B(ein[439]), .Z(n41187) );
  XOR U43864 ( .A(ein[42]), .B(n41188), .Z(ereg_next[43]) );
  AND U43865 ( .A(mul_pow), .B(n41189), .Z(n41188) );
  XOR U43866 ( .A(ein[43]), .B(ein[42]), .Z(n41189) );
  XOR U43867 ( .A(ein[438]), .B(n41190), .Z(ereg_next[439]) );
  AND U43868 ( .A(mul_pow), .B(n41191), .Z(n41190) );
  XOR U43869 ( .A(ein[439]), .B(ein[438]), .Z(n41191) );
  XOR U43870 ( .A(ein[437]), .B(n41192), .Z(ereg_next[438]) );
  AND U43871 ( .A(mul_pow), .B(n41193), .Z(n41192) );
  XOR U43872 ( .A(ein[438]), .B(ein[437]), .Z(n41193) );
  XOR U43873 ( .A(ein[436]), .B(n41194), .Z(ereg_next[437]) );
  AND U43874 ( .A(mul_pow), .B(n41195), .Z(n41194) );
  XOR U43875 ( .A(ein[437]), .B(ein[436]), .Z(n41195) );
  XOR U43876 ( .A(ein[435]), .B(n41196), .Z(ereg_next[436]) );
  AND U43877 ( .A(mul_pow), .B(n41197), .Z(n41196) );
  XOR U43878 ( .A(ein[436]), .B(ein[435]), .Z(n41197) );
  XOR U43879 ( .A(ein[434]), .B(n41198), .Z(ereg_next[435]) );
  AND U43880 ( .A(mul_pow), .B(n41199), .Z(n41198) );
  XOR U43881 ( .A(ein[435]), .B(ein[434]), .Z(n41199) );
  XOR U43882 ( .A(ein[433]), .B(n41200), .Z(ereg_next[434]) );
  AND U43883 ( .A(mul_pow), .B(n41201), .Z(n41200) );
  XOR U43884 ( .A(ein[434]), .B(ein[433]), .Z(n41201) );
  XOR U43885 ( .A(ein[432]), .B(n41202), .Z(ereg_next[433]) );
  AND U43886 ( .A(mul_pow), .B(n41203), .Z(n41202) );
  XOR U43887 ( .A(ein[433]), .B(ein[432]), .Z(n41203) );
  XOR U43888 ( .A(ein[431]), .B(n41204), .Z(ereg_next[432]) );
  AND U43889 ( .A(mul_pow), .B(n41205), .Z(n41204) );
  XOR U43890 ( .A(ein[432]), .B(ein[431]), .Z(n41205) );
  XOR U43891 ( .A(ein[430]), .B(n41206), .Z(ereg_next[431]) );
  AND U43892 ( .A(mul_pow), .B(n41207), .Z(n41206) );
  XOR U43893 ( .A(ein[431]), .B(ein[430]), .Z(n41207) );
  XOR U43894 ( .A(ein[429]), .B(n41208), .Z(ereg_next[430]) );
  AND U43895 ( .A(mul_pow), .B(n41209), .Z(n41208) );
  XOR U43896 ( .A(ein[430]), .B(ein[429]), .Z(n41209) );
  XOR U43897 ( .A(ein[41]), .B(n41210), .Z(ereg_next[42]) );
  AND U43898 ( .A(mul_pow), .B(n41211), .Z(n41210) );
  XOR U43899 ( .A(ein[42]), .B(ein[41]), .Z(n41211) );
  XOR U43900 ( .A(ein[428]), .B(n41212), .Z(ereg_next[429]) );
  AND U43901 ( .A(mul_pow), .B(n41213), .Z(n41212) );
  XOR U43902 ( .A(ein[429]), .B(ein[428]), .Z(n41213) );
  XOR U43903 ( .A(ein[427]), .B(n41214), .Z(ereg_next[428]) );
  AND U43904 ( .A(mul_pow), .B(n41215), .Z(n41214) );
  XOR U43905 ( .A(ein[428]), .B(ein[427]), .Z(n41215) );
  XOR U43906 ( .A(ein[426]), .B(n41216), .Z(ereg_next[427]) );
  AND U43907 ( .A(mul_pow), .B(n41217), .Z(n41216) );
  XOR U43908 ( .A(ein[427]), .B(ein[426]), .Z(n41217) );
  XOR U43909 ( .A(ein[425]), .B(n41218), .Z(ereg_next[426]) );
  AND U43910 ( .A(mul_pow), .B(n41219), .Z(n41218) );
  XOR U43911 ( .A(ein[426]), .B(ein[425]), .Z(n41219) );
  XOR U43912 ( .A(ein[424]), .B(n41220), .Z(ereg_next[425]) );
  AND U43913 ( .A(mul_pow), .B(n41221), .Z(n41220) );
  XOR U43914 ( .A(ein[425]), .B(ein[424]), .Z(n41221) );
  XOR U43915 ( .A(ein[423]), .B(n41222), .Z(ereg_next[424]) );
  AND U43916 ( .A(mul_pow), .B(n41223), .Z(n41222) );
  XOR U43917 ( .A(ein[424]), .B(ein[423]), .Z(n41223) );
  XOR U43918 ( .A(ein[422]), .B(n41224), .Z(ereg_next[423]) );
  AND U43919 ( .A(mul_pow), .B(n41225), .Z(n41224) );
  XOR U43920 ( .A(ein[423]), .B(ein[422]), .Z(n41225) );
  XOR U43921 ( .A(ein[421]), .B(n41226), .Z(ereg_next[422]) );
  AND U43922 ( .A(mul_pow), .B(n41227), .Z(n41226) );
  XOR U43923 ( .A(ein[422]), .B(ein[421]), .Z(n41227) );
  XOR U43924 ( .A(ein[420]), .B(n41228), .Z(ereg_next[421]) );
  AND U43925 ( .A(mul_pow), .B(n41229), .Z(n41228) );
  XOR U43926 ( .A(ein[421]), .B(ein[420]), .Z(n41229) );
  XOR U43927 ( .A(ein[419]), .B(n41230), .Z(ereg_next[420]) );
  AND U43928 ( .A(mul_pow), .B(n41231), .Z(n41230) );
  XOR U43929 ( .A(ein[420]), .B(ein[419]), .Z(n41231) );
  XOR U43930 ( .A(ein[40]), .B(n41232), .Z(ereg_next[41]) );
  AND U43931 ( .A(mul_pow), .B(n41233), .Z(n41232) );
  XOR U43932 ( .A(ein[41]), .B(ein[40]), .Z(n41233) );
  XOR U43933 ( .A(ein[418]), .B(n41234), .Z(ereg_next[419]) );
  AND U43934 ( .A(mul_pow), .B(n41235), .Z(n41234) );
  XOR U43935 ( .A(ein[419]), .B(ein[418]), .Z(n41235) );
  XOR U43936 ( .A(ein[417]), .B(n41236), .Z(ereg_next[418]) );
  AND U43937 ( .A(mul_pow), .B(n41237), .Z(n41236) );
  XOR U43938 ( .A(ein[418]), .B(ein[417]), .Z(n41237) );
  XOR U43939 ( .A(ein[416]), .B(n41238), .Z(ereg_next[417]) );
  AND U43940 ( .A(mul_pow), .B(n41239), .Z(n41238) );
  XOR U43941 ( .A(ein[417]), .B(ein[416]), .Z(n41239) );
  XOR U43942 ( .A(ein[415]), .B(n41240), .Z(ereg_next[416]) );
  AND U43943 ( .A(mul_pow), .B(n41241), .Z(n41240) );
  XOR U43944 ( .A(ein[416]), .B(ein[415]), .Z(n41241) );
  XOR U43945 ( .A(ein[414]), .B(n41242), .Z(ereg_next[415]) );
  AND U43946 ( .A(mul_pow), .B(n41243), .Z(n41242) );
  XOR U43947 ( .A(ein[415]), .B(ein[414]), .Z(n41243) );
  XOR U43948 ( .A(ein[413]), .B(n41244), .Z(ereg_next[414]) );
  AND U43949 ( .A(mul_pow), .B(n41245), .Z(n41244) );
  XOR U43950 ( .A(ein[414]), .B(ein[413]), .Z(n41245) );
  XOR U43951 ( .A(ein[412]), .B(n41246), .Z(ereg_next[413]) );
  AND U43952 ( .A(mul_pow), .B(n41247), .Z(n41246) );
  XOR U43953 ( .A(ein[413]), .B(ein[412]), .Z(n41247) );
  XOR U43954 ( .A(ein[411]), .B(n41248), .Z(ereg_next[412]) );
  AND U43955 ( .A(mul_pow), .B(n41249), .Z(n41248) );
  XOR U43956 ( .A(ein[412]), .B(ein[411]), .Z(n41249) );
  XOR U43957 ( .A(ein[410]), .B(n41250), .Z(ereg_next[411]) );
  AND U43958 ( .A(mul_pow), .B(n41251), .Z(n41250) );
  XOR U43959 ( .A(ein[411]), .B(ein[410]), .Z(n41251) );
  XOR U43960 ( .A(ein[409]), .B(n41252), .Z(ereg_next[410]) );
  AND U43961 ( .A(mul_pow), .B(n41253), .Z(n41252) );
  XOR U43962 ( .A(ein[410]), .B(ein[409]), .Z(n41253) );
  XOR U43963 ( .A(ein[39]), .B(n41254), .Z(ereg_next[40]) );
  AND U43964 ( .A(mul_pow), .B(n41255), .Z(n41254) );
  XOR U43965 ( .A(ein[40]), .B(ein[39]), .Z(n41255) );
  XOR U43966 ( .A(ein[408]), .B(n41256), .Z(ereg_next[409]) );
  AND U43967 ( .A(mul_pow), .B(n41257), .Z(n41256) );
  XOR U43968 ( .A(ein[409]), .B(ein[408]), .Z(n41257) );
  XOR U43969 ( .A(ein[407]), .B(n41258), .Z(ereg_next[408]) );
  AND U43970 ( .A(mul_pow), .B(n41259), .Z(n41258) );
  XOR U43971 ( .A(ein[408]), .B(ein[407]), .Z(n41259) );
  XOR U43972 ( .A(ein[406]), .B(n41260), .Z(ereg_next[407]) );
  AND U43973 ( .A(mul_pow), .B(n41261), .Z(n41260) );
  XOR U43974 ( .A(ein[407]), .B(ein[406]), .Z(n41261) );
  XOR U43975 ( .A(ein[405]), .B(n41262), .Z(ereg_next[406]) );
  AND U43976 ( .A(mul_pow), .B(n41263), .Z(n41262) );
  XOR U43977 ( .A(ein[406]), .B(ein[405]), .Z(n41263) );
  XOR U43978 ( .A(ein[404]), .B(n41264), .Z(ereg_next[405]) );
  AND U43979 ( .A(mul_pow), .B(n41265), .Z(n41264) );
  XOR U43980 ( .A(ein[405]), .B(ein[404]), .Z(n41265) );
  XOR U43981 ( .A(ein[403]), .B(n41266), .Z(ereg_next[404]) );
  AND U43982 ( .A(mul_pow), .B(n41267), .Z(n41266) );
  XOR U43983 ( .A(ein[404]), .B(ein[403]), .Z(n41267) );
  XOR U43984 ( .A(ein[402]), .B(n41268), .Z(ereg_next[403]) );
  AND U43985 ( .A(mul_pow), .B(n41269), .Z(n41268) );
  XOR U43986 ( .A(ein[403]), .B(ein[402]), .Z(n41269) );
  XOR U43987 ( .A(ein[401]), .B(n41270), .Z(ereg_next[402]) );
  AND U43988 ( .A(mul_pow), .B(n41271), .Z(n41270) );
  XOR U43989 ( .A(ein[402]), .B(ein[401]), .Z(n41271) );
  XOR U43990 ( .A(ein[400]), .B(n41272), .Z(ereg_next[401]) );
  AND U43991 ( .A(mul_pow), .B(n41273), .Z(n41272) );
  XOR U43992 ( .A(ein[401]), .B(ein[400]), .Z(n41273) );
  XOR U43993 ( .A(ein[399]), .B(n41274), .Z(ereg_next[400]) );
  AND U43994 ( .A(mul_pow), .B(n41275), .Z(n41274) );
  XOR U43995 ( .A(ein[400]), .B(ein[399]), .Z(n41275) );
  XOR U43996 ( .A(ein[2]), .B(n41276), .Z(ereg_next[3]) );
  AND U43997 ( .A(mul_pow), .B(n41277), .Z(n41276) );
  XOR U43998 ( .A(ein[3]), .B(ein[2]), .Z(n41277) );
  XOR U43999 ( .A(ein[38]), .B(n41278), .Z(ereg_next[39]) );
  AND U44000 ( .A(mul_pow), .B(n41279), .Z(n41278) );
  XOR U44001 ( .A(ein[39]), .B(ein[38]), .Z(n41279) );
  XOR U44002 ( .A(ein[398]), .B(n41280), .Z(ereg_next[399]) );
  AND U44003 ( .A(mul_pow), .B(n41281), .Z(n41280) );
  XOR U44004 ( .A(ein[399]), .B(ein[398]), .Z(n41281) );
  XOR U44005 ( .A(ein[397]), .B(n41282), .Z(ereg_next[398]) );
  AND U44006 ( .A(mul_pow), .B(n41283), .Z(n41282) );
  XOR U44007 ( .A(ein[398]), .B(ein[397]), .Z(n41283) );
  XOR U44008 ( .A(ein[396]), .B(n41284), .Z(ereg_next[397]) );
  AND U44009 ( .A(mul_pow), .B(n41285), .Z(n41284) );
  XOR U44010 ( .A(ein[397]), .B(ein[396]), .Z(n41285) );
  XOR U44011 ( .A(ein[395]), .B(n41286), .Z(ereg_next[396]) );
  AND U44012 ( .A(mul_pow), .B(n41287), .Z(n41286) );
  XOR U44013 ( .A(ein[396]), .B(ein[395]), .Z(n41287) );
  XOR U44014 ( .A(ein[394]), .B(n41288), .Z(ereg_next[395]) );
  AND U44015 ( .A(mul_pow), .B(n41289), .Z(n41288) );
  XOR U44016 ( .A(ein[395]), .B(ein[394]), .Z(n41289) );
  XOR U44017 ( .A(ein[393]), .B(n41290), .Z(ereg_next[394]) );
  AND U44018 ( .A(mul_pow), .B(n41291), .Z(n41290) );
  XOR U44019 ( .A(ein[394]), .B(ein[393]), .Z(n41291) );
  XOR U44020 ( .A(ein[392]), .B(n41292), .Z(ereg_next[393]) );
  AND U44021 ( .A(mul_pow), .B(n41293), .Z(n41292) );
  XOR U44022 ( .A(ein[393]), .B(ein[392]), .Z(n41293) );
  XOR U44023 ( .A(ein[391]), .B(n41294), .Z(ereg_next[392]) );
  AND U44024 ( .A(mul_pow), .B(n41295), .Z(n41294) );
  XOR U44025 ( .A(ein[392]), .B(ein[391]), .Z(n41295) );
  XOR U44026 ( .A(ein[390]), .B(n41296), .Z(ereg_next[391]) );
  AND U44027 ( .A(mul_pow), .B(n41297), .Z(n41296) );
  XOR U44028 ( .A(ein[391]), .B(ein[390]), .Z(n41297) );
  XOR U44029 ( .A(ein[389]), .B(n41298), .Z(ereg_next[390]) );
  AND U44030 ( .A(mul_pow), .B(n41299), .Z(n41298) );
  XOR U44031 ( .A(ein[390]), .B(ein[389]), .Z(n41299) );
  XOR U44032 ( .A(ein[37]), .B(n41300), .Z(ereg_next[38]) );
  AND U44033 ( .A(mul_pow), .B(n41301), .Z(n41300) );
  XOR U44034 ( .A(ein[38]), .B(ein[37]), .Z(n41301) );
  XOR U44035 ( .A(ein[388]), .B(n41302), .Z(ereg_next[389]) );
  AND U44036 ( .A(mul_pow), .B(n41303), .Z(n41302) );
  XOR U44037 ( .A(ein[389]), .B(ein[388]), .Z(n41303) );
  XOR U44038 ( .A(ein[387]), .B(n41304), .Z(ereg_next[388]) );
  AND U44039 ( .A(mul_pow), .B(n41305), .Z(n41304) );
  XOR U44040 ( .A(ein[388]), .B(ein[387]), .Z(n41305) );
  XOR U44041 ( .A(ein[386]), .B(n41306), .Z(ereg_next[387]) );
  AND U44042 ( .A(mul_pow), .B(n41307), .Z(n41306) );
  XOR U44043 ( .A(ein[387]), .B(ein[386]), .Z(n41307) );
  XOR U44044 ( .A(ein[385]), .B(n41308), .Z(ereg_next[386]) );
  AND U44045 ( .A(mul_pow), .B(n41309), .Z(n41308) );
  XOR U44046 ( .A(ein[386]), .B(ein[385]), .Z(n41309) );
  XOR U44047 ( .A(ein[384]), .B(n41310), .Z(ereg_next[385]) );
  AND U44048 ( .A(mul_pow), .B(n41311), .Z(n41310) );
  XOR U44049 ( .A(ein[385]), .B(ein[384]), .Z(n41311) );
  XOR U44050 ( .A(ein[383]), .B(n41312), .Z(ereg_next[384]) );
  AND U44051 ( .A(mul_pow), .B(n41313), .Z(n41312) );
  XOR U44052 ( .A(ein[384]), .B(ein[383]), .Z(n41313) );
  XOR U44053 ( .A(ein[382]), .B(n41314), .Z(ereg_next[383]) );
  AND U44054 ( .A(mul_pow), .B(n41315), .Z(n41314) );
  XOR U44055 ( .A(ein[383]), .B(ein[382]), .Z(n41315) );
  XOR U44056 ( .A(ein[381]), .B(n41316), .Z(ereg_next[382]) );
  AND U44057 ( .A(mul_pow), .B(n41317), .Z(n41316) );
  XOR U44058 ( .A(ein[382]), .B(ein[381]), .Z(n41317) );
  XOR U44059 ( .A(ein[380]), .B(n41318), .Z(ereg_next[381]) );
  AND U44060 ( .A(mul_pow), .B(n41319), .Z(n41318) );
  XOR U44061 ( .A(ein[381]), .B(ein[380]), .Z(n41319) );
  XOR U44062 ( .A(ein[379]), .B(n41320), .Z(ereg_next[380]) );
  AND U44063 ( .A(mul_pow), .B(n41321), .Z(n41320) );
  XOR U44064 ( .A(ein[380]), .B(ein[379]), .Z(n41321) );
  XOR U44065 ( .A(ein[36]), .B(n41322), .Z(ereg_next[37]) );
  AND U44066 ( .A(mul_pow), .B(n41323), .Z(n41322) );
  XOR U44067 ( .A(ein[37]), .B(ein[36]), .Z(n41323) );
  XOR U44068 ( .A(ein[378]), .B(n41324), .Z(ereg_next[379]) );
  AND U44069 ( .A(mul_pow), .B(n41325), .Z(n41324) );
  XOR U44070 ( .A(ein[379]), .B(ein[378]), .Z(n41325) );
  XOR U44071 ( .A(ein[377]), .B(n41326), .Z(ereg_next[378]) );
  AND U44072 ( .A(mul_pow), .B(n41327), .Z(n41326) );
  XOR U44073 ( .A(ein[378]), .B(ein[377]), .Z(n41327) );
  XOR U44074 ( .A(ein[376]), .B(n41328), .Z(ereg_next[377]) );
  AND U44075 ( .A(mul_pow), .B(n41329), .Z(n41328) );
  XOR U44076 ( .A(ein[377]), .B(ein[376]), .Z(n41329) );
  XOR U44077 ( .A(ein[375]), .B(n41330), .Z(ereg_next[376]) );
  AND U44078 ( .A(mul_pow), .B(n41331), .Z(n41330) );
  XOR U44079 ( .A(ein[376]), .B(ein[375]), .Z(n41331) );
  XOR U44080 ( .A(ein[374]), .B(n41332), .Z(ereg_next[375]) );
  AND U44081 ( .A(mul_pow), .B(n41333), .Z(n41332) );
  XOR U44082 ( .A(ein[375]), .B(ein[374]), .Z(n41333) );
  XOR U44083 ( .A(ein[373]), .B(n41334), .Z(ereg_next[374]) );
  AND U44084 ( .A(mul_pow), .B(n41335), .Z(n41334) );
  XOR U44085 ( .A(ein[374]), .B(ein[373]), .Z(n41335) );
  XOR U44086 ( .A(ein[372]), .B(n41336), .Z(ereg_next[373]) );
  AND U44087 ( .A(mul_pow), .B(n41337), .Z(n41336) );
  XOR U44088 ( .A(ein[373]), .B(ein[372]), .Z(n41337) );
  XOR U44089 ( .A(ein[371]), .B(n41338), .Z(ereg_next[372]) );
  AND U44090 ( .A(mul_pow), .B(n41339), .Z(n41338) );
  XOR U44091 ( .A(ein[372]), .B(ein[371]), .Z(n41339) );
  XOR U44092 ( .A(ein[370]), .B(n41340), .Z(ereg_next[371]) );
  AND U44093 ( .A(mul_pow), .B(n41341), .Z(n41340) );
  XOR U44094 ( .A(ein[371]), .B(ein[370]), .Z(n41341) );
  XOR U44095 ( .A(ein[369]), .B(n41342), .Z(ereg_next[370]) );
  AND U44096 ( .A(mul_pow), .B(n41343), .Z(n41342) );
  XOR U44097 ( .A(ein[370]), .B(ein[369]), .Z(n41343) );
  XOR U44098 ( .A(ein[35]), .B(n41344), .Z(ereg_next[36]) );
  AND U44099 ( .A(mul_pow), .B(n41345), .Z(n41344) );
  XOR U44100 ( .A(ein[36]), .B(ein[35]), .Z(n41345) );
  XOR U44101 ( .A(ein[368]), .B(n41346), .Z(ereg_next[369]) );
  AND U44102 ( .A(mul_pow), .B(n41347), .Z(n41346) );
  XOR U44103 ( .A(ein[369]), .B(ein[368]), .Z(n41347) );
  XOR U44104 ( .A(ein[367]), .B(n41348), .Z(ereg_next[368]) );
  AND U44105 ( .A(mul_pow), .B(n41349), .Z(n41348) );
  XOR U44106 ( .A(ein[368]), .B(ein[367]), .Z(n41349) );
  XOR U44107 ( .A(ein[366]), .B(n41350), .Z(ereg_next[367]) );
  AND U44108 ( .A(mul_pow), .B(n41351), .Z(n41350) );
  XOR U44109 ( .A(ein[367]), .B(ein[366]), .Z(n41351) );
  XOR U44110 ( .A(ein[365]), .B(n41352), .Z(ereg_next[366]) );
  AND U44111 ( .A(mul_pow), .B(n41353), .Z(n41352) );
  XOR U44112 ( .A(ein[366]), .B(ein[365]), .Z(n41353) );
  XOR U44113 ( .A(ein[364]), .B(n41354), .Z(ereg_next[365]) );
  AND U44114 ( .A(mul_pow), .B(n41355), .Z(n41354) );
  XOR U44115 ( .A(ein[365]), .B(ein[364]), .Z(n41355) );
  XOR U44116 ( .A(ein[363]), .B(n41356), .Z(ereg_next[364]) );
  AND U44117 ( .A(mul_pow), .B(n41357), .Z(n41356) );
  XOR U44118 ( .A(ein[364]), .B(ein[363]), .Z(n41357) );
  XOR U44119 ( .A(ein[362]), .B(n41358), .Z(ereg_next[363]) );
  AND U44120 ( .A(mul_pow), .B(n41359), .Z(n41358) );
  XOR U44121 ( .A(ein[363]), .B(ein[362]), .Z(n41359) );
  XOR U44122 ( .A(ein[361]), .B(n41360), .Z(ereg_next[362]) );
  AND U44123 ( .A(mul_pow), .B(n41361), .Z(n41360) );
  XOR U44124 ( .A(ein[362]), .B(ein[361]), .Z(n41361) );
  XOR U44125 ( .A(ein[360]), .B(n41362), .Z(ereg_next[361]) );
  AND U44126 ( .A(mul_pow), .B(n41363), .Z(n41362) );
  XOR U44127 ( .A(ein[361]), .B(ein[360]), .Z(n41363) );
  XOR U44128 ( .A(ein[359]), .B(n41364), .Z(ereg_next[360]) );
  AND U44129 ( .A(mul_pow), .B(n41365), .Z(n41364) );
  XOR U44130 ( .A(ein[360]), .B(ein[359]), .Z(n41365) );
  XOR U44131 ( .A(ein[34]), .B(n41366), .Z(ereg_next[35]) );
  AND U44132 ( .A(mul_pow), .B(n41367), .Z(n41366) );
  XOR U44133 ( .A(ein[35]), .B(ein[34]), .Z(n41367) );
  XOR U44134 ( .A(ein[358]), .B(n41368), .Z(ereg_next[359]) );
  AND U44135 ( .A(mul_pow), .B(n41369), .Z(n41368) );
  XOR U44136 ( .A(ein[359]), .B(ein[358]), .Z(n41369) );
  XOR U44137 ( .A(ein[357]), .B(n41370), .Z(ereg_next[358]) );
  AND U44138 ( .A(mul_pow), .B(n41371), .Z(n41370) );
  XOR U44139 ( .A(ein[358]), .B(ein[357]), .Z(n41371) );
  XOR U44140 ( .A(ein[356]), .B(n41372), .Z(ereg_next[357]) );
  AND U44141 ( .A(mul_pow), .B(n41373), .Z(n41372) );
  XOR U44142 ( .A(ein[357]), .B(ein[356]), .Z(n41373) );
  XOR U44143 ( .A(ein[355]), .B(n41374), .Z(ereg_next[356]) );
  AND U44144 ( .A(mul_pow), .B(n41375), .Z(n41374) );
  XOR U44145 ( .A(ein[356]), .B(ein[355]), .Z(n41375) );
  XOR U44146 ( .A(ein[354]), .B(n41376), .Z(ereg_next[355]) );
  AND U44147 ( .A(mul_pow), .B(n41377), .Z(n41376) );
  XOR U44148 ( .A(ein[355]), .B(ein[354]), .Z(n41377) );
  XOR U44149 ( .A(ein[353]), .B(n41378), .Z(ereg_next[354]) );
  AND U44150 ( .A(mul_pow), .B(n41379), .Z(n41378) );
  XOR U44151 ( .A(ein[354]), .B(ein[353]), .Z(n41379) );
  XOR U44152 ( .A(ein[352]), .B(n41380), .Z(ereg_next[353]) );
  AND U44153 ( .A(mul_pow), .B(n41381), .Z(n41380) );
  XOR U44154 ( .A(ein[353]), .B(ein[352]), .Z(n41381) );
  XOR U44155 ( .A(ein[351]), .B(n41382), .Z(ereg_next[352]) );
  AND U44156 ( .A(mul_pow), .B(n41383), .Z(n41382) );
  XOR U44157 ( .A(ein[352]), .B(ein[351]), .Z(n41383) );
  XOR U44158 ( .A(ein[350]), .B(n41384), .Z(ereg_next[351]) );
  AND U44159 ( .A(mul_pow), .B(n41385), .Z(n41384) );
  XOR U44160 ( .A(ein[351]), .B(ein[350]), .Z(n41385) );
  XOR U44161 ( .A(ein[349]), .B(n41386), .Z(ereg_next[350]) );
  AND U44162 ( .A(mul_pow), .B(n41387), .Z(n41386) );
  XOR U44163 ( .A(ein[350]), .B(ein[349]), .Z(n41387) );
  XOR U44164 ( .A(ein[33]), .B(n41388), .Z(ereg_next[34]) );
  AND U44165 ( .A(mul_pow), .B(n41389), .Z(n41388) );
  XOR U44166 ( .A(ein[34]), .B(ein[33]), .Z(n41389) );
  XOR U44167 ( .A(ein[348]), .B(n41390), .Z(ereg_next[349]) );
  AND U44168 ( .A(mul_pow), .B(n41391), .Z(n41390) );
  XOR U44169 ( .A(ein[349]), .B(ein[348]), .Z(n41391) );
  XOR U44170 ( .A(ein[347]), .B(n41392), .Z(ereg_next[348]) );
  AND U44171 ( .A(mul_pow), .B(n41393), .Z(n41392) );
  XOR U44172 ( .A(ein[348]), .B(ein[347]), .Z(n41393) );
  XOR U44173 ( .A(ein[346]), .B(n41394), .Z(ereg_next[347]) );
  AND U44174 ( .A(mul_pow), .B(n41395), .Z(n41394) );
  XOR U44175 ( .A(ein[347]), .B(ein[346]), .Z(n41395) );
  XOR U44176 ( .A(ein[345]), .B(n41396), .Z(ereg_next[346]) );
  AND U44177 ( .A(mul_pow), .B(n41397), .Z(n41396) );
  XOR U44178 ( .A(ein[346]), .B(ein[345]), .Z(n41397) );
  XOR U44179 ( .A(ein[344]), .B(n41398), .Z(ereg_next[345]) );
  AND U44180 ( .A(mul_pow), .B(n41399), .Z(n41398) );
  XOR U44181 ( .A(ein[345]), .B(ein[344]), .Z(n41399) );
  XOR U44182 ( .A(ein[343]), .B(n41400), .Z(ereg_next[344]) );
  AND U44183 ( .A(mul_pow), .B(n41401), .Z(n41400) );
  XOR U44184 ( .A(ein[344]), .B(ein[343]), .Z(n41401) );
  XOR U44185 ( .A(ein[342]), .B(n41402), .Z(ereg_next[343]) );
  AND U44186 ( .A(mul_pow), .B(n41403), .Z(n41402) );
  XOR U44187 ( .A(ein[343]), .B(ein[342]), .Z(n41403) );
  XOR U44188 ( .A(ein[341]), .B(n41404), .Z(ereg_next[342]) );
  AND U44189 ( .A(mul_pow), .B(n41405), .Z(n41404) );
  XOR U44190 ( .A(ein[342]), .B(ein[341]), .Z(n41405) );
  XOR U44191 ( .A(ein[340]), .B(n41406), .Z(ereg_next[341]) );
  AND U44192 ( .A(mul_pow), .B(n41407), .Z(n41406) );
  XOR U44193 ( .A(ein[341]), .B(ein[340]), .Z(n41407) );
  XOR U44194 ( .A(ein[339]), .B(n41408), .Z(ereg_next[340]) );
  AND U44195 ( .A(mul_pow), .B(n41409), .Z(n41408) );
  XOR U44196 ( .A(ein[340]), .B(ein[339]), .Z(n41409) );
  XOR U44197 ( .A(ein[32]), .B(n41410), .Z(ereg_next[33]) );
  AND U44198 ( .A(mul_pow), .B(n41411), .Z(n41410) );
  XOR U44199 ( .A(ein[33]), .B(ein[32]), .Z(n41411) );
  XOR U44200 ( .A(ein[338]), .B(n41412), .Z(ereg_next[339]) );
  AND U44201 ( .A(mul_pow), .B(n41413), .Z(n41412) );
  XOR U44202 ( .A(ein[339]), .B(ein[338]), .Z(n41413) );
  XOR U44203 ( .A(ein[337]), .B(n41414), .Z(ereg_next[338]) );
  AND U44204 ( .A(mul_pow), .B(n41415), .Z(n41414) );
  XOR U44205 ( .A(ein[338]), .B(ein[337]), .Z(n41415) );
  XOR U44206 ( .A(ein[336]), .B(n41416), .Z(ereg_next[337]) );
  AND U44207 ( .A(mul_pow), .B(n41417), .Z(n41416) );
  XOR U44208 ( .A(ein[337]), .B(ein[336]), .Z(n41417) );
  XOR U44209 ( .A(ein[335]), .B(n41418), .Z(ereg_next[336]) );
  AND U44210 ( .A(mul_pow), .B(n41419), .Z(n41418) );
  XOR U44211 ( .A(ein[336]), .B(ein[335]), .Z(n41419) );
  XOR U44212 ( .A(ein[334]), .B(n41420), .Z(ereg_next[335]) );
  AND U44213 ( .A(mul_pow), .B(n41421), .Z(n41420) );
  XOR U44214 ( .A(ein[335]), .B(ein[334]), .Z(n41421) );
  XOR U44215 ( .A(ein[333]), .B(n41422), .Z(ereg_next[334]) );
  AND U44216 ( .A(mul_pow), .B(n41423), .Z(n41422) );
  XOR U44217 ( .A(ein[334]), .B(ein[333]), .Z(n41423) );
  XOR U44218 ( .A(ein[332]), .B(n41424), .Z(ereg_next[333]) );
  AND U44219 ( .A(mul_pow), .B(n41425), .Z(n41424) );
  XOR U44220 ( .A(ein[333]), .B(ein[332]), .Z(n41425) );
  XOR U44221 ( .A(ein[331]), .B(n41426), .Z(ereg_next[332]) );
  AND U44222 ( .A(mul_pow), .B(n41427), .Z(n41426) );
  XOR U44223 ( .A(ein[332]), .B(ein[331]), .Z(n41427) );
  XOR U44224 ( .A(ein[330]), .B(n41428), .Z(ereg_next[331]) );
  AND U44225 ( .A(mul_pow), .B(n41429), .Z(n41428) );
  XOR U44226 ( .A(ein[331]), .B(ein[330]), .Z(n41429) );
  XOR U44227 ( .A(ein[329]), .B(n41430), .Z(ereg_next[330]) );
  AND U44228 ( .A(mul_pow), .B(n41431), .Z(n41430) );
  XOR U44229 ( .A(ein[330]), .B(ein[329]), .Z(n41431) );
  XOR U44230 ( .A(ein[31]), .B(n41432), .Z(ereg_next[32]) );
  AND U44231 ( .A(mul_pow), .B(n41433), .Z(n41432) );
  XOR U44232 ( .A(ein[32]), .B(ein[31]), .Z(n41433) );
  XOR U44233 ( .A(ein[328]), .B(n41434), .Z(ereg_next[329]) );
  AND U44234 ( .A(mul_pow), .B(n41435), .Z(n41434) );
  XOR U44235 ( .A(ein[329]), .B(ein[328]), .Z(n41435) );
  XOR U44236 ( .A(ein[327]), .B(n41436), .Z(ereg_next[328]) );
  AND U44237 ( .A(mul_pow), .B(n41437), .Z(n41436) );
  XOR U44238 ( .A(ein[328]), .B(ein[327]), .Z(n41437) );
  XOR U44239 ( .A(ein[326]), .B(n41438), .Z(ereg_next[327]) );
  AND U44240 ( .A(mul_pow), .B(n41439), .Z(n41438) );
  XOR U44241 ( .A(ein[327]), .B(ein[326]), .Z(n41439) );
  XOR U44242 ( .A(ein[325]), .B(n41440), .Z(ereg_next[326]) );
  AND U44243 ( .A(mul_pow), .B(n41441), .Z(n41440) );
  XOR U44244 ( .A(ein[326]), .B(ein[325]), .Z(n41441) );
  XOR U44245 ( .A(ein[324]), .B(n41442), .Z(ereg_next[325]) );
  AND U44246 ( .A(mul_pow), .B(n41443), .Z(n41442) );
  XOR U44247 ( .A(ein[325]), .B(ein[324]), .Z(n41443) );
  XOR U44248 ( .A(ein[323]), .B(n41444), .Z(ereg_next[324]) );
  AND U44249 ( .A(mul_pow), .B(n41445), .Z(n41444) );
  XOR U44250 ( .A(ein[324]), .B(ein[323]), .Z(n41445) );
  XOR U44251 ( .A(ein[322]), .B(n41446), .Z(ereg_next[323]) );
  AND U44252 ( .A(mul_pow), .B(n41447), .Z(n41446) );
  XOR U44253 ( .A(ein[323]), .B(ein[322]), .Z(n41447) );
  XOR U44254 ( .A(ein[321]), .B(n41448), .Z(ereg_next[322]) );
  AND U44255 ( .A(mul_pow), .B(n41449), .Z(n41448) );
  XOR U44256 ( .A(ein[322]), .B(ein[321]), .Z(n41449) );
  XOR U44257 ( .A(ein[320]), .B(n41450), .Z(ereg_next[321]) );
  AND U44258 ( .A(mul_pow), .B(n41451), .Z(n41450) );
  XOR U44259 ( .A(ein[321]), .B(ein[320]), .Z(n41451) );
  XOR U44260 ( .A(ein[319]), .B(n41452), .Z(ereg_next[320]) );
  AND U44261 ( .A(mul_pow), .B(n41453), .Z(n41452) );
  XOR U44262 ( .A(ein[320]), .B(ein[319]), .Z(n41453) );
  XOR U44263 ( .A(ein[30]), .B(n41454), .Z(ereg_next[31]) );
  AND U44264 ( .A(mul_pow), .B(n41455), .Z(n41454) );
  XOR U44265 ( .A(ein[31]), .B(ein[30]), .Z(n41455) );
  XOR U44266 ( .A(ein[318]), .B(n41456), .Z(ereg_next[319]) );
  AND U44267 ( .A(mul_pow), .B(n41457), .Z(n41456) );
  XOR U44268 ( .A(ein[319]), .B(ein[318]), .Z(n41457) );
  XOR U44269 ( .A(ein[317]), .B(n41458), .Z(ereg_next[318]) );
  AND U44270 ( .A(mul_pow), .B(n41459), .Z(n41458) );
  XOR U44271 ( .A(ein[318]), .B(ein[317]), .Z(n41459) );
  XOR U44272 ( .A(ein[316]), .B(n41460), .Z(ereg_next[317]) );
  AND U44273 ( .A(mul_pow), .B(n41461), .Z(n41460) );
  XOR U44274 ( .A(ein[317]), .B(ein[316]), .Z(n41461) );
  XOR U44275 ( .A(ein[315]), .B(n41462), .Z(ereg_next[316]) );
  AND U44276 ( .A(mul_pow), .B(n41463), .Z(n41462) );
  XOR U44277 ( .A(ein[316]), .B(ein[315]), .Z(n41463) );
  XOR U44278 ( .A(ein[314]), .B(n41464), .Z(ereg_next[315]) );
  AND U44279 ( .A(mul_pow), .B(n41465), .Z(n41464) );
  XOR U44280 ( .A(ein[315]), .B(ein[314]), .Z(n41465) );
  XOR U44281 ( .A(ein[313]), .B(n41466), .Z(ereg_next[314]) );
  AND U44282 ( .A(mul_pow), .B(n41467), .Z(n41466) );
  XOR U44283 ( .A(ein[314]), .B(ein[313]), .Z(n41467) );
  XOR U44284 ( .A(ein[312]), .B(n41468), .Z(ereg_next[313]) );
  AND U44285 ( .A(mul_pow), .B(n41469), .Z(n41468) );
  XOR U44286 ( .A(ein[313]), .B(ein[312]), .Z(n41469) );
  XOR U44287 ( .A(ein[311]), .B(n41470), .Z(ereg_next[312]) );
  AND U44288 ( .A(mul_pow), .B(n41471), .Z(n41470) );
  XOR U44289 ( .A(ein[312]), .B(ein[311]), .Z(n41471) );
  XOR U44290 ( .A(ein[310]), .B(n41472), .Z(ereg_next[311]) );
  AND U44291 ( .A(mul_pow), .B(n41473), .Z(n41472) );
  XOR U44292 ( .A(ein[311]), .B(ein[310]), .Z(n41473) );
  XOR U44293 ( .A(ein[309]), .B(n41474), .Z(ereg_next[310]) );
  AND U44294 ( .A(mul_pow), .B(n41475), .Z(n41474) );
  XOR U44295 ( .A(ein[310]), .B(ein[309]), .Z(n41475) );
  XOR U44296 ( .A(ein[29]), .B(n41476), .Z(ereg_next[30]) );
  AND U44297 ( .A(mul_pow), .B(n41477), .Z(n41476) );
  XOR U44298 ( .A(ein[30]), .B(ein[29]), .Z(n41477) );
  XOR U44299 ( .A(ein[308]), .B(n41478), .Z(ereg_next[309]) );
  AND U44300 ( .A(mul_pow), .B(n41479), .Z(n41478) );
  XOR U44301 ( .A(ein[309]), .B(ein[308]), .Z(n41479) );
  XOR U44302 ( .A(ein[307]), .B(n41480), .Z(ereg_next[308]) );
  AND U44303 ( .A(mul_pow), .B(n41481), .Z(n41480) );
  XOR U44304 ( .A(ein[308]), .B(ein[307]), .Z(n41481) );
  XOR U44305 ( .A(ein[306]), .B(n41482), .Z(ereg_next[307]) );
  AND U44306 ( .A(mul_pow), .B(n41483), .Z(n41482) );
  XOR U44307 ( .A(ein[307]), .B(ein[306]), .Z(n41483) );
  XOR U44308 ( .A(ein[305]), .B(n41484), .Z(ereg_next[306]) );
  AND U44309 ( .A(mul_pow), .B(n41485), .Z(n41484) );
  XOR U44310 ( .A(ein[306]), .B(ein[305]), .Z(n41485) );
  XOR U44311 ( .A(ein[304]), .B(n41486), .Z(ereg_next[305]) );
  AND U44312 ( .A(mul_pow), .B(n41487), .Z(n41486) );
  XOR U44313 ( .A(ein[305]), .B(ein[304]), .Z(n41487) );
  XOR U44314 ( .A(ein[303]), .B(n41488), .Z(ereg_next[304]) );
  AND U44315 ( .A(mul_pow), .B(n41489), .Z(n41488) );
  XOR U44316 ( .A(ein[304]), .B(ein[303]), .Z(n41489) );
  XOR U44317 ( .A(ein[302]), .B(n41490), .Z(ereg_next[303]) );
  AND U44318 ( .A(mul_pow), .B(n41491), .Z(n41490) );
  XOR U44319 ( .A(ein[303]), .B(ein[302]), .Z(n41491) );
  XOR U44320 ( .A(ein[301]), .B(n41492), .Z(ereg_next[302]) );
  AND U44321 ( .A(mul_pow), .B(n41493), .Z(n41492) );
  XOR U44322 ( .A(ein[302]), .B(ein[301]), .Z(n41493) );
  XOR U44323 ( .A(ein[300]), .B(n41494), .Z(ereg_next[301]) );
  AND U44324 ( .A(mul_pow), .B(n41495), .Z(n41494) );
  XOR U44325 ( .A(ein[301]), .B(ein[300]), .Z(n41495) );
  XOR U44326 ( .A(ein[299]), .B(n41496), .Z(ereg_next[300]) );
  AND U44327 ( .A(mul_pow), .B(n41497), .Z(n41496) );
  XOR U44328 ( .A(ein[300]), .B(ein[299]), .Z(n41497) );
  XOR U44329 ( .A(ein[1]), .B(n41498), .Z(ereg_next[2]) );
  AND U44330 ( .A(mul_pow), .B(n41499), .Z(n41498) );
  XOR U44331 ( .A(ein[2]), .B(ein[1]), .Z(n41499) );
  XOR U44332 ( .A(ein[28]), .B(n41500), .Z(ereg_next[29]) );
  AND U44333 ( .A(mul_pow), .B(n41501), .Z(n41500) );
  XOR U44334 ( .A(ein[29]), .B(ein[28]), .Z(n41501) );
  XOR U44335 ( .A(ein[298]), .B(n41502), .Z(ereg_next[299]) );
  AND U44336 ( .A(mul_pow), .B(n41503), .Z(n41502) );
  XOR U44337 ( .A(ein[299]), .B(ein[298]), .Z(n41503) );
  XOR U44338 ( .A(ein[297]), .B(n41504), .Z(ereg_next[298]) );
  AND U44339 ( .A(mul_pow), .B(n41505), .Z(n41504) );
  XOR U44340 ( .A(ein[298]), .B(ein[297]), .Z(n41505) );
  XOR U44341 ( .A(ein[296]), .B(n41506), .Z(ereg_next[297]) );
  AND U44342 ( .A(mul_pow), .B(n41507), .Z(n41506) );
  XOR U44343 ( .A(ein[297]), .B(ein[296]), .Z(n41507) );
  XOR U44344 ( .A(ein[295]), .B(n41508), .Z(ereg_next[296]) );
  AND U44345 ( .A(mul_pow), .B(n41509), .Z(n41508) );
  XOR U44346 ( .A(ein[296]), .B(ein[295]), .Z(n41509) );
  XOR U44347 ( .A(ein[294]), .B(n41510), .Z(ereg_next[295]) );
  AND U44348 ( .A(mul_pow), .B(n41511), .Z(n41510) );
  XOR U44349 ( .A(ein[295]), .B(ein[294]), .Z(n41511) );
  XOR U44350 ( .A(ein[293]), .B(n41512), .Z(ereg_next[294]) );
  AND U44351 ( .A(mul_pow), .B(n41513), .Z(n41512) );
  XOR U44352 ( .A(ein[294]), .B(ein[293]), .Z(n41513) );
  XOR U44353 ( .A(ein[292]), .B(n41514), .Z(ereg_next[293]) );
  AND U44354 ( .A(mul_pow), .B(n41515), .Z(n41514) );
  XOR U44355 ( .A(ein[293]), .B(ein[292]), .Z(n41515) );
  XOR U44356 ( .A(ein[291]), .B(n41516), .Z(ereg_next[292]) );
  AND U44357 ( .A(mul_pow), .B(n41517), .Z(n41516) );
  XOR U44358 ( .A(ein[292]), .B(ein[291]), .Z(n41517) );
  XOR U44359 ( .A(ein[290]), .B(n41518), .Z(ereg_next[291]) );
  AND U44360 ( .A(mul_pow), .B(n41519), .Z(n41518) );
  XOR U44361 ( .A(ein[291]), .B(ein[290]), .Z(n41519) );
  XOR U44362 ( .A(ein[289]), .B(n41520), .Z(ereg_next[290]) );
  AND U44363 ( .A(mul_pow), .B(n41521), .Z(n41520) );
  XOR U44364 ( .A(ein[290]), .B(ein[289]), .Z(n41521) );
  XOR U44365 ( .A(ein[27]), .B(n41522), .Z(ereg_next[28]) );
  AND U44366 ( .A(mul_pow), .B(n41523), .Z(n41522) );
  XOR U44367 ( .A(ein[28]), .B(ein[27]), .Z(n41523) );
  XOR U44368 ( .A(ein[288]), .B(n41524), .Z(ereg_next[289]) );
  AND U44369 ( .A(mul_pow), .B(n41525), .Z(n41524) );
  XOR U44370 ( .A(ein[289]), .B(ein[288]), .Z(n41525) );
  XOR U44371 ( .A(ein[287]), .B(n41526), .Z(ereg_next[288]) );
  AND U44372 ( .A(mul_pow), .B(n41527), .Z(n41526) );
  XOR U44373 ( .A(ein[288]), .B(ein[287]), .Z(n41527) );
  XOR U44374 ( .A(ein[286]), .B(n41528), .Z(ereg_next[287]) );
  AND U44375 ( .A(mul_pow), .B(n41529), .Z(n41528) );
  XOR U44376 ( .A(ein[287]), .B(ein[286]), .Z(n41529) );
  XOR U44377 ( .A(ein[285]), .B(n41530), .Z(ereg_next[286]) );
  AND U44378 ( .A(mul_pow), .B(n41531), .Z(n41530) );
  XOR U44379 ( .A(ein[286]), .B(ein[285]), .Z(n41531) );
  XOR U44380 ( .A(ein[284]), .B(n41532), .Z(ereg_next[285]) );
  AND U44381 ( .A(mul_pow), .B(n41533), .Z(n41532) );
  XOR U44382 ( .A(ein[285]), .B(ein[284]), .Z(n41533) );
  XOR U44383 ( .A(ein[283]), .B(n41534), .Z(ereg_next[284]) );
  AND U44384 ( .A(mul_pow), .B(n41535), .Z(n41534) );
  XOR U44385 ( .A(ein[284]), .B(ein[283]), .Z(n41535) );
  XOR U44386 ( .A(ein[282]), .B(n41536), .Z(ereg_next[283]) );
  AND U44387 ( .A(mul_pow), .B(n41537), .Z(n41536) );
  XOR U44388 ( .A(ein[283]), .B(ein[282]), .Z(n41537) );
  XOR U44389 ( .A(ein[281]), .B(n41538), .Z(ereg_next[282]) );
  AND U44390 ( .A(mul_pow), .B(n41539), .Z(n41538) );
  XOR U44391 ( .A(ein[282]), .B(ein[281]), .Z(n41539) );
  XOR U44392 ( .A(ein[280]), .B(n41540), .Z(ereg_next[281]) );
  AND U44393 ( .A(mul_pow), .B(n41541), .Z(n41540) );
  XOR U44394 ( .A(ein[281]), .B(ein[280]), .Z(n41541) );
  XOR U44395 ( .A(ein[279]), .B(n41542), .Z(ereg_next[280]) );
  AND U44396 ( .A(mul_pow), .B(n41543), .Z(n41542) );
  XOR U44397 ( .A(ein[280]), .B(ein[279]), .Z(n41543) );
  XOR U44398 ( .A(ein[26]), .B(n41544), .Z(ereg_next[27]) );
  AND U44399 ( .A(mul_pow), .B(n41545), .Z(n41544) );
  XOR U44400 ( .A(ein[27]), .B(ein[26]), .Z(n41545) );
  XOR U44401 ( .A(ein[278]), .B(n41546), .Z(ereg_next[279]) );
  AND U44402 ( .A(mul_pow), .B(n41547), .Z(n41546) );
  XOR U44403 ( .A(ein[279]), .B(ein[278]), .Z(n41547) );
  XOR U44404 ( .A(ein[277]), .B(n41548), .Z(ereg_next[278]) );
  AND U44405 ( .A(mul_pow), .B(n41549), .Z(n41548) );
  XOR U44406 ( .A(ein[278]), .B(ein[277]), .Z(n41549) );
  XOR U44407 ( .A(ein[276]), .B(n41550), .Z(ereg_next[277]) );
  AND U44408 ( .A(mul_pow), .B(n41551), .Z(n41550) );
  XOR U44409 ( .A(ein[277]), .B(ein[276]), .Z(n41551) );
  XOR U44410 ( .A(ein[275]), .B(n41552), .Z(ereg_next[276]) );
  AND U44411 ( .A(mul_pow), .B(n41553), .Z(n41552) );
  XOR U44412 ( .A(ein[276]), .B(ein[275]), .Z(n41553) );
  XOR U44413 ( .A(ein[274]), .B(n41554), .Z(ereg_next[275]) );
  AND U44414 ( .A(mul_pow), .B(n41555), .Z(n41554) );
  XOR U44415 ( .A(ein[275]), .B(ein[274]), .Z(n41555) );
  XOR U44416 ( .A(ein[273]), .B(n41556), .Z(ereg_next[274]) );
  AND U44417 ( .A(mul_pow), .B(n41557), .Z(n41556) );
  XOR U44418 ( .A(ein[274]), .B(ein[273]), .Z(n41557) );
  XOR U44419 ( .A(ein[272]), .B(n41558), .Z(ereg_next[273]) );
  AND U44420 ( .A(mul_pow), .B(n41559), .Z(n41558) );
  XOR U44421 ( .A(ein[273]), .B(ein[272]), .Z(n41559) );
  XOR U44422 ( .A(ein[271]), .B(n41560), .Z(ereg_next[272]) );
  AND U44423 ( .A(mul_pow), .B(n41561), .Z(n41560) );
  XOR U44424 ( .A(ein[272]), .B(ein[271]), .Z(n41561) );
  XOR U44425 ( .A(ein[270]), .B(n41562), .Z(ereg_next[271]) );
  AND U44426 ( .A(mul_pow), .B(n41563), .Z(n41562) );
  XOR U44427 ( .A(ein[271]), .B(ein[270]), .Z(n41563) );
  XOR U44428 ( .A(ein[269]), .B(n41564), .Z(ereg_next[270]) );
  AND U44429 ( .A(mul_pow), .B(n41565), .Z(n41564) );
  XOR U44430 ( .A(ein[270]), .B(ein[269]), .Z(n41565) );
  XOR U44431 ( .A(ein[25]), .B(n41566), .Z(ereg_next[26]) );
  AND U44432 ( .A(mul_pow), .B(n41567), .Z(n41566) );
  XOR U44433 ( .A(ein[26]), .B(ein[25]), .Z(n41567) );
  XOR U44434 ( .A(ein[268]), .B(n41568), .Z(ereg_next[269]) );
  AND U44435 ( .A(mul_pow), .B(n41569), .Z(n41568) );
  XOR U44436 ( .A(ein[269]), .B(ein[268]), .Z(n41569) );
  XOR U44437 ( .A(ein[267]), .B(n41570), .Z(ereg_next[268]) );
  AND U44438 ( .A(mul_pow), .B(n41571), .Z(n41570) );
  XOR U44439 ( .A(ein[268]), .B(ein[267]), .Z(n41571) );
  XOR U44440 ( .A(ein[266]), .B(n41572), .Z(ereg_next[267]) );
  AND U44441 ( .A(mul_pow), .B(n41573), .Z(n41572) );
  XOR U44442 ( .A(ein[267]), .B(ein[266]), .Z(n41573) );
  XOR U44443 ( .A(ein[265]), .B(n41574), .Z(ereg_next[266]) );
  AND U44444 ( .A(mul_pow), .B(n41575), .Z(n41574) );
  XOR U44445 ( .A(ein[266]), .B(ein[265]), .Z(n41575) );
  XOR U44446 ( .A(ein[264]), .B(n41576), .Z(ereg_next[265]) );
  AND U44447 ( .A(mul_pow), .B(n41577), .Z(n41576) );
  XOR U44448 ( .A(ein[265]), .B(ein[264]), .Z(n41577) );
  XOR U44449 ( .A(ein[263]), .B(n41578), .Z(ereg_next[264]) );
  AND U44450 ( .A(mul_pow), .B(n41579), .Z(n41578) );
  XOR U44451 ( .A(ein[264]), .B(ein[263]), .Z(n41579) );
  XOR U44452 ( .A(ein[262]), .B(n41580), .Z(ereg_next[263]) );
  AND U44453 ( .A(mul_pow), .B(n41581), .Z(n41580) );
  XOR U44454 ( .A(ein[263]), .B(ein[262]), .Z(n41581) );
  XOR U44455 ( .A(ein[261]), .B(n41582), .Z(ereg_next[262]) );
  AND U44456 ( .A(mul_pow), .B(n41583), .Z(n41582) );
  XOR U44457 ( .A(ein[262]), .B(ein[261]), .Z(n41583) );
  XOR U44458 ( .A(ein[260]), .B(n41584), .Z(ereg_next[261]) );
  AND U44459 ( .A(mul_pow), .B(n41585), .Z(n41584) );
  XOR U44460 ( .A(ein[261]), .B(ein[260]), .Z(n41585) );
  XOR U44461 ( .A(ein[259]), .B(n41586), .Z(ereg_next[260]) );
  AND U44462 ( .A(mul_pow), .B(n41587), .Z(n41586) );
  XOR U44463 ( .A(ein[260]), .B(ein[259]), .Z(n41587) );
  XOR U44464 ( .A(ein[24]), .B(n41588), .Z(ereg_next[25]) );
  AND U44465 ( .A(mul_pow), .B(n41589), .Z(n41588) );
  XOR U44466 ( .A(ein[25]), .B(ein[24]), .Z(n41589) );
  XOR U44467 ( .A(ein[258]), .B(n41590), .Z(ereg_next[259]) );
  AND U44468 ( .A(mul_pow), .B(n41591), .Z(n41590) );
  XOR U44469 ( .A(ein[259]), .B(ein[258]), .Z(n41591) );
  XOR U44470 ( .A(ein[257]), .B(n41592), .Z(ereg_next[258]) );
  AND U44471 ( .A(mul_pow), .B(n41593), .Z(n41592) );
  XOR U44472 ( .A(ein[258]), .B(ein[257]), .Z(n41593) );
  XOR U44473 ( .A(ein[256]), .B(n41594), .Z(ereg_next[257]) );
  AND U44474 ( .A(mul_pow), .B(n41595), .Z(n41594) );
  XOR U44475 ( .A(ein[257]), .B(ein[256]), .Z(n41595) );
  XOR U44476 ( .A(ein[255]), .B(n41596), .Z(ereg_next[256]) );
  AND U44477 ( .A(mul_pow), .B(n41597), .Z(n41596) );
  XOR U44478 ( .A(ein[256]), .B(ein[255]), .Z(n41597) );
  XOR U44479 ( .A(ein[254]), .B(n41598), .Z(ereg_next[255]) );
  AND U44480 ( .A(mul_pow), .B(n41599), .Z(n41598) );
  XOR U44481 ( .A(ein[255]), .B(ein[254]), .Z(n41599) );
  XOR U44482 ( .A(ein[253]), .B(n41600), .Z(ereg_next[254]) );
  AND U44483 ( .A(mul_pow), .B(n41601), .Z(n41600) );
  XOR U44484 ( .A(ein[254]), .B(ein[253]), .Z(n41601) );
  XOR U44485 ( .A(ein[252]), .B(n41602), .Z(ereg_next[253]) );
  AND U44486 ( .A(mul_pow), .B(n41603), .Z(n41602) );
  XOR U44487 ( .A(ein[253]), .B(ein[252]), .Z(n41603) );
  XOR U44488 ( .A(ein[251]), .B(n41604), .Z(ereg_next[252]) );
  AND U44489 ( .A(mul_pow), .B(n41605), .Z(n41604) );
  XOR U44490 ( .A(ein[252]), .B(ein[251]), .Z(n41605) );
  XOR U44491 ( .A(ein[250]), .B(n41606), .Z(ereg_next[251]) );
  AND U44492 ( .A(mul_pow), .B(n41607), .Z(n41606) );
  XOR U44493 ( .A(ein[251]), .B(ein[250]), .Z(n41607) );
  XOR U44494 ( .A(ein[249]), .B(n41608), .Z(ereg_next[250]) );
  AND U44495 ( .A(mul_pow), .B(n41609), .Z(n41608) );
  XOR U44496 ( .A(ein[250]), .B(ein[249]), .Z(n41609) );
  XOR U44497 ( .A(ein[23]), .B(n41610), .Z(ereg_next[24]) );
  AND U44498 ( .A(mul_pow), .B(n41611), .Z(n41610) );
  XOR U44499 ( .A(ein[24]), .B(ein[23]), .Z(n41611) );
  XOR U44500 ( .A(ein[248]), .B(n41612), .Z(ereg_next[249]) );
  AND U44501 ( .A(mul_pow), .B(n41613), .Z(n41612) );
  XOR U44502 ( .A(ein[249]), .B(ein[248]), .Z(n41613) );
  XOR U44503 ( .A(ein[247]), .B(n41614), .Z(ereg_next[248]) );
  AND U44504 ( .A(mul_pow), .B(n41615), .Z(n41614) );
  XOR U44505 ( .A(ein[248]), .B(ein[247]), .Z(n41615) );
  XOR U44506 ( .A(ein[246]), .B(n41616), .Z(ereg_next[247]) );
  AND U44507 ( .A(mul_pow), .B(n41617), .Z(n41616) );
  XOR U44508 ( .A(ein[247]), .B(ein[246]), .Z(n41617) );
  XOR U44509 ( .A(ein[245]), .B(n41618), .Z(ereg_next[246]) );
  AND U44510 ( .A(mul_pow), .B(n41619), .Z(n41618) );
  XOR U44511 ( .A(ein[246]), .B(ein[245]), .Z(n41619) );
  XOR U44512 ( .A(ein[244]), .B(n41620), .Z(ereg_next[245]) );
  AND U44513 ( .A(mul_pow), .B(n41621), .Z(n41620) );
  XOR U44514 ( .A(ein[245]), .B(ein[244]), .Z(n41621) );
  XOR U44515 ( .A(ein[243]), .B(n41622), .Z(ereg_next[244]) );
  AND U44516 ( .A(mul_pow), .B(n41623), .Z(n41622) );
  XOR U44517 ( .A(ein[244]), .B(ein[243]), .Z(n41623) );
  XOR U44518 ( .A(ein[242]), .B(n41624), .Z(ereg_next[243]) );
  AND U44519 ( .A(mul_pow), .B(n41625), .Z(n41624) );
  XOR U44520 ( .A(ein[243]), .B(ein[242]), .Z(n41625) );
  XOR U44521 ( .A(ein[241]), .B(n41626), .Z(ereg_next[242]) );
  AND U44522 ( .A(mul_pow), .B(n41627), .Z(n41626) );
  XOR U44523 ( .A(ein[242]), .B(ein[241]), .Z(n41627) );
  XOR U44524 ( .A(ein[240]), .B(n41628), .Z(ereg_next[241]) );
  AND U44525 ( .A(mul_pow), .B(n41629), .Z(n41628) );
  XOR U44526 ( .A(ein[241]), .B(ein[240]), .Z(n41629) );
  XOR U44527 ( .A(ein[239]), .B(n41630), .Z(ereg_next[240]) );
  AND U44528 ( .A(mul_pow), .B(n41631), .Z(n41630) );
  XOR U44529 ( .A(ein[240]), .B(ein[239]), .Z(n41631) );
  XOR U44530 ( .A(ein[22]), .B(n41632), .Z(ereg_next[23]) );
  AND U44531 ( .A(mul_pow), .B(n41633), .Z(n41632) );
  XOR U44532 ( .A(ein[23]), .B(ein[22]), .Z(n41633) );
  XOR U44533 ( .A(ein[238]), .B(n41634), .Z(ereg_next[239]) );
  AND U44534 ( .A(mul_pow), .B(n41635), .Z(n41634) );
  XOR U44535 ( .A(ein[239]), .B(ein[238]), .Z(n41635) );
  XOR U44536 ( .A(ein[237]), .B(n41636), .Z(ereg_next[238]) );
  AND U44537 ( .A(mul_pow), .B(n41637), .Z(n41636) );
  XOR U44538 ( .A(ein[238]), .B(ein[237]), .Z(n41637) );
  XOR U44539 ( .A(ein[236]), .B(n41638), .Z(ereg_next[237]) );
  AND U44540 ( .A(mul_pow), .B(n41639), .Z(n41638) );
  XOR U44541 ( .A(ein[237]), .B(ein[236]), .Z(n41639) );
  XOR U44542 ( .A(ein[235]), .B(n41640), .Z(ereg_next[236]) );
  AND U44543 ( .A(mul_pow), .B(n41641), .Z(n41640) );
  XOR U44544 ( .A(ein[236]), .B(ein[235]), .Z(n41641) );
  XOR U44545 ( .A(ein[234]), .B(n41642), .Z(ereg_next[235]) );
  AND U44546 ( .A(mul_pow), .B(n41643), .Z(n41642) );
  XOR U44547 ( .A(ein[235]), .B(ein[234]), .Z(n41643) );
  XOR U44548 ( .A(ein[233]), .B(n41644), .Z(ereg_next[234]) );
  AND U44549 ( .A(mul_pow), .B(n41645), .Z(n41644) );
  XOR U44550 ( .A(ein[234]), .B(ein[233]), .Z(n41645) );
  XOR U44551 ( .A(ein[232]), .B(n41646), .Z(ereg_next[233]) );
  AND U44552 ( .A(mul_pow), .B(n41647), .Z(n41646) );
  XOR U44553 ( .A(ein[233]), .B(ein[232]), .Z(n41647) );
  XOR U44554 ( .A(ein[231]), .B(n41648), .Z(ereg_next[232]) );
  AND U44555 ( .A(mul_pow), .B(n41649), .Z(n41648) );
  XOR U44556 ( .A(ein[232]), .B(ein[231]), .Z(n41649) );
  XOR U44557 ( .A(ein[230]), .B(n41650), .Z(ereg_next[231]) );
  AND U44558 ( .A(mul_pow), .B(n41651), .Z(n41650) );
  XOR U44559 ( .A(ein[231]), .B(ein[230]), .Z(n41651) );
  XOR U44560 ( .A(ein[229]), .B(n41652), .Z(ereg_next[230]) );
  AND U44561 ( .A(mul_pow), .B(n41653), .Z(n41652) );
  XOR U44562 ( .A(ein[230]), .B(ein[229]), .Z(n41653) );
  XOR U44563 ( .A(ein[21]), .B(n41654), .Z(ereg_next[22]) );
  AND U44564 ( .A(mul_pow), .B(n41655), .Z(n41654) );
  XOR U44565 ( .A(ein[22]), .B(ein[21]), .Z(n41655) );
  XOR U44566 ( .A(ein[228]), .B(n41656), .Z(ereg_next[229]) );
  AND U44567 ( .A(mul_pow), .B(n41657), .Z(n41656) );
  XOR U44568 ( .A(ein[229]), .B(ein[228]), .Z(n41657) );
  XOR U44569 ( .A(ein[227]), .B(n41658), .Z(ereg_next[228]) );
  AND U44570 ( .A(mul_pow), .B(n41659), .Z(n41658) );
  XOR U44571 ( .A(ein[228]), .B(ein[227]), .Z(n41659) );
  XOR U44572 ( .A(ein[226]), .B(n41660), .Z(ereg_next[227]) );
  AND U44573 ( .A(mul_pow), .B(n41661), .Z(n41660) );
  XOR U44574 ( .A(ein[227]), .B(ein[226]), .Z(n41661) );
  XOR U44575 ( .A(ein[225]), .B(n41662), .Z(ereg_next[226]) );
  AND U44576 ( .A(mul_pow), .B(n41663), .Z(n41662) );
  XOR U44577 ( .A(ein[226]), .B(ein[225]), .Z(n41663) );
  XOR U44578 ( .A(ein[224]), .B(n41664), .Z(ereg_next[225]) );
  AND U44579 ( .A(mul_pow), .B(n41665), .Z(n41664) );
  XOR U44580 ( .A(ein[225]), .B(ein[224]), .Z(n41665) );
  XOR U44581 ( .A(ein[223]), .B(n41666), .Z(ereg_next[224]) );
  AND U44582 ( .A(mul_pow), .B(n41667), .Z(n41666) );
  XOR U44583 ( .A(ein[224]), .B(ein[223]), .Z(n41667) );
  XOR U44584 ( .A(ein[222]), .B(n41668), .Z(ereg_next[223]) );
  AND U44585 ( .A(mul_pow), .B(n41669), .Z(n41668) );
  XOR U44586 ( .A(ein[223]), .B(ein[222]), .Z(n41669) );
  XOR U44587 ( .A(ein[221]), .B(n41670), .Z(ereg_next[222]) );
  AND U44588 ( .A(mul_pow), .B(n41671), .Z(n41670) );
  XOR U44589 ( .A(ein[222]), .B(ein[221]), .Z(n41671) );
  XOR U44590 ( .A(ein[220]), .B(n41672), .Z(ereg_next[221]) );
  AND U44591 ( .A(mul_pow), .B(n41673), .Z(n41672) );
  XOR U44592 ( .A(ein[221]), .B(ein[220]), .Z(n41673) );
  XOR U44593 ( .A(ein[219]), .B(n41674), .Z(ereg_next[220]) );
  AND U44594 ( .A(mul_pow), .B(n41675), .Z(n41674) );
  XOR U44595 ( .A(ein[220]), .B(ein[219]), .Z(n41675) );
  XOR U44596 ( .A(ein[20]), .B(n41676), .Z(ereg_next[21]) );
  AND U44597 ( .A(mul_pow), .B(n41677), .Z(n41676) );
  XOR U44598 ( .A(ein[21]), .B(ein[20]), .Z(n41677) );
  XOR U44599 ( .A(ein[218]), .B(n41678), .Z(ereg_next[219]) );
  AND U44600 ( .A(mul_pow), .B(n41679), .Z(n41678) );
  XOR U44601 ( .A(ein[219]), .B(ein[218]), .Z(n41679) );
  XOR U44602 ( .A(ein[217]), .B(n41680), .Z(ereg_next[218]) );
  AND U44603 ( .A(mul_pow), .B(n41681), .Z(n41680) );
  XOR U44604 ( .A(ein[218]), .B(ein[217]), .Z(n41681) );
  XOR U44605 ( .A(ein[216]), .B(n41682), .Z(ereg_next[217]) );
  AND U44606 ( .A(mul_pow), .B(n41683), .Z(n41682) );
  XOR U44607 ( .A(ein[217]), .B(ein[216]), .Z(n41683) );
  XOR U44608 ( .A(ein[215]), .B(n41684), .Z(ereg_next[216]) );
  AND U44609 ( .A(mul_pow), .B(n41685), .Z(n41684) );
  XOR U44610 ( .A(ein[216]), .B(ein[215]), .Z(n41685) );
  XOR U44611 ( .A(ein[214]), .B(n41686), .Z(ereg_next[215]) );
  AND U44612 ( .A(mul_pow), .B(n41687), .Z(n41686) );
  XOR U44613 ( .A(ein[215]), .B(ein[214]), .Z(n41687) );
  XOR U44614 ( .A(ein[213]), .B(n41688), .Z(ereg_next[214]) );
  AND U44615 ( .A(mul_pow), .B(n41689), .Z(n41688) );
  XOR U44616 ( .A(ein[214]), .B(ein[213]), .Z(n41689) );
  XOR U44617 ( .A(ein[212]), .B(n41690), .Z(ereg_next[213]) );
  AND U44618 ( .A(mul_pow), .B(n41691), .Z(n41690) );
  XOR U44619 ( .A(ein[213]), .B(ein[212]), .Z(n41691) );
  XOR U44620 ( .A(ein[211]), .B(n41692), .Z(ereg_next[212]) );
  AND U44621 ( .A(mul_pow), .B(n41693), .Z(n41692) );
  XOR U44622 ( .A(ein[212]), .B(ein[211]), .Z(n41693) );
  XOR U44623 ( .A(ein[210]), .B(n41694), .Z(ereg_next[211]) );
  AND U44624 ( .A(mul_pow), .B(n41695), .Z(n41694) );
  XOR U44625 ( .A(ein[211]), .B(ein[210]), .Z(n41695) );
  XOR U44626 ( .A(ein[209]), .B(n41696), .Z(ereg_next[210]) );
  AND U44627 ( .A(mul_pow), .B(n41697), .Z(n41696) );
  XOR U44628 ( .A(ein[210]), .B(ein[209]), .Z(n41697) );
  XOR U44629 ( .A(ein[19]), .B(n41698), .Z(ereg_next[20]) );
  AND U44630 ( .A(mul_pow), .B(n41699), .Z(n41698) );
  XOR U44631 ( .A(ein[20]), .B(ein[19]), .Z(n41699) );
  XOR U44632 ( .A(ein[208]), .B(n41700), .Z(ereg_next[209]) );
  AND U44633 ( .A(mul_pow), .B(n41701), .Z(n41700) );
  XOR U44634 ( .A(ein[209]), .B(ein[208]), .Z(n41701) );
  XOR U44635 ( .A(ein[207]), .B(n41702), .Z(ereg_next[208]) );
  AND U44636 ( .A(mul_pow), .B(n41703), .Z(n41702) );
  XOR U44637 ( .A(ein[208]), .B(ein[207]), .Z(n41703) );
  XOR U44638 ( .A(ein[206]), .B(n41704), .Z(ereg_next[207]) );
  AND U44639 ( .A(mul_pow), .B(n41705), .Z(n41704) );
  XOR U44640 ( .A(ein[207]), .B(ein[206]), .Z(n41705) );
  XOR U44641 ( .A(ein[205]), .B(n41706), .Z(ereg_next[206]) );
  AND U44642 ( .A(mul_pow), .B(n41707), .Z(n41706) );
  XOR U44643 ( .A(ein[206]), .B(ein[205]), .Z(n41707) );
  XOR U44644 ( .A(ein[204]), .B(n41708), .Z(ereg_next[205]) );
  AND U44645 ( .A(mul_pow), .B(n41709), .Z(n41708) );
  XOR U44646 ( .A(ein[205]), .B(ein[204]), .Z(n41709) );
  XOR U44647 ( .A(ein[203]), .B(n41710), .Z(ereg_next[204]) );
  AND U44648 ( .A(mul_pow), .B(n41711), .Z(n41710) );
  XOR U44649 ( .A(ein[204]), .B(ein[203]), .Z(n41711) );
  XOR U44650 ( .A(ein[202]), .B(n41712), .Z(ereg_next[203]) );
  AND U44651 ( .A(mul_pow), .B(n41713), .Z(n41712) );
  XOR U44652 ( .A(ein[203]), .B(ein[202]), .Z(n41713) );
  XOR U44653 ( .A(ein[201]), .B(n41714), .Z(ereg_next[202]) );
  AND U44654 ( .A(mul_pow), .B(n41715), .Z(n41714) );
  XOR U44655 ( .A(ein[202]), .B(ein[201]), .Z(n41715) );
  XOR U44656 ( .A(ein[200]), .B(n41716), .Z(ereg_next[201]) );
  AND U44657 ( .A(mul_pow), .B(n41717), .Z(n41716) );
  XOR U44658 ( .A(ein[201]), .B(ein[200]), .Z(n41717) );
  XOR U44659 ( .A(ein[199]), .B(n41718), .Z(ereg_next[200]) );
  AND U44660 ( .A(mul_pow), .B(n41719), .Z(n41718) );
  XOR U44661 ( .A(ein[200]), .B(ein[199]), .Z(n41719) );
  XOR U44662 ( .A(ein[0]), .B(n41720), .Z(ereg_next[1]) );
  AND U44663 ( .A(mul_pow), .B(n41721), .Z(n41720) );
  XOR U44664 ( .A(ein[1]), .B(ein[0]), .Z(n41721) );
  XOR U44665 ( .A(ein[18]), .B(n41722), .Z(ereg_next[19]) );
  AND U44666 ( .A(mul_pow), .B(n41723), .Z(n41722) );
  XOR U44667 ( .A(ein[19]), .B(ein[18]), .Z(n41723) );
  XOR U44668 ( .A(ein[198]), .B(n41724), .Z(ereg_next[199]) );
  AND U44669 ( .A(mul_pow), .B(n41725), .Z(n41724) );
  XOR U44670 ( .A(ein[199]), .B(ein[198]), .Z(n41725) );
  XOR U44671 ( .A(ein[197]), .B(n41726), .Z(ereg_next[198]) );
  AND U44672 ( .A(mul_pow), .B(n41727), .Z(n41726) );
  XOR U44673 ( .A(ein[198]), .B(ein[197]), .Z(n41727) );
  XOR U44674 ( .A(ein[196]), .B(n41728), .Z(ereg_next[197]) );
  AND U44675 ( .A(mul_pow), .B(n41729), .Z(n41728) );
  XOR U44676 ( .A(ein[197]), .B(ein[196]), .Z(n41729) );
  XOR U44677 ( .A(ein[195]), .B(n41730), .Z(ereg_next[196]) );
  AND U44678 ( .A(mul_pow), .B(n41731), .Z(n41730) );
  XOR U44679 ( .A(ein[196]), .B(ein[195]), .Z(n41731) );
  XOR U44680 ( .A(ein[194]), .B(n41732), .Z(ereg_next[195]) );
  AND U44681 ( .A(mul_pow), .B(n41733), .Z(n41732) );
  XOR U44682 ( .A(ein[195]), .B(ein[194]), .Z(n41733) );
  XOR U44683 ( .A(ein[193]), .B(n41734), .Z(ereg_next[194]) );
  AND U44684 ( .A(mul_pow), .B(n41735), .Z(n41734) );
  XOR U44685 ( .A(ein[194]), .B(ein[193]), .Z(n41735) );
  XOR U44686 ( .A(ein[192]), .B(n41736), .Z(ereg_next[193]) );
  AND U44687 ( .A(mul_pow), .B(n41737), .Z(n41736) );
  XOR U44688 ( .A(ein[193]), .B(ein[192]), .Z(n41737) );
  XOR U44689 ( .A(ein[191]), .B(n41738), .Z(ereg_next[192]) );
  AND U44690 ( .A(mul_pow), .B(n41739), .Z(n41738) );
  XOR U44691 ( .A(ein[192]), .B(ein[191]), .Z(n41739) );
  XOR U44692 ( .A(ein[190]), .B(n41740), .Z(ereg_next[191]) );
  AND U44693 ( .A(mul_pow), .B(n41741), .Z(n41740) );
  XOR U44694 ( .A(ein[191]), .B(ein[190]), .Z(n41741) );
  XOR U44695 ( .A(ein[189]), .B(n41742), .Z(ereg_next[190]) );
  AND U44696 ( .A(mul_pow), .B(n41743), .Z(n41742) );
  XOR U44697 ( .A(ein[190]), .B(ein[189]), .Z(n41743) );
  XOR U44698 ( .A(ein[17]), .B(n41744), .Z(ereg_next[18]) );
  AND U44699 ( .A(mul_pow), .B(n41745), .Z(n41744) );
  XOR U44700 ( .A(ein[18]), .B(ein[17]), .Z(n41745) );
  XOR U44701 ( .A(ein[188]), .B(n41746), .Z(ereg_next[189]) );
  AND U44702 ( .A(mul_pow), .B(n41747), .Z(n41746) );
  XOR U44703 ( .A(ein[189]), .B(ein[188]), .Z(n41747) );
  XOR U44704 ( .A(ein[187]), .B(n41748), .Z(ereg_next[188]) );
  AND U44705 ( .A(mul_pow), .B(n41749), .Z(n41748) );
  XOR U44706 ( .A(ein[188]), .B(ein[187]), .Z(n41749) );
  XOR U44707 ( .A(ein[186]), .B(n41750), .Z(ereg_next[187]) );
  AND U44708 ( .A(mul_pow), .B(n41751), .Z(n41750) );
  XOR U44709 ( .A(ein[187]), .B(ein[186]), .Z(n41751) );
  XOR U44710 ( .A(ein[185]), .B(n41752), .Z(ereg_next[186]) );
  AND U44711 ( .A(mul_pow), .B(n41753), .Z(n41752) );
  XOR U44712 ( .A(ein[186]), .B(ein[185]), .Z(n41753) );
  XOR U44713 ( .A(ein[184]), .B(n41754), .Z(ereg_next[185]) );
  AND U44714 ( .A(mul_pow), .B(n41755), .Z(n41754) );
  XOR U44715 ( .A(ein[185]), .B(ein[184]), .Z(n41755) );
  XOR U44716 ( .A(ein[183]), .B(n41756), .Z(ereg_next[184]) );
  AND U44717 ( .A(mul_pow), .B(n41757), .Z(n41756) );
  XOR U44718 ( .A(ein[184]), .B(ein[183]), .Z(n41757) );
  XOR U44719 ( .A(ein[182]), .B(n41758), .Z(ereg_next[183]) );
  AND U44720 ( .A(mul_pow), .B(n41759), .Z(n41758) );
  XOR U44721 ( .A(ein[183]), .B(ein[182]), .Z(n41759) );
  XOR U44722 ( .A(ein[181]), .B(n41760), .Z(ereg_next[182]) );
  AND U44723 ( .A(mul_pow), .B(n41761), .Z(n41760) );
  XOR U44724 ( .A(ein[182]), .B(ein[181]), .Z(n41761) );
  XOR U44725 ( .A(ein[180]), .B(n41762), .Z(ereg_next[181]) );
  AND U44726 ( .A(mul_pow), .B(n41763), .Z(n41762) );
  XOR U44727 ( .A(ein[181]), .B(ein[180]), .Z(n41763) );
  XOR U44728 ( .A(ein[179]), .B(n41764), .Z(ereg_next[180]) );
  AND U44729 ( .A(mul_pow), .B(n41765), .Z(n41764) );
  XOR U44730 ( .A(ein[180]), .B(ein[179]), .Z(n41765) );
  XOR U44731 ( .A(ein[16]), .B(n41766), .Z(ereg_next[17]) );
  AND U44732 ( .A(mul_pow), .B(n41767), .Z(n41766) );
  XOR U44733 ( .A(ein[17]), .B(ein[16]), .Z(n41767) );
  XOR U44734 ( .A(ein[178]), .B(n41768), .Z(ereg_next[179]) );
  AND U44735 ( .A(mul_pow), .B(n41769), .Z(n41768) );
  XOR U44736 ( .A(ein[179]), .B(ein[178]), .Z(n41769) );
  XOR U44737 ( .A(ein[177]), .B(n41770), .Z(ereg_next[178]) );
  AND U44738 ( .A(mul_pow), .B(n41771), .Z(n41770) );
  XOR U44739 ( .A(ein[178]), .B(ein[177]), .Z(n41771) );
  XOR U44740 ( .A(ein[176]), .B(n41772), .Z(ereg_next[177]) );
  AND U44741 ( .A(mul_pow), .B(n41773), .Z(n41772) );
  XOR U44742 ( .A(ein[177]), .B(ein[176]), .Z(n41773) );
  XOR U44743 ( .A(ein[175]), .B(n41774), .Z(ereg_next[176]) );
  AND U44744 ( .A(mul_pow), .B(n41775), .Z(n41774) );
  XOR U44745 ( .A(ein[176]), .B(ein[175]), .Z(n41775) );
  XOR U44746 ( .A(ein[174]), .B(n41776), .Z(ereg_next[175]) );
  AND U44747 ( .A(mul_pow), .B(n41777), .Z(n41776) );
  XOR U44748 ( .A(ein[175]), .B(ein[174]), .Z(n41777) );
  XOR U44749 ( .A(ein[173]), .B(n41778), .Z(ereg_next[174]) );
  AND U44750 ( .A(mul_pow), .B(n41779), .Z(n41778) );
  XOR U44751 ( .A(ein[174]), .B(ein[173]), .Z(n41779) );
  XOR U44752 ( .A(ein[172]), .B(n41780), .Z(ereg_next[173]) );
  AND U44753 ( .A(mul_pow), .B(n41781), .Z(n41780) );
  XOR U44754 ( .A(ein[173]), .B(ein[172]), .Z(n41781) );
  XOR U44755 ( .A(ein[171]), .B(n41782), .Z(ereg_next[172]) );
  AND U44756 ( .A(mul_pow), .B(n41783), .Z(n41782) );
  XOR U44757 ( .A(ein[172]), .B(ein[171]), .Z(n41783) );
  XOR U44758 ( .A(ein[170]), .B(n41784), .Z(ereg_next[171]) );
  AND U44759 ( .A(mul_pow), .B(n41785), .Z(n41784) );
  XOR U44760 ( .A(ein[171]), .B(ein[170]), .Z(n41785) );
  XOR U44761 ( .A(ein[169]), .B(n41786), .Z(ereg_next[170]) );
  AND U44762 ( .A(mul_pow), .B(n41787), .Z(n41786) );
  XOR U44763 ( .A(ein[170]), .B(ein[169]), .Z(n41787) );
  XOR U44764 ( .A(ein[15]), .B(n41788), .Z(ereg_next[16]) );
  AND U44765 ( .A(mul_pow), .B(n41789), .Z(n41788) );
  XOR U44766 ( .A(ein[16]), .B(ein[15]), .Z(n41789) );
  XOR U44767 ( .A(ein[168]), .B(n41790), .Z(ereg_next[169]) );
  AND U44768 ( .A(mul_pow), .B(n41791), .Z(n41790) );
  XOR U44769 ( .A(ein[169]), .B(ein[168]), .Z(n41791) );
  XOR U44770 ( .A(ein[167]), .B(n41792), .Z(ereg_next[168]) );
  AND U44771 ( .A(mul_pow), .B(n41793), .Z(n41792) );
  XOR U44772 ( .A(ein[168]), .B(ein[167]), .Z(n41793) );
  XOR U44773 ( .A(ein[166]), .B(n41794), .Z(ereg_next[167]) );
  AND U44774 ( .A(mul_pow), .B(n41795), .Z(n41794) );
  XOR U44775 ( .A(ein[167]), .B(ein[166]), .Z(n41795) );
  XOR U44776 ( .A(ein[165]), .B(n41796), .Z(ereg_next[166]) );
  AND U44777 ( .A(mul_pow), .B(n41797), .Z(n41796) );
  XOR U44778 ( .A(ein[166]), .B(ein[165]), .Z(n41797) );
  XOR U44779 ( .A(ein[164]), .B(n41798), .Z(ereg_next[165]) );
  AND U44780 ( .A(mul_pow), .B(n41799), .Z(n41798) );
  XOR U44781 ( .A(ein[165]), .B(ein[164]), .Z(n41799) );
  XOR U44782 ( .A(ein[163]), .B(n41800), .Z(ereg_next[164]) );
  AND U44783 ( .A(mul_pow), .B(n41801), .Z(n41800) );
  XOR U44784 ( .A(ein[164]), .B(ein[163]), .Z(n41801) );
  XOR U44785 ( .A(ein[162]), .B(n41802), .Z(ereg_next[163]) );
  AND U44786 ( .A(mul_pow), .B(n41803), .Z(n41802) );
  XOR U44787 ( .A(ein[163]), .B(ein[162]), .Z(n41803) );
  XOR U44788 ( .A(ein[161]), .B(n41804), .Z(ereg_next[162]) );
  AND U44789 ( .A(mul_pow), .B(n41805), .Z(n41804) );
  XOR U44790 ( .A(ein[162]), .B(ein[161]), .Z(n41805) );
  XOR U44791 ( .A(ein[160]), .B(n41806), .Z(ereg_next[161]) );
  AND U44792 ( .A(mul_pow), .B(n41807), .Z(n41806) );
  XOR U44793 ( .A(ein[161]), .B(ein[160]), .Z(n41807) );
  XOR U44794 ( .A(ein[159]), .B(n41808), .Z(ereg_next[160]) );
  AND U44795 ( .A(mul_pow), .B(n41809), .Z(n41808) );
  XOR U44796 ( .A(ein[160]), .B(ein[159]), .Z(n41809) );
  XOR U44797 ( .A(ein[14]), .B(n41810), .Z(ereg_next[15]) );
  AND U44798 ( .A(mul_pow), .B(n41811), .Z(n41810) );
  XOR U44799 ( .A(ein[15]), .B(ein[14]), .Z(n41811) );
  XOR U44800 ( .A(ein[158]), .B(n41812), .Z(ereg_next[159]) );
  AND U44801 ( .A(mul_pow), .B(n41813), .Z(n41812) );
  XOR U44802 ( .A(ein[159]), .B(ein[158]), .Z(n41813) );
  XOR U44803 ( .A(ein[157]), .B(n41814), .Z(ereg_next[158]) );
  AND U44804 ( .A(mul_pow), .B(n41815), .Z(n41814) );
  XOR U44805 ( .A(ein[158]), .B(ein[157]), .Z(n41815) );
  XOR U44806 ( .A(ein[156]), .B(n41816), .Z(ereg_next[157]) );
  AND U44807 ( .A(mul_pow), .B(n41817), .Z(n41816) );
  XOR U44808 ( .A(ein[157]), .B(ein[156]), .Z(n41817) );
  XOR U44809 ( .A(ein[155]), .B(n41818), .Z(ereg_next[156]) );
  AND U44810 ( .A(mul_pow), .B(n41819), .Z(n41818) );
  XOR U44811 ( .A(ein[156]), .B(ein[155]), .Z(n41819) );
  XOR U44812 ( .A(ein[154]), .B(n41820), .Z(ereg_next[155]) );
  AND U44813 ( .A(mul_pow), .B(n41821), .Z(n41820) );
  XOR U44814 ( .A(ein[155]), .B(ein[154]), .Z(n41821) );
  XOR U44815 ( .A(ein[153]), .B(n41822), .Z(ereg_next[154]) );
  AND U44816 ( .A(mul_pow), .B(n41823), .Z(n41822) );
  XOR U44817 ( .A(ein[154]), .B(ein[153]), .Z(n41823) );
  XOR U44818 ( .A(ein[152]), .B(n41824), .Z(ereg_next[153]) );
  AND U44819 ( .A(mul_pow), .B(n41825), .Z(n41824) );
  XOR U44820 ( .A(ein[153]), .B(ein[152]), .Z(n41825) );
  XOR U44821 ( .A(ein[151]), .B(n41826), .Z(ereg_next[152]) );
  AND U44822 ( .A(mul_pow), .B(n41827), .Z(n41826) );
  XOR U44823 ( .A(ein[152]), .B(ein[151]), .Z(n41827) );
  XOR U44824 ( .A(ein[150]), .B(n41828), .Z(ereg_next[151]) );
  AND U44825 ( .A(mul_pow), .B(n41829), .Z(n41828) );
  XOR U44826 ( .A(ein[151]), .B(ein[150]), .Z(n41829) );
  XOR U44827 ( .A(ein[149]), .B(n41830), .Z(ereg_next[150]) );
  AND U44828 ( .A(mul_pow), .B(n41831), .Z(n41830) );
  XOR U44829 ( .A(ein[150]), .B(ein[149]), .Z(n41831) );
  XOR U44830 ( .A(ein[13]), .B(n41832), .Z(ereg_next[14]) );
  AND U44831 ( .A(mul_pow), .B(n41833), .Z(n41832) );
  XOR U44832 ( .A(ein[14]), .B(ein[13]), .Z(n41833) );
  XOR U44833 ( .A(ein[148]), .B(n41834), .Z(ereg_next[149]) );
  AND U44834 ( .A(mul_pow), .B(n41835), .Z(n41834) );
  XOR U44835 ( .A(ein[149]), .B(ein[148]), .Z(n41835) );
  XOR U44836 ( .A(ein[147]), .B(n41836), .Z(ereg_next[148]) );
  AND U44837 ( .A(mul_pow), .B(n41837), .Z(n41836) );
  XOR U44838 ( .A(ein[148]), .B(ein[147]), .Z(n41837) );
  XOR U44839 ( .A(ein[146]), .B(n41838), .Z(ereg_next[147]) );
  AND U44840 ( .A(mul_pow), .B(n41839), .Z(n41838) );
  XOR U44841 ( .A(ein[147]), .B(ein[146]), .Z(n41839) );
  XOR U44842 ( .A(ein[145]), .B(n41840), .Z(ereg_next[146]) );
  AND U44843 ( .A(mul_pow), .B(n41841), .Z(n41840) );
  XOR U44844 ( .A(ein[146]), .B(ein[145]), .Z(n41841) );
  XOR U44845 ( .A(ein[144]), .B(n41842), .Z(ereg_next[145]) );
  AND U44846 ( .A(mul_pow), .B(n41843), .Z(n41842) );
  XOR U44847 ( .A(ein[145]), .B(ein[144]), .Z(n41843) );
  XOR U44848 ( .A(ein[143]), .B(n41844), .Z(ereg_next[144]) );
  AND U44849 ( .A(mul_pow), .B(n41845), .Z(n41844) );
  XOR U44850 ( .A(ein[144]), .B(ein[143]), .Z(n41845) );
  XOR U44851 ( .A(ein[142]), .B(n41846), .Z(ereg_next[143]) );
  AND U44852 ( .A(mul_pow), .B(n41847), .Z(n41846) );
  XOR U44853 ( .A(ein[143]), .B(ein[142]), .Z(n41847) );
  XOR U44854 ( .A(ein[141]), .B(n41848), .Z(ereg_next[142]) );
  AND U44855 ( .A(mul_pow), .B(n41849), .Z(n41848) );
  XOR U44856 ( .A(ein[142]), .B(ein[141]), .Z(n41849) );
  XOR U44857 ( .A(ein[140]), .B(n41850), .Z(ereg_next[141]) );
  AND U44858 ( .A(mul_pow), .B(n41851), .Z(n41850) );
  XOR U44859 ( .A(ein[141]), .B(ein[140]), .Z(n41851) );
  XOR U44860 ( .A(ein[139]), .B(n41852), .Z(ereg_next[140]) );
  AND U44861 ( .A(mul_pow), .B(n41853), .Z(n41852) );
  XOR U44862 ( .A(ein[140]), .B(ein[139]), .Z(n41853) );
  XOR U44863 ( .A(ein[12]), .B(n41854), .Z(ereg_next[13]) );
  AND U44864 ( .A(mul_pow), .B(n41855), .Z(n41854) );
  XOR U44865 ( .A(ein[13]), .B(ein[12]), .Z(n41855) );
  XOR U44866 ( .A(ein[138]), .B(n41856), .Z(ereg_next[139]) );
  AND U44867 ( .A(mul_pow), .B(n41857), .Z(n41856) );
  XOR U44868 ( .A(ein[139]), .B(ein[138]), .Z(n41857) );
  XOR U44869 ( .A(ein[137]), .B(n41858), .Z(ereg_next[138]) );
  AND U44870 ( .A(mul_pow), .B(n41859), .Z(n41858) );
  XOR U44871 ( .A(ein[138]), .B(ein[137]), .Z(n41859) );
  XOR U44872 ( .A(ein[136]), .B(n41860), .Z(ereg_next[137]) );
  AND U44873 ( .A(mul_pow), .B(n41861), .Z(n41860) );
  XOR U44874 ( .A(ein[137]), .B(ein[136]), .Z(n41861) );
  XOR U44875 ( .A(ein[135]), .B(n41862), .Z(ereg_next[136]) );
  AND U44876 ( .A(mul_pow), .B(n41863), .Z(n41862) );
  XOR U44877 ( .A(ein[136]), .B(ein[135]), .Z(n41863) );
  XOR U44878 ( .A(ein[134]), .B(n41864), .Z(ereg_next[135]) );
  AND U44879 ( .A(mul_pow), .B(n41865), .Z(n41864) );
  XOR U44880 ( .A(ein[135]), .B(ein[134]), .Z(n41865) );
  XOR U44881 ( .A(ein[133]), .B(n41866), .Z(ereg_next[134]) );
  AND U44882 ( .A(mul_pow), .B(n41867), .Z(n41866) );
  XOR U44883 ( .A(ein[134]), .B(ein[133]), .Z(n41867) );
  XOR U44884 ( .A(ein[132]), .B(n41868), .Z(ereg_next[133]) );
  AND U44885 ( .A(mul_pow), .B(n41869), .Z(n41868) );
  XOR U44886 ( .A(ein[133]), .B(ein[132]), .Z(n41869) );
  XOR U44887 ( .A(ein[131]), .B(n41870), .Z(ereg_next[132]) );
  AND U44888 ( .A(mul_pow), .B(n41871), .Z(n41870) );
  XOR U44889 ( .A(ein[132]), .B(ein[131]), .Z(n41871) );
  XOR U44890 ( .A(ein[130]), .B(n41872), .Z(ereg_next[131]) );
  AND U44891 ( .A(mul_pow), .B(n41873), .Z(n41872) );
  XOR U44892 ( .A(ein[131]), .B(ein[130]), .Z(n41873) );
  XOR U44893 ( .A(ein[129]), .B(n41874), .Z(ereg_next[130]) );
  AND U44894 ( .A(mul_pow), .B(n41875), .Z(n41874) );
  XOR U44895 ( .A(ein[130]), .B(ein[129]), .Z(n41875) );
  XOR U44896 ( .A(ein[11]), .B(n41876), .Z(ereg_next[12]) );
  AND U44897 ( .A(mul_pow), .B(n41877), .Z(n41876) );
  XOR U44898 ( .A(ein[12]), .B(ein[11]), .Z(n41877) );
  XOR U44899 ( .A(ein[128]), .B(n41878), .Z(ereg_next[129]) );
  AND U44900 ( .A(mul_pow), .B(n41879), .Z(n41878) );
  XOR U44901 ( .A(ein[129]), .B(ein[128]), .Z(n41879) );
  XOR U44902 ( .A(ein[127]), .B(n41880), .Z(ereg_next[128]) );
  AND U44903 ( .A(mul_pow), .B(n41881), .Z(n41880) );
  XOR U44904 ( .A(ein[128]), .B(ein[127]), .Z(n41881) );
  XOR U44905 ( .A(ein[126]), .B(n41882), .Z(ereg_next[127]) );
  AND U44906 ( .A(mul_pow), .B(n41883), .Z(n41882) );
  XOR U44907 ( .A(ein[127]), .B(ein[126]), .Z(n41883) );
  XOR U44908 ( .A(ein[125]), .B(n41884), .Z(ereg_next[126]) );
  AND U44909 ( .A(mul_pow), .B(n41885), .Z(n41884) );
  XOR U44910 ( .A(ein[126]), .B(ein[125]), .Z(n41885) );
  XOR U44911 ( .A(ein[124]), .B(n41886), .Z(ereg_next[125]) );
  AND U44912 ( .A(mul_pow), .B(n41887), .Z(n41886) );
  XOR U44913 ( .A(ein[125]), .B(ein[124]), .Z(n41887) );
  XOR U44914 ( .A(ein[123]), .B(n41888), .Z(ereg_next[124]) );
  AND U44915 ( .A(mul_pow), .B(n41889), .Z(n41888) );
  XOR U44916 ( .A(ein[124]), .B(ein[123]), .Z(n41889) );
  XOR U44917 ( .A(ein[122]), .B(n41890), .Z(ereg_next[123]) );
  AND U44918 ( .A(mul_pow), .B(n41891), .Z(n41890) );
  XOR U44919 ( .A(ein[123]), .B(ein[122]), .Z(n41891) );
  XOR U44920 ( .A(ein[121]), .B(n41892), .Z(ereg_next[122]) );
  AND U44921 ( .A(mul_pow), .B(n41893), .Z(n41892) );
  XOR U44922 ( .A(ein[122]), .B(ein[121]), .Z(n41893) );
  XOR U44923 ( .A(ein[120]), .B(n41894), .Z(ereg_next[121]) );
  AND U44924 ( .A(mul_pow), .B(n41895), .Z(n41894) );
  XOR U44925 ( .A(ein[121]), .B(ein[120]), .Z(n41895) );
  XOR U44926 ( .A(ein[119]), .B(n41896), .Z(ereg_next[120]) );
  AND U44927 ( .A(mul_pow), .B(n41897), .Z(n41896) );
  XOR U44928 ( .A(ein[120]), .B(ein[119]), .Z(n41897) );
  XOR U44929 ( .A(ein[10]), .B(n41898), .Z(ereg_next[11]) );
  AND U44930 ( .A(mul_pow), .B(n41899), .Z(n41898) );
  XOR U44931 ( .A(ein[11]), .B(ein[10]), .Z(n41899) );
  XOR U44932 ( .A(ein[118]), .B(n41900), .Z(ereg_next[119]) );
  AND U44933 ( .A(mul_pow), .B(n41901), .Z(n41900) );
  XOR U44934 ( .A(ein[119]), .B(ein[118]), .Z(n41901) );
  XOR U44935 ( .A(ein[117]), .B(n41902), .Z(ereg_next[118]) );
  AND U44936 ( .A(mul_pow), .B(n41903), .Z(n41902) );
  XOR U44937 ( .A(ein[118]), .B(ein[117]), .Z(n41903) );
  XOR U44938 ( .A(ein[116]), .B(n41904), .Z(ereg_next[117]) );
  AND U44939 ( .A(mul_pow), .B(n41905), .Z(n41904) );
  XOR U44940 ( .A(ein[117]), .B(ein[116]), .Z(n41905) );
  XOR U44941 ( .A(ein[115]), .B(n41906), .Z(ereg_next[116]) );
  AND U44942 ( .A(mul_pow), .B(n41907), .Z(n41906) );
  XOR U44943 ( .A(ein[116]), .B(ein[115]), .Z(n41907) );
  XOR U44944 ( .A(ein[114]), .B(n41908), .Z(ereg_next[115]) );
  AND U44945 ( .A(mul_pow), .B(n41909), .Z(n41908) );
  XOR U44946 ( .A(ein[115]), .B(ein[114]), .Z(n41909) );
  XOR U44947 ( .A(ein[113]), .B(n41910), .Z(ereg_next[114]) );
  AND U44948 ( .A(mul_pow), .B(n41911), .Z(n41910) );
  XOR U44949 ( .A(ein[114]), .B(ein[113]), .Z(n41911) );
  XOR U44950 ( .A(ein[112]), .B(n41912), .Z(ereg_next[113]) );
  AND U44951 ( .A(mul_pow), .B(n41913), .Z(n41912) );
  XOR U44952 ( .A(ein[113]), .B(ein[112]), .Z(n41913) );
  XOR U44953 ( .A(ein[111]), .B(n41914), .Z(ereg_next[112]) );
  AND U44954 ( .A(mul_pow), .B(n41915), .Z(n41914) );
  XOR U44955 ( .A(ein[112]), .B(ein[111]), .Z(n41915) );
  XOR U44956 ( .A(ein[110]), .B(n41916), .Z(ereg_next[111]) );
  AND U44957 ( .A(mul_pow), .B(n41917), .Z(n41916) );
  XOR U44958 ( .A(ein[111]), .B(ein[110]), .Z(n41917) );
  XOR U44959 ( .A(ein[109]), .B(n41918), .Z(ereg_next[110]) );
  AND U44960 ( .A(mul_pow), .B(n41919), .Z(n41918) );
  XOR U44961 ( .A(ein[110]), .B(ein[109]), .Z(n41919) );
  XOR U44962 ( .A(ein[9]), .B(n41920), .Z(ereg_next[10]) );
  AND U44963 ( .A(mul_pow), .B(n41921), .Z(n41920) );
  XOR U44964 ( .A(ein[9]), .B(ein[10]), .Z(n41921) );
  XOR U44965 ( .A(ein[108]), .B(n41922), .Z(ereg_next[109]) );
  AND U44966 ( .A(mul_pow), .B(n41923), .Z(n41922) );
  XOR U44967 ( .A(ein[109]), .B(ein[108]), .Z(n41923) );
  XOR U44968 ( .A(ein[107]), .B(n41924), .Z(ereg_next[108]) );
  AND U44969 ( .A(mul_pow), .B(n41925), .Z(n41924) );
  XOR U44970 ( .A(ein[108]), .B(ein[107]), .Z(n41925) );
  XOR U44971 ( .A(ein[106]), .B(n41926), .Z(ereg_next[107]) );
  AND U44972 ( .A(mul_pow), .B(n41927), .Z(n41926) );
  XOR U44973 ( .A(ein[107]), .B(ein[106]), .Z(n41927) );
  XOR U44974 ( .A(ein[105]), .B(n41928), .Z(ereg_next[106]) );
  AND U44975 ( .A(mul_pow), .B(n41929), .Z(n41928) );
  XOR U44976 ( .A(ein[106]), .B(ein[105]), .Z(n41929) );
  XOR U44977 ( .A(ein[104]), .B(n41930), .Z(ereg_next[105]) );
  AND U44978 ( .A(mul_pow), .B(n41931), .Z(n41930) );
  XOR U44979 ( .A(ein[105]), .B(ein[104]), .Z(n41931) );
  XOR U44980 ( .A(ein[103]), .B(n41932), .Z(ereg_next[104]) );
  AND U44981 ( .A(mul_pow), .B(n41933), .Z(n41932) );
  XOR U44982 ( .A(ein[104]), .B(ein[103]), .Z(n41933) );
  XOR U44983 ( .A(ein[102]), .B(n41934), .Z(ereg_next[103]) );
  AND U44984 ( .A(mul_pow), .B(n41935), .Z(n41934) );
  XOR U44985 ( .A(ein[103]), .B(ein[102]), .Z(n41935) );
  XOR U44986 ( .A(ein[101]), .B(n41936), .Z(ereg_next[102]) );
  AND U44987 ( .A(mul_pow), .B(n41937), .Z(n41936) );
  XOR U44988 ( .A(ein[102]), .B(ein[101]), .Z(n41937) );
  XOR U44989 ( .A(ein[1022]), .B(n41938), .Z(ereg_next[1023]) );
  AND U44990 ( .A(mul_pow), .B(n41939), .Z(n41938) );
  XOR U44991 ( .A(ein[1023]), .B(ein[1022]), .Z(n41939) );
  XOR U44992 ( .A(ein[1021]), .B(n41940), .Z(ereg_next[1022]) );
  AND U44993 ( .A(mul_pow), .B(n41941), .Z(n41940) );
  XOR U44994 ( .A(ein[1022]), .B(ein[1021]), .Z(n41941) );
  XOR U44995 ( .A(ein[1020]), .B(n41942), .Z(ereg_next[1021]) );
  AND U44996 ( .A(mul_pow), .B(n41943), .Z(n41942) );
  XOR U44997 ( .A(ein[1021]), .B(ein[1020]), .Z(n41943) );
  XOR U44998 ( .A(ein[1019]), .B(n41944), .Z(ereg_next[1020]) );
  AND U44999 ( .A(mul_pow), .B(n41945), .Z(n41944) );
  XOR U45000 ( .A(ein[1020]), .B(ein[1019]), .Z(n41945) );
  XOR U45001 ( .A(ein[100]), .B(n41946), .Z(ereg_next[101]) );
  AND U45002 ( .A(mul_pow), .B(n41947), .Z(n41946) );
  XOR U45003 ( .A(ein[101]), .B(ein[100]), .Z(n41947) );
  XOR U45004 ( .A(ein[1018]), .B(n41948), .Z(ereg_next[1019]) );
  AND U45005 ( .A(mul_pow), .B(n41949), .Z(n41948) );
  XOR U45006 ( .A(ein[1019]), .B(ein[1018]), .Z(n41949) );
  XOR U45007 ( .A(ein[1017]), .B(n41950), .Z(ereg_next[1018]) );
  AND U45008 ( .A(mul_pow), .B(n41951), .Z(n41950) );
  XOR U45009 ( .A(ein[1018]), .B(ein[1017]), .Z(n41951) );
  XOR U45010 ( .A(ein[1016]), .B(n41952), .Z(ereg_next[1017]) );
  AND U45011 ( .A(mul_pow), .B(n41953), .Z(n41952) );
  XOR U45012 ( .A(ein[1017]), .B(ein[1016]), .Z(n41953) );
  XOR U45013 ( .A(ein[1015]), .B(n41954), .Z(ereg_next[1016]) );
  AND U45014 ( .A(mul_pow), .B(n41955), .Z(n41954) );
  XOR U45015 ( .A(ein[1016]), .B(ein[1015]), .Z(n41955) );
  XOR U45016 ( .A(ein[1014]), .B(n41956), .Z(ereg_next[1015]) );
  AND U45017 ( .A(mul_pow), .B(n41957), .Z(n41956) );
  XOR U45018 ( .A(ein[1015]), .B(ein[1014]), .Z(n41957) );
  XOR U45019 ( .A(ein[1013]), .B(n41958), .Z(ereg_next[1014]) );
  AND U45020 ( .A(mul_pow), .B(n41959), .Z(n41958) );
  XOR U45021 ( .A(ein[1014]), .B(ein[1013]), .Z(n41959) );
  XOR U45022 ( .A(ein[1012]), .B(n41960), .Z(ereg_next[1013]) );
  AND U45023 ( .A(mul_pow), .B(n41961), .Z(n41960) );
  XOR U45024 ( .A(ein[1013]), .B(ein[1012]), .Z(n41961) );
  XOR U45025 ( .A(ein[1011]), .B(n41962), .Z(ereg_next[1012]) );
  AND U45026 ( .A(mul_pow), .B(n41963), .Z(n41962) );
  XOR U45027 ( .A(ein[1012]), .B(ein[1011]), .Z(n41963) );
  XOR U45028 ( .A(ein[1010]), .B(n41964), .Z(ereg_next[1011]) );
  AND U45029 ( .A(mul_pow), .B(n41965), .Z(n41964) );
  XOR U45030 ( .A(ein[1011]), .B(ein[1010]), .Z(n41965) );
  XOR U45031 ( .A(ein[1009]), .B(n41966), .Z(ereg_next[1010]) );
  AND U45032 ( .A(mul_pow), .B(n41967), .Z(n41966) );
  XOR U45033 ( .A(ein[1010]), .B(ein[1009]), .Z(n41967) );
  XOR U45034 ( .A(ein[99]), .B(n41968), .Z(ereg_next[100]) );
  AND U45035 ( .A(mul_pow), .B(n41969), .Z(n41968) );
  XOR U45036 ( .A(ein[99]), .B(ein[100]), .Z(n41969) );
  XOR U45037 ( .A(ein[1008]), .B(n41970), .Z(ereg_next[1009]) );
  AND U45038 ( .A(mul_pow), .B(n41971), .Z(n41970) );
  XOR U45039 ( .A(ein[1009]), .B(ein[1008]), .Z(n41971) );
  XOR U45040 ( .A(ein[1007]), .B(n41972), .Z(ereg_next[1008]) );
  AND U45041 ( .A(mul_pow), .B(n41973), .Z(n41972) );
  XOR U45042 ( .A(ein[1008]), .B(ein[1007]), .Z(n41973) );
  XOR U45043 ( .A(ein[1006]), .B(n41974), .Z(ereg_next[1007]) );
  AND U45044 ( .A(mul_pow), .B(n41975), .Z(n41974) );
  XOR U45045 ( .A(ein[1007]), .B(ein[1006]), .Z(n41975) );
  XOR U45046 ( .A(ein[1005]), .B(n41976), .Z(ereg_next[1006]) );
  AND U45047 ( .A(mul_pow), .B(n41977), .Z(n41976) );
  XOR U45048 ( .A(ein[1006]), .B(ein[1005]), .Z(n41977) );
  XOR U45049 ( .A(ein[1004]), .B(n41978), .Z(ereg_next[1005]) );
  AND U45050 ( .A(mul_pow), .B(n41979), .Z(n41978) );
  XOR U45051 ( .A(ein[1005]), .B(ein[1004]), .Z(n41979) );
  XOR U45052 ( .A(ein[1003]), .B(n41980), .Z(ereg_next[1004]) );
  AND U45053 ( .A(mul_pow), .B(n41981), .Z(n41980) );
  XOR U45054 ( .A(ein[1004]), .B(ein[1003]), .Z(n41981) );
  XOR U45055 ( .A(ein[1002]), .B(n41982), .Z(ereg_next[1003]) );
  AND U45056 ( .A(mul_pow), .B(n41983), .Z(n41982) );
  XOR U45057 ( .A(ein[1003]), .B(ein[1002]), .Z(n41983) );
  XOR U45058 ( .A(ein[1001]), .B(n41984), .Z(ereg_next[1002]) );
  AND U45059 ( .A(mul_pow), .B(n41985), .Z(n41984) );
  XOR U45060 ( .A(ein[1002]), .B(ein[1001]), .Z(n41985) );
  XOR U45061 ( .A(ein[1000]), .B(n41986), .Z(ereg_next[1001]) );
  AND U45062 ( .A(mul_pow), .B(n41987), .Z(n41986) );
  XOR U45063 ( .A(ein[1001]), .B(ein[1000]), .Z(n41987) );
  XOR U45064 ( .A(ein[999]), .B(n41988), .Z(ereg_next[1000]) );
  AND U45065 ( .A(mul_pow), .B(n41989), .Z(n41988) );
  XOR U45066 ( .A(ein[999]), .B(ein[1000]), .Z(n41989) );
  AND U45067 ( .A(ein[0]), .B(mul_pow), .Z(ereg_next[0]) );
endmodule

