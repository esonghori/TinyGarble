module MixColumns(
x,
z);

	input [127:0] x;
	output [127:0] z;
	wire w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687;

	assign {w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127} = x;

	assign z = {w164, w165, w166, w167, w168, w169, w170, w171, w196, w197, w198, w199, w200, w201, w202, w203, w228, w229, w230, w231, w232, w233, w234, w235, w260, w261, w262, w263, w264, w265, w266, w267, w304, w305, w306, w307, w308, w309, w310, w311, w336, w337, w338, w339, w340, w341, w342, w343, w368, w369, w370, w371, w372, w373, w374, w375, w400, w401, w402, w403, w404, w405, w406, w407, w444, w445, w446, w447, w448, w449, w450, w451, w476, w477, w478, w479, w480, w481, w482, w483, w508, w509, w510, w511, w512, w513, w514, w515, w540, w541, w542, w543, w544, w545, w546, w547, w584, w585, w586, w587, w588, w589, w590, w591, w616, w617, w618, w619, w620, w621, w622, w623, w648, w649, w650, w651, w652, w653, w654, w655, w680, w681, w682, w683, w684, w685, w686, w687};

	XOR U0 ( .A(w7), .B(w2), .Z(w128) );
	XOR U1 ( .A(w7), .B(w3), .Z(w129) );
	XOR U2 ( .A(w7), .B(w0), .Z(w130) );
	XOR U3 ( .A(w15), .B(w10), .Z(w131) );
	XOR U4 ( .A(w15), .B(w11), .Z(w132) );
	XOR U5 ( .A(w15), .B(w8), .Z(w133) );
	XOR U6 ( .A(w23), .B(w18), .Z(w134) );
	XOR U7 ( .A(w23), .B(w19), .Z(w135) );
	XOR U8 ( .A(w23), .B(w16), .Z(w136) );
	XOR U9 ( .A(w31), .B(w26), .Z(w137) );
	XOR U10 ( .A(w31), .B(w27), .Z(w138) );
	XOR U11 ( .A(w31), .B(w24), .Z(w139) );
	XOR U12 ( .A(w7), .B(w15), .Z(w140) );
	XOR U13 ( .A(w130), .B(w133), .Z(w141) );
	XOR U14 ( .A(w1), .B(w9), .Z(w142) );
	XOR U15 ( .A(w128), .B(w131), .Z(w143) );
	XOR U16 ( .A(w129), .B(w132), .Z(w144) );
	XOR U17 ( .A(w4), .B(w12), .Z(w145) );
	XOR U18 ( .A(w5), .B(w13), .Z(w146) );
	XOR U19 ( .A(w6), .B(w14), .Z(w147) );
	XOR U20 ( .A(w140), .B(w8), .Z(w148) );
	XOR U21 ( .A(w141), .B(w9), .Z(w149) );
	XOR U22 ( .A(w142), .B(w10), .Z(w150) );
	XOR U23 ( .A(w143), .B(w11), .Z(w151) );
	XOR U24 ( .A(w144), .B(w12), .Z(w152) );
	XOR U25 ( .A(w145), .B(w13), .Z(w153) );
	XOR U26 ( .A(w146), .B(w14), .Z(w154) );
	XOR U27 ( .A(w147), .B(w15), .Z(w155) );
	XOR U28 ( .A(w148), .B(w16), .Z(w156) );
	XOR U29 ( .A(w149), .B(w17), .Z(w157) );
	XOR U30 ( .A(w150), .B(w18), .Z(w158) );
	XOR U31 ( .A(w151), .B(w19), .Z(w159) );
	XOR U32 ( .A(w152), .B(w20), .Z(w160) );
	XOR U33 ( .A(w153), .B(w21), .Z(w161) );
	XOR U34 ( .A(w154), .B(w22), .Z(w162) );
	XOR U35 ( .A(w155), .B(w23), .Z(w163) );
	XOR U36 ( .A(w156), .B(w24), .Z(w164) );
	XOR U37 ( .A(w157), .B(w25), .Z(w165) );
	XOR U38 ( .A(w158), .B(w26), .Z(w166) );
	XOR U39 ( .A(w159), .B(w27), .Z(w167) );
	XOR U40 ( .A(w160), .B(w28), .Z(w168) );
	XOR U41 ( .A(w161), .B(w29), .Z(w169) );
	XOR U42 ( .A(w162), .B(w30), .Z(w170) );
	XOR U43 ( .A(w163), .B(w31), .Z(w171) );
	XOR U44 ( .A(w15), .B(w23), .Z(w172) );
	XOR U45 ( .A(w133), .B(w136), .Z(w173) );
	XOR U46 ( .A(w9), .B(w17), .Z(w174) );
	XOR U47 ( .A(w131), .B(w134), .Z(w175) );
	XOR U48 ( .A(w132), .B(w135), .Z(w176) );
	XOR U49 ( .A(w12), .B(w20), .Z(w177) );
	XOR U50 ( .A(w13), .B(w21), .Z(w178) );
	XOR U51 ( .A(w14), .B(w22), .Z(w179) );
	XOR U52 ( .A(w172), .B(w16), .Z(w180) );
	XOR U53 ( .A(w173), .B(w17), .Z(w181) );
	XOR U54 ( .A(w174), .B(w18), .Z(w182) );
	XOR U55 ( .A(w175), .B(w19), .Z(w183) );
	XOR U56 ( .A(w176), .B(w20), .Z(w184) );
	XOR U57 ( .A(w177), .B(w21), .Z(w185) );
	XOR U58 ( .A(w178), .B(w22), .Z(w186) );
	XOR U59 ( .A(w179), .B(w23), .Z(w187) );
	XOR U60 ( .A(w180), .B(w24), .Z(w188) );
	XOR U61 ( .A(w181), .B(w25), .Z(w189) );
	XOR U62 ( .A(w182), .B(w26), .Z(w190) );
	XOR U63 ( .A(w183), .B(w27), .Z(w191) );
	XOR U64 ( .A(w184), .B(w28), .Z(w192) );
	XOR U65 ( .A(w185), .B(w29), .Z(w193) );
	XOR U66 ( .A(w186), .B(w30), .Z(w194) );
	XOR U67 ( .A(w187), .B(w31), .Z(w195) );
	XOR U68 ( .A(w188), .B(w0), .Z(w196) );
	XOR U69 ( .A(w189), .B(w1), .Z(w197) );
	XOR U70 ( .A(w190), .B(w2), .Z(w198) );
	XOR U71 ( .A(w191), .B(w3), .Z(w199) );
	XOR U72 ( .A(w192), .B(w4), .Z(w200) );
	XOR U73 ( .A(w193), .B(w5), .Z(w201) );
	XOR U74 ( .A(w194), .B(w6), .Z(w202) );
	XOR U75 ( .A(w195), .B(w7), .Z(w203) );
	XOR U76 ( .A(w23), .B(w31), .Z(w204) );
	XOR U77 ( .A(w136), .B(w139), .Z(w205) );
	XOR U78 ( .A(w17), .B(w25), .Z(w206) );
	XOR U79 ( .A(w134), .B(w137), .Z(w207) );
	XOR U80 ( .A(w135), .B(w138), .Z(w208) );
	XOR U81 ( .A(w20), .B(w28), .Z(w209) );
	XOR U82 ( .A(w21), .B(w29), .Z(w210) );
	XOR U83 ( .A(w22), .B(w30), .Z(w211) );
	XOR U84 ( .A(w204), .B(w24), .Z(w212) );
	XOR U85 ( .A(w205), .B(w25), .Z(w213) );
	XOR U86 ( .A(w206), .B(w26), .Z(w214) );
	XOR U87 ( .A(w207), .B(w27), .Z(w215) );
	XOR U88 ( .A(w208), .B(w28), .Z(w216) );
	XOR U89 ( .A(w209), .B(w29), .Z(w217) );
	XOR U90 ( .A(w210), .B(w30), .Z(w218) );
	XOR U91 ( .A(w211), .B(w31), .Z(w219) );
	XOR U92 ( .A(w212), .B(w0), .Z(w220) );
	XOR U93 ( .A(w213), .B(w1), .Z(w221) );
	XOR U94 ( .A(w214), .B(w2), .Z(w222) );
	XOR U95 ( .A(w215), .B(w3), .Z(w223) );
	XOR U96 ( .A(w216), .B(w4), .Z(w224) );
	XOR U97 ( .A(w217), .B(w5), .Z(w225) );
	XOR U98 ( .A(w218), .B(w6), .Z(w226) );
	XOR U99 ( .A(w219), .B(w7), .Z(w227) );
	XOR U100 ( .A(w220), .B(w8), .Z(w228) );
	XOR U101 ( .A(w221), .B(w9), .Z(w229) );
	XOR U102 ( .A(w222), .B(w10), .Z(w230) );
	XOR U103 ( .A(w223), .B(w11), .Z(w231) );
	XOR U104 ( .A(w224), .B(w12), .Z(w232) );
	XOR U105 ( .A(w225), .B(w13), .Z(w233) );
	XOR U106 ( .A(w226), .B(w14), .Z(w234) );
	XOR U107 ( .A(w227), .B(w15), .Z(w235) );
	XOR U108 ( .A(w31), .B(w7), .Z(w236) );
	XOR U109 ( .A(w139), .B(w130), .Z(w237) );
	XOR U110 ( .A(w25), .B(w1), .Z(w238) );
	XOR U111 ( .A(w137), .B(w128), .Z(w239) );
	XOR U112 ( .A(w138), .B(w129), .Z(w240) );
	XOR U113 ( .A(w28), .B(w4), .Z(w241) );
	XOR U114 ( .A(w29), .B(w5), .Z(w242) );
	XOR U115 ( .A(w30), .B(w6), .Z(w243) );
	XOR U116 ( .A(w236), .B(w0), .Z(w244) );
	XOR U117 ( .A(w237), .B(w1), .Z(w245) );
	XOR U118 ( .A(w238), .B(w2), .Z(w246) );
	XOR U119 ( .A(w239), .B(w3), .Z(w247) );
	XOR U120 ( .A(w240), .B(w4), .Z(w248) );
	XOR U121 ( .A(w241), .B(w5), .Z(w249) );
	XOR U122 ( .A(w242), .B(w6), .Z(w250) );
	XOR U123 ( .A(w243), .B(w7), .Z(w251) );
	XOR U124 ( .A(w244), .B(w8), .Z(w252) );
	XOR U125 ( .A(w245), .B(w9), .Z(w253) );
	XOR U126 ( .A(w246), .B(w10), .Z(w254) );
	XOR U127 ( .A(w247), .B(w11), .Z(w255) );
	XOR U128 ( .A(w248), .B(w12), .Z(w256) );
	XOR U129 ( .A(w249), .B(w13), .Z(w257) );
	XOR U130 ( .A(w250), .B(w14), .Z(w258) );
	XOR U131 ( .A(w251), .B(w15), .Z(w259) );
	XOR U132 ( .A(w252), .B(w16), .Z(w260) );
	XOR U133 ( .A(w253), .B(w17), .Z(w261) );
	XOR U134 ( .A(w254), .B(w18), .Z(w262) );
	XOR U135 ( .A(w255), .B(w19), .Z(w263) );
	XOR U136 ( .A(w256), .B(w20), .Z(w264) );
	XOR U137 ( .A(w257), .B(w21), .Z(w265) );
	XOR U138 ( .A(w258), .B(w22), .Z(w266) );
	XOR U139 ( .A(w259), .B(w23), .Z(w267) );
	XOR U140 ( .A(w39), .B(w34), .Z(w268) );
	XOR U141 ( .A(w39), .B(w35), .Z(w269) );
	XOR U142 ( .A(w39), .B(w32), .Z(w270) );
	XOR U143 ( .A(w47), .B(w42), .Z(w271) );
	XOR U144 ( .A(w47), .B(w43), .Z(w272) );
	XOR U145 ( .A(w47), .B(w40), .Z(w273) );
	XOR U146 ( .A(w55), .B(w50), .Z(w274) );
	XOR U147 ( .A(w55), .B(w51), .Z(w275) );
	XOR U148 ( .A(w55), .B(w48), .Z(w276) );
	XOR U149 ( .A(w63), .B(w58), .Z(w277) );
	XOR U150 ( .A(w63), .B(w59), .Z(w278) );
	XOR U151 ( .A(w63), .B(w56), .Z(w279) );
	XOR U152 ( .A(w39), .B(w47), .Z(w280) );
	XOR U153 ( .A(w270), .B(w273), .Z(w281) );
	XOR U154 ( .A(w33), .B(w41), .Z(w282) );
	XOR U155 ( .A(w268), .B(w271), .Z(w283) );
	XOR U156 ( .A(w269), .B(w272), .Z(w284) );
	XOR U157 ( .A(w36), .B(w44), .Z(w285) );
	XOR U158 ( .A(w37), .B(w45), .Z(w286) );
	XOR U159 ( .A(w38), .B(w46), .Z(w287) );
	XOR U160 ( .A(w280), .B(w40), .Z(w288) );
	XOR U161 ( .A(w281), .B(w41), .Z(w289) );
	XOR U162 ( .A(w282), .B(w42), .Z(w290) );
	XOR U163 ( .A(w283), .B(w43), .Z(w291) );
	XOR U164 ( .A(w284), .B(w44), .Z(w292) );
	XOR U165 ( .A(w285), .B(w45), .Z(w293) );
	XOR U166 ( .A(w286), .B(w46), .Z(w294) );
	XOR U167 ( .A(w287), .B(w47), .Z(w295) );
	XOR U168 ( .A(w288), .B(w48), .Z(w296) );
	XOR U169 ( .A(w289), .B(w49), .Z(w297) );
	XOR U170 ( .A(w290), .B(w50), .Z(w298) );
	XOR U171 ( .A(w291), .B(w51), .Z(w299) );
	XOR U172 ( .A(w292), .B(w52), .Z(w300) );
	XOR U173 ( .A(w293), .B(w53), .Z(w301) );
	XOR U174 ( .A(w294), .B(w54), .Z(w302) );
	XOR U175 ( .A(w295), .B(w55), .Z(w303) );
	XOR U176 ( .A(w296), .B(w56), .Z(w304) );
	XOR U177 ( .A(w297), .B(w57), .Z(w305) );
	XOR U178 ( .A(w298), .B(w58), .Z(w306) );
	XOR U179 ( .A(w299), .B(w59), .Z(w307) );
	XOR U180 ( .A(w300), .B(w60), .Z(w308) );
	XOR U181 ( .A(w301), .B(w61), .Z(w309) );
	XOR U182 ( .A(w302), .B(w62), .Z(w310) );
	XOR U183 ( .A(w303), .B(w63), .Z(w311) );
	XOR U184 ( .A(w47), .B(w55), .Z(w312) );
	XOR U185 ( .A(w273), .B(w276), .Z(w313) );
	XOR U186 ( .A(w41), .B(w49), .Z(w314) );
	XOR U187 ( .A(w271), .B(w274), .Z(w315) );
	XOR U188 ( .A(w272), .B(w275), .Z(w316) );
	XOR U189 ( .A(w44), .B(w52), .Z(w317) );
	XOR U190 ( .A(w45), .B(w53), .Z(w318) );
	XOR U191 ( .A(w46), .B(w54), .Z(w319) );
	XOR U192 ( .A(w312), .B(w48), .Z(w320) );
	XOR U193 ( .A(w313), .B(w49), .Z(w321) );
	XOR U194 ( .A(w314), .B(w50), .Z(w322) );
	XOR U195 ( .A(w315), .B(w51), .Z(w323) );
	XOR U196 ( .A(w316), .B(w52), .Z(w324) );
	XOR U197 ( .A(w317), .B(w53), .Z(w325) );
	XOR U198 ( .A(w318), .B(w54), .Z(w326) );
	XOR U199 ( .A(w319), .B(w55), .Z(w327) );
	XOR U200 ( .A(w320), .B(w56), .Z(w328) );
	XOR U201 ( .A(w321), .B(w57), .Z(w329) );
	XOR U202 ( .A(w322), .B(w58), .Z(w330) );
	XOR U203 ( .A(w323), .B(w59), .Z(w331) );
	XOR U204 ( .A(w324), .B(w60), .Z(w332) );
	XOR U205 ( .A(w325), .B(w61), .Z(w333) );
	XOR U206 ( .A(w326), .B(w62), .Z(w334) );
	XOR U207 ( .A(w327), .B(w63), .Z(w335) );
	XOR U208 ( .A(w328), .B(w32), .Z(w336) );
	XOR U209 ( .A(w329), .B(w33), .Z(w337) );
	XOR U210 ( .A(w330), .B(w34), .Z(w338) );
	XOR U211 ( .A(w331), .B(w35), .Z(w339) );
	XOR U212 ( .A(w332), .B(w36), .Z(w340) );
	XOR U213 ( .A(w333), .B(w37), .Z(w341) );
	XOR U214 ( .A(w334), .B(w38), .Z(w342) );
	XOR U215 ( .A(w335), .B(w39), .Z(w343) );
	XOR U216 ( .A(w55), .B(w63), .Z(w344) );
	XOR U217 ( .A(w276), .B(w279), .Z(w345) );
	XOR U218 ( .A(w49), .B(w57), .Z(w346) );
	XOR U219 ( .A(w274), .B(w277), .Z(w347) );
	XOR U220 ( .A(w275), .B(w278), .Z(w348) );
	XOR U221 ( .A(w52), .B(w60), .Z(w349) );
	XOR U222 ( .A(w53), .B(w61), .Z(w350) );
	XOR U223 ( .A(w54), .B(w62), .Z(w351) );
	XOR U224 ( .A(w344), .B(w56), .Z(w352) );
	XOR U225 ( .A(w345), .B(w57), .Z(w353) );
	XOR U226 ( .A(w346), .B(w58), .Z(w354) );
	XOR U227 ( .A(w347), .B(w59), .Z(w355) );
	XOR U228 ( .A(w348), .B(w60), .Z(w356) );
	XOR U229 ( .A(w349), .B(w61), .Z(w357) );
	XOR U230 ( .A(w350), .B(w62), .Z(w358) );
	XOR U231 ( .A(w351), .B(w63), .Z(w359) );
	XOR U232 ( .A(w352), .B(w32), .Z(w360) );
	XOR U233 ( .A(w353), .B(w33), .Z(w361) );
	XOR U234 ( .A(w354), .B(w34), .Z(w362) );
	XOR U235 ( .A(w355), .B(w35), .Z(w363) );
	XOR U236 ( .A(w356), .B(w36), .Z(w364) );
	XOR U237 ( .A(w357), .B(w37), .Z(w365) );
	XOR U238 ( .A(w358), .B(w38), .Z(w366) );
	XOR U239 ( .A(w359), .B(w39), .Z(w367) );
	XOR U240 ( .A(w360), .B(w40), .Z(w368) );
	XOR U241 ( .A(w361), .B(w41), .Z(w369) );
	XOR U242 ( .A(w362), .B(w42), .Z(w370) );
	XOR U243 ( .A(w363), .B(w43), .Z(w371) );
	XOR U244 ( .A(w364), .B(w44), .Z(w372) );
	XOR U245 ( .A(w365), .B(w45), .Z(w373) );
	XOR U246 ( .A(w366), .B(w46), .Z(w374) );
	XOR U247 ( .A(w367), .B(w47), .Z(w375) );
	XOR U248 ( .A(w63), .B(w39), .Z(w376) );
	XOR U249 ( .A(w279), .B(w270), .Z(w377) );
	XOR U250 ( .A(w57), .B(w33), .Z(w378) );
	XOR U251 ( .A(w277), .B(w268), .Z(w379) );
	XOR U252 ( .A(w278), .B(w269), .Z(w380) );
	XOR U253 ( .A(w60), .B(w36), .Z(w381) );
	XOR U254 ( .A(w61), .B(w37), .Z(w382) );
	XOR U255 ( .A(w62), .B(w38), .Z(w383) );
	XOR U256 ( .A(w376), .B(w32), .Z(w384) );
	XOR U257 ( .A(w377), .B(w33), .Z(w385) );
	XOR U258 ( .A(w378), .B(w34), .Z(w386) );
	XOR U259 ( .A(w379), .B(w35), .Z(w387) );
	XOR U260 ( .A(w380), .B(w36), .Z(w388) );
	XOR U261 ( .A(w381), .B(w37), .Z(w389) );
	XOR U262 ( .A(w382), .B(w38), .Z(w390) );
	XOR U263 ( .A(w383), .B(w39), .Z(w391) );
	XOR U264 ( .A(w384), .B(w40), .Z(w392) );
	XOR U265 ( .A(w385), .B(w41), .Z(w393) );
	XOR U266 ( .A(w386), .B(w42), .Z(w394) );
	XOR U267 ( .A(w387), .B(w43), .Z(w395) );
	XOR U268 ( .A(w388), .B(w44), .Z(w396) );
	XOR U269 ( .A(w389), .B(w45), .Z(w397) );
	XOR U270 ( .A(w390), .B(w46), .Z(w398) );
	XOR U271 ( .A(w391), .B(w47), .Z(w399) );
	XOR U272 ( .A(w392), .B(w48), .Z(w400) );
	XOR U273 ( .A(w393), .B(w49), .Z(w401) );
	XOR U274 ( .A(w394), .B(w50), .Z(w402) );
	XOR U275 ( .A(w395), .B(w51), .Z(w403) );
	XOR U276 ( .A(w396), .B(w52), .Z(w404) );
	XOR U277 ( .A(w397), .B(w53), .Z(w405) );
	XOR U278 ( .A(w398), .B(w54), .Z(w406) );
	XOR U279 ( .A(w399), .B(w55), .Z(w407) );
	XOR U280 ( .A(w71), .B(w66), .Z(w408) );
	XOR U281 ( .A(w71), .B(w67), .Z(w409) );
	XOR U282 ( .A(w71), .B(w64), .Z(w410) );
	XOR U283 ( .A(w79), .B(w74), .Z(w411) );
	XOR U284 ( .A(w79), .B(w75), .Z(w412) );
	XOR U285 ( .A(w79), .B(w72), .Z(w413) );
	XOR U286 ( .A(w87), .B(w82), .Z(w414) );
	XOR U287 ( .A(w87), .B(w83), .Z(w415) );
	XOR U288 ( .A(w87), .B(w80), .Z(w416) );
	XOR U289 ( .A(w95), .B(w90), .Z(w417) );
	XOR U290 ( .A(w95), .B(w91), .Z(w418) );
	XOR U291 ( .A(w95), .B(w88), .Z(w419) );
	XOR U292 ( .A(w71), .B(w79), .Z(w420) );
	XOR U293 ( .A(w410), .B(w413), .Z(w421) );
	XOR U294 ( .A(w65), .B(w73), .Z(w422) );
	XOR U295 ( .A(w408), .B(w411), .Z(w423) );
	XOR U296 ( .A(w409), .B(w412), .Z(w424) );
	XOR U297 ( .A(w68), .B(w76), .Z(w425) );
	XOR U298 ( .A(w69), .B(w77), .Z(w426) );
	XOR U299 ( .A(w70), .B(w78), .Z(w427) );
	XOR U300 ( .A(w420), .B(w72), .Z(w428) );
	XOR U301 ( .A(w421), .B(w73), .Z(w429) );
	XOR U302 ( .A(w422), .B(w74), .Z(w430) );
	XOR U303 ( .A(w423), .B(w75), .Z(w431) );
	XOR U304 ( .A(w424), .B(w76), .Z(w432) );
	XOR U305 ( .A(w425), .B(w77), .Z(w433) );
	XOR U306 ( .A(w426), .B(w78), .Z(w434) );
	XOR U307 ( .A(w427), .B(w79), .Z(w435) );
	XOR U308 ( .A(w428), .B(w80), .Z(w436) );
	XOR U309 ( .A(w429), .B(w81), .Z(w437) );
	XOR U310 ( .A(w430), .B(w82), .Z(w438) );
	XOR U311 ( .A(w431), .B(w83), .Z(w439) );
	XOR U312 ( .A(w432), .B(w84), .Z(w440) );
	XOR U313 ( .A(w433), .B(w85), .Z(w441) );
	XOR U314 ( .A(w434), .B(w86), .Z(w442) );
	XOR U315 ( .A(w435), .B(w87), .Z(w443) );
	XOR U316 ( .A(w436), .B(w88), .Z(w444) );
	XOR U317 ( .A(w437), .B(w89), .Z(w445) );
	XOR U318 ( .A(w438), .B(w90), .Z(w446) );
	XOR U319 ( .A(w439), .B(w91), .Z(w447) );
	XOR U320 ( .A(w440), .B(w92), .Z(w448) );
	XOR U321 ( .A(w441), .B(w93), .Z(w449) );
	XOR U322 ( .A(w442), .B(w94), .Z(w450) );
	XOR U323 ( .A(w443), .B(w95), .Z(w451) );
	XOR U324 ( .A(w79), .B(w87), .Z(w452) );
	XOR U325 ( .A(w413), .B(w416), .Z(w453) );
	XOR U326 ( .A(w73), .B(w81), .Z(w454) );
	XOR U327 ( .A(w411), .B(w414), .Z(w455) );
	XOR U328 ( .A(w412), .B(w415), .Z(w456) );
	XOR U329 ( .A(w76), .B(w84), .Z(w457) );
	XOR U330 ( .A(w77), .B(w85), .Z(w458) );
	XOR U331 ( .A(w78), .B(w86), .Z(w459) );
	XOR U332 ( .A(w452), .B(w80), .Z(w460) );
	XOR U333 ( .A(w453), .B(w81), .Z(w461) );
	XOR U334 ( .A(w454), .B(w82), .Z(w462) );
	XOR U335 ( .A(w455), .B(w83), .Z(w463) );
	XOR U336 ( .A(w456), .B(w84), .Z(w464) );
	XOR U337 ( .A(w457), .B(w85), .Z(w465) );
	XOR U338 ( .A(w458), .B(w86), .Z(w466) );
	XOR U339 ( .A(w459), .B(w87), .Z(w467) );
	XOR U340 ( .A(w460), .B(w88), .Z(w468) );
	XOR U341 ( .A(w461), .B(w89), .Z(w469) );
	XOR U342 ( .A(w462), .B(w90), .Z(w470) );
	XOR U343 ( .A(w463), .B(w91), .Z(w471) );
	XOR U344 ( .A(w464), .B(w92), .Z(w472) );
	XOR U345 ( .A(w465), .B(w93), .Z(w473) );
	XOR U346 ( .A(w466), .B(w94), .Z(w474) );
	XOR U347 ( .A(w467), .B(w95), .Z(w475) );
	XOR U348 ( .A(w468), .B(w64), .Z(w476) );
	XOR U349 ( .A(w469), .B(w65), .Z(w477) );
	XOR U350 ( .A(w470), .B(w66), .Z(w478) );
	XOR U351 ( .A(w471), .B(w67), .Z(w479) );
	XOR U352 ( .A(w472), .B(w68), .Z(w480) );
	XOR U353 ( .A(w473), .B(w69), .Z(w481) );
	XOR U354 ( .A(w474), .B(w70), .Z(w482) );
	XOR U355 ( .A(w475), .B(w71), .Z(w483) );
	XOR U356 ( .A(w87), .B(w95), .Z(w484) );
	XOR U357 ( .A(w416), .B(w419), .Z(w485) );
	XOR U358 ( .A(w81), .B(w89), .Z(w486) );
	XOR U359 ( .A(w414), .B(w417), .Z(w487) );
	XOR U360 ( .A(w415), .B(w418), .Z(w488) );
	XOR U361 ( .A(w84), .B(w92), .Z(w489) );
	XOR U362 ( .A(w85), .B(w93), .Z(w490) );
	XOR U363 ( .A(w86), .B(w94), .Z(w491) );
	XOR U364 ( .A(w484), .B(w88), .Z(w492) );
	XOR U365 ( .A(w485), .B(w89), .Z(w493) );
	XOR U366 ( .A(w486), .B(w90), .Z(w494) );
	XOR U367 ( .A(w487), .B(w91), .Z(w495) );
	XOR U368 ( .A(w488), .B(w92), .Z(w496) );
	XOR U369 ( .A(w489), .B(w93), .Z(w497) );
	XOR U370 ( .A(w490), .B(w94), .Z(w498) );
	XOR U371 ( .A(w491), .B(w95), .Z(w499) );
	XOR U372 ( .A(w492), .B(w64), .Z(w500) );
	XOR U373 ( .A(w493), .B(w65), .Z(w501) );
	XOR U374 ( .A(w494), .B(w66), .Z(w502) );
	XOR U375 ( .A(w495), .B(w67), .Z(w503) );
	XOR U376 ( .A(w496), .B(w68), .Z(w504) );
	XOR U377 ( .A(w497), .B(w69), .Z(w505) );
	XOR U378 ( .A(w498), .B(w70), .Z(w506) );
	XOR U379 ( .A(w499), .B(w71), .Z(w507) );
	XOR U380 ( .A(w500), .B(w72), .Z(w508) );
	XOR U381 ( .A(w501), .B(w73), .Z(w509) );
	XOR U382 ( .A(w502), .B(w74), .Z(w510) );
	XOR U383 ( .A(w503), .B(w75), .Z(w511) );
	XOR U384 ( .A(w504), .B(w76), .Z(w512) );
	XOR U385 ( .A(w505), .B(w77), .Z(w513) );
	XOR U386 ( .A(w506), .B(w78), .Z(w514) );
	XOR U387 ( .A(w507), .B(w79), .Z(w515) );
	XOR U388 ( .A(w95), .B(w71), .Z(w516) );
	XOR U389 ( .A(w419), .B(w410), .Z(w517) );
	XOR U390 ( .A(w89), .B(w65), .Z(w518) );
	XOR U391 ( .A(w417), .B(w408), .Z(w519) );
	XOR U392 ( .A(w418), .B(w409), .Z(w520) );
	XOR U393 ( .A(w92), .B(w68), .Z(w521) );
	XOR U394 ( .A(w93), .B(w69), .Z(w522) );
	XOR U395 ( .A(w94), .B(w70), .Z(w523) );
	XOR U396 ( .A(w516), .B(w64), .Z(w524) );
	XOR U397 ( .A(w517), .B(w65), .Z(w525) );
	XOR U398 ( .A(w518), .B(w66), .Z(w526) );
	XOR U399 ( .A(w519), .B(w67), .Z(w527) );
	XOR U400 ( .A(w520), .B(w68), .Z(w528) );
	XOR U401 ( .A(w521), .B(w69), .Z(w529) );
	XOR U402 ( .A(w522), .B(w70), .Z(w530) );
	XOR U403 ( .A(w523), .B(w71), .Z(w531) );
	XOR U404 ( .A(w524), .B(w72), .Z(w532) );
	XOR U405 ( .A(w525), .B(w73), .Z(w533) );
	XOR U406 ( .A(w526), .B(w74), .Z(w534) );
	XOR U407 ( .A(w527), .B(w75), .Z(w535) );
	XOR U408 ( .A(w528), .B(w76), .Z(w536) );
	XOR U409 ( .A(w529), .B(w77), .Z(w537) );
	XOR U410 ( .A(w530), .B(w78), .Z(w538) );
	XOR U411 ( .A(w531), .B(w79), .Z(w539) );
	XOR U412 ( .A(w532), .B(w80), .Z(w540) );
	XOR U413 ( .A(w533), .B(w81), .Z(w541) );
	XOR U414 ( .A(w534), .B(w82), .Z(w542) );
	XOR U415 ( .A(w535), .B(w83), .Z(w543) );
	XOR U416 ( .A(w536), .B(w84), .Z(w544) );
	XOR U417 ( .A(w537), .B(w85), .Z(w545) );
	XOR U418 ( .A(w538), .B(w86), .Z(w546) );
	XOR U419 ( .A(w539), .B(w87), .Z(w547) );
	XOR U420 ( .A(w103), .B(w98), .Z(w548) );
	XOR U421 ( .A(w103), .B(w99), .Z(w549) );
	XOR U422 ( .A(w103), .B(w96), .Z(w550) );
	XOR U423 ( .A(w111), .B(w106), .Z(w551) );
	XOR U424 ( .A(w111), .B(w107), .Z(w552) );
	XOR U425 ( .A(w111), .B(w104), .Z(w553) );
	XOR U426 ( .A(w119), .B(w114), .Z(w554) );
	XOR U427 ( .A(w119), .B(w115), .Z(w555) );
	XOR U428 ( .A(w119), .B(w112), .Z(w556) );
	XOR U429 ( .A(w127), .B(w122), .Z(w557) );
	XOR U430 ( .A(w127), .B(w123), .Z(w558) );
	XOR U431 ( .A(w127), .B(w120), .Z(w559) );
	XOR U432 ( .A(w103), .B(w111), .Z(w560) );
	XOR U433 ( .A(w550), .B(w553), .Z(w561) );
	XOR U434 ( .A(w97), .B(w105), .Z(w562) );
	XOR U435 ( .A(w548), .B(w551), .Z(w563) );
	XOR U436 ( .A(w549), .B(w552), .Z(w564) );
	XOR U437 ( .A(w100), .B(w108), .Z(w565) );
	XOR U438 ( .A(w101), .B(w109), .Z(w566) );
	XOR U439 ( .A(w102), .B(w110), .Z(w567) );
	XOR U440 ( .A(w560), .B(w104), .Z(w568) );
	XOR U441 ( .A(w561), .B(w105), .Z(w569) );
	XOR U442 ( .A(w562), .B(w106), .Z(w570) );
	XOR U443 ( .A(w563), .B(w107), .Z(w571) );
	XOR U444 ( .A(w564), .B(w108), .Z(w572) );
	XOR U445 ( .A(w565), .B(w109), .Z(w573) );
	XOR U446 ( .A(w566), .B(w110), .Z(w574) );
	XOR U447 ( .A(w567), .B(w111), .Z(w575) );
	XOR U448 ( .A(w568), .B(w112), .Z(w576) );
	XOR U449 ( .A(w569), .B(w113), .Z(w577) );
	XOR U450 ( .A(w570), .B(w114), .Z(w578) );
	XOR U451 ( .A(w571), .B(w115), .Z(w579) );
	XOR U452 ( .A(w572), .B(w116), .Z(w580) );
	XOR U453 ( .A(w573), .B(w117), .Z(w581) );
	XOR U454 ( .A(w574), .B(w118), .Z(w582) );
	XOR U455 ( .A(w575), .B(w119), .Z(w583) );
	XOR U456 ( .A(w576), .B(w120), .Z(w584) );
	XOR U457 ( .A(w577), .B(w121), .Z(w585) );
	XOR U458 ( .A(w578), .B(w122), .Z(w586) );
	XOR U459 ( .A(w579), .B(w123), .Z(w587) );
	XOR U460 ( .A(w580), .B(w124), .Z(w588) );
	XOR U461 ( .A(w581), .B(w125), .Z(w589) );
	XOR U462 ( .A(w582), .B(w126), .Z(w590) );
	XOR U463 ( .A(w583), .B(w127), .Z(w591) );
	XOR U464 ( .A(w111), .B(w119), .Z(w592) );
	XOR U465 ( .A(w553), .B(w556), .Z(w593) );
	XOR U466 ( .A(w105), .B(w113), .Z(w594) );
	XOR U467 ( .A(w551), .B(w554), .Z(w595) );
	XOR U468 ( .A(w552), .B(w555), .Z(w596) );
	XOR U469 ( .A(w108), .B(w116), .Z(w597) );
	XOR U470 ( .A(w109), .B(w117), .Z(w598) );
	XOR U471 ( .A(w110), .B(w118), .Z(w599) );
	XOR U472 ( .A(w592), .B(w112), .Z(w600) );
	XOR U473 ( .A(w593), .B(w113), .Z(w601) );
	XOR U474 ( .A(w594), .B(w114), .Z(w602) );
	XOR U475 ( .A(w595), .B(w115), .Z(w603) );
	XOR U476 ( .A(w596), .B(w116), .Z(w604) );
	XOR U477 ( .A(w597), .B(w117), .Z(w605) );
	XOR U478 ( .A(w598), .B(w118), .Z(w606) );
	XOR U479 ( .A(w599), .B(w119), .Z(w607) );
	XOR U480 ( .A(w600), .B(w120), .Z(w608) );
	XOR U481 ( .A(w601), .B(w121), .Z(w609) );
	XOR U482 ( .A(w602), .B(w122), .Z(w610) );
	XOR U483 ( .A(w603), .B(w123), .Z(w611) );
	XOR U484 ( .A(w604), .B(w124), .Z(w612) );
	XOR U485 ( .A(w605), .B(w125), .Z(w613) );
	XOR U486 ( .A(w606), .B(w126), .Z(w614) );
	XOR U487 ( .A(w607), .B(w127), .Z(w615) );
	XOR U488 ( .A(w608), .B(w96), .Z(w616) );
	XOR U489 ( .A(w609), .B(w97), .Z(w617) );
	XOR U490 ( .A(w610), .B(w98), .Z(w618) );
	XOR U491 ( .A(w611), .B(w99), .Z(w619) );
	XOR U492 ( .A(w612), .B(w100), .Z(w620) );
	XOR U493 ( .A(w613), .B(w101), .Z(w621) );
	XOR U494 ( .A(w614), .B(w102), .Z(w622) );
	XOR U495 ( .A(w615), .B(w103), .Z(w623) );
	XOR U496 ( .A(w119), .B(w127), .Z(w624) );
	XOR U497 ( .A(w556), .B(w559), .Z(w625) );
	XOR U498 ( .A(w113), .B(w121), .Z(w626) );
	XOR U499 ( .A(w554), .B(w557), .Z(w627) );
	XOR U500 ( .A(w555), .B(w558), .Z(w628) );
	XOR U501 ( .A(w116), .B(w124), .Z(w629) );
	XOR U502 ( .A(w117), .B(w125), .Z(w630) );
	XOR U503 ( .A(w118), .B(w126), .Z(w631) );
	XOR U504 ( .A(w624), .B(w120), .Z(w632) );
	XOR U505 ( .A(w625), .B(w121), .Z(w633) );
	XOR U506 ( .A(w626), .B(w122), .Z(w634) );
	XOR U507 ( .A(w627), .B(w123), .Z(w635) );
	XOR U508 ( .A(w628), .B(w124), .Z(w636) );
	XOR U509 ( .A(w629), .B(w125), .Z(w637) );
	XOR U510 ( .A(w630), .B(w126), .Z(w638) );
	XOR U511 ( .A(w631), .B(w127), .Z(w639) );
	XOR U512 ( .A(w632), .B(w96), .Z(w640) );
	XOR U513 ( .A(w633), .B(w97), .Z(w641) );
	XOR U514 ( .A(w634), .B(w98), .Z(w642) );
	XOR U515 ( .A(w635), .B(w99), .Z(w643) );
	XOR U516 ( .A(w636), .B(w100), .Z(w644) );
	XOR U517 ( .A(w637), .B(w101), .Z(w645) );
	XOR U518 ( .A(w638), .B(w102), .Z(w646) );
	XOR U519 ( .A(w639), .B(w103), .Z(w647) );
	XOR U520 ( .A(w640), .B(w104), .Z(w648) );
	XOR U521 ( .A(w641), .B(w105), .Z(w649) );
	XOR U522 ( .A(w642), .B(w106), .Z(w650) );
	XOR U523 ( .A(w643), .B(w107), .Z(w651) );
	XOR U524 ( .A(w644), .B(w108), .Z(w652) );
	XOR U525 ( .A(w645), .B(w109), .Z(w653) );
	XOR U526 ( .A(w646), .B(w110), .Z(w654) );
	XOR U527 ( .A(w647), .B(w111), .Z(w655) );
	XOR U528 ( .A(w127), .B(w103), .Z(w656) );
	XOR U529 ( .A(w559), .B(w550), .Z(w657) );
	XOR U530 ( .A(w121), .B(w97), .Z(w658) );
	XOR U531 ( .A(w557), .B(w548), .Z(w659) );
	XOR U532 ( .A(w558), .B(w549), .Z(w660) );
	XOR U533 ( .A(w124), .B(w100), .Z(w661) );
	XOR U534 ( .A(w125), .B(w101), .Z(w662) );
	XOR U535 ( .A(w126), .B(w102), .Z(w663) );
	XOR U536 ( .A(w656), .B(w96), .Z(w664) );
	XOR U537 ( .A(w657), .B(w97), .Z(w665) );
	XOR U538 ( .A(w658), .B(w98), .Z(w666) );
	XOR U539 ( .A(w659), .B(w99), .Z(w667) );
	XOR U540 ( .A(w660), .B(w100), .Z(w668) );
	XOR U541 ( .A(w661), .B(w101), .Z(w669) );
	XOR U542 ( .A(w662), .B(w102), .Z(w670) );
	XOR U543 ( .A(w663), .B(w103), .Z(w671) );
	XOR U544 ( .A(w664), .B(w104), .Z(w672) );
	XOR U545 ( .A(w665), .B(w105), .Z(w673) );
	XOR U546 ( .A(w666), .B(w106), .Z(w674) );
	XOR U547 ( .A(w667), .B(w107), .Z(w675) );
	XOR U548 ( .A(w668), .B(w108), .Z(w676) );
	XOR U549 ( .A(w669), .B(w109), .Z(w677) );
	XOR U550 ( .A(w670), .B(w110), .Z(w678) );
	XOR U551 ( .A(w671), .B(w111), .Z(w679) );
	XOR U552 ( .A(w672), .B(w112), .Z(w680) );
	XOR U553 ( .A(w673), .B(w113), .Z(w681) );
	XOR U554 ( .A(w674), .B(w114), .Z(w682) );
	XOR U555 ( .A(w675), .B(w115), .Z(w683) );
	XOR U556 ( .A(w676), .B(w116), .Z(w684) );
	XOR U557 ( .A(w677), .B(w117), .Z(w685) );
	XOR U558 ( .A(w678), .B(w118), .Z(w686) );
	XOR U559 ( .A(w679), .B(w119), .Z(w687) );
endmodule

