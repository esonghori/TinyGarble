
module mult_N64_CC16 ( clk, rst, a, b, c );
  input [63:0] a;
  input [3:0] b;
  output [127:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765;
  wire   [127:0] sreg;

  DFF \sreg_reg[123]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(sreg[123]) );
  DFF \sreg_reg[122]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(sreg[122]) );
  DFF \sreg_reg[121]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(sreg[121]) );
  DFF \sreg_reg[120]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(sreg[120]) );
  DFF \sreg_reg[119]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(sreg[119]) );
  DFF \sreg_reg[118]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(sreg[118]) );
  DFF \sreg_reg[117]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(sreg[117]) );
  DFF \sreg_reg[116]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(sreg[116]) );
  DFF \sreg_reg[115]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(sreg[115]) );
  DFF \sreg_reg[114]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(sreg[114]) );
  DFF \sreg_reg[113]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(sreg[113]) );
  DFF \sreg_reg[112]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(sreg[112]) );
  DFF \sreg_reg[111]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(sreg[111]) );
  DFF \sreg_reg[110]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(sreg[110]) );
  DFF \sreg_reg[109]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(sreg[109]) );
  DFF \sreg_reg[108]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(sreg[108]) );
  DFF \sreg_reg[107]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(sreg[107]) );
  DFF \sreg_reg[106]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(sreg[106]) );
  DFF \sreg_reg[105]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(sreg[105]) );
  DFF \sreg_reg[104]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(sreg[104]) );
  DFF \sreg_reg[103]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(sreg[103]) );
  DFF \sreg_reg[102]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(sreg[102]) );
  DFF \sreg_reg[101]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(sreg[101]) );
  DFF \sreg_reg[100]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(sreg[100]) );
  DFF \sreg_reg[99]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(sreg[99]) );
  DFF \sreg_reg[98]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(sreg[98]) );
  DFF \sreg_reg[97]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(sreg[97]) );
  DFF \sreg_reg[96]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(sreg[96]) );
  DFF \sreg_reg[95]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(sreg[95]) );
  DFF \sreg_reg[94]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(sreg[94]) );
  DFF \sreg_reg[93]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(sreg[93]) );
  DFF \sreg_reg[92]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(sreg[92]) );
  DFF \sreg_reg[91]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(sreg[91]) );
  DFF \sreg_reg[90]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(sreg[90]) );
  DFF \sreg_reg[89]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(sreg[89]) );
  DFF \sreg_reg[88]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(sreg[88]) );
  DFF \sreg_reg[87]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(sreg[87]) );
  DFF \sreg_reg[86]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(sreg[86]) );
  DFF \sreg_reg[85]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(sreg[85]) );
  DFF \sreg_reg[84]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(sreg[84]) );
  DFF \sreg_reg[83]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(sreg[83]) );
  DFF \sreg_reg[82]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(sreg[82]) );
  DFF \sreg_reg[81]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(sreg[81]) );
  DFF \sreg_reg[80]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(sreg[80]) );
  DFF \sreg_reg[79]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(sreg[79]) );
  DFF \sreg_reg[78]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(sreg[78]) );
  DFF \sreg_reg[77]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(sreg[77]) );
  DFF \sreg_reg[76]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(sreg[76]) );
  DFF \sreg_reg[75]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(sreg[75]) );
  DFF \sreg_reg[74]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(sreg[74]) );
  DFF \sreg_reg[73]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(sreg[73]) );
  DFF \sreg_reg[72]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(sreg[72]) );
  DFF \sreg_reg[71]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(sreg[71]) );
  DFF \sreg_reg[70]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(sreg[70]) );
  DFF \sreg_reg[69]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(sreg[69]) );
  DFF \sreg_reg[68]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(sreg[68]) );
  DFF \sreg_reg[67]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(sreg[67]) );
  DFF \sreg_reg[66]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(sreg[66]) );
  DFF \sreg_reg[65]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(sreg[65]) );
  DFF \sreg_reg[64]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(sreg[64]) );
  DFF \sreg_reg[63]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(sreg[63]) );
  DFF \sreg_reg[62]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(sreg[62]) );
  DFF \sreg_reg[61]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(sreg[61]) );
  DFF \sreg_reg[60]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(sreg[60]) );
  DFF \sreg_reg[59]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[58]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[57]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[56]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[55]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[54]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[53]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[52]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[51]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[50]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[49]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[48]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[47]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[46]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[45]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[44]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[43]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[42]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[41]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[40]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[39]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[38]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[37]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[36]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[35]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[34]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[33]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[32]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[31]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[7]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[6]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[5]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[4]), .CLK(clk), .RST(rst), .Q(c[0]) );
  AND U7 ( .A(n578), .B(n579), .Z(n602) );
  XOR U8 ( .A(n607), .B(n608), .Z(n1) );
  NANDN U9 ( .A(n609), .B(n1), .Z(n2) );
  NAND U10 ( .A(n607), .B(n608), .Z(n3) );
  AND U11 ( .A(n2), .B(n3), .Z(n632) );
  NAND U12 ( .A(n624), .B(n625), .Z(n4) );
  XOR U13 ( .A(n624), .B(n625), .Z(n5) );
  NANDN U14 ( .A(n623), .B(n5), .Z(n6) );
  NAND U15 ( .A(n4), .B(n6), .Z(n651) );
  XOR U16 ( .A(n1702), .B(n1703), .Z(n7) );
  NANDN U17 ( .A(n1704), .B(n7), .Z(n8) );
  NAND U18 ( .A(n1702), .B(n1703), .Z(n9) );
  AND U19 ( .A(n8), .B(n9), .Z(n1724) );
  XOR U20 ( .A(n1732), .B(n1733), .Z(n10) );
  NANDN U21 ( .A(n1734), .B(n10), .Z(n11) );
  NAND U22 ( .A(n1732), .B(n1733), .Z(n12) );
  AND U23 ( .A(n11), .B(n12), .Z(n1748) );
  NAND U24 ( .A(n584), .B(n585), .Z(n13) );
  XOR U25 ( .A(n584), .B(n585), .Z(n14) );
  NANDN U26 ( .A(n583), .B(n14), .Z(n15) );
  NAND U27 ( .A(n13), .B(n15), .Z(n600) );
  NAND U28 ( .A(n627), .B(n629), .Z(n16) );
  XOR U29 ( .A(n627), .B(n629), .Z(n17) );
  NAND U30 ( .A(n17), .B(n628), .Z(n18) );
  NAND U31 ( .A(n16), .B(n18), .Z(n646) );
  XOR U32 ( .A(sreg[64]), .B(n619), .Z(n19) );
  NANDN U33 ( .A(n620), .B(n19), .Z(n20) );
  NAND U34 ( .A(sreg[64]), .B(n619), .Z(n21) );
  AND U35 ( .A(n20), .B(n21), .Z(n635) );
  NAND U36 ( .A(n692), .B(n691), .Z(n22) );
  XOR U37 ( .A(n692), .B(n691), .Z(n23) );
  NANDN U38 ( .A(sreg[68]), .B(n23), .Z(n24) );
  NAND U39 ( .A(n22), .B(n24), .Z(n711) );
  NAND U40 ( .A(n768), .B(n767), .Z(n25) );
  XOR U41 ( .A(n768), .B(n767), .Z(n26) );
  NANDN U42 ( .A(sreg[72]), .B(n26), .Z(n27) );
  NAND U43 ( .A(n25), .B(n27), .Z(n787) );
  NAND U44 ( .A(n844), .B(n843), .Z(n28) );
  XOR U45 ( .A(n844), .B(n843), .Z(n29) );
  NANDN U46 ( .A(sreg[76]), .B(n29), .Z(n30) );
  NAND U47 ( .A(n28), .B(n30), .Z(n863) );
  NAND U48 ( .A(n920), .B(n919), .Z(n31) );
  XOR U49 ( .A(n920), .B(n919), .Z(n32) );
  NANDN U50 ( .A(sreg[80]), .B(n32), .Z(n33) );
  NAND U51 ( .A(n31), .B(n33), .Z(n939) );
  NAND U52 ( .A(n996), .B(n995), .Z(n34) );
  XOR U53 ( .A(n996), .B(n995), .Z(n35) );
  NANDN U54 ( .A(sreg[84]), .B(n35), .Z(n36) );
  NAND U55 ( .A(n34), .B(n36), .Z(n1015) );
  NAND U56 ( .A(n1072), .B(n1071), .Z(n37) );
  XOR U57 ( .A(n1072), .B(n1071), .Z(n38) );
  NANDN U58 ( .A(sreg[88]), .B(n38), .Z(n39) );
  NAND U59 ( .A(n37), .B(n39), .Z(n1091) );
  NAND U60 ( .A(n1148), .B(n1147), .Z(n40) );
  XOR U61 ( .A(n1148), .B(n1147), .Z(n41) );
  NANDN U62 ( .A(sreg[92]), .B(n41), .Z(n42) );
  NAND U63 ( .A(n40), .B(n42), .Z(n1167) );
  NAND U64 ( .A(n1224), .B(n1223), .Z(n43) );
  XOR U65 ( .A(n1224), .B(n1223), .Z(n44) );
  NANDN U66 ( .A(sreg[96]), .B(n44), .Z(n45) );
  NAND U67 ( .A(n43), .B(n45), .Z(n1243) );
  NAND U68 ( .A(n1300), .B(n1299), .Z(n46) );
  XOR U69 ( .A(n1300), .B(n1299), .Z(n47) );
  NANDN U70 ( .A(sreg[100]), .B(n47), .Z(n48) );
  NAND U71 ( .A(n46), .B(n48), .Z(n1319) );
  NAND U72 ( .A(n1376), .B(n1375), .Z(n49) );
  XOR U73 ( .A(n1376), .B(n1375), .Z(n50) );
  NANDN U74 ( .A(sreg[104]), .B(n50), .Z(n51) );
  NAND U75 ( .A(n49), .B(n51), .Z(n1395) );
  NAND U76 ( .A(n1452), .B(n1451), .Z(n52) );
  XOR U77 ( .A(n1452), .B(n1451), .Z(n53) );
  NANDN U78 ( .A(sreg[108]), .B(n53), .Z(n54) );
  NAND U79 ( .A(n52), .B(n54), .Z(n1471) );
  NAND U80 ( .A(n1528), .B(n1527), .Z(n55) );
  XOR U81 ( .A(n1528), .B(n1527), .Z(n56) );
  NANDN U82 ( .A(sreg[112]), .B(n56), .Z(n57) );
  NAND U83 ( .A(n55), .B(n57), .Z(n1547) );
  NAND U84 ( .A(n1604), .B(n1603), .Z(n58) );
  XOR U85 ( .A(n1604), .B(n1603), .Z(n59) );
  NANDN U86 ( .A(sreg[116]), .B(n59), .Z(n60) );
  NAND U87 ( .A(n58), .B(n60), .Z(n1623) );
  NAND U88 ( .A(n1680), .B(n1679), .Z(n61) );
  XOR U89 ( .A(n1680), .B(n1679), .Z(n62) );
  NANDN U90 ( .A(sreg[120]), .B(n62), .Z(n63) );
  NAND U91 ( .A(n61), .B(n63), .Z(n1699) );
  AND U92 ( .A(n594), .B(n595), .Z(n609) );
  XOR U93 ( .A(n676), .B(n677), .Z(n64) );
  NANDN U94 ( .A(n678), .B(n64), .Z(n65) );
  NAND U95 ( .A(n676), .B(n677), .Z(n66) );
  AND U96 ( .A(n65), .B(n66), .Z(n708) );
  XOR U97 ( .A(n695), .B(n696), .Z(n67) );
  NANDN U98 ( .A(n697), .B(n67), .Z(n68) );
  NAND U99 ( .A(n695), .B(n696), .Z(n69) );
  AND U100 ( .A(n68), .B(n69), .Z(n727) );
  XOR U101 ( .A(n752), .B(n753), .Z(n70) );
  NANDN U102 ( .A(n754), .B(n70), .Z(n71) );
  NAND U103 ( .A(n752), .B(n753), .Z(n72) );
  AND U104 ( .A(n71), .B(n72), .Z(n784) );
  XOR U105 ( .A(n771), .B(n772), .Z(n73) );
  NANDN U106 ( .A(n773), .B(n73), .Z(n74) );
  NAND U107 ( .A(n771), .B(n772), .Z(n75) );
  AND U108 ( .A(n74), .B(n75), .Z(n803) );
  XOR U109 ( .A(n828), .B(n829), .Z(n76) );
  NANDN U110 ( .A(n830), .B(n76), .Z(n77) );
  NAND U111 ( .A(n828), .B(n829), .Z(n78) );
  AND U112 ( .A(n77), .B(n78), .Z(n860) );
  XOR U113 ( .A(n847), .B(n848), .Z(n79) );
  NANDN U114 ( .A(n849), .B(n79), .Z(n80) );
  NAND U115 ( .A(n847), .B(n848), .Z(n81) );
  AND U116 ( .A(n80), .B(n81), .Z(n879) );
  XOR U117 ( .A(n904), .B(n905), .Z(n82) );
  NANDN U118 ( .A(n906), .B(n82), .Z(n83) );
  NAND U119 ( .A(n904), .B(n905), .Z(n84) );
  AND U120 ( .A(n83), .B(n84), .Z(n936) );
  XOR U121 ( .A(n923), .B(n924), .Z(n85) );
  NANDN U122 ( .A(n925), .B(n85), .Z(n86) );
  NAND U123 ( .A(n923), .B(n924), .Z(n87) );
  AND U124 ( .A(n86), .B(n87), .Z(n955) );
  XOR U125 ( .A(n980), .B(n981), .Z(n88) );
  NANDN U126 ( .A(n982), .B(n88), .Z(n89) );
  NAND U127 ( .A(n980), .B(n981), .Z(n90) );
  AND U128 ( .A(n89), .B(n90), .Z(n1012) );
  XOR U129 ( .A(n999), .B(n1000), .Z(n91) );
  NANDN U130 ( .A(n1001), .B(n91), .Z(n92) );
  NAND U131 ( .A(n999), .B(n1000), .Z(n93) );
  AND U132 ( .A(n92), .B(n93), .Z(n1031) );
  XOR U133 ( .A(n1056), .B(n1057), .Z(n94) );
  NANDN U134 ( .A(n1058), .B(n94), .Z(n95) );
  NAND U135 ( .A(n1056), .B(n1057), .Z(n96) );
  AND U136 ( .A(n95), .B(n96), .Z(n1088) );
  XOR U137 ( .A(n1075), .B(n1076), .Z(n97) );
  NANDN U138 ( .A(n1077), .B(n97), .Z(n98) );
  NAND U139 ( .A(n1075), .B(n1076), .Z(n99) );
  AND U140 ( .A(n98), .B(n99), .Z(n1107) );
  XOR U141 ( .A(n1132), .B(n1133), .Z(n100) );
  NANDN U142 ( .A(n1134), .B(n100), .Z(n101) );
  NAND U143 ( .A(n1132), .B(n1133), .Z(n102) );
  AND U144 ( .A(n101), .B(n102), .Z(n1164) );
  XOR U145 ( .A(n1151), .B(n1152), .Z(n103) );
  NANDN U146 ( .A(n1153), .B(n103), .Z(n104) );
  NAND U147 ( .A(n1151), .B(n1152), .Z(n105) );
  AND U148 ( .A(n104), .B(n105), .Z(n1183) );
  XOR U149 ( .A(n1208), .B(n1209), .Z(n106) );
  NANDN U150 ( .A(n1210), .B(n106), .Z(n107) );
  NAND U151 ( .A(n1208), .B(n1209), .Z(n108) );
  AND U152 ( .A(n107), .B(n108), .Z(n1240) );
  XOR U153 ( .A(n1227), .B(n1228), .Z(n109) );
  NANDN U154 ( .A(n1229), .B(n109), .Z(n110) );
  NAND U155 ( .A(n1227), .B(n1228), .Z(n111) );
  AND U156 ( .A(n110), .B(n111), .Z(n1259) );
  XOR U157 ( .A(n1284), .B(n1285), .Z(n112) );
  NANDN U158 ( .A(n1286), .B(n112), .Z(n113) );
  NAND U159 ( .A(n1284), .B(n1285), .Z(n114) );
  AND U160 ( .A(n113), .B(n114), .Z(n1316) );
  XOR U161 ( .A(n1303), .B(n1304), .Z(n115) );
  NANDN U162 ( .A(n1305), .B(n115), .Z(n116) );
  NAND U163 ( .A(n1303), .B(n1304), .Z(n117) );
  AND U164 ( .A(n116), .B(n117), .Z(n1335) );
  XOR U165 ( .A(n1360), .B(n1361), .Z(n118) );
  NANDN U166 ( .A(n1362), .B(n118), .Z(n119) );
  NAND U167 ( .A(n1360), .B(n1361), .Z(n120) );
  AND U168 ( .A(n119), .B(n120), .Z(n1392) );
  XOR U169 ( .A(n1379), .B(n1380), .Z(n121) );
  NANDN U170 ( .A(n1381), .B(n121), .Z(n122) );
  NAND U171 ( .A(n1379), .B(n1380), .Z(n123) );
  AND U172 ( .A(n122), .B(n123), .Z(n1411) );
  XOR U173 ( .A(n1436), .B(n1437), .Z(n124) );
  NANDN U174 ( .A(n1438), .B(n124), .Z(n125) );
  NAND U175 ( .A(n1436), .B(n1437), .Z(n126) );
  AND U176 ( .A(n125), .B(n126), .Z(n1468) );
  XOR U177 ( .A(n1455), .B(n1456), .Z(n127) );
  NANDN U178 ( .A(n1457), .B(n127), .Z(n128) );
  NAND U179 ( .A(n1455), .B(n1456), .Z(n129) );
  AND U180 ( .A(n128), .B(n129), .Z(n1487) );
  XOR U181 ( .A(n1512), .B(n1513), .Z(n130) );
  NANDN U182 ( .A(n1514), .B(n130), .Z(n131) );
  NAND U183 ( .A(n1512), .B(n1513), .Z(n132) );
  AND U184 ( .A(n131), .B(n132), .Z(n1544) );
  XOR U185 ( .A(n1531), .B(n1532), .Z(n133) );
  NANDN U186 ( .A(n1533), .B(n133), .Z(n134) );
  NAND U187 ( .A(n1531), .B(n1532), .Z(n135) );
  AND U188 ( .A(n134), .B(n135), .Z(n1563) );
  XOR U189 ( .A(n1588), .B(n1589), .Z(n136) );
  NANDN U190 ( .A(n1590), .B(n136), .Z(n137) );
  NAND U191 ( .A(n1588), .B(n1589), .Z(n138) );
  AND U192 ( .A(n137), .B(n138), .Z(n1620) );
  XOR U193 ( .A(n1607), .B(n1608), .Z(n139) );
  NANDN U194 ( .A(n1609), .B(n139), .Z(n140) );
  NAND U195 ( .A(n1607), .B(n1608), .Z(n141) );
  AND U196 ( .A(n140), .B(n141), .Z(n1639) );
  XOR U197 ( .A(n1664), .B(n1665), .Z(n142) );
  NANDN U198 ( .A(n1666), .B(n142), .Z(n143) );
  NAND U199 ( .A(n1664), .B(n1665), .Z(n144) );
  AND U200 ( .A(n143), .B(n144), .Z(n1696) );
  XOR U201 ( .A(n1683), .B(n1684), .Z(n145) );
  NANDN U202 ( .A(n1685), .B(n145), .Z(n146) );
  NAND U203 ( .A(n1683), .B(n1684), .Z(n147) );
  AND U204 ( .A(n146), .B(n147), .Z(n1715) );
  NANDN U205 ( .A(n601), .B(n624), .Z(n148) );
  ANDN U206 ( .B(n148), .A(n602), .Z(n612) );
  NAND U207 ( .A(n1741), .B(n1739), .Z(n149) );
  XOR U208 ( .A(n1741), .B(n1739), .Z(n150) );
  NANDN U209 ( .A(n1740), .B(n150), .Z(n151) );
  NAND U210 ( .A(n149), .B(n151), .Z(n1752) );
  NAND U211 ( .A(n635), .B(n634), .Z(n152) );
  XOR U212 ( .A(n635), .B(n634), .Z(n153) );
  NANDN U213 ( .A(sreg[65]), .B(n153), .Z(n154) );
  NAND U214 ( .A(n152), .B(n154), .Z(n654) );
  NAND U215 ( .A(n711), .B(n710), .Z(n155) );
  XOR U216 ( .A(n711), .B(n710), .Z(n156) );
  NANDN U217 ( .A(sreg[69]), .B(n156), .Z(n157) );
  NAND U218 ( .A(n155), .B(n157), .Z(n730) );
  NAND U219 ( .A(n787), .B(n786), .Z(n158) );
  XOR U220 ( .A(n787), .B(n786), .Z(n159) );
  NANDN U221 ( .A(sreg[73]), .B(n159), .Z(n160) );
  NAND U222 ( .A(n158), .B(n160), .Z(n806) );
  NAND U223 ( .A(n863), .B(n862), .Z(n161) );
  XOR U224 ( .A(n863), .B(n862), .Z(n162) );
  NANDN U225 ( .A(sreg[77]), .B(n162), .Z(n163) );
  NAND U226 ( .A(n161), .B(n163), .Z(n882) );
  NAND U227 ( .A(n939), .B(n938), .Z(n164) );
  XOR U228 ( .A(n939), .B(n938), .Z(n165) );
  NANDN U229 ( .A(sreg[81]), .B(n165), .Z(n166) );
  NAND U230 ( .A(n164), .B(n166), .Z(n958) );
  NAND U231 ( .A(n1015), .B(n1014), .Z(n167) );
  XOR U232 ( .A(n1015), .B(n1014), .Z(n168) );
  NANDN U233 ( .A(sreg[85]), .B(n168), .Z(n169) );
  NAND U234 ( .A(n167), .B(n169), .Z(n1034) );
  NAND U235 ( .A(n1091), .B(n1090), .Z(n170) );
  XOR U236 ( .A(n1091), .B(n1090), .Z(n171) );
  NANDN U237 ( .A(sreg[89]), .B(n171), .Z(n172) );
  NAND U238 ( .A(n170), .B(n172), .Z(n1110) );
  NAND U239 ( .A(n1167), .B(n1166), .Z(n173) );
  XOR U240 ( .A(n1167), .B(n1166), .Z(n174) );
  NANDN U241 ( .A(sreg[93]), .B(n174), .Z(n175) );
  NAND U242 ( .A(n173), .B(n175), .Z(n1186) );
  NAND U243 ( .A(n1243), .B(n1242), .Z(n176) );
  XOR U244 ( .A(n1243), .B(n1242), .Z(n177) );
  NANDN U245 ( .A(sreg[97]), .B(n177), .Z(n178) );
  NAND U246 ( .A(n176), .B(n178), .Z(n1262) );
  NAND U247 ( .A(n1319), .B(n1318), .Z(n179) );
  XOR U248 ( .A(n1319), .B(n1318), .Z(n180) );
  NANDN U249 ( .A(sreg[101]), .B(n180), .Z(n181) );
  NAND U250 ( .A(n179), .B(n181), .Z(n1338) );
  NAND U251 ( .A(n1395), .B(n1394), .Z(n182) );
  XOR U252 ( .A(n1395), .B(n1394), .Z(n183) );
  NANDN U253 ( .A(sreg[105]), .B(n183), .Z(n184) );
  NAND U254 ( .A(n182), .B(n184), .Z(n1414) );
  NAND U255 ( .A(n1471), .B(n1470), .Z(n185) );
  XOR U256 ( .A(n1471), .B(n1470), .Z(n186) );
  NANDN U257 ( .A(sreg[109]), .B(n186), .Z(n187) );
  NAND U258 ( .A(n185), .B(n187), .Z(n1490) );
  NAND U259 ( .A(n1547), .B(n1546), .Z(n188) );
  XOR U260 ( .A(n1547), .B(n1546), .Z(n189) );
  NANDN U261 ( .A(sreg[113]), .B(n189), .Z(n190) );
  NAND U262 ( .A(n188), .B(n190), .Z(n1566) );
  NAND U263 ( .A(n1623), .B(n1622), .Z(n191) );
  XOR U264 ( .A(n1623), .B(n1622), .Z(n192) );
  NANDN U265 ( .A(sreg[117]), .B(n192), .Z(n193) );
  NAND U266 ( .A(n191), .B(n193), .Z(n1642) );
  NAND U267 ( .A(n1699), .B(n1698), .Z(n194) );
  XOR U268 ( .A(n1699), .B(n1698), .Z(n195) );
  NANDN U269 ( .A(sreg[121]), .B(n195), .Z(n196) );
  NAND U270 ( .A(n194), .B(n196), .Z(n1718) );
  XOR U271 ( .A(n638), .B(n639), .Z(n197) );
  NANDN U272 ( .A(n640), .B(n197), .Z(n198) );
  NAND U273 ( .A(n638), .B(n639), .Z(n199) );
  AND U274 ( .A(n198), .B(n199), .Z(n670) );
  XOR U275 ( .A(n657), .B(n658), .Z(n200) );
  NANDN U276 ( .A(n659), .B(n200), .Z(n201) );
  NAND U277 ( .A(n657), .B(n658), .Z(n202) );
  AND U278 ( .A(n201), .B(n202), .Z(n689) );
  XOR U279 ( .A(n714), .B(n715), .Z(n203) );
  NANDN U280 ( .A(n716), .B(n203), .Z(n204) );
  NAND U281 ( .A(n714), .B(n715), .Z(n205) );
  AND U282 ( .A(n204), .B(n205), .Z(n746) );
  XOR U283 ( .A(n733), .B(n734), .Z(n206) );
  NANDN U284 ( .A(n735), .B(n206), .Z(n207) );
  NAND U285 ( .A(n733), .B(n734), .Z(n208) );
  AND U286 ( .A(n207), .B(n208), .Z(n765) );
  XOR U287 ( .A(n790), .B(n791), .Z(n209) );
  NANDN U288 ( .A(n792), .B(n209), .Z(n210) );
  NAND U289 ( .A(n790), .B(n791), .Z(n211) );
  AND U290 ( .A(n210), .B(n211), .Z(n822) );
  XOR U291 ( .A(n809), .B(n810), .Z(n212) );
  NANDN U292 ( .A(n811), .B(n212), .Z(n213) );
  NAND U293 ( .A(n809), .B(n810), .Z(n214) );
  AND U294 ( .A(n213), .B(n214), .Z(n841) );
  XOR U295 ( .A(n866), .B(n867), .Z(n215) );
  NANDN U296 ( .A(n868), .B(n215), .Z(n216) );
  NAND U297 ( .A(n866), .B(n867), .Z(n217) );
  AND U298 ( .A(n216), .B(n217), .Z(n898) );
  XOR U299 ( .A(n885), .B(n886), .Z(n218) );
  NANDN U300 ( .A(n887), .B(n218), .Z(n219) );
  NAND U301 ( .A(n885), .B(n886), .Z(n220) );
  AND U302 ( .A(n219), .B(n220), .Z(n917) );
  XOR U303 ( .A(n942), .B(n943), .Z(n221) );
  NANDN U304 ( .A(n944), .B(n221), .Z(n222) );
  NAND U305 ( .A(n942), .B(n943), .Z(n223) );
  AND U306 ( .A(n222), .B(n223), .Z(n974) );
  XOR U307 ( .A(n961), .B(n962), .Z(n224) );
  NANDN U308 ( .A(n963), .B(n224), .Z(n225) );
  NAND U309 ( .A(n961), .B(n962), .Z(n226) );
  AND U310 ( .A(n225), .B(n226), .Z(n993) );
  XOR U311 ( .A(n1018), .B(n1019), .Z(n227) );
  NANDN U312 ( .A(n1020), .B(n227), .Z(n228) );
  NAND U313 ( .A(n1018), .B(n1019), .Z(n229) );
  AND U314 ( .A(n228), .B(n229), .Z(n1050) );
  XOR U315 ( .A(n1037), .B(n1038), .Z(n230) );
  NANDN U316 ( .A(n1039), .B(n230), .Z(n231) );
  NAND U317 ( .A(n1037), .B(n1038), .Z(n232) );
  AND U318 ( .A(n231), .B(n232), .Z(n1069) );
  XOR U319 ( .A(n1094), .B(n1095), .Z(n233) );
  NANDN U320 ( .A(n1096), .B(n233), .Z(n234) );
  NAND U321 ( .A(n1094), .B(n1095), .Z(n235) );
  AND U322 ( .A(n234), .B(n235), .Z(n1126) );
  XOR U323 ( .A(n1113), .B(n1114), .Z(n236) );
  NANDN U324 ( .A(n1115), .B(n236), .Z(n237) );
  NAND U325 ( .A(n1113), .B(n1114), .Z(n238) );
  AND U326 ( .A(n237), .B(n238), .Z(n1145) );
  XOR U327 ( .A(n1170), .B(n1171), .Z(n239) );
  NANDN U328 ( .A(n1172), .B(n239), .Z(n240) );
  NAND U329 ( .A(n1170), .B(n1171), .Z(n241) );
  AND U330 ( .A(n240), .B(n241), .Z(n1202) );
  XOR U331 ( .A(n1189), .B(n1190), .Z(n242) );
  NANDN U332 ( .A(n1191), .B(n242), .Z(n243) );
  NAND U333 ( .A(n1189), .B(n1190), .Z(n244) );
  AND U334 ( .A(n243), .B(n244), .Z(n1221) );
  XOR U335 ( .A(n1246), .B(n1247), .Z(n245) );
  NANDN U336 ( .A(n1248), .B(n245), .Z(n246) );
  NAND U337 ( .A(n1246), .B(n1247), .Z(n247) );
  AND U338 ( .A(n246), .B(n247), .Z(n1278) );
  XOR U339 ( .A(n1265), .B(n1266), .Z(n248) );
  NANDN U340 ( .A(n1267), .B(n248), .Z(n249) );
  NAND U341 ( .A(n1265), .B(n1266), .Z(n250) );
  AND U342 ( .A(n249), .B(n250), .Z(n1297) );
  XOR U343 ( .A(n1322), .B(n1323), .Z(n251) );
  NANDN U344 ( .A(n1324), .B(n251), .Z(n252) );
  NAND U345 ( .A(n1322), .B(n1323), .Z(n253) );
  AND U346 ( .A(n252), .B(n253), .Z(n1354) );
  XOR U347 ( .A(n1341), .B(n1342), .Z(n254) );
  NANDN U348 ( .A(n1343), .B(n254), .Z(n255) );
  NAND U349 ( .A(n1341), .B(n1342), .Z(n256) );
  AND U350 ( .A(n255), .B(n256), .Z(n1373) );
  XOR U351 ( .A(n1398), .B(n1399), .Z(n257) );
  NANDN U352 ( .A(n1400), .B(n257), .Z(n258) );
  NAND U353 ( .A(n1398), .B(n1399), .Z(n259) );
  AND U354 ( .A(n258), .B(n259), .Z(n1430) );
  XOR U355 ( .A(n1417), .B(n1418), .Z(n260) );
  NANDN U356 ( .A(n1419), .B(n260), .Z(n261) );
  NAND U357 ( .A(n1417), .B(n1418), .Z(n262) );
  AND U358 ( .A(n261), .B(n262), .Z(n1449) );
  XOR U359 ( .A(n1474), .B(n1475), .Z(n263) );
  NANDN U360 ( .A(n1476), .B(n263), .Z(n264) );
  NAND U361 ( .A(n1474), .B(n1475), .Z(n265) );
  AND U362 ( .A(n264), .B(n265), .Z(n1506) );
  XOR U363 ( .A(n1493), .B(n1494), .Z(n266) );
  NANDN U364 ( .A(n1495), .B(n266), .Z(n267) );
  NAND U365 ( .A(n1493), .B(n1494), .Z(n268) );
  AND U366 ( .A(n267), .B(n268), .Z(n1525) );
  XOR U367 ( .A(n1550), .B(n1551), .Z(n269) );
  NANDN U368 ( .A(n1552), .B(n269), .Z(n270) );
  NAND U369 ( .A(n1550), .B(n1551), .Z(n271) );
  AND U370 ( .A(n270), .B(n271), .Z(n1582) );
  XOR U371 ( .A(n1569), .B(n1570), .Z(n272) );
  NANDN U372 ( .A(n1571), .B(n272), .Z(n273) );
  NAND U373 ( .A(n1569), .B(n1570), .Z(n274) );
  AND U374 ( .A(n273), .B(n274), .Z(n1601) );
  XOR U375 ( .A(n1626), .B(n1627), .Z(n275) );
  NANDN U376 ( .A(n1628), .B(n275), .Z(n276) );
  NAND U377 ( .A(n1626), .B(n1627), .Z(n277) );
  AND U378 ( .A(n276), .B(n277), .Z(n1658) );
  XOR U379 ( .A(n1645), .B(n1646), .Z(n278) );
  NANDN U380 ( .A(n1647), .B(n278), .Z(n279) );
  NAND U381 ( .A(n1645), .B(n1646), .Z(n280) );
  AND U382 ( .A(n279), .B(n280), .Z(n1677) );
  NAND U383 ( .A(n613), .B(n614), .Z(n281) );
  XOR U384 ( .A(n613), .B(n614), .Z(n282) );
  NANDN U385 ( .A(n612), .B(n282), .Z(n283) );
  NAND U386 ( .A(n281), .B(n283), .Z(n629) );
  NAND U387 ( .A(n631), .B(n632), .Z(n284) );
  XOR U388 ( .A(n631), .B(n632), .Z(n285) );
  NANDN U389 ( .A(n630), .B(n285), .Z(n286) );
  NAND U390 ( .A(n284), .B(n286), .Z(n644) );
  NAND U391 ( .A(n707), .B(n708), .Z(n287) );
  XOR U392 ( .A(n707), .B(n708), .Z(n288) );
  NANDN U393 ( .A(n706), .B(n288), .Z(n289) );
  NAND U394 ( .A(n287), .B(n289), .Z(n720) );
  NAND U395 ( .A(n783), .B(n784), .Z(n290) );
  XOR U396 ( .A(n783), .B(n784), .Z(n291) );
  NANDN U397 ( .A(n782), .B(n291), .Z(n292) );
  NAND U398 ( .A(n290), .B(n292), .Z(n796) );
  NAND U399 ( .A(n859), .B(n860), .Z(n293) );
  XOR U400 ( .A(n859), .B(n860), .Z(n294) );
  NANDN U401 ( .A(n858), .B(n294), .Z(n295) );
  NAND U402 ( .A(n293), .B(n295), .Z(n872) );
  NAND U403 ( .A(n935), .B(n936), .Z(n296) );
  XOR U404 ( .A(n935), .B(n936), .Z(n297) );
  NANDN U405 ( .A(n934), .B(n297), .Z(n298) );
  NAND U406 ( .A(n296), .B(n298), .Z(n948) );
  NAND U407 ( .A(n1011), .B(n1012), .Z(n299) );
  XOR U408 ( .A(n1011), .B(n1012), .Z(n300) );
  NANDN U409 ( .A(n1010), .B(n300), .Z(n301) );
  NAND U410 ( .A(n299), .B(n301), .Z(n1024) );
  NAND U411 ( .A(n1087), .B(n1088), .Z(n302) );
  XOR U412 ( .A(n1087), .B(n1088), .Z(n303) );
  NANDN U413 ( .A(n1086), .B(n303), .Z(n304) );
  NAND U414 ( .A(n302), .B(n304), .Z(n1100) );
  NAND U415 ( .A(n1163), .B(n1164), .Z(n305) );
  XOR U416 ( .A(n1163), .B(n1164), .Z(n306) );
  NANDN U417 ( .A(n1162), .B(n306), .Z(n307) );
  NAND U418 ( .A(n305), .B(n307), .Z(n1176) );
  NAND U419 ( .A(n1239), .B(n1240), .Z(n308) );
  XOR U420 ( .A(n1239), .B(n1240), .Z(n309) );
  NANDN U421 ( .A(n1238), .B(n309), .Z(n310) );
  NAND U422 ( .A(n308), .B(n310), .Z(n1252) );
  NAND U423 ( .A(n1315), .B(n1316), .Z(n311) );
  XOR U424 ( .A(n1315), .B(n1316), .Z(n312) );
  NANDN U425 ( .A(n1314), .B(n312), .Z(n313) );
  NAND U426 ( .A(n311), .B(n313), .Z(n1328) );
  NAND U427 ( .A(n1391), .B(n1392), .Z(n314) );
  XOR U428 ( .A(n1391), .B(n1392), .Z(n315) );
  NANDN U429 ( .A(n1390), .B(n315), .Z(n316) );
  NAND U430 ( .A(n314), .B(n316), .Z(n1404) );
  NAND U431 ( .A(n1467), .B(n1468), .Z(n317) );
  XOR U432 ( .A(n1467), .B(n1468), .Z(n318) );
  NANDN U433 ( .A(n1466), .B(n318), .Z(n319) );
  NAND U434 ( .A(n317), .B(n319), .Z(n1480) );
  NAND U435 ( .A(n1543), .B(n1544), .Z(n320) );
  XOR U436 ( .A(n1543), .B(n1544), .Z(n321) );
  NANDN U437 ( .A(n1542), .B(n321), .Z(n322) );
  NAND U438 ( .A(n320), .B(n322), .Z(n1556) );
  NAND U439 ( .A(n1619), .B(n1620), .Z(n323) );
  XOR U440 ( .A(n1619), .B(n1620), .Z(n324) );
  NANDN U441 ( .A(n1618), .B(n324), .Z(n325) );
  NAND U442 ( .A(n323), .B(n325), .Z(n1632) );
  NAND U443 ( .A(n1695), .B(n1696), .Z(n326) );
  XOR U444 ( .A(n1695), .B(n1696), .Z(n327) );
  NANDN U445 ( .A(n1694), .B(n327), .Z(n328) );
  NAND U446 ( .A(n326), .B(n328), .Z(n1708) );
  NAND U447 ( .A(n1723), .B(n1724), .Z(n329) );
  XOR U448 ( .A(n1723), .B(n1724), .Z(n330) );
  NANDN U449 ( .A(n1722), .B(n330), .Z(n331) );
  NAND U450 ( .A(n329), .B(n331), .Z(n1739) );
  XOR U451 ( .A(n1748), .B(n1747), .Z(n332) );
  NANDN U452 ( .A(n1746), .B(n332), .Z(n333) );
  NAND U453 ( .A(n1748), .B(n1747), .Z(n334) );
  AND U454 ( .A(n333), .B(n334), .Z(n1750) );
  XOR U455 ( .A(sreg[63]), .B(n604), .Z(n335) );
  NANDN U456 ( .A(n605), .B(n335), .Z(n336) );
  NAND U457 ( .A(sreg[63]), .B(n604), .Z(n337) );
  AND U458 ( .A(n336), .B(n337), .Z(n620) );
  NAND U459 ( .A(n673), .B(n672), .Z(n338) );
  XOR U460 ( .A(n673), .B(n672), .Z(n339) );
  NANDN U461 ( .A(sreg[67]), .B(n339), .Z(n340) );
  NAND U462 ( .A(n338), .B(n340), .Z(n692) );
  NAND U463 ( .A(n749), .B(n748), .Z(n341) );
  XOR U464 ( .A(n749), .B(n748), .Z(n342) );
  NANDN U465 ( .A(sreg[71]), .B(n342), .Z(n343) );
  NAND U466 ( .A(n341), .B(n343), .Z(n768) );
  NAND U467 ( .A(n825), .B(n824), .Z(n344) );
  XOR U468 ( .A(n825), .B(n824), .Z(n345) );
  NANDN U469 ( .A(sreg[75]), .B(n345), .Z(n346) );
  NAND U470 ( .A(n344), .B(n346), .Z(n844) );
  NAND U471 ( .A(n901), .B(n900), .Z(n347) );
  XOR U472 ( .A(n901), .B(n900), .Z(n348) );
  NANDN U473 ( .A(sreg[79]), .B(n348), .Z(n349) );
  NAND U474 ( .A(n347), .B(n349), .Z(n920) );
  NAND U475 ( .A(n977), .B(n976), .Z(n350) );
  XOR U476 ( .A(n977), .B(n976), .Z(n351) );
  NANDN U477 ( .A(sreg[83]), .B(n351), .Z(n352) );
  NAND U478 ( .A(n350), .B(n352), .Z(n996) );
  NAND U479 ( .A(n1053), .B(n1052), .Z(n353) );
  XOR U480 ( .A(n1053), .B(n1052), .Z(n354) );
  NANDN U481 ( .A(sreg[87]), .B(n354), .Z(n355) );
  NAND U482 ( .A(n353), .B(n355), .Z(n1072) );
  NAND U483 ( .A(n1129), .B(n1128), .Z(n356) );
  XOR U484 ( .A(n1129), .B(n1128), .Z(n357) );
  NANDN U485 ( .A(sreg[91]), .B(n357), .Z(n358) );
  NAND U486 ( .A(n356), .B(n358), .Z(n1148) );
  NAND U487 ( .A(n1205), .B(n1204), .Z(n359) );
  XOR U488 ( .A(n1205), .B(n1204), .Z(n360) );
  NANDN U489 ( .A(sreg[95]), .B(n360), .Z(n361) );
  NAND U490 ( .A(n359), .B(n361), .Z(n1224) );
  NAND U491 ( .A(n1281), .B(n1280), .Z(n362) );
  XOR U492 ( .A(n1281), .B(n1280), .Z(n363) );
  NANDN U493 ( .A(sreg[99]), .B(n363), .Z(n364) );
  NAND U494 ( .A(n362), .B(n364), .Z(n1300) );
  NAND U495 ( .A(n1357), .B(n1356), .Z(n365) );
  XOR U496 ( .A(n1357), .B(n1356), .Z(n366) );
  NANDN U497 ( .A(sreg[103]), .B(n366), .Z(n367) );
  NAND U498 ( .A(n365), .B(n367), .Z(n1376) );
  NAND U499 ( .A(n1433), .B(n1432), .Z(n368) );
  XOR U500 ( .A(n1433), .B(n1432), .Z(n369) );
  NANDN U501 ( .A(sreg[107]), .B(n369), .Z(n370) );
  NAND U502 ( .A(n368), .B(n370), .Z(n1452) );
  NAND U503 ( .A(n1509), .B(n1508), .Z(n371) );
  XOR U504 ( .A(n1509), .B(n1508), .Z(n372) );
  NANDN U505 ( .A(sreg[111]), .B(n372), .Z(n373) );
  NAND U506 ( .A(n371), .B(n373), .Z(n1528) );
  NAND U507 ( .A(n1585), .B(n1584), .Z(n374) );
  XOR U508 ( .A(n1585), .B(n1584), .Z(n375) );
  NANDN U509 ( .A(sreg[115]), .B(n375), .Z(n376) );
  NAND U510 ( .A(n374), .B(n376), .Z(n1604) );
  NAND U511 ( .A(n1661), .B(n1660), .Z(n377) );
  XOR U512 ( .A(n1661), .B(n1660), .Z(n378) );
  NANDN U513 ( .A(sreg[119]), .B(n378), .Z(n379) );
  NAND U514 ( .A(n377), .B(n379), .Z(n1680) );
  NAND U515 ( .A(n1721), .B(n1720), .Z(n380) );
  XOR U516 ( .A(n1721), .B(n1720), .Z(n381) );
  NANDN U517 ( .A(sreg[123]), .B(n381), .Z(n382) );
  NAND U518 ( .A(n380), .B(n382), .Z(n1737) );
  NAND U519 ( .A(n599), .B(n600), .Z(n383) );
  XOR U520 ( .A(n599), .B(n600), .Z(n384) );
  NANDN U521 ( .A(n598), .B(n384), .Z(n385) );
  NAND U522 ( .A(n383), .B(n385), .Z(n613) );
  NAND U523 ( .A(n616), .B(n617), .Z(n386) );
  XOR U524 ( .A(n616), .B(n617), .Z(n387) );
  NANDN U525 ( .A(n615), .B(n387), .Z(n388) );
  NAND U526 ( .A(n386), .B(n388), .Z(n628) );
  NAND U527 ( .A(n650), .B(n651), .Z(n389) );
  XOR U528 ( .A(n650), .B(n651), .Z(n390) );
  NANDN U529 ( .A(n649), .B(n390), .Z(n391) );
  NAND U530 ( .A(n389), .B(n391), .Z(n663) );
  NAND U531 ( .A(n669), .B(n670), .Z(n392) );
  XOR U532 ( .A(n669), .B(n670), .Z(n393) );
  NANDN U533 ( .A(n668), .B(n393), .Z(n394) );
  NAND U534 ( .A(n392), .B(n394), .Z(n682) );
  NAND U535 ( .A(n688), .B(n689), .Z(n395) );
  XOR U536 ( .A(n688), .B(n689), .Z(n396) );
  NANDN U537 ( .A(n687), .B(n396), .Z(n397) );
  NAND U538 ( .A(n395), .B(n397), .Z(n701) );
  NAND U539 ( .A(n726), .B(n727), .Z(n398) );
  XOR U540 ( .A(n726), .B(n727), .Z(n399) );
  NANDN U541 ( .A(n725), .B(n399), .Z(n400) );
  NAND U542 ( .A(n398), .B(n400), .Z(n739) );
  NAND U543 ( .A(n745), .B(n746), .Z(n401) );
  XOR U544 ( .A(n745), .B(n746), .Z(n402) );
  NANDN U545 ( .A(n744), .B(n402), .Z(n403) );
  NAND U546 ( .A(n401), .B(n403), .Z(n758) );
  NAND U547 ( .A(n764), .B(n765), .Z(n404) );
  XOR U548 ( .A(n764), .B(n765), .Z(n405) );
  NANDN U549 ( .A(n763), .B(n405), .Z(n406) );
  NAND U550 ( .A(n404), .B(n406), .Z(n777) );
  NAND U551 ( .A(n802), .B(n803), .Z(n407) );
  XOR U552 ( .A(n802), .B(n803), .Z(n408) );
  NANDN U553 ( .A(n801), .B(n408), .Z(n409) );
  NAND U554 ( .A(n407), .B(n409), .Z(n815) );
  NAND U555 ( .A(n821), .B(n822), .Z(n410) );
  XOR U556 ( .A(n821), .B(n822), .Z(n411) );
  NANDN U557 ( .A(n820), .B(n411), .Z(n412) );
  NAND U558 ( .A(n410), .B(n412), .Z(n834) );
  NAND U559 ( .A(n840), .B(n841), .Z(n413) );
  XOR U560 ( .A(n840), .B(n841), .Z(n414) );
  NANDN U561 ( .A(n839), .B(n414), .Z(n415) );
  NAND U562 ( .A(n413), .B(n415), .Z(n853) );
  NAND U563 ( .A(n878), .B(n879), .Z(n416) );
  XOR U564 ( .A(n878), .B(n879), .Z(n417) );
  NANDN U565 ( .A(n877), .B(n417), .Z(n418) );
  NAND U566 ( .A(n416), .B(n418), .Z(n891) );
  NAND U567 ( .A(n897), .B(n898), .Z(n419) );
  XOR U568 ( .A(n897), .B(n898), .Z(n420) );
  NANDN U569 ( .A(n896), .B(n420), .Z(n421) );
  NAND U570 ( .A(n419), .B(n421), .Z(n910) );
  NAND U571 ( .A(n916), .B(n917), .Z(n422) );
  XOR U572 ( .A(n916), .B(n917), .Z(n423) );
  NANDN U573 ( .A(n915), .B(n423), .Z(n424) );
  NAND U574 ( .A(n422), .B(n424), .Z(n929) );
  NAND U575 ( .A(n954), .B(n955), .Z(n425) );
  XOR U576 ( .A(n954), .B(n955), .Z(n426) );
  NANDN U577 ( .A(n953), .B(n426), .Z(n427) );
  NAND U578 ( .A(n425), .B(n427), .Z(n967) );
  NAND U579 ( .A(n973), .B(n974), .Z(n428) );
  XOR U580 ( .A(n973), .B(n974), .Z(n429) );
  NANDN U581 ( .A(n972), .B(n429), .Z(n430) );
  NAND U582 ( .A(n428), .B(n430), .Z(n986) );
  NAND U583 ( .A(n992), .B(n993), .Z(n431) );
  XOR U584 ( .A(n992), .B(n993), .Z(n432) );
  NANDN U585 ( .A(n991), .B(n432), .Z(n433) );
  NAND U586 ( .A(n431), .B(n433), .Z(n1005) );
  NAND U587 ( .A(n1030), .B(n1031), .Z(n434) );
  XOR U588 ( .A(n1030), .B(n1031), .Z(n435) );
  NANDN U589 ( .A(n1029), .B(n435), .Z(n436) );
  NAND U590 ( .A(n434), .B(n436), .Z(n1043) );
  NAND U591 ( .A(n1049), .B(n1050), .Z(n437) );
  XOR U592 ( .A(n1049), .B(n1050), .Z(n438) );
  NANDN U593 ( .A(n1048), .B(n438), .Z(n439) );
  NAND U594 ( .A(n437), .B(n439), .Z(n1062) );
  NAND U595 ( .A(n1068), .B(n1069), .Z(n440) );
  XOR U596 ( .A(n1068), .B(n1069), .Z(n441) );
  NANDN U597 ( .A(n1067), .B(n441), .Z(n442) );
  NAND U598 ( .A(n440), .B(n442), .Z(n1081) );
  NAND U599 ( .A(n1106), .B(n1107), .Z(n443) );
  XOR U600 ( .A(n1106), .B(n1107), .Z(n444) );
  NANDN U601 ( .A(n1105), .B(n444), .Z(n445) );
  NAND U602 ( .A(n443), .B(n445), .Z(n1119) );
  NAND U603 ( .A(n1125), .B(n1126), .Z(n446) );
  XOR U604 ( .A(n1125), .B(n1126), .Z(n447) );
  NANDN U605 ( .A(n1124), .B(n447), .Z(n448) );
  NAND U606 ( .A(n446), .B(n448), .Z(n1138) );
  NAND U607 ( .A(n1144), .B(n1145), .Z(n449) );
  XOR U608 ( .A(n1144), .B(n1145), .Z(n450) );
  NANDN U609 ( .A(n1143), .B(n450), .Z(n451) );
  NAND U610 ( .A(n449), .B(n451), .Z(n1157) );
  NAND U611 ( .A(n1182), .B(n1183), .Z(n452) );
  XOR U612 ( .A(n1182), .B(n1183), .Z(n453) );
  NANDN U613 ( .A(n1181), .B(n453), .Z(n454) );
  NAND U614 ( .A(n452), .B(n454), .Z(n1195) );
  NAND U615 ( .A(n1201), .B(n1202), .Z(n455) );
  XOR U616 ( .A(n1201), .B(n1202), .Z(n456) );
  NANDN U617 ( .A(n1200), .B(n456), .Z(n457) );
  NAND U618 ( .A(n455), .B(n457), .Z(n1214) );
  NAND U619 ( .A(n1220), .B(n1221), .Z(n458) );
  XOR U620 ( .A(n1220), .B(n1221), .Z(n459) );
  NANDN U621 ( .A(n1219), .B(n459), .Z(n460) );
  NAND U622 ( .A(n458), .B(n460), .Z(n1233) );
  NAND U623 ( .A(n1258), .B(n1259), .Z(n461) );
  XOR U624 ( .A(n1258), .B(n1259), .Z(n462) );
  NANDN U625 ( .A(n1257), .B(n462), .Z(n463) );
  NAND U626 ( .A(n461), .B(n463), .Z(n1271) );
  NAND U627 ( .A(n1277), .B(n1278), .Z(n464) );
  XOR U628 ( .A(n1277), .B(n1278), .Z(n465) );
  NANDN U629 ( .A(n1276), .B(n465), .Z(n466) );
  NAND U630 ( .A(n464), .B(n466), .Z(n1290) );
  NAND U631 ( .A(n1296), .B(n1297), .Z(n467) );
  XOR U632 ( .A(n1296), .B(n1297), .Z(n468) );
  NANDN U633 ( .A(n1295), .B(n468), .Z(n469) );
  NAND U634 ( .A(n467), .B(n469), .Z(n1309) );
  NAND U635 ( .A(n1334), .B(n1335), .Z(n470) );
  XOR U636 ( .A(n1334), .B(n1335), .Z(n471) );
  NANDN U637 ( .A(n1333), .B(n471), .Z(n472) );
  NAND U638 ( .A(n470), .B(n472), .Z(n1347) );
  NAND U639 ( .A(n1353), .B(n1354), .Z(n473) );
  XOR U640 ( .A(n1353), .B(n1354), .Z(n474) );
  NANDN U641 ( .A(n1352), .B(n474), .Z(n475) );
  NAND U642 ( .A(n473), .B(n475), .Z(n1366) );
  NAND U643 ( .A(n1372), .B(n1373), .Z(n476) );
  XOR U644 ( .A(n1372), .B(n1373), .Z(n477) );
  NANDN U645 ( .A(n1371), .B(n477), .Z(n478) );
  NAND U646 ( .A(n476), .B(n478), .Z(n1385) );
  NAND U647 ( .A(n1410), .B(n1411), .Z(n479) );
  XOR U648 ( .A(n1410), .B(n1411), .Z(n480) );
  NANDN U649 ( .A(n1409), .B(n480), .Z(n481) );
  NAND U650 ( .A(n479), .B(n481), .Z(n1423) );
  NAND U651 ( .A(n1429), .B(n1430), .Z(n482) );
  XOR U652 ( .A(n1429), .B(n1430), .Z(n483) );
  NANDN U653 ( .A(n1428), .B(n483), .Z(n484) );
  NAND U654 ( .A(n482), .B(n484), .Z(n1442) );
  NAND U655 ( .A(n1448), .B(n1449), .Z(n485) );
  XOR U656 ( .A(n1448), .B(n1449), .Z(n486) );
  NANDN U657 ( .A(n1447), .B(n486), .Z(n487) );
  NAND U658 ( .A(n485), .B(n487), .Z(n1461) );
  NAND U659 ( .A(n1486), .B(n1487), .Z(n488) );
  XOR U660 ( .A(n1486), .B(n1487), .Z(n489) );
  NANDN U661 ( .A(n1485), .B(n489), .Z(n490) );
  NAND U662 ( .A(n488), .B(n490), .Z(n1499) );
  NAND U663 ( .A(n1505), .B(n1506), .Z(n491) );
  XOR U664 ( .A(n1505), .B(n1506), .Z(n492) );
  NANDN U665 ( .A(n1504), .B(n492), .Z(n493) );
  NAND U666 ( .A(n491), .B(n493), .Z(n1518) );
  NAND U667 ( .A(n1524), .B(n1525), .Z(n494) );
  XOR U668 ( .A(n1524), .B(n1525), .Z(n495) );
  NANDN U669 ( .A(n1523), .B(n495), .Z(n496) );
  NAND U670 ( .A(n494), .B(n496), .Z(n1537) );
  NAND U671 ( .A(n1562), .B(n1563), .Z(n497) );
  XOR U672 ( .A(n1562), .B(n1563), .Z(n498) );
  NANDN U673 ( .A(n1561), .B(n498), .Z(n499) );
  NAND U674 ( .A(n497), .B(n499), .Z(n1575) );
  NAND U675 ( .A(n1581), .B(n1582), .Z(n500) );
  XOR U676 ( .A(n1581), .B(n1582), .Z(n501) );
  NANDN U677 ( .A(n1580), .B(n501), .Z(n502) );
  NAND U678 ( .A(n500), .B(n502), .Z(n1594) );
  NAND U679 ( .A(n1600), .B(n1601), .Z(n503) );
  XOR U680 ( .A(n1600), .B(n1601), .Z(n504) );
  NANDN U681 ( .A(n1599), .B(n504), .Z(n505) );
  NAND U682 ( .A(n503), .B(n505), .Z(n1613) );
  NAND U683 ( .A(n1638), .B(n1639), .Z(n506) );
  XOR U684 ( .A(n1638), .B(n1639), .Z(n507) );
  NANDN U685 ( .A(n1637), .B(n507), .Z(n508) );
  NAND U686 ( .A(n506), .B(n508), .Z(n1651) );
  NAND U687 ( .A(n1657), .B(n1658), .Z(n509) );
  XOR U688 ( .A(n1657), .B(n1658), .Z(n510) );
  NANDN U689 ( .A(n1656), .B(n510), .Z(n511) );
  NAND U690 ( .A(n509), .B(n511), .Z(n1670) );
  NAND U691 ( .A(n1676), .B(n1677), .Z(n512) );
  XOR U692 ( .A(n1676), .B(n1677), .Z(n513) );
  NANDN U693 ( .A(n1675), .B(n513), .Z(n514) );
  NAND U694 ( .A(n512), .B(n514), .Z(n1689) );
  NAND U695 ( .A(n1714), .B(n1715), .Z(n515) );
  XOR U696 ( .A(n1714), .B(n1715), .Z(n516) );
  NANDN U697 ( .A(n1713), .B(n516), .Z(n517) );
  NAND U698 ( .A(n515), .B(n517), .Z(n1727) );
  NAND U699 ( .A(n654), .B(n653), .Z(n518) );
  XOR U700 ( .A(n654), .B(n653), .Z(n519) );
  NANDN U701 ( .A(sreg[66]), .B(n519), .Z(n520) );
  NAND U702 ( .A(n518), .B(n520), .Z(n673) );
  NAND U703 ( .A(n730), .B(n729), .Z(n521) );
  XOR U704 ( .A(n730), .B(n729), .Z(n522) );
  NANDN U705 ( .A(sreg[70]), .B(n522), .Z(n523) );
  NAND U706 ( .A(n521), .B(n523), .Z(n749) );
  NAND U707 ( .A(n806), .B(n805), .Z(n524) );
  XOR U708 ( .A(n806), .B(n805), .Z(n525) );
  NANDN U709 ( .A(sreg[74]), .B(n525), .Z(n526) );
  NAND U710 ( .A(n524), .B(n526), .Z(n825) );
  NAND U711 ( .A(n882), .B(n881), .Z(n527) );
  XOR U712 ( .A(n882), .B(n881), .Z(n528) );
  NANDN U713 ( .A(sreg[78]), .B(n528), .Z(n529) );
  NAND U714 ( .A(n527), .B(n529), .Z(n901) );
  NAND U715 ( .A(n958), .B(n957), .Z(n530) );
  XOR U716 ( .A(n958), .B(n957), .Z(n531) );
  NANDN U717 ( .A(sreg[82]), .B(n531), .Z(n532) );
  NAND U718 ( .A(n530), .B(n532), .Z(n977) );
  NAND U719 ( .A(n1034), .B(n1033), .Z(n533) );
  XOR U720 ( .A(n1034), .B(n1033), .Z(n534) );
  NANDN U721 ( .A(sreg[86]), .B(n534), .Z(n535) );
  NAND U722 ( .A(n533), .B(n535), .Z(n1053) );
  NAND U723 ( .A(n1110), .B(n1109), .Z(n536) );
  XOR U724 ( .A(n1110), .B(n1109), .Z(n537) );
  NANDN U725 ( .A(sreg[90]), .B(n537), .Z(n538) );
  NAND U726 ( .A(n536), .B(n538), .Z(n1129) );
  NAND U727 ( .A(n1186), .B(n1185), .Z(n539) );
  XOR U728 ( .A(n1186), .B(n1185), .Z(n540) );
  NANDN U729 ( .A(sreg[94]), .B(n540), .Z(n541) );
  NAND U730 ( .A(n539), .B(n541), .Z(n1205) );
  NAND U731 ( .A(n1262), .B(n1261), .Z(n542) );
  XOR U732 ( .A(n1262), .B(n1261), .Z(n543) );
  NANDN U733 ( .A(sreg[98]), .B(n543), .Z(n544) );
  NAND U734 ( .A(n542), .B(n544), .Z(n1281) );
  NAND U735 ( .A(n1338), .B(n1337), .Z(n545) );
  XOR U736 ( .A(n1338), .B(n1337), .Z(n546) );
  NANDN U737 ( .A(sreg[102]), .B(n546), .Z(n547) );
  NAND U738 ( .A(n545), .B(n547), .Z(n1357) );
  NAND U739 ( .A(n1414), .B(n1413), .Z(n548) );
  XOR U740 ( .A(n1414), .B(n1413), .Z(n549) );
  NANDN U741 ( .A(sreg[106]), .B(n549), .Z(n550) );
  NAND U742 ( .A(n548), .B(n550), .Z(n1433) );
  NAND U743 ( .A(n1490), .B(n1489), .Z(n551) );
  XOR U744 ( .A(n1490), .B(n1489), .Z(n552) );
  NANDN U745 ( .A(sreg[110]), .B(n552), .Z(n553) );
  NAND U746 ( .A(n551), .B(n553), .Z(n1509) );
  NAND U747 ( .A(n1566), .B(n1565), .Z(n554) );
  XOR U748 ( .A(n1566), .B(n1565), .Z(n555) );
  NANDN U749 ( .A(sreg[114]), .B(n555), .Z(n556) );
  NAND U750 ( .A(n554), .B(n556), .Z(n1585) );
  NAND U751 ( .A(n1642), .B(n1641), .Z(n557) );
  XOR U752 ( .A(n1642), .B(n1641), .Z(n558) );
  NANDN U753 ( .A(sreg[118]), .B(n558), .Z(n559) );
  NAND U754 ( .A(n557), .B(n559), .Z(n1661) );
  NAND U755 ( .A(n1718), .B(n1717), .Z(n560) );
  XOR U756 ( .A(n1718), .B(n1717), .Z(n561) );
  NANDN U757 ( .A(sreg[122]), .B(n561), .Z(n562) );
  NAND U758 ( .A(n560), .B(n562), .Z(n1721) );
  NANDN U759 ( .A(n1750), .B(n1751), .Z(n563) );
  XNOR U760 ( .A(n1750), .B(n1751), .Z(n564) );
  NAND U761 ( .A(n1752), .B(n564), .Z(n565) );
  AND U762 ( .A(n563), .B(n565), .Z(n566) );
  XNOR U763 ( .A(n1761), .B(n566), .Z(n1758) );
  AND U764 ( .A(a[0]), .B(b[0]), .Z(n567) );
  XOR U765 ( .A(n567), .B(sreg[60]), .Z(c[60]) );
  NAND U766 ( .A(b[1]), .B(a[0]), .Z(n601) );
  AND U767 ( .A(b[0]), .B(a[1]), .Z(n569) );
  XOR U768 ( .A(n601), .B(n569), .Z(n573) );
  NAND U769 ( .A(n567), .B(sreg[60]), .Z(n572) );
  IV U770 ( .A(n572), .Z(n571) );
  XOR U771 ( .A(sreg[61]), .B(n571), .Z(n568) );
  XNOR U772 ( .A(n573), .B(n568), .Z(c[61]) );
  NAND U773 ( .A(a[0]), .B(b[2]), .Z(n583) );
  ANDN U774 ( .B(n569), .A(n601), .Z(n585) );
  AND U775 ( .A(b[0]), .B(a[2]), .Z(n579) );
  AND U776 ( .A(b[1]), .B(a[1]), .Z(n578) );
  XOR U777 ( .A(n579), .B(n578), .Z(n584) );
  XNOR U778 ( .A(n585), .B(n584), .Z(n570) );
  XOR U779 ( .A(n583), .B(n570), .Z(n589) );
  IV U780 ( .A(n589), .Z(n587) );
  OR U781 ( .A(sreg[61]), .B(n571), .Z(n576) );
  ANDN U782 ( .B(sreg[61]), .A(n572), .Z(n574) );
  NANDN U783 ( .A(n574), .B(n573), .Z(n575) );
  AND U784 ( .A(n576), .B(n575), .Z(n588) );
  XOR U785 ( .A(n587), .B(n588), .Z(n577) );
  XNOR U786 ( .A(sreg[62]), .B(n577), .Z(c[62]) );
  AND U787 ( .A(a[1]), .B(b[2]), .Z(n595) );
  AND U788 ( .A(b[0]), .B(a[3]), .Z(n594) );
  XOR U789 ( .A(n595), .B(n594), .Z(n599) );
  AND U790 ( .A(a[2]), .B(b[1]), .Z(n581) );
  AND U791 ( .A(a[0]), .B(b[3]), .Z(n580) );
  XNOR U792 ( .A(n581), .B(n580), .Z(n582) );
  XOR U793 ( .A(n602), .B(n582), .Z(n598) );
  XNOR U794 ( .A(n598), .B(n600), .Z(n586) );
  XOR U795 ( .A(n599), .B(n586), .Z(n604) );
  NANDN U796 ( .A(n587), .B(n588), .Z(n592) );
  NOR U797 ( .A(n589), .B(n588), .Z(n590) );
  NANDN U798 ( .A(n590), .B(sreg[62]), .Z(n591) );
  AND U799 ( .A(n592), .B(n591), .Z(n605) );
  XNOR U800 ( .A(n605), .B(sreg[63]), .Z(n593) );
  XOR U801 ( .A(n604), .B(n593), .Z(c[63]) );
  NAND U802 ( .A(a[2]), .B(b[2]), .Z(n608) );
  NAND U803 ( .A(b[3]), .B(a[1]), .Z(n607) );
  XOR U804 ( .A(n609), .B(n607), .Z(n596) );
  XOR U805 ( .A(n608), .B(n596), .Z(n616) );
  AND U806 ( .A(b[1]), .B(a[3]), .Z(n617) );
  NAND U807 ( .A(b[0]), .B(a[4]), .Z(n615) );
  XOR U808 ( .A(n617), .B(n615), .Z(n597) );
  XNOR U809 ( .A(n616), .B(n597), .Z(n614) );
  AND U810 ( .A(b[3]), .B(a[2]), .Z(n624) );
  XNOR U811 ( .A(n613), .B(n612), .Z(n603) );
  XOR U812 ( .A(n614), .B(n603), .Z(n619) );
  XNOR U813 ( .A(n620), .B(sreg[64]), .Z(n606) );
  XOR U814 ( .A(n619), .B(n606), .Z(c[64]) );
  NAND U815 ( .A(b[0]), .B(a[5]), .Z(n630) );
  NAND U816 ( .A(b[2]), .B(a[3]), .Z(n623) );
  AND U817 ( .A(b[1]), .B(a[4]), .Z(n625) );
  XNOR U818 ( .A(n624), .B(n625), .Z(n610) );
  XOR U819 ( .A(n623), .B(n610), .Z(n631) );
  XNOR U820 ( .A(n632), .B(n631), .Z(n611) );
  XOR U821 ( .A(n630), .B(n611), .Z(n627) );
  XNOR U822 ( .A(n629), .B(n628), .Z(n618) );
  XOR U823 ( .A(n627), .B(n618), .Z(n634) );
  XNOR U824 ( .A(n635), .B(sreg[65]), .Z(n621) );
  XNOR U825 ( .A(n634), .B(n621), .Z(c[65]) );
  NAND U826 ( .A(b[2]), .B(a[4]), .Z(n639) );
  AND U827 ( .A(b[1]), .B(a[5]), .Z(n640) );
  NAND U828 ( .A(b[3]), .B(a[3]), .Z(n638) );
  XOR U829 ( .A(n640), .B(n638), .Z(n622) );
  XOR U830 ( .A(n639), .B(n622), .Z(n650) );
  NAND U831 ( .A(b[0]), .B(a[6]), .Z(n649) );
  XOR U832 ( .A(n651), .B(n649), .Z(n626) );
  XOR U833 ( .A(n650), .B(n626), .Z(n643) );
  IV U834 ( .A(n643), .Z(n642) );
  XNOR U835 ( .A(n646), .B(n644), .Z(n633) );
  XOR U836 ( .A(n642), .B(n633), .Z(n653) );
  XNOR U837 ( .A(n654), .B(sreg[66]), .Z(n636) );
  XNOR U838 ( .A(n653), .B(n636), .Z(c[66]) );
  NAND U839 ( .A(b[2]), .B(a[5]), .Z(n658) );
  AND U840 ( .A(b[1]), .B(a[6]), .Z(n659) );
  NAND U841 ( .A(b[3]), .B(a[4]), .Z(n657) );
  XOR U842 ( .A(n659), .B(n657), .Z(n637) );
  XOR U843 ( .A(n658), .B(n637), .Z(n669) );
  NAND U844 ( .A(b[0]), .B(a[7]), .Z(n668) );
  XOR U845 ( .A(n670), .B(n668), .Z(n641) );
  XOR U846 ( .A(n669), .B(n641), .Z(n662) );
  IV U847 ( .A(n662), .Z(n661) );
  OR U848 ( .A(n644), .B(n642), .Z(n648) );
  ANDN U849 ( .B(n644), .A(n643), .Z(n645) );
  OR U850 ( .A(n646), .B(n645), .Z(n647) );
  AND U851 ( .A(n648), .B(n647), .Z(n665) );
  XNOR U852 ( .A(n665), .B(n663), .Z(n652) );
  XOR U853 ( .A(n661), .B(n652), .Z(n672) );
  XNOR U854 ( .A(n673), .B(sreg[67]), .Z(n655) );
  XNOR U855 ( .A(n672), .B(n655), .Z(c[67]) );
  NAND U856 ( .A(b[2]), .B(a[6]), .Z(n677) );
  AND U857 ( .A(b[1]), .B(a[7]), .Z(n678) );
  NAND U858 ( .A(b[3]), .B(a[5]), .Z(n676) );
  XOR U859 ( .A(n678), .B(n676), .Z(n656) );
  XOR U860 ( .A(n677), .B(n656), .Z(n688) );
  NAND U861 ( .A(b[0]), .B(a[8]), .Z(n687) );
  XOR U862 ( .A(n689), .B(n687), .Z(n660) );
  XOR U863 ( .A(n688), .B(n660), .Z(n681) );
  IV U864 ( .A(n681), .Z(n680) );
  OR U865 ( .A(n663), .B(n661), .Z(n667) );
  ANDN U866 ( .B(n663), .A(n662), .Z(n664) );
  OR U867 ( .A(n665), .B(n664), .Z(n666) );
  AND U868 ( .A(n667), .B(n666), .Z(n684) );
  XNOR U869 ( .A(n684), .B(n682), .Z(n671) );
  XOR U870 ( .A(n680), .B(n671), .Z(n691) );
  XNOR U871 ( .A(n692), .B(sreg[68]), .Z(n674) );
  XNOR U872 ( .A(n691), .B(n674), .Z(c[68]) );
  NAND U873 ( .A(b[2]), .B(a[7]), .Z(n696) );
  AND U874 ( .A(b[1]), .B(a[8]), .Z(n697) );
  NAND U875 ( .A(b[3]), .B(a[6]), .Z(n695) );
  XOR U876 ( .A(n697), .B(n695), .Z(n675) );
  XOR U877 ( .A(n696), .B(n675), .Z(n707) );
  NAND U878 ( .A(b[0]), .B(a[9]), .Z(n706) );
  XOR U879 ( .A(n708), .B(n706), .Z(n679) );
  XOR U880 ( .A(n707), .B(n679), .Z(n700) );
  IV U881 ( .A(n700), .Z(n699) );
  OR U882 ( .A(n682), .B(n680), .Z(n686) );
  ANDN U883 ( .B(n682), .A(n681), .Z(n683) );
  OR U884 ( .A(n684), .B(n683), .Z(n685) );
  AND U885 ( .A(n686), .B(n685), .Z(n703) );
  XNOR U886 ( .A(n703), .B(n701), .Z(n690) );
  XOR U887 ( .A(n699), .B(n690), .Z(n710) );
  XNOR U888 ( .A(n711), .B(sreg[69]), .Z(n693) );
  XNOR U889 ( .A(n710), .B(n693), .Z(c[69]) );
  NAND U890 ( .A(b[2]), .B(a[8]), .Z(n715) );
  AND U891 ( .A(b[1]), .B(a[9]), .Z(n716) );
  NAND U892 ( .A(b[3]), .B(a[7]), .Z(n714) );
  XOR U893 ( .A(n716), .B(n714), .Z(n694) );
  XOR U894 ( .A(n715), .B(n694), .Z(n726) );
  NAND U895 ( .A(b[0]), .B(a[10]), .Z(n725) );
  XOR U896 ( .A(n727), .B(n725), .Z(n698) );
  XOR U897 ( .A(n726), .B(n698), .Z(n719) );
  IV U898 ( .A(n719), .Z(n718) );
  OR U899 ( .A(n701), .B(n699), .Z(n705) );
  ANDN U900 ( .B(n701), .A(n700), .Z(n702) );
  OR U901 ( .A(n703), .B(n702), .Z(n704) );
  AND U902 ( .A(n705), .B(n704), .Z(n722) );
  XNOR U903 ( .A(n722), .B(n720), .Z(n709) );
  XOR U904 ( .A(n718), .B(n709), .Z(n729) );
  XNOR U905 ( .A(n730), .B(sreg[70]), .Z(n712) );
  XNOR U906 ( .A(n729), .B(n712), .Z(c[70]) );
  NAND U907 ( .A(b[2]), .B(a[9]), .Z(n734) );
  AND U908 ( .A(b[1]), .B(a[10]), .Z(n735) );
  NAND U909 ( .A(b[3]), .B(a[8]), .Z(n733) );
  XOR U910 ( .A(n735), .B(n733), .Z(n713) );
  XOR U911 ( .A(n734), .B(n713), .Z(n745) );
  NAND U912 ( .A(b[0]), .B(a[11]), .Z(n744) );
  XOR U913 ( .A(n746), .B(n744), .Z(n717) );
  XOR U914 ( .A(n745), .B(n717), .Z(n738) );
  IV U915 ( .A(n738), .Z(n737) );
  OR U916 ( .A(n720), .B(n718), .Z(n724) );
  ANDN U917 ( .B(n720), .A(n719), .Z(n721) );
  OR U918 ( .A(n722), .B(n721), .Z(n723) );
  AND U919 ( .A(n724), .B(n723), .Z(n741) );
  XNOR U920 ( .A(n741), .B(n739), .Z(n728) );
  XOR U921 ( .A(n737), .B(n728), .Z(n748) );
  XNOR U922 ( .A(n749), .B(sreg[71]), .Z(n731) );
  XNOR U923 ( .A(n748), .B(n731), .Z(c[71]) );
  NAND U924 ( .A(b[2]), .B(a[10]), .Z(n753) );
  AND U925 ( .A(b[1]), .B(a[11]), .Z(n754) );
  NAND U926 ( .A(b[3]), .B(a[9]), .Z(n752) );
  XOR U927 ( .A(n754), .B(n752), .Z(n732) );
  XOR U928 ( .A(n753), .B(n732), .Z(n764) );
  NAND U929 ( .A(b[0]), .B(a[12]), .Z(n763) );
  XOR U930 ( .A(n765), .B(n763), .Z(n736) );
  XOR U931 ( .A(n764), .B(n736), .Z(n757) );
  IV U932 ( .A(n757), .Z(n756) );
  OR U933 ( .A(n739), .B(n737), .Z(n743) );
  ANDN U934 ( .B(n739), .A(n738), .Z(n740) );
  OR U935 ( .A(n741), .B(n740), .Z(n742) );
  AND U936 ( .A(n743), .B(n742), .Z(n760) );
  XNOR U937 ( .A(n760), .B(n758), .Z(n747) );
  XOR U938 ( .A(n756), .B(n747), .Z(n767) );
  XNOR U939 ( .A(n768), .B(sreg[72]), .Z(n750) );
  XNOR U940 ( .A(n767), .B(n750), .Z(c[72]) );
  NAND U941 ( .A(b[2]), .B(a[11]), .Z(n772) );
  AND U942 ( .A(b[1]), .B(a[12]), .Z(n773) );
  NAND U943 ( .A(b[3]), .B(a[10]), .Z(n771) );
  XOR U944 ( .A(n773), .B(n771), .Z(n751) );
  XOR U945 ( .A(n772), .B(n751), .Z(n783) );
  NAND U946 ( .A(b[0]), .B(a[13]), .Z(n782) );
  XOR U947 ( .A(n784), .B(n782), .Z(n755) );
  XOR U948 ( .A(n783), .B(n755), .Z(n776) );
  IV U949 ( .A(n776), .Z(n775) );
  OR U950 ( .A(n758), .B(n756), .Z(n762) );
  ANDN U951 ( .B(n758), .A(n757), .Z(n759) );
  OR U952 ( .A(n760), .B(n759), .Z(n761) );
  AND U953 ( .A(n762), .B(n761), .Z(n779) );
  XNOR U954 ( .A(n779), .B(n777), .Z(n766) );
  XOR U955 ( .A(n775), .B(n766), .Z(n786) );
  XNOR U956 ( .A(n787), .B(sreg[73]), .Z(n769) );
  XNOR U957 ( .A(n786), .B(n769), .Z(c[73]) );
  NAND U958 ( .A(b[2]), .B(a[12]), .Z(n791) );
  AND U959 ( .A(b[1]), .B(a[13]), .Z(n792) );
  NAND U960 ( .A(b[3]), .B(a[11]), .Z(n790) );
  XOR U961 ( .A(n792), .B(n790), .Z(n770) );
  XOR U962 ( .A(n791), .B(n770), .Z(n802) );
  NAND U963 ( .A(b[0]), .B(a[14]), .Z(n801) );
  XOR U964 ( .A(n803), .B(n801), .Z(n774) );
  XOR U965 ( .A(n802), .B(n774), .Z(n795) );
  IV U966 ( .A(n795), .Z(n794) );
  OR U967 ( .A(n777), .B(n775), .Z(n781) );
  ANDN U968 ( .B(n777), .A(n776), .Z(n778) );
  OR U969 ( .A(n779), .B(n778), .Z(n780) );
  AND U970 ( .A(n781), .B(n780), .Z(n798) );
  XNOR U971 ( .A(n798), .B(n796), .Z(n785) );
  XOR U972 ( .A(n794), .B(n785), .Z(n805) );
  XNOR U973 ( .A(n806), .B(sreg[74]), .Z(n788) );
  XNOR U974 ( .A(n805), .B(n788), .Z(c[74]) );
  NAND U975 ( .A(b[2]), .B(a[13]), .Z(n810) );
  AND U976 ( .A(b[1]), .B(a[14]), .Z(n811) );
  NAND U977 ( .A(b[3]), .B(a[12]), .Z(n809) );
  XOR U978 ( .A(n811), .B(n809), .Z(n789) );
  XOR U979 ( .A(n810), .B(n789), .Z(n821) );
  NAND U980 ( .A(b[0]), .B(a[15]), .Z(n820) );
  XOR U981 ( .A(n822), .B(n820), .Z(n793) );
  XOR U982 ( .A(n821), .B(n793), .Z(n814) );
  IV U983 ( .A(n814), .Z(n813) );
  OR U984 ( .A(n796), .B(n794), .Z(n800) );
  ANDN U985 ( .B(n796), .A(n795), .Z(n797) );
  OR U986 ( .A(n798), .B(n797), .Z(n799) );
  AND U987 ( .A(n800), .B(n799), .Z(n817) );
  XNOR U988 ( .A(n817), .B(n815), .Z(n804) );
  XOR U989 ( .A(n813), .B(n804), .Z(n824) );
  XNOR U990 ( .A(n825), .B(sreg[75]), .Z(n807) );
  XNOR U991 ( .A(n824), .B(n807), .Z(c[75]) );
  NAND U992 ( .A(b[2]), .B(a[14]), .Z(n829) );
  AND U993 ( .A(b[1]), .B(a[15]), .Z(n830) );
  NAND U994 ( .A(b[3]), .B(a[13]), .Z(n828) );
  XOR U995 ( .A(n830), .B(n828), .Z(n808) );
  XOR U996 ( .A(n829), .B(n808), .Z(n840) );
  NAND U997 ( .A(b[0]), .B(a[16]), .Z(n839) );
  XOR U998 ( .A(n841), .B(n839), .Z(n812) );
  XOR U999 ( .A(n840), .B(n812), .Z(n833) );
  IV U1000 ( .A(n833), .Z(n832) );
  OR U1001 ( .A(n815), .B(n813), .Z(n819) );
  ANDN U1002 ( .B(n815), .A(n814), .Z(n816) );
  OR U1003 ( .A(n817), .B(n816), .Z(n818) );
  AND U1004 ( .A(n819), .B(n818), .Z(n836) );
  XNOR U1005 ( .A(n836), .B(n834), .Z(n823) );
  XOR U1006 ( .A(n832), .B(n823), .Z(n843) );
  XNOR U1007 ( .A(n844), .B(sreg[76]), .Z(n826) );
  XNOR U1008 ( .A(n843), .B(n826), .Z(c[76]) );
  NAND U1009 ( .A(b[2]), .B(a[15]), .Z(n848) );
  AND U1010 ( .A(b[1]), .B(a[16]), .Z(n849) );
  NAND U1011 ( .A(b[3]), .B(a[14]), .Z(n847) );
  XOR U1012 ( .A(n849), .B(n847), .Z(n827) );
  XOR U1013 ( .A(n848), .B(n827), .Z(n859) );
  NAND U1014 ( .A(b[0]), .B(a[17]), .Z(n858) );
  XOR U1015 ( .A(n860), .B(n858), .Z(n831) );
  XOR U1016 ( .A(n859), .B(n831), .Z(n852) );
  IV U1017 ( .A(n852), .Z(n851) );
  OR U1018 ( .A(n834), .B(n832), .Z(n838) );
  ANDN U1019 ( .B(n834), .A(n833), .Z(n835) );
  OR U1020 ( .A(n836), .B(n835), .Z(n837) );
  AND U1021 ( .A(n838), .B(n837), .Z(n855) );
  XNOR U1022 ( .A(n855), .B(n853), .Z(n842) );
  XOR U1023 ( .A(n851), .B(n842), .Z(n862) );
  XNOR U1024 ( .A(n863), .B(sreg[77]), .Z(n845) );
  XNOR U1025 ( .A(n862), .B(n845), .Z(c[77]) );
  NAND U1026 ( .A(b[2]), .B(a[16]), .Z(n867) );
  AND U1027 ( .A(b[1]), .B(a[17]), .Z(n868) );
  NAND U1028 ( .A(b[3]), .B(a[15]), .Z(n866) );
  XOR U1029 ( .A(n868), .B(n866), .Z(n846) );
  XOR U1030 ( .A(n867), .B(n846), .Z(n878) );
  NAND U1031 ( .A(b[0]), .B(a[18]), .Z(n877) );
  XOR U1032 ( .A(n879), .B(n877), .Z(n850) );
  XOR U1033 ( .A(n878), .B(n850), .Z(n871) );
  IV U1034 ( .A(n871), .Z(n870) );
  OR U1035 ( .A(n853), .B(n851), .Z(n857) );
  ANDN U1036 ( .B(n853), .A(n852), .Z(n854) );
  OR U1037 ( .A(n855), .B(n854), .Z(n856) );
  AND U1038 ( .A(n857), .B(n856), .Z(n874) );
  XNOR U1039 ( .A(n874), .B(n872), .Z(n861) );
  XOR U1040 ( .A(n870), .B(n861), .Z(n881) );
  XNOR U1041 ( .A(n882), .B(sreg[78]), .Z(n864) );
  XNOR U1042 ( .A(n881), .B(n864), .Z(c[78]) );
  NAND U1043 ( .A(b[2]), .B(a[17]), .Z(n886) );
  AND U1044 ( .A(b[1]), .B(a[18]), .Z(n887) );
  NAND U1045 ( .A(b[3]), .B(a[16]), .Z(n885) );
  XOR U1046 ( .A(n887), .B(n885), .Z(n865) );
  XOR U1047 ( .A(n886), .B(n865), .Z(n897) );
  NAND U1048 ( .A(b[0]), .B(a[19]), .Z(n896) );
  XOR U1049 ( .A(n898), .B(n896), .Z(n869) );
  XOR U1050 ( .A(n897), .B(n869), .Z(n890) );
  IV U1051 ( .A(n890), .Z(n889) );
  OR U1052 ( .A(n872), .B(n870), .Z(n876) );
  ANDN U1053 ( .B(n872), .A(n871), .Z(n873) );
  OR U1054 ( .A(n874), .B(n873), .Z(n875) );
  AND U1055 ( .A(n876), .B(n875), .Z(n893) );
  XNOR U1056 ( .A(n893), .B(n891), .Z(n880) );
  XOR U1057 ( .A(n889), .B(n880), .Z(n900) );
  XNOR U1058 ( .A(n901), .B(sreg[79]), .Z(n883) );
  XNOR U1059 ( .A(n900), .B(n883), .Z(c[79]) );
  NAND U1060 ( .A(b[2]), .B(a[18]), .Z(n905) );
  AND U1061 ( .A(b[1]), .B(a[19]), .Z(n906) );
  NAND U1062 ( .A(b[3]), .B(a[17]), .Z(n904) );
  XOR U1063 ( .A(n906), .B(n904), .Z(n884) );
  XOR U1064 ( .A(n905), .B(n884), .Z(n916) );
  NAND U1065 ( .A(b[0]), .B(a[20]), .Z(n915) );
  XOR U1066 ( .A(n917), .B(n915), .Z(n888) );
  XOR U1067 ( .A(n916), .B(n888), .Z(n909) );
  IV U1068 ( .A(n909), .Z(n908) );
  OR U1069 ( .A(n891), .B(n889), .Z(n895) );
  ANDN U1070 ( .B(n891), .A(n890), .Z(n892) );
  OR U1071 ( .A(n893), .B(n892), .Z(n894) );
  AND U1072 ( .A(n895), .B(n894), .Z(n912) );
  XNOR U1073 ( .A(n912), .B(n910), .Z(n899) );
  XOR U1074 ( .A(n908), .B(n899), .Z(n919) );
  XNOR U1075 ( .A(n920), .B(sreg[80]), .Z(n902) );
  XNOR U1076 ( .A(n919), .B(n902), .Z(c[80]) );
  NAND U1077 ( .A(b[2]), .B(a[19]), .Z(n924) );
  AND U1078 ( .A(b[1]), .B(a[20]), .Z(n925) );
  NAND U1079 ( .A(b[3]), .B(a[18]), .Z(n923) );
  XOR U1080 ( .A(n925), .B(n923), .Z(n903) );
  XOR U1081 ( .A(n924), .B(n903), .Z(n935) );
  NAND U1082 ( .A(b[0]), .B(a[21]), .Z(n934) );
  XOR U1083 ( .A(n936), .B(n934), .Z(n907) );
  XOR U1084 ( .A(n935), .B(n907), .Z(n928) );
  IV U1085 ( .A(n928), .Z(n927) );
  OR U1086 ( .A(n910), .B(n908), .Z(n914) );
  ANDN U1087 ( .B(n910), .A(n909), .Z(n911) );
  OR U1088 ( .A(n912), .B(n911), .Z(n913) );
  AND U1089 ( .A(n914), .B(n913), .Z(n931) );
  XNOR U1090 ( .A(n931), .B(n929), .Z(n918) );
  XOR U1091 ( .A(n927), .B(n918), .Z(n938) );
  XNOR U1092 ( .A(n939), .B(sreg[81]), .Z(n921) );
  XNOR U1093 ( .A(n938), .B(n921), .Z(c[81]) );
  NAND U1094 ( .A(b[2]), .B(a[20]), .Z(n943) );
  AND U1095 ( .A(b[1]), .B(a[21]), .Z(n944) );
  NAND U1096 ( .A(b[3]), .B(a[19]), .Z(n942) );
  XOR U1097 ( .A(n944), .B(n942), .Z(n922) );
  XOR U1098 ( .A(n943), .B(n922), .Z(n954) );
  NAND U1099 ( .A(b[0]), .B(a[22]), .Z(n953) );
  XOR U1100 ( .A(n955), .B(n953), .Z(n926) );
  XOR U1101 ( .A(n954), .B(n926), .Z(n947) );
  IV U1102 ( .A(n947), .Z(n946) );
  OR U1103 ( .A(n929), .B(n927), .Z(n933) );
  ANDN U1104 ( .B(n929), .A(n928), .Z(n930) );
  OR U1105 ( .A(n931), .B(n930), .Z(n932) );
  AND U1106 ( .A(n933), .B(n932), .Z(n950) );
  XNOR U1107 ( .A(n950), .B(n948), .Z(n937) );
  XOR U1108 ( .A(n946), .B(n937), .Z(n957) );
  XNOR U1109 ( .A(n958), .B(sreg[82]), .Z(n940) );
  XNOR U1110 ( .A(n957), .B(n940), .Z(c[82]) );
  NAND U1111 ( .A(b[2]), .B(a[21]), .Z(n962) );
  AND U1112 ( .A(b[1]), .B(a[22]), .Z(n963) );
  NAND U1113 ( .A(b[3]), .B(a[20]), .Z(n961) );
  XOR U1114 ( .A(n963), .B(n961), .Z(n941) );
  XOR U1115 ( .A(n962), .B(n941), .Z(n973) );
  NAND U1116 ( .A(b[0]), .B(a[23]), .Z(n972) );
  XOR U1117 ( .A(n974), .B(n972), .Z(n945) );
  XOR U1118 ( .A(n973), .B(n945), .Z(n966) );
  IV U1119 ( .A(n966), .Z(n965) );
  OR U1120 ( .A(n948), .B(n946), .Z(n952) );
  ANDN U1121 ( .B(n948), .A(n947), .Z(n949) );
  OR U1122 ( .A(n950), .B(n949), .Z(n951) );
  AND U1123 ( .A(n952), .B(n951), .Z(n969) );
  XNOR U1124 ( .A(n969), .B(n967), .Z(n956) );
  XOR U1125 ( .A(n965), .B(n956), .Z(n976) );
  XNOR U1126 ( .A(n977), .B(sreg[83]), .Z(n959) );
  XNOR U1127 ( .A(n976), .B(n959), .Z(c[83]) );
  NAND U1128 ( .A(b[2]), .B(a[22]), .Z(n981) );
  AND U1129 ( .A(b[1]), .B(a[23]), .Z(n982) );
  NAND U1130 ( .A(b[3]), .B(a[21]), .Z(n980) );
  XOR U1131 ( .A(n982), .B(n980), .Z(n960) );
  XOR U1132 ( .A(n981), .B(n960), .Z(n992) );
  NAND U1133 ( .A(b[0]), .B(a[24]), .Z(n991) );
  XOR U1134 ( .A(n993), .B(n991), .Z(n964) );
  XOR U1135 ( .A(n992), .B(n964), .Z(n985) );
  IV U1136 ( .A(n985), .Z(n984) );
  OR U1137 ( .A(n967), .B(n965), .Z(n971) );
  ANDN U1138 ( .B(n967), .A(n966), .Z(n968) );
  OR U1139 ( .A(n969), .B(n968), .Z(n970) );
  AND U1140 ( .A(n971), .B(n970), .Z(n988) );
  XNOR U1141 ( .A(n988), .B(n986), .Z(n975) );
  XOR U1142 ( .A(n984), .B(n975), .Z(n995) );
  XNOR U1143 ( .A(n996), .B(sreg[84]), .Z(n978) );
  XNOR U1144 ( .A(n995), .B(n978), .Z(c[84]) );
  NAND U1145 ( .A(b[2]), .B(a[23]), .Z(n1000) );
  AND U1146 ( .A(b[1]), .B(a[24]), .Z(n1001) );
  NAND U1147 ( .A(b[3]), .B(a[22]), .Z(n999) );
  XOR U1148 ( .A(n1001), .B(n999), .Z(n979) );
  XOR U1149 ( .A(n1000), .B(n979), .Z(n1011) );
  NAND U1150 ( .A(b[0]), .B(a[25]), .Z(n1010) );
  XOR U1151 ( .A(n1012), .B(n1010), .Z(n983) );
  XOR U1152 ( .A(n1011), .B(n983), .Z(n1004) );
  IV U1153 ( .A(n1004), .Z(n1003) );
  OR U1154 ( .A(n986), .B(n984), .Z(n990) );
  ANDN U1155 ( .B(n986), .A(n985), .Z(n987) );
  OR U1156 ( .A(n988), .B(n987), .Z(n989) );
  AND U1157 ( .A(n990), .B(n989), .Z(n1007) );
  XNOR U1158 ( .A(n1007), .B(n1005), .Z(n994) );
  XOR U1159 ( .A(n1003), .B(n994), .Z(n1014) );
  XNOR U1160 ( .A(n1015), .B(sreg[85]), .Z(n997) );
  XNOR U1161 ( .A(n1014), .B(n997), .Z(c[85]) );
  NAND U1162 ( .A(b[2]), .B(a[24]), .Z(n1019) );
  AND U1163 ( .A(b[1]), .B(a[25]), .Z(n1020) );
  NAND U1164 ( .A(b[3]), .B(a[23]), .Z(n1018) );
  XOR U1165 ( .A(n1020), .B(n1018), .Z(n998) );
  XOR U1166 ( .A(n1019), .B(n998), .Z(n1030) );
  NAND U1167 ( .A(b[0]), .B(a[26]), .Z(n1029) );
  XOR U1168 ( .A(n1031), .B(n1029), .Z(n1002) );
  XOR U1169 ( .A(n1030), .B(n1002), .Z(n1023) );
  IV U1170 ( .A(n1023), .Z(n1022) );
  OR U1171 ( .A(n1005), .B(n1003), .Z(n1009) );
  ANDN U1172 ( .B(n1005), .A(n1004), .Z(n1006) );
  OR U1173 ( .A(n1007), .B(n1006), .Z(n1008) );
  AND U1174 ( .A(n1009), .B(n1008), .Z(n1026) );
  XNOR U1175 ( .A(n1026), .B(n1024), .Z(n1013) );
  XOR U1176 ( .A(n1022), .B(n1013), .Z(n1033) );
  XNOR U1177 ( .A(n1034), .B(sreg[86]), .Z(n1016) );
  XNOR U1178 ( .A(n1033), .B(n1016), .Z(c[86]) );
  NAND U1179 ( .A(b[2]), .B(a[25]), .Z(n1038) );
  AND U1180 ( .A(b[1]), .B(a[26]), .Z(n1039) );
  NAND U1181 ( .A(b[3]), .B(a[24]), .Z(n1037) );
  XOR U1182 ( .A(n1039), .B(n1037), .Z(n1017) );
  XOR U1183 ( .A(n1038), .B(n1017), .Z(n1049) );
  NAND U1184 ( .A(b[0]), .B(a[27]), .Z(n1048) );
  XOR U1185 ( .A(n1050), .B(n1048), .Z(n1021) );
  XOR U1186 ( .A(n1049), .B(n1021), .Z(n1042) );
  IV U1187 ( .A(n1042), .Z(n1041) );
  OR U1188 ( .A(n1024), .B(n1022), .Z(n1028) );
  ANDN U1189 ( .B(n1024), .A(n1023), .Z(n1025) );
  OR U1190 ( .A(n1026), .B(n1025), .Z(n1027) );
  AND U1191 ( .A(n1028), .B(n1027), .Z(n1045) );
  XNOR U1192 ( .A(n1045), .B(n1043), .Z(n1032) );
  XOR U1193 ( .A(n1041), .B(n1032), .Z(n1052) );
  XNOR U1194 ( .A(n1053), .B(sreg[87]), .Z(n1035) );
  XNOR U1195 ( .A(n1052), .B(n1035), .Z(c[87]) );
  NAND U1196 ( .A(b[2]), .B(a[26]), .Z(n1057) );
  AND U1197 ( .A(b[1]), .B(a[27]), .Z(n1058) );
  NAND U1198 ( .A(b[3]), .B(a[25]), .Z(n1056) );
  XOR U1199 ( .A(n1058), .B(n1056), .Z(n1036) );
  XOR U1200 ( .A(n1057), .B(n1036), .Z(n1068) );
  NAND U1201 ( .A(b[0]), .B(a[28]), .Z(n1067) );
  XOR U1202 ( .A(n1069), .B(n1067), .Z(n1040) );
  XOR U1203 ( .A(n1068), .B(n1040), .Z(n1061) );
  IV U1204 ( .A(n1061), .Z(n1060) );
  OR U1205 ( .A(n1043), .B(n1041), .Z(n1047) );
  ANDN U1206 ( .B(n1043), .A(n1042), .Z(n1044) );
  OR U1207 ( .A(n1045), .B(n1044), .Z(n1046) );
  AND U1208 ( .A(n1047), .B(n1046), .Z(n1064) );
  XNOR U1209 ( .A(n1064), .B(n1062), .Z(n1051) );
  XOR U1210 ( .A(n1060), .B(n1051), .Z(n1071) );
  XNOR U1211 ( .A(n1072), .B(sreg[88]), .Z(n1054) );
  XNOR U1212 ( .A(n1071), .B(n1054), .Z(c[88]) );
  NAND U1213 ( .A(b[2]), .B(a[27]), .Z(n1076) );
  AND U1214 ( .A(b[1]), .B(a[28]), .Z(n1077) );
  NAND U1215 ( .A(b[3]), .B(a[26]), .Z(n1075) );
  XOR U1216 ( .A(n1077), .B(n1075), .Z(n1055) );
  XOR U1217 ( .A(n1076), .B(n1055), .Z(n1087) );
  NAND U1218 ( .A(b[0]), .B(a[29]), .Z(n1086) );
  XOR U1219 ( .A(n1088), .B(n1086), .Z(n1059) );
  XOR U1220 ( .A(n1087), .B(n1059), .Z(n1080) );
  IV U1221 ( .A(n1080), .Z(n1079) );
  OR U1222 ( .A(n1062), .B(n1060), .Z(n1066) );
  ANDN U1223 ( .B(n1062), .A(n1061), .Z(n1063) );
  OR U1224 ( .A(n1064), .B(n1063), .Z(n1065) );
  AND U1225 ( .A(n1066), .B(n1065), .Z(n1083) );
  XNOR U1226 ( .A(n1083), .B(n1081), .Z(n1070) );
  XOR U1227 ( .A(n1079), .B(n1070), .Z(n1090) );
  XNOR U1228 ( .A(n1091), .B(sreg[89]), .Z(n1073) );
  XNOR U1229 ( .A(n1090), .B(n1073), .Z(c[89]) );
  NAND U1230 ( .A(b[2]), .B(a[28]), .Z(n1095) );
  AND U1231 ( .A(b[1]), .B(a[29]), .Z(n1096) );
  NAND U1232 ( .A(b[3]), .B(a[27]), .Z(n1094) );
  XOR U1233 ( .A(n1096), .B(n1094), .Z(n1074) );
  XOR U1234 ( .A(n1095), .B(n1074), .Z(n1106) );
  NAND U1235 ( .A(b[0]), .B(a[30]), .Z(n1105) );
  XOR U1236 ( .A(n1107), .B(n1105), .Z(n1078) );
  XOR U1237 ( .A(n1106), .B(n1078), .Z(n1099) );
  IV U1238 ( .A(n1099), .Z(n1098) );
  OR U1239 ( .A(n1081), .B(n1079), .Z(n1085) );
  ANDN U1240 ( .B(n1081), .A(n1080), .Z(n1082) );
  OR U1241 ( .A(n1083), .B(n1082), .Z(n1084) );
  AND U1242 ( .A(n1085), .B(n1084), .Z(n1102) );
  XNOR U1243 ( .A(n1102), .B(n1100), .Z(n1089) );
  XOR U1244 ( .A(n1098), .B(n1089), .Z(n1109) );
  XNOR U1245 ( .A(n1110), .B(sreg[90]), .Z(n1092) );
  XNOR U1246 ( .A(n1109), .B(n1092), .Z(c[90]) );
  NAND U1247 ( .A(b[2]), .B(a[29]), .Z(n1114) );
  AND U1248 ( .A(b[1]), .B(a[30]), .Z(n1115) );
  NAND U1249 ( .A(b[3]), .B(a[28]), .Z(n1113) );
  XOR U1250 ( .A(n1115), .B(n1113), .Z(n1093) );
  XOR U1251 ( .A(n1114), .B(n1093), .Z(n1125) );
  NAND U1252 ( .A(b[0]), .B(a[31]), .Z(n1124) );
  XOR U1253 ( .A(n1126), .B(n1124), .Z(n1097) );
  XOR U1254 ( .A(n1125), .B(n1097), .Z(n1118) );
  IV U1255 ( .A(n1118), .Z(n1117) );
  OR U1256 ( .A(n1100), .B(n1098), .Z(n1104) );
  ANDN U1257 ( .B(n1100), .A(n1099), .Z(n1101) );
  OR U1258 ( .A(n1102), .B(n1101), .Z(n1103) );
  AND U1259 ( .A(n1104), .B(n1103), .Z(n1121) );
  XNOR U1260 ( .A(n1121), .B(n1119), .Z(n1108) );
  XOR U1261 ( .A(n1117), .B(n1108), .Z(n1128) );
  XNOR U1262 ( .A(n1129), .B(sreg[91]), .Z(n1111) );
  XNOR U1263 ( .A(n1128), .B(n1111), .Z(c[91]) );
  NAND U1264 ( .A(b[2]), .B(a[30]), .Z(n1133) );
  AND U1265 ( .A(b[1]), .B(a[31]), .Z(n1134) );
  NAND U1266 ( .A(b[3]), .B(a[29]), .Z(n1132) );
  XOR U1267 ( .A(n1134), .B(n1132), .Z(n1112) );
  XOR U1268 ( .A(n1133), .B(n1112), .Z(n1144) );
  NAND U1269 ( .A(b[0]), .B(a[32]), .Z(n1143) );
  XOR U1270 ( .A(n1145), .B(n1143), .Z(n1116) );
  XOR U1271 ( .A(n1144), .B(n1116), .Z(n1137) );
  IV U1272 ( .A(n1137), .Z(n1136) );
  OR U1273 ( .A(n1119), .B(n1117), .Z(n1123) );
  ANDN U1274 ( .B(n1119), .A(n1118), .Z(n1120) );
  OR U1275 ( .A(n1121), .B(n1120), .Z(n1122) );
  AND U1276 ( .A(n1123), .B(n1122), .Z(n1140) );
  XNOR U1277 ( .A(n1140), .B(n1138), .Z(n1127) );
  XOR U1278 ( .A(n1136), .B(n1127), .Z(n1147) );
  XNOR U1279 ( .A(n1148), .B(sreg[92]), .Z(n1130) );
  XNOR U1280 ( .A(n1147), .B(n1130), .Z(c[92]) );
  NAND U1281 ( .A(b[2]), .B(a[31]), .Z(n1152) );
  AND U1282 ( .A(b[1]), .B(a[32]), .Z(n1153) );
  NAND U1283 ( .A(b[3]), .B(a[30]), .Z(n1151) );
  XOR U1284 ( .A(n1153), .B(n1151), .Z(n1131) );
  XOR U1285 ( .A(n1152), .B(n1131), .Z(n1163) );
  NAND U1286 ( .A(b[0]), .B(a[33]), .Z(n1162) );
  XOR U1287 ( .A(n1164), .B(n1162), .Z(n1135) );
  XOR U1288 ( .A(n1163), .B(n1135), .Z(n1156) );
  IV U1289 ( .A(n1156), .Z(n1155) );
  OR U1290 ( .A(n1138), .B(n1136), .Z(n1142) );
  ANDN U1291 ( .B(n1138), .A(n1137), .Z(n1139) );
  OR U1292 ( .A(n1140), .B(n1139), .Z(n1141) );
  AND U1293 ( .A(n1142), .B(n1141), .Z(n1159) );
  XNOR U1294 ( .A(n1159), .B(n1157), .Z(n1146) );
  XOR U1295 ( .A(n1155), .B(n1146), .Z(n1166) );
  XNOR U1296 ( .A(n1167), .B(sreg[93]), .Z(n1149) );
  XNOR U1297 ( .A(n1166), .B(n1149), .Z(c[93]) );
  NAND U1298 ( .A(b[2]), .B(a[32]), .Z(n1171) );
  AND U1299 ( .A(b[1]), .B(a[33]), .Z(n1172) );
  NAND U1300 ( .A(b[3]), .B(a[31]), .Z(n1170) );
  XOR U1301 ( .A(n1172), .B(n1170), .Z(n1150) );
  XOR U1302 ( .A(n1171), .B(n1150), .Z(n1182) );
  NAND U1303 ( .A(b[0]), .B(a[34]), .Z(n1181) );
  XOR U1304 ( .A(n1183), .B(n1181), .Z(n1154) );
  XOR U1305 ( .A(n1182), .B(n1154), .Z(n1175) );
  IV U1306 ( .A(n1175), .Z(n1174) );
  OR U1307 ( .A(n1157), .B(n1155), .Z(n1161) );
  ANDN U1308 ( .B(n1157), .A(n1156), .Z(n1158) );
  OR U1309 ( .A(n1159), .B(n1158), .Z(n1160) );
  AND U1310 ( .A(n1161), .B(n1160), .Z(n1178) );
  XNOR U1311 ( .A(n1178), .B(n1176), .Z(n1165) );
  XOR U1312 ( .A(n1174), .B(n1165), .Z(n1185) );
  XNOR U1313 ( .A(n1186), .B(sreg[94]), .Z(n1168) );
  XNOR U1314 ( .A(n1185), .B(n1168), .Z(c[94]) );
  NAND U1315 ( .A(b[2]), .B(a[33]), .Z(n1190) );
  AND U1316 ( .A(b[1]), .B(a[34]), .Z(n1191) );
  NAND U1317 ( .A(b[3]), .B(a[32]), .Z(n1189) );
  XOR U1318 ( .A(n1191), .B(n1189), .Z(n1169) );
  XOR U1319 ( .A(n1190), .B(n1169), .Z(n1201) );
  NAND U1320 ( .A(b[0]), .B(a[35]), .Z(n1200) );
  XOR U1321 ( .A(n1202), .B(n1200), .Z(n1173) );
  XOR U1322 ( .A(n1201), .B(n1173), .Z(n1194) );
  IV U1323 ( .A(n1194), .Z(n1193) );
  OR U1324 ( .A(n1176), .B(n1174), .Z(n1180) );
  ANDN U1325 ( .B(n1176), .A(n1175), .Z(n1177) );
  OR U1326 ( .A(n1178), .B(n1177), .Z(n1179) );
  AND U1327 ( .A(n1180), .B(n1179), .Z(n1197) );
  XNOR U1328 ( .A(n1197), .B(n1195), .Z(n1184) );
  XOR U1329 ( .A(n1193), .B(n1184), .Z(n1204) );
  XNOR U1330 ( .A(n1205), .B(sreg[95]), .Z(n1187) );
  XNOR U1331 ( .A(n1204), .B(n1187), .Z(c[95]) );
  NAND U1332 ( .A(b[2]), .B(a[34]), .Z(n1209) );
  AND U1333 ( .A(b[1]), .B(a[35]), .Z(n1210) );
  NAND U1334 ( .A(b[3]), .B(a[33]), .Z(n1208) );
  XOR U1335 ( .A(n1210), .B(n1208), .Z(n1188) );
  XOR U1336 ( .A(n1209), .B(n1188), .Z(n1220) );
  NAND U1337 ( .A(b[0]), .B(a[36]), .Z(n1219) );
  XOR U1338 ( .A(n1221), .B(n1219), .Z(n1192) );
  XOR U1339 ( .A(n1220), .B(n1192), .Z(n1213) );
  IV U1340 ( .A(n1213), .Z(n1212) );
  OR U1341 ( .A(n1195), .B(n1193), .Z(n1199) );
  ANDN U1342 ( .B(n1195), .A(n1194), .Z(n1196) );
  OR U1343 ( .A(n1197), .B(n1196), .Z(n1198) );
  AND U1344 ( .A(n1199), .B(n1198), .Z(n1216) );
  XNOR U1345 ( .A(n1216), .B(n1214), .Z(n1203) );
  XOR U1346 ( .A(n1212), .B(n1203), .Z(n1223) );
  XNOR U1347 ( .A(n1224), .B(sreg[96]), .Z(n1206) );
  XNOR U1348 ( .A(n1223), .B(n1206), .Z(c[96]) );
  NAND U1349 ( .A(b[2]), .B(a[35]), .Z(n1228) );
  AND U1350 ( .A(b[1]), .B(a[36]), .Z(n1229) );
  NAND U1351 ( .A(b[3]), .B(a[34]), .Z(n1227) );
  XOR U1352 ( .A(n1229), .B(n1227), .Z(n1207) );
  XOR U1353 ( .A(n1228), .B(n1207), .Z(n1239) );
  NAND U1354 ( .A(b[0]), .B(a[37]), .Z(n1238) );
  XOR U1355 ( .A(n1240), .B(n1238), .Z(n1211) );
  XOR U1356 ( .A(n1239), .B(n1211), .Z(n1232) );
  IV U1357 ( .A(n1232), .Z(n1231) );
  OR U1358 ( .A(n1214), .B(n1212), .Z(n1218) );
  ANDN U1359 ( .B(n1214), .A(n1213), .Z(n1215) );
  OR U1360 ( .A(n1216), .B(n1215), .Z(n1217) );
  AND U1361 ( .A(n1218), .B(n1217), .Z(n1235) );
  XNOR U1362 ( .A(n1235), .B(n1233), .Z(n1222) );
  XOR U1363 ( .A(n1231), .B(n1222), .Z(n1242) );
  XNOR U1364 ( .A(n1243), .B(sreg[97]), .Z(n1225) );
  XNOR U1365 ( .A(n1242), .B(n1225), .Z(c[97]) );
  NAND U1366 ( .A(b[2]), .B(a[36]), .Z(n1247) );
  AND U1367 ( .A(b[1]), .B(a[37]), .Z(n1248) );
  NAND U1368 ( .A(b[3]), .B(a[35]), .Z(n1246) );
  XOR U1369 ( .A(n1248), .B(n1246), .Z(n1226) );
  XOR U1370 ( .A(n1247), .B(n1226), .Z(n1258) );
  NAND U1371 ( .A(b[0]), .B(a[38]), .Z(n1257) );
  XOR U1372 ( .A(n1259), .B(n1257), .Z(n1230) );
  XOR U1373 ( .A(n1258), .B(n1230), .Z(n1251) );
  IV U1374 ( .A(n1251), .Z(n1250) );
  OR U1375 ( .A(n1233), .B(n1231), .Z(n1237) );
  ANDN U1376 ( .B(n1233), .A(n1232), .Z(n1234) );
  OR U1377 ( .A(n1235), .B(n1234), .Z(n1236) );
  AND U1378 ( .A(n1237), .B(n1236), .Z(n1254) );
  XNOR U1379 ( .A(n1254), .B(n1252), .Z(n1241) );
  XOR U1380 ( .A(n1250), .B(n1241), .Z(n1261) );
  XNOR U1381 ( .A(n1262), .B(sreg[98]), .Z(n1244) );
  XNOR U1382 ( .A(n1261), .B(n1244), .Z(c[98]) );
  NAND U1383 ( .A(b[2]), .B(a[37]), .Z(n1266) );
  AND U1384 ( .A(b[1]), .B(a[38]), .Z(n1267) );
  NAND U1385 ( .A(b[3]), .B(a[36]), .Z(n1265) );
  XOR U1386 ( .A(n1267), .B(n1265), .Z(n1245) );
  XOR U1387 ( .A(n1266), .B(n1245), .Z(n1277) );
  NAND U1388 ( .A(b[0]), .B(a[39]), .Z(n1276) );
  XOR U1389 ( .A(n1278), .B(n1276), .Z(n1249) );
  XOR U1390 ( .A(n1277), .B(n1249), .Z(n1270) );
  IV U1391 ( .A(n1270), .Z(n1269) );
  OR U1392 ( .A(n1252), .B(n1250), .Z(n1256) );
  ANDN U1393 ( .B(n1252), .A(n1251), .Z(n1253) );
  OR U1394 ( .A(n1254), .B(n1253), .Z(n1255) );
  AND U1395 ( .A(n1256), .B(n1255), .Z(n1273) );
  XNOR U1396 ( .A(n1273), .B(n1271), .Z(n1260) );
  XOR U1397 ( .A(n1269), .B(n1260), .Z(n1280) );
  XNOR U1398 ( .A(n1281), .B(sreg[99]), .Z(n1263) );
  XNOR U1399 ( .A(n1280), .B(n1263), .Z(c[99]) );
  NAND U1400 ( .A(b[2]), .B(a[38]), .Z(n1285) );
  AND U1401 ( .A(b[1]), .B(a[39]), .Z(n1286) );
  NAND U1402 ( .A(b[3]), .B(a[37]), .Z(n1284) );
  XOR U1403 ( .A(n1286), .B(n1284), .Z(n1264) );
  XOR U1404 ( .A(n1285), .B(n1264), .Z(n1296) );
  NAND U1405 ( .A(b[0]), .B(a[40]), .Z(n1295) );
  XOR U1406 ( .A(n1297), .B(n1295), .Z(n1268) );
  XOR U1407 ( .A(n1296), .B(n1268), .Z(n1289) );
  IV U1408 ( .A(n1289), .Z(n1288) );
  OR U1409 ( .A(n1271), .B(n1269), .Z(n1275) );
  ANDN U1410 ( .B(n1271), .A(n1270), .Z(n1272) );
  OR U1411 ( .A(n1273), .B(n1272), .Z(n1274) );
  AND U1412 ( .A(n1275), .B(n1274), .Z(n1292) );
  XNOR U1413 ( .A(n1292), .B(n1290), .Z(n1279) );
  XOR U1414 ( .A(n1288), .B(n1279), .Z(n1299) );
  XNOR U1415 ( .A(n1300), .B(sreg[100]), .Z(n1282) );
  XNOR U1416 ( .A(n1299), .B(n1282), .Z(c[100]) );
  NAND U1417 ( .A(b[2]), .B(a[39]), .Z(n1304) );
  AND U1418 ( .A(b[1]), .B(a[40]), .Z(n1305) );
  NAND U1419 ( .A(b[3]), .B(a[38]), .Z(n1303) );
  XOR U1420 ( .A(n1305), .B(n1303), .Z(n1283) );
  XOR U1421 ( .A(n1304), .B(n1283), .Z(n1315) );
  NAND U1422 ( .A(b[0]), .B(a[41]), .Z(n1314) );
  XOR U1423 ( .A(n1316), .B(n1314), .Z(n1287) );
  XOR U1424 ( .A(n1315), .B(n1287), .Z(n1308) );
  IV U1425 ( .A(n1308), .Z(n1307) );
  OR U1426 ( .A(n1290), .B(n1288), .Z(n1294) );
  ANDN U1427 ( .B(n1290), .A(n1289), .Z(n1291) );
  OR U1428 ( .A(n1292), .B(n1291), .Z(n1293) );
  AND U1429 ( .A(n1294), .B(n1293), .Z(n1311) );
  XNOR U1430 ( .A(n1311), .B(n1309), .Z(n1298) );
  XOR U1431 ( .A(n1307), .B(n1298), .Z(n1318) );
  XNOR U1432 ( .A(n1319), .B(sreg[101]), .Z(n1301) );
  XNOR U1433 ( .A(n1318), .B(n1301), .Z(c[101]) );
  NAND U1434 ( .A(b[2]), .B(a[40]), .Z(n1323) );
  AND U1435 ( .A(b[1]), .B(a[41]), .Z(n1324) );
  NAND U1436 ( .A(b[3]), .B(a[39]), .Z(n1322) );
  XOR U1437 ( .A(n1324), .B(n1322), .Z(n1302) );
  XOR U1438 ( .A(n1323), .B(n1302), .Z(n1334) );
  NAND U1439 ( .A(b[0]), .B(a[42]), .Z(n1333) );
  XOR U1440 ( .A(n1335), .B(n1333), .Z(n1306) );
  XOR U1441 ( .A(n1334), .B(n1306), .Z(n1327) );
  IV U1442 ( .A(n1327), .Z(n1326) );
  OR U1443 ( .A(n1309), .B(n1307), .Z(n1313) );
  ANDN U1444 ( .B(n1309), .A(n1308), .Z(n1310) );
  OR U1445 ( .A(n1311), .B(n1310), .Z(n1312) );
  AND U1446 ( .A(n1313), .B(n1312), .Z(n1330) );
  XNOR U1447 ( .A(n1330), .B(n1328), .Z(n1317) );
  XOR U1448 ( .A(n1326), .B(n1317), .Z(n1337) );
  XNOR U1449 ( .A(n1338), .B(sreg[102]), .Z(n1320) );
  XNOR U1450 ( .A(n1337), .B(n1320), .Z(c[102]) );
  NAND U1451 ( .A(b[2]), .B(a[41]), .Z(n1342) );
  AND U1452 ( .A(b[1]), .B(a[42]), .Z(n1343) );
  NAND U1453 ( .A(b[3]), .B(a[40]), .Z(n1341) );
  XOR U1454 ( .A(n1343), .B(n1341), .Z(n1321) );
  XOR U1455 ( .A(n1342), .B(n1321), .Z(n1353) );
  NAND U1456 ( .A(b[0]), .B(a[43]), .Z(n1352) );
  XOR U1457 ( .A(n1354), .B(n1352), .Z(n1325) );
  XOR U1458 ( .A(n1353), .B(n1325), .Z(n1346) );
  IV U1459 ( .A(n1346), .Z(n1345) );
  OR U1460 ( .A(n1328), .B(n1326), .Z(n1332) );
  ANDN U1461 ( .B(n1328), .A(n1327), .Z(n1329) );
  OR U1462 ( .A(n1330), .B(n1329), .Z(n1331) );
  AND U1463 ( .A(n1332), .B(n1331), .Z(n1349) );
  XNOR U1464 ( .A(n1349), .B(n1347), .Z(n1336) );
  XOR U1465 ( .A(n1345), .B(n1336), .Z(n1356) );
  XNOR U1466 ( .A(n1357), .B(sreg[103]), .Z(n1339) );
  XNOR U1467 ( .A(n1356), .B(n1339), .Z(c[103]) );
  NAND U1468 ( .A(b[2]), .B(a[42]), .Z(n1361) );
  AND U1469 ( .A(b[1]), .B(a[43]), .Z(n1362) );
  NAND U1470 ( .A(b[3]), .B(a[41]), .Z(n1360) );
  XOR U1471 ( .A(n1362), .B(n1360), .Z(n1340) );
  XOR U1472 ( .A(n1361), .B(n1340), .Z(n1372) );
  NAND U1473 ( .A(b[0]), .B(a[44]), .Z(n1371) );
  XOR U1474 ( .A(n1373), .B(n1371), .Z(n1344) );
  XOR U1475 ( .A(n1372), .B(n1344), .Z(n1365) );
  IV U1476 ( .A(n1365), .Z(n1364) );
  OR U1477 ( .A(n1347), .B(n1345), .Z(n1351) );
  ANDN U1478 ( .B(n1347), .A(n1346), .Z(n1348) );
  OR U1479 ( .A(n1349), .B(n1348), .Z(n1350) );
  AND U1480 ( .A(n1351), .B(n1350), .Z(n1368) );
  XNOR U1481 ( .A(n1368), .B(n1366), .Z(n1355) );
  XOR U1482 ( .A(n1364), .B(n1355), .Z(n1375) );
  XNOR U1483 ( .A(n1376), .B(sreg[104]), .Z(n1358) );
  XNOR U1484 ( .A(n1375), .B(n1358), .Z(c[104]) );
  NAND U1485 ( .A(b[2]), .B(a[43]), .Z(n1380) );
  AND U1486 ( .A(b[1]), .B(a[44]), .Z(n1381) );
  NAND U1487 ( .A(b[3]), .B(a[42]), .Z(n1379) );
  XOR U1488 ( .A(n1381), .B(n1379), .Z(n1359) );
  XOR U1489 ( .A(n1380), .B(n1359), .Z(n1391) );
  NAND U1490 ( .A(b[0]), .B(a[45]), .Z(n1390) );
  XOR U1491 ( .A(n1392), .B(n1390), .Z(n1363) );
  XOR U1492 ( .A(n1391), .B(n1363), .Z(n1384) );
  IV U1493 ( .A(n1384), .Z(n1383) );
  OR U1494 ( .A(n1366), .B(n1364), .Z(n1370) );
  ANDN U1495 ( .B(n1366), .A(n1365), .Z(n1367) );
  OR U1496 ( .A(n1368), .B(n1367), .Z(n1369) );
  AND U1497 ( .A(n1370), .B(n1369), .Z(n1387) );
  XNOR U1498 ( .A(n1387), .B(n1385), .Z(n1374) );
  XOR U1499 ( .A(n1383), .B(n1374), .Z(n1394) );
  XNOR U1500 ( .A(n1395), .B(sreg[105]), .Z(n1377) );
  XNOR U1501 ( .A(n1394), .B(n1377), .Z(c[105]) );
  NAND U1502 ( .A(b[2]), .B(a[44]), .Z(n1399) );
  AND U1503 ( .A(b[1]), .B(a[45]), .Z(n1400) );
  NAND U1504 ( .A(b[3]), .B(a[43]), .Z(n1398) );
  XOR U1505 ( .A(n1400), .B(n1398), .Z(n1378) );
  XOR U1506 ( .A(n1399), .B(n1378), .Z(n1410) );
  NAND U1507 ( .A(b[0]), .B(a[46]), .Z(n1409) );
  XOR U1508 ( .A(n1411), .B(n1409), .Z(n1382) );
  XOR U1509 ( .A(n1410), .B(n1382), .Z(n1403) );
  IV U1510 ( .A(n1403), .Z(n1402) );
  OR U1511 ( .A(n1385), .B(n1383), .Z(n1389) );
  ANDN U1512 ( .B(n1385), .A(n1384), .Z(n1386) );
  OR U1513 ( .A(n1387), .B(n1386), .Z(n1388) );
  AND U1514 ( .A(n1389), .B(n1388), .Z(n1406) );
  XNOR U1515 ( .A(n1406), .B(n1404), .Z(n1393) );
  XOR U1516 ( .A(n1402), .B(n1393), .Z(n1413) );
  XNOR U1517 ( .A(n1414), .B(sreg[106]), .Z(n1396) );
  XNOR U1518 ( .A(n1413), .B(n1396), .Z(c[106]) );
  NAND U1519 ( .A(b[2]), .B(a[45]), .Z(n1418) );
  AND U1520 ( .A(b[1]), .B(a[46]), .Z(n1419) );
  NAND U1521 ( .A(b[3]), .B(a[44]), .Z(n1417) );
  XOR U1522 ( .A(n1419), .B(n1417), .Z(n1397) );
  XOR U1523 ( .A(n1418), .B(n1397), .Z(n1429) );
  NAND U1524 ( .A(b[0]), .B(a[47]), .Z(n1428) );
  XOR U1525 ( .A(n1430), .B(n1428), .Z(n1401) );
  XOR U1526 ( .A(n1429), .B(n1401), .Z(n1422) );
  IV U1527 ( .A(n1422), .Z(n1421) );
  OR U1528 ( .A(n1404), .B(n1402), .Z(n1408) );
  ANDN U1529 ( .B(n1404), .A(n1403), .Z(n1405) );
  OR U1530 ( .A(n1406), .B(n1405), .Z(n1407) );
  AND U1531 ( .A(n1408), .B(n1407), .Z(n1425) );
  XNOR U1532 ( .A(n1425), .B(n1423), .Z(n1412) );
  XOR U1533 ( .A(n1421), .B(n1412), .Z(n1432) );
  XNOR U1534 ( .A(n1433), .B(sreg[107]), .Z(n1415) );
  XNOR U1535 ( .A(n1432), .B(n1415), .Z(c[107]) );
  NAND U1536 ( .A(b[2]), .B(a[46]), .Z(n1437) );
  AND U1537 ( .A(b[1]), .B(a[47]), .Z(n1438) );
  NAND U1538 ( .A(b[3]), .B(a[45]), .Z(n1436) );
  XOR U1539 ( .A(n1438), .B(n1436), .Z(n1416) );
  XOR U1540 ( .A(n1437), .B(n1416), .Z(n1448) );
  NAND U1541 ( .A(b[0]), .B(a[48]), .Z(n1447) );
  XOR U1542 ( .A(n1449), .B(n1447), .Z(n1420) );
  XOR U1543 ( .A(n1448), .B(n1420), .Z(n1441) );
  IV U1544 ( .A(n1441), .Z(n1440) );
  OR U1545 ( .A(n1423), .B(n1421), .Z(n1427) );
  ANDN U1546 ( .B(n1423), .A(n1422), .Z(n1424) );
  OR U1547 ( .A(n1425), .B(n1424), .Z(n1426) );
  AND U1548 ( .A(n1427), .B(n1426), .Z(n1444) );
  XNOR U1549 ( .A(n1444), .B(n1442), .Z(n1431) );
  XOR U1550 ( .A(n1440), .B(n1431), .Z(n1451) );
  XNOR U1551 ( .A(n1452), .B(sreg[108]), .Z(n1434) );
  XNOR U1552 ( .A(n1451), .B(n1434), .Z(c[108]) );
  NAND U1553 ( .A(b[2]), .B(a[47]), .Z(n1456) );
  AND U1554 ( .A(b[1]), .B(a[48]), .Z(n1457) );
  NAND U1555 ( .A(b[3]), .B(a[46]), .Z(n1455) );
  XOR U1556 ( .A(n1457), .B(n1455), .Z(n1435) );
  XOR U1557 ( .A(n1456), .B(n1435), .Z(n1467) );
  NAND U1558 ( .A(b[0]), .B(a[49]), .Z(n1466) );
  XOR U1559 ( .A(n1468), .B(n1466), .Z(n1439) );
  XOR U1560 ( .A(n1467), .B(n1439), .Z(n1460) );
  IV U1561 ( .A(n1460), .Z(n1459) );
  OR U1562 ( .A(n1442), .B(n1440), .Z(n1446) );
  ANDN U1563 ( .B(n1442), .A(n1441), .Z(n1443) );
  OR U1564 ( .A(n1444), .B(n1443), .Z(n1445) );
  AND U1565 ( .A(n1446), .B(n1445), .Z(n1463) );
  XNOR U1566 ( .A(n1463), .B(n1461), .Z(n1450) );
  XOR U1567 ( .A(n1459), .B(n1450), .Z(n1470) );
  XNOR U1568 ( .A(n1471), .B(sreg[109]), .Z(n1453) );
  XNOR U1569 ( .A(n1470), .B(n1453), .Z(c[109]) );
  NAND U1570 ( .A(b[2]), .B(a[48]), .Z(n1475) );
  AND U1571 ( .A(b[1]), .B(a[49]), .Z(n1476) );
  NAND U1572 ( .A(b[3]), .B(a[47]), .Z(n1474) );
  XOR U1573 ( .A(n1476), .B(n1474), .Z(n1454) );
  XOR U1574 ( .A(n1475), .B(n1454), .Z(n1486) );
  NAND U1575 ( .A(b[0]), .B(a[50]), .Z(n1485) );
  XOR U1576 ( .A(n1487), .B(n1485), .Z(n1458) );
  XOR U1577 ( .A(n1486), .B(n1458), .Z(n1479) );
  IV U1578 ( .A(n1479), .Z(n1478) );
  OR U1579 ( .A(n1461), .B(n1459), .Z(n1465) );
  ANDN U1580 ( .B(n1461), .A(n1460), .Z(n1462) );
  OR U1581 ( .A(n1463), .B(n1462), .Z(n1464) );
  AND U1582 ( .A(n1465), .B(n1464), .Z(n1482) );
  XNOR U1583 ( .A(n1482), .B(n1480), .Z(n1469) );
  XOR U1584 ( .A(n1478), .B(n1469), .Z(n1489) );
  XNOR U1585 ( .A(n1490), .B(sreg[110]), .Z(n1472) );
  XNOR U1586 ( .A(n1489), .B(n1472), .Z(c[110]) );
  NAND U1587 ( .A(b[2]), .B(a[49]), .Z(n1494) );
  AND U1588 ( .A(b[1]), .B(a[50]), .Z(n1495) );
  NAND U1589 ( .A(b[3]), .B(a[48]), .Z(n1493) );
  XOR U1590 ( .A(n1495), .B(n1493), .Z(n1473) );
  XOR U1591 ( .A(n1494), .B(n1473), .Z(n1505) );
  NAND U1592 ( .A(b[0]), .B(a[51]), .Z(n1504) );
  XOR U1593 ( .A(n1506), .B(n1504), .Z(n1477) );
  XOR U1594 ( .A(n1505), .B(n1477), .Z(n1498) );
  IV U1595 ( .A(n1498), .Z(n1497) );
  OR U1596 ( .A(n1480), .B(n1478), .Z(n1484) );
  ANDN U1597 ( .B(n1480), .A(n1479), .Z(n1481) );
  OR U1598 ( .A(n1482), .B(n1481), .Z(n1483) );
  AND U1599 ( .A(n1484), .B(n1483), .Z(n1501) );
  XNOR U1600 ( .A(n1501), .B(n1499), .Z(n1488) );
  XOR U1601 ( .A(n1497), .B(n1488), .Z(n1508) );
  XNOR U1602 ( .A(n1509), .B(sreg[111]), .Z(n1491) );
  XNOR U1603 ( .A(n1508), .B(n1491), .Z(c[111]) );
  NAND U1604 ( .A(b[2]), .B(a[50]), .Z(n1513) );
  AND U1605 ( .A(b[1]), .B(a[51]), .Z(n1514) );
  NAND U1606 ( .A(b[3]), .B(a[49]), .Z(n1512) );
  XOR U1607 ( .A(n1514), .B(n1512), .Z(n1492) );
  XOR U1608 ( .A(n1513), .B(n1492), .Z(n1524) );
  NAND U1609 ( .A(b[0]), .B(a[52]), .Z(n1523) );
  XOR U1610 ( .A(n1525), .B(n1523), .Z(n1496) );
  XOR U1611 ( .A(n1524), .B(n1496), .Z(n1517) );
  IV U1612 ( .A(n1517), .Z(n1516) );
  OR U1613 ( .A(n1499), .B(n1497), .Z(n1503) );
  ANDN U1614 ( .B(n1499), .A(n1498), .Z(n1500) );
  OR U1615 ( .A(n1501), .B(n1500), .Z(n1502) );
  AND U1616 ( .A(n1503), .B(n1502), .Z(n1520) );
  XNOR U1617 ( .A(n1520), .B(n1518), .Z(n1507) );
  XOR U1618 ( .A(n1516), .B(n1507), .Z(n1527) );
  XNOR U1619 ( .A(n1528), .B(sreg[112]), .Z(n1510) );
  XNOR U1620 ( .A(n1527), .B(n1510), .Z(c[112]) );
  NAND U1621 ( .A(b[2]), .B(a[51]), .Z(n1532) );
  AND U1622 ( .A(b[1]), .B(a[52]), .Z(n1533) );
  NAND U1623 ( .A(b[3]), .B(a[50]), .Z(n1531) );
  XOR U1624 ( .A(n1533), .B(n1531), .Z(n1511) );
  XOR U1625 ( .A(n1532), .B(n1511), .Z(n1543) );
  NAND U1626 ( .A(b[0]), .B(a[53]), .Z(n1542) );
  XOR U1627 ( .A(n1544), .B(n1542), .Z(n1515) );
  XOR U1628 ( .A(n1543), .B(n1515), .Z(n1536) );
  IV U1629 ( .A(n1536), .Z(n1535) );
  OR U1630 ( .A(n1518), .B(n1516), .Z(n1522) );
  ANDN U1631 ( .B(n1518), .A(n1517), .Z(n1519) );
  OR U1632 ( .A(n1520), .B(n1519), .Z(n1521) );
  AND U1633 ( .A(n1522), .B(n1521), .Z(n1539) );
  XNOR U1634 ( .A(n1539), .B(n1537), .Z(n1526) );
  XOR U1635 ( .A(n1535), .B(n1526), .Z(n1546) );
  XNOR U1636 ( .A(n1547), .B(sreg[113]), .Z(n1529) );
  XNOR U1637 ( .A(n1546), .B(n1529), .Z(c[113]) );
  NAND U1638 ( .A(b[2]), .B(a[52]), .Z(n1551) );
  AND U1639 ( .A(b[1]), .B(a[53]), .Z(n1552) );
  NAND U1640 ( .A(b[3]), .B(a[51]), .Z(n1550) );
  XOR U1641 ( .A(n1552), .B(n1550), .Z(n1530) );
  XOR U1642 ( .A(n1551), .B(n1530), .Z(n1562) );
  NAND U1643 ( .A(b[0]), .B(a[54]), .Z(n1561) );
  XOR U1644 ( .A(n1563), .B(n1561), .Z(n1534) );
  XOR U1645 ( .A(n1562), .B(n1534), .Z(n1555) );
  IV U1646 ( .A(n1555), .Z(n1554) );
  OR U1647 ( .A(n1537), .B(n1535), .Z(n1541) );
  ANDN U1648 ( .B(n1537), .A(n1536), .Z(n1538) );
  OR U1649 ( .A(n1539), .B(n1538), .Z(n1540) );
  AND U1650 ( .A(n1541), .B(n1540), .Z(n1558) );
  XNOR U1651 ( .A(n1558), .B(n1556), .Z(n1545) );
  XOR U1652 ( .A(n1554), .B(n1545), .Z(n1565) );
  XNOR U1653 ( .A(n1566), .B(sreg[114]), .Z(n1548) );
  XNOR U1654 ( .A(n1565), .B(n1548), .Z(c[114]) );
  NAND U1655 ( .A(b[2]), .B(a[53]), .Z(n1570) );
  AND U1656 ( .A(b[1]), .B(a[54]), .Z(n1571) );
  NAND U1657 ( .A(b[3]), .B(a[52]), .Z(n1569) );
  XOR U1658 ( .A(n1571), .B(n1569), .Z(n1549) );
  XOR U1659 ( .A(n1570), .B(n1549), .Z(n1581) );
  NAND U1660 ( .A(b[0]), .B(a[55]), .Z(n1580) );
  XOR U1661 ( .A(n1582), .B(n1580), .Z(n1553) );
  XOR U1662 ( .A(n1581), .B(n1553), .Z(n1574) );
  IV U1663 ( .A(n1574), .Z(n1573) );
  OR U1664 ( .A(n1556), .B(n1554), .Z(n1560) );
  ANDN U1665 ( .B(n1556), .A(n1555), .Z(n1557) );
  OR U1666 ( .A(n1558), .B(n1557), .Z(n1559) );
  AND U1667 ( .A(n1560), .B(n1559), .Z(n1577) );
  XNOR U1668 ( .A(n1577), .B(n1575), .Z(n1564) );
  XOR U1669 ( .A(n1573), .B(n1564), .Z(n1584) );
  XNOR U1670 ( .A(n1585), .B(sreg[115]), .Z(n1567) );
  XNOR U1671 ( .A(n1584), .B(n1567), .Z(c[115]) );
  NAND U1672 ( .A(b[2]), .B(a[54]), .Z(n1589) );
  AND U1673 ( .A(b[1]), .B(a[55]), .Z(n1590) );
  NAND U1674 ( .A(b[3]), .B(a[53]), .Z(n1588) );
  XOR U1675 ( .A(n1590), .B(n1588), .Z(n1568) );
  XOR U1676 ( .A(n1589), .B(n1568), .Z(n1600) );
  NAND U1677 ( .A(b[0]), .B(a[56]), .Z(n1599) );
  XOR U1678 ( .A(n1601), .B(n1599), .Z(n1572) );
  XOR U1679 ( .A(n1600), .B(n1572), .Z(n1593) );
  IV U1680 ( .A(n1593), .Z(n1592) );
  OR U1681 ( .A(n1575), .B(n1573), .Z(n1579) );
  ANDN U1682 ( .B(n1575), .A(n1574), .Z(n1576) );
  OR U1683 ( .A(n1577), .B(n1576), .Z(n1578) );
  AND U1684 ( .A(n1579), .B(n1578), .Z(n1596) );
  XNOR U1685 ( .A(n1596), .B(n1594), .Z(n1583) );
  XOR U1686 ( .A(n1592), .B(n1583), .Z(n1603) );
  XNOR U1687 ( .A(n1604), .B(sreg[116]), .Z(n1586) );
  XNOR U1688 ( .A(n1603), .B(n1586), .Z(c[116]) );
  NAND U1689 ( .A(b[2]), .B(a[55]), .Z(n1608) );
  AND U1690 ( .A(b[1]), .B(a[56]), .Z(n1609) );
  NAND U1691 ( .A(b[3]), .B(a[54]), .Z(n1607) );
  XOR U1692 ( .A(n1609), .B(n1607), .Z(n1587) );
  XOR U1693 ( .A(n1608), .B(n1587), .Z(n1619) );
  NAND U1694 ( .A(b[0]), .B(a[57]), .Z(n1618) );
  XOR U1695 ( .A(n1620), .B(n1618), .Z(n1591) );
  XOR U1696 ( .A(n1619), .B(n1591), .Z(n1612) );
  IV U1697 ( .A(n1612), .Z(n1611) );
  OR U1698 ( .A(n1594), .B(n1592), .Z(n1598) );
  ANDN U1699 ( .B(n1594), .A(n1593), .Z(n1595) );
  OR U1700 ( .A(n1596), .B(n1595), .Z(n1597) );
  AND U1701 ( .A(n1598), .B(n1597), .Z(n1615) );
  XNOR U1702 ( .A(n1615), .B(n1613), .Z(n1602) );
  XOR U1703 ( .A(n1611), .B(n1602), .Z(n1622) );
  XNOR U1704 ( .A(n1623), .B(sreg[117]), .Z(n1605) );
  XNOR U1705 ( .A(n1622), .B(n1605), .Z(c[117]) );
  NAND U1706 ( .A(b[2]), .B(a[56]), .Z(n1627) );
  AND U1707 ( .A(b[1]), .B(a[57]), .Z(n1628) );
  NAND U1708 ( .A(b[3]), .B(a[55]), .Z(n1626) );
  XOR U1709 ( .A(n1628), .B(n1626), .Z(n1606) );
  XOR U1710 ( .A(n1627), .B(n1606), .Z(n1638) );
  NAND U1711 ( .A(b[0]), .B(a[58]), .Z(n1637) );
  XOR U1712 ( .A(n1639), .B(n1637), .Z(n1610) );
  XOR U1713 ( .A(n1638), .B(n1610), .Z(n1631) );
  IV U1714 ( .A(n1631), .Z(n1630) );
  OR U1715 ( .A(n1613), .B(n1611), .Z(n1617) );
  ANDN U1716 ( .B(n1613), .A(n1612), .Z(n1614) );
  OR U1717 ( .A(n1615), .B(n1614), .Z(n1616) );
  AND U1718 ( .A(n1617), .B(n1616), .Z(n1634) );
  XNOR U1719 ( .A(n1634), .B(n1632), .Z(n1621) );
  XOR U1720 ( .A(n1630), .B(n1621), .Z(n1641) );
  XNOR U1721 ( .A(n1642), .B(sreg[118]), .Z(n1624) );
  XNOR U1722 ( .A(n1641), .B(n1624), .Z(c[118]) );
  NAND U1723 ( .A(b[2]), .B(a[57]), .Z(n1646) );
  AND U1724 ( .A(b[1]), .B(a[58]), .Z(n1647) );
  NAND U1725 ( .A(b[3]), .B(a[56]), .Z(n1645) );
  XOR U1726 ( .A(n1647), .B(n1645), .Z(n1625) );
  XOR U1727 ( .A(n1646), .B(n1625), .Z(n1657) );
  NAND U1728 ( .A(b[0]), .B(a[59]), .Z(n1656) );
  XOR U1729 ( .A(n1658), .B(n1656), .Z(n1629) );
  XOR U1730 ( .A(n1657), .B(n1629), .Z(n1650) );
  IV U1731 ( .A(n1650), .Z(n1649) );
  OR U1732 ( .A(n1632), .B(n1630), .Z(n1636) );
  ANDN U1733 ( .B(n1632), .A(n1631), .Z(n1633) );
  OR U1734 ( .A(n1634), .B(n1633), .Z(n1635) );
  AND U1735 ( .A(n1636), .B(n1635), .Z(n1653) );
  XNOR U1736 ( .A(n1653), .B(n1651), .Z(n1640) );
  XOR U1737 ( .A(n1649), .B(n1640), .Z(n1660) );
  XNOR U1738 ( .A(n1661), .B(sreg[119]), .Z(n1643) );
  XNOR U1739 ( .A(n1660), .B(n1643), .Z(c[119]) );
  NAND U1740 ( .A(b[2]), .B(a[58]), .Z(n1665) );
  AND U1741 ( .A(b[1]), .B(a[59]), .Z(n1666) );
  NAND U1742 ( .A(b[3]), .B(a[57]), .Z(n1664) );
  XOR U1743 ( .A(n1666), .B(n1664), .Z(n1644) );
  XOR U1744 ( .A(n1665), .B(n1644), .Z(n1676) );
  NAND U1745 ( .A(b[0]), .B(a[60]), .Z(n1675) );
  XOR U1746 ( .A(n1677), .B(n1675), .Z(n1648) );
  XOR U1747 ( .A(n1676), .B(n1648), .Z(n1669) );
  IV U1748 ( .A(n1669), .Z(n1668) );
  OR U1749 ( .A(n1651), .B(n1649), .Z(n1655) );
  ANDN U1750 ( .B(n1651), .A(n1650), .Z(n1652) );
  OR U1751 ( .A(n1653), .B(n1652), .Z(n1654) );
  AND U1752 ( .A(n1655), .B(n1654), .Z(n1672) );
  XNOR U1753 ( .A(n1672), .B(n1670), .Z(n1659) );
  XOR U1754 ( .A(n1668), .B(n1659), .Z(n1679) );
  XNOR U1755 ( .A(n1680), .B(sreg[120]), .Z(n1662) );
  XNOR U1756 ( .A(n1679), .B(n1662), .Z(c[120]) );
  NAND U1757 ( .A(b[2]), .B(a[59]), .Z(n1684) );
  AND U1758 ( .A(b[1]), .B(a[60]), .Z(n1685) );
  NAND U1759 ( .A(b[3]), .B(a[58]), .Z(n1683) );
  XOR U1760 ( .A(n1685), .B(n1683), .Z(n1663) );
  XOR U1761 ( .A(n1684), .B(n1663), .Z(n1695) );
  NAND U1762 ( .A(b[0]), .B(a[61]), .Z(n1694) );
  XOR U1763 ( .A(n1696), .B(n1694), .Z(n1667) );
  XOR U1764 ( .A(n1695), .B(n1667), .Z(n1688) );
  IV U1765 ( .A(n1688), .Z(n1687) );
  OR U1766 ( .A(n1670), .B(n1668), .Z(n1674) );
  ANDN U1767 ( .B(n1670), .A(n1669), .Z(n1671) );
  OR U1768 ( .A(n1672), .B(n1671), .Z(n1673) );
  AND U1769 ( .A(n1674), .B(n1673), .Z(n1691) );
  XNOR U1770 ( .A(n1691), .B(n1689), .Z(n1678) );
  XOR U1771 ( .A(n1687), .B(n1678), .Z(n1698) );
  XNOR U1772 ( .A(n1699), .B(sreg[121]), .Z(n1681) );
  XNOR U1773 ( .A(n1698), .B(n1681), .Z(c[121]) );
  NAND U1774 ( .A(b[2]), .B(a[60]), .Z(n1703) );
  AND U1775 ( .A(b[1]), .B(a[61]), .Z(n1704) );
  NAND U1776 ( .A(b[3]), .B(a[59]), .Z(n1702) );
  XOR U1777 ( .A(n1704), .B(n1702), .Z(n1682) );
  XOR U1778 ( .A(n1703), .B(n1682), .Z(n1714) );
  NAND U1779 ( .A(b[0]), .B(a[62]), .Z(n1713) );
  XOR U1780 ( .A(n1715), .B(n1713), .Z(n1686) );
  XOR U1781 ( .A(n1714), .B(n1686), .Z(n1707) );
  IV U1782 ( .A(n1707), .Z(n1706) );
  OR U1783 ( .A(n1689), .B(n1687), .Z(n1693) );
  ANDN U1784 ( .B(n1689), .A(n1688), .Z(n1690) );
  OR U1785 ( .A(n1691), .B(n1690), .Z(n1692) );
  AND U1786 ( .A(n1693), .B(n1692), .Z(n1710) );
  XNOR U1787 ( .A(n1710), .B(n1708), .Z(n1697) );
  XOR U1788 ( .A(n1706), .B(n1697), .Z(n1717) );
  XNOR U1789 ( .A(n1718), .B(sreg[122]), .Z(n1700) );
  XNOR U1790 ( .A(n1717), .B(n1700), .Z(c[122]) );
  NAND U1791 ( .A(b[2]), .B(a[61]), .Z(n1733) );
  AND U1792 ( .A(b[1]), .B(a[62]), .Z(n1734) );
  NAND U1793 ( .A(b[3]), .B(a[60]), .Z(n1732) );
  XOR U1794 ( .A(n1734), .B(n1732), .Z(n1701) );
  XOR U1795 ( .A(n1733), .B(n1701), .Z(n1723) );
  NAND U1796 ( .A(a[63]), .B(b[0]), .Z(n1722) );
  XOR U1797 ( .A(n1724), .B(n1722), .Z(n1705) );
  XOR U1798 ( .A(n1723), .B(n1705), .Z(n1726) );
  IV U1799 ( .A(n1726), .Z(n1725) );
  OR U1800 ( .A(n1708), .B(n1706), .Z(n1712) );
  ANDN U1801 ( .B(n1708), .A(n1707), .Z(n1709) );
  OR U1802 ( .A(n1710), .B(n1709), .Z(n1711) );
  AND U1803 ( .A(n1712), .B(n1711), .Z(n1729) );
  XNOR U1804 ( .A(n1729), .B(n1727), .Z(n1716) );
  XOR U1805 ( .A(n1725), .B(n1716), .Z(n1720) );
  XNOR U1806 ( .A(n1721), .B(sreg[123]), .Z(n1719) );
  XNOR U1807 ( .A(n1720), .B(n1719), .Z(c[123]) );
  OR U1808 ( .A(n1727), .B(n1725), .Z(n1731) );
  ANDN U1809 ( .B(n1727), .A(n1726), .Z(n1728) );
  OR U1810 ( .A(n1729), .B(n1728), .Z(n1730) );
  AND U1811 ( .A(n1731), .B(n1730), .Z(n1741) );
  AND U1812 ( .A(b[3]), .B(a[61]), .Z(n1747) );
  AND U1813 ( .A(b[2]), .B(a[62]), .Z(n1759) );
  AND U1814 ( .A(a[63]), .B(b[1]), .Z(n1753) );
  XNOR U1815 ( .A(n1759), .B(n1753), .Z(n1746) );
  XOR U1816 ( .A(n1747), .B(n1746), .Z(n1735) );
  XOR U1817 ( .A(n1748), .B(n1735), .Z(n1740) );
  XOR U1818 ( .A(n1741), .B(n1740), .Z(n1736) );
  XNOR U1819 ( .A(n1739), .B(n1736), .Z(n1738) );
  XNOR U1820 ( .A(n1737), .B(n1738), .Z(c[124]) );
  ANDN U1821 ( .B(n1738), .A(n1737), .Z(n1757) );
  AND U1822 ( .A(n1759), .B(n1753), .Z(n1745) );
  AND U1823 ( .A(b[2]), .B(a[63]), .Z(n1743) );
  NAND U1824 ( .A(a[62]), .B(b[3]), .Z(n1742) );
  XNOR U1825 ( .A(n1743), .B(n1742), .Z(n1744) );
  XOR U1826 ( .A(n1745), .B(n1744), .Z(n1751) );
  XOR U1827 ( .A(n1751), .B(n1750), .Z(n1749) );
  XNOR U1828 ( .A(n1752), .B(n1749), .Z(n1756) );
  XOR U1829 ( .A(n1757), .B(n1756), .Z(c[125]) );
  AND U1830 ( .A(b[3]), .B(a[63]), .Z(n1761) );
  OR U1831 ( .A(n1761), .B(n1753), .Z(n1754) );
  AND U1832 ( .A(n1759), .B(n1754), .Z(n1755) );
  XNOR U1833 ( .A(n1758), .B(n1755), .Z(n1763) );
  AND U1834 ( .A(n1757), .B(n1756), .Z(n1762) );
  XNOR U1835 ( .A(n1763), .B(n1762), .Z(c[126]) );
  NANDN U1836 ( .A(n1759), .B(n1758), .Z(n1760) );
  AND U1837 ( .A(n1761), .B(n1760), .Z(n1765) );
  NANDN U1838 ( .A(n1763), .B(n1762), .Z(n1764) );
  NANDN U1839 ( .A(n1765), .B(n1764), .Z(c[127]) );
endmodule

