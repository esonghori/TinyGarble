
module mult_N64_CC2 ( clk, rst, a, b, c );
  input [63:0] a;
  input [31:0] b;
  output [127:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926;
  wire   [127:0] sreg;

  DFF \sreg_reg[95]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(sreg[95]) );
  DFF \sreg_reg[94]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(sreg[94]) );
  DFF \sreg_reg[93]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(sreg[93]) );
  DFF \sreg_reg[92]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(sreg[92]) );
  DFF \sreg_reg[91]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(sreg[91]) );
  DFF \sreg_reg[90]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(sreg[90]) );
  DFF \sreg_reg[89]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(sreg[89]) );
  DFF \sreg_reg[88]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(sreg[88]) );
  DFF \sreg_reg[87]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(sreg[87]) );
  DFF \sreg_reg[86]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(sreg[86]) );
  DFF \sreg_reg[85]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(sreg[85]) );
  DFF \sreg_reg[84]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(sreg[84]) );
  DFF \sreg_reg[83]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(sreg[83]) );
  DFF \sreg_reg[82]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(sreg[82]) );
  DFF \sreg_reg[81]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(sreg[81]) );
  DFF \sreg_reg[80]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(sreg[80]) );
  DFF \sreg_reg[79]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(sreg[79]) );
  DFF \sreg_reg[78]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(sreg[78]) );
  DFF \sreg_reg[77]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(sreg[77]) );
  DFF \sreg_reg[76]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(sreg[76]) );
  DFF \sreg_reg[75]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(sreg[75]) );
  DFF \sreg_reg[74]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(sreg[74]) );
  DFF \sreg_reg[73]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(sreg[73]) );
  DFF \sreg_reg[72]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(sreg[72]) );
  DFF \sreg_reg[71]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(sreg[71]) );
  DFF \sreg_reg[70]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(sreg[70]) );
  DFF \sreg_reg[69]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(sreg[69]) );
  DFF \sreg_reg[68]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(sreg[68]) );
  DFF \sreg_reg[67]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(sreg[67]) );
  DFF \sreg_reg[66]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(sreg[66]) );
  DFF \sreg_reg[65]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(sreg[65]) );
  DFF \sreg_reg[64]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(sreg[64]) );
  DFF \sreg_reg[63]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(sreg[63]) );
  DFF \sreg_reg[62]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(sreg[62]) );
  DFF \sreg_reg[61]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(sreg[61]) );
  DFF \sreg_reg[60]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(sreg[60]) );
  DFF \sreg_reg[59]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(sreg[59]) );
  DFF \sreg_reg[58]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(sreg[58]) );
  DFF \sreg_reg[57]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(sreg[57]) );
  DFF \sreg_reg[56]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(sreg[56]) );
  DFF \sreg_reg[55]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(sreg[55]) );
  DFF \sreg_reg[54]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(sreg[54]) );
  DFF \sreg_reg[53]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(sreg[53]) );
  DFF \sreg_reg[52]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(sreg[52]) );
  DFF \sreg_reg[51]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(sreg[51]) );
  DFF \sreg_reg[50]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(sreg[50]) );
  DFF \sreg_reg[49]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(sreg[49]) );
  DFF \sreg_reg[48]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(sreg[48]) );
  DFF \sreg_reg[47]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(sreg[47]) );
  DFF \sreg_reg[46]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(sreg[46]) );
  DFF \sreg_reg[45]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(sreg[45]) );
  DFF \sreg_reg[44]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(sreg[44]) );
  DFF \sreg_reg[43]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(sreg[43]) );
  DFF \sreg_reg[42]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(sreg[42]) );
  DFF \sreg_reg[41]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(sreg[41]) );
  DFF \sreg_reg[40]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(sreg[40]) );
  DFF \sreg_reg[39]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(sreg[39]) );
  DFF \sreg_reg[38]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(sreg[38]) );
  DFF \sreg_reg[37]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(sreg[37]) );
  DFF \sreg_reg[36]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(sreg[36]) );
  DFF \sreg_reg[35]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(sreg[35]) );
  DFF \sreg_reg[34]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(sreg[34]) );
  DFF \sreg_reg[33]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(sreg[33]) );
  DFF \sreg_reg[32]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(sreg[32]) );
  DFF \sreg_reg[31]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[0]) );
  NANDN U35 ( .A(n7596), .B(n7597), .Z(n1) );
  NANDN U36 ( .A(n7594), .B(n7595), .Z(n2) );
  NAND U37 ( .A(n1), .B(n2), .Z(n7669) );
  XOR U38 ( .A(n7765), .B(n7764), .Z(n7766) );
  NANDN U39 ( .A(n7706), .B(n7707), .Z(n3) );
  NANDN U40 ( .A(n7708), .B(n7709), .Z(n4) );
  AND U41 ( .A(n3), .B(n4), .Z(n7802) );
  NANDN U42 ( .A(n7794), .B(n7795), .Z(n5) );
  NANDN U43 ( .A(n7797), .B(n7796), .Z(n6) );
  NAND U44 ( .A(n5), .B(n6), .Z(n7873) );
  NANDN U45 ( .A(n7843), .B(n7844), .Z(n7) );
  NANDN U46 ( .A(n7841), .B(n7842), .Z(n8) );
  NAND U47 ( .A(n7), .B(n8), .Z(n7870) );
  NANDN U48 ( .A(n8013), .B(n8014), .Z(n9) );
  NANDN U49 ( .A(n8011), .B(n8012), .Z(n10) );
  NAND U50 ( .A(n9), .B(n10), .Z(n8126) );
  NANDN U51 ( .A(n8015), .B(n8016), .Z(n11) );
  NANDN U52 ( .A(n8017), .B(n8018), .Z(n12) );
  AND U53 ( .A(n11), .B(n12), .Z(n8201) );
  NAND U54 ( .A(n8196), .B(n8195), .Z(n13) );
  NANDN U55 ( .A(n8193), .B(n8194), .Z(n14) );
  NAND U56 ( .A(n13), .B(n14), .Z(n8232) );
  NANDN U57 ( .A(n8418), .B(n8419), .Z(n15) );
  NANDN U58 ( .A(n8421), .B(n8420), .Z(n16) );
  NAND U59 ( .A(n15), .B(n16), .Z(n8511) );
  NANDN U60 ( .A(n8504), .B(n8505), .Z(n17) );
  NANDN U61 ( .A(n8502), .B(n8503), .Z(n18) );
  NAND U62 ( .A(n17), .B(n18), .Z(n8616) );
  NANDN U63 ( .A(n8237), .B(n8238), .Z(n19) );
  NANDN U64 ( .A(n8236), .B(n8235), .Z(n20) );
  AND U65 ( .A(n19), .B(n20), .Z(n8337) );
  NANDN U66 ( .A(n8446), .B(n8447), .Z(n21) );
  NANDN U67 ( .A(n8448), .B(n8449), .Z(n22) );
  AND U68 ( .A(n21), .B(n22), .Z(n8549) );
  NANDN U69 ( .A(n8736), .B(n8737), .Z(n23) );
  NANDN U70 ( .A(n8734), .B(n8735), .Z(n24) );
  NAND U71 ( .A(n23), .B(n24), .Z(n8754) );
  NANDN U72 ( .A(n8972), .B(n8973), .Z(n25) );
  NANDN U73 ( .A(n8970), .B(n8971), .Z(n26) );
  NAND U74 ( .A(n25), .B(n26), .Z(n9022) );
  NANDN U75 ( .A(n9347), .B(n9348), .Z(n27) );
  NANDN U76 ( .A(n9349), .B(n9350), .Z(n28) );
  AND U77 ( .A(n27), .B(n28), .Z(n9407) );
  NANDN U78 ( .A(n7507), .B(n7508), .Z(n29) );
  NANDN U79 ( .A(n7506), .B(n7505), .Z(n30) );
  NAND U80 ( .A(n29), .B(n30), .Z(n7621) );
  OR U81 ( .A(n7727), .B(n7726), .Z(n31) );
  NANDN U82 ( .A(n7728), .B(n7729), .Z(n32) );
  NAND U83 ( .A(n31), .B(n32), .Z(n7748) );
  NANDN U84 ( .A(n7762), .B(n7763), .Z(n33) );
  NANDN U85 ( .A(n7761), .B(n7760), .Z(n34) );
  AND U86 ( .A(n33), .B(n34), .Z(n7866) );
  NANDN U87 ( .A(n7986), .B(n7987), .Z(n35) );
  NANDN U88 ( .A(n7988), .B(n7989), .Z(n36) );
  AND U89 ( .A(n35), .B(n36), .Z(n8111) );
  NANDN U90 ( .A(n8669), .B(n8670), .Z(n37) );
  NANDN U91 ( .A(n8668), .B(n8667), .Z(n38) );
  AND U92 ( .A(n37), .B(n38), .Z(n8822) );
  NANDN U93 ( .A(n8891), .B(n8892), .Z(n39) );
  NANDN U94 ( .A(n8890), .B(n8889), .Z(n40) );
  AND U95 ( .A(n39), .B(n40), .Z(n8933) );
  NAND U96 ( .A(n8905), .B(n8904), .Z(n41) );
  NANDN U97 ( .A(n8906), .B(n8907), .Z(n42) );
  AND U98 ( .A(n41), .B(n42), .Z(n8929) );
  NANDN U99 ( .A(n9161), .B(n9162), .Z(n43) );
  NANDN U100 ( .A(n9159), .B(n9160), .Z(n44) );
  NAND U101 ( .A(n43), .B(n44), .Z(n9182) );
  NANDN U102 ( .A(n9310), .B(n9311), .Z(n45) );
  NANDN U103 ( .A(n9309), .B(n9308), .Z(n46) );
  NAND U104 ( .A(n45), .B(n46), .Z(n9331) );
  NANDN U105 ( .A(n9338), .B(n9339), .Z(n47) );
  NANDN U106 ( .A(n9340), .B(n9341), .Z(n48) );
  AND U107 ( .A(n47), .B(n48), .Z(n9401) );
  NANDN U108 ( .A(n9409), .B(n9410), .Z(n49) );
  NANDN U109 ( .A(n9411), .B(n9412), .Z(n50) );
  AND U110 ( .A(n49), .B(n50), .Z(n9502) );
  NANDN U111 ( .A(n9460), .B(n9461), .Z(n51) );
  NANDN U112 ( .A(n9462), .B(n9463), .Z(n52) );
  AND U113 ( .A(n51), .B(n52), .Z(n9558) );
  NAND U114 ( .A(n9523), .B(n9524), .Z(n53) );
  NANDN U115 ( .A(n9521), .B(n9522), .Z(n54) );
  AND U116 ( .A(n53), .B(n54), .Z(n9579) );
  NAND U117 ( .A(n9557), .B(n9556), .Z(n55) );
  NANDN U118 ( .A(n9554), .B(n9555), .Z(n56) );
  NAND U119 ( .A(n55), .B(n56), .Z(n9575) );
  XOR U120 ( .A(n7767), .B(n7766), .Z(n7805) );
  NANDN U121 ( .A(n7921), .B(n7922), .Z(n57) );
  NANDN U122 ( .A(n7919), .B(n7920), .Z(n58) );
  NAND U123 ( .A(n57), .B(n58), .Z(n8028) );
  NAND U124 ( .A(n8416), .B(n8417), .Z(n59) );
  NANDN U125 ( .A(n8414), .B(n8415), .Z(n60) );
  AND U126 ( .A(n59), .B(n60), .Z(n8510) );
  NANDN U127 ( .A(n8498), .B(n8499), .Z(n61) );
  NANDN U128 ( .A(n8500), .B(n8501), .Z(n62) );
  AND U129 ( .A(n61), .B(n62), .Z(n8615) );
  NANDN U130 ( .A(n7652), .B(n7653), .Z(n63) );
  NANDN U131 ( .A(n7654), .B(n7655), .Z(n64) );
  AND U132 ( .A(n63), .B(n64), .Z(n7850) );
  NANDN U133 ( .A(n7925), .B(n7926), .Z(n65) );
  NANDN U134 ( .A(n7923), .B(n7924), .Z(n66) );
  NAND U135 ( .A(n65), .B(n66), .Z(n8080) );
  NANDN U136 ( .A(n8126), .B(n8127), .Z(n67) );
  NANDN U137 ( .A(n8125), .B(n8124), .Z(n68) );
  AND U138 ( .A(n67), .B(n68), .Z(n8251) );
  NANDN U139 ( .A(n8122), .B(n8123), .Z(n69) );
  NANDN U140 ( .A(n8121), .B(n8120), .Z(n70) );
  AND U141 ( .A(n69), .B(n70), .Z(n8229) );
  NANDN U142 ( .A(n8234), .B(n8233), .Z(n71) );
  NANDN U143 ( .A(n8231), .B(n8232), .Z(n72) );
  AND U144 ( .A(n71), .B(n72), .Z(n8339) );
  NANDN U145 ( .A(n8347), .B(n8348), .Z(n73) );
  NANDN U146 ( .A(n8349), .B(n8350), .Z(n74) );
  AND U147 ( .A(n73), .B(n74), .Z(n8443) );
  NANDN U148 ( .A(n8627), .B(n8628), .Z(n75) );
  NANDN U149 ( .A(n8626), .B(n8625), .Z(n76) );
  NAND U150 ( .A(n75), .B(n76), .Z(n8678) );
  NAND U151 ( .A(n8814), .B(n8813), .Z(n77) );
  NANDN U152 ( .A(n8811), .B(n8812), .Z(n78) );
  AND U153 ( .A(n77), .B(n78), .Z(n8905) );
  NANDN U154 ( .A(n8885), .B(n8886), .Z(n79) );
  NANDN U155 ( .A(n8887), .B(n8888), .Z(n80) );
  AND U156 ( .A(n79), .B(n80), .Z(n8996) );
  NANDN U157 ( .A(n8936), .B(n8937), .Z(n81) );
  NANDN U158 ( .A(n8938), .B(n8939), .Z(n82) );
  AND U159 ( .A(n81), .B(n82), .Z(n9024) );
  NANDN U160 ( .A(n7504), .B(n7503), .Z(n83) );
  NANDN U161 ( .A(n7501), .B(n7502), .Z(n84) );
  AND U162 ( .A(n83), .B(n84), .Z(n7620) );
  NANDN U163 ( .A(n7722), .B(n7723), .Z(n85) );
  NANDN U164 ( .A(n7724), .B(n7725), .Z(n86) );
  AND U165 ( .A(n85), .B(n86), .Z(n7749) );
  NANDN U166 ( .A(n7962), .B(n7963), .Z(n87) );
  NANDN U167 ( .A(n7964), .B(n7965), .Z(n88) );
  AND U168 ( .A(n87), .B(n88), .Z(n8090) );
  NANDN U169 ( .A(n7985), .B(n7984), .Z(n89) );
  NANDN U170 ( .A(n7982), .B(n7983), .Z(n90) );
  AND U171 ( .A(n89), .B(n90), .Z(n8110) );
  NANDN U172 ( .A(n8248), .B(n8247), .Z(n91) );
  NANDN U173 ( .A(n8245), .B(n8246), .Z(n92) );
  AND U174 ( .A(n91), .B(n92), .Z(n8334) );
  NANDN U175 ( .A(n8422), .B(n8423), .Z(n93) );
  NANDN U176 ( .A(n8425), .B(n8424), .Z(n94) );
  NAND U177 ( .A(n93), .B(n94), .Z(n8533) );
  NANDN U178 ( .A(n8548), .B(n8549), .Z(n95) );
  NANDN U179 ( .A(n8550), .B(n8551), .Z(n96) );
  AND U180 ( .A(n95), .B(n96), .Z(n8662) );
  NANDN U181 ( .A(n8666), .B(n8665), .Z(n97) );
  NANDN U182 ( .A(n8663), .B(n8664), .Z(n98) );
  AND U183 ( .A(n97), .B(n98), .Z(n8824) );
  NANDN U184 ( .A(n8805), .B(n8806), .Z(n99) );
  NANDN U185 ( .A(n8804), .B(n8803), .Z(n100) );
  AND U186 ( .A(n99), .B(n100), .Z(n8838) );
  NAND U187 ( .A(n8756), .B(n8757), .Z(n101) );
  NANDN U188 ( .A(n8754), .B(n8755), .Z(n102) );
  AND U189 ( .A(n101), .B(n102), .Z(n8908) );
  OR U190 ( .A(n8900), .B(n8901), .Z(n103) );
  NANDN U191 ( .A(n8902), .B(n8903), .Z(n104) );
  AND U192 ( .A(n103), .B(n104), .Z(n8928) );
  NANDN U193 ( .A(n9062), .B(n9063), .Z(n105) );
  NANDN U194 ( .A(n9065), .B(n9064), .Z(n106) );
  NAND U195 ( .A(n105), .B(n106), .Z(n9163) );
  NAND U196 ( .A(n9029), .B(n9028), .Z(n107) );
  NANDN U197 ( .A(n9026), .B(n9027), .Z(n108) );
  NAND U198 ( .A(n107), .B(n108), .Z(n9099) );
  NANDN U199 ( .A(n9155), .B(n9156), .Z(n109) );
  NANDN U200 ( .A(n9157), .B(n9158), .Z(n110) );
  AND U201 ( .A(n109), .B(n110), .Z(n9181) );
  NANDN U202 ( .A(n9244), .B(n9243), .Z(n111) );
  NANDN U203 ( .A(n9241), .B(n9242), .Z(n112) );
  AND U204 ( .A(n111), .B(n112), .Z(n9257) );
  NANDN U205 ( .A(n9306), .B(n9307), .Z(n113) );
  NANDN U206 ( .A(n9305), .B(n9304), .Z(n114) );
  AND U207 ( .A(n113), .B(n114), .Z(n9330) );
  NANDN U208 ( .A(n9336), .B(n9337), .Z(n115) );
  NANDN U209 ( .A(n9335), .B(n9334), .Z(n116) );
  AND U210 ( .A(n115), .B(n116), .Z(n9403) );
  NANDN U211 ( .A(n9405), .B(n9406), .Z(n117) );
  NANDN U212 ( .A(n9407), .B(n9408), .Z(n118) );
  AND U213 ( .A(n117), .B(n118), .Z(n9504) );
  NANDN U214 ( .A(n9493), .B(n9494), .Z(n119) );
  NANDN U215 ( .A(n9491), .B(n9492), .Z(n120) );
  NAND U216 ( .A(n119), .B(n120), .Z(n9517) );
  NANDN U217 ( .A(n9589), .B(n9590), .Z(n121) );
  NANDN U218 ( .A(n9588), .B(n9611), .Z(n122) );
  AND U219 ( .A(n121), .B(n122), .Z(n9623) );
  NANDN U220 ( .A(n9649), .B(n9650), .Z(n123) );
  NANDN U221 ( .A(n9647), .B(n9648), .Z(n124) );
  NAND U222 ( .A(n123), .B(n124), .Z(n9677) );
  NAND U223 ( .A(n9658), .B(n9657), .Z(n125) );
  NANDN U224 ( .A(n9655), .B(n9656), .Z(n126) );
  NAND U225 ( .A(n125), .B(n126), .Z(n9672) );
  OR U226 ( .A(n9726), .B(n9698), .Z(n127) );
  NANDN U227 ( .A(n9700), .B(n9699), .Z(n128) );
  NAND U228 ( .A(n127), .B(n128), .Z(n9713) );
  NANDN U229 ( .A(n7493), .B(n7494), .Z(n129) );
  NANDN U230 ( .A(n7495), .B(n7496), .Z(n130) );
  AND U231 ( .A(n129), .B(n130), .Z(n7738) );
  NANDN U232 ( .A(n7752), .B(n7753), .Z(n131) );
  NANDN U233 ( .A(n7755), .B(n7754), .Z(n132) );
  NAND U234 ( .A(n131), .B(n132), .Z(n7971) );
  NANDN U235 ( .A(n9558), .B(n9559), .Z(n133) );
  NANDN U236 ( .A(n9560), .B(n9561), .Z(n134) );
  AND U237 ( .A(n133), .B(n134), .Z(n9571) );
  NANDN U238 ( .A(n9578), .B(n9579), .Z(n135) );
  NANDN U239 ( .A(n9580), .B(n9581), .Z(n136) );
  AND U240 ( .A(n135), .B(n136), .Z(n9618) );
  OR U241 ( .A(n9858), .B(n9830), .Z(n137) );
  NANDN U242 ( .A(n9832), .B(n9831), .Z(n138) );
  AND U243 ( .A(n137), .B(n138), .Z(n9866) );
  NANDN U244 ( .A(n7773), .B(n7772), .Z(n139) );
  NANDN U245 ( .A(n7770), .B(n7771), .Z(n140) );
  AND U246 ( .A(n139), .B(n140), .Z(n7961) );
  NANDN U247 ( .A(n7790), .B(n7791), .Z(n141) );
  NANDN U248 ( .A(n7792), .B(n7793), .Z(n142) );
  AND U249 ( .A(n141), .B(n142), .Z(n7874) );
  NANDN U250 ( .A(n7515), .B(n7516), .Z(n143) );
  NANDN U251 ( .A(n7517), .B(n7518), .Z(n144) );
  AND U252 ( .A(n143), .B(n144), .Z(n7719) );
  NANDN U253 ( .A(n7558), .B(n7559), .Z(n145) );
  NANDN U254 ( .A(n7557), .B(n7556), .Z(n146) );
  AND U255 ( .A(n145), .B(n146), .Z(n7722) );
  NANDN U256 ( .A(n7668), .B(n7669), .Z(n147) );
  NANDN U257 ( .A(n7670), .B(n7671), .Z(n148) );
  AND U258 ( .A(n147), .B(n148), .Z(n7758) );
  NANDN U259 ( .A(n7929), .B(n7930), .Z(n149) );
  NANDN U260 ( .A(n7927), .B(n7928), .Z(n150) );
  NAND U261 ( .A(n149), .B(n150), .Z(n8082) );
  NANDN U262 ( .A(n8207), .B(n8208), .Z(n151) );
  NANDN U263 ( .A(n8206), .B(n8205), .Z(n152) );
  AND U264 ( .A(n151), .B(n152), .Z(n8245) );
  NANDN U265 ( .A(n8995), .B(n8994), .Z(n153) );
  NANDN U266 ( .A(n8992), .B(n8993), .Z(n154) );
  AND U267 ( .A(n153), .B(n154), .Z(n9028) );
  NANDN U268 ( .A(n8197), .B(n8198), .Z(n155) );
  NANDN U269 ( .A(n8199), .B(n8200), .Z(n156) );
  AND U270 ( .A(n155), .B(n156), .Z(n8321) );
  NANDN U271 ( .A(n8229), .B(n8230), .Z(n157) );
  NANDN U272 ( .A(n8228), .B(n8227), .Z(n158) );
  AND U273 ( .A(n157), .B(n158), .Z(n8335) );
  NANDN U274 ( .A(n8370), .B(n8371), .Z(n159) );
  NANDN U275 ( .A(n8372), .B(n8373), .Z(n160) );
  AND U276 ( .A(n159), .B(n160), .Z(n8526) );
  NANDN U277 ( .A(n8340), .B(n8339), .Z(n161) );
  NANDN U278 ( .A(n8337), .B(n8338), .Z(n162) );
  AND U279 ( .A(n161), .B(n162), .Z(n8534) );
  NAND U280 ( .A(n8443), .B(n8442), .Z(n163) );
  NANDN U281 ( .A(n8444), .B(n8445), .Z(n164) );
  AND U282 ( .A(n163), .B(n164), .Z(n8631) );
  NAND U283 ( .A(n8507), .B(n8506), .Z(n165) );
  NANDN U284 ( .A(n8508), .B(n8509), .Z(n166) );
  AND U285 ( .A(n165), .B(n166), .Z(n8636) );
  NAND U286 ( .A(n8613), .B(n8614), .Z(n167) );
  NANDN U287 ( .A(n8611), .B(n8612), .Z(n168) );
  AND U288 ( .A(n167), .B(n168), .Z(n8655) );
  NANDN U289 ( .A(n8680), .B(n8679), .Z(n169) );
  NANDN U290 ( .A(n8677), .B(n8678), .Z(n170) );
  AND U291 ( .A(n169), .B(n170), .Z(n8826) );
  NANDN U292 ( .A(n8750), .B(n8751), .Z(n171) );
  NANDN U293 ( .A(n8752), .B(n8753), .Z(n172) );
  AND U294 ( .A(n171), .B(n172), .Z(n8910) );
  NANDN U295 ( .A(n9004), .B(n9005), .Z(n173) );
  NANDN U296 ( .A(n9002), .B(n9003), .Z(n174) );
  NAND U297 ( .A(n173), .B(n174), .Z(n9018) );
  NANDN U298 ( .A(n9025), .B(n9024), .Z(n175) );
  NANDN U299 ( .A(n9022), .B(n9023), .Z(n176) );
  AND U300 ( .A(n175), .B(n176), .Z(n9100) );
  NANDN U301 ( .A(n9653), .B(n9654), .Z(n177) );
  NANDN U302 ( .A(n9651), .B(n9652), .Z(n178) );
  AND U303 ( .A(n177), .B(n178), .Z(n9671) );
  NANDN U304 ( .A(n9744), .B(n9743), .Z(n179) );
  NANDN U305 ( .A(n9741), .B(n9742), .Z(n180) );
  AND U306 ( .A(n179), .B(n180), .Z(n9777) );
  NANDN U307 ( .A(n9758), .B(n9759), .Z(n181) );
  NANDN U308 ( .A(n9757), .B(n9767), .Z(n182) );
  AND U309 ( .A(n181), .B(n182), .Z(n9793) );
  NAND U310 ( .A(n9808), .B(n582), .Z(n183) );
  AND U311 ( .A(n9809), .B(n183), .Z(n9830) );
  NANDN U312 ( .A(n7620), .B(n7621), .Z(n184) );
  NANDN U313 ( .A(n7622), .B(n7623), .Z(n185) );
  AND U314 ( .A(n184), .B(n185), .Z(n7855) );
  NANDN U315 ( .A(n7969), .B(n7968), .Z(n186) );
  NANDN U316 ( .A(n7966), .B(n7967), .Z(n187) );
  AND U317 ( .A(n186), .B(n187), .Z(n8094) );
  NANDN U318 ( .A(n8084), .B(n8085), .Z(n188) );
  NANDN U319 ( .A(n8086), .B(n8087), .Z(n189) );
  AND U320 ( .A(n188), .B(n189), .Z(n8106) );
  NANDN U321 ( .A(n8110), .B(n8111), .Z(n190) );
  NANDN U322 ( .A(n8112), .B(n8113), .Z(n191) );
  AND U323 ( .A(n190), .B(n191), .Z(n8225) );
  NAND U324 ( .A(n8429), .B(n8428), .Z(n192) );
  NANDN U325 ( .A(n8426), .B(n8427), .Z(n193) );
  NAND U326 ( .A(n192), .B(n193), .Z(n8536) );
  OR U327 ( .A(n8659), .B(n8660), .Z(n194) );
  NANDN U328 ( .A(n8661), .B(n8662), .Z(n195) );
  AND U329 ( .A(n194), .B(n195), .Z(n8747) );
  NANDN U330 ( .A(n8825), .B(n8824), .Z(n196) );
  NANDN U331 ( .A(n8822), .B(n8823), .Z(n197) );
  AND U332 ( .A(n196), .B(n197), .Z(n8912) );
  NANDN U333 ( .A(n8841), .B(n8840), .Z(n198) );
  NANDN U334 ( .A(n8838), .B(n8839), .Z(n199) );
  AND U335 ( .A(n198), .B(n199), .Z(n8925) );
  NANDN U336 ( .A(n8932), .B(n8933), .Z(n200) );
  NANDN U337 ( .A(n8934), .B(n8935), .Z(n201) );
  AND U338 ( .A(n200), .B(n201), .Z(n9015) );
  NANDN U339 ( .A(n9181), .B(n9182), .Z(n202) );
  NANDN U340 ( .A(n9183), .B(n9184), .Z(n203) );
  AND U341 ( .A(n202), .B(n203), .Z(n9255) );
  NAND U342 ( .A(n9258), .B(n9257), .Z(n204) );
  NANDN U343 ( .A(n9259), .B(n9260), .Z(n205) );
  NAND U344 ( .A(n204), .B(n205), .Z(n9329) );
  NANDN U345 ( .A(n9330), .B(n9331), .Z(n206) );
  NANDN U346 ( .A(n9332), .B(n9333), .Z(n207) );
  AND U347 ( .A(n206), .B(n207), .Z(n9393) );
  NANDN U348 ( .A(n9404), .B(n9403), .Z(n208) );
  NANDN U349 ( .A(n9401), .B(n9402), .Z(n209) );
  AND U350 ( .A(n208), .B(n209), .Z(n9457) );
  NAND U351 ( .A(n9504), .B(n9503), .Z(n210) );
  NANDN U352 ( .A(n9501), .B(n9502), .Z(n211) );
  NAND U353 ( .A(n210), .B(n211), .Z(n9515) );
  NANDN U354 ( .A(n9520), .B(n9519), .Z(n212) );
  NANDN U355 ( .A(n9517), .B(n9518), .Z(n213) );
  AND U356 ( .A(n212), .B(n213), .Z(n9572) );
  NANDN U357 ( .A(n9577), .B(n9576), .Z(n214) );
  NANDN U358 ( .A(n9574), .B(n9575), .Z(n215) );
  AND U359 ( .A(n214), .B(n215), .Z(n9621) );
  NANDN U360 ( .A(n9624), .B(n9625), .Z(n216) );
  NANDN U361 ( .A(n9622), .B(n9623), .Z(n217) );
  NAND U362 ( .A(n216), .B(n217), .Z(n9669) );
  NANDN U363 ( .A(n9677), .B(n9678), .Z(n218) );
  NANDN U364 ( .A(n9676), .B(n9675), .Z(n219) );
  AND U365 ( .A(n218), .B(n219), .Z(n9709) );
  NANDN U366 ( .A(n9813), .B(n9812), .Z(n220) );
  NANDN U367 ( .A(n9810), .B(n9811), .Z(n221) );
  AND U368 ( .A(n220), .B(n221), .Z(n9840) );
  NANDN U369 ( .A(n7973), .B(n7972), .Z(n222) );
  NANDN U370 ( .A(n7970), .B(n7971), .Z(n223) );
  AND U371 ( .A(n222), .B(n223), .Z(n7976) );
  NANDN U372 ( .A(n9854), .B(n9853), .Z(n224) );
  NANDN U373 ( .A(n9851), .B(n9852), .Z(n225) );
  AND U374 ( .A(n224), .B(n225), .Z(n9889) );
  NANDN U375 ( .A(n7618), .B(n7619), .Z(n226) );
  NANDN U376 ( .A(n7616), .B(n7617), .Z(n227) );
  NAND U377 ( .A(n226), .B(n227), .Z(n7746) );
  NANDN U378 ( .A(n2832), .B(n2833), .Z(n228) );
  NANDN U379 ( .A(n2831), .B(n2830), .Z(n229) );
  AND U380 ( .A(n228), .B(n229), .Z(n3017) );
  NANDN U381 ( .A(n3461), .B(n3462), .Z(n230) );
  NANDN U382 ( .A(n3460), .B(n3459), .Z(n231) );
  AND U383 ( .A(n230), .B(n231), .Z(n3503) );
  OR U384 ( .A(n7532), .B(n7533), .Z(n232) );
  NANDN U385 ( .A(n7530), .B(n7531), .Z(n233) );
  NAND U386 ( .A(n232), .B(n233), .Z(n7675) );
  NANDN U387 ( .A(n7590), .B(n7591), .Z(n234) );
  NANDN U388 ( .A(n7592), .B(n7593), .Z(n235) );
  AND U389 ( .A(n234), .B(n235), .Z(n7668) );
  OR U390 ( .A(n7632), .B(n7633), .Z(n236) );
  NANDN U391 ( .A(n7630), .B(n7631), .Z(n237) );
  AND U392 ( .A(n236), .B(n237), .Z(n7847) );
  NANDN U393 ( .A(n7837), .B(n7838), .Z(n238) );
  NANDN U394 ( .A(n7839), .B(n7840), .Z(n239) );
  AND U395 ( .A(n238), .B(n239), .Z(n7869) );
  NANDN U396 ( .A(n8048), .B(n8049), .Z(n240) );
  NANDN U397 ( .A(n8051), .B(n8050), .Z(n241) );
  NAND U398 ( .A(n240), .B(n241), .Z(n8207) );
  NANDN U399 ( .A(n8285), .B(n8284), .Z(n242) );
  NANDN U400 ( .A(n8282), .B(n8283), .Z(n243) );
  AND U401 ( .A(n242), .B(n243), .Z(n8374) );
  NANDN U402 ( .A(n8729), .B(n8730), .Z(n244) );
  NANDN U403 ( .A(n8727), .B(n8728), .Z(n245) );
  NAND U404 ( .A(n244), .B(n245), .Z(n8760) );
  NANDN U405 ( .A(n1598), .B(n1599), .Z(n246) );
  NANDN U406 ( .A(n1597), .B(n1596), .Z(n247) );
  AND U407 ( .A(n246), .B(n247), .Z(n1706) );
  NANDN U408 ( .A(n7381), .B(n7380), .Z(n248) );
  NANDN U409 ( .A(n7378), .B(n7379), .Z(n249) );
  AND U410 ( .A(n248), .B(n249), .Z(n7599) );
  NANDN U411 ( .A(n7555), .B(n7554), .Z(n250) );
  NANDN U412 ( .A(n7552), .B(n7553), .Z(n251) );
  AND U413 ( .A(n250), .B(n251), .Z(n7724) );
  NANDN U414 ( .A(n7666), .B(n7667), .Z(n252) );
  NANDN U415 ( .A(n7664), .B(n7665), .Z(n253) );
  NAND U416 ( .A(n252), .B(n253), .Z(n7851) );
  NANDN U417 ( .A(n7805), .B(n7804), .Z(n254) );
  NANDN U418 ( .A(n7802), .B(n7803), .Z(n255) );
  AND U419 ( .A(n254), .B(n255), .Z(n7897) );
  OR U420 ( .A(n7959), .B(n7958), .Z(n256) );
  NANDN U421 ( .A(n7960), .B(n7961), .Z(n257) );
  NAND U422 ( .A(n256), .B(n257), .Z(n7988) );
  NAND U423 ( .A(n7876), .B(n7875), .Z(n258) );
  NANDN U424 ( .A(n7873), .B(n7874), .Z(n259) );
  NAND U425 ( .A(n258), .B(n259), .Z(n7983) );
  XOR U426 ( .A(n8316), .B(n8315), .Z(n8318) );
  NANDN U427 ( .A(n8253), .B(n8254), .Z(n260) );
  NANDN U428 ( .A(n8255), .B(n8256), .Z(n261) );
  AND U429 ( .A(n260), .B(n261), .Z(n8371) );
  NAND U430 ( .A(n8563), .B(n8564), .Z(n262) );
  NANDN U431 ( .A(n8561), .B(n8562), .Z(n263) );
  AND U432 ( .A(n262), .B(n263), .Z(n8667) );
  NANDN U433 ( .A(n8782), .B(n8783), .Z(n264) );
  NANDN U434 ( .A(n8780), .B(n8781), .Z(n265) );
  NAND U435 ( .A(n264), .B(n265), .Z(n8895) );
  NAND U436 ( .A(n8802), .B(n8801), .Z(n266) );
  NANDN U437 ( .A(n8799), .B(n8800), .Z(n267) );
  NAND U438 ( .A(n266), .B(n267), .Z(n8891) );
  OR U439 ( .A(n8943), .B(n8846), .Z(n268) );
  NANDN U440 ( .A(n8848), .B(n8847), .Z(n269) );
  AND U441 ( .A(n268), .B(n269), .Z(n8976) );
  NANDN U442 ( .A(n9077), .B(n9076), .Z(n270) );
  NANDN U443 ( .A(n9074), .B(n9075), .Z(n271) );
  AND U444 ( .A(n270), .B(n271), .Z(n9156) );
  NANDN U445 ( .A(n9153), .B(n9154), .Z(n272) );
  NANDN U446 ( .A(n9151), .B(n9152), .Z(n273) );
  NAND U447 ( .A(n272), .B(n273), .Z(n9242) );
  NANDN U448 ( .A(n9109), .B(n9110), .Z(n274) );
  NANDN U449 ( .A(n9112), .B(n9111), .Z(n275) );
  NAND U450 ( .A(n274), .B(n275), .Z(n9239) );
  NANDN U451 ( .A(n9201), .B(n9202), .Z(n276) );
  NANDN U452 ( .A(n9203), .B(n9204), .Z(n277) );
  AND U453 ( .A(n276), .B(n277), .Z(n9308) );
  NANDN U454 ( .A(n7720), .B(n7721), .Z(n278) );
  NANDN U455 ( .A(n7718), .B(n7719), .Z(n279) );
  NAND U456 ( .A(n278), .B(n279), .Z(n7752) );
  NANDN U457 ( .A(n8082), .B(n8083), .Z(n280) );
  NANDN U458 ( .A(n8080), .B(n8081), .Z(n281) );
  NAND U459 ( .A(n280), .B(n281), .Z(n8114) );
  NANDN U460 ( .A(n8249), .B(n8250), .Z(n282) );
  NANDN U461 ( .A(n8251), .B(n8252), .Z(n283) );
  AND U462 ( .A(n282), .B(n283), .Z(n8429) );
  NANDN U463 ( .A(n9591), .B(n9592), .Z(n284) );
  NANDN U464 ( .A(n9593), .B(n9594), .Z(n285) );
  AND U465 ( .A(n284), .B(n285), .Z(n9629) );
  NANDN U466 ( .A(n9681), .B(n9682), .Z(n286) );
  NANDN U467 ( .A(n9679), .B(n9680), .Z(n287) );
  NAND U468 ( .A(n286), .B(n287), .Z(n9715) );
  NANDN U469 ( .A(n7497), .B(n7498), .Z(n288) );
  NANDN U470 ( .A(n7500), .B(n7499), .Z(n289) );
  NAND U471 ( .A(n288), .B(n289), .Z(n7736) );
  NAND U472 ( .A(n7867), .B(n7868), .Z(n290) );
  NANDN U473 ( .A(n7865), .B(n7866), .Z(n291) );
  AND U474 ( .A(n290), .B(n291), .Z(n8096) );
  NANDN U475 ( .A(n8321), .B(n8322), .Z(n292) );
  NANDN U476 ( .A(n8324), .B(n8323), .Z(n293) );
  NAND U477 ( .A(n292), .B(n293), .Z(n8432) );
  NANDN U478 ( .A(n8333), .B(n8334), .Z(n294) );
  NANDN U479 ( .A(n8335), .B(n8336), .Z(n295) );
  AND U480 ( .A(n294), .B(n295), .Z(n8538) );
  NANDN U481 ( .A(n8534), .B(n8535), .Z(n296) );
  NANDN U482 ( .A(n8532), .B(n8533), .Z(n297) );
  NAND U483 ( .A(n296), .B(n297), .Z(n8641) );
  NANDN U484 ( .A(n8637), .B(n8638), .Z(n298) );
  NANDN U485 ( .A(n8635), .B(n8636), .Z(n299) );
  NAND U486 ( .A(n298), .B(n299), .Z(n8653) );
  NANDN U487 ( .A(n8658), .B(n8657), .Z(n300) );
  NANDN U488 ( .A(n8655), .B(n8656), .Z(n301) );
  AND U489 ( .A(n300), .B(n301), .Z(n8748) );
  NAND U490 ( .A(n8829), .B(n8828), .Z(n302) );
  NANDN U491 ( .A(n8826), .B(n8827), .Z(n303) );
  NAND U492 ( .A(n302), .B(n303), .Z(n8914) );
  NANDN U493 ( .A(n8910), .B(n8911), .Z(n304) );
  NANDN U494 ( .A(n8908), .B(n8909), .Z(n305) );
  NAND U495 ( .A(n304), .B(n305), .Z(n8926) );
  NAND U496 ( .A(n8930), .B(n8931), .Z(n306) );
  NANDN U497 ( .A(n8928), .B(n8929), .Z(n307) );
  AND U498 ( .A(n306), .B(n307), .Z(n9017) );
  NANDN U499 ( .A(n9018), .B(n9019), .Z(n308) );
  NANDN U500 ( .A(n9021), .B(n9020), .Z(n309) );
  NAND U501 ( .A(n308), .B(n309), .Z(n9095) );
  NANDN U502 ( .A(n9099), .B(n9100), .Z(n310) );
  NANDN U503 ( .A(n9101), .B(n9102), .Z(n311) );
  AND U504 ( .A(n310), .B(n311), .Z(n9179) );
  NANDN U505 ( .A(n9381), .B(n9382), .Z(n312) );
  NANDN U506 ( .A(n9384), .B(n9383), .Z(n313) );
  NAND U507 ( .A(n312), .B(n313), .Z(n9391) );
  NANDN U508 ( .A(n9399), .B(n9400), .Z(n314) );
  NANDN U509 ( .A(n9398), .B(n9397), .Z(n315) );
  AND U510 ( .A(n314), .B(n315), .Z(n9458) );
  NANDN U511 ( .A(n9674), .B(n9673), .Z(n316) );
  NANDN U512 ( .A(n9671), .B(n9672), .Z(n317) );
  AND U513 ( .A(n316), .B(n317), .Z(n9711) );
  NANDN U514 ( .A(n9721), .B(n9722), .Z(n318) );
  NANDN U515 ( .A(n9719), .B(n9720), .Z(n319) );
  NAND U516 ( .A(n318), .B(n319), .Z(n9754) );
  NANDN U517 ( .A(n9775), .B(n9776), .Z(n320) );
  NANDN U518 ( .A(n9773), .B(n9774), .Z(n321) );
  NAND U519 ( .A(n320), .B(n321), .Z(n9815) );
  NANDN U520 ( .A(n9794), .B(n9793), .Z(n322) );
  NANDN U521 ( .A(n9791), .B(n9792), .Z(n323) );
  AND U522 ( .A(n322), .B(n323), .Z(n9841) );
  NANDN U523 ( .A(n9829), .B(n9828), .Z(n324) );
  NANDN U524 ( .A(n9826), .B(n9827), .Z(n325) );
  AND U525 ( .A(n324), .B(n325), .Z(n9868) );
  NANDN U526 ( .A(n7604), .B(n7605), .Z(n326) );
  NANDN U527 ( .A(n7602), .B(n7603), .Z(n327) );
  NAND U528 ( .A(n326), .B(n327), .Z(n7617) );
  NANDN U529 ( .A(n8109), .B(n8108), .Z(n328) );
  NANDN U530 ( .A(n8106), .B(n8107), .Z(n329) );
  AND U531 ( .A(n328), .B(n329), .Z(n8218) );
  NANDN U532 ( .A(n9255), .B(n9256), .Z(n330) );
  NANDN U533 ( .A(n9254), .B(n9253), .Z(n331) );
  NAND U534 ( .A(n330), .B(n331), .Z(n9320) );
  NAND U535 ( .A(n9327), .B(n9326), .Z(n332) );
  NANDN U536 ( .A(n9328), .B(n9329), .Z(n333) );
  AND U537 ( .A(n332), .B(n333), .Z(n9387) );
  NANDN U538 ( .A(n9513), .B(n9514), .Z(n334) );
  NANDN U539 ( .A(n9515), .B(n9516), .Z(n335) );
  AND U540 ( .A(n334), .B(n335), .Z(n9565) );
  NANDN U541 ( .A(n9572), .B(n9573), .Z(n336) );
  NANDN U542 ( .A(n9570), .B(n9571), .Z(n337) );
  NAND U543 ( .A(n336), .B(n337), .Z(n9615) );
  NAND U544 ( .A(n9621), .B(n9620), .Z(n338) );
  NANDN U545 ( .A(n9618), .B(n9619), .Z(n339) );
  NAND U546 ( .A(n338), .B(n339), .Z(n9661) );
  NAND U547 ( .A(n621), .B(n622), .Z(n340) );
  XOR U548 ( .A(n621), .B(n622), .Z(n341) );
  NANDN U549 ( .A(n620), .B(n341), .Z(n342) );
  NAND U550 ( .A(n340), .B(n342), .Z(n635) );
  NANDN U551 ( .A(n7861), .B(n7862), .Z(n343) );
  NANDN U552 ( .A(n7864), .B(n7863), .Z(n344) );
  NAND U553 ( .A(n343), .B(n344), .Z(n7978) );
  NANDN U554 ( .A(n9887), .B(n9888), .Z(n345) );
  NANDN U555 ( .A(n9889), .B(n9890), .Z(n346) );
  AND U556 ( .A(n345), .B(n346), .Z(n9891) );
  NAND U557 ( .A(n2762), .B(n2763), .Z(n347) );
  XOR U558 ( .A(n2762), .B(n2763), .Z(n348) );
  NAND U559 ( .A(n348), .B(sreg[62]), .Z(n349) );
  NAND U560 ( .A(n347), .B(n349), .Z(n2902) );
  NANDN U561 ( .A(b[0]), .B(a[63]), .Z(n350) );
  AND U562 ( .A(b[1]), .B(n350), .Z(n7772) );
  NANDN U563 ( .A(n2658), .B(n2659), .Z(n351) );
  NANDN U564 ( .A(n2657), .B(n2656), .Z(n352) );
  NAND U565 ( .A(n351), .B(n352), .Z(n2776) );
  NANDN U566 ( .A(n4017), .B(n4018), .Z(n353) );
  NANDN U567 ( .A(n4016), .B(n4015), .Z(n354) );
  AND U568 ( .A(n353), .B(n354), .Z(n4207) );
  NANDN U569 ( .A(n5058), .B(n5059), .Z(n355) );
  NANDN U570 ( .A(n5057), .B(n5056), .Z(n356) );
  AND U571 ( .A(n355), .B(n356), .Z(n5252) );
  NANDN U572 ( .A(n5193), .B(n5194), .Z(n357) );
  NANDN U573 ( .A(n5192), .B(n5191), .Z(n358) );
  AND U574 ( .A(n357), .B(n358), .Z(n5399) );
  NANDN U575 ( .A(n5340), .B(n5341), .Z(n359) );
  NANDN U576 ( .A(n5339), .B(n5338), .Z(n360) );
  AND U577 ( .A(n359), .B(n360), .Z(n5548) );
  NANDN U578 ( .A(n5946), .B(n5947), .Z(n361) );
  NANDN U579 ( .A(n5945), .B(n5944), .Z(n362) );
  AND U580 ( .A(n361), .B(n362), .Z(n6134) );
  NANDN U581 ( .A(n6075), .B(n6076), .Z(n363) );
  NANDN U582 ( .A(n6074), .B(n6073), .Z(n364) );
  AND U583 ( .A(n363), .B(n364), .Z(n6289) );
  NANDN U584 ( .A(n6389), .B(n6390), .Z(n365) );
  NANDN U585 ( .A(n6388), .B(n6387), .Z(n366) );
  AND U586 ( .A(n365), .B(n366), .Z(n6585) );
  OR U587 ( .A(n7358), .B(n7359), .Z(n367) );
  NANDN U588 ( .A(n7356), .B(n7357), .Z(n368) );
  AND U589 ( .A(n367), .B(n368), .Z(n7558) );
  NANDN U590 ( .A(n7436), .B(n7437), .Z(n369) );
  NANDN U591 ( .A(n7439), .B(n7438), .Z(n370) );
  NAND U592 ( .A(n369), .B(n370), .Z(n7553) );
  NANDN U593 ( .A(n7932), .B(n7933), .Z(n371) );
  NANDN U594 ( .A(b[1]), .B(n7931), .Z(n372) );
  AND U595 ( .A(n371), .B(n372), .Z(n8076) );
  NANDN U596 ( .A(n7798), .B(n7799), .Z(n373) );
  NANDN U597 ( .A(n7800), .B(n7801), .Z(n374) );
  AND U598 ( .A(n373), .B(n374), .Z(n7875) );
  NANDN U599 ( .A(n7891), .B(n7892), .Z(n375) );
  NANDN U600 ( .A(n7893), .B(n7894), .Z(n376) );
  AND U601 ( .A(n375), .B(n376), .Z(n7992) );
  NANDN U602 ( .A(n8070), .B(n8071), .Z(n377) );
  NANDN U603 ( .A(n8072), .B(n8073), .Z(n378) );
  AND U604 ( .A(n377), .B(n378), .Z(n8211) );
  NANDN U605 ( .A(n8166), .B(n8167), .Z(n379) );
  NANDN U606 ( .A(n8168), .B(n8169), .Z(n380) );
  AND U607 ( .A(n379), .B(n380), .Z(n8241) );
  NANDN U608 ( .A(n8149), .B(n8150), .Z(n381) );
  NANDN U609 ( .A(n8147), .B(n8148), .Z(n382) );
  NAND U610 ( .A(n381), .B(n382), .Z(n8237) );
  NANDN U611 ( .A(n8192), .B(n8191), .Z(n383) );
  NANDN U612 ( .A(n8189), .B(n8190), .Z(n384) );
  AND U613 ( .A(n383), .B(n384), .Z(n8231) );
  NANDN U614 ( .A(n8351), .B(n8352), .Z(n385) );
  NANDN U615 ( .A(n8353), .B(n8354), .Z(n386) );
  AND U616 ( .A(n385), .B(n386), .Z(n8516) );
  NANDN U617 ( .A(n8595), .B(n8596), .Z(n387) );
  NANDN U618 ( .A(n8597), .B(n8598), .Z(n388) );
  AND U619 ( .A(n387), .B(n388), .Z(n8683) );
  NANDN U620 ( .A(n2074), .B(n2075), .Z(n389) );
  NANDN U621 ( .A(n2073), .B(n2072), .Z(n390) );
  AND U622 ( .A(n389), .B(n390), .Z(n2230) );
  NANDN U623 ( .A(n2878), .B(n2879), .Z(n391) );
  NANDN U624 ( .A(n2881), .B(n2880), .Z(n392) );
  NAND U625 ( .A(n391), .B(n392), .Z(n3027) );
  NANDN U626 ( .A(n3356), .B(n3355), .Z(n393) );
  NANDN U627 ( .A(n3353), .B(n3354), .Z(n394) );
  AND U628 ( .A(n393), .B(n394), .Z(n3628) );
  NANDN U629 ( .A(n7283), .B(n7284), .Z(n395) );
  NANDN U630 ( .A(n7282), .B(n7281), .Z(n396) );
  AND U631 ( .A(n395), .B(n396), .Z(n7461) );
  NANDN U632 ( .A(n7528), .B(n7529), .Z(n397) );
  NANDN U633 ( .A(n7526), .B(n7527), .Z(n398) );
  NAND U634 ( .A(n397), .B(n398), .Z(n7720) );
  NANDN U635 ( .A(n7847), .B(n7848), .Z(n399) );
  NANDN U636 ( .A(n7846), .B(n7845), .Z(n400) );
  AND U637 ( .A(n399), .B(n400), .Z(n7895) );
  NANDN U638 ( .A(n7869), .B(n7870), .Z(n401) );
  NANDN U639 ( .A(n7871), .B(n7872), .Z(n402) );
  AND U640 ( .A(n401), .B(n402), .Z(n7984) );
  NANDN U641 ( .A(n8028), .B(n8029), .Z(n403) );
  NANDN U642 ( .A(n8027), .B(n8026), .Z(n404) );
  NAND U643 ( .A(n403), .B(n404), .Z(n8198) );
  NANDN U644 ( .A(n8185), .B(n8186), .Z(n405) );
  NANDN U645 ( .A(n8187), .B(n8188), .Z(n406) );
  AND U646 ( .A(n405), .B(n406), .Z(n8317) );
  NANDN U647 ( .A(n8204), .B(n8203), .Z(n407) );
  NANDN U648 ( .A(n8201), .B(n8202), .Z(n408) );
  AND U649 ( .A(n407), .B(n408), .Z(n8247) );
  NANDN U650 ( .A(n8259), .B(n8260), .Z(n409) );
  NANDN U651 ( .A(n8257), .B(n8258), .Z(n410) );
  NAND U652 ( .A(n409), .B(n410), .Z(n8370) );
  NANDN U653 ( .A(n8313), .B(n8314), .Z(n411) );
  NANDN U654 ( .A(n8311), .B(n8312), .Z(n412) );
  NAND U655 ( .A(n411), .B(n412), .Z(n8422) );
  NANDN U656 ( .A(n8374), .B(n8375), .Z(n413) );
  NANDN U657 ( .A(n8377), .B(n8376), .Z(n414) );
  NAND U658 ( .A(n413), .B(n414), .Z(n8509) );
  NANDN U659 ( .A(n8473), .B(n8474), .Z(n415) );
  NANDN U660 ( .A(n8471), .B(n8472), .Z(n416) );
  NAND U661 ( .A(n415), .B(n416), .Z(n8550) );
  NANDN U662 ( .A(n8510), .B(n8511), .Z(n417) );
  NANDN U663 ( .A(n8512), .B(n8513), .Z(n418) );
  AND U664 ( .A(n417), .B(n418), .Z(n8614) );
  NANDN U665 ( .A(n8567), .B(n8568), .Z(n419) );
  NANDN U666 ( .A(n8565), .B(n8566), .Z(n420) );
  NAND U667 ( .A(n419), .B(n420), .Z(n8669) );
  NANDN U668 ( .A(n8591), .B(n8592), .Z(n421) );
  NANDN U669 ( .A(n8593), .B(n8594), .Z(n422) );
  AND U670 ( .A(n421), .B(n422), .Z(n8663) );
  OR U671 ( .A(n8617), .B(n8618), .Z(n423) );
  NANDN U672 ( .A(n8615), .B(n8616), .Z(n424) );
  AND U673 ( .A(n423), .B(n424), .Z(n8679) );
  NANDN U674 ( .A(n8709), .B(n8710), .Z(n425) );
  NANDN U675 ( .A(n8707), .B(n8708), .Z(n426) );
  NAND U676 ( .A(n425), .B(n426), .Z(n8805) );
  NANDN U677 ( .A(n8732), .B(n8733), .Z(n427) );
  NANDN U678 ( .A(n8731), .B(n8811), .Z(n428) );
  AND U679 ( .A(n427), .B(n428), .Z(n8755) );
  NANDN U680 ( .A(n8807), .B(n8808), .Z(n429) );
  NANDN U681 ( .A(n8809), .B(n8810), .Z(n430) );
  AND U682 ( .A(n429), .B(n430), .Z(n8907) );
  NANDN U683 ( .A(n8760), .B(n8761), .Z(n431) );
  NANDN U684 ( .A(n8759), .B(n8758), .Z(n432) );
  AND U685 ( .A(n431), .B(n432), .Z(n8903) );
  NANDN U686 ( .A(n8869), .B(n8868), .Z(n433) );
  NANDN U687 ( .A(n8866), .B(n8867), .Z(n434) );
  AND U688 ( .A(n433), .B(n434), .Z(n9002) );
  NANDN U689 ( .A(n8842), .B(n8843), .Z(n435) );
  NANDN U690 ( .A(n8844), .B(n8845), .Z(n436) );
  AND U691 ( .A(n435), .B(n436), .Z(n8998) );
  NANDN U692 ( .A(n9054), .B(n9055), .Z(n437) );
  NANDN U693 ( .A(n9052), .B(n9053), .Z(n438) );
  NAND U694 ( .A(n437), .B(n438), .Z(n9159) );
  NANDN U695 ( .A(n9116), .B(n9078), .Z(n439) );
  NANDN U696 ( .A(n9080), .B(n9079), .Z(n440) );
  NAND U697 ( .A(n439), .B(n440), .Z(n9157) );
  NANDN U698 ( .A(n9147), .B(n9148), .Z(n441) );
  NANDN U699 ( .A(n9149), .B(n9150), .Z(n442) );
  AND U700 ( .A(n441), .B(n442), .Z(n9241) );
  NANDN U701 ( .A(n9207), .B(n9208), .Z(n443) );
  NANDN U702 ( .A(n9205), .B(n9206), .Z(n444) );
  NAND U703 ( .A(n443), .B(n444), .Z(n9310) );
  NANDN U704 ( .A(n9279), .B(n9280), .Z(n445) );
  NANDN U705 ( .A(n9277), .B(n9278), .Z(n446) );
  NAND U706 ( .A(n445), .B(n446), .Z(n9336) );
  NANDN U707 ( .A(n9300), .B(n9301), .Z(n447) );
  NANDN U708 ( .A(n9302), .B(n9303), .Z(n448) );
  AND U709 ( .A(n447), .B(n448), .Z(n9377) );
  NAND U710 ( .A(n9415), .B(n9416), .Z(n449) );
  NANDN U711 ( .A(n9413), .B(n9414), .Z(n450) );
  AND U712 ( .A(n449), .B(n450), .Z(n9493) );
  NANDN U713 ( .A(n1153), .B(n1154), .Z(n451) );
  NANDN U714 ( .A(n1152), .B(n1151), .Z(n452) );
  NAND U715 ( .A(n451), .B(n452), .Z(n1177) );
  NANDN U716 ( .A(n1595), .B(n1594), .Z(n453) );
  NANDN U717 ( .A(n1592), .B(n1593), .Z(n454) );
  AND U718 ( .A(n453), .B(n454), .Z(n1694) );
  NANDN U719 ( .A(n1707), .B(n1708), .Z(n455) );
  NANDN U720 ( .A(n1706), .B(n1705), .Z(n456) );
  AND U721 ( .A(n455), .B(n456), .Z(n1788) );
  NANDN U722 ( .A(n2020), .B(n2021), .Z(n457) );
  NANDN U723 ( .A(n2019), .B(n2018), .Z(n458) );
  AND U724 ( .A(n457), .B(n458), .Z(n2138) );
  NANDN U725 ( .A(n7600), .B(n7601), .Z(n459) );
  NANDN U726 ( .A(n7598), .B(n7599), .Z(n460) );
  NAND U727 ( .A(n459), .B(n460), .Z(n7730) );
  NANDN U728 ( .A(n7849), .B(n7850), .Z(n461) );
  NANDN U729 ( .A(n7851), .B(n7852), .Z(n462) );
  AND U730 ( .A(n461), .B(n462), .Z(n7967) );
  NANDN U731 ( .A(n7756), .B(n7757), .Z(n463) );
  NANDN U732 ( .A(n7758), .B(n7759), .Z(n464) );
  AND U733 ( .A(n463), .B(n464), .Z(n7865) );
  XOR U734 ( .A(n8089), .B(n8088), .Z(n8091) );
  NANDN U735 ( .A(n9240), .B(n9239), .Z(n465) );
  NANDN U736 ( .A(n9237), .B(n9238), .Z(n466) );
  AND U737 ( .A(n465), .B(n466), .Z(n9258) );
  NAND U738 ( .A(n9283), .B(n9284), .Z(n467) );
  NANDN U739 ( .A(n9281), .B(n9282), .Z(n468) );
  AND U740 ( .A(n467), .B(n468), .Z(n9381) );
  NANDN U741 ( .A(n9444), .B(n9445), .Z(n469) );
  NANDN U742 ( .A(n9446), .B(n9447), .Z(n470) );
  AND U743 ( .A(n469), .B(n470), .Z(n9495) );
  NANDN U744 ( .A(n9465), .B(n9466), .Z(n471) );
  NANDN U745 ( .A(n9464), .B(n9486), .Z(n472) );
  NAND U746 ( .A(n471), .B(n472), .Z(n9559) );
  NANDN U747 ( .A(n9487), .B(n9488), .Z(n473) );
  NANDN U748 ( .A(n9489), .B(n9490), .Z(n474) );
  AND U749 ( .A(n473), .B(n474), .Z(n9518) );
  NANDN U750 ( .A(n9534), .B(n9535), .Z(n475) );
  NANDN U751 ( .A(n9532), .B(n9533), .Z(n476) );
  NAND U752 ( .A(n475), .B(n476), .Z(n9580) );
  NANDN U753 ( .A(n7748), .B(n7749), .Z(n477) );
  NANDN U754 ( .A(n7750), .B(n7751), .Z(n478) );
  AND U755 ( .A(n477), .B(n478), .Z(n7972) );
  NANDN U756 ( .A(n9081), .B(n9082), .Z(n479) );
  NANDN U757 ( .A(n9084), .B(n9083), .Z(n480) );
  NAND U758 ( .A(n479), .B(n480), .Z(n9093) );
  ANDN U759 ( .B(n7951), .A(n609), .Z(n8180) );
  NANDN U760 ( .A(n635), .B(n634), .Z(n481) );
  NANDN U761 ( .A(n632), .B(n633), .Z(n482) );
  AND U762 ( .A(n481), .B(n482), .Z(n666) );
  NANDN U763 ( .A(n8225), .B(n8226), .Z(n483) );
  NANDN U764 ( .A(n8223), .B(n8224), .Z(n484) );
  NAND U765 ( .A(n483), .B(n484), .Z(n8327) );
  NANDN U766 ( .A(n8430), .B(n8431), .Z(n485) );
  NANDN U767 ( .A(n8432), .B(n8433), .Z(n486) );
  AND U768 ( .A(n485), .B(n486), .Z(n8436) );
  NANDN U769 ( .A(n8538), .B(n8539), .Z(n487) );
  NANDN U770 ( .A(n8537), .B(n8536), .Z(n488) );
  AND U771 ( .A(n487), .B(n488), .Z(n8542) );
  NANDN U772 ( .A(n8641), .B(n8642), .Z(n489) );
  NANDN U773 ( .A(n8640), .B(n8639), .Z(n490) );
  AND U774 ( .A(n489), .B(n490), .Z(n8645) );
  NANDN U775 ( .A(n8651), .B(n8652), .Z(n491) );
  NANDN U776 ( .A(n8653), .B(n8654), .Z(n492) );
  AND U777 ( .A(n491), .B(n492), .Z(n8741) );
  NANDN U778 ( .A(n8748), .B(n8749), .Z(n493) );
  NANDN U779 ( .A(n8746), .B(n8747), .Z(n494) );
  NAND U780 ( .A(n493), .B(n494), .Z(n8832) );
  NANDN U781 ( .A(n8914), .B(n8915), .Z(n495) );
  NANDN U782 ( .A(n8913), .B(n8912), .Z(n496) );
  AND U783 ( .A(n495), .B(n496), .Z(n8918) );
  NANDN U784 ( .A(n8924), .B(n8925), .Z(n497) );
  NANDN U785 ( .A(n8926), .B(n8927), .Z(n498) );
  AND U786 ( .A(n497), .B(n498), .Z(n9009) );
  NAND U787 ( .A(n9015), .B(n9014), .Z(n499) );
  NANDN U788 ( .A(n9016), .B(n9017), .Z(n500) );
  NAND U789 ( .A(n499), .B(n500), .Z(n9087) );
  NANDN U790 ( .A(n9179), .B(n9180), .Z(n501) );
  NANDN U791 ( .A(n9178), .B(n9177), .Z(n502) );
  AND U792 ( .A(n501), .B(n502), .Z(n9248) );
  NANDN U793 ( .A(n9458), .B(n9459), .Z(n503) );
  NANDN U794 ( .A(n9456), .B(n9457), .Z(n504) );
  NAND U795 ( .A(n503), .B(n504), .Z(n9507) );
  NANDN U796 ( .A(n9667), .B(n9668), .Z(n505) );
  NANDN U797 ( .A(n9670), .B(n9669), .Z(n506) );
  NAND U798 ( .A(n505), .B(n506), .Z(n9703) );
  NANDN U799 ( .A(n9711), .B(n9712), .Z(n507) );
  NANDN U800 ( .A(n9710), .B(n9709), .Z(n508) );
  AND U801 ( .A(n507), .B(n508), .Z(n9748) );
  NANDN U802 ( .A(n9753), .B(n9754), .Z(n509) );
  NANDN U803 ( .A(n9756), .B(n9755), .Z(n510) );
  NAND U804 ( .A(n509), .B(n510), .Z(n9785) );
  NANDN U805 ( .A(n9814), .B(n9815), .Z(n511) );
  NANDN U806 ( .A(n9816), .B(n9817), .Z(n512) );
  AND U807 ( .A(n511), .B(n512), .Z(n9820) );
  NANDN U808 ( .A(n9841), .B(n9842), .Z(n513) );
  NANDN U809 ( .A(n9839), .B(n9840), .Z(n514) );
  NAND U810 ( .A(n513), .B(n514), .Z(n9845) );
  NAND U811 ( .A(n9857), .B(n9858), .Z(n515) );
  NANDN U812 ( .A(n9855), .B(n9856), .Z(n516) );
  AND U813 ( .A(n515), .B(n516), .Z(n9887) );
  NANDN U814 ( .A(n9866), .B(n9867), .Z(n517) );
  NANDN U815 ( .A(n9868), .B(n9869), .Z(n518) );
  AND U816 ( .A(n517), .B(n518), .Z(n9872) );
  NAND U817 ( .A(n619), .B(n618), .Z(n519) );
  XOR U818 ( .A(n619), .B(n618), .Z(n520) );
  NANDN U819 ( .A(sreg[35]), .B(n520), .Z(n521) );
  NAND U820 ( .A(n519), .B(n521), .Z(n653) );
  NANDN U821 ( .A(n7744), .B(n7745), .Z(n522) );
  NANDN U822 ( .A(n7747), .B(n7746), .Z(n523) );
  NAND U823 ( .A(n522), .B(n523), .Z(n7863) );
  NANDN U824 ( .A(n8102), .B(n8103), .Z(n524) );
  NANDN U825 ( .A(n8105), .B(n8104), .Z(n525) );
  NAND U826 ( .A(n524), .B(n525), .Z(n8219) );
  NANDN U827 ( .A(n9387), .B(n9388), .Z(n526) );
  NANDN U828 ( .A(n9390), .B(n9389), .Z(n527) );
  NAND U829 ( .A(n526), .B(n527), .Z(n9452) );
  NANDN U830 ( .A(n9614), .B(n9615), .Z(n528) );
  NANDN U831 ( .A(n9617), .B(n9616), .Z(n529) );
  NAND U832 ( .A(n528), .B(n529), .Z(n9663) );
  NAND U833 ( .A(n1406), .B(n1407), .Z(n530) );
  XOR U834 ( .A(n1406), .B(n1407), .Z(n531) );
  NAND U835 ( .A(n531), .B(sreg[50]), .Z(n532) );
  NAND U836 ( .A(n530), .B(n532), .Z(n1495) );
  NAND U837 ( .A(n3047), .B(n3046), .Z(n533) );
  XOR U838 ( .A(n3047), .B(n3046), .Z(n534) );
  NANDN U839 ( .A(sreg[64]), .B(n534), .Z(n535) );
  NAND U840 ( .A(n533), .B(n535), .Z(n3338) );
  NAND U841 ( .A(n3487), .B(n3488), .Z(n536) );
  XOR U842 ( .A(n3487), .B(n3488), .Z(n537) );
  NAND U843 ( .A(n537), .B(sreg[67]), .Z(n538) );
  NAND U844 ( .A(n536), .B(n538), .Z(n3779) );
  AND U845 ( .A(n9920), .B(n9921), .Z(n539) );
  NANDN U846 ( .A(n9921), .B(n9917), .Z(n540) );
  NANDN U847 ( .A(n9919), .B(n539), .Z(n541) );
  XNOR U848 ( .A(n539), .B(n9919), .Z(n542) );
  NAND U849 ( .A(n542), .B(n9918), .Z(n543) );
  NAND U850 ( .A(n541), .B(n543), .Z(n544) );
  AND U851 ( .A(n540), .B(n544), .Z(n545) );
  NAND U852 ( .A(n9924), .B(n9925), .Z(n546) );
  NAND U853 ( .A(n9922), .B(n9923), .Z(n547) );
  AND U854 ( .A(n546), .B(n547), .Z(n548) );
  XNOR U855 ( .A(a[62]), .B(a[63]), .Z(n549) );
  XNOR U856 ( .A(n9926), .B(n549), .Z(n550) );
  NAND U857 ( .A(n550), .B(b[31]), .Z(n551) );
  XNOR U858 ( .A(n545), .B(n548), .Z(n552) );
  XNOR U859 ( .A(n551), .B(n552), .Z(c[127]) );
  NAND U860 ( .A(n1080), .B(n8853), .Z(n553) );
  NAND U861 ( .A(n1340), .B(n9195), .Z(n554) );
  XNOR U862 ( .A(b[18]), .B(b[17]), .Z(n555) );
  NAND U863 ( .A(n1753), .B(n9480), .Z(n556) );
  NAND U864 ( .A(n1209), .B(n9067), .Z(n557) );
  NAND U865 ( .A(n747), .B(n8290), .Z(n558) );
  NAND U866 ( .A(n2702), .B(n9796), .Z(n559) );
  NAND U867 ( .A(n623), .B(n7784), .Z(n560) );
  NAND U868 ( .A(n675), .B(n8041), .Z(n561) );
  NAND U869 ( .A(n945), .B(n8701), .Z(n562) );
  NAND U870 ( .A(n1978), .B(n9605), .Z(n563) );
  NAND U871 ( .A(n840), .B(n8485), .Z(n564) );
  NAND U872 ( .A(n2467), .B(n9692), .Z(n565) );
  NAND U873 ( .A(n2158), .B(n9684), .Z(n566) );
  IV U874 ( .A(n561), .Z(n567) );
  IV U875 ( .A(n560), .Z(n568) );
  IV U876 ( .A(n558), .Z(n569) );
  IV U877 ( .A(n564), .Z(n570) );
  IV U878 ( .A(n562), .Z(n571) );
  IV U879 ( .A(n553), .Z(n572) );
  IV U880 ( .A(n557), .Z(n573) );
  IV U881 ( .A(n9046), .Z(n574) );
  IV U882 ( .A(n555), .Z(n575) );
  IV U883 ( .A(n554), .Z(n576) );
  IV U884 ( .A(n556), .Z(n577) );
  IV U885 ( .A(n563), .Z(n578) );
  IV U886 ( .A(n566), .Z(n579) );
  IV U887 ( .A(n9764), .Z(n580) );
  IV U888 ( .A(n9796), .Z(n581) );
  IV U889 ( .A(n565), .Z(n582) );
  IV U890 ( .A(n559), .Z(n583) );
  IV U891 ( .A(n9904), .Z(n584) );
  AND U892 ( .A(b[0]), .B(a[0]), .Z(n585) );
  XOR U893 ( .A(n585), .B(sreg[32]), .Z(c[32]) );
  AND U894 ( .A(b[1]), .B(a[0]), .Z(n603) );
  NAND U895 ( .A(b[0]), .B(a[1]), .Z(n592) );
  XOR U896 ( .A(n603), .B(n592), .Z(n586) );
  XNOR U897 ( .A(sreg[33]), .B(n586), .Z(n588) );
  AND U898 ( .A(n585), .B(sreg[32]), .Z(n587) );
  XOR U899 ( .A(n588), .B(n587), .Z(c[33]) );
  NANDN U900 ( .A(n586), .B(sreg[33]), .Z(n590) );
  NAND U901 ( .A(n588), .B(n587), .Z(n589) );
  AND U902 ( .A(n590), .B(n589), .Z(n612) );
  XNOR U903 ( .A(n612), .B(sreg[34]), .Z(n614) );
  NAND U904 ( .A(a[0]), .B(b[2]), .Z(n591) );
  XNOR U905 ( .A(b[1]), .B(n591), .Z(n594) );
  OR U906 ( .A(a[0]), .B(n592), .Z(n593) );
  NAND U907 ( .A(n594), .B(n593), .Z(n599) );
  AND U908 ( .A(b[0]), .B(a[2]), .Z(n595) );
  XOR U909 ( .A(b[1]), .B(n595), .Z(n597) );
  NANDN U910 ( .A(b[0]), .B(a[1]), .Z(n596) );
  AND U911 ( .A(n597), .B(n596), .Z(n598) );
  XNOR U912 ( .A(n599), .B(n598), .Z(n613) );
  XOR U913 ( .A(n614), .B(n613), .Z(c[34]) );
  NANDN U914 ( .A(n599), .B(n598), .Z(n622) );
  NAND U915 ( .A(b[0]), .B(a[3]), .Z(n600) );
  XNOR U916 ( .A(b[1]), .B(n600), .Z(n602) );
  NANDN U917 ( .A(b[0]), .B(a[2]), .Z(n601) );
  NAND U918 ( .A(n602), .B(n601), .Z(n630) );
  XNOR U919 ( .A(b[2]), .B(b[1]), .Z(n7784) );
  IV U920 ( .A(n7784), .Z(n7245) );
  XOR U921 ( .A(b[3]), .B(a[1]), .Z(n624) );
  NAND U922 ( .A(n7245), .B(n624), .Z(n608) );
  ANDN U923 ( .B(b[3]), .A(b[2]), .Z(n609) );
  OR U924 ( .A(n603), .B(n609), .Z(n605) );
  NAND U925 ( .A(a[0]), .B(b[3]), .Z(n604) );
  AND U926 ( .A(n605), .B(n604), .Z(n606) );
  NANDN U927 ( .A(n7245), .B(n606), .Z(n607) );
  AND U928 ( .A(n608), .B(n607), .Z(n631) );
  XNOR U929 ( .A(n630), .B(n631), .Z(n621) );
  NAND U930 ( .A(n7245), .B(a[0]), .Z(n610) );
  NAND U931 ( .A(n7245), .B(b[3]), .Z(n7951) );
  ANDN U932 ( .B(n610), .A(n8180), .Z(n620) );
  XOR U933 ( .A(n621), .B(n620), .Z(n611) );
  XNOR U934 ( .A(n622), .B(n611), .Z(n618) );
  NANDN U935 ( .A(n612), .B(sreg[34]), .Z(n616) );
  NAND U936 ( .A(n614), .B(n613), .Z(n615) );
  AND U937 ( .A(n616), .B(n615), .Z(n619) );
  XNOR U938 ( .A(sreg[35]), .B(n619), .Z(n617) );
  XNOR U939 ( .A(n618), .B(n617), .Z(c[35]) );
  XNOR U940 ( .A(n653), .B(sreg[36]), .Z(n655) );
  XOR U941 ( .A(b[2]), .B(b[3]), .Z(n623) );
  NAND U942 ( .A(n568), .B(n624), .Z(n626) );
  XOR U943 ( .A(b[3]), .B(a[2]), .Z(n636) );
  NAND U944 ( .A(n7245), .B(n636), .Z(n625) );
  AND U945 ( .A(n626), .B(n625), .Z(n650) );
  XNOR U946 ( .A(b[4]), .B(b[3]), .Z(n8041) );
  IV U947 ( .A(n8041), .Z(n7235) );
  AND U948 ( .A(a[0]), .B(n7235), .Z(n647) );
  NAND U949 ( .A(b[0]), .B(a[4]), .Z(n627) );
  XNOR U950 ( .A(b[1]), .B(n627), .Z(n629) );
  NANDN U951 ( .A(b[0]), .B(a[3]), .Z(n628) );
  NAND U952 ( .A(n629), .B(n628), .Z(n648) );
  XNOR U953 ( .A(n647), .B(n648), .Z(n649) );
  XNOR U954 ( .A(n650), .B(n649), .Z(n633) );
  OR U955 ( .A(n631), .B(n630), .Z(n632) );
  XNOR U956 ( .A(n633), .B(n632), .Z(n634) );
  XNOR U957 ( .A(n635), .B(n634), .Z(n654) );
  XOR U958 ( .A(n655), .B(n654), .Z(c[36]) );
  NAND U959 ( .A(n568), .B(n636), .Z(n638) );
  XOR U960 ( .A(b[3]), .B(a[3]), .Z(n669) );
  NAND U961 ( .A(n7245), .B(n669), .Z(n637) );
  AND U962 ( .A(n638), .B(n637), .Z(n682) );
  NANDN U963 ( .A(b[4]), .B(b[5]), .Z(n639) );
  NAND U964 ( .A(n7235), .B(b[5]), .Z(n8165) );
  NAND U965 ( .A(n639), .B(n8165), .Z(n8365) );
  ANDN U966 ( .B(n8365), .A(n647), .Z(n681) );
  XNOR U967 ( .A(n682), .B(n681), .Z(n684) );
  NAND U968 ( .A(b[0]), .B(a[5]), .Z(n640) );
  XNOR U969 ( .A(b[1]), .B(n640), .Z(n642) );
  NANDN U970 ( .A(b[0]), .B(a[4]), .Z(n641) );
  NAND U971 ( .A(n642), .B(n641), .Z(n679) );
  XOR U972 ( .A(b[5]), .B(b[4]), .Z(n675) );
  XOR U973 ( .A(b[5]), .B(a[0]), .Z(n643) );
  NAND U974 ( .A(n675), .B(n643), .Z(n644) );
  NANDN U975 ( .A(n644), .B(n8041), .Z(n646) );
  XOR U976 ( .A(b[5]), .B(a[1]), .Z(n676) );
  NANDN U977 ( .A(n8041), .B(n676), .Z(n645) );
  NAND U978 ( .A(n646), .B(n645), .Z(n680) );
  XNOR U979 ( .A(n679), .B(n680), .Z(n683) );
  XOR U980 ( .A(n684), .B(n683), .Z(n664) );
  NANDN U981 ( .A(n648), .B(n647), .Z(n652) );
  NANDN U982 ( .A(n650), .B(n649), .Z(n651) );
  AND U983 ( .A(n652), .B(n651), .Z(n663) );
  XNOR U984 ( .A(n664), .B(n663), .Z(n665) );
  XOR U985 ( .A(n666), .B(n665), .Z(n658) );
  XNOR U986 ( .A(n658), .B(sreg[37]), .Z(n660) );
  NANDN U987 ( .A(n653), .B(sreg[36]), .Z(n657) );
  NAND U988 ( .A(n655), .B(n654), .Z(n656) );
  NAND U989 ( .A(n657), .B(n656), .Z(n659) );
  XOR U990 ( .A(n660), .B(n659), .Z(c[37]) );
  NANDN U991 ( .A(n658), .B(sreg[37]), .Z(n662) );
  NAND U992 ( .A(n660), .B(n659), .Z(n661) );
  AND U993 ( .A(n662), .B(n661), .Z(n719) );
  XNOR U994 ( .A(n719), .B(sreg[38]), .Z(n721) );
  NANDN U995 ( .A(n664), .B(n663), .Z(n668) );
  NAND U996 ( .A(n666), .B(n665), .Z(n667) );
  AND U997 ( .A(n668), .B(n667), .Z(n689) );
  NAND U998 ( .A(n568), .B(n669), .Z(n671) );
  XOR U999 ( .A(b[3]), .B(a[4]), .Z(n704) );
  NAND U1000 ( .A(n7245), .B(n704), .Z(n670) );
  AND U1001 ( .A(n671), .B(n670), .Z(n710) );
  XNOR U1002 ( .A(b[6]), .B(b[5]), .Z(n8290) );
  IV U1003 ( .A(n8290), .Z(n7819) );
  AND U1004 ( .A(a[0]), .B(n7819), .Z(n707) );
  NAND U1005 ( .A(b[0]), .B(a[6]), .Z(n672) );
  XNOR U1006 ( .A(b[1]), .B(n672), .Z(n674) );
  NANDN U1007 ( .A(b[0]), .B(a[5]), .Z(n673) );
  NAND U1008 ( .A(n674), .B(n673), .Z(n708) );
  XNOR U1009 ( .A(n707), .B(n708), .Z(n709) );
  XNOR U1010 ( .A(n710), .B(n709), .Z(n716) );
  NAND U1011 ( .A(n567), .B(n676), .Z(n678) );
  XOR U1012 ( .A(b[5]), .B(a[2]), .Z(n693) );
  NAND U1013 ( .A(n7235), .B(n693), .Z(n677) );
  AND U1014 ( .A(n678), .B(n677), .Z(n714) );
  ANDN U1015 ( .B(n680), .A(n679), .Z(n713) );
  XNOR U1016 ( .A(n714), .B(n713), .Z(n715) );
  XOR U1017 ( .A(n716), .B(n715), .Z(n688) );
  NANDN U1018 ( .A(n682), .B(n681), .Z(n686) );
  NAND U1019 ( .A(n684), .B(n683), .Z(n685) );
  AND U1020 ( .A(n686), .B(n685), .Z(n687) );
  XOR U1021 ( .A(n688), .B(n687), .Z(n690) );
  XNOR U1022 ( .A(n689), .B(n690), .Z(n720) );
  XOR U1023 ( .A(n721), .B(n720), .Z(c[38]) );
  NANDN U1024 ( .A(n688), .B(n687), .Z(n692) );
  OR U1025 ( .A(n690), .B(n689), .Z(n691) );
  AND U1026 ( .A(n692), .B(n691), .Z(n731) );
  NAND U1027 ( .A(n567), .B(n693), .Z(n695) );
  XOR U1028 ( .A(b[5]), .B(a[3]), .Z(n759) );
  NAND U1029 ( .A(n7235), .B(n759), .Z(n694) );
  AND U1030 ( .A(n695), .B(n694), .Z(n754) );
  XOR U1031 ( .A(b[7]), .B(b[6]), .Z(n747) );
  XOR U1032 ( .A(b[7]), .B(a[0]), .Z(n696) );
  NAND U1033 ( .A(n747), .B(n696), .Z(n697) );
  NANDN U1034 ( .A(n697), .B(n8290), .Z(n699) );
  XOR U1035 ( .A(b[7]), .B(a[1]), .Z(n748) );
  NANDN U1036 ( .A(n8290), .B(n748), .Z(n698) );
  AND U1037 ( .A(n699), .B(n698), .Z(n755) );
  XOR U1038 ( .A(n754), .B(n755), .Z(n744) );
  NANDN U1039 ( .A(b[6]), .B(b[7]), .Z(n700) );
  NAND U1040 ( .A(n7819), .B(b[7]), .Z(n8413) );
  NAND U1041 ( .A(n700), .B(n8413), .Z(n8491) );
  ANDN U1042 ( .B(n8491), .A(n707), .Z(n742) );
  NAND U1043 ( .A(b[0]), .B(a[7]), .Z(n701) );
  XNOR U1044 ( .A(b[1]), .B(n701), .Z(n703) );
  NANDN U1045 ( .A(b[0]), .B(a[6]), .Z(n702) );
  NAND U1046 ( .A(n703), .B(n702), .Z(n741) );
  XNOR U1047 ( .A(n742), .B(n741), .Z(n743) );
  XNOR U1048 ( .A(n744), .B(n743), .Z(n735) );
  NANDN U1049 ( .A(n560), .B(n704), .Z(n706) );
  XNOR U1050 ( .A(b[3]), .B(a[5]), .Z(n751) );
  OR U1051 ( .A(n751), .B(n7784), .Z(n705) );
  NAND U1052 ( .A(n706), .B(n705), .Z(n736) );
  XNOR U1053 ( .A(n735), .B(n736), .Z(n737) );
  NANDN U1054 ( .A(n708), .B(n707), .Z(n712) );
  NANDN U1055 ( .A(n710), .B(n709), .Z(n711) );
  NAND U1056 ( .A(n712), .B(n711), .Z(n738) );
  XNOR U1057 ( .A(n737), .B(n738), .Z(n729) );
  NANDN U1058 ( .A(n714), .B(n713), .Z(n718) );
  NAND U1059 ( .A(n716), .B(n715), .Z(n717) );
  NAND U1060 ( .A(n718), .B(n717), .Z(n730) );
  XOR U1061 ( .A(n729), .B(n730), .Z(n732) );
  XOR U1062 ( .A(n731), .B(n732), .Z(n724) );
  XNOR U1063 ( .A(n724), .B(sreg[39]), .Z(n726) );
  NANDN U1064 ( .A(n719), .B(sreg[38]), .Z(n723) );
  NAND U1065 ( .A(n721), .B(n720), .Z(n722) );
  NAND U1066 ( .A(n723), .B(n722), .Z(n725) );
  XOR U1067 ( .A(n726), .B(n725), .Z(c[39]) );
  NANDN U1068 ( .A(n724), .B(sreg[39]), .Z(n728) );
  NAND U1069 ( .A(n726), .B(n725), .Z(n727) );
  AND U1070 ( .A(n728), .B(n727), .Z(n803) );
  XNOR U1071 ( .A(n803), .B(sreg[40]), .Z(n805) );
  NANDN U1072 ( .A(n730), .B(n729), .Z(n734) );
  OR U1073 ( .A(n732), .B(n731), .Z(n733) );
  AND U1074 ( .A(n734), .B(n733), .Z(n799) );
  NANDN U1075 ( .A(n736), .B(n735), .Z(n740) );
  NANDN U1076 ( .A(n738), .B(n737), .Z(n739) );
  AND U1077 ( .A(n740), .B(n739), .Z(n798) );
  NANDN U1078 ( .A(n742), .B(n741), .Z(n746) );
  NANDN U1079 ( .A(n744), .B(n743), .Z(n745) );
  AND U1080 ( .A(n746), .B(n745), .Z(n765) );
  NAND U1081 ( .A(n569), .B(n748), .Z(n750) );
  XOR U1082 ( .A(b[7]), .B(a[2]), .Z(n779) );
  NAND U1083 ( .A(n7819), .B(n779), .Z(n749) );
  AND U1084 ( .A(n750), .B(n749), .Z(n769) );
  OR U1085 ( .A(n751), .B(n560), .Z(n753) );
  XOR U1086 ( .A(b[3]), .B(a[6]), .Z(n794) );
  NAND U1087 ( .A(n7245), .B(n794), .Z(n752) );
  NAND U1088 ( .A(n753), .B(n752), .Z(n768) );
  XNOR U1089 ( .A(n769), .B(n768), .Z(n771) );
  NOR U1090 ( .A(n755), .B(n754), .Z(n770) );
  XOR U1091 ( .A(n771), .B(n770), .Z(n763) );
  NAND U1092 ( .A(b[0]), .B(a[8]), .Z(n756) );
  XNOR U1093 ( .A(b[1]), .B(n756), .Z(n758) );
  NANDN U1094 ( .A(b[0]), .B(a[7]), .Z(n757) );
  NAND U1095 ( .A(n758), .B(n757), .Z(n776) );
  XNOR U1096 ( .A(b[8]), .B(b[7]), .Z(n8485) );
  IV U1097 ( .A(n8485), .Z(n8037) );
  AND U1098 ( .A(a[0]), .B(n8037), .Z(n787) );
  NAND U1099 ( .A(n567), .B(n759), .Z(n761) );
  XOR U1100 ( .A(b[5]), .B(a[4]), .Z(n788) );
  NAND U1101 ( .A(n7235), .B(n788), .Z(n760) );
  AND U1102 ( .A(n761), .B(n760), .Z(n774) );
  XOR U1103 ( .A(n787), .B(n774), .Z(n775) );
  XNOR U1104 ( .A(n776), .B(n775), .Z(n762) );
  XNOR U1105 ( .A(n763), .B(n762), .Z(n764) );
  XNOR U1106 ( .A(n765), .B(n764), .Z(n797) );
  XOR U1107 ( .A(n798), .B(n797), .Z(n800) );
  XNOR U1108 ( .A(n799), .B(n800), .Z(n804) );
  XOR U1109 ( .A(n805), .B(n804), .Z(c[40]) );
  NANDN U1110 ( .A(n763), .B(n762), .Z(n767) );
  NANDN U1111 ( .A(n765), .B(n764), .Z(n766) );
  AND U1112 ( .A(n767), .B(n766), .Z(n813) );
  NANDN U1113 ( .A(n769), .B(n768), .Z(n773) );
  NAND U1114 ( .A(n771), .B(n770), .Z(n772) );
  AND U1115 ( .A(n773), .B(n772), .Z(n852) );
  NANDN U1116 ( .A(n774), .B(n787), .Z(n778) );
  OR U1117 ( .A(n776), .B(n775), .Z(n777) );
  AND U1118 ( .A(n778), .B(n777), .Z(n850) );
  NAND U1119 ( .A(n569), .B(n779), .Z(n781) );
  XOR U1120 ( .A(b[7]), .B(a[3]), .Z(n834) );
  NAND U1121 ( .A(n7819), .B(n834), .Z(n780) );
  AND U1122 ( .A(n781), .B(n780), .Z(n844) );
  XOR U1123 ( .A(b[9]), .B(b[8]), .Z(n840) );
  XOR U1124 ( .A(b[9]), .B(a[0]), .Z(n782) );
  NAND U1125 ( .A(n840), .B(n782), .Z(n783) );
  NANDN U1126 ( .A(n783), .B(n8485), .Z(n785) );
  XOR U1127 ( .A(b[9]), .B(a[1]), .Z(n841) );
  NANDN U1128 ( .A(n8485), .B(n841), .Z(n784) );
  NAND U1129 ( .A(n785), .B(n784), .Z(n845) );
  XOR U1130 ( .A(n844), .B(n845), .Z(n821) );
  NANDN U1131 ( .A(b[8]), .B(b[9]), .Z(n786) );
  NAND U1132 ( .A(n8037), .B(b[9]), .Z(n8604) );
  NAND U1133 ( .A(n786), .B(n8604), .Z(n8726) );
  ANDN U1134 ( .B(n8726), .A(n787), .Z(n820) );
  NAND U1135 ( .A(n567), .B(n788), .Z(n790) );
  XOR U1136 ( .A(b[5]), .B(a[5]), .Z(n837) );
  NAND U1137 ( .A(n7235), .B(n837), .Z(n789) );
  AND U1138 ( .A(n790), .B(n789), .Z(n819) );
  XOR U1139 ( .A(n820), .B(n819), .Z(n822) );
  XOR U1140 ( .A(n821), .B(n822), .Z(n828) );
  NAND U1141 ( .A(b[0]), .B(a[9]), .Z(n791) );
  XNOR U1142 ( .A(b[1]), .B(n791), .Z(n793) );
  NANDN U1143 ( .A(b[0]), .B(a[8]), .Z(n792) );
  NAND U1144 ( .A(n793), .B(n792), .Z(n826) );
  NAND U1145 ( .A(n568), .B(n794), .Z(n796) );
  XOR U1146 ( .A(b[3]), .B(a[7]), .Z(n846) );
  NAND U1147 ( .A(n7245), .B(n846), .Z(n795) );
  NAND U1148 ( .A(n796), .B(n795), .Z(n825) );
  XNOR U1149 ( .A(n826), .B(n825), .Z(n827) );
  XOR U1150 ( .A(n828), .B(n827), .Z(n849) );
  XNOR U1151 ( .A(n850), .B(n849), .Z(n851) );
  XOR U1152 ( .A(n852), .B(n851), .Z(n814) );
  XNOR U1153 ( .A(n813), .B(n814), .Z(n815) );
  NANDN U1154 ( .A(n798), .B(n797), .Z(n802) );
  OR U1155 ( .A(n800), .B(n799), .Z(n801) );
  NAND U1156 ( .A(n802), .B(n801), .Z(n816) );
  XOR U1157 ( .A(n815), .B(n816), .Z(n808) );
  XNOR U1158 ( .A(sreg[41]), .B(n808), .Z(n810) );
  NANDN U1159 ( .A(n803), .B(sreg[40]), .Z(n807) );
  NAND U1160 ( .A(n805), .B(n804), .Z(n806) );
  NAND U1161 ( .A(n807), .B(n806), .Z(n809) );
  XOR U1162 ( .A(n810), .B(n809), .Z(c[41]) );
  NANDN U1163 ( .A(n808), .B(sreg[41]), .Z(n812) );
  NAND U1164 ( .A(n810), .B(n809), .Z(n811) );
  AND U1165 ( .A(n812), .B(n811), .Z(n855) );
  XNOR U1166 ( .A(n855), .B(sreg[42]), .Z(n857) );
  NANDN U1167 ( .A(n814), .B(n813), .Z(n818) );
  NANDN U1168 ( .A(n816), .B(n815), .Z(n817) );
  AND U1169 ( .A(n818), .B(n817), .Z(n863) );
  NANDN U1170 ( .A(n820), .B(n819), .Z(n824) );
  NANDN U1171 ( .A(n822), .B(n821), .Z(n823) );
  AND U1172 ( .A(n824), .B(n823), .Z(n905) );
  NANDN U1173 ( .A(n826), .B(n825), .Z(n830) );
  NAND U1174 ( .A(n828), .B(n827), .Z(n829) );
  AND U1175 ( .A(n830), .B(n829), .Z(n904) );
  XNOR U1176 ( .A(n905), .B(n904), .Z(n906) );
  NAND U1177 ( .A(b[0]), .B(a[10]), .Z(n831) );
  XNOR U1178 ( .A(b[1]), .B(n831), .Z(n833) );
  NANDN U1179 ( .A(b[0]), .B(a[9]), .Z(n832) );
  NAND U1180 ( .A(n833), .B(n832), .Z(n874) );
  XNOR U1181 ( .A(b[10]), .B(b[9]), .Z(n8701) );
  IV U1182 ( .A(n8701), .Z(n8135) );
  AND U1183 ( .A(a[0]), .B(n8135), .Z(n897) );
  NAND U1184 ( .A(n569), .B(n834), .Z(n836) );
  XOR U1185 ( .A(b[7]), .B(a[4]), .Z(n898) );
  NAND U1186 ( .A(n7819), .B(n898), .Z(n835) );
  AND U1187 ( .A(n836), .B(n835), .Z(n872) );
  XOR U1188 ( .A(n897), .B(n872), .Z(n873) );
  XOR U1189 ( .A(n874), .B(n873), .Z(n869) );
  NAND U1190 ( .A(n567), .B(n837), .Z(n839) );
  XOR U1191 ( .A(b[5]), .B(a[6]), .Z(n893) );
  NAND U1192 ( .A(n7235), .B(n893), .Z(n838) );
  AND U1193 ( .A(n839), .B(n838), .Z(n878) );
  NAND U1194 ( .A(n570), .B(n841), .Z(n843) );
  XOR U1195 ( .A(b[9]), .B(a[2]), .Z(n887) );
  NAND U1196 ( .A(n8037), .B(n887), .Z(n842) );
  NAND U1197 ( .A(n843), .B(n842), .Z(n877) );
  XNOR U1198 ( .A(n878), .B(n877), .Z(n880) );
  ANDN U1199 ( .B(n845), .A(n844), .Z(n879) );
  XOR U1200 ( .A(n880), .B(n879), .Z(n867) );
  NANDN U1201 ( .A(n560), .B(n846), .Z(n848) );
  XNOR U1202 ( .A(b[3]), .B(a[8]), .Z(n901) );
  OR U1203 ( .A(n901), .B(n7784), .Z(n847) );
  AND U1204 ( .A(n848), .B(n847), .Z(n866) );
  XNOR U1205 ( .A(n867), .B(n866), .Z(n868) );
  XOR U1206 ( .A(n869), .B(n868), .Z(n907) );
  XNOR U1207 ( .A(n906), .B(n907), .Z(n860) );
  NANDN U1208 ( .A(n850), .B(n849), .Z(n854) );
  NANDN U1209 ( .A(n852), .B(n851), .Z(n853) );
  NAND U1210 ( .A(n854), .B(n853), .Z(n861) );
  XNOR U1211 ( .A(n860), .B(n861), .Z(n862) );
  XNOR U1212 ( .A(n863), .B(n862), .Z(n856) );
  XOR U1213 ( .A(n857), .B(n856), .Z(c[42]) );
  NANDN U1214 ( .A(n855), .B(sreg[42]), .Z(n859) );
  NAND U1215 ( .A(n857), .B(n856), .Z(n858) );
  AND U1216 ( .A(n859), .B(n858), .Z(n912) );
  NANDN U1217 ( .A(n861), .B(n860), .Z(n865) );
  NAND U1218 ( .A(n863), .B(n862), .Z(n864) );
  AND U1219 ( .A(n865), .B(n864), .Z(n918) );
  NANDN U1220 ( .A(n867), .B(n866), .Z(n871) );
  NANDN U1221 ( .A(n869), .B(n868), .Z(n870) );
  AND U1222 ( .A(n871), .B(n870), .Z(n963) );
  NANDN U1223 ( .A(n872), .B(n897), .Z(n876) );
  OR U1224 ( .A(n874), .B(n873), .Z(n875) );
  AND U1225 ( .A(n876), .B(n875), .Z(n961) );
  NANDN U1226 ( .A(n878), .B(n877), .Z(n882) );
  NAND U1227 ( .A(n880), .B(n879), .Z(n881) );
  AND U1228 ( .A(n882), .B(n881), .Z(n924) );
  XOR U1229 ( .A(b[11]), .B(b[10]), .Z(n945) );
  XOR U1230 ( .A(b[11]), .B(a[0]), .Z(n883) );
  NAND U1231 ( .A(n945), .B(n883), .Z(n884) );
  NANDN U1232 ( .A(n884), .B(n8701), .Z(n886) );
  XOR U1233 ( .A(b[11]), .B(a[1]), .Z(n946) );
  NANDN U1234 ( .A(n8701), .B(n946), .Z(n885) );
  AND U1235 ( .A(n886), .B(n885), .Z(n953) );
  NAND U1236 ( .A(n570), .B(n887), .Z(n889) );
  XOR U1237 ( .A(b[9]), .B(a[3]), .Z(n936) );
  NAND U1238 ( .A(n8037), .B(n936), .Z(n888) );
  AND U1239 ( .A(n889), .B(n888), .Z(n952) );
  XOR U1240 ( .A(n953), .B(n952), .Z(n941) );
  NAND U1241 ( .A(b[0]), .B(a[11]), .Z(n890) );
  XNOR U1242 ( .A(b[1]), .B(n890), .Z(n892) );
  NANDN U1243 ( .A(b[0]), .B(a[10]), .Z(n891) );
  NAND U1244 ( .A(n892), .B(n891), .Z(n939) );
  NANDN U1245 ( .A(n561), .B(n893), .Z(n895) );
  XNOR U1246 ( .A(b[5]), .B(a[7]), .Z(n949) );
  OR U1247 ( .A(n949), .B(n8041), .Z(n894) );
  NAND U1248 ( .A(n895), .B(n894), .Z(n940) );
  XOR U1249 ( .A(n939), .B(n940), .Z(n942) );
  XOR U1250 ( .A(n941), .B(n942), .Z(n922) );
  NANDN U1251 ( .A(b[10]), .B(b[11]), .Z(n896) );
  NAND U1252 ( .A(n8135), .B(b[11]), .Z(n8798) );
  NAND U1253 ( .A(n896), .B(n8798), .Z(n8865) );
  IV U1254 ( .A(n8865), .Z(n8941) );
  NOR U1255 ( .A(n8941), .B(n897), .Z(n928) );
  NANDN U1256 ( .A(n558), .B(n898), .Z(n900) );
  XNOR U1257 ( .A(b[7]), .B(a[5]), .Z(n957) );
  OR U1258 ( .A(n957), .B(n8290), .Z(n899) );
  NAND U1259 ( .A(n900), .B(n899), .Z(n927) );
  XOR U1260 ( .A(n928), .B(n927), .Z(n930) );
  OR U1261 ( .A(n901), .B(n560), .Z(n903) );
  XNOR U1262 ( .A(b[3]), .B(a[9]), .Z(n954) );
  OR U1263 ( .A(n954), .B(n7784), .Z(n902) );
  NAND U1264 ( .A(n903), .B(n902), .Z(n929) );
  XOR U1265 ( .A(n930), .B(n929), .Z(n921) );
  XNOR U1266 ( .A(n922), .B(n921), .Z(n923) );
  XNOR U1267 ( .A(n924), .B(n923), .Z(n960) );
  XNOR U1268 ( .A(n961), .B(n960), .Z(n962) );
  XOR U1269 ( .A(n963), .B(n962), .Z(n916) );
  NANDN U1270 ( .A(n905), .B(n904), .Z(n909) );
  NANDN U1271 ( .A(n907), .B(n906), .Z(n908) );
  NAND U1272 ( .A(n909), .B(n908), .Z(n915) );
  XNOR U1273 ( .A(n916), .B(n915), .Z(n917) );
  XNOR U1274 ( .A(n918), .B(n917), .Z(n910) );
  XNOR U1275 ( .A(sreg[43]), .B(n910), .Z(n911) );
  XNOR U1276 ( .A(n912), .B(n911), .Z(c[43]) );
  NANDN U1277 ( .A(sreg[43]), .B(n910), .Z(n914) );
  NAND U1278 ( .A(n912), .B(n911), .Z(n913) );
  NAND U1279 ( .A(n914), .B(n913), .Z(n1025) );
  XNOR U1280 ( .A(sreg[44]), .B(n1025), .Z(n1027) );
  NANDN U1281 ( .A(n916), .B(n915), .Z(n920) );
  NANDN U1282 ( .A(n918), .B(n917), .Z(n919) );
  AND U1283 ( .A(n920), .B(n919), .Z(n968) );
  NANDN U1284 ( .A(n922), .B(n921), .Z(n926) );
  NANDN U1285 ( .A(n924), .B(n923), .Z(n925) );
  AND U1286 ( .A(n926), .B(n925), .Z(n1020) );
  NAND U1287 ( .A(n928), .B(n927), .Z(n932) );
  NAND U1288 ( .A(n930), .B(n929), .Z(n931) );
  NAND U1289 ( .A(n932), .B(n931), .Z(n1019) );
  XNOR U1290 ( .A(n1020), .B(n1019), .Z(n1022) );
  NAND U1291 ( .A(b[0]), .B(a[12]), .Z(n933) );
  XNOR U1292 ( .A(b[1]), .B(n933), .Z(n935) );
  NANDN U1293 ( .A(b[0]), .B(a[11]), .Z(n934) );
  NAND U1294 ( .A(n935), .B(n934), .Z(n1010) );
  XNOR U1295 ( .A(b[12]), .B(b[11]), .Z(n8853) );
  IV U1296 ( .A(n8853), .Z(n8585) );
  AND U1297 ( .A(a[0]), .B(n8585), .Z(n1007) );
  NAND U1298 ( .A(n570), .B(n936), .Z(n938) );
  XOR U1299 ( .A(b[9]), .B(a[4]), .Z(n1000) );
  NAND U1300 ( .A(n8037), .B(n1000), .Z(n937) );
  AND U1301 ( .A(n938), .B(n937), .Z(n1008) );
  XNOR U1302 ( .A(n1007), .B(n1008), .Z(n1009) );
  XNOR U1303 ( .A(n1010), .B(n1009), .Z(n972) );
  NANDN U1304 ( .A(n940), .B(n939), .Z(n944) );
  OR U1305 ( .A(n942), .B(n941), .Z(n943) );
  NAND U1306 ( .A(n944), .B(n943), .Z(n973) );
  XNOR U1307 ( .A(n972), .B(n973), .Z(n974) );
  NAND U1308 ( .A(n571), .B(n946), .Z(n948) );
  XOR U1309 ( .A(b[11]), .B(a[2]), .Z(n990) );
  NAND U1310 ( .A(n8135), .B(n990), .Z(n947) );
  AND U1311 ( .A(n948), .B(n947), .Z(n981) );
  OR U1312 ( .A(n949), .B(n561), .Z(n951) );
  XOR U1313 ( .A(b[5]), .B(a[8]), .Z(n1004) );
  NAND U1314 ( .A(n7235), .B(n1004), .Z(n950) );
  AND U1315 ( .A(n951), .B(n950), .Z(n979) );
  NOR U1316 ( .A(n953), .B(n952), .Z(n1015) );
  OR U1317 ( .A(n954), .B(n560), .Z(n956) );
  XNOR U1318 ( .A(b[3]), .B(a[10]), .Z(n997) );
  OR U1319 ( .A(n997), .B(n7784), .Z(n955) );
  AND U1320 ( .A(n956), .B(n955), .Z(n1013) );
  OR U1321 ( .A(n957), .B(n558), .Z(n959) );
  XNOR U1322 ( .A(b[7]), .B(a[6]), .Z(n987) );
  OR U1323 ( .A(n987), .B(n8290), .Z(n958) );
  NAND U1324 ( .A(n959), .B(n958), .Z(n1014) );
  XOR U1325 ( .A(n1013), .B(n1014), .Z(n1016) );
  XNOR U1326 ( .A(n1015), .B(n1016), .Z(n978) );
  XNOR U1327 ( .A(n979), .B(n978), .Z(n980) );
  XOR U1328 ( .A(n981), .B(n980), .Z(n975) );
  XNOR U1329 ( .A(n974), .B(n975), .Z(n1021) );
  XOR U1330 ( .A(n1022), .B(n1021), .Z(n967) );
  NANDN U1331 ( .A(n961), .B(n960), .Z(n965) );
  NAND U1332 ( .A(n963), .B(n962), .Z(n964) );
  AND U1333 ( .A(n965), .B(n964), .Z(n966) );
  XOR U1334 ( .A(n967), .B(n966), .Z(n969) );
  XNOR U1335 ( .A(n968), .B(n969), .Z(n1026) );
  XOR U1336 ( .A(n1027), .B(n1026), .Z(c[44]) );
  NANDN U1337 ( .A(n967), .B(n966), .Z(n971) );
  OR U1338 ( .A(n969), .B(n968), .Z(n970) );
  AND U1339 ( .A(n971), .B(n970), .Z(n1037) );
  NANDN U1340 ( .A(n973), .B(n972), .Z(n977) );
  NANDN U1341 ( .A(n975), .B(n974), .Z(n976) );
  AND U1342 ( .A(n977), .B(n976), .Z(n1091) );
  NANDN U1343 ( .A(n979), .B(n978), .Z(n983) );
  NANDN U1344 ( .A(n981), .B(n980), .Z(n982) );
  AND U1345 ( .A(n983), .B(n982), .Z(n1090) );
  NAND U1346 ( .A(b[0]), .B(a[13]), .Z(n984) );
  XNOR U1347 ( .A(b[1]), .B(n984), .Z(n986) );
  NANDN U1348 ( .A(b[0]), .B(a[12]), .Z(n985) );
  NAND U1349 ( .A(n986), .B(n985), .Z(n1075) );
  OR U1350 ( .A(n987), .B(n558), .Z(n989) );
  XOR U1351 ( .A(b[7]), .B(a[7]), .Z(n1068) );
  NAND U1352 ( .A(n7819), .B(n1068), .Z(n988) );
  NAND U1353 ( .A(n989), .B(n988), .Z(n1074) );
  XNOR U1354 ( .A(n1075), .B(n1074), .Z(n1077) );
  NAND U1355 ( .A(n571), .B(n990), .Z(n992) );
  XOR U1356 ( .A(b[11]), .B(a[3]), .Z(n1062) );
  NAND U1357 ( .A(n8135), .B(n1062), .Z(n991) );
  AND U1358 ( .A(n992), .B(n991), .Z(n1088) );
  XOR U1359 ( .A(b[13]), .B(b[12]), .Z(n1080) );
  XOR U1360 ( .A(b[13]), .B(a[0]), .Z(n993) );
  NAND U1361 ( .A(n1080), .B(n993), .Z(n994) );
  NANDN U1362 ( .A(n994), .B(n8853), .Z(n996) );
  XOR U1363 ( .A(b[13]), .B(a[1]), .Z(n1081) );
  NANDN U1364 ( .A(n8853), .B(n1081), .Z(n995) );
  NAND U1365 ( .A(n996), .B(n995), .Z(n1087) );
  XNOR U1366 ( .A(n1088), .B(n1087), .Z(n1076) );
  XOR U1367 ( .A(n1077), .B(n1076), .Z(n1049) );
  OR U1368 ( .A(n997), .B(n560), .Z(n999) );
  XOR U1369 ( .A(b[3]), .B(a[11]), .Z(n1071) );
  NAND U1370 ( .A(n7245), .B(n1071), .Z(n998) );
  AND U1371 ( .A(n999), .B(n998), .Z(n1054) );
  NAND U1372 ( .A(n570), .B(n1000), .Z(n1002) );
  XOR U1373 ( .A(b[9]), .B(a[5]), .Z(n1084) );
  NAND U1374 ( .A(n8037), .B(n1084), .Z(n1001) );
  NAND U1375 ( .A(n1002), .B(n1001), .Z(n1053) );
  XNOR U1376 ( .A(n1054), .B(n1053), .Z(n1056) );
  NANDN U1377 ( .A(b[12]), .B(b[13]), .Z(n1003) );
  NAND U1378 ( .A(n8585), .B(b[13]), .Z(n8982) );
  NAND U1379 ( .A(n1003), .B(n8982), .Z(n9073) );
  IV U1380 ( .A(n9073), .Z(n9114) );
  NOR U1381 ( .A(n9114), .B(n1007), .Z(n1055) );
  XOR U1382 ( .A(n1056), .B(n1055), .Z(n1048) );
  NANDN U1383 ( .A(n561), .B(n1004), .Z(n1006) );
  XNOR U1384 ( .A(b[5]), .B(a[9]), .Z(n1065) );
  OR U1385 ( .A(n1065), .B(n8041), .Z(n1005) );
  AND U1386 ( .A(n1006), .B(n1005), .Z(n1047) );
  XOR U1387 ( .A(n1048), .B(n1047), .Z(n1050) );
  XOR U1388 ( .A(n1049), .B(n1050), .Z(n1044) );
  NANDN U1389 ( .A(n1008), .B(n1007), .Z(n1012) );
  NANDN U1390 ( .A(n1010), .B(n1009), .Z(n1011) );
  AND U1391 ( .A(n1012), .B(n1011), .Z(n1042) );
  NANDN U1392 ( .A(n1014), .B(n1013), .Z(n1018) );
  OR U1393 ( .A(n1016), .B(n1015), .Z(n1017) );
  AND U1394 ( .A(n1018), .B(n1017), .Z(n1041) );
  XNOR U1395 ( .A(n1042), .B(n1041), .Z(n1043) );
  XNOR U1396 ( .A(n1044), .B(n1043), .Z(n1089) );
  XOR U1397 ( .A(n1090), .B(n1089), .Z(n1092) );
  XOR U1398 ( .A(n1091), .B(n1092), .Z(n1036) );
  NANDN U1399 ( .A(n1020), .B(n1019), .Z(n1024) );
  NAND U1400 ( .A(n1022), .B(n1021), .Z(n1023) );
  AND U1401 ( .A(n1024), .B(n1023), .Z(n1035) );
  XOR U1402 ( .A(n1036), .B(n1035), .Z(n1038) );
  XOR U1403 ( .A(n1037), .B(n1038), .Z(n1030) );
  XNOR U1404 ( .A(n1030), .B(sreg[45]), .Z(n1032) );
  NANDN U1405 ( .A(n1025), .B(sreg[44]), .Z(n1029) );
  NAND U1406 ( .A(n1027), .B(n1026), .Z(n1028) );
  NAND U1407 ( .A(n1029), .B(n1028), .Z(n1031) );
  XOR U1408 ( .A(n1032), .B(n1031), .Z(c[45]) );
  NANDN U1409 ( .A(n1030), .B(sreg[45]), .Z(n1034) );
  NAND U1410 ( .A(n1032), .B(n1031), .Z(n1033) );
  AND U1411 ( .A(n1034), .B(n1033), .Z(n1161) );
  XNOR U1412 ( .A(sreg[46]), .B(n1161), .Z(n1163) );
  NANDN U1413 ( .A(n1036), .B(n1035), .Z(n1040) );
  OR U1414 ( .A(n1038), .B(n1037), .Z(n1039) );
  AND U1415 ( .A(n1040), .B(n1039), .Z(n1098) );
  NANDN U1416 ( .A(n1042), .B(n1041), .Z(n1046) );
  NANDN U1417 ( .A(n1044), .B(n1043), .Z(n1045) );
  AND U1418 ( .A(n1046), .B(n1045), .Z(n1157) );
  NANDN U1419 ( .A(n1048), .B(n1047), .Z(n1052) );
  OR U1420 ( .A(n1050), .B(n1049), .Z(n1051) );
  AND U1421 ( .A(n1052), .B(n1051), .Z(n1155) );
  NANDN U1422 ( .A(n1054), .B(n1053), .Z(n1058) );
  NAND U1423 ( .A(n1056), .B(n1055), .Z(n1057) );
  AND U1424 ( .A(n1058), .B(n1057), .Z(n1142) );
  NAND U1425 ( .A(b[0]), .B(a[14]), .Z(n1059) );
  XNOR U1426 ( .A(b[1]), .B(n1059), .Z(n1061) );
  NANDN U1427 ( .A(b[0]), .B(a[13]), .Z(n1060) );
  NAND U1428 ( .A(n1061), .B(n1060), .Z(n1148) );
  XNOR U1429 ( .A(b[14]), .B(b[13]), .Z(n9067) );
  IV U1430 ( .A(n9067), .Z(n8694) );
  AND U1431 ( .A(a[0]), .B(n8694), .Z(n1145) );
  NAND U1432 ( .A(n571), .B(n1062), .Z(n1064) );
  XOR U1433 ( .A(b[11]), .B(a[4]), .Z(n1116) );
  NAND U1434 ( .A(n8135), .B(n1116), .Z(n1063) );
  AND U1435 ( .A(n1064), .B(n1063), .Z(n1146) );
  XNOR U1436 ( .A(n1145), .B(n1146), .Z(n1147) );
  XNOR U1437 ( .A(n1148), .B(n1147), .Z(n1139) );
  OR U1438 ( .A(n1065), .B(n561), .Z(n1067) );
  XOR U1439 ( .A(b[5]), .B(a[10]), .Z(n1110) );
  NAND U1440 ( .A(n7235), .B(n1110), .Z(n1066) );
  AND U1441 ( .A(n1067), .B(n1066), .Z(n1136) );
  NAND U1442 ( .A(n569), .B(n1068), .Z(n1070) );
  XOR U1443 ( .A(b[7]), .B(a[8]), .Z(n1107) );
  NAND U1444 ( .A(n7819), .B(n1107), .Z(n1069) );
  AND U1445 ( .A(n1070), .B(n1069), .Z(n1134) );
  NAND U1446 ( .A(n568), .B(n1071), .Z(n1073) );
  XOR U1447 ( .A(b[3]), .B(a[12]), .Z(n1113) );
  NAND U1448 ( .A(n7245), .B(n1113), .Z(n1072) );
  NAND U1449 ( .A(n1073), .B(n1072), .Z(n1133) );
  XNOR U1450 ( .A(n1134), .B(n1133), .Z(n1135) );
  XOR U1451 ( .A(n1136), .B(n1135), .Z(n1140) );
  XNOR U1452 ( .A(n1139), .B(n1140), .Z(n1141) );
  XNOR U1453 ( .A(n1142), .B(n1141), .Z(n1103) );
  NANDN U1454 ( .A(n1075), .B(n1074), .Z(n1079) );
  NAND U1455 ( .A(n1077), .B(n1076), .Z(n1078) );
  AND U1456 ( .A(n1079), .B(n1078), .Z(n1102) );
  NAND U1457 ( .A(n572), .B(n1081), .Z(n1083) );
  XOR U1458 ( .A(b[13]), .B(a[2]), .Z(n1130) );
  NAND U1459 ( .A(n8585), .B(n1130), .Z(n1082) );
  AND U1460 ( .A(n1083), .B(n1082), .Z(n1152) );
  NAND U1461 ( .A(n570), .B(n1084), .Z(n1086) );
  XOR U1462 ( .A(b[9]), .B(a[6]), .Z(n1123) );
  NAND U1463 ( .A(n8037), .B(n1123), .Z(n1085) );
  NAND U1464 ( .A(n1086), .B(n1085), .Z(n1151) );
  XNOR U1465 ( .A(n1152), .B(n1151), .Z(n1154) );
  NANDN U1466 ( .A(n1088), .B(n1087), .Z(n1153) );
  XNOR U1467 ( .A(n1154), .B(n1153), .Z(n1101) );
  XOR U1468 ( .A(n1102), .B(n1101), .Z(n1104) );
  XOR U1469 ( .A(n1103), .B(n1104), .Z(n1156) );
  XOR U1470 ( .A(n1155), .B(n1156), .Z(n1158) );
  XOR U1471 ( .A(n1157), .B(n1158), .Z(n1096) );
  NANDN U1472 ( .A(n1090), .B(n1089), .Z(n1094) );
  OR U1473 ( .A(n1092), .B(n1091), .Z(n1093) );
  AND U1474 ( .A(n1094), .B(n1093), .Z(n1095) );
  XNOR U1475 ( .A(n1096), .B(n1095), .Z(n1097) );
  XNOR U1476 ( .A(n1098), .B(n1097), .Z(n1162) );
  XNOR U1477 ( .A(n1163), .B(n1162), .Z(c[46]) );
  NANDN U1478 ( .A(n1096), .B(n1095), .Z(n1100) );
  NANDN U1479 ( .A(n1098), .B(n1097), .Z(n1099) );
  AND U1480 ( .A(n1100), .B(n1099), .Z(n1173) );
  NANDN U1481 ( .A(n1102), .B(n1101), .Z(n1106) );
  NANDN U1482 ( .A(n1104), .B(n1103), .Z(n1105) );
  AND U1483 ( .A(n1106), .B(n1105), .Z(n1235) );
  NAND U1484 ( .A(n569), .B(n1107), .Z(n1109) );
  XOR U1485 ( .A(b[7]), .B(a[9]), .Z(n1203) );
  NAND U1486 ( .A(n7819), .B(n1203), .Z(n1108) );
  AND U1487 ( .A(n1109), .B(n1108), .Z(n1190) );
  NAND U1488 ( .A(n567), .B(n1110), .Z(n1112) );
  XOR U1489 ( .A(b[5]), .B(a[11]), .Z(n1213) );
  NAND U1490 ( .A(n7235), .B(n1213), .Z(n1111) );
  AND U1491 ( .A(n1112), .B(n1111), .Z(n1219) );
  NAND U1492 ( .A(n568), .B(n1113), .Z(n1115) );
  XOR U1493 ( .A(b[3]), .B(a[13]), .Z(n1197) );
  NAND U1494 ( .A(n7245), .B(n1197), .Z(n1114) );
  AND U1495 ( .A(n1115), .B(n1114), .Z(n1217) );
  NAND U1496 ( .A(n571), .B(n1116), .Z(n1118) );
  XOR U1497 ( .A(b[11]), .B(a[5]), .Z(n1206) );
  NAND U1498 ( .A(n8135), .B(n1206), .Z(n1117) );
  NAND U1499 ( .A(n1118), .B(n1117), .Z(n1216) );
  XNOR U1500 ( .A(n1217), .B(n1216), .Z(n1218) );
  XNOR U1501 ( .A(n1219), .B(n1218), .Z(n1189) );
  XNOR U1502 ( .A(n1190), .B(n1189), .Z(n1192) );
  NANDN U1503 ( .A(b[14]), .B(b[15]), .Z(n1119) );
  NAND U1504 ( .A(n8694), .B(b[15]), .Z(n9121) );
  NAND U1505 ( .A(n1119), .B(n9121), .Z(n9272) );
  ANDN U1506 ( .B(n9272), .A(n1145), .Z(n1191) );
  XOR U1507 ( .A(n1192), .B(n1191), .Z(n1185) );
  NAND U1508 ( .A(b[0]), .B(a[15]), .Z(n1120) );
  XNOR U1509 ( .A(b[1]), .B(n1120), .Z(n1122) );
  NANDN U1510 ( .A(b[0]), .B(a[14]), .Z(n1121) );
  NAND U1511 ( .A(n1122), .B(n1121), .Z(n1223) );
  NAND U1512 ( .A(n570), .B(n1123), .Z(n1125) );
  XOR U1513 ( .A(b[9]), .B(a[7]), .Z(n1200) );
  NAND U1514 ( .A(n8037), .B(n1200), .Z(n1124) );
  NAND U1515 ( .A(n1125), .B(n1124), .Z(n1222) );
  XNOR U1516 ( .A(n1223), .B(n1222), .Z(n1225) );
  XOR U1517 ( .A(b[15]), .B(b[14]), .Z(n1209) );
  XOR U1518 ( .A(b[15]), .B(a[0]), .Z(n1126) );
  NAND U1519 ( .A(n1209), .B(n1126), .Z(n1127) );
  NANDN U1520 ( .A(n1127), .B(n9067), .Z(n1129) );
  XOR U1521 ( .A(b[15]), .B(a[1]), .Z(n1210) );
  NANDN U1522 ( .A(n9067), .B(n1210), .Z(n1128) );
  AND U1523 ( .A(n1129), .B(n1128), .Z(n1195) );
  NAND U1524 ( .A(n572), .B(n1130), .Z(n1132) );
  XOR U1525 ( .A(b[13]), .B(a[3]), .Z(n1231) );
  NAND U1526 ( .A(n8585), .B(n1231), .Z(n1131) );
  NAND U1527 ( .A(n1132), .B(n1131), .Z(n1196) );
  XNOR U1528 ( .A(n1195), .B(n1196), .Z(n1224) );
  XOR U1529 ( .A(n1225), .B(n1224), .Z(n1184) );
  NANDN U1530 ( .A(n1134), .B(n1133), .Z(n1138) );
  NANDN U1531 ( .A(n1136), .B(n1135), .Z(n1137) );
  AND U1532 ( .A(n1138), .B(n1137), .Z(n1183) );
  XOR U1533 ( .A(n1184), .B(n1183), .Z(n1186) );
  XNOR U1534 ( .A(n1185), .B(n1186), .Z(n1234) );
  XNOR U1535 ( .A(n1235), .B(n1234), .Z(n1237) );
  NANDN U1536 ( .A(n1140), .B(n1139), .Z(n1144) );
  NANDN U1537 ( .A(n1142), .B(n1141), .Z(n1143) );
  AND U1538 ( .A(n1144), .B(n1143), .Z(n1180) );
  NANDN U1539 ( .A(n1146), .B(n1145), .Z(n1150) );
  NANDN U1540 ( .A(n1148), .B(n1147), .Z(n1149) );
  AND U1541 ( .A(n1150), .B(n1149), .Z(n1178) );
  XNOR U1542 ( .A(n1178), .B(n1177), .Z(n1179) );
  XNOR U1543 ( .A(n1180), .B(n1179), .Z(n1236) );
  XOR U1544 ( .A(n1237), .B(n1236), .Z(n1172) );
  NANDN U1545 ( .A(n1156), .B(n1155), .Z(n1160) );
  OR U1546 ( .A(n1158), .B(n1157), .Z(n1159) );
  AND U1547 ( .A(n1160), .B(n1159), .Z(n1171) );
  XOR U1548 ( .A(n1172), .B(n1171), .Z(n1174) );
  XOR U1549 ( .A(n1173), .B(n1174), .Z(n1166) );
  XNOR U1550 ( .A(n1166), .B(sreg[47]), .Z(n1168) );
  NANDN U1551 ( .A(sreg[46]), .B(n1161), .Z(n1165) );
  NAND U1552 ( .A(n1163), .B(n1162), .Z(n1164) );
  AND U1553 ( .A(n1165), .B(n1164), .Z(n1167) );
  XOR U1554 ( .A(n1168), .B(n1167), .Z(c[47]) );
  NANDN U1555 ( .A(n1166), .B(sreg[47]), .Z(n1170) );
  NAND U1556 ( .A(n1168), .B(n1167), .Z(n1169) );
  AND U1557 ( .A(n1170), .B(n1169), .Z(n1317) );
  XNOR U1558 ( .A(sreg[48]), .B(n1317), .Z(n1319) );
  NANDN U1559 ( .A(n1172), .B(n1171), .Z(n1176) );
  OR U1560 ( .A(n1174), .B(n1173), .Z(n1175) );
  AND U1561 ( .A(n1176), .B(n1175), .Z(n1243) );
  NANDN U1562 ( .A(n1178), .B(n1177), .Z(n1182) );
  NANDN U1563 ( .A(n1180), .B(n1179), .Z(n1181) );
  AND U1564 ( .A(n1182), .B(n1181), .Z(n1313) );
  NANDN U1565 ( .A(n1184), .B(n1183), .Z(n1188) );
  OR U1566 ( .A(n1186), .B(n1185), .Z(n1187) );
  AND U1567 ( .A(n1188), .B(n1187), .Z(n1311) );
  NANDN U1568 ( .A(n1190), .B(n1189), .Z(n1194) );
  NAND U1569 ( .A(n1192), .B(n1191), .Z(n1193) );
  AND U1570 ( .A(n1194), .B(n1193), .Z(n1306) );
  ANDN U1571 ( .B(n1196), .A(n1195), .Z(n1280) );
  NANDN U1572 ( .A(n560), .B(n1197), .Z(n1199) );
  XNOR U1573 ( .A(b[3]), .B(a[14]), .Z(n1263) );
  OR U1574 ( .A(n1263), .B(n7784), .Z(n1198) );
  AND U1575 ( .A(n1199), .B(n1198), .Z(n1278) );
  NANDN U1576 ( .A(n564), .B(n1200), .Z(n1202) );
  XNOR U1577 ( .A(b[9]), .B(a[8]), .Z(n1260) );
  OR U1578 ( .A(n1260), .B(n8485), .Z(n1201) );
  NAND U1579 ( .A(n1202), .B(n1201), .Z(n1279) );
  XOR U1580 ( .A(n1278), .B(n1279), .Z(n1281) );
  XOR U1581 ( .A(n1280), .B(n1281), .Z(n1275) );
  NAND U1582 ( .A(n569), .B(n1203), .Z(n1205) );
  XOR U1583 ( .A(b[7]), .B(a[10]), .Z(n1290) );
  NAND U1584 ( .A(n7819), .B(n1290), .Z(n1204) );
  AND U1585 ( .A(n1205), .B(n1204), .Z(n1273) );
  NAND U1586 ( .A(n571), .B(n1206), .Z(n1208) );
  XOR U1587 ( .A(b[11]), .B(a[6]), .Z(n1284) );
  NAND U1588 ( .A(n8135), .B(n1284), .Z(n1207) );
  AND U1589 ( .A(n1208), .B(n1207), .Z(n1296) );
  NAND U1590 ( .A(n573), .B(n1210), .Z(n1212) );
  XOR U1591 ( .A(b[15]), .B(a[2]), .Z(n1251) );
  NAND U1592 ( .A(n8694), .B(n1251), .Z(n1211) );
  AND U1593 ( .A(n1212), .B(n1211), .Z(n1294) );
  NAND U1594 ( .A(n567), .B(n1213), .Z(n1215) );
  XOR U1595 ( .A(b[5]), .B(a[12]), .Z(n1269) );
  NAND U1596 ( .A(n7235), .B(n1269), .Z(n1214) );
  NAND U1597 ( .A(n1215), .B(n1214), .Z(n1293) );
  XNOR U1598 ( .A(n1294), .B(n1293), .Z(n1295) );
  XNOR U1599 ( .A(n1296), .B(n1295), .Z(n1272) );
  XNOR U1600 ( .A(n1273), .B(n1272), .Z(n1274) );
  XNOR U1601 ( .A(n1275), .B(n1274), .Z(n1305) );
  XNOR U1602 ( .A(n1306), .B(n1305), .Z(n1307) );
  NANDN U1603 ( .A(n1217), .B(n1216), .Z(n1221) );
  NANDN U1604 ( .A(n1219), .B(n1218), .Z(n1220) );
  AND U1605 ( .A(n1221), .B(n1220), .Z(n1302) );
  NANDN U1606 ( .A(n1223), .B(n1222), .Z(n1227) );
  NAND U1607 ( .A(n1225), .B(n1224), .Z(n1226) );
  AND U1608 ( .A(n1227), .B(n1226), .Z(n1300) );
  NAND U1609 ( .A(b[0]), .B(a[16]), .Z(n1228) );
  XNOR U1610 ( .A(b[1]), .B(n1228), .Z(n1230) );
  NANDN U1611 ( .A(b[0]), .B(a[15]), .Z(n1229) );
  NAND U1612 ( .A(n1230), .B(n1229), .Z(n1248) );
  XNOR U1613 ( .A(b[16]), .B(b[15]), .Z(n9195) );
  IV U1614 ( .A(n9195), .Z(n9141) );
  AND U1615 ( .A(a[0]), .B(n9141), .Z(n1259) );
  NAND U1616 ( .A(n572), .B(n1231), .Z(n1233) );
  XOR U1617 ( .A(b[13]), .B(a[4]), .Z(n1287) );
  NAND U1618 ( .A(n8585), .B(n1287), .Z(n1232) );
  AND U1619 ( .A(n1233), .B(n1232), .Z(n1246) );
  XNOR U1620 ( .A(n1259), .B(n1246), .Z(n1247) );
  XNOR U1621 ( .A(n1248), .B(n1247), .Z(n1299) );
  XNOR U1622 ( .A(n1300), .B(n1299), .Z(n1301) );
  XOR U1623 ( .A(n1302), .B(n1301), .Z(n1308) );
  XOR U1624 ( .A(n1307), .B(n1308), .Z(n1312) );
  XOR U1625 ( .A(n1311), .B(n1312), .Z(n1314) );
  XOR U1626 ( .A(n1313), .B(n1314), .Z(n1241) );
  NANDN U1627 ( .A(n1235), .B(n1234), .Z(n1239) );
  NAND U1628 ( .A(n1237), .B(n1236), .Z(n1238) );
  AND U1629 ( .A(n1239), .B(n1238), .Z(n1240) );
  XNOR U1630 ( .A(n1241), .B(n1240), .Z(n1242) );
  XNOR U1631 ( .A(n1243), .B(n1242), .Z(n1318) );
  XNOR U1632 ( .A(n1319), .B(n1318), .Z(c[48]) );
  NANDN U1633 ( .A(n1241), .B(n1240), .Z(n1245) );
  NANDN U1634 ( .A(n1243), .B(n1242), .Z(n1244) );
  AND U1635 ( .A(n1245), .B(n1244), .Z(n1325) );
  NANDN U1636 ( .A(n1246), .B(n1259), .Z(n1250) );
  NANDN U1637 ( .A(n1248), .B(n1247), .Z(n1249) );
  AND U1638 ( .A(n1250), .B(n1249), .Z(n1384) );
  NAND U1639 ( .A(n573), .B(n1251), .Z(n1253) );
  XOR U1640 ( .A(b[15]), .B(a[3]), .Z(n1352) );
  NAND U1641 ( .A(n8694), .B(n1352), .Z(n1252) );
  AND U1642 ( .A(n1253), .B(n1252), .Z(n1347) );
  XOR U1643 ( .A(b[17]), .B(b[16]), .Z(n1340) );
  XOR U1644 ( .A(b[17]), .B(a[0]), .Z(n1254) );
  NAND U1645 ( .A(n1340), .B(n1254), .Z(n1255) );
  NANDN U1646 ( .A(n1255), .B(n9195), .Z(n1257) );
  XOR U1647 ( .A(b[17]), .B(a[1]), .Z(n1341) );
  NANDN U1648 ( .A(n9195), .B(n1341), .Z(n1256) );
  AND U1649 ( .A(n1257), .B(n1256), .Z(n1348) );
  XOR U1650 ( .A(n1347), .B(n1348), .Z(n1336) );
  NANDN U1651 ( .A(b[16]), .B(b[17]), .Z(n1258) );
  NAND U1652 ( .A(n9141), .B(b[17]), .Z(n9299) );
  NAND U1653 ( .A(n1258), .B(n9299), .Z(n9373) );
  ANDN U1654 ( .B(n9373), .A(n1259), .Z(n1335) );
  OR U1655 ( .A(n1260), .B(n564), .Z(n1262) );
  XNOR U1656 ( .A(b[9]), .B(a[9]), .Z(n1367) );
  OR U1657 ( .A(n1367), .B(n8485), .Z(n1261) );
  AND U1658 ( .A(n1262), .B(n1261), .Z(n1334) );
  XOR U1659 ( .A(n1335), .B(n1334), .Z(n1337) );
  XOR U1660 ( .A(n1336), .B(n1337), .Z(n1383) );
  OR U1661 ( .A(n1263), .B(n560), .Z(n1265) );
  XOR U1662 ( .A(b[3]), .B(a[15]), .Z(n1373) );
  NAND U1663 ( .A(n7245), .B(n1373), .Z(n1264) );
  AND U1664 ( .A(n1265), .B(n1264), .Z(n1379) );
  NAND U1665 ( .A(b[0]), .B(a[17]), .Z(n1266) );
  XNOR U1666 ( .A(b[1]), .B(n1266), .Z(n1268) );
  NANDN U1667 ( .A(b[0]), .B(a[16]), .Z(n1267) );
  NAND U1668 ( .A(n1268), .B(n1267), .Z(n1377) );
  NAND U1669 ( .A(n567), .B(n1269), .Z(n1271) );
  XOR U1670 ( .A(b[5]), .B(a[13]), .Z(n1361) );
  NAND U1671 ( .A(n7235), .B(n1361), .Z(n1270) );
  NAND U1672 ( .A(n1271), .B(n1270), .Z(n1376) );
  XNOR U1673 ( .A(n1377), .B(n1376), .Z(n1378) );
  XNOR U1674 ( .A(n1379), .B(n1378), .Z(n1382) );
  XOR U1675 ( .A(n1383), .B(n1382), .Z(n1385) );
  XOR U1676 ( .A(n1384), .B(n1385), .Z(n1329) );
  NANDN U1677 ( .A(n1273), .B(n1272), .Z(n1277) );
  NANDN U1678 ( .A(n1275), .B(n1274), .Z(n1276) );
  AND U1679 ( .A(n1277), .B(n1276), .Z(n1328) );
  XNOR U1680 ( .A(n1329), .B(n1328), .Z(n1330) );
  NANDN U1681 ( .A(n1279), .B(n1278), .Z(n1283) );
  OR U1682 ( .A(n1281), .B(n1280), .Z(n1282) );
  AND U1683 ( .A(n1283), .B(n1282), .Z(n1389) );
  NAND U1684 ( .A(n571), .B(n1284), .Z(n1286) );
  XOR U1685 ( .A(b[11]), .B(a[7]), .Z(n1344) );
  NAND U1686 ( .A(n8135), .B(n1344), .Z(n1285) );
  AND U1687 ( .A(n1286), .B(n1285), .Z(n1357) );
  NAND U1688 ( .A(n572), .B(n1287), .Z(n1289) );
  XOR U1689 ( .A(b[13]), .B(a[5]), .Z(n1370) );
  NAND U1690 ( .A(n8585), .B(n1370), .Z(n1288) );
  AND U1691 ( .A(n1289), .B(n1288), .Z(n1356) );
  NAND U1692 ( .A(n569), .B(n1290), .Z(n1292) );
  XOR U1693 ( .A(b[7]), .B(a[11]), .Z(n1364) );
  NAND U1694 ( .A(n7819), .B(n1364), .Z(n1291) );
  NAND U1695 ( .A(n1292), .B(n1291), .Z(n1355) );
  XOR U1696 ( .A(n1356), .B(n1355), .Z(n1358) );
  XNOR U1697 ( .A(n1357), .B(n1358), .Z(n1388) );
  XNOR U1698 ( .A(n1389), .B(n1388), .Z(n1390) );
  NANDN U1699 ( .A(n1294), .B(n1293), .Z(n1298) );
  NANDN U1700 ( .A(n1296), .B(n1295), .Z(n1297) );
  NAND U1701 ( .A(n1298), .B(n1297), .Z(n1391) );
  XOR U1702 ( .A(n1390), .B(n1391), .Z(n1331) );
  XNOR U1703 ( .A(n1330), .B(n1331), .Z(n1396) );
  NANDN U1704 ( .A(n1300), .B(n1299), .Z(n1304) );
  NANDN U1705 ( .A(n1302), .B(n1301), .Z(n1303) );
  AND U1706 ( .A(n1304), .B(n1303), .Z(n1394) );
  NANDN U1707 ( .A(n1306), .B(n1305), .Z(n1310) );
  NANDN U1708 ( .A(n1308), .B(n1307), .Z(n1309) );
  NAND U1709 ( .A(n1310), .B(n1309), .Z(n1395) );
  XOR U1710 ( .A(n1394), .B(n1395), .Z(n1397) );
  XNOR U1711 ( .A(n1396), .B(n1397), .Z(n1322) );
  NANDN U1712 ( .A(n1312), .B(n1311), .Z(n1316) );
  OR U1713 ( .A(n1314), .B(n1313), .Z(n1315) );
  NAND U1714 ( .A(n1316), .B(n1315), .Z(n1323) );
  XNOR U1715 ( .A(n1322), .B(n1323), .Z(n1324) );
  XNOR U1716 ( .A(n1325), .B(n1324), .Z(n1400) );
  XNOR U1717 ( .A(sreg[49]), .B(n1400), .Z(n1402) );
  NANDN U1718 ( .A(sreg[48]), .B(n1317), .Z(n1321) );
  NAND U1719 ( .A(n1319), .B(n1318), .Z(n1320) );
  NAND U1720 ( .A(n1321), .B(n1320), .Z(n1401) );
  XNOR U1721 ( .A(n1402), .B(n1401), .Z(c[49]) );
  NANDN U1722 ( .A(n1323), .B(n1322), .Z(n1327) );
  NANDN U1723 ( .A(n1325), .B(n1324), .Z(n1326) );
  AND U1724 ( .A(n1327), .B(n1326), .Z(n1410) );
  NANDN U1725 ( .A(n1329), .B(n1328), .Z(n1333) );
  NANDN U1726 ( .A(n1331), .B(n1330), .Z(n1332) );
  AND U1727 ( .A(n1333), .B(n1332), .Z(n1491) );
  NANDN U1728 ( .A(n1335), .B(n1334), .Z(n1339) );
  OR U1729 ( .A(n1337), .B(n1336), .Z(n1338) );
  AND U1730 ( .A(n1339), .B(n1338), .Z(n1478) );
  NAND U1731 ( .A(n576), .B(n1341), .Z(n1343) );
  XOR U1732 ( .A(b[17]), .B(a[2]), .Z(n1462) );
  NAND U1733 ( .A(n9141), .B(n1462), .Z(n1342) );
  AND U1734 ( .A(n1343), .B(n1342), .Z(n1453) );
  NAND U1735 ( .A(n571), .B(n1344), .Z(n1346) );
  XOR U1736 ( .A(b[11]), .B(a[8]), .Z(n1449) );
  NAND U1737 ( .A(n8135), .B(n1449), .Z(n1345) );
  NAND U1738 ( .A(n1346), .B(n1345), .Z(n1452) );
  XNOR U1739 ( .A(n1453), .B(n1452), .Z(n1455) );
  NOR U1740 ( .A(n1348), .B(n1347), .Z(n1454) );
  XOR U1741 ( .A(n1455), .B(n1454), .Z(n1477) );
  NAND U1742 ( .A(b[0]), .B(a[18]), .Z(n1349) );
  XNOR U1743 ( .A(b[1]), .B(n1349), .Z(n1351) );
  NANDN U1744 ( .A(b[0]), .B(a[17]), .Z(n1350) );
  NAND U1745 ( .A(n1351), .B(n1350), .Z(n1428) );
  AND U1746 ( .A(a[0]), .B(n575), .Z(n1466) );
  NAND U1747 ( .A(n573), .B(n1352), .Z(n1354) );
  XOR U1748 ( .A(b[15]), .B(a[4]), .Z(n1437) );
  NAND U1749 ( .A(n8694), .B(n1437), .Z(n1353) );
  NAND U1750 ( .A(n1354), .B(n1353), .Z(n1426) );
  XOR U1751 ( .A(n1466), .B(n1426), .Z(n1427) );
  XOR U1752 ( .A(n1428), .B(n1427), .Z(n1476) );
  XOR U1753 ( .A(n1477), .B(n1476), .Z(n1479) );
  XOR U1754 ( .A(n1478), .B(n1479), .Z(n1484) );
  NANDN U1755 ( .A(n1356), .B(n1355), .Z(n1360) );
  OR U1756 ( .A(n1358), .B(n1357), .Z(n1359) );
  AND U1757 ( .A(n1360), .B(n1359), .Z(n1483) );
  NAND U1758 ( .A(n567), .B(n1361), .Z(n1363) );
  XOR U1759 ( .A(b[5]), .B(a[14]), .Z(n1440) );
  NAND U1760 ( .A(n7235), .B(n1440), .Z(n1362) );
  AND U1761 ( .A(n1363), .B(n1362), .Z(n1421) );
  NAND U1762 ( .A(n569), .B(n1364), .Z(n1366) );
  XOR U1763 ( .A(b[7]), .B(a[12]), .Z(n1431) );
  NAND U1764 ( .A(n7819), .B(n1431), .Z(n1365) );
  NAND U1765 ( .A(n1366), .B(n1365), .Z(n1420) );
  XNOR U1766 ( .A(n1421), .B(n1420), .Z(n1422) );
  OR U1767 ( .A(n1367), .B(n564), .Z(n1369) );
  XOR U1768 ( .A(b[9]), .B(a[10]), .Z(n1467) );
  NAND U1769 ( .A(n8037), .B(n1467), .Z(n1368) );
  AND U1770 ( .A(n1369), .B(n1368), .Z(n1473) );
  NAND U1771 ( .A(n572), .B(n1370), .Z(n1372) );
  XOR U1772 ( .A(b[13]), .B(a[6]), .Z(n1434) );
  NAND U1773 ( .A(n8585), .B(n1434), .Z(n1371) );
  AND U1774 ( .A(n1372), .B(n1371), .Z(n1471) );
  NAND U1775 ( .A(n568), .B(n1373), .Z(n1375) );
  XOR U1776 ( .A(b[3]), .B(a[16]), .Z(n1443) );
  NAND U1777 ( .A(n7245), .B(n1443), .Z(n1374) );
  NAND U1778 ( .A(n1375), .B(n1374), .Z(n1470) );
  XNOR U1779 ( .A(n1471), .B(n1470), .Z(n1472) );
  XOR U1780 ( .A(n1473), .B(n1472), .Z(n1423) );
  XNOR U1781 ( .A(n1422), .B(n1423), .Z(n1482) );
  XOR U1782 ( .A(n1483), .B(n1482), .Z(n1485) );
  XOR U1783 ( .A(n1484), .B(n1485), .Z(n1416) );
  NANDN U1784 ( .A(n1377), .B(n1376), .Z(n1381) );
  NANDN U1785 ( .A(n1379), .B(n1378), .Z(n1380) );
  AND U1786 ( .A(n1381), .B(n1380), .Z(n1414) );
  NANDN U1787 ( .A(n1383), .B(n1382), .Z(n1387) );
  OR U1788 ( .A(n1385), .B(n1384), .Z(n1386) );
  NAND U1789 ( .A(n1387), .B(n1386), .Z(n1415) );
  XOR U1790 ( .A(n1414), .B(n1415), .Z(n1417) );
  XOR U1791 ( .A(n1416), .B(n1417), .Z(n1489) );
  NANDN U1792 ( .A(n1389), .B(n1388), .Z(n1393) );
  NANDN U1793 ( .A(n1391), .B(n1390), .Z(n1392) );
  AND U1794 ( .A(n1393), .B(n1392), .Z(n1488) );
  XNOR U1795 ( .A(n1489), .B(n1488), .Z(n1490) );
  XOR U1796 ( .A(n1491), .B(n1490), .Z(n1409) );
  NANDN U1797 ( .A(n1395), .B(n1394), .Z(n1399) );
  NANDN U1798 ( .A(n1397), .B(n1396), .Z(n1398) );
  NAND U1799 ( .A(n1399), .B(n1398), .Z(n1408) );
  XOR U1800 ( .A(n1409), .B(n1408), .Z(n1411) );
  XNOR U1801 ( .A(n1410), .B(n1411), .Z(n1407) );
  NANDN U1802 ( .A(sreg[49]), .B(n1400), .Z(n1404) );
  NAND U1803 ( .A(n1402), .B(n1401), .Z(n1403) );
  AND U1804 ( .A(n1404), .B(n1403), .Z(n1406) );
  XNOR U1805 ( .A(sreg[50]), .B(n1406), .Z(n1405) );
  XNOR U1806 ( .A(n1407), .B(n1405), .Z(c[50]) );
  NANDN U1807 ( .A(n1409), .B(n1408), .Z(n1413) );
  OR U1808 ( .A(n1411), .B(n1410), .Z(n1412) );
  AND U1809 ( .A(n1413), .B(n1412), .Z(n1502) );
  NANDN U1810 ( .A(n1415), .B(n1414), .Z(n1419) );
  OR U1811 ( .A(n1417), .B(n1416), .Z(n1418) );
  AND U1812 ( .A(n1419), .B(n1418), .Z(n1583) );
  NANDN U1813 ( .A(n1421), .B(n1420), .Z(n1425) );
  NANDN U1814 ( .A(n1423), .B(n1422), .Z(n1424) );
  NAND U1815 ( .A(n1425), .B(n1424), .Z(n1506) );
  NAND U1816 ( .A(n1466), .B(n1426), .Z(n1430) );
  NANDN U1817 ( .A(n1428), .B(n1427), .Z(n1429) );
  NAND U1818 ( .A(n1430), .B(n1429), .Z(n1505) );
  XOR U1819 ( .A(n1506), .B(n1505), .Z(n1508) );
  NAND U1820 ( .A(n569), .B(n1431), .Z(n1433) );
  XOR U1821 ( .A(b[7]), .B(a[13]), .Z(n1532) );
  NAND U1822 ( .A(n7819), .B(n1532), .Z(n1432) );
  AND U1823 ( .A(n1433), .B(n1432), .Z(n1575) );
  NAND U1824 ( .A(n572), .B(n1434), .Z(n1436) );
  XOR U1825 ( .A(b[13]), .B(a[7]), .Z(n1565) );
  NAND U1826 ( .A(n8585), .B(n1565), .Z(n1435) );
  AND U1827 ( .A(n1436), .B(n1435), .Z(n1520) );
  NAND U1828 ( .A(n573), .B(n1437), .Z(n1439) );
  XOR U1829 ( .A(b[15]), .B(a[5]), .Z(n1562) );
  NAND U1830 ( .A(n8694), .B(n1562), .Z(n1438) );
  AND U1831 ( .A(n1439), .B(n1438), .Z(n1518) );
  NAND U1832 ( .A(n567), .B(n1440), .Z(n1442) );
  XOR U1833 ( .A(b[5]), .B(a[15]), .Z(n1529) );
  NAND U1834 ( .A(n7235), .B(n1529), .Z(n1441) );
  NAND U1835 ( .A(n1442), .B(n1441), .Z(n1517) );
  XNOR U1836 ( .A(n1518), .B(n1517), .Z(n1519) );
  XNOR U1837 ( .A(n1520), .B(n1519), .Z(n1574) );
  XNOR U1838 ( .A(n1575), .B(n1574), .Z(n1576) );
  NAND U1839 ( .A(n568), .B(n1443), .Z(n1445) );
  XOR U1840 ( .A(b[3]), .B(a[17]), .Z(n1535) );
  NAND U1841 ( .A(n7245), .B(n1535), .Z(n1444) );
  AND U1842 ( .A(n1445), .B(n1444), .Z(n1547) );
  NAND U1843 ( .A(b[0]), .B(a[19]), .Z(n1446) );
  XNOR U1844 ( .A(b[1]), .B(n1446), .Z(n1448) );
  NANDN U1845 ( .A(b[0]), .B(a[18]), .Z(n1447) );
  NAND U1846 ( .A(n1448), .B(n1447), .Z(n1545) );
  NAND U1847 ( .A(n571), .B(n1449), .Z(n1451) );
  XOR U1848 ( .A(b[11]), .B(a[9]), .Z(n1554) );
  NAND U1849 ( .A(n8135), .B(n1554), .Z(n1450) );
  NAND U1850 ( .A(n1451), .B(n1450), .Z(n1544) );
  XNOR U1851 ( .A(n1545), .B(n1544), .Z(n1546) );
  XOR U1852 ( .A(n1547), .B(n1546), .Z(n1577) );
  XNOR U1853 ( .A(n1576), .B(n1577), .Z(n1507) );
  XOR U1854 ( .A(n1508), .B(n1507), .Z(n1514) );
  NANDN U1855 ( .A(n1453), .B(n1452), .Z(n1457) );
  NAND U1856 ( .A(n1455), .B(n1454), .Z(n1456) );
  AND U1857 ( .A(n1457), .B(n1456), .Z(n1570) );
  XOR U1858 ( .A(b[19]), .B(b[18]), .Z(n1550) );
  XOR U1859 ( .A(b[19]), .B(a[0]), .Z(n1458) );
  NAND U1860 ( .A(n1550), .B(n1458), .Z(n1459) );
  NANDN U1861 ( .A(n1459), .B(n555), .Z(n1461) );
  XOR U1862 ( .A(b[19]), .B(a[1]), .Z(n1551) );
  NANDN U1863 ( .A(n555), .B(n1551), .Z(n1460) );
  AND U1864 ( .A(n1461), .B(n1460), .Z(n1558) );
  NAND U1865 ( .A(n576), .B(n1462), .Z(n1464) );
  XOR U1866 ( .A(b[17]), .B(a[3]), .Z(n1526) );
  NAND U1867 ( .A(n9141), .B(n1526), .Z(n1463) );
  AND U1868 ( .A(n1464), .B(n1463), .Z(n1557) );
  XOR U1869 ( .A(n1558), .B(n1557), .Z(n1540) );
  NANDN U1870 ( .A(b[18]), .B(b[19]), .Z(n1465) );
  NAND U1871 ( .A(n575), .B(b[19]), .Z(n9428) );
  NAND U1872 ( .A(n1465), .B(n9428), .Z(n9521) );
  ANDN U1873 ( .B(n9521), .A(n1466), .Z(n1539) );
  NANDN U1874 ( .A(n564), .B(n1467), .Z(n1469) );
  XNOR U1875 ( .A(b[9]), .B(a[11]), .Z(n1559) );
  OR U1876 ( .A(n1559), .B(n8485), .Z(n1468) );
  AND U1877 ( .A(n1469), .B(n1468), .Z(n1538) );
  XOR U1878 ( .A(n1539), .B(n1538), .Z(n1541) );
  XOR U1879 ( .A(n1540), .B(n1541), .Z(n1569) );
  NANDN U1880 ( .A(n1471), .B(n1470), .Z(n1475) );
  NANDN U1881 ( .A(n1473), .B(n1472), .Z(n1474) );
  NAND U1882 ( .A(n1475), .B(n1474), .Z(n1568) );
  XOR U1883 ( .A(n1569), .B(n1568), .Z(n1571) );
  XOR U1884 ( .A(n1570), .B(n1571), .Z(n1512) );
  NANDN U1885 ( .A(n1477), .B(n1476), .Z(n1481) );
  OR U1886 ( .A(n1479), .B(n1478), .Z(n1480) );
  NAND U1887 ( .A(n1481), .B(n1480), .Z(n1511) );
  XNOR U1888 ( .A(n1512), .B(n1511), .Z(n1513) );
  XNOR U1889 ( .A(n1514), .B(n1513), .Z(n1580) );
  NANDN U1890 ( .A(n1483), .B(n1482), .Z(n1487) );
  OR U1891 ( .A(n1485), .B(n1484), .Z(n1486) );
  NAND U1892 ( .A(n1487), .B(n1486), .Z(n1581) );
  XNOR U1893 ( .A(n1580), .B(n1581), .Z(n1582) );
  XNOR U1894 ( .A(n1583), .B(n1582), .Z(n1499) );
  NANDN U1895 ( .A(n1489), .B(n1488), .Z(n1493) );
  NAND U1896 ( .A(n1491), .B(n1490), .Z(n1492) );
  NAND U1897 ( .A(n1493), .B(n1492), .Z(n1500) );
  XNOR U1898 ( .A(n1499), .B(n1500), .Z(n1501) );
  XOR U1899 ( .A(n1502), .B(n1501), .Z(n1494) );
  XNOR U1900 ( .A(sreg[51]), .B(n1494), .Z(n1496) );
  XNOR U1901 ( .A(n1495), .B(n1496), .Z(c[51]) );
  OR U1902 ( .A(sreg[51]), .B(n1494), .Z(n1498) );
  OR U1903 ( .A(n1496), .B(n1495), .Z(n1497) );
  NAND U1904 ( .A(n1498), .B(n1497), .Z(n1677) );
  XNOR U1905 ( .A(sreg[52]), .B(n1677), .Z(n1679) );
  NANDN U1906 ( .A(n1500), .B(n1499), .Z(n1504) );
  NANDN U1907 ( .A(n1502), .B(n1501), .Z(n1503) );
  AND U1908 ( .A(n1504), .B(n1503), .Z(n1589) );
  NAND U1909 ( .A(n1506), .B(n1505), .Z(n1510) );
  NAND U1910 ( .A(n1508), .B(n1507), .Z(n1509) );
  AND U1911 ( .A(n1510), .B(n1509), .Z(n1672) );
  NANDN U1912 ( .A(n1512), .B(n1511), .Z(n1516) );
  NANDN U1913 ( .A(n1514), .B(n1513), .Z(n1515) );
  AND U1914 ( .A(n1516), .B(n1515), .Z(n1671) );
  XNOR U1915 ( .A(n1672), .B(n1671), .Z(n1674) );
  NANDN U1916 ( .A(n1518), .B(n1517), .Z(n1522) );
  NANDN U1917 ( .A(n1520), .B(n1519), .Z(n1521) );
  AND U1918 ( .A(n1522), .B(n1521), .Z(n1655) );
  NAND U1919 ( .A(b[0]), .B(a[20]), .Z(n1523) );
  XNOR U1920 ( .A(b[1]), .B(n1523), .Z(n1525) );
  NANDN U1921 ( .A(b[0]), .B(a[19]), .Z(n1524) );
  NAND U1922 ( .A(n1525), .B(n1524), .Z(n1638) );
  XNOR U1923 ( .A(b[20]), .B(b[19]), .Z(n9480) );
  IV U1924 ( .A(n9480), .Z(n9216) );
  AND U1925 ( .A(a[0]), .B(n9216), .Z(n1635) );
  NAND U1926 ( .A(n576), .B(n1526), .Z(n1528) );
  XOR U1927 ( .A(b[17]), .B(a[4]), .Z(n1609) );
  NAND U1928 ( .A(n9141), .B(n1609), .Z(n1527) );
  AND U1929 ( .A(n1528), .B(n1527), .Z(n1636) );
  XNOR U1930 ( .A(n1635), .B(n1636), .Z(n1637) );
  XNOR U1931 ( .A(n1638), .B(n1637), .Z(n1653) );
  NAND U1932 ( .A(n567), .B(n1529), .Z(n1531) );
  XOR U1933 ( .A(b[5]), .B(a[16]), .Z(n1603) );
  NAND U1934 ( .A(n7235), .B(n1603), .Z(n1530) );
  AND U1935 ( .A(n1531), .B(n1530), .Z(n1650) );
  NAND U1936 ( .A(n569), .B(n1532), .Z(n1534) );
  XOR U1937 ( .A(b[7]), .B(a[14]), .Z(n1600) );
  NAND U1938 ( .A(n7819), .B(n1600), .Z(n1533) );
  AND U1939 ( .A(n1534), .B(n1533), .Z(n1648) );
  NAND U1940 ( .A(n568), .B(n1535), .Z(n1537) );
  XOR U1941 ( .A(b[3]), .B(a[18]), .Z(n1615) );
  NAND U1942 ( .A(n7245), .B(n1615), .Z(n1536) );
  NAND U1943 ( .A(n1537), .B(n1536), .Z(n1647) );
  XNOR U1944 ( .A(n1648), .B(n1647), .Z(n1649) );
  XOR U1945 ( .A(n1650), .B(n1649), .Z(n1654) );
  XOR U1946 ( .A(n1653), .B(n1654), .Z(n1656) );
  XOR U1947 ( .A(n1655), .B(n1656), .Z(n1661) );
  NANDN U1948 ( .A(n1539), .B(n1538), .Z(n1543) );
  OR U1949 ( .A(n1541), .B(n1540), .Z(n1542) );
  AND U1950 ( .A(n1543), .B(n1542), .Z(n1660) );
  NANDN U1951 ( .A(n1545), .B(n1544), .Z(n1549) );
  NANDN U1952 ( .A(n1547), .B(n1546), .Z(n1548) );
  AND U1953 ( .A(n1549), .B(n1548), .Z(n1595) );
  AND U1954 ( .A(n1550), .B(n555), .Z(n9046) );
  NAND U1955 ( .A(n9046), .B(n1551), .Z(n1553) );
  XOR U1956 ( .A(b[19]), .B(a[2]), .Z(n1628) );
  NAND U1957 ( .A(n575), .B(n1628), .Z(n1552) );
  AND U1958 ( .A(n1553), .B(n1552), .Z(n1597) );
  NAND U1959 ( .A(n571), .B(n1554), .Z(n1556) );
  XOR U1960 ( .A(b[11]), .B(a[10]), .Z(n1632) );
  NAND U1961 ( .A(n8135), .B(n1632), .Z(n1555) );
  NAND U1962 ( .A(n1556), .B(n1555), .Z(n1596) );
  XNOR U1963 ( .A(n1597), .B(n1596), .Z(n1599) );
  OR U1964 ( .A(n1558), .B(n1557), .Z(n1598) );
  XNOR U1965 ( .A(n1599), .B(n1598), .Z(n1593) );
  OR U1966 ( .A(n1559), .B(n564), .Z(n1561) );
  XNOR U1967 ( .A(b[9]), .B(a[12]), .Z(n1621) );
  OR U1968 ( .A(n1621), .B(n8485), .Z(n1560) );
  NAND U1969 ( .A(n1561), .B(n1560), .Z(n1642) );
  NAND U1970 ( .A(n573), .B(n1562), .Z(n1564) );
  XOR U1971 ( .A(b[15]), .B(a[6]), .Z(n1612) );
  NAND U1972 ( .A(n8694), .B(n1612), .Z(n1563) );
  NAND U1973 ( .A(n1564), .B(n1563), .Z(n1641) );
  XOR U1974 ( .A(n1642), .B(n1641), .Z(n1644) );
  NANDN U1975 ( .A(n553), .B(n1565), .Z(n1567) );
  XNOR U1976 ( .A(b[13]), .B(a[8]), .Z(n1606) );
  OR U1977 ( .A(n1606), .B(n8853), .Z(n1566) );
  NAND U1978 ( .A(n1567), .B(n1566), .Z(n1643) );
  XNOR U1979 ( .A(n1644), .B(n1643), .Z(n1592) );
  XNOR U1980 ( .A(n1593), .B(n1592), .Z(n1594) );
  XOR U1981 ( .A(n1595), .B(n1594), .Z(n1659) );
  XOR U1982 ( .A(n1660), .B(n1659), .Z(n1662) );
  XOR U1983 ( .A(n1661), .B(n1662), .Z(n1668) );
  NANDN U1984 ( .A(n1569), .B(n1568), .Z(n1573) );
  OR U1985 ( .A(n1571), .B(n1570), .Z(n1572) );
  AND U1986 ( .A(n1573), .B(n1572), .Z(n1666) );
  NANDN U1987 ( .A(n1575), .B(n1574), .Z(n1579) );
  NANDN U1988 ( .A(n1577), .B(n1576), .Z(n1578) );
  NAND U1989 ( .A(n1579), .B(n1578), .Z(n1665) );
  XNOR U1990 ( .A(n1666), .B(n1665), .Z(n1667) );
  XNOR U1991 ( .A(n1668), .B(n1667), .Z(n1673) );
  XOR U1992 ( .A(n1674), .B(n1673), .Z(n1587) );
  NANDN U1993 ( .A(n1581), .B(n1580), .Z(n1585) );
  NANDN U1994 ( .A(n1583), .B(n1582), .Z(n1584) );
  NAND U1995 ( .A(n1585), .B(n1584), .Z(n1586) );
  XNOR U1996 ( .A(n1587), .B(n1586), .Z(n1588) );
  XNOR U1997 ( .A(n1589), .B(n1588), .Z(n1678) );
  XNOR U1998 ( .A(n1679), .B(n1678), .Z(c[52]) );
  NANDN U1999 ( .A(n1587), .B(n1586), .Z(n1591) );
  NANDN U2000 ( .A(n1589), .B(n1588), .Z(n1590) );
  AND U2001 ( .A(n1591), .B(n1590), .Z(n1689) );
  NAND U2002 ( .A(n569), .B(n1600), .Z(n1602) );
  XOR U2003 ( .A(b[7]), .B(a[15]), .Z(n1741) );
  NAND U2004 ( .A(n7819), .B(n1741), .Z(n1601) );
  AND U2005 ( .A(n1602), .B(n1601), .Z(n1716) );
  NAND U2006 ( .A(n567), .B(n1603), .Z(n1605) );
  XOR U2007 ( .A(b[5]), .B(a[17]), .Z(n1744) );
  NAND U2008 ( .A(n7235), .B(n1744), .Z(n1604) );
  NAND U2009 ( .A(n1605), .B(n1604), .Z(n1715) );
  XNOR U2010 ( .A(n1716), .B(n1715), .Z(n1717) );
  OR U2011 ( .A(n1606), .B(n553), .Z(n1608) );
  XOR U2012 ( .A(b[13]), .B(a[9]), .Z(n1730) );
  NAND U2013 ( .A(n8585), .B(n1730), .Z(n1607) );
  AND U2014 ( .A(n1608), .B(n1607), .Z(n1766) );
  NAND U2015 ( .A(n576), .B(n1609), .Z(n1611) );
  XOR U2016 ( .A(b[17]), .B(a[5]), .Z(n1750) );
  NAND U2017 ( .A(n9141), .B(n1750), .Z(n1610) );
  AND U2018 ( .A(n1611), .B(n1610), .Z(n1764) );
  NAND U2019 ( .A(n573), .B(n1612), .Z(n1614) );
  XOR U2020 ( .A(b[15]), .B(a[7]), .Z(n1747) );
  NAND U2021 ( .A(n8694), .B(n1747), .Z(n1613) );
  NAND U2022 ( .A(n1614), .B(n1613), .Z(n1763) );
  XNOR U2023 ( .A(n1764), .B(n1763), .Z(n1765) );
  XOR U2024 ( .A(n1766), .B(n1765), .Z(n1718) );
  XNOR U2025 ( .A(n1717), .B(n1718), .Z(n1705) );
  XNOR U2026 ( .A(n1706), .B(n1705), .Z(n1708) );
  NAND U2027 ( .A(n568), .B(n1615), .Z(n1617) );
  XOR U2028 ( .A(b[3]), .B(a[19]), .Z(n1727) );
  NAND U2029 ( .A(n7245), .B(n1727), .Z(n1616) );
  AND U2030 ( .A(n1617), .B(n1616), .Z(n1772) );
  NAND U2031 ( .A(b[0]), .B(a[21]), .Z(n1618) );
  XNOR U2032 ( .A(b[1]), .B(n1618), .Z(n1620) );
  NANDN U2033 ( .A(b[0]), .B(a[20]), .Z(n1619) );
  NAND U2034 ( .A(n1620), .B(n1619), .Z(n1770) );
  OR U2035 ( .A(n1621), .B(n564), .Z(n1623) );
  XOR U2036 ( .A(b[9]), .B(a[13]), .Z(n1757) );
  NAND U2037 ( .A(n8037), .B(n1757), .Z(n1622) );
  NAND U2038 ( .A(n1623), .B(n1622), .Z(n1769) );
  XNOR U2039 ( .A(n1770), .B(n1769), .Z(n1771) );
  XNOR U2040 ( .A(n1772), .B(n1771), .Z(n1710) );
  XOR U2041 ( .A(b[21]), .B(b[20]), .Z(n1753) );
  XOR U2042 ( .A(b[21]), .B(a[0]), .Z(n1624) );
  NAND U2043 ( .A(n1753), .B(n1624), .Z(n1625) );
  NANDN U2044 ( .A(n1625), .B(n9480), .Z(n1627) );
  XOR U2045 ( .A(b[21]), .B(a[1]), .Z(n1754) );
  NANDN U2046 ( .A(n9480), .B(n1754), .Z(n1626) );
  AND U2047 ( .A(n1627), .B(n1626), .Z(n1734) );
  NAND U2048 ( .A(n9046), .B(n1628), .Z(n1630) );
  XOR U2049 ( .A(b[19]), .B(a[3]), .Z(n1738) );
  NAND U2050 ( .A(n575), .B(n1738), .Z(n1629) );
  AND U2051 ( .A(n1630), .B(n1629), .Z(n1733) );
  XOR U2052 ( .A(n1734), .B(n1733), .Z(n1724) );
  NANDN U2053 ( .A(b[20]), .B(b[21]), .Z(n1631) );
  NAND U2054 ( .A(n9216), .B(b[21]), .Z(n9541) );
  NAND U2055 ( .A(n1631), .B(n9541), .Z(n9651) );
  ANDN U2056 ( .B(n9651), .A(n1635), .Z(n1722) );
  NANDN U2057 ( .A(n562), .B(n1632), .Z(n1634) );
  XNOR U2058 ( .A(b[11]), .B(a[11]), .Z(n1760) );
  OR U2059 ( .A(n1760), .B(n8701), .Z(n1633) );
  AND U2060 ( .A(n1634), .B(n1633), .Z(n1721) );
  XNOR U2061 ( .A(n1722), .B(n1721), .Z(n1723) );
  XOR U2062 ( .A(n1724), .B(n1723), .Z(n1709) );
  XOR U2063 ( .A(n1710), .B(n1709), .Z(n1712) );
  NANDN U2064 ( .A(n1636), .B(n1635), .Z(n1640) );
  NANDN U2065 ( .A(n1638), .B(n1637), .Z(n1639) );
  NAND U2066 ( .A(n1640), .B(n1639), .Z(n1711) );
  XNOR U2067 ( .A(n1712), .B(n1711), .Z(n1707) );
  XNOR U2068 ( .A(n1708), .B(n1707), .Z(n1693) );
  XNOR U2069 ( .A(n1694), .B(n1693), .Z(n1696) );
  NAND U2070 ( .A(n1642), .B(n1641), .Z(n1646) );
  NAND U2071 ( .A(n1644), .B(n1643), .Z(n1645) );
  NAND U2072 ( .A(n1646), .B(n1645), .Z(n1700) );
  NANDN U2073 ( .A(n1648), .B(n1647), .Z(n1652) );
  NANDN U2074 ( .A(n1650), .B(n1649), .Z(n1651) );
  NAND U2075 ( .A(n1652), .B(n1651), .Z(n1699) );
  XOR U2076 ( .A(n1700), .B(n1699), .Z(n1702) );
  NANDN U2077 ( .A(n1654), .B(n1653), .Z(n1658) );
  OR U2078 ( .A(n1656), .B(n1655), .Z(n1657) );
  NAND U2079 ( .A(n1658), .B(n1657), .Z(n1701) );
  XOR U2080 ( .A(n1702), .B(n1701), .Z(n1695) );
  XOR U2081 ( .A(n1696), .B(n1695), .Z(n1776) );
  NANDN U2082 ( .A(n1660), .B(n1659), .Z(n1664) );
  OR U2083 ( .A(n1662), .B(n1661), .Z(n1663) );
  NAND U2084 ( .A(n1664), .B(n1663), .Z(n1775) );
  XNOR U2085 ( .A(n1776), .B(n1775), .Z(n1777) );
  NANDN U2086 ( .A(n1666), .B(n1665), .Z(n1670) );
  NANDN U2087 ( .A(n1668), .B(n1667), .Z(n1669) );
  NAND U2088 ( .A(n1670), .B(n1669), .Z(n1778) );
  XNOR U2089 ( .A(n1777), .B(n1778), .Z(n1687) );
  NANDN U2090 ( .A(n1672), .B(n1671), .Z(n1676) );
  NAND U2091 ( .A(n1674), .B(n1673), .Z(n1675) );
  NAND U2092 ( .A(n1676), .B(n1675), .Z(n1688) );
  XOR U2093 ( .A(n1687), .B(n1688), .Z(n1690) );
  XOR U2094 ( .A(n1689), .B(n1690), .Z(n1682) );
  XNOR U2095 ( .A(n1682), .B(sreg[53]), .Z(n1684) );
  NANDN U2096 ( .A(sreg[52]), .B(n1677), .Z(n1681) );
  NAND U2097 ( .A(n1679), .B(n1678), .Z(n1680) );
  AND U2098 ( .A(n1681), .B(n1680), .Z(n1683) );
  XOR U2099 ( .A(n1684), .B(n1683), .Z(c[53]) );
  NANDN U2100 ( .A(n1682), .B(sreg[53]), .Z(n1686) );
  NAND U2101 ( .A(n1684), .B(n1683), .Z(n1685) );
  AND U2102 ( .A(n1686), .B(n1685), .Z(n1885) );
  XNOR U2103 ( .A(sreg[54]), .B(n1885), .Z(n1887) );
  NANDN U2104 ( .A(n1688), .B(n1687), .Z(n1692) );
  OR U2105 ( .A(n1690), .B(n1689), .Z(n1691) );
  AND U2106 ( .A(n1692), .B(n1691), .Z(n1784) );
  NANDN U2107 ( .A(n1694), .B(n1693), .Z(n1698) );
  NAND U2108 ( .A(n1696), .B(n1695), .Z(n1697) );
  AND U2109 ( .A(n1698), .B(n1697), .Z(n1880) );
  NAND U2110 ( .A(n1700), .B(n1699), .Z(n1704) );
  NAND U2111 ( .A(n1702), .B(n1701), .Z(n1703) );
  NAND U2112 ( .A(n1704), .B(n1703), .Z(n1879) );
  XNOR U2113 ( .A(n1880), .B(n1879), .Z(n1882) );
  NAND U2114 ( .A(n1710), .B(n1709), .Z(n1714) );
  NAND U2115 ( .A(n1712), .B(n1711), .Z(n1713) );
  NAND U2116 ( .A(n1714), .B(n1713), .Z(n1787) );
  XNOR U2117 ( .A(n1788), .B(n1787), .Z(n1789) );
  NANDN U2118 ( .A(n1716), .B(n1715), .Z(n1720) );
  NANDN U2119 ( .A(n1718), .B(n1717), .Z(n1719) );
  AND U2120 ( .A(n1720), .B(n1719), .Z(n1794) );
  NANDN U2121 ( .A(n1722), .B(n1721), .Z(n1726) );
  NANDN U2122 ( .A(n1724), .B(n1723), .Z(n1725) );
  AND U2123 ( .A(n1726), .B(n1725), .Z(n1801) );
  NAND U2124 ( .A(n568), .B(n1727), .Z(n1729) );
  XOR U2125 ( .A(b[3]), .B(a[20]), .Z(n1822) );
  NAND U2126 ( .A(n7245), .B(n1822), .Z(n1728) );
  AND U2127 ( .A(n1729), .B(n1728), .Z(n1862) );
  NAND U2128 ( .A(n572), .B(n1730), .Z(n1732) );
  XOR U2129 ( .A(b[13]), .B(a[10]), .Z(n1836) );
  NAND U2130 ( .A(n8585), .B(n1836), .Z(n1731) );
  NAND U2131 ( .A(n1732), .B(n1731), .Z(n1861) );
  XNOR U2132 ( .A(n1862), .B(n1861), .Z(n1864) );
  NOR U2133 ( .A(n1734), .B(n1733), .Z(n1863) );
  XOR U2134 ( .A(n1864), .B(n1863), .Z(n1800) );
  NAND U2135 ( .A(b[0]), .B(a[22]), .Z(n1735) );
  XNOR U2136 ( .A(b[1]), .B(n1735), .Z(n1737) );
  NANDN U2137 ( .A(b[0]), .B(a[21]), .Z(n1736) );
  NAND U2138 ( .A(n1737), .B(n1736), .Z(n1819) );
  XNOR U2139 ( .A(b[22]), .B(b[21]), .Z(n9605) );
  IV U2140 ( .A(n9605), .Z(n9268) );
  AND U2141 ( .A(a[0]), .B(n9268), .Z(n1829) );
  NAND U2142 ( .A(n9046), .B(n1738), .Z(n1740) );
  XOR U2143 ( .A(b[19]), .B(a[4]), .Z(n1833) );
  NAND U2144 ( .A(n575), .B(n1833), .Z(n1739) );
  AND U2145 ( .A(n1740), .B(n1739), .Z(n1817) );
  XOR U2146 ( .A(n1829), .B(n1817), .Z(n1818) );
  XNOR U2147 ( .A(n1819), .B(n1818), .Z(n1799) );
  XOR U2148 ( .A(n1800), .B(n1799), .Z(n1802) );
  XNOR U2149 ( .A(n1801), .B(n1802), .Z(n1793) );
  XNOR U2150 ( .A(n1794), .B(n1793), .Z(n1795) );
  NAND U2151 ( .A(n569), .B(n1741), .Z(n1743) );
  XOR U2152 ( .A(b[7]), .B(a[16]), .Z(n1852) );
  NAND U2153 ( .A(n7819), .B(n1852), .Z(n1742) );
  AND U2154 ( .A(n1743), .B(n1742), .Z(n1875) );
  NAND U2155 ( .A(n567), .B(n1744), .Z(n1746) );
  XOR U2156 ( .A(b[5]), .B(a[18]), .Z(n1858) );
  NAND U2157 ( .A(n7235), .B(n1858), .Z(n1745) );
  AND U2158 ( .A(n1746), .B(n1745), .Z(n1874) );
  NAND U2159 ( .A(n573), .B(n1747), .Z(n1749) );
  XOR U2160 ( .A(b[15]), .B(a[8]), .Z(n1825) );
  NAND U2161 ( .A(n8694), .B(n1825), .Z(n1748) );
  NAND U2162 ( .A(n1749), .B(n1748), .Z(n1873) );
  XOR U2163 ( .A(n1874), .B(n1873), .Z(n1876) );
  XOR U2164 ( .A(n1875), .B(n1876), .Z(n1813) );
  NAND U2165 ( .A(n576), .B(n1750), .Z(n1752) );
  XOR U2166 ( .A(b[17]), .B(a[6]), .Z(n1830) );
  NAND U2167 ( .A(n9141), .B(n1830), .Z(n1751) );
  AND U2168 ( .A(n1752), .B(n1751), .Z(n1869) );
  NAND U2169 ( .A(n577), .B(n1754), .Z(n1756) );
  XOR U2170 ( .A(b[21]), .B(a[2]), .Z(n1845) );
  NAND U2171 ( .A(n9216), .B(n1845), .Z(n1755) );
  AND U2172 ( .A(n1756), .B(n1755), .Z(n1868) );
  NAND U2173 ( .A(n570), .B(n1757), .Z(n1759) );
  XOR U2174 ( .A(b[9]), .B(a[14]), .Z(n1855) );
  NAND U2175 ( .A(n8037), .B(n1855), .Z(n1758) );
  NAND U2176 ( .A(n1759), .B(n1758), .Z(n1867) );
  XOR U2177 ( .A(n1868), .B(n1867), .Z(n1870) );
  XOR U2178 ( .A(n1869), .B(n1870), .Z(n1812) );
  OR U2179 ( .A(n1760), .B(n562), .Z(n1762) );
  XNOR U2180 ( .A(b[11]), .B(a[12]), .Z(n1842) );
  OR U2181 ( .A(n1842), .B(n8701), .Z(n1761) );
  AND U2182 ( .A(n1762), .B(n1761), .Z(n1811) );
  XOR U2183 ( .A(n1812), .B(n1811), .Z(n1814) );
  XOR U2184 ( .A(n1813), .B(n1814), .Z(n1808) );
  NANDN U2185 ( .A(n1764), .B(n1763), .Z(n1768) );
  NANDN U2186 ( .A(n1766), .B(n1765), .Z(n1767) );
  AND U2187 ( .A(n1768), .B(n1767), .Z(n1806) );
  NANDN U2188 ( .A(n1770), .B(n1769), .Z(n1774) );
  NANDN U2189 ( .A(n1772), .B(n1771), .Z(n1773) );
  NAND U2190 ( .A(n1774), .B(n1773), .Z(n1805) );
  XNOR U2191 ( .A(n1806), .B(n1805), .Z(n1807) );
  XOR U2192 ( .A(n1808), .B(n1807), .Z(n1796) );
  XOR U2193 ( .A(n1795), .B(n1796), .Z(n1790) );
  XNOR U2194 ( .A(n1789), .B(n1790), .Z(n1881) );
  XOR U2195 ( .A(n1882), .B(n1881), .Z(n1782) );
  NANDN U2196 ( .A(n1776), .B(n1775), .Z(n1780) );
  NANDN U2197 ( .A(n1778), .B(n1777), .Z(n1779) );
  NAND U2198 ( .A(n1780), .B(n1779), .Z(n1781) );
  XNOR U2199 ( .A(n1782), .B(n1781), .Z(n1783) );
  XNOR U2200 ( .A(n1784), .B(n1783), .Z(n1886) );
  XNOR U2201 ( .A(n1887), .B(n1886), .Z(c[54]) );
  NANDN U2202 ( .A(n1782), .B(n1781), .Z(n1786) );
  NANDN U2203 ( .A(n1784), .B(n1783), .Z(n1785) );
  AND U2204 ( .A(n1786), .B(n1785), .Z(n1898) );
  NANDN U2205 ( .A(n1788), .B(n1787), .Z(n1792) );
  NANDN U2206 ( .A(n1790), .B(n1789), .Z(n1791) );
  AND U2207 ( .A(n1792), .B(n1791), .Z(n1996) );
  NANDN U2208 ( .A(n1794), .B(n1793), .Z(n1798) );
  NANDN U2209 ( .A(n1796), .B(n1795), .Z(n1797) );
  AND U2210 ( .A(n1798), .B(n1797), .Z(n1904) );
  NANDN U2211 ( .A(n1800), .B(n1799), .Z(n1804) );
  OR U2212 ( .A(n1802), .B(n1801), .Z(n1803) );
  AND U2213 ( .A(n1804), .B(n1803), .Z(n1902) );
  NANDN U2214 ( .A(n1806), .B(n1805), .Z(n1810) );
  NANDN U2215 ( .A(n1808), .B(n1807), .Z(n1809) );
  AND U2216 ( .A(n1810), .B(n1809), .Z(n1901) );
  XNOR U2217 ( .A(n1902), .B(n1901), .Z(n1903) );
  XOR U2218 ( .A(n1904), .B(n1903), .Z(n1995) );
  NANDN U2219 ( .A(n1812), .B(n1811), .Z(n1816) );
  OR U2220 ( .A(n1814), .B(n1813), .Z(n1815) );
  AND U2221 ( .A(n1816), .B(n1815), .Z(n1907) );
  NANDN U2222 ( .A(n1817), .B(n1829), .Z(n1821) );
  OR U2223 ( .A(n1819), .B(n1818), .Z(n1820) );
  AND U2224 ( .A(n1821), .B(n1820), .Z(n1991) );
  NAND U2225 ( .A(n568), .B(n1822), .Z(n1824) );
  XOR U2226 ( .A(b[3]), .B(a[21]), .Z(n1930) );
  NAND U2227 ( .A(n7245), .B(n1930), .Z(n1823) );
  AND U2228 ( .A(n1824), .B(n1823), .Z(n1942) );
  NAND U2229 ( .A(n573), .B(n1825), .Z(n1827) );
  XOR U2230 ( .A(b[15]), .B(a[9]), .Z(n1966) );
  NAND U2231 ( .A(n8694), .B(n1966), .Z(n1826) );
  AND U2232 ( .A(n1827), .B(n1826), .Z(n1940) );
  NANDN U2233 ( .A(b[22]), .B(b[23]), .Z(n1828) );
  NAND U2234 ( .A(n9268), .B(b[23]), .Z(n9646) );
  NAND U2235 ( .A(n1828), .B(n9646), .Z(n9690) );
  IV U2236 ( .A(n9690), .Z(n9724) );
  NOR U2237 ( .A(n9724), .B(n1829), .Z(n1939) );
  XNOR U2238 ( .A(n1940), .B(n1939), .Z(n1941) );
  XNOR U2239 ( .A(n1942), .B(n1941), .Z(n1988) );
  NAND U2240 ( .A(n576), .B(n1830), .Z(n1832) );
  XOR U2241 ( .A(b[17]), .B(a[7]), .Z(n1963) );
  NAND U2242 ( .A(n9141), .B(n1963), .Z(n1831) );
  AND U2243 ( .A(n1832), .B(n1831), .Z(n1922) );
  NAND U2244 ( .A(n9046), .B(n1833), .Z(n1835) );
  XOR U2245 ( .A(b[19]), .B(a[5]), .Z(n1975) );
  NAND U2246 ( .A(n575), .B(n1975), .Z(n1834) );
  AND U2247 ( .A(n1835), .B(n1834), .Z(n1920) );
  NAND U2248 ( .A(n572), .B(n1836), .Z(n1838) );
  XOR U2249 ( .A(b[13]), .B(a[11]), .Z(n1927) );
  NAND U2250 ( .A(n8585), .B(n1927), .Z(n1837) );
  NAND U2251 ( .A(n1838), .B(n1837), .Z(n1919) );
  XNOR U2252 ( .A(n1920), .B(n1919), .Z(n1921) );
  XOR U2253 ( .A(n1922), .B(n1921), .Z(n1989) );
  XNOR U2254 ( .A(n1988), .B(n1989), .Z(n1990) );
  XOR U2255 ( .A(n1991), .B(n1990), .Z(n1908) );
  XNOR U2256 ( .A(n1907), .B(n1908), .Z(n1909) );
  NAND U2257 ( .A(b[0]), .B(a[23]), .Z(n1839) );
  XNOR U2258 ( .A(b[1]), .B(n1839), .Z(n1841) );
  NANDN U2259 ( .A(b[0]), .B(a[22]), .Z(n1840) );
  NAND U2260 ( .A(n1841), .B(n1840), .Z(n1934) );
  OR U2261 ( .A(n1842), .B(n562), .Z(n1844) );
  XOR U2262 ( .A(b[11]), .B(a[13]), .Z(n1969) );
  NAND U2263 ( .A(n8135), .B(n1969), .Z(n1843) );
  NAND U2264 ( .A(n1844), .B(n1843), .Z(n1933) );
  XNOR U2265 ( .A(n1934), .B(n1933), .Z(n1935) );
  NAND U2266 ( .A(n577), .B(n1845), .Z(n1847) );
  XOR U2267 ( .A(b[21]), .B(a[3]), .Z(n1951) );
  NAND U2268 ( .A(n9216), .B(n1951), .Z(n1846) );
  AND U2269 ( .A(n1847), .B(n1846), .Z(n1925) );
  XOR U2270 ( .A(b[23]), .B(b[22]), .Z(n1978) );
  XOR U2271 ( .A(b[23]), .B(a[0]), .Z(n1848) );
  NAND U2272 ( .A(n1978), .B(n1848), .Z(n1849) );
  NANDN U2273 ( .A(n1849), .B(n9605), .Z(n1851) );
  XOR U2274 ( .A(b[23]), .B(a[1]), .Z(n1979) );
  NANDN U2275 ( .A(n9605), .B(n1979), .Z(n1850) );
  NAND U2276 ( .A(n1851), .B(n1850), .Z(n1926) );
  XOR U2277 ( .A(n1925), .B(n1926), .Z(n1936) );
  XNOR U2278 ( .A(n1935), .B(n1936), .Z(n1983) );
  NAND U2279 ( .A(n569), .B(n1852), .Z(n1854) );
  XOR U2280 ( .A(b[7]), .B(a[17]), .Z(n1957) );
  NAND U2281 ( .A(n7819), .B(n1957), .Z(n1853) );
  AND U2282 ( .A(n1854), .B(n1853), .Z(n1947) );
  NAND U2283 ( .A(n570), .B(n1855), .Z(n1857) );
  XOR U2284 ( .A(b[9]), .B(a[15]), .Z(n1972) );
  NAND U2285 ( .A(n8037), .B(n1972), .Z(n1856) );
  AND U2286 ( .A(n1857), .B(n1856), .Z(n1946) );
  NAND U2287 ( .A(n567), .B(n1858), .Z(n1860) );
  XOR U2288 ( .A(b[5]), .B(a[19]), .Z(n1960) );
  NAND U2289 ( .A(n7235), .B(n1960), .Z(n1859) );
  NAND U2290 ( .A(n1860), .B(n1859), .Z(n1945) );
  XOR U2291 ( .A(n1946), .B(n1945), .Z(n1948) );
  XOR U2292 ( .A(n1947), .B(n1948), .Z(n1982) );
  XOR U2293 ( .A(n1983), .B(n1982), .Z(n1985) );
  NANDN U2294 ( .A(n1862), .B(n1861), .Z(n1866) );
  NAND U2295 ( .A(n1864), .B(n1863), .Z(n1865) );
  NAND U2296 ( .A(n1866), .B(n1865), .Z(n1984) );
  XOR U2297 ( .A(n1985), .B(n1984), .Z(n1915) );
  NANDN U2298 ( .A(n1868), .B(n1867), .Z(n1872) );
  OR U2299 ( .A(n1870), .B(n1869), .Z(n1871) );
  AND U2300 ( .A(n1872), .B(n1871), .Z(n1914) );
  NANDN U2301 ( .A(n1874), .B(n1873), .Z(n1878) );
  OR U2302 ( .A(n1876), .B(n1875), .Z(n1877) );
  NAND U2303 ( .A(n1878), .B(n1877), .Z(n1913) );
  XOR U2304 ( .A(n1914), .B(n1913), .Z(n1916) );
  XOR U2305 ( .A(n1915), .B(n1916), .Z(n1910) );
  XNOR U2306 ( .A(n1909), .B(n1910), .Z(n1994) );
  XOR U2307 ( .A(n1995), .B(n1994), .Z(n1997) );
  XOR U2308 ( .A(n1996), .B(n1997), .Z(n1896) );
  NANDN U2309 ( .A(n1880), .B(n1879), .Z(n1884) );
  NAND U2310 ( .A(n1882), .B(n1881), .Z(n1883) );
  AND U2311 ( .A(n1884), .B(n1883), .Z(n1895) );
  XNOR U2312 ( .A(n1896), .B(n1895), .Z(n1897) );
  XNOR U2313 ( .A(n1898), .B(n1897), .Z(n1890) );
  XNOR U2314 ( .A(sreg[55]), .B(n1890), .Z(n1892) );
  NANDN U2315 ( .A(sreg[54]), .B(n1885), .Z(n1889) );
  NAND U2316 ( .A(n1887), .B(n1886), .Z(n1888) );
  NAND U2317 ( .A(n1889), .B(n1888), .Z(n1891) );
  XNOR U2318 ( .A(n1892), .B(n1891), .Z(c[55]) );
  NANDN U2319 ( .A(sreg[55]), .B(n1890), .Z(n1894) );
  NAND U2320 ( .A(n1892), .B(n1891), .Z(n1893) );
  NAND U2321 ( .A(n1894), .B(n1893), .Z(n2109) );
  XNOR U2322 ( .A(sreg[56]), .B(n2109), .Z(n2111) );
  NANDN U2323 ( .A(n1896), .B(n1895), .Z(n1900) );
  NANDN U2324 ( .A(n1898), .B(n1897), .Z(n1899) );
  AND U2325 ( .A(n1900), .B(n1899), .Z(n2003) );
  NANDN U2326 ( .A(n1902), .B(n1901), .Z(n1906) );
  NAND U2327 ( .A(n1904), .B(n1903), .Z(n1905) );
  AND U2328 ( .A(n1906), .B(n1905), .Z(n2009) );
  NANDN U2329 ( .A(n1908), .B(n1907), .Z(n1912) );
  NANDN U2330 ( .A(n1910), .B(n1909), .Z(n1911) );
  AND U2331 ( .A(n1912), .B(n1911), .Z(n2006) );
  NANDN U2332 ( .A(n1914), .B(n1913), .Z(n1918) );
  NANDN U2333 ( .A(n1916), .B(n1915), .Z(n1917) );
  AND U2334 ( .A(n1918), .B(n1917), .Z(n2105) );
  NANDN U2335 ( .A(n1920), .B(n1919), .Z(n1924) );
  NANDN U2336 ( .A(n1922), .B(n1921), .Z(n1923) );
  AND U2337 ( .A(n1924), .B(n1923), .Z(n2022) );
  ANDN U2338 ( .B(n1926), .A(n1925), .Z(n2063) );
  NANDN U2339 ( .A(n553), .B(n1927), .Z(n1929) );
  XNOR U2340 ( .A(b[13]), .B(a[12]), .Z(n2049) );
  OR U2341 ( .A(n2049), .B(n8853), .Z(n1928) );
  AND U2342 ( .A(n1929), .B(n1928), .Z(n2060) );
  NANDN U2343 ( .A(n560), .B(n1930), .Z(n1932) );
  XNOR U2344 ( .A(b[3]), .B(a[22]), .Z(n2052) );
  OR U2345 ( .A(n2052), .B(n7784), .Z(n1931) );
  NAND U2346 ( .A(n1932), .B(n1931), .Z(n2061) );
  XNOR U2347 ( .A(n2060), .B(n2061), .Z(n2062) );
  XOR U2348 ( .A(n2063), .B(n2062), .Z(n2023) );
  XNOR U2349 ( .A(n2022), .B(n2023), .Z(n2025) );
  NANDN U2350 ( .A(n1934), .B(n1933), .Z(n1938) );
  NANDN U2351 ( .A(n1936), .B(n1935), .Z(n1937) );
  AND U2352 ( .A(n1938), .B(n1937), .Z(n2024) );
  XOR U2353 ( .A(n2025), .B(n2024), .Z(n2104) );
  NANDN U2354 ( .A(n1940), .B(n1939), .Z(n1944) );
  NANDN U2355 ( .A(n1942), .B(n1941), .Z(n1943) );
  AND U2356 ( .A(n1944), .B(n1943), .Z(n2019) );
  NANDN U2357 ( .A(n1946), .B(n1945), .Z(n1950) );
  OR U2358 ( .A(n1948), .B(n1947), .Z(n1949) );
  NAND U2359 ( .A(n1950), .B(n1949), .Z(n2018) );
  XNOR U2360 ( .A(n2019), .B(n2018), .Z(n2021) );
  XNOR U2361 ( .A(b[24]), .B(b[23]), .Z(n9684) );
  IV U2362 ( .A(n9684), .Z(n9364) );
  AND U2363 ( .A(a[0]), .B(n9364), .Z(n2059) );
  NAND U2364 ( .A(n577), .B(n1951), .Z(n1953) );
  XOR U2365 ( .A(b[21]), .B(a[4]), .Z(n2094) );
  NAND U2366 ( .A(n9216), .B(n2094), .Z(n1952) );
  AND U2367 ( .A(n1953), .B(n1952), .Z(n2034) );
  XNOR U2368 ( .A(n2059), .B(n2034), .Z(n2035) );
  NAND U2369 ( .A(b[0]), .B(a[24]), .Z(n1954) );
  XNOR U2370 ( .A(b[1]), .B(n1954), .Z(n1956) );
  NANDN U2371 ( .A(b[0]), .B(a[23]), .Z(n1955) );
  NAND U2372 ( .A(n1956), .B(n1955), .Z(n2036) );
  XNOR U2373 ( .A(n2035), .B(n2036), .Z(n2028) );
  NAND U2374 ( .A(n569), .B(n1957), .Z(n1959) );
  XOR U2375 ( .A(b[7]), .B(a[18]), .Z(n2082) );
  NAND U2376 ( .A(n7819), .B(n2082), .Z(n1958) );
  AND U2377 ( .A(n1959), .B(n1958), .Z(n2079) );
  NAND U2378 ( .A(n567), .B(n1960), .Z(n1962) );
  XOR U2379 ( .A(b[5]), .B(a[20]), .Z(n2085) );
  NAND U2380 ( .A(n7235), .B(n2085), .Z(n1961) );
  AND U2381 ( .A(n1962), .B(n1961), .Z(n2077) );
  NAND U2382 ( .A(n576), .B(n1963), .Z(n1965) );
  XOR U2383 ( .A(b[17]), .B(a[8]), .Z(n2088) );
  NAND U2384 ( .A(n9141), .B(n2088), .Z(n1964) );
  NAND U2385 ( .A(n1965), .B(n1964), .Z(n2076) );
  XNOR U2386 ( .A(n2077), .B(n2076), .Z(n2078) );
  XOR U2387 ( .A(n2079), .B(n2078), .Z(n2029) );
  XNOR U2388 ( .A(n2028), .B(n2029), .Z(n2030) );
  NAND U2389 ( .A(n573), .B(n1966), .Z(n1968) );
  XOR U2390 ( .A(b[15]), .B(a[10]), .Z(n2055) );
  NAND U2391 ( .A(n8694), .B(n2055), .Z(n1967) );
  AND U2392 ( .A(n1968), .B(n1967), .Z(n2073) );
  NAND U2393 ( .A(n571), .B(n1969), .Z(n1971) );
  XOR U2394 ( .A(b[11]), .B(a[14]), .Z(n2100) );
  NAND U2395 ( .A(n8135), .B(n2100), .Z(n1970) );
  NAND U2396 ( .A(n1971), .B(n1970), .Z(n2072) );
  XNOR U2397 ( .A(n2073), .B(n2072), .Z(n2075) );
  NANDN U2398 ( .A(n564), .B(n1972), .Z(n1974) );
  XNOR U2399 ( .A(b[9]), .B(a[16]), .Z(n2097) );
  OR U2400 ( .A(n2097), .B(n8485), .Z(n1973) );
  NAND U2401 ( .A(n1974), .B(n1973), .Z(n2068) );
  NANDN U2402 ( .A(n574), .B(n1975), .Z(n1977) );
  XNOR U2403 ( .A(b[19]), .B(a[6]), .Z(n2091) );
  OR U2404 ( .A(n2091), .B(n555), .Z(n1976) );
  NAND U2405 ( .A(n1977), .B(n1976), .Z(n2067) );
  NAND U2406 ( .A(n578), .B(n1979), .Z(n1981) );
  XOR U2407 ( .A(b[23]), .B(a[2]), .Z(n2039) );
  NAND U2408 ( .A(n9268), .B(n2039), .Z(n1980) );
  NAND U2409 ( .A(n1981), .B(n1980), .Z(n2066) );
  XOR U2410 ( .A(n2067), .B(n2066), .Z(n2069) );
  XNOR U2411 ( .A(n2068), .B(n2069), .Z(n2074) );
  XNOR U2412 ( .A(n2075), .B(n2074), .Z(n2031) );
  XNOR U2413 ( .A(n2030), .B(n2031), .Z(n2020) );
  XNOR U2414 ( .A(n2021), .B(n2020), .Z(n2103) );
  XOR U2415 ( .A(n2104), .B(n2103), .Z(n2106) );
  XOR U2416 ( .A(n2105), .B(n2106), .Z(n2015) );
  NAND U2417 ( .A(n1983), .B(n1982), .Z(n1987) );
  NAND U2418 ( .A(n1985), .B(n1984), .Z(n1986) );
  AND U2419 ( .A(n1987), .B(n1986), .Z(n2012) );
  NANDN U2420 ( .A(n1989), .B(n1988), .Z(n1993) );
  NANDN U2421 ( .A(n1991), .B(n1990), .Z(n1992) );
  NAND U2422 ( .A(n1993), .B(n1992), .Z(n2013) );
  XNOR U2423 ( .A(n2012), .B(n2013), .Z(n2014) );
  XOR U2424 ( .A(n2015), .B(n2014), .Z(n2007) );
  XNOR U2425 ( .A(n2006), .B(n2007), .Z(n2008) );
  XNOR U2426 ( .A(n2009), .B(n2008), .Z(n2000) );
  NANDN U2427 ( .A(n1995), .B(n1994), .Z(n1999) );
  OR U2428 ( .A(n1997), .B(n1996), .Z(n1998) );
  NAND U2429 ( .A(n1999), .B(n1998), .Z(n2001) );
  XNOR U2430 ( .A(n2000), .B(n2001), .Z(n2002) );
  XNOR U2431 ( .A(n2003), .B(n2002), .Z(n2110) );
  XNOR U2432 ( .A(n2111), .B(n2110), .Z(c[56]) );
  NANDN U2433 ( .A(n2001), .B(n2000), .Z(n2005) );
  NANDN U2434 ( .A(n2003), .B(n2002), .Z(n2004) );
  AND U2435 ( .A(n2005), .B(n2004), .Z(n2122) );
  NANDN U2436 ( .A(n2007), .B(n2006), .Z(n2011) );
  NANDN U2437 ( .A(n2009), .B(n2008), .Z(n2010) );
  AND U2438 ( .A(n2011), .B(n2010), .Z(n2120) );
  NANDN U2439 ( .A(n2013), .B(n2012), .Z(n2017) );
  NANDN U2440 ( .A(n2015), .B(n2014), .Z(n2016) );
  AND U2441 ( .A(n2017), .B(n2016), .Z(n2128) );
  NANDN U2442 ( .A(n2023), .B(n2022), .Z(n2027) );
  NAND U2443 ( .A(n2025), .B(n2024), .Z(n2026) );
  AND U2444 ( .A(n2027), .B(n2026), .Z(n2137) );
  XNOR U2445 ( .A(n2138), .B(n2137), .Z(n2140) );
  NANDN U2446 ( .A(n2029), .B(n2028), .Z(n2033) );
  NAND U2447 ( .A(n2031), .B(n2030), .Z(n2032) );
  AND U2448 ( .A(n2033), .B(n2032), .Z(n2132) );
  NANDN U2449 ( .A(n2034), .B(n2059), .Z(n2038) );
  NANDN U2450 ( .A(n2036), .B(n2035), .Z(n2037) );
  AND U2451 ( .A(n2038), .B(n2037), .Z(n2145) );
  NAND U2452 ( .A(n578), .B(n2039), .Z(n2041) );
  XOR U2453 ( .A(b[23]), .B(a[3]), .Z(n2180) );
  NAND U2454 ( .A(n9268), .B(n2180), .Z(n2040) );
  AND U2455 ( .A(n2041), .B(n2040), .Z(n2198) );
  XOR U2456 ( .A(b[25]), .B(b[24]), .Z(n2158) );
  XOR U2457 ( .A(b[25]), .B(a[0]), .Z(n2042) );
  NAND U2458 ( .A(n2158), .B(n2042), .Z(n2043) );
  NANDN U2459 ( .A(n2043), .B(n9684), .Z(n2045) );
  XOR U2460 ( .A(b[25]), .B(a[1]), .Z(n2159) );
  NANDN U2461 ( .A(n9684), .B(n2159), .Z(n2044) );
  AND U2462 ( .A(n2045), .B(n2044), .Z(n2199) );
  XOR U2463 ( .A(n2198), .B(n2199), .Z(n2151) );
  NAND U2464 ( .A(b[0]), .B(a[25]), .Z(n2046) );
  XNOR U2465 ( .A(b[1]), .B(n2046), .Z(n2048) );
  NANDN U2466 ( .A(b[0]), .B(a[24]), .Z(n2047) );
  NAND U2467 ( .A(n2048), .B(n2047), .Z(n2149) );
  OR U2468 ( .A(n2049), .B(n553), .Z(n2051) );
  XNOR U2469 ( .A(b[13]), .B(a[13]), .Z(n2206) );
  OR U2470 ( .A(n2206), .B(n8853), .Z(n2050) );
  NAND U2471 ( .A(n2051), .B(n2050), .Z(n2150) );
  XOR U2472 ( .A(n2149), .B(n2150), .Z(n2152) );
  XOR U2473 ( .A(n2151), .B(n2152), .Z(n2144) );
  OR U2474 ( .A(n2052), .B(n560), .Z(n2054) );
  XOR U2475 ( .A(b[3]), .B(a[23]), .Z(n2203) );
  NAND U2476 ( .A(n7245), .B(n2203), .Z(n2053) );
  AND U2477 ( .A(n2054), .B(n2053), .Z(n2168) );
  NAND U2478 ( .A(n573), .B(n2055), .Z(n2057) );
  XOR U2479 ( .A(b[15]), .B(a[11]), .Z(n2200) );
  NAND U2480 ( .A(n8694), .B(n2200), .Z(n2056) );
  AND U2481 ( .A(n2057), .B(n2056), .Z(n2166) );
  NANDN U2482 ( .A(b[24]), .B(b[25]), .Z(n2058) );
  NAND U2483 ( .A(n9364), .B(b[25]), .Z(n9740) );
  NAND U2484 ( .A(n2058), .B(n9740), .Z(n9768) );
  IV U2485 ( .A(n9768), .Z(n9800) );
  NOR U2486 ( .A(n9800), .B(n2059), .Z(n2165) );
  XNOR U2487 ( .A(n2166), .B(n2165), .Z(n2167) );
  XNOR U2488 ( .A(n2168), .B(n2167), .Z(n2143) );
  XOR U2489 ( .A(n2144), .B(n2143), .Z(n2146) );
  XOR U2490 ( .A(n2145), .B(n2146), .Z(n2223) );
  NANDN U2491 ( .A(n2061), .B(n2060), .Z(n2065) );
  NANDN U2492 ( .A(n2063), .B(n2062), .Z(n2064) );
  AND U2493 ( .A(n2065), .B(n2064), .Z(n2222) );
  NAND U2494 ( .A(n2067), .B(n2066), .Z(n2071) );
  NAND U2495 ( .A(n2069), .B(n2068), .Z(n2070) );
  AND U2496 ( .A(n2071), .B(n2070), .Z(n2221) );
  XOR U2497 ( .A(n2222), .B(n2221), .Z(n2224) );
  XNOR U2498 ( .A(n2223), .B(n2224), .Z(n2131) );
  XNOR U2499 ( .A(n2132), .B(n2131), .Z(n2133) );
  NANDN U2500 ( .A(n2077), .B(n2076), .Z(n2081) );
  NANDN U2501 ( .A(n2079), .B(n2078), .Z(n2080) );
  AND U2502 ( .A(n2081), .B(n2080), .Z(n2228) );
  NAND U2503 ( .A(n569), .B(n2082), .Z(n2084) );
  XOR U2504 ( .A(b[7]), .B(a[19]), .Z(n2189) );
  NAND U2505 ( .A(n7819), .B(n2189), .Z(n2083) );
  AND U2506 ( .A(n2084), .B(n2083), .Z(n2194) );
  NAND U2507 ( .A(n567), .B(n2085), .Z(n2087) );
  XOR U2508 ( .A(b[5]), .B(a[21]), .Z(n2212) );
  NAND U2509 ( .A(n7235), .B(n2212), .Z(n2086) );
  AND U2510 ( .A(n2087), .B(n2086), .Z(n2193) );
  NAND U2511 ( .A(n576), .B(n2088), .Z(n2090) );
  XOR U2512 ( .A(b[17]), .B(a[9]), .Z(n2162) );
  NAND U2513 ( .A(n9141), .B(n2162), .Z(n2089) );
  NAND U2514 ( .A(n2090), .B(n2089), .Z(n2192) );
  XOR U2515 ( .A(n2193), .B(n2192), .Z(n2195) );
  XOR U2516 ( .A(n2194), .B(n2195), .Z(n2217) );
  OR U2517 ( .A(n2091), .B(n574), .Z(n2093) );
  XOR U2518 ( .A(b[19]), .B(a[7]), .Z(n2209) );
  NAND U2519 ( .A(n575), .B(n2209), .Z(n2092) );
  AND U2520 ( .A(n2093), .B(n2092), .Z(n2173) );
  NAND U2521 ( .A(n577), .B(n2094), .Z(n2096) );
  XOR U2522 ( .A(b[21]), .B(a[5]), .Z(n2155) );
  NAND U2523 ( .A(n9216), .B(n2155), .Z(n2095) );
  AND U2524 ( .A(n2096), .B(n2095), .Z(n2172) );
  OR U2525 ( .A(n2097), .B(n564), .Z(n2099) );
  XOR U2526 ( .A(b[9]), .B(a[17]), .Z(n2183) );
  NAND U2527 ( .A(n8037), .B(n2183), .Z(n2098) );
  NAND U2528 ( .A(n2099), .B(n2098), .Z(n2171) );
  XOR U2529 ( .A(n2172), .B(n2171), .Z(n2174) );
  XOR U2530 ( .A(n2173), .B(n2174), .Z(n2216) );
  NANDN U2531 ( .A(n562), .B(n2100), .Z(n2102) );
  XNOR U2532 ( .A(b[11]), .B(a[15]), .Z(n2186) );
  OR U2533 ( .A(n2186), .B(n8701), .Z(n2101) );
  AND U2534 ( .A(n2102), .B(n2101), .Z(n2215) );
  XOR U2535 ( .A(n2216), .B(n2215), .Z(n2218) );
  XNOR U2536 ( .A(n2217), .B(n2218), .Z(n2227) );
  XNOR U2537 ( .A(n2228), .B(n2227), .Z(n2229) );
  XOR U2538 ( .A(n2230), .B(n2229), .Z(n2134) );
  XNOR U2539 ( .A(n2133), .B(n2134), .Z(n2139) );
  XOR U2540 ( .A(n2140), .B(n2139), .Z(n2126) );
  NANDN U2541 ( .A(n2104), .B(n2103), .Z(n2108) );
  OR U2542 ( .A(n2106), .B(n2105), .Z(n2107) );
  AND U2543 ( .A(n2108), .B(n2107), .Z(n2125) );
  XNOR U2544 ( .A(n2126), .B(n2125), .Z(n2127) );
  XNOR U2545 ( .A(n2128), .B(n2127), .Z(n2119) );
  XNOR U2546 ( .A(n2120), .B(n2119), .Z(n2121) );
  XNOR U2547 ( .A(n2122), .B(n2121), .Z(n2114) );
  XNOR U2548 ( .A(sreg[57]), .B(n2114), .Z(n2116) );
  NANDN U2549 ( .A(sreg[56]), .B(n2109), .Z(n2113) );
  NAND U2550 ( .A(n2111), .B(n2110), .Z(n2112) );
  NAND U2551 ( .A(n2113), .B(n2112), .Z(n2115) );
  XNOR U2552 ( .A(n2116), .B(n2115), .Z(c[57]) );
  NANDN U2553 ( .A(sreg[57]), .B(n2114), .Z(n2118) );
  NAND U2554 ( .A(n2116), .B(n2115), .Z(n2117) );
  NAND U2555 ( .A(n2118), .B(n2117), .Z(n2355) );
  XNOR U2556 ( .A(sreg[58]), .B(n2355), .Z(n2357) );
  NANDN U2557 ( .A(n2120), .B(n2119), .Z(n2124) );
  NANDN U2558 ( .A(n2122), .B(n2121), .Z(n2123) );
  AND U2559 ( .A(n2124), .B(n2123), .Z(n2236) );
  NANDN U2560 ( .A(n2126), .B(n2125), .Z(n2130) );
  NANDN U2561 ( .A(n2128), .B(n2127), .Z(n2129) );
  AND U2562 ( .A(n2130), .B(n2129), .Z(n2234) );
  NANDN U2563 ( .A(n2132), .B(n2131), .Z(n2136) );
  NANDN U2564 ( .A(n2134), .B(n2133), .Z(n2135) );
  AND U2565 ( .A(n2136), .B(n2135), .Z(n2239) );
  NANDN U2566 ( .A(n2138), .B(n2137), .Z(n2142) );
  NAND U2567 ( .A(n2140), .B(n2139), .Z(n2141) );
  NAND U2568 ( .A(n2142), .B(n2141), .Z(n2240) );
  XNOR U2569 ( .A(n2239), .B(n2240), .Z(n2241) );
  NANDN U2570 ( .A(n2144), .B(n2143), .Z(n2148) );
  OR U2571 ( .A(n2146), .B(n2145), .Z(n2147) );
  AND U2572 ( .A(n2148), .B(n2147), .Z(n2258) );
  NANDN U2573 ( .A(n2150), .B(n2149), .Z(n2154) );
  OR U2574 ( .A(n2152), .B(n2151), .Z(n2153) );
  AND U2575 ( .A(n2154), .B(n2153), .Z(n2338) );
  NAND U2576 ( .A(n577), .B(n2155), .Z(n2157) );
  XOR U2577 ( .A(b[21]), .B(a[6]), .Z(n2322) );
  NAND U2578 ( .A(n9216), .B(n2322), .Z(n2156) );
  AND U2579 ( .A(n2157), .B(n2156), .Z(n2293) );
  NAND U2580 ( .A(n579), .B(n2159), .Z(n2161) );
  XOR U2581 ( .A(b[25]), .B(a[2]), .Z(n2269) );
  NAND U2582 ( .A(n9364), .B(n2269), .Z(n2160) );
  AND U2583 ( .A(n2161), .B(n2160), .Z(n2292) );
  NAND U2584 ( .A(n576), .B(n2162), .Z(n2164) );
  XOR U2585 ( .A(b[17]), .B(a[10]), .Z(n2319) );
  NAND U2586 ( .A(n9141), .B(n2319), .Z(n2163) );
  NAND U2587 ( .A(n2164), .B(n2163), .Z(n2291) );
  XOR U2588 ( .A(n2292), .B(n2291), .Z(n2294) );
  XNOR U2589 ( .A(n2293), .B(n2294), .Z(n2337) );
  XNOR U2590 ( .A(n2338), .B(n2337), .Z(n2340) );
  NANDN U2591 ( .A(n2166), .B(n2165), .Z(n2170) );
  NANDN U2592 ( .A(n2168), .B(n2167), .Z(n2169) );
  AND U2593 ( .A(n2170), .B(n2169), .Z(n2339) );
  XNOR U2594 ( .A(n2340), .B(n2339), .Z(n2257) );
  XNOR U2595 ( .A(n2258), .B(n2257), .Z(n2260) );
  NANDN U2596 ( .A(n2172), .B(n2171), .Z(n2176) );
  OR U2597 ( .A(n2174), .B(n2173), .Z(n2175) );
  AND U2598 ( .A(n2176), .B(n2175), .Z(n2346) );
  NAND U2599 ( .A(b[0]), .B(a[26]), .Z(n2177) );
  XNOR U2600 ( .A(b[1]), .B(n2177), .Z(n2179) );
  NANDN U2601 ( .A(b[0]), .B(a[25]), .Z(n2178) );
  NAND U2602 ( .A(n2179), .B(n2178), .Z(n2305) );
  XNOR U2603 ( .A(b[26]), .B(b[25]), .Z(n9692) );
  IV U2604 ( .A(n9692), .Z(n9770) );
  AND U2605 ( .A(a[0]), .B(n9770), .Z(n2315) );
  NAND U2606 ( .A(n578), .B(n2180), .Z(n2182) );
  XOR U2607 ( .A(b[23]), .B(a[4]), .Z(n2325) );
  NAND U2608 ( .A(n9268), .B(n2325), .Z(n2181) );
  AND U2609 ( .A(n2182), .B(n2181), .Z(n2303) );
  XNOR U2610 ( .A(n2315), .B(n2303), .Z(n2304) );
  XNOR U2611 ( .A(n2305), .B(n2304), .Z(n2343) );
  NAND U2612 ( .A(n570), .B(n2183), .Z(n2185) );
  XOR U2613 ( .A(b[9]), .B(a[18]), .Z(n2328) );
  NAND U2614 ( .A(n8037), .B(n2328), .Z(n2184) );
  AND U2615 ( .A(n2185), .B(n2184), .Z(n2300) );
  OR U2616 ( .A(n2186), .B(n562), .Z(n2188) );
  XOR U2617 ( .A(b[11]), .B(a[16]), .Z(n2316) );
  NAND U2618 ( .A(n8135), .B(n2316), .Z(n2187) );
  AND U2619 ( .A(n2188), .B(n2187), .Z(n2298) );
  NAND U2620 ( .A(n569), .B(n2189), .Z(n2191) );
  XOR U2621 ( .A(b[7]), .B(a[20]), .Z(n2276) );
  NAND U2622 ( .A(n7819), .B(n2276), .Z(n2190) );
  NAND U2623 ( .A(n2191), .B(n2190), .Z(n2297) );
  XNOR U2624 ( .A(n2298), .B(n2297), .Z(n2299) );
  XOR U2625 ( .A(n2300), .B(n2299), .Z(n2344) );
  XNOR U2626 ( .A(n2343), .B(n2344), .Z(n2345) );
  XNOR U2627 ( .A(n2346), .B(n2345), .Z(n2252) );
  NANDN U2628 ( .A(n2193), .B(n2192), .Z(n2197) );
  OR U2629 ( .A(n2195), .B(n2194), .Z(n2196) );
  AND U2630 ( .A(n2197), .B(n2196), .Z(n2351) );
  NOR U2631 ( .A(n2199), .B(n2198), .Z(n2287) );
  NANDN U2632 ( .A(n557), .B(n2200), .Z(n2202) );
  XNOR U2633 ( .A(b[15]), .B(a[12]), .Z(n2311) );
  OR U2634 ( .A(n2311), .B(n9067), .Z(n2201) );
  AND U2635 ( .A(n2202), .B(n2201), .Z(n2285) );
  NANDN U2636 ( .A(n560), .B(n2203), .Z(n2205) );
  XNOR U2637 ( .A(b[3]), .B(a[24]), .Z(n2308) );
  OR U2638 ( .A(n2308), .B(n7784), .Z(n2204) );
  NAND U2639 ( .A(n2205), .B(n2204), .Z(n2286) );
  XOR U2640 ( .A(n2285), .B(n2286), .Z(n2288) );
  XOR U2641 ( .A(n2287), .B(n2288), .Z(n2350) );
  OR U2642 ( .A(n2206), .B(n553), .Z(n2208) );
  XOR U2643 ( .A(b[13]), .B(a[14]), .Z(n2263) );
  NAND U2644 ( .A(n8585), .B(n2263), .Z(n2207) );
  AND U2645 ( .A(n2208), .B(n2207), .Z(n2334) );
  NAND U2646 ( .A(n9046), .B(n2209), .Z(n2211) );
  XOR U2647 ( .A(b[19]), .B(a[8]), .Z(n2282) );
  NAND U2648 ( .A(n575), .B(n2282), .Z(n2210) );
  AND U2649 ( .A(n2211), .B(n2210), .Z(n2332) );
  NAND U2650 ( .A(n567), .B(n2212), .Z(n2214) );
  XOR U2651 ( .A(b[5]), .B(a[22]), .Z(n2279) );
  NAND U2652 ( .A(n7235), .B(n2279), .Z(n2213) );
  NAND U2653 ( .A(n2214), .B(n2213), .Z(n2331) );
  XNOR U2654 ( .A(n2332), .B(n2331), .Z(n2333) );
  XNOR U2655 ( .A(n2334), .B(n2333), .Z(n2349) );
  XOR U2656 ( .A(n2350), .B(n2349), .Z(n2352) );
  XOR U2657 ( .A(n2351), .B(n2352), .Z(n2251) );
  XOR U2658 ( .A(n2252), .B(n2251), .Z(n2254) );
  NANDN U2659 ( .A(n2216), .B(n2215), .Z(n2220) );
  OR U2660 ( .A(n2218), .B(n2217), .Z(n2219) );
  AND U2661 ( .A(n2220), .B(n2219), .Z(n2253) );
  XOR U2662 ( .A(n2254), .B(n2253), .Z(n2259) );
  XOR U2663 ( .A(n2260), .B(n2259), .Z(n2248) );
  NANDN U2664 ( .A(n2222), .B(n2221), .Z(n2226) );
  OR U2665 ( .A(n2224), .B(n2223), .Z(n2225) );
  AND U2666 ( .A(n2226), .B(n2225), .Z(n2246) );
  NANDN U2667 ( .A(n2228), .B(n2227), .Z(n2232) );
  NANDN U2668 ( .A(n2230), .B(n2229), .Z(n2231) );
  AND U2669 ( .A(n2232), .B(n2231), .Z(n2245) );
  XNOR U2670 ( .A(n2246), .B(n2245), .Z(n2247) );
  XOR U2671 ( .A(n2248), .B(n2247), .Z(n2242) );
  XNOR U2672 ( .A(n2241), .B(n2242), .Z(n2233) );
  XNOR U2673 ( .A(n2234), .B(n2233), .Z(n2235) );
  XNOR U2674 ( .A(n2236), .B(n2235), .Z(n2356) );
  XNOR U2675 ( .A(n2357), .B(n2356), .Z(c[58]) );
  NANDN U2676 ( .A(n2234), .B(n2233), .Z(n2238) );
  NANDN U2677 ( .A(n2236), .B(n2235), .Z(n2237) );
  AND U2678 ( .A(n2238), .B(n2237), .Z(n2368) );
  NANDN U2679 ( .A(n2240), .B(n2239), .Z(n2244) );
  NANDN U2680 ( .A(n2242), .B(n2241), .Z(n2243) );
  AND U2681 ( .A(n2244), .B(n2243), .Z(n2366) );
  NANDN U2682 ( .A(n2246), .B(n2245), .Z(n2250) );
  NANDN U2683 ( .A(n2248), .B(n2247), .Z(n2249) );
  AND U2684 ( .A(n2250), .B(n2249), .Z(n2374) );
  NAND U2685 ( .A(n2252), .B(n2251), .Z(n2256) );
  NAND U2686 ( .A(n2254), .B(n2253), .Z(n2255) );
  AND U2687 ( .A(n2256), .B(n2255), .Z(n2371) );
  NANDN U2688 ( .A(n2258), .B(n2257), .Z(n2262) );
  NAND U2689 ( .A(n2260), .B(n2259), .Z(n2261) );
  AND U2690 ( .A(n2262), .B(n2261), .Z(n2484) );
  NAND U2691 ( .A(n572), .B(n2263), .Z(n2265) );
  XOR U2692 ( .A(b[13]), .B(a[15]), .Z(n2401) );
  NAND U2693 ( .A(n8585), .B(n2401), .Z(n2264) );
  NAND U2694 ( .A(n2265), .B(n2264), .Z(n2404) );
  NAND U2695 ( .A(b[0]), .B(a[27]), .Z(n2266) );
  XNOR U2696 ( .A(b[1]), .B(n2266), .Z(n2268) );
  NANDN U2697 ( .A(b[0]), .B(a[26]), .Z(n2267) );
  NAND U2698 ( .A(n2268), .B(n2267), .Z(n2405) );
  XNOR U2699 ( .A(n2404), .B(n2405), .Z(n2406) );
  NAND U2700 ( .A(n579), .B(n2269), .Z(n2271) );
  XOR U2701 ( .A(b[25]), .B(a[3]), .Z(n2464) );
  NAND U2702 ( .A(n9364), .B(n2464), .Z(n2270) );
  AND U2703 ( .A(n2271), .B(n2270), .Z(n2474) );
  XOR U2704 ( .A(b[27]), .B(b[26]), .Z(n2467) );
  XOR U2705 ( .A(b[27]), .B(a[0]), .Z(n2272) );
  NAND U2706 ( .A(n2467), .B(n2272), .Z(n2273) );
  NANDN U2707 ( .A(n2273), .B(n9692), .Z(n2275) );
  XOR U2708 ( .A(b[27]), .B(a[1]), .Z(n2468) );
  NANDN U2709 ( .A(n9692), .B(n2468), .Z(n2274) );
  NAND U2710 ( .A(n2275), .B(n2274), .Z(n2475) );
  XOR U2711 ( .A(n2474), .B(n2475), .Z(n2407) );
  XNOR U2712 ( .A(n2406), .B(n2407), .Z(n2437) );
  NAND U2713 ( .A(n569), .B(n2276), .Z(n2278) );
  XOR U2714 ( .A(b[7]), .B(a[21]), .Z(n2431) );
  NAND U2715 ( .A(n7819), .B(n2431), .Z(n2277) );
  AND U2716 ( .A(n2278), .B(n2277), .Z(n2458) );
  NAND U2717 ( .A(n567), .B(n2279), .Z(n2281) );
  XOR U2718 ( .A(b[5]), .B(a[23]), .Z(n2422) );
  NAND U2719 ( .A(n7235), .B(n2422), .Z(n2280) );
  AND U2720 ( .A(n2281), .B(n2280), .Z(n2456) );
  NAND U2721 ( .A(n9046), .B(n2282), .Z(n2284) );
  XOR U2722 ( .A(b[19]), .B(a[9]), .Z(n2416) );
  NAND U2723 ( .A(n575), .B(n2416), .Z(n2283) );
  NAND U2724 ( .A(n2284), .B(n2283), .Z(n2455) );
  XNOR U2725 ( .A(n2456), .B(n2455), .Z(n2457) );
  XOR U2726 ( .A(n2458), .B(n2457), .Z(n2438) );
  XNOR U2727 ( .A(n2437), .B(n2438), .Z(n2439) );
  NANDN U2728 ( .A(n2286), .B(n2285), .Z(n2290) );
  OR U2729 ( .A(n2288), .B(n2287), .Z(n2289) );
  NAND U2730 ( .A(n2290), .B(n2289), .Z(n2440) );
  XNOR U2731 ( .A(n2439), .B(n2440), .Z(n2386) );
  NANDN U2732 ( .A(n2292), .B(n2291), .Z(n2296) );
  OR U2733 ( .A(n2294), .B(n2293), .Z(n2295) );
  NAND U2734 ( .A(n2296), .B(n2295), .Z(n2384) );
  NANDN U2735 ( .A(n2298), .B(n2297), .Z(n2302) );
  NANDN U2736 ( .A(n2300), .B(n2299), .Z(n2301) );
  NAND U2737 ( .A(n2302), .B(n2301), .Z(n2383) );
  XOR U2738 ( .A(n2384), .B(n2383), .Z(n2385) );
  XOR U2739 ( .A(n2386), .B(n2385), .Z(n2392) );
  NANDN U2740 ( .A(n2303), .B(n2315), .Z(n2307) );
  NANDN U2741 ( .A(n2305), .B(n2304), .Z(n2306) );
  AND U2742 ( .A(n2307), .B(n2306), .Z(n2444) );
  OR U2743 ( .A(n2308), .B(n560), .Z(n2310) );
  XOR U2744 ( .A(b[3]), .B(a[25]), .Z(n2395) );
  NAND U2745 ( .A(n7245), .B(n2395), .Z(n2309) );
  AND U2746 ( .A(n2310), .B(n2309), .Z(n2477) );
  OR U2747 ( .A(n2311), .B(n557), .Z(n2313) );
  XOR U2748 ( .A(b[15]), .B(a[13]), .Z(n2471) );
  NAND U2749 ( .A(n8694), .B(n2471), .Z(n2312) );
  NAND U2750 ( .A(n2313), .B(n2312), .Z(n2476) );
  XNOR U2751 ( .A(n2477), .B(n2476), .Z(n2478) );
  NANDN U2752 ( .A(b[26]), .B(b[27]), .Z(n2314) );
  NAND U2753 ( .A(n9770), .B(b[27]), .Z(n9809) );
  NAND U2754 ( .A(n2314), .B(n9809), .Z(n9855) );
  ANDN U2755 ( .B(n9855), .A(n2315), .Z(n2479) );
  XOR U2756 ( .A(n2478), .B(n2479), .Z(n2443) );
  XNOR U2757 ( .A(n2444), .B(n2443), .Z(n2446) );
  NAND U2758 ( .A(n571), .B(n2316), .Z(n2318) );
  XOR U2759 ( .A(b[11]), .B(a[17]), .Z(n2425) );
  NAND U2760 ( .A(n8135), .B(n2425), .Z(n2317) );
  AND U2761 ( .A(n2318), .B(n2317), .Z(n2450) );
  NAND U2762 ( .A(n576), .B(n2319), .Z(n2321) );
  XOR U2763 ( .A(b[17]), .B(a[11]), .Z(n2428) );
  NAND U2764 ( .A(n9141), .B(n2428), .Z(n2320) );
  NAND U2765 ( .A(n2321), .B(n2320), .Z(n2449) );
  XNOR U2766 ( .A(n2450), .B(n2449), .Z(n2451) );
  NAND U2767 ( .A(n577), .B(n2322), .Z(n2324) );
  XOR U2768 ( .A(b[21]), .B(a[7]), .Z(n2419) );
  NAND U2769 ( .A(n9216), .B(n2419), .Z(n2323) );
  AND U2770 ( .A(n2324), .B(n2323), .Z(n2413) );
  NAND U2771 ( .A(n578), .B(n2325), .Z(n2327) );
  XOR U2772 ( .A(b[23]), .B(a[5]), .Z(n2398) );
  NAND U2773 ( .A(n9268), .B(n2398), .Z(n2326) );
  AND U2774 ( .A(n2327), .B(n2326), .Z(n2411) );
  NAND U2775 ( .A(n570), .B(n2328), .Z(n2330) );
  XOR U2776 ( .A(b[9]), .B(a[19]), .Z(n2434) );
  NAND U2777 ( .A(n8037), .B(n2434), .Z(n2329) );
  NAND U2778 ( .A(n2330), .B(n2329), .Z(n2410) );
  XNOR U2779 ( .A(n2411), .B(n2410), .Z(n2412) );
  XOR U2780 ( .A(n2413), .B(n2412), .Z(n2452) );
  XNOR U2781 ( .A(n2451), .B(n2452), .Z(n2445) );
  XOR U2782 ( .A(n2446), .B(n2445), .Z(n2390) );
  NANDN U2783 ( .A(n2332), .B(n2331), .Z(n2336) );
  NANDN U2784 ( .A(n2334), .B(n2333), .Z(n2335) );
  AND U2785 ( .A(n2336), .B(n2335), .Z(n2389) );
  XNOR U2786 ( .A(n2390), .B(n2389), .Z(n2391) );
  XNOR U2787 ( .A(n2392), .B(n2391), .Z(n2482) );
  NANDN U2788 ( .A(n2338), .B(n2337), .Z(n2342) );
  NAND U2789 ( .A(n2340), .B(n2339), .Z(n2341) );
  AND U2790 ( .A(n2342), .B(n2341), .Z(n2380) );
  NANDN U2791 ( .A(n2344), .B(n2343), .Z(n2348) );
  NANDN U2792 ( .A(n2346), .B(n2345), .Z(n2347) );
  AND U2793 ( .A(n2348), .B(n2347), .Z(n2377) );
  NANDN U2794 ( .A(n2350), .B(n2349), .Z(n2354) );
  OR U2795 ( .A(n2352), .B(n2351), .Z(n2353) );
  NAND U2796 ( .A(n2354), .B(n2353), .Z(n2378) );
  XNOR U2797 ( .A(n2377), .B(n2378), .Z(n2379) );
  XOR U2798 ( .A(n2380), .B(n2379), .Z(n2483) );
  XOR U2799 ( .A(n2482), .B(n2483), .Z(n2485) );
  XOR U2800 ( .A(n2484), .B(n2485), .Z(n2372) );
  XNOR U2801 ( .A(n2371), .B(n2372), .Z(n2373) );
  XNOR U2802 ( .A(n2374), .B(n2373), .Z(n2365) );
  XNOR U2803 ( .A(n2366), .B(n2365), .Z(n2367) );
  XNOR U2804 ( .A(n2368), .B(n2367), .Z(n2360) );
  XNOR U2805 ( .A(sreg[59]), .B(n2360), .Z(n2362) );
  NANDN U2806 ( .A(sreg[58]), .B(n2355), .Z(n2359) );
  NAND U2807 ( .A(n2357), .B(n2356), .Z(n2358) );
  NAND U2808 ( .A(n2359), .B(n2358), .Z(n2361) );
  XNOR U2809 ( .A(n2362), .B(n2361), .Z(c[59]) );
  NANDN U2810 ( .A(sreg[59]), .B(n2360), .Z(n2364) );
  NAND U2811 ( .A(n2362), .B(n2361), .Z(n2363) );
  NAND U2812 ( .A(n2364), .B(n2363), .Z(n2621) );
  XNOR U2813 ( .A(sreg[60]), .B(n2621), .Z(n2623) );
  NANDN U2814 ( .A(n2366), .B(n2365), .Z(n2370) );
  NANDN U2815 ( .A(n2368), .B(n2367), .Z(n2369) );
  AND U2816 ( .A(n2370), .B(n2369), .Z(n2491) );
  NANDN U2817 ( .A(n2372), .B(n2371), .Z(n2376) );
  NANDN U2818 ( .A(n2374), .B(n2373), .Z(n2375) );
  AND U2819 ( .A(n2376), .B(n2375), .Z(n2489) );
  NANDN U2820 ( .A(n2378), .B(n2377), .Z(n2382) );
  NANDN U2821 ( .A(n2380), .B(n2379), .Z(n2381) );
  AND U2822 ( .A(n2382), .B(n2381), .Z(n2497) );
  NAND U2823 ( .A(n2384), .B(n2383), .Z(n2388) );
  NAND U2824 ( .A(n2386), .B(n2385), .Z(n2387) );
  AND U2825 ( .A(n2388), .B(n2387), .Z(n2495) );
  NANDN U2826 ( .A(n2390), .B(n2389), .Z(n2394) );
  NANDN U2827 ( .A(n2392), .B(n2391), .Z(n2393) );
  AND U2828 ( .A(n2394), .B(n2393), .Z(n2494) );
  XNOR U2829 ( .A(n2495), .B(n2494), .Z(n2496) );
  XOR U2830 ( .A(n2497), .B(n2496), .Z(n2618) );
  NAND U2831 ( .A(n568), .B(n2395), .Z(n2397) );
  XOR U2832 ( .A(b[3]), .B(a[26]), .Z(n2558) );
  NAND U2833 ( .A(n7245), .B(n2558), .Z(n2396) );
  AND U2834 ( .A(n2397), .B(n2396), .Z(n2539) );
  NAND U2835 ( .A(n578), .B(n2398), .Z(n2400) );
  XOR U2836 ( .A(b[23]), .B(a[6]), .Z(n2564) );
  NAND U2837 ( .A(n9268), .B(n2564), .Z(n2399) );
  AND U2838 ( .A(n2400), .B(n2399), .Z(n2538) );
  NAND U2839 ( .A(n572), .B(n2401), .Z(n2403) );
  XOR U2840 ( .A(b[13]), .B(a[16]), .Z(n2528) );
  NAND U2841 ( .A(n8585), .B(n2528), .Z(n2402) );
  NAND U2842 ( .A(n2403), .B(n2402), .Z(n2537) );
  XOR U2843 ( .A(n2538), .B(n2537), .Z(n2540) );
  XOR U2844 ( .A(n2539), .B(n2540), .Z(n2592) );
  NANDN U2845 ( .A(n2405), .B(n2404), .Z(n2409) );
  NANDN U2846 ( .A(n2407), .B(n2406), .Z(n2408) );
  AND U2847 ( .A(n2409), .B(n2408), .Z(n2591) );
  XNOR U2848 ( .A(n2592), .B(n2591), .Z(n2593) );
  NANDN U2849 ( .A(n2411), .B(n2410), .Z(n2415) );
  NANDN U2850 ( .A(n2413), .B(n2412), .Z(n2414) );
  NAND U2851 ( .A(n2415), .B(n2414), .Z(n2594) );
  XNOR U2852 ( .A(n2593), .B(n2594), .Z(n2609) );
  NAND U2853 ( .A(n9046), .B(n2416), .Z(n2418) );
  XOR U2854 ( .A(b[19]), .B(a[10]), .Z(n2531) );
  NAND U2855 ( .A(n575), .B(n2531), .Z(n2417) );
  AND U2856 ( .A(n2418), .B(n2417), .Z(n2545) );
  NAND U2857 ( .A(n577), .B(n2419), .Z(n2421) );
  XOR U2858 ( .A(b[21]), .B(a[8]), .Z(n2552) );
  NAND U2859 ( .A(n9216), .B(n2552), .Z(n2420) );
  AND U2860 ( .A(n2421), .B(n2420), .Z(n2544) );
  NAND U2861 ( .A(n567), .B(n2422), .Z(n2424) );
  XOR U2862 ( .A(b[5]), .B(a[24]), .Z(n2555) );
  NAND U2863 ( .A(n7235), .B(n2555), .Z(n2423) );
  NAND U2864 ( .A(n2424), .B(n2423), .Z(n2543) );
  XOR U2865 ( .A(n2544), .B(n2543), .Z(n2546) );
  XOR U2866 ( .A(n2545), .B(n2546), .Z(n2606) );
  NAND U2867 ( .A(n571), .B(n2425), .Z(n2427) );
  XOR U2868 ( .A(b[11]), .B(a[18]), .Z(n2534) );
  NAND U2869 ( .A(n8135), .B(n2534), .Z(n2426) );
  AND U2870 ( .A(n2427), .B(n2426), .Z(n2581) );
  NAND U2871 ( .A(n576), .B(n2428), .Z(n2430) );
  XOR U2872 ( .A(b[17]), .B(a[12]), .Z(n2561) );
  NAND U2873 ( .A(n9141), .B(n2561), .Z(n2429) );
  AND U2874 ( .A(n2430), .B(n2429), .Z(n2580) );
  NAND U2875 ( .A(n569), .B(n2431), .Z(n2433) );
  XOR U2876 ( .A(b[7]), .B(a[22]), .Z(n2549) );
  NAND U2877 ( .A(n7819), .B(n2549), .Z(n2432) );
  NAND U2878 ( .A(n2433), .B(n2432), .Z(n2579) );
  XOR U2879 ( .A(n2580), .B(n2579), .Z(n2582) );
  XOR U2880 ( .A(n2581), .B(n2582), .Z(n2604) );
  NANDN U2881 ( .A(n564), .B(n2434), .Z(n2436) );
  XNOR U2882 ( .A(b[9]), .B(a[20]), .Z(n2570) );
  OR U2883 ( .A(n2570), .B(n8485), .Z(n2435) );
  AND U2884 ( .A(n2436), .B(n2435), .Z(n2603) );
  XNOR U2885 ( .A(n2604), .B(n2603), .Z(n2605) );
  XOR U2886 ( .A(n2606), .B(n2605), .Z(n2610) );
  XNOR U2887 ( .A(n2609), .B(n2610), .Z(n2612) );
  NANDN U2888 ( .A(n2438), .B(n2437), .Z(n2442) );
  NANDN U2889 ( .A(n2440), .B(n2439), .Z(n2441) );
  AND U2890 ( .A(n2442), .B(n2441), .Z(n2611) );
  XOR U2891 ( .A(n2612), .B(n2611), .Z(n2502) );
  NANDN U2892 ( .A(n2444), .B(n2443), .Z(n2448) );
  NAND U2893 ( .A(n2446), .B(n2445), .Z(n2447) );
  AND U2894 ( .A(n2448), .B(n2447), .Z(n2501) );
  NANDN U2895 ( .A(n2450), .B(n2449), .Z(n2454) );
  NANDN U2896 ( .A(n2452), .B(n2451), .Z(n2453) );
  AND U2897 ( .A(n2454), .B(n2453), .Z(n2588) );
  NANDN U2898 ( .A(n2456), .B(n2455), .Z(n2460) );
  NANDN U2899 ( .A(n2458), .B(n2457), .Z(n2459) );
  AND U2900 ( .A(n2460), .B(n2459), .Z(n2600) );
  NAND U2901 ( .A(b[0]), .B(a[28]), .Z(n2461) );
  XNOR U2902 ( .A(b[1]), .B(n2461), .Z(n2463) );
  NANDN U2903 ( .A(b[0]), .B(a[27]), .Z(n2462) );
  NAND U2904 ( .A(n2463), .B(n2462), .Z(n2576) );
  XNOR U2905 ( .A(b[27]), .B(b[28]), .Z(n9796) );
  AND U2906 ( .A(a[0]), .B(n581), .Z(n2573) );
  NAND U2907 ( .A(n579), .B(n2464), .Z(n2466) );
  XOR U2908 ( .A(b[25]), .B(a[4]), .Z(n2567) );
  NAND U2909 ( .A(n9364), .B(n2567), .Z(n2465) );
  AND U2910 ( .A(n2466), .B(n2465), .Z(n2574) );
  XOR U2911 ( .A(n2573), .B(n2574), .Z(n2575) );
  XOR U2912 ( .A(n2576), .B(n2575), .Z(n2598) );
  NAND U2913 ( .A(n582), .B(n2468), .Z(n2470) );
  XOR U2914 ( .A(b[27]), .B(a[2]), .Z(n2512) );
  NAND U2915 ( .A(n9770), .B(n2512), .Z(n2469) );
  AND U2916 ( .A(n2470), .B(n2469), .Z(n2507) );
  NAND U2917 ( .A(n573), .B(n2471), .Z(n2473) );
  XOR U2918 ( .A(b[15]), .B(a[14]), .Z(n2525) );
  NAND U2919 ( .A(n8694), .B(n2525), .Z(n2472) );
  NAND U2920 ( .A(n2473), .B(n2472), .Z(n2506) );
  XNOR U2921 ( .A(n2507), .B(n2506), .Z(n2509) );
  ANDN U2922 ( .B(n2475), .A(n2474), .Z(n2508) );
  XNOR U2923 ( .A(n2509), .B(n2508), .Z(n2597) );
  XNOR U2924 ( .A(n2598), .B(n2597), .Z(n2599) );
  XOR U2925 ( .A(n2600), .B(n2599), .Z(n2586) );
  NANDN U2926 ( .A(n2477), .B(n2476), .Z(n2481) );
  NAND U2927 ( .A(n2479), .B(n2478), .Z(n2480) );
  NAND U2928 ( .A(n2481), .B(n2480), .Z(n2585) );
  XNOR U2929 ( .A(n2586), .B(n2585), .Z(n2587) );
  XNOR U2930 ( .A(n2588), .B(n2587), .Z(n2500) );
  XOR U2931 ( .A(n2501), .B(n2500), .Z(n2503) );
  XOR U2932 ( .A(n2502), .B(n2503), .Z(n2616) );
  NANDN U2933 ( .A(n2483), .B(n2482), .Z(n2487) );
  NANDN U2934 ( .A(n2485), .B(n2484), .Z(n2486) );
  NAND U2935 ( .A(n2487), .B(n2486), .Z(n2615) );
  XNOR U2936 ( .A(n2616), .B(n2615), .Z(n2617) );
  XNOR U2937 ( .A(n2618), .B(n2617), .Z(n2488) );
  XNOR U2938 ( .A(n2489), .B(n2488), .Z(n2490) );
  XNOR U2939 ( .A(n2491), .B(n2490), .Z(n2622) );
  XNOR U2940 ( .A(n2623), .B(n2622), .Z(c[60]) );
  NANDN U2941 ( .A(n2489), .B(n2488), .Z(n2493) );
  NANDN U2942 ( .A(n2491), .B(n2490), .Z(n2492) );
  AND U2943 ( .A(n2493), .B(n2492), .Z(n2629) );
  NANDN U2944 ( .A(n2495), .B(n2494), .Z(n2499) );
  NAND U2945 ( .A(n2497), .B(n2496), .Z(n2498) );
  AND U2946 ( .A(n2499), .B(n2498), .Z(n2752) );
  NANDN U2947 ( .A(n2501), .B(n2500), .Z(n2505) );
  OR U2948 ( .A(n2503), .B(n2502), .Z(n2504) );
  AND U2949 ( .A(n2505), .B(n2504), .Z(n2751) );
  NANDN U2950 ( .A(n2507), .B(n2506), .Z(n2511) );
  NAND U2951 ( .A(n2509), .B(n2508), .Z(n2510) );
  AND U2952 ( .A(n2511), .B(n2510), .Z(n2741) );
  NAND U2953 ( .A(n582), .B(n2512), .Z(n2514) );
  XOR U2954 ( .A(b[27]), .B(a[3]), .Z(n2666) );
  NAND U2955 ( .A(n9770), .B(n2666), .Z(n2513) );
  AND U2956 ( .A(n2514), .B(n2513), .Z(n2709) );
  XOR U2957 ( .A(b[29]), .B(a[1]), .Z(n2703) );
  NAND U2958 ( .A(n581), .B(n2703), .Z(n2521) );
  ANDN U2959 ( .B(b[28]), .A(b[29]), .Z(n2515) );
  NAND U2960 ( .A(n2515), .B(a[0]), .Z(n2518) );
  NAND U2961 ( .A(b[27]), .B(b[28]), .Z(n2516) );
  NAND U2962 ( .A(b[29]), .B(n2516), .Z(n9909) );
  OR U2963 ( .A(a[0]), .B(n9909), .Z(n2517) );
  NAND U2964 ( .A(n2518), .B(n2517), .Z(n2519) );
  NANDN U2965 ( .A(n581), .B(n2519), .Z(n2520) );
  AND U2966 ( .A(n2521), .B(n2520), .Z(n2710) );
  XOR U2967 ( .A(n2709), .B(n2710), .Z(n2734) );
  NAND U2968 ( .A(b[0]), .B(a[29]), .Z(n2522) );
  XNOR U2969 ( .A(b[1]), .B(n2522), .Z(n2524) );
  NANDN U2970 ( .A(b[0]), .B(a[28]), .Z(n2523) );
  NAND U2971 ( .A(n2524), .B(n2523), .Z(n2732) );
  NANDN U2972 ( .A(n557), .B(n2525), .Z(n2527) );
  XNOR U2973 ( .A(b[15]), .B(a[15]), .Z(n2699) );
  OR U2974 ( .A(n2699), .B(n9067), .Z(n2526) );
  NAND U2975 ( .A(n2527), .B(n2526), .Z(n2733) );
  XOR U2976 ( .A(n2732), .B(n2733), .Z(n2735) );
  XOR U2977 ( .A(n2734), .B(n2735), .Z(n2739) );
  NAND U2978 ( .A(n572), .B(n2528), .Z(n2530) );
  XOR U2979 ( .A(b[13]), .B(a[17]), .Z(n2717) );
  NAND U2980 ( .A(n8585), .B(n2717), .Z(n2529) );
  AND U2981 ( .A(n2530), .B(n2529), .Z(n2729) );
  NAND U2982 ( .A(n9046), .B(n2531), .Z(n2533) );
  XOR U2983 ( .A(b[19]), .B(a[11]), .Z(n2720) );
  NAND U2984 ( .A(n575), .B(n2720), .Z(n2532) );
  AND U2985 ( .A(n2533), .B(n2532), .Z(n2727) );
  NAND U2986 ( .A(n571), .B(n2534), .Z(n2536) );
  XOR U2987 ( .A(b[11]), .B(a[19]), .Z(n2711) );
  NAND U2988 ( .A(n8135), .B(n2711), .Z(n2535) );
  NAND U2989 ( .A(n2536), .B(n2535), .Z(n2726) );
  XNOR U2990 ( .A(n2727), .B(n2726), .Z(n2728) );
  XNOR U2991 ( .A(n2729), .B(n2728), .Z(n2738) );
  XNOR U2992 ( .A(n2739), .B(n2738), .Z(n2740) );
  XNOR U2993 ( .A(n2741), .B(n2740), .Z(n2641) );
  NANDN U2994 ( .A(n2538), .B(n2537), .Z(n2542) );
  OR U2995 ( .A(n2540), .B(n2539), .Z(n2541) );
  AND U2996 ( .A(n2542), .B(n2541), .Z(n2639) );
  NANDN U2997 ( .A(n2544), .B(n2543), .Z(n2548) );
  OR U2998 ( .A(n2546), .B(n2545), .Z(n2547) );
  AND U2999 ( .A(n2548), .B(n2547), .Z(n2647) );
  NAND U3000 ( .A(n569), .B(n2549), .Z(n2551) );
  XOR U3001 ( .A(b[7]), .B(a[23]), .Z(n2723) );
  NAND U3002 ( .A(n7819), .B(n2723), .Z(n2550) );
  AND U3003 ( .A(n2551), .B(n2550), .Z(n2657) );
  NAND U3004 ( .A(n577), .B(n2552), .Z(n2554) );
  XOR U3005 ( .A(b[21]), .B(a[9]), .Z(n2678) );
  NAND U3006 ( .A(n9216), .B(n2678), .Z(n2553) );
  NAND U3007 ( .A(n2554), .B(n2553), .Z(n2656) );
  XNOR U3008 ( .A(n2657), .B(n2656), .Z(n2659) );
  OR U3009 ( .A(n9909), .B(n2573), .Z(n2658) );
  XNOR U3010 ( .A(n2659), .B(n2658), .Z(n2644) );
  NAND U3011 ( .A(n567), .B(n2555), .Z(n2557) );
  XOR U3012 ( .A(b[5]), .B(a[25]), .Z(n2693) );
  NAND U3013 ( .A(n7235), .B(n2693), .Z(n2556) );
  AND U3014 ( .A(n2557), .B(n2556), .Z(n2663) );
  NAND U3015 ( .A(n568), .B(n2558), .Z(n2560) );
  XOR U3016 ( .A(b[3]), .B(a[27]), .Z(n2696) );
  NAND U3017 ( .A(n7245), .B(n2696), .Z(n2559) );
  AND U3018 ( .A(n2560), .B(n2559), .Z(n2661) );
  NAND U3019 ( .A(n576), .B(n2561), .Z(n2563) );
  XOR U3020 ( .A(b[17]), .B(a[13]), .Z(n2706) );
  NAND U3021 ( .A(n9141), .B(n2706), .Z(n2562) );
  NAND U3022 ( .A(n2563), .B(n2562), .Z(n2660) );
  XNOR U3023 ( .A(n2661), .B(n2660), .Z(n2662) );
  XOR U3024 ( .A(n2663), .B(n2662), .Z(n2645) );
  XNOR U3025 ( .A(n2644), .B(n2645), .Z(n2646) );
  XNOR U3026 ( .A(n2647), .B(n2646), .Z(n2638) );
  XNOR U3027 ( .A(n2639), .B(n2638), .Z(n2640) );
  XOR U3028 ( .A(n2641), .B(n2640), .Z(n2745) );
  NAND U3029 ( .A(n578), .B(n2564), .Z(n2566) );
  XOR U3030 ( .A(b[23]), .B(a[7]), .Z(n2672) );
  NAND U3031 ( .A(n9268), .B(n2672), .Z(n2565) );
  AND U3032 ( .A(n2566), .B(n2565), .Z(n2652) );
  NAND U3033 ( .A(n579), .B(n2567), .Z(n2569) );
  XOR U3034 ( .A(b[25]), .B(a[5]), .Z(n2675) );
  NAND U3035 ( .A(n9364), .B(n2675), .Z(n2568) );
  AND U3036 ( .A(n2569), .B(n2568), .Z(n2651) );
  OR U3037 ( .A(n2570), .B(n564), .Z(n2572) );
  XOR U3038 ( .A(b[9]), .B(a[21]), .Z(n2714) );
  NAND U3039 ( .A(n8037), .B(n2714), .Z(n2571) );
  NAND U3040 ( .A(n2572), .B(n2571), .Z(n2650) );
  XOR U3041 ( .A(n2651), .B(n2650), .Z(n2653) );
  XOR U3042 ( .A(n2652), .B(n2653), .Z(n2688) );
  NANDN U3043 ( .A(n2574), .B(n2573), .Z(n2578) );
  OR U3044 ( .A(n2576), .B(n2575), .Z(n2577) );
  AND U3045 ( .A(n2578), .B(n2577), .Z(n2687) );
  XNOR U3046 ( .A(n2688), .B(n2687), .Z(n2689) );
  NANDN U3047 ( .A(n2580), .B(n2579), .Z(n2584) );
  OR U3048 ( .A(n2582), .B(n2581), .Z(n2583) );
  NAND U3049 ( .A(n2584), .B(n2583), .Z(n2690) );
  XNOR U3050 ( .A(n2689), .B(n2690), .Z(n2744) );
  XNOR U3051 ( .A(n2745), .B(n2744), .Z(n2747) );
  NANDN U3052 ( .A(n2586), .B(n2585), .Z(n2590) );
  NANDN U3053 ( .A(n2588), .B(n2587), .Z(n2589) );
  AND U3054 ( .A(n2590), .B(n2589), .Z(n2746) );
  XOR U3055 ( .A(n2747), .B(n2746), .Z(n2635) );
  NANDN U3056 ( .A(n2592), .B(n2591), .Z(n2596) );
  NANDN U3057 ( .A(n2594), .B(n2593), .Z(n2595) );
  AND U3058 ( .A(n2596), .B(n2595), .Z(n2683) );
  NANDN U3059 ( .A(n2598), .B(n2597), .Z(n2602) );
  NAND U3060 ( .A(n2600), .B(n2599), .Z(n2601) );
  AND U3061 ( .A(n2602), .B(n2601), .Z(n2682) );
  NANDN U3062 ( .A(n2604), .B(n2603), .Z(n2608) );
  NANDN U3063 ( .A(n2606), .B(n2605), .Z(n2607) );
  NAND U3064 ( .A(n2608), .B(n2607), .Z(n2681) );
  XOR U3065 ( .A(n2682), .B(n2681), .Z(n2684) );
  XOR U3066 ( .A(n2683), .B(n2684), .Z(n2633) );
  NANDN U3067 ( .A(n2610), .B(n2609), .Z(n2614) );
  NAND U3068 ( .A(n2612), .B(n2611), .Z(n2613) );
  AND U3069 ( .A(n2614), .B(n2613), .Z(n2632) );
  XNOR U3070 ( .A(n2633), .B(n2632), .Z(n2634) );
  XNOR U3071 ( .A(n2635), .B(n2634), .Z(n2750) );
  XOR U3072 ( .A(n2751), .B(n2750), .Z(n2753) );
  XOR U3073 ( .A(n2752), .B(n2753), .Z(n2627) );
  NANDN U3074 ( .A(n2616), .B(n2615), .Z(n2620) );
  NANDN U3075 ( .A(n2618), .B(n2617), .Z(n2619) );
  NAND U3076 ( .A(n2620), .B(n2619), .Z(n2626) );
  XNOR U3077 ( .A(n2627), .B(n2626), .Z(n2628) );
  XNOR U3078 ( .A(n2629), .B(n2628), .Z(n2756) );
  XNOR U3079 ( .A(sreg[61]), .B(n2756), .Z(n2758) );
  NANDN U3080 ( .A(sreg[60]), .B(n2621), .Z(n2625) );
  NAND U3081 ( .A(n2623), .B(n2622), .Z(n2624) );
  NAND U3082 ( .A(n2625), .B(n2624), .Z(n2757) );
  XNOR U3083 ( .A(n2758), .B(n2757), .Z(c[61]) );
  NANDN U3084 ( .A(n2627), .B(n2626), .Z(n2631) );
  NANDN U3085 ( .A(n2629), .B(n2628), .Z(n2630) );
  AND U3086 ( .A(n2631), .B(n2630), .Z(n2766) );
  NANDN U3087 ( .A(n2633), .B(n2632), .Z(n2637) );
  NANDN U3088 ( .A(n2635), .B(n2634), .Z(n2636) );
  AND U3089 ( .A(n2637), .B(n2636), .Z(n2896) );
  NANDN U3090 ( .A(n2639), .B(n2638), .Z(n2643) );
  NAND U3091 ( .A(n2641), .B(n2640), .Z(n2642) );
  AND U3092 ( .A(n2643), .B(n2642), .Z(n2890) );
  NANDN U3093 ( .A(n2645), .B(n2644), .Z(n2649) );
  NANDN U3094 ( .A(n2647), .B(n2646), .Z(n2648) );
  AND U3095 ( .A(n2649), .B(n2648), .Z(n2889) );
  NANDN U3096 ( .A(n2651), .B(n2650), .Z(n2655) );
  OR U3097 ( .A(n2653), .B(n2652), .Z(n2654) );
  AND U3098 ( .A(n2655), .B(n2654), .Z(n2777) );
  XNOR U3099 ( .A(n2777), .B(n2776), .Z(n2778) );
  NANDN U3100 ( .A(n2661), .B(n2660), .Z(n2665) );
  NANDN U3101 ( .A(n2663), .B(n2662), .Z(n2664) );
  AND U3102 ( .A(n2665), .B(n2664), .Z(n2875) );
  XNOR U3103 ( .A(b[30]), .B(b[29]), .Z(n9904) );
  AND U3104 ( .A(a[0]), .B(n584), .Z(n2849) );
  NAND U3105 ( .A(n582), .B(n2666), .Z(n2668) );
  XOR U3106 ( .A(b[27]), .B(a[4]), .Z(n2857) );
  NAND U3107 ( .A(n9770), .B(n2857), .Z(n2667) );
  AND U3108 ( .A(n2668), .B(n2667), .Z(n2807) );
  XNOR U3109 ( .A(n2849), .B(n2807), .Z(n2808) );
  NAND U3110 ( .A(b[0]), .B(a[30]), .Z(n2669) );
  XNOR U3111 ( .A(b[1]), .B(n2669), .Z(n2671) );
  NANDN U3112 ( .A(b[0]), .B(a[29]), .Z(n2670) );
  NAND U3113 ( .A(n2671), .B(n2670), .Z(n2809) );
  XNOR U3114 ( .A(n2808), .B(n2809), .Z(n2872) );
  NAND U3115 ( .A(n578), .B(n2672), .Z(n2674) );
  XOR U3116 ( .A(b[23]), .B(a[8]), .Z(n2851) );
  NAND U3117 ( .A(n9268), .B(n2851), .Z(n2673) );
  AND U3118 ( .A(n2674), .B(n2673), .Z(n2821) );
  NAND U3119 ( .A(n579), .B(n2675), .Z(n2677) );
  XOR U3120 ( .A(b[25]), .B(a[6]), .Z(n2854) );
  NAND U3121 ( .A(n9364), .B(n2854), .Z(n2676) );
  AND U3122 ( .A(n2677), .B(n2676), .Z(n2819) );
  NAND U3123 ( .A(n577), .B(n2678), .Z(n2680) );
  XOR U3124 ( .A(b[21]), .B(a[10]), .Z(n2863) );
  NAND U3125 ( .A(n9216), .B(n2863), .Z(n2679) );
  NAND U3126 ( .A(n2680), .B(n2679), .Z(n2818) );
  XNOR U3127 ( .A(n2819), .B(n2818), .Z(n2820) );
  XOR U3128 ( .A(n2821), .B(n2820), .Z(n2873) );
  XNOR U3129 ( .A(n2872), .B(n2873), .Z(n2874) );
  XOR U3130 ( .A(n2875), .B(n2874), .Z(n2779) );
  XNOR U3131 ( .A(n2778), .B(n2779), .Z(n2888) );
  XOR U3132 ( .A(n2889), .B(n2888), .Z(n2891) );
  XOR U3133 ( .A(n2890), .B(n2891), .Z(n2772) );
  NANDN U3134 ( .A(n2682), .B(n2681), .Z(n2686) );
  OR U3135 ( .A(n2684), .B(n2683), .Z(n2685) );
  AND U3136 ( .A(n2686), .B(n2685), .Z(n2771) );
  NANDN U3137 ( .A(n2688), .B(n2687), .Z(n2692) );
  NANDN U3138 ( .A(n2690), .B(n2689), .Z(n2691) );
  AND U3139 ( .A(n2692), .B(n2691), .Z(n2885) );
  NAND U3140 ( .A(n567), .B(n2693), .Z(n2695) );
  XOR U3141 ( .A(b[5]), .B(a[26]), .Z(n2837) );
  NAND U3142 ( .A(n7235), .B(n2837), .Z(n2694) );
  AND U3143 ( .A(n2695), .B(n2694), .Z(n2827) );
  NAND U3144 ( .A(n568), .B(n2696), .Z(n2698) );
  XOR U3145 ( .A(b[3]), .B(a[28]), .Z(n2843) );
  NAND U3146 ( .A(n7245), .B(n2843), .Z(n2697) );
  AND U3147 ( .A(n2698), .B(n2697), .Z(n2825) );
  OR U3148 ( .A(n2699), .B(n557), .Z(n2701) );
  XOR U3149 ( .A(b[15]), .B(a[16]), .Z(n2804) );
  NAND U3150 ( .A(n8694), .B(n2804), .Z(n2700) );
  NAND U3151 ( .A(n2701), .B(n2700), .Z(n2824) );
  XNOR U3152 ( .A(n2825), .B(n2824), .Z(n2826) );
  XNOR U3153 ( .A(n2827), .B(n2826), .Z(n2879) );
  XOR U3154 ( .A(b[28]), .B(b[29]), .Z(n2702) );
  NAND U3155 ( .A(n583), .B(n2703), .Z(n2705) );
  XOR U3156 ( .A(b[29]), .B(a[2]), .Z(n2794) );
  NAND U3157 ( .A(n581), .B(n2794), .Z(n2704) );
  AND U3158 ( .A(n2705), .B(n2704), .Z(n2831) );
  NAND U3159 ( .A(n576), .B(n2706), .Z(n2708) );
  XOR U3160 ( .A(b[17]), .B(a[14]), .Z(n2846) );
  NAND U3161 ( .A(n9141), .B(n2846), .Z(n2707) );
  NAND U3162 ( .A(n2708), .B(n2707), .Z(n2830) );
  XNOR U3163 ( .A(n2831), .B(n2830), .Z(n2833) );
  OR U3164 ( .A(n2710), .B(n2709), .Z(n2832) );
  XOR U3165 ( .A(n2833), .B(n2832), .Z(n2878) );
  XNOR U3166 ( .A(n2879), .B(n2878), .Z(n2880) );
  NAND U3167 ( .A(n571), .B(n2711), .Z(n2713) );
  XOR U3168 ( .A(b[11]), .B(a[20]), .Z(n2869) );
  NAND U3169 ( .A(n8135), .B(n2869), .Z(n2712) );
  AND U3170 ( .A(n2713), .B(n2712), .Z(n2813) );
  NAND U3171 ( .A(n570), .B(n2714), .Z(n2716) );
  XOR U3172 ( .A(b[9]), .B(a[22]), .Z(n2866) );
  NAND U3173 ( .A(n8037), .B(n2866), .Z(n2715) );
  NAND U3174 ( .A(n2716), .B(n2715), .Z(n2812) );
  XNOR U3175 ( .A(n2813), .B(n2812), .Z(n2814) );
  NAND U3176 ( .A(n572), .B(n2717), .Z(n2719) );
  XOR U3177 ( .A(b[13]), .B(a[18]), .Z(n2860) );
  NAND U3178 ( .A(n8585), .B(n2860), .Z(n2718) );
  AND U3179 ( .A(n2719), .B(n2718), .Z(n2791) );
  NAND U3180 ( .A(n9046), .B(n2720), .Z(n2722) );
  XOR U3181 ( .A(b[19]), .B(a[12]), .Z(n2840) );
  NAND U3182 ( .A(n575), .B(n2840), .Z(n2721) );
  AND U3183 ( .A(n2722), .B(n2721), .Z(n2789) );
  NAND U3184 ( .A(n569), .B(n2723), .Z(n2725) );
  XOR U3185 ( .A(b[7]), .B(a[24]), .Z(n2834) );
  NAND U3186 ( .A(n7819), .B(n2834), .Z(n2724) );
  NAND U3187 ( .A(n2725), .B(n2724), .Z(n2788) );
  XNOR U3188 ( .A(n2789), .B(n2788), .Z(n2790) );
  XOR U3189 ( .A(n2791), .B(n2790), .Z(n2815) );
  XOR U3190 ( .A(n2814), .B(n2815), .Z(n2881) );
  XNOR U3191 ( .A(n2880), .B(n2881), .Z(n2785) );
  NANDN U3192 ( .A(n2727), .B(n2726), .Z(n2731) );
  NANDN U3193 ( .A(n2729), .B(n2728), .Z(n2730) );
  AND U3194 ( .A(n2731), .B(n2730), .Z(n2783) );
  NANDN U3195 ( .A(n2733), .B(n2732), .Z(n2737) );
  OR U3196 ( .A(n2735), .B(n2734), .Z(n2736) );
  AND U3197 ( .A(n2737), .B(n2736), .Z(n2782) );
  XNOR U3198 ( .A(n2783), .B(n2782), .Z(n2784) );
  XOR U3199 ( .A(n2785), .B(n2784), .Z(n2883) );
  NANDN U3200 ( .A(n2739), .B(n2738), .Z(n2743) );
  NANDN U3201 ( .A(n2741), .B(n2740), .Z(n2742) );
  AND U3202 ( .A(n2743), .B(n2742), .Z(n2882) );
  XNOR U3203 ( .A(n2883), .B(n2882), .Z(n2884) );
  XNOR U3204 ( .A(n2885), .B(n2884), .Z(n2770) );
  XOR U3205 ( .A(n2771), .B(n2770), .Z(n2773) );
  XOR U3206 ( .A(n2772), .B(n2773), .Z(n2895) );
  NANDN U3207 ( .A(n2745), .B(n2744), .Z(n2749) );
  NAND U3208 ( .A(n2747), .B(n2746), .Z(n2748) );
  AND U3209 ( .A(n2749), .B(n2748), .Z(n2894) );
  XOR U3210 ( .A(n2895), .B(n2894), .Z(n2897) );
  XOR U3211 ( .A(n2896), .B(n2897), .Z(n2765) );
  NANDN U3212 ( .A(n2751), .B(n2750), .Z(n2755) );
  OR U3213 ( .A(n2753), .B(n2752), .Z(n2754) );
  AND U3214 ( .A(n2755), .B(n2754), .Z(n2764) );
  XOR U3215 ( .A(n2765), .B(n2764), .Z(n2767) );
  XNOR U3216 ( .A(n2766), .B(n2767), .Z(n2763) );
  NANDN U3217 ( .A(sreg[61]), .B(n2756), .Z(n2760) );
  NAND U3218 ( .A(n2758), .B(n2757), .Z(n2759) );
  AND U3219 ( .A(n2760), .B(n2759), .Z(n2762) );
  XNOR U3220 ( .A(sreg[62]), .B(n2762), .Z(n2761) );
  XNOR U3221 ( .A(n2763), .B(n2761), .Z(c[62]) );
  NANDN U3222 ( .A(n2765), .B(n2764), .Z(n2769) );
  OR U3223 ( .A(n2767), .B(n2766), .Z(n2768) );
  AND U3224 ( .A(n2769), .B(n2768), .Z(n2908) );
  NANDN U3225 ( .A(n2771), .B(n2770), .Z(n2775) );
  OR U3226 ( .A(n2773), .B(n2772), .Z(n2774) );
  AND U3227 ( .A(n2775), .B(n2774), .Z(n3042) );
  NANDN U3228 ( .A(n2777), .B(n2776), .Z(n2781) );
  NANDN U3229 ( .A(n2779), .B(n2778), .Z(n2780) );
  AND U3230 ( .A(n2781), .B(n2780), .Z(n2920) );
  NANDN U3231 ( .A(n2783), .B(n2782), .Z(n2787) );
  NAND U3232 ( .A(n2785), .B(n2784), .Z(n2786) );
  AND U3233 ( .A(n2787), .B(n2786), .Z(n2918) );
  NANDN U3234 ( .A(n2789), .B(n2788), .Z(n2793) );
  NANDN U3235 ( .A(n2791), .B(n2790), .Z(n2792) );
  AND U3236 ( .A(n2793), .B(n2792), .Z(n3024) );
  NAND U3237 ( .A(n583), .B(n2794), .Z(n2796) );
  XOR U3238 ( .A(b[29]), .B(a[3]), .Z(n3006) );
  NAND U3239 ( .A(n581), .B(n3006), .Z(n2795) );
  AND U3240 ( .A(n2796), .B(n2795), .Z(n2960) );
  XOR U3241 ( .A(b[30]), .B(b[31]), .Z(n2797) );
  AND U3242 ( .A(n2797), .B(n9904), .Z(n9764) );
  XOR U3243 ( .A(a[0]), .B(b[31]), .Z(n2798) );
  NAND U3244 ( .A(n9764), .B(n2798), .Z(n2800) );
  XOR U3245 ( .A(b[31]), .B(a[1]), .Z(n2970) );
  AND U3246 ( .A(n2970), .B(n584), .Z(n2799) );
  ANDN U3247 ( .B(n2800), .A(n2799), .Z(n2959) );
  XOR U3248 ( .A(n2960), .B(n2959), .Z(n2990) );
  NAND U3249 ( .A(b[0]), .B(a[31]), .Z(n2801) );
  XNOR U3250 ( .A(b[1]), .B(n2801), .Z(n2803) );
  NANDN U3251 ( .A(b[0]), .B(a[30]), .Z(n2802) );
  NAND U3252 ( .A(n2803), .B(n2802), .Z(n2988) );
  NANDN U3253 ( .A(n557), .B(n2804), .Z(n2806) );
  XNOR U3254 ( .A(b[15]), .B(a[17]), .Z(n2997) );
  OR U3255 ( .A(n2997), .B(n9067), .Z(n2805) );
  NAND U3256 ( .A(n2806), .B(n2805), .Z(n2989) );
  XOR U3257 ( .A(n2988), .B(n2989), .Z(n2991) );
  XOR U3258 ( .A(n2990), .B(n2991), .Z(n3022) );
  NANDN U3259 ( .A(n2807), .B(n2849), .Z(n2811) );
  NANDN U3260 ( .A(n2809), .B(n2808), .Z(n2810) );
  NAND U3261 ( .A(n2811), .B(n2810), .Z(n3021) );
  XNOR U3262 ( .A(n3022), .B(n3021), .Z(n3023) );
  XNOR U3263 ( .A(n3024), .B(n3023), .Z(n2917) );
  XNOR U3264 ( .A(n2918), .B(n2917), .Z(n2919) );
  XNOR U3265 ( .A(n2920), .B(n2919), .Z(n2914) );
  NANDN U3266 ( .A(n2813), .B(n2812), .Z(n2817) );
  NANDN U3267 ( .A(n2815), .B(n2814), .Z(n2816) );
  AND U3268 ( .A(n2817), .B(n2816), .Z(n2978) );
  NANDN U3269 ( .A(n2819), .B(n2818), .Z(n2823) );
  NANDN U3270 ( .A(n2821), .B(n2820), .Z(n2822) );
  AND U3271 ( .A(n2823), .B(n2822), .Z(n2977) );
  NANDN U3272 ( .A(n2825), .B(n2824), .Z(n2829) );
  NANDN U3273 ( .A(n2827), .B(n2826), .Z(n2828) );
  NAND U3274 ( .A(n2829), .B(n2828), .Z(n2976) );
  XOR U3275 ( .A(n2977), .B(n2976), .Z(n2979) );
  XOR U3276 ( .A(n2978), .B(n2979), .Z(n3035) );
  NAND U3277 ( .A(n569), .B(n2834), .Z(n2836) );
  XOR U3278 ( .A(b[7]), .B(a[25]), .Z(n2938) );
  NAND U3279 ( .A(n7819), .B(n2938), .Z(n2835) );
  AND U3280 ( .A(n2836), .B(n2835), .Z(n2956) );
  NAND U3281 ( .A(n567), .B(n2837), .Z(n2839) );
  XOR U3282 ( .A(b[5]), .B(a[27]), .Z(n2941) );
  NAND U3283 ( .A(n7235), .B(n2941), .Z(n2838) );
  AND U3284 ( .A(n2839), .B(n2838), .Z(n2954) );
  NAND U3285 ( .A(n9046), .B(n2840), .Z(n2842) );
  XOR U3286 ( .A(b[19]), .B(a[13]), .Z(n2944) );
  NAND U3287 ( .A(n575), .B(n2944), .Z(n2841) );
  NAND U3288 ( .A(n2842), .B(n2841), .Z(n2953) );
  XNOR U3289 ( .A(n2954), .B(n2953), .Z(n2955) );
  XNOR U3290 ( .A(n2956), .B(n2955), .Z(n3015) );
  NAND U3291 ( .A(n568), .B(n2843), .Z(n2845) );
  XOR U3292 ( .A(b[3]), .B(a[29]), .Z(n2961) );
  NAND U3293 ( .A(n7245), .B(n2961), .Z(n2844) );
  AND U3294 ( .A(n2845), .B(n2844), .Z(n2985) );
  NAND U3295 ( .A(n576), .B(n2846), .Z(n2848) );
  XOR U3296 ( .A(b[17]), .B(a[15]), .Z(n2964) );
  NAND U3297 ( .A(n9141), .B(n2964), .Z(n2847) );
  AND U3298 ( .A(n2848), .B(n2847), .Z(n2983) );
  NAND U3299 ( .A(b[30]), .B(b[29]), .Z(n9926) );
  ANDN U3300 ( .B(n9926), .A(n2849), .Z(n2850) );
  AND U3301 ( .A(b[31]), .B(n2850), .Z(n2982) );
  XNOR U3302 ( .A(n2983), .B(n2982), .Z(n2984) );
  XOR U3303 ( .A(n2985), .B(n2984), .Z(n3016) );
  XOR U3304 ( .A(n3015), .B(n3016), .Z(n3018) );
  XOR U3305 ( .A(n3017), .B(n3018), .Z(n3034) );
  NAND U3306 ( .A(n578), .B(n2851), .Z(n2853) );
  XOR U3307 ( .A(b[23]), .B(a[9]), .Z(n2973) );
  NAND U3308 ( .A(n9268), .B(n2973), .Z(n2852) );
  AND U3309 ( .A(n2853), .B(n2852), .Z(n2949) );
  NAND U3310 ( .A(n579), .B(n2854), .Z(n2856) );
  XOR U3311 ( .A(b[25]), .B(a[7]), .Z(n2929) );
  NAND U3312 ( .A(n9364), .B(n2929), .Z(n2855) );
  AND U3313 ( .A(n2856), .B(n2855), .Z(n2948) );
  NAND U3314 ( .A(n582), .B(n2857), .Z(n2859) );
  XOR U3315 ( .A(b[27]), .B(a[5]), .Z(n2932) );
  NAND U3316 ( .A(n9770), .B(n2932), .Z(n2858) );
  NAND U3317 ( .A(n2859), .B(n2858), .Z(n2947) );
  XOR U3318 ( .A(n2948), .B(n2947), .Z(n2950) );
  XOR U3319 ( .A(n2949), .B(n2950), .Z(n2926) );
  NAND U3320 ( .A(n572), .B(n2860), .Z(n2862) );
  XOR U3321 ( .A(b[13]), .B(a[19]), .Z(n3000) );
  NAND U3322 ( .A(n8585), .B(n3000), .Z(n2861) );
  AND U3323 ( .A(n2862), .B(n2861), .Z(n3011) );
  NAND U3324 ( .A(n577), .B(n2863), .Z(n2865) );
  XOR U3325 ( .A(b[21]), .B(a[11]), .Z(n2994) );
  NAND U3326 ( .A(n9216), .B(n2994), .Z(n2864) );
  AND U3327 ( .A(n2865), .B(n2864), .Z(n3010) );
  NAND U3328 ( .A(n570), .B(n2866), .Z(n2868) );
  XOR U3329 ( .A(b[9]), .B(a[23]), .Z(n2967) );
  NAND U3330 ( .A(n8037), .B(n2967), .Z(n2867) );
  NAND U3331 ( .A(n2868), .B(n2867), .Z(n3009) );
  XOR U3332 ( .A(n3010), .B(n3009), .Z(n3012) );
  XOR U3333 ( .A(n3011), .B(n3012), .Z(n2924) );
  NANDN U3334 ( .A(n562), .B(n2869), .Z(n2871) );
  XNOR U3335 ( .A(b[11]), .B(a[21]), .Z(n2935) );
  OR U3336 ( .A(n2935), .B(n8701), .Z(n2870) );
  AND U3337 ( .A(n2871), .B(n2870), .Z(n2923) );
  XNOR U3338 ( .A(n2924), .B(n2923), .Z(n2925) );
  XNOR U3339 ( .A(n2926), .B(n2925), .Z(n3033) );
  XOR U3340 ( .A(n3034), .B(n3033), .Z(n3036) );
  XOR U3341 ( .A(n3035), .B(n3036), .Z(n3030) );
  NANDN U3342 ( .A(n2873), .B(n2872), .Z(n2877) );
  NANDN U3343 ( .A(n2875), .B(n2874), .Z(n2876) );
  AND U3344 ( .A(n2877), .B(n2876), .Z(n3028) );
  XNOR U3345 ( .A(n3028), .B(n3027), .Z(n3029) );
  XNOR U3346 ( .A(n3030), .B(n3029), .Z(n2911) );
  NANDN U3347 ( .A(n2883), .B(n2882), .Z(n2887) );
  NANDN U3348 ( .A(n2885), .B(n2884), .Z(n2886) );
  NAND U3349 ( .A(n2887), .B(n2886), .Z(n2912) );
  XNOR U3350 ( .A(n2911), .B(n2912), .Z(n2913) );
  XOR U3351 ( .A(n2914), .B(n2913), .Z(n3040) );
  NANDN U3352 ( .A(n2889), .B(n2888), .Z(n2893) );
  OR U3353 ( .A(n2891), .B(n2890), .Z(n2892) );
  AND U3354 ( .A(n2893), .B(n2892), .Z(n3039) );
  XNOR U3355 ( .A(n3040), .B(n3039), .Z(n3041) );
  XNOR U3356 ( .A(n3042), .B(n3041), .Z(n2905) );
  NANDN U3357 ( .A(n2895), .B(n2894), .Z(n2899) );
  OR U3358 ( .A(n2897), .B(n2896), .Z(n2898) );
  NAND U3359 ( .A(n2899), .B(n2898), .Z(n2906) );
  XNOR U3360 ( .A(n2905), .B(n2906), .Z(n2907) );
  XNOR U3361 ( .A(n2908), .B(n2907), .Z(n2900) );
  XNOR U3362 ( .A(sreg[63]), .B(n2900), .Z(n2901) );
  XOR U3363 ( .A(n2902), .B(n2901), .Z(c[63]) );
  NANDN U3364 ( .A(sreg[63]), .B(n2900), .Z(n2904) );
  NANDN U3365 ( .A(n2902), .B(n2901), .Z(n2903) );
  NAND U3366 ( .A(n2904), .B(n2903), .Z(n3046) );
  NANDN U3367 ( .A(n2906), .B(n2905), .Z(n2910) );
  NANDN U3368 ( .A(n2908), .B(n2907), .Z(n2909) );
  AND U3369 ( .A(n2910), .B(n2909), .Z(n3051) );
  NANDN U3370 ( .A(n2912), .B(n2911), .Z(n2916) );
  NAND U3371 ( .A(n2914), .B(n2913), .Z(n2915) );
  AND U3372 ( .A(n2916), .B(n2915), .Z(n3188) );
  NANDN U3373 ( .A(n2918), .B(n2917), .Z(n2922) );
  NANDN U3374 ( .A(n2920), .B(n2919), .Z(n2921) );
  AND U3375 ( .A(n2922), .B(n2921), .Z(n3187) );
  NANDN U3376 ( .A(n2924), .B(n2923), .Z(n2928) );
  NANDN U3377 ( .A(n2926), .B(n2925), .Z(n2927) );
  AND U3378 ( .A(n2928), .B(n2927), .Z(n3087) );
  NAND U3379 ( .A(n579), .B(n2929), .Z(n2931) );
  XOR U3380 ( .A(b[25]), .B(a[8]), .Z(n3111) );
  NAND U3381 ( .A(n9364), .B(n3111), .Z(n2930) );
  AND U3382 ( .A(n2931), .B(n2930), .Z(n3131) );
  NAND U3383 ( .A(n582), .B(n2932), .Z(n2934) );
  XOR U3384 ( .A(b[27]), .B(a[6]), .Z(n3120) );
  NAND U3385 ( .A(n9770), .B(n3120), .Z(n2933) );
  AND U3386 ( .A(n2934), .B(n2933), .Z(n3130) );
  OR U3387 ( .A(n2935), .B(n562), .Z(n2937) );
  XOR U3388 ( .A(b[11]), .B(a[22]), .Z(n3105) );
  NAND U3389 ( .A(n8135), .B(n3105), .Z(n2936) );
  NAND U3390 ( .A(n2937), .B(n2936), .Z(n3129) );
  XOR U3391 ( .A(n3130), .B(n3129), .Z(n3132) );
  XOR U3392 ( .A(n3131), .B(n3132), .Z(n3067) );
  NAND U3393 ( .A(n569), .B(n2938), .Z(n2940) );
  XOR U3394 ( .A(b[7]), .B(a[26]), .Z(n3096) );
  NAND U3395 ( .A(n7819), .B(n3096), .Z(n2939) );
  AND U3396 ( .A(n2940), .B(n2939), .Z(n3158) );
  NAND U3397 ( .A(n567), .B(n2941), .Z(n2943) );
  XOR U3398 ( .A(b[5]), .B(a[28]), .Z(n3099) );
  NAND U3399 ( .A(n7235), .B(n3099), .Z(n2942) );
  AND U3400 ( .A(n2943), .B(n2942), .Z(n3157) );
  NAND U3401 ( .A(n9046), .B(n2944), .Z(n2946) );
  XOR U3402 ( .A(b[19]), .B(a[14]), .Z(n3147) );
  NAND U3403 ( .A(n575), .B(n3147), .Z(n2945) );
  NAND U3404 ( .A(n2946), .B(n2945), .Z(n3156) );
  XOR U3405 ( .A(n3157), .B(n3156), .Z(n3159) );
  XNOR U3406 ( .A(n3158), .B(n3159), .Z(n3066) );
  XNOR U3407 ( .A(n3067), .B(n3066), .Z(n3069) );
  NANDN U3408 ( .A(n2948), .B(n2947), .Z(n2952) );
  OR U3409 ( .A(n2950), .B(n2949), .Z(n2951) );
  AND U3410 ( .A(n2952), .B(n2951), .Z(n3068) );
  XOR U3411 ( .A(n3069), .B(n3068), .Z(n3085) );
  NANDN U3412 ( .A(n2954), .B(n2953), .Z(n2958) );
  NANDN U3413 ( .A(n2956), .B(n2955), .Z(n2957) );
  AND U3414 ( .A(n2958), .B(n2957), .Z(n3075) );
  NOR U3415 ( .A(n2960), .B(n2959), .Z(n3093) );
  NANDN U3416 ( .A(n560), .B(n2961), .Z(n2963) );
  XNOR U3417 ( .A(b[3]), .B(a[30]), .Z(n3108) );
  OR U3418 ( .A(n3108), .B(n7784), .Z(n2962) );
  AND U3419 ( .A(n2963), .B(n2962), .Z(n3091) );
  NANDN U3420 ( .A(n554), .B(n2964), .Z(n2966) );
  XNOR U3421 ( .A(b[17]), .B(a[16]), .Z(n3126) );
  OR U3422 ( .A(n3126), .B(n9195), .Z(n2965) );
  AND U3423 ( .A(n2966), .B(n2965), .Z(n3090) );
  XOR U3424 ( .A(n3091), .B(n3090), .Z(n3092) );
  XOR U3425 ( .A(n3093), .B(n3092), .Z(n3073) );
  NAND U3426 ( .A(n570), .B(n2967), .Z(n2969) );
  XOR U3427 ( .A(b[9]), .B(a[24]), .Z(n3102) );
  NAND U3428 ( .A(n8037), .B(n3102), .Z(n2968) );
  AND U3429 ( .A(n2969), .B(n2968), .Z(n3171) );
  NAND U3430 ( .A(n9764), .B(n2970), .Z(n2972) );
  XOR U3431 ( .A(b[31]), .B(a[2]), .Z(n3123) );
  NAND U3432 ( .A(n584), .B(n3123), .Z(n2971) );
  AND U3433 ( .A(n2972), .B(n2971), .Z(n3169) );
  NAND U3434 ( .A(n578), .B(n2973), .Z(n2975) );
  XOR U3435 ( .A(b[23]), .B(a[10]), .Z(n3144) );
  NAND U3436 ( .A(n9268), .B(n3144), .Z(n2974) );
  NAND U3437 ( .A(n2975), .B(n2974), .Z(n3168) );
  XNOR U3438 ( .A(n3169), .B(n3168), .Z(n3170) );
  XNOR U3439 ( .A(n3171), .B(n3170), .Z(n3072) );
  XOR U3440 ( .A(n3073), .B(n3072), .Z(n3074) );
  XNOR U3441 ( .A(n3075), .B(n3074), .Z(n3084) );
  XNOR U3442 ( .A(n3085), .B(n3084), .Z(n3086) );
  XOR U3443 ( .A(n3087), .B(n3086), .Z(n3055) );
  NANDN U3444 ( .A(n2977), .B(n2976), .Z(n2981) );
  OR U3445 ( .A(n2979), .B(n2978), .Z(n2980) );
  AND U3446 ( .A(n2981), .B(n2980), .Z(n3054) );
  XNOR U3447 ( .A(n3055), .B(n3054), .Z(n3057) );
  NANDN U3448 ( .A(n2983), .B(n2982), .Z(n2987) );
  NANDN U3449 ( .A(n2985), .B(n2984), .Z(n2986) );
  AND U3450 ( .A(n2987), .B(n2986), .Z(n3079) );
  NANDN U3451 ( .A(n2989), .B(n2988), .Z(n2993) );
  OR U3452 ( .A(n2991), .B(n2990), .Z(n2992) );
  AND U3453 ( .A(n2993), .B(n2992), .Z(n3078) );
  XNOR U3454 ( .A(n3079), .B(n3078), .Z(n3081) );
  NAND U3455 ( .A(n577), .B(n2994), .Z(n2996) );
  XOR U3456 ( .A(b[21]), .B(a[12]), .Z(n3141) );
  NAND U3457 ( .A(n9216), .B(n3141), .Z(n2995) );
  AND U3458 ( .A(n2996), .B(n2995), .Z(n3138) );
  OR U3459 ( .A(n2997), .B(n557), .Z(n2999) );
  XOR U3460 ( .A(b[15]), .B(a[18]), .Z(n3150) );
  NAND U3461 ( .A(n8694), .B(n3150), .Z(n2998) );
  AND U3462 ( .A(n2999), .B(n2998), .Z(n3136) );
  NAND U3463 ( .A(n572), .B(n3000), .Z(n3002) );
  XOR U3464 ( .A(b[13]), .B(a[20]), .Z(n3117) );
  NAND U3465 ( .A(n8585), .B(n3117), .Z(n3001) );
  NAND U3466 ( .A(n3002), .B(n3001), .Z(n3135) );
  XNOR U3467 ( .A(n3136), .B(n3135), .Z(n3137) );
  XNOR U3468 ( .A(n3138), .B(n3137), .Z(n3175) );
  NAND U3469 ( .A(b[0]), .B(a[32]), .Z(n3003) );
  XNOR U3470 ( .A(b[1]), .B(n3003), .Z(n3005) );
  NANDN U3471 ( .A(b[0]), .B(a[31]), .Z(n3004) );
  NAND U3472 ( .A(n3005), .B(n3004), .Z(n3165) );
  NAND U3473 ( .A(n583), .B(n3006), .Z(n3008) );
  XOR U3474 ( .A(b[29]), .B(a[4]), .Z(n3153) );
  NAND U3475 ( .A(n581), .B(n3153), .Z(n3007) );
  AND U3476 ( .A(n3008), .B(n3007), .Z(n3163) );
  AND U3477 ( .A(b[31]), .B(a[0]), .Z(n3162) );
  XOR U3478 ( .A(n3163), .B(n3162), .Z(n3164) );
  XOR U3479 ( .A(n3165), .B(n3164), .Z(n3174) );
  XOR U3480 ( .A(n3175), .B(n3174), .Z(n3177) );
  NANDN U3481 ( .A(n3010), .B(n3009), .Z(n3014) );
  OR U3482 ( .A(n3012), .B(n3011), .Z(n3013) );
  NAND U3483 ( .A(n3014), .B(n3013), .Z(n3176) );
  XOR U3484 ( .A(n3177), .B(n3176), .Z(n3080) );
  XOR U3485 ( .A(n3081), .B(n3080), .Z(n3061) );
  NANDN U3486 ( .A(n3016), .B(n3015), .Z(n3020) );
  OR U3487 ( .A(n3018), .B(n3017), .Z(n3019) );
  AND U3488 ( .A(n3020), .B(n3019), .Z(n3060) );
  XNOR U3489 ( .A(n3061), .B(n3060), .Z(n3062) );
  NANDN U3490 ( .A(n3022), .B(n3021), .Z(n3026) );
  NANDN U3491 ( .A(n3024), .B(n3023), .Z(n3025) );
  NAND U3492 ( .A(n3026), .B(n3025), .Z(n3063) );
  XNOR U3493 ( .A(n3062), .B(n3063), .Z(n3056) );
  XOR U3494 ( .A(n3057), .B(n3056), .Z(n3183) );
  NANDN U3495 ( .A(n3028), .B(n3027), .Z(n3032) );
  NANDN U3496 ( .A(n3030), .B(n3029), .Z(n3031) );
  AND U3497 ( .A(n3032), .B(n3031), .Z(n3181) );
  NANDN U3498 ( .A(n3034), .B(n3033), .Z(n3038) );
  OR U3499 ( .A(n3036), .B(n3035), .Z(n3037) );
  AND U3500 ( .A(n3038), .B(n3037), .Z(n3180) );
  XNOR U3501 ( .A(n3181), .B(n3180), .Z(n3182) );
  XNOR U3502 ( .A(n3183), .B(n3182), .Z(n3186) );
  XOR U3503 ( .A(n3187), .B(n3186), .Z(n3189) );
  XOR U3504 ( .A(n3188), .B(n3189), .Z(n3049) );
  NANDN U3505 ( .A(n3040), .B(n3039), .Z(n3044) );
  NANDN U3506 ( .A(n3042), .B(n3041), .Z(n3043) );
  NAND U3507 ( .A(n3044), .B(n3043), .Z(n3048) );
  XNOR U3508 ( .A(n3049), .B(n3048), .Z(n3050) );
  XNOR U3509 ( .A(n3051), .B(n3050), .Z(n3047) );
  XNOR U3510 ( .A(sreg[64]), .B(n3047), .Z(n3045) );
  XNOR U3511 ( .A(n3046), .B(n3045), .Z(c[64]) );
  NANDN U3512 ( .A(n3049), .B(n3048), .Z(n3053) );
  NANDN U3513 ( .A(n3051), .B(n3050), .Z(n3052) );
  AND U3514 ( .A(n3053), .B(n3052), .Z(n3195) );
  NANDN U3515 ( .A(n3055), .B(n3054), .Z(n3059) );
  NAND U3516 ( .A(n3057), .B(n3056), .Z(n3058) );
  AND U3517 ( .A(n3059), .B(n3058), .Z(n3207) );
  NANDN U3518 ( .A(n3061), .B(n3060), .Z(n3065) );
  NANDN U3519 ( .A(n3063), .B(n3062), .Z(n3064) );
  AND U3520 ( .A(n3065), .B(n3064), .Z(n3205) );
  NANDN U3521 ( .A(n3067), .B(n3066), .Z(n3071) );
  NAND U3522 ( .A(n3069), .B(n3068), .Z(n3070) );
  AND U3523 ( .A(n3071), .B(n3070), .Z(n3217) );
  NAND U3524 ( .A(n3073), .B(n3072), .Z(n3077) );
  NANDN U3525 ( .A(n3075), .B(n3074), .Z(n3076) );
  AND U3526 ( .A(n3077), .B(n3076), .Z(n3216) );
  XNOR U3527 ( .A(n3217), .B(n3216), .Z(n3218) );
  NANDN U3528 ( .A(n3079), .B(n3078), .Z(n3083) );
  NAND U3529 ( .A(n3081), .B(n3080), .Z(n3082) );
  NAND U3530 ( .A(n3083), .B(n3082), .Z(n3219) );
  XNOR U3531 ( .A(n3218), .B(n3219), .Z(n3204) );
  XNOR U3532 ( .A(n3205), .B(n3204), .Z(n3206) );
  XNOR U3533 ( .A(n3207), .B(n3206), .Z(n3198) );
  NANDN U3534 ( .A(n3085), .B(n3084), .Z(n3089) );
  NAND U3535 ( .A(n3087), .B(n3086), .Z(n3088) );
  AND U3536 ( .A(n3089), .B(n3088), .Z(n3332) );
  NAND U3537 ( .A(n3091), .B(n3090), .Z(n3095) );
  NANDN U3538 ( .A(n3093), .B(n3092), .Z(n3094) );
  AND U3539 ( .A(n3095), .B(n3094), .Z(n3210) );
  NAND U3540 ( .A(n569), .B(n3096), .Z(n3098) );
  XOR U3541 ( .A(b[7]), .B(a[27]), .Z(n3309) );
  NAND U3542 ( .A(n7819), .B(n3309), .Z(n3097) );
  AND U3543 ( .A(n3098), .B(n3097), .Z(n3241) );
  NAND U3544 ( .A(n567), .B(n3099), .Z(n3101) );
  XOR U3545 ( .A(b[5]), .B(a[29]), .Z(n3258) );
  NAND U3546 ( .A(n7235), .B(n3258), .Z(n3100) );
  NAND U3547 ( .A(n3101), .B(n3100), .Z(n3240) );
  XNOR U3548 ( .A(n3241), .B(n3240), .Z(n3243) );
  NAND U3549 ( .A(n570), .B(n3102), .Z(n3104) );
  XOR U3550 ( .A(b[9]), .B(a[25]), .Z(n3327) );
  NAND U3551 ( .A(n8037), .B(n3327), .Z(n3103) );
  AND U3552 ( .A(n3104), .B(n3103), .Z(n3237) );
  NAND U3553 ( .A(n571), .B(n3105), .Z(n3107) );
  XOR U3554 ( .A(b[11]), .B(a[23]), .Z(n3318) );
  NAND U3555 ( .A(n8135), .B(n3318), .Z(n3106) );
  AND U3556 ( .A(n3107), .B(n3106), .Z(n3235) );
  OR U3557 ( .A(n3108), .B(n560), .Z(n3110) );
  XOR U3558 ( .A(b[3]), .B(a[31]), .Z(n3249) );
  NAND U3559 ( .A(n7245), .B(n3249), .Z(n3109) );
  NAND U3560 ( .A(n3110), .B(n3109), .Z(n3234) );
  XNOR U3561 ( .A(n3235), .B(n3234), .Z(n3236) );
  XNOR U3562 ( .A(n3237), .B(n3236), .Z(n3242) );
  XOR U3563 ( .A(n3243), .B(n3242), .Z(n3284) );
  NAND U3564 ( .A(n579), .B(n3111), .Z(n3113) );
  XOR U3565 ( .A(b[25]), .B(a[9]), .Z(n3312) );
  NAND U3566 ( .A(n9364), .B(n3312), .Z(n3112) );
  AND U3567 ( .A(n3113), .B(n3112), .Z(n3290) );
  NAND U3568 ( .A(b[0]), .B(a[33]), .Z(n3114) );
  XNOR U3569 ( .A(b[1]), .B(n3114), .Z(n3116) );
  NANDN U3570 ( .A(b[0]), .B(a[32]), .Z(n3115) );
  NAND U3571 ( .A(n3116), .B(n3115), .Z(n3289) );
  NAND U3572 ( .A(n572), .B(n3117), .Z(n3119) );
  XOR U3573 ( .A(b[13]), .B(a[21]), .Z(n3315) );
  NAND U3574 ( .A(n8585), .B(n3315), .Z(n3118) );
  NAND U3575 ( .A(n3119), .B(n3118), .Z(n3288) );
  XOR U3576 ( .A(n3289), .B(n3288), .Z(n3291) );
  XOR U3577 ( .A(n3290), .B(n3291), .Z(n3283) );
  NAND U3578 ( .A(n582), .B(n3120), .Z(n3122) );
  XOR U3579 ( .A(b[27]), .B(a[7]), .Z(n3255) );
  NAND U3580 ( .A(n9770), .B(n3255), .Z(n3121) );
  AND U3581 ( .A(n3122), .B(n3121), .Z(n3230) );
  NAND U3582 ( .A(n9764), .B(n3123), .Z(n3125) );
  XOR U3583 ( .A(b[31]), .B(a[3]), .Z(n3246) );
  NAND U3584 ( .A(n584), .B(n3246), .Z(n3124) );
  AND U3585 ( .A(n3125), .B(n3124), .Z(n3229) );
  OR U3586 ( .A(n3126), .B(n554), .Z(n3128) );
  XOR U3587 ( .A(b[17]), .B(a[17]), .Z(n3252) );
  NAND U3588 ( .A(n9141), .B(n3252), .Z(n3127) );
  NAND U3589 ( .A(n3128), .B(n3127), .Z(n3228) );
  XOR U3590 ( .A(n3229), .B(n3228), .Z(n3231) );
  XNOR U3591 ( .A(n3230), .B(n3231), .Z(n3282) );
  XOR U3592 ( .A(n3283), .B(n3282), .Z(n3285) );
  XOR U3593 ( .A(n3284), .B(n3285), .Z(n3273) );
  NANDN U3594 ( .A(n3130), .B(n3129), .Z(n3134) );
  OR U3595 ( .A(n3132), .B(n3131), .Z(n3133) );
  AND U3596 ( .A(n3134), .B(n3133), .Z(n3271) );
  NANDN U3597 ( .A(n3136), .B(n3135), .Z(n3140) );
  NANDN U3598 ( .A(n3138), .B(n3137), .Z(n3139) );
  NAND U3599 ( .A(n3140), .B(n3139), .Z(n3270) );
  XNOR U3600 ( .A(n3271), .B(n3270), .Z(n3272) );
  XOR U3601 ( .A(n3273), .B(n3272), .Z(n3211) );
  XNOR U3602 ( .A(n3210), .B(n3211), .Z(n3213) );
  NAND U3603 ( .A(n577), .B(n3141), .Z(n3143) );
  XOR U3604 ( .A(b[21]), .B(a[13]), .Z(n3324) );
  NAND U3605 ( .A(n9216), .B(n3324), .Z(n3142) );
  AND U3606 ( .A(n3143), .B(n3142), .Z(n3296) );
  NAND U3607 ( .A(n578), .B(n3144), .Z(n3146) );
  XOR U3608 ( .A(b[23]), .B(a[11]), .Z(n3306) );
  NAND U3609 ( .A(n9268), .B(n3306), .Z(n3145) );
  AND U3610 ( .A(n3146), .B(n3145), .Z(n3295) );
  NAND U3611 ( .A(n9046), .B(n3147), .Z(n3149) );
  XOR U3612 ( .A(b[19]), .B(a[15]), .Z(n3261) );
  NAND U3613 ( .A(n575), .B(n3261), .Z(n3148) );
  NAND U3614 ( .A(n3149), .B(n3148), .Z(n3294) );
  XOR U3615 ( .A(n3295), .B(n3294), .Z(n3297) );
  XOR U3616 ( .A(n3296), .B(n3297), .Z(n3223) );
  NAND U3617 ( .A(n573), .B(n3150), .Z(n3152) );
  XOR U3618 ( .A(b[15]), .B(a[19]), .Z(n3321) );
  NAND U3619 ( .A(n8694), .B(n3321), .Z(n3151) );
  AND U3620 ( .A(n3152), .B(n3151), .Z(n3266) );
  NAND U3621 ( .A(n583), .B(n3153), .Z(n3155) );
  XOR U3622 ( .A(b[29]), .B(a[5]), .Z(n3300) );
  NAND U3623 ( .A(n581), .B(n3300), .Z(n3154) );
  AND U3624 ( .A(n3155), .B(n3154), .Z(n3265) );
  AND U3625 ( .A(b[31]), .B(a[1]), .Z(n3264) );
  XOR U3626 ( .A(n3265), .B(n3264), .Z(n3267) );
  XNOR U3627 ( .A(n3266), .B(n3267), .Z(n3222) );
  XNOR U3628 ( .A(n3223), .B(n3222), .Z(n3225) );
  NANDN U3629 ( .A(n3157), .B(n3156), .Z(n3161) );
  OR U3630 ( .A(n3159), .B(n3158), .Z(n3160) );
  AND U3631 ( .A(n3161), .B(n3160), .Z(n3224) );
  XOR U3632 ( .A(n3225), .B(n3224), .Z(n3279) );
  NANDN U3633 ( .A(n3163), .B(n3162), .Z(n3167) );
  OR U3634 ( .A(n3165), .B(n3164), .Z(n3166) );
  AND U3635 ( .A(n3167), .B(n3166), .Z(n3277) );
  NANDN U3636 ( .A(n3169), .B(n3168), .Z(n3173) );
  NANDN U3637 ( .A(n3171), .B(n3170), .Z(n3172) );
  NAND U3638 ( .A(n3173), .B(n3172), .Z(n3276) );
  XNOR U3639 ( .A(n3277), .B(n3276), .Z(n3278) );
  XNOR U3640 ( .A(n3279), .B(n3278), .Z(n3212) );
  XOR U3641 ( .A(n3213), .B(n3212), .Z(n3331) );
  NAND U3642 ( .A(n3175), .B(n3174), .Z(n3179) );
  NAND U3643 ( .A(n3177), .B(n3176), .Z(n3178) );
  AND U3644 ( .A(n3179), .B(n3178), .Z(n3330) );
  XOR U3645 ( .A(n3331), .B(n3330), .Z(n3333) );
  XOR U3646 ( .A(n3332), .B(n3333), .Z(n3199) );
  XNOR U3647 ( .A(n3198), .B(n3199), .Z(n3200) );
  NANDN U3648 ( .A(n3181), .B(n3180), .Z(n3185) );
  NANDN U3649 ( .A(n3183), .B(n3182), .Z(n3184) );
  NAND U3650 ( .A(n3185), .B(n3184), .Z(n3201) );
  XNOR U3651 ( .A(n3200), .B(n3201), .Z(n3192) );
  NANDN U3652 ( .A(n3187), .B(n3186), .Z(n3191) );
  OR U3653 ( .A(n3189), .B(n3188), .Z(n3190) );
  NAND U3654 ( .A(n3191), .B(n3190), .Z(n3193) );
  XNOR U3655 ( .A(n3192), .B(n3193), .Z(n3194) );
  XNOR U3656 ( .A(n3195), .B(n3194), .Z(n3336) );
  XNOR U3657 ( .A(sreg[65]), .B(n3336), .Z(n3337) );
  XNOR U3658 ( .A(n3338), .B(n3337), .Z(c[65]) );
  NANDN U3659 ( .A(n3193), .B(n3192), .Z(n3197) );
  NANDN U3660 ( .A(n3195), .B(n3194), .Z(n3196) );
  AND U3661 ( .A(n3197), .B(n3196), .Z(n3344) );
  NANDN U3662 ( .A(n3199), .B(n3198), .Z(n3203) );
  NANDN U3663 ( .A(n3201), .B(n3200), .Z(n3202) );
  AND U3664 ( .A(n3203), .B(n3202), .Z(n3342) );
  NANDN U3665 ( .A(n3205), .B(n3204), .Z(n3209) );
  NANDN U3666 ( .A(n3207), .B(n3206), .Z(n3208) );
  AND U3667 ( .A(n3209), .B(n3208), .Z(n3350) );
  NANDN U3668 ( .A(n3211), .B(n3210), .Z(n3215) );
  NAND U3669 ( .A(n3213), .B(n3212), .Z(n3214) );
  AND U3670 ( .A(n3215), .B(n3214), .Z(n3476) );
  NANDN U3671 ( .A(n3217), .B(n3216), .Z(n3221) );
  NANDN U3672 ( .A(n3219), .B(n3218), .Z(n3220) );
  AND U3673 ( .A(n3221), .B(n3220), .Z(n3475) );
  XNOR U3674 ( .A(n3476), .B(n3475), .Z(n3478) );
  NANDN U3675 ( .A(n3223), .B(n3222), .Z(n3227) );
  NAND U3676 ( .A(n3225), .B(n3224), .Z(n3226) );
  AND U3677 ( .A(n3227), .B(n3226), .Z(n3359) );
  NANDN U3678 ( .A(n3229), .B(n3228), .Z(n3233) );
  OR U3679 ( .A(n3231), .B(n3230), .Z(n3232) );
  AND U3680 ( .A(n3233), .B(n3232), .Z(n3463) );
  NANDN U3681 ( .A(n3235), .B(n3234), .Z(n3239) );
  NANDN U3682 ( .A(n3237), .B(n3236), .Z(n3238) );
  NAND U3683 ( .A(n3239), .B(n3238), .Z(n3464) );
  XNOR U3684 ( .A(n3463), .B(n3464), .Z(n3465) );
  NANDN U3685 ( .A(n3241), .B(n3240), .Z(n3245) );
  NAND U3686 ( .A(n3243), .B(n3242), .Z(n3244) );
  NAND U3687 ( .A(n3245), .B(n3244), .Z(n3466) );
  XNOR U3688 ( .A(n3465), .B(n3466), .Z(n3357) );
  NAND U3689 ( .A(n9764), .B(n3246), .Z(n3248) );
  XOR U3690 ( .A(b[31]), .B(a[4]), .Z(n3378) );
  NAND U3691 ( .A(n584), .B(n3378), .Z(n3247) );
  AND U3692 ( .A(n3248), .B(n3247), .Z(n3389) );
  NAND U3693 ( .A(n568), .B(n3249), .Z(n3251) );
  XOR U3694 ( .A(b[3]), .B(a[32]), .Z(n3381) );
  NAND U3695 ( .A(n7245), .B(n3381), .Z(n3250) );
  AND U3696 ( .A(n3251), .B(n3250), .Z(n3388) );
  NAND U3697 ( .A(n576), .B(n3252), .Z(n3254) );
  XOR U3698 ( .A(b[17]), .B(a[18]), .Z(n3384) );
  NAND U3699 ( .A(n9141), .B(n3384), .Z(n3253) );
  NAND U3700 ( .A(n3254), .B(n3253), .Z(n3387) );
  XOR U3701 ( .A(n3388), .B(n3387), .Z(n3390) );
  XOR U3702 ( .A(n3389), .B(n3390), .Z(n3454) );
  NAND U3703 ( .A(n582), .B(n3255), .Z(n3257) );
  XOR U3704 ( .A(b[27]), .B(a[8]), .Z(n3369) );
  NAND U3705 ( .A(n9770), .B(n3369), .Z(n3256) );
  AND U3706 ( .A(n3257), .B(n3256), .Z(n3413) );
  NAND U3707 ( .A(n567), .B(n3258), .Z(n3260) );
  XOR U3708 ( .A(b[5]), .B(a[30]), .Z(n3372) );
  NAND U3709 ( .A(n7235), .B(n3372), .Z(n3259) );
  AND U3710 ( .A(n3260), .B(n3259), .Z(n3412) );
  NAND U3711 ( .A(n9046), .B(n3261), .Z(n3263) );
  XOR U3712 ( .A(b[19]), .B(a[16]), .Z(n3375) );
  NAND U3713 ( .A(n575), .B(n3375), .Z(n3262) );
  NAND U3714 ( .A(n3263), .B(n3262), .Z(n3411) );
  XOR U3715 ( .A(n3412), .B(n3411), .Z(n3414) );
  XNOR U3716 ( .A(n3413), .B(n3414), .Z(n3453) );
  XNOR U3717 ( .A(n3454), .B(n3453), .Z(n3455) );
  NANDN U3718 ( .A(n3265), .B(n3264), .Z(n3269) );
  OR U3719 ( .A(n3267), .B(n3266), .Z(n3268) );
  NAND U3720 ( .A(n3269), .B(n3268), .Z(n3456) );
  XOR U3721 ( .A(n3455), .B(n3456), .Z(n3358) );
  XOR U3722 ( .A(n3357), .B(n3358), .Z(n3360) );
  XOR U3723 ( .A(n3359), .B(n3360), .Z(n3472) );
  NANDN U3724 ( .A(n3271), .B(n3270), .Z(n3275) );
  NANDN U3725 ( .A(n3273), .B(n3272), .Z(n3274) );
  AND U3726 ( .A(n3275), .B(n3274), .Z(n3470) );
  NANDN U3727 ( .A(n3277), .B(n3276), .Z(n3281) );
  NANDN U3728 ( .A(n3279), .B(n3278), .Z(n3280) );
  AND U3729 ( .A(n3281), .B(n3280), .Z(n3356) );
  NANDN U3730 ( .A(n3283), .B(n3282), .Z(n3287) );
  OR U3731 ( .A(n3285), .B(n3284), .Z(n3286) );
  AND U3732 ( .A(n3287), .B(n3286), .Z(n3354) );
  NANDN U3733 ( .A(n3289), .B(n3288), .Z(n3293) );
  OR U3734 ( .A(n3291), .B(n3290), .Z(n3292) );
  AND U3735 ( .A(n3293), .B(n3292), .Z(n3460) );
  NANDN U3736 ( .A(n3295), .B(n3294), .Z(n3299) );
  OR U3737 ( .A(n3297), .B(n3296), .Z(n3298) );
  NAND U3738 ( .A(n3299), .B(n3298), .Z(n3459) );
  XNOR U3739 ( .A(n3460), .B(n3459), .Z(n3462) );
  NAND U3740 ( .A(n583), .B(n3300), .Z(n3302) );
  XOR U3741 ( .A(b[29]), .B(a[6]), .Z(n3426) );
  NAND U3742 ( .A(n581), .B(n3426), .Z(n3301) );
  AND U3743 ( .A(n3302), .B(n3301), .Z(n3364) );
  AND U3744 ( .A(b[31]), .B(a[2]), .Z(n3363) );
  XNOR U3745 ( .A(n3364), .B(n3363), .Z(n3365) );
  NAND U3746 ( .A(b[0]), .B(a[34]), .Z(n3303) );
  XNOR U3747 ( .A(b[1]), .B(n3303), .Z(n3305) );
  NANDN U3748 ( .A(b[0]), .B(a[33]), .Z(n3304) );
  NAND U3749 ( .A(n3305), .B(n3304), .Z(n3366) );
  XNOR U3750 ( .A(n3365), .B(n3366), .Z(n3406) );
  NAND U3751 ( .A(n578), .B(n3306), .Z(n3308) );
  XOR U3752 ( .A(b[23]), .B(a[12]), .Z(n3429) );
  NAND U3753 ( .A(n9268), .B(n3429), .Z(n3307) );
  AND U3754 ( .A(n3308), .B(n3307), .Z(n3419) );
  NAND U3755 ( .A(n569), .B(n3309), .Z(n3311) );
  XOR U3756 ( .A(b[7]), .B(a[28]), .Z(n3432) );
  NAND U3757 ( .A(n7819), .B(n3432), .Z(n3310) );
  AND U3758 ( .A(n3311), .B(n3310), .Z(n3418) );
  NAND U3759 ( .A(n579), .B(n3312), .Z(n3314) );
  XOR U3760 ( .A(b[25]), .B(a[10]), .Z(n3435) );
  NAND U3761 ( .A(n9364), .B(n3435), .Z(n3313) );
  NAND U3762 ( .A(n3314), .B(n3313), .Z(n3417) );
  XOR U3763 ( .A(n3418), .B(n3417), .Z(n3420) );
  XOR U3764 ( .A(n3419), .B(n3420), .Z(n3405) );
  XOR U3765 ( .A(n3406), .B(n3405), .Z(n3408) );
  NAND U3766 ( .A(n572), .B(n3315), .Z(n3317) );
  XOR U3767 ( .A(b[13]), .B(a[22]), .Z(n3438) );
  NAND U3768 ( .A(n8585), .B(n3438), .Z(n3316) );
  AND U3769 ( .A(n3317), .B(n3316), .Z(n3400) );
  NAND U3770 ( .A(n571), .B(n3318), .Z(n3320) );
  XOR U3771 ( .A(b[11]), .B(a[24]), .Z(n3441) );
  NAND U3772 ( .A(n8135), .B(n3441), .Z(n3319) );
  NAND U3773 ( .A(n3320), .B(n3319), .Z(n3399) );
  XNOR U3774 ( .A(n3400), .B(n3399), .Z(n3402) );
  NAND U3775 ( .A(n573), .B(n3321), .Z(n3323) );
  XOR U3776 ( .A(b[15]), .B(a[20]), .Z(n3444) );
  NAND U3777 ( .A(n8694), .B(n3444), .Z(n3322) );
  AND U3778 ( .A(n3323), .B(n3322), .Z(n3396) );
  NAND U3779 ( .A(n577), .B(n3324), .Z(n3326) );
  XOR U3780 ( .A(b[21]), .B(a[14]), .Z(n3447) );
  NAND U3781 ( .A(n9216), .B(n3447), .Z(n3325) );
  AND U3782 ( .A(n3326), .B(n3325), .Z(n3394) );
  NAND U3783 ( .A(n570), .B(n3327), .Z(n3329) );
  XOR U3784 ( .A(b[9]), .B(a[26]), .Z(n3450) );
  NAND U3785 ( .A(n8037), .B(n3450), .Z(n3328) );
  NAND U3786 ( .A(n3329), .B(n3328), .Z(n3393) );
  XNOR U3787 ( .A(n3394), .B(n3393), .Z(n3395) );
  XNOR U3788 ( .A(n3396), .B(n3395), .Z(n3401) );
  XOR U3789 ( .A(n3402), .B(n3401), .Z(n3407) );
  XNOR U3790 ( .A(n3408), .B(n3407), .Z(n3461) );
  XOR U3791 ( .A(n3462), .B(n3461), .Z(n3353) );
  XNOR U3792 ( .A(n3354), .B(n3353), .Z(n3355) );
  XNOR U3793 ( .A(n3356), .B(n3355), .Z(n3469) );
  XNOR U3794 ( .A(n3470), .B(n3469), .Z(n3471) );
  XNOR U3795 ( .A(n3472), .B(n3471), .Z(n3477) );
  XOR U3796 ( .A(n3478), .B(n3477), .Z(n3348) );
  NANDN U3797 ( .A(n3331), .B(n3330), .Z(n3335) );
  NANDN U3798 ( .A(n3333), .B(n3332), .Z(n3334) );
  NAND U3799 ( .A(n3335), .B(n3334), .Z(n3347) );
  XNOR U3800 ( .A(n3348), .B(n3347), .Z(n3349) );
  XNOR U3801 ( .A(n3350), .B(n3349), .Z(n3341) );
  XNOR U3802 ( .A(n3342), .B(n3341), .Z(n3343) );
  XNOR U3803 ( .A(n3344), .B(n3343), .Z(n3481) );
  XNOR U3804 ( .A(sreg[66]), .B(n3481), .Z(n3483) );
  NANDN U3805 ( .A(sreg[65]), .B(n3336), .Z(n3340) );
  NAND U3806 ( .A(n3338), .B(n3337), .Z(n3339) );
  NAND U3807 ( .A(n3340), .B(n3339), .Z(n3482) );
  XNOR U3808 ( .A(n3483), .B(n3482), .Z(c[66]) );
  NANDN U3809 ( .A(n3342), .B(n3341), .Z(n3346) );
  NANDN U3810 ( .A(n3344), .B(n3343), .Z(n3345) );
  AND U3811 ( .A(n3346), .B(n3345), .Z(n3491) );
  NANDN U3812 ( .A(n3348), .B(n3347), .Z(n3352) );
  NANDN U3813 ( .A(n3350), .B(n3349), .Z(n3351) );
  AND U3814 ( .A(n3352), .B(n3351), .Z(n3490) );
  NANDN U3815 ( .A(n3358), .B(n3357), .Z(n3362) );
  OR U3816 ( .A(n3360), .B(n3359), .Z(n3361) );
  AND U3817 ( .A(n3362), .B(n3361), .Z(n3627) );
  XNOR U3818 ( .A(n3628), .B(n3627), .Z(n3630) );
  NANDN U3819 ( .A(n3364), .B(n3363), .Z(n3368) );
  NANDN U3820 ( .A(n3366), .B(n3365), .Z(n3367) );
  AND U3821 ( .A(n3368), .B(n3367), .Z(n3575) );
  NAND U3822 ( .A(n582), .B(n3369), .Z(n3371) );
  XOR U3823 ( .A(b[27]), .B(a[9]), .Z(n3519) );
  NAND U3824 ( .A(n9770), .B(n3519), .Z(n3370) );
  AND U3825 ( .A(n3371), .B(n3370), .Z(n3582) );
  NAND U3826 ( .A(n567), .B(n3372), .Z(n3374) );
  XOR U3827 ( .A(b[5]), .B(a[31]), .Z(n3522) );
  NAND U3828 ( .A(n7235), .B(n3522), .Z(n3373) );
  AND U3829 ( .A(n3374), .B(n3373), .Z(n3580) );
  NAND U3830 ( .A(n9046), .B(n3375), .Z(n3377) );
  XOR U3831 ( .A(b[19]), .B(a[17]), .Z(n3525) );
  NAND U3832 ( .A(n575), .B(n3525), .Z(n3376) );
  NAND U3833 ( .A(n3377), .B(n3376), .Z(n3579) );
  XNOR U3834 ( .A(n3580), .B(n3579), .Z(n3581) );
  XNOR U3835 ( .A(n3582), .B(n3581), .Z(n3573) );
  NAND U3836 ( .A(n9764), .B(n3378), .Z(n3380) );
  XOR U3837 ( .A(b[31]), .B(a[5]), .Z(n3528) );
  NAND U3838 ( .A(n584), .B(n3528), .Z(n3379) );
  AND U3839 ( .A(n3380), .B(n3379), .Z(n3540) );
  NAND U3840 ( .A(n568), .B(n3381), .Z(n3383) );
  XOR U3841 ( .A(b[3]), .B(a[33]), .Z(n3531) );
  NAND U3842 ( .A(n7245), .B(n3531), .Z(n3382) );
  AND U3843 ( .A(n3383), .B(n3382), .Z(n3538) );
  NAND U3844 ( .A(n576), .B(n3384), .Z(n3386) );
  XOR U3845 ( .A(b[17]), .B(a[19]), .Z(n3534) );
  NAND U3846 ( .A(n9141), .B(n3534), .Z(n3385) );
  NAND U3847 ( .A(n3386), .B(n3385), .Z(n3537) );
  XNOR U3848 ( .A(n3538), .B(n3537), .Z(n3539) );
  XOR U3849 ( .A(n3540), .B(n3539), .Z(n3574) );
  XOR U3850 ( .A(n3573), .B(n3574), .Z(n3576) );
  XOR U3851 ( .A(n3575), .B(n3576), .Z(n3508) );
  NANDN U3852 ( .A(n3388), .B(n3387), .Z(n3392) );
  OR U3853 ( .A(n3390), .B(n3389), .Z(n3391) );
  AND U3854 ( .A(n3392), .B(n3391), .Z(n3561) );
  NANDN U3855 ( .A(n3394), .B(n3393), .Z(n3398) );
  NANDN U3856 ( .A(n3396), .B(n3395), .Z(n3397) );
  NAND U3857 ( .A(n3398), .B(n3397), .Z(n3562) );
  XNOR U3858 ( .A(n3561), .B(n3562), .Z(n3563) );
  NANDN U3859 ( .A(n3400), .B(n3399), .Z(n3404) );
  NAND U3860 ( .A(n3402), .B(n3401), .Z(n3403) );
  NAND U3861 ( .A(n3404), .B(n3403), .Z(n3564) );
  XNOR U3862 ( .A(n3563), .B(n3564), .Z(n3507) );
  XNOR U3863 ( .A(n3508), .B(n3507), .Z(n3510) );
  NAND U3864 ( .A(n3406), .B(n3405), .Z(n3410) );
  NAND U3865 ( .A(n3408), .B(n3407), .Z(n3409) );
  AND U3866 ( .A(n3410), .B(n3409), .Z(n3509) );
  XOR U3867 ( .A(n3510), .B(n3509), .Z(n3624) );
  NANDN U3868 ( .A(n3412), .B(n3411), .Z(n3416) );
  OR U3869 ( .A(n3414), .B(n3413), .Z(n3415) );
  AND U3870 ( .A(n3416), .B(n3415), .Z(n3568) );
  NANDN U3871 ( .A(n3418), .B(n3417), .Z(n3422) );
  OR U3872 ( .A(n3420), .B(n3419), .Z(n3421) );
  NAND U3873 ( .A(n3422), .B(n3421), .Z(n3567) );
  XNOR U3874 ( .A(n3568), .B(n3567), .Z(n3570) );
  NAND U3875 ( .A(b[0]), .B(a[35]), .Z(n3423) );
  XNOR U3876 ( .A(b[1]), .B(n3423), .Z(n3425) );
  NANDN U3877 ( .A(b[0]), .B(a[34]), .Z(n3424) );
  NAND U3878 ( .A(n3425), .B(n3424), .Z(n3516) );
  NAND U3879 ( .A(n583), .B(n3426), .Z(n3428) );
  XOR U3880 ( .A(b[29]), .B(a[7]), .Z(n3594) );
  NAND U3881 ( .A(n581), .B(n3594), .Z(n3427) );
  AND U3882 ( .A(n3428), .B(n3427), .Z(n3514) );
  AND U3883 ( .A(b[31]), .B(a[3]), .Z(n3513) );
  XNOR U3884 ( .A(n3514), .B(n3513), .Z(n3515) );
  XNOR U3885 ( .A(n3516), .B(n3515), .Z(n3555) );
  NAND U3886 ( .A(n578), .B(n3429), .Z(n3431) );
  XOR U3887 ( .A(b[23]), .B(a[13]), .Z(n3597) );
  NAND U3888 ( .A(n9268), .B(n3597), .Z(n3430) );
  AND U3889 ( .A(n3431), .B(n3430), .Z(n3588) );
  NAND U3890 ( .A(n569), .B(n3432), .Z(n3434) );
  XOR U3891 ( .A(b[7]), .B(a[29]), .Z(n3600) );
  NAND U3892 ( .A(n7819), .B(n3600), .Z(n3433) );
  AND U3893 ( .A(n3434), .B(n3433), .Z(n3586) );
  NAND U3894 ( .A(n579), .B(n3435), .Z(n3437) );
  XOR U3895 ( .A(b[25]), .B(a[11]), .Z(n3603) );
  NAND U3896 ( .A(n9364), .B(n3603), .Z(n3436) );
  NAND U3897 ( .A(n3437), .B(n3436), .Z(n3585) );
  XNOR U3898 ( .A(n3586), .B(n3585), .Z(n3587) );
  XOR U3899 ( .A(n3588), .B(n3587), .Z(n3556) );
  XNOR U3900 ( .A(n3555), .B(n3556), .Z(n3557) );
  NAND U3901 ( .A(n572), .B(n3438), .Z(n3440) );
  XOR U3902 ( .A(b[13]), .B(a[23]), .Z(n3606) );
  NAND U3903 ( .A(n8585), .B(n3606), .Z(n3439) );
  AND U3904 ( .A(n3440), .B(n3439), .Z(n3550) );
  NAND U3905 ( .A(n571), .B(n3441), .Z(n3443) );
  XOR U3906 ( .A(b[11]), .B(a[25]), .Z(n3609) );
  NAND U3907 ( .A(n8135), .B(n3609), .Z(n3442) );
  NAND U3908 ( .A(n3443), .B(n3442), .Z(n3549) );
  XNOR U3909 ( .A(n3550), .B(n3549), .Z(n3551) );
  NAND U3910 ( .A(n573), .B(n3444), .Z(n3446) );
  XOR U3911 ( .A(b[15]), .B(a[21]), .Z(n3612) );
  NAND U3912 ( .A(n8694), .B(n3612), .Z(n3445) );
  AND U3913 ( .A(n3446), .B(n3445), .Z(n3546) );
  NAND U3914 ( .A(n577), .B(n3447), .Z(n3449) );
  XOR U3915 ( .A(b[21]), .B(a[15]), .Z(n3615) );
  NAND U3916 ( .A(n9216), .B(n3615), .Z(n3448) );
  AND U3917 ( .A(n3449), .B(n3448), .Z(n3544) );
  NAND U3918 ( .A(n570), .B(n3450), .Z(n3452) );
  XOR U3919 ( .A(b[9]), .B(a[27]), .Z(n3618) );
  NAND U3920 ( .A(n8037), .B(n3618), .Z(n3451) );
  NAND U3921 ( .A(n3452), .B(n3451), .Z(n3543) );
  XNOR U3922 ( .A(n3544), .B(n3543), .Z(n3545) );
  XOR U3923 ( .A(n3546), .B(n3545), .Z(n3552) );
  XOR U3924 ( .A(n3551), .B(n3552), .Z(n3558) );
  XNOR U3925 ( .A(n3557), .B(n3558), .Z(n3569) );
  XOR U3926 ( .A(n3570), .B(n3569), .Z(n3502) );
  NANDN U3927 ( .A(n3454), .B(n3453), .Z(n3458) );
  NANDN U3928 ( .A(n3456), .B(n3455), .Z(n3457) );
  NAND U3929 ( .A(n3458), .B(n3457), .Z(n3501) );
  XNOR U3930 ( .A(n3502), .B(n3501), .Z(n3504) );
  XOR U3931 ( .A(n3504), .B(n3503), .Z(n3622) );
  NANDN U3932 ( .A(n3464), .B(n3463), .Z(n3468) );
  NANDN U3933 ( .A(n3466), .B(n3465), .Z(n3467) );
  AND U3934 ( .A(n3468), .B(n3467), .Z(n3621) );
  XNOR U3935 ( .A(n3622), .B(n3621), .Z(n3623) );
  XNOR U3936 ( .A(n3624), .B(n3623), .Z(n3629) );
  XOR U3937 ( .A(n3630), .B(n3629), .Z(n3496) );
  NANDN U3938 ( .A(n3470), .B(n3469), .Z(n3474) );
  NANDN U3939 ( .A(n3472), .B(n3471), .Z(n3473) );
  AND U3940 ( .A(n3474), .B(n3473), .Z(n3495) );
  XNOR U3941 ( .A(n3496), .B(n3495), .Z(n3497) );
  NANDN U3942 ( .A(n3476), .B(n3475), .Z(n3480) );
  NAND U3943 ( .A(n3478), .B(n3477), .Z(n3479) );
  NAND U3944 ( .A(n3480), .B(n3479), .Z(n3498) );
  XNOR U3945 ( .A(n3497), .B(n3498), .Z(n3489) );
  XOR U3946 ( .A(n3490), .B(n3489), .Z(n3492) );
  XNOR U3947 ( .A(n3491), .B(n3492), .Z(n3487) );
  NANDN U3948 ( .A(sreg[66]), .B(n3481), .Z(n3485) );
  NAND U3949 ( .A(n3483), .B(n3482), .Z(n3484) );
  AND U3950 ( .A(n3485), .B(n3484), .Z(n3488) );
  XNOR U3951 ( .A(sreg[67]), .B(n3488), .Z(n3486) );
  XNOR U3952 ( .A(n3487), .B(n3486), .Z(c[67]) );
  NANDN U3953 ( .A(n3490), .B(n3489), .Z(n3494) );
  OR U3954 ( .A(n3492), .B(n3491), .Z(n3493) );
  AND U3955 ( .A(n3494), .B(n3493), .Z(n3636) );
  NANDN U3956 ( .A(n3496), .B(n3495), .Z(n3500) );
  NANDN U3957 ( .A(n3498), .B(n3497), .Z(n3499) );
  AND U3958 ( .A(n3500), .B(n3499), .Z(n3634) );
  NANDN U3959 ( .A(n3502), .B(n3501), .Z(n3506) );
  NAND U3960 ( .A(n3504), .B(n3503), .Z(n3505) );
  AND U3961 ( .A(n3506), .B(n3505), .Z(n3771) );
  NANDN U3962 ( .A(n3508), .B(n3507), .Z(n3512) );
  NAND U3963 ( .A(n3510), .B(n3509), .Z(n3511) );
  NAND U3964 ( .A(n3512), .B(n3511), .Z(n3772) );
  XNOR U3965 ( .A(n3771), .B(n3772), .Z(n3774) );
  NANDN U3966 ( .A(n3514), .B(n3513), .Z(n3518) );
  NANDN U3967 ( .A(n3516), .B(n3515), .Z(n3517) );
  AND U3968 ( .A(n3518), .B(n3517), .Z(n3719) );
  NAND U3969 ( .A(n582), .B(n3519), .Z(n3521) );
  XOR U3970 ( .A(b[27]), .B(a[10]), .Z(n3663) );
  NAND U3971 ( .A(n9770), .B(n3663), .Z(n3520) );
  AND U3972 ( .A(n3521), .B(n3520), .Z(n3726) );
  NAND U3973 ( .A(n567), .B(n3522), .Z(n3524) );
  XOR U3974 ( .A(b[5]), .B(a[32]), .Z(n3666) );
  NAND U3975 ( .A(n7235), .B(n3666), .Z(n3523) );
  AND U3976 ( .A(n3524), .B(n3523), .Z(n3724) );
  NAND U3977 ( .A(n9046), .B(n3525), .Z(n3527) );
  XOR U3978 ( .A(b[19]), .B(a[18]), .Z(n3669) );
  NAND U3979 ( .A(n575), .B(n3669), .Z(n3526) );
  NAND U3980 ( .A(n3527), .B(n3526), .Z(n3723) );
  XNOR U3981 ( .A(n3724), .B(n3723), .Z(n3725) );
  XNOR U3982 ( .A(n3726), .B(n3725), .Z(n3717) );
  NAND U3983 ( .A(n9764), .B(n3528), .Z(n3530) );
  XOR U3984 ( .A(b[31]), .B(a[6]), .Z(n3672) );
  NAND U3985 ( .A(n584), .B(n3672), .Z(n3529) );
  AND U3986 ( .A(n3530), .B(n3529), .Z(n3684) );
  NAND U3987 ( .A(n568), .B(n3531), .Z(n3533) );
  XOR U3988 ( .A(b[3]), .B(a[34]), .Z(n3675) );
  NAND U3989 ( .A(n7245), .B(n3675), .Z(n3532) );
  AND U3990 ( .A(n3533), .B(n3532), .Z(n3682) );
  NAND U3991 ( .A(n576), .B(n3534), .Z(n3536) );
  XOR U3992 ( .A(b[17]), .B(a[20]), .Z(n3678) );
  NAND U3993 ( .A(n9141), .B(n3678), .Z(n3535) );
  NAND U3994 ( .A(n3536), .B(n3535), .Z(n3681) );
  XNOR U3995 ( .A(n3682), .B(n3681), .Z(n3683) );
  XOR U3996 ( .A(n3684), .B(n3683), .Z(n3718) );
  XOR U3997 ( .A(n3717), .B(n3718), .Z(n3720) );
  XOR U3998 ( .A(n3719), .B(n3720), .Z(n3652) );
  NANDN U3999 ( .A(n3538), .B(n3537), .Z(n3542) );
  NANDN U4000 ( .A(n3540), .B(n3539), .Z(n3541) );
  AND U4001 ( .A(n3542), .B(n3541), .Z(n3705) );
  NANDN U4002 ( .A(n3544), .B(n3543), .Z(n3548) );
  NANDN U4003 ( .A(n3546), .B(n3545), .Z(n3547) );
  NAND U4004 ( .A(n3548), .B(n3547), .Z(n3706) );
  XNOR U4005 ( .A(n3705), .B(n3706), .Z(n3707) );
  NANDN U4006 ( .A(n3550), .B(n3549), .Z(n3554) );
  NANDN U4007 ( .A(n3552), .B(n3551), .Z(n3553) );
  NAND U4008 ( .A(n3554), .B(n3553), .Z(n3708) );
  XNOR U4009 ( .A(n3707), .B(n3708), .Z(n3651) );
  XNOR U4010 ( .A(n3652), .B(n3651), .Z(n3654) );
  NANDN U4011 ( .A(n3556), .B(n3555), .Z(n3560) );
  NANDN U4012 ( .A(n3558), .B(n3557), .Z(n3559) );
  AND U4013 ( .A(n3560), .B(n3559), .Z(n3653) );
  XOR U4014 ( .A(n3654), .B(n3653), .Z(n3768) );
  NANDN U4015 ( .A(n3562), .B(n3561), .Z(n3566) );
  NANDN U4016 ( .A(n3564), .B(n3563), .Z(n3565) );
  AND U4017 ( .A(n3566), .B(n3565), .Z(n3765) );
  NANDN U4018 ( .A(n3568), .B(n3567), .Z(n3572) );
  NAND U4019 ( .A(n3570), .B(n3569), .Z(n3571) );
  AND U4020 ( .A(n3572), .B(n3571), .Z(n3648) );
  NANDN U4021 ( .A(n3574), .B(n3573), .Z(n3578) );
  OR U4022 ( .A(n3576), .B(n3575), .Z(n3577) );
  AND U4023 ( .A(n3578), .B(n3577), .Z(n3646) );
  NANDN U4024 ( .A(n3580), .B(n3579), .Z(n3584) );
  NANDN U4025 ( .A(n3582), .B(n3581), .Z(n3583) );
  AND U4026 ( .A(n3584), .B(n3583), .Z(n3712) );
  NANDN U4027 ( .A(n3586), .B(n3585), .Z(n3590) );
  NANDN U4028 ( .A(n3588), .B(n3587), .Z(n3589) );
  NAND U4029 ( .A(n3590), .B(n3589), .Z(n3711) );
  XNOR U4030 ( .A(n3712), .B(n3711), .Z(n3713) );
  NAND U4031 ( .A(b[0]), .B(a[36]), .Z(n3591) );
  XNOR U4032 ( .A(b[1]), .B(n3591), .Z(n3593) );
  NANDN U4033 ( .A(b[0]), .B(a[35]), .Z(n3592) );
  NAND U4034 ( .A(n3593), .B(n3592), .Z(n3660) );
  NAND U4035 ( .A(n583), .B(n3594), .Z(n3596) );
  XOR U4036 ( .A(b[29]), .B(a[8]), .Z(n3735) );
  NAND U4037 ( .A(n581), .B(n3735), .Z(n3595) );
  AND U4038 ( .A(n3596), .B(n3595), .Z(n3658) );
  AND U4039 ( .A(b[31]), .B(a[4]), .Z(n3657) );
  XNOR U4040 ( .A(n3658), .B(n3657), .Z(n3659) );
  XNOR U4041 ( .A(n3660), .B(n3659), .Z(n3699) );
  NAND U4042 ( .A(n578), .B(n3597), .Z(n3599) );
  XOR U4043 ( .A(b[23]), .B(a[14]), .Z(n3741) );
  NAND U4044 ( .A(n9268), .B(n3741), .Z(n3598) );
  AND U4045 ( .A(n3599), .B(n3598), .Z(n3732) );
  NAND U4046 ( .A(n569), .B(n3600), .Z(n3602) );
  XOR U4047 ( .A(b[7]), .B(a[30]), .Z(n3744) );
  NAND U4048 ( .A(n7819), .B(n3744), .Z(n3601) );
  AND U4049 ( .A(n3602), .B(n3601), .Z(n3730) );
  NAND U4050 ( .A(n579), .B(n3603), .Z(n3605) );
  XOR U4051 ( .A(b[25]), .B(a[12]), .Z(n3747) );
  NAND U4052 ( .A(n9364), .B(n3747), .Z(n3604) );
  NAND U4053 ( .A(n3605), .B(n3604), .Z(n3729) );
  XNOR U4054 ( .A(n3730), .B(n3729), .Z(n3731) );
  XOR U4055 ( .A(n3732), .B(n3731), .Z(n3700) );
  XNOR U4056 ( .A(n3699), .B(n3700), .Z(n3701) );
  NAND U4057 ( .A(n572), .B(n3606), .Z(n3608) );
  XOR U4058 ( .A(b[13]), .B(a[24]), .Z(n3750) );
  NAND U4059 ( .A(n8585), .B(n3750), .Z(n3607) );
  AND U4060 ( .A(n3608), .B(n3607), .Z(n3694) );
  NAND U4061 ( .A(n571), .B(n3609), .Z(n3611) );
  XOR U4062 ( .A(b[11]), .B(a[26]), .Z(n3753) );
  NAND U4063 ( .A(n8135), .B(n3753), .Z(n3610) );
  NAND U4064 ( .A(n3611), .B(n3610), .Z(n3693) );
  XNOR U4065 ( .A(n3694), .B(n3693), .Z(n3695) );
  NAND U4066 ( .A(n573), .B(n3612), .Z(n3614) );
  XOR U4067 ( .A(b[15]), .B(a[22]), .Z(n3756) );
  NAND U4068 ( .A(n8694), .B(n3756), .Z(n3613) );
  AND U4069 ( .A(n3614), .B(n3613), .Z(n3690) );
  NAND U4070 ( .A(n577), .B(n3615), .Z(n3617) );
  XOR U4071 ( .A(b[21]), .B(a[16]), .Z(n3759) );
  NAND U4072 ( .A(n9216), .B(n3759), .Z(n3616) );
  AND U4073 ( .A(n3617), .B(n3616), .Z(n3688) );
  NAND U4074 ( .A(n570), .B(n3618), .Z(n3620) );
  XOR U4075 ( .A(b[9]), .B(a[28]), .Z(n3762) );
  NAND U4076 ( .A(n8037), .B(n3762), .Z(n3619) );
  NAND U4077 ( .A(n3620), .B(n3619), .Z(n3687) );
  XNOR U4078 ( .A(n3688), .B(n3687), .Z(n3689) );
  XOR U4079 ( .A(n3690), .B(n3689), .Z(n3696) );
  XOR U4080 ( .A(n3695), .B(n3696), .Z(n3702) );
  XOR U4081 ( .A(n3701), .B(n3702), .Z(n3714) );
  XNOR U4082 ( .A(n3713), .B(n3714), .Z(n3645) );
  XNOR U4083 ( .A(n3646), .B(n3645), .Z(n3647) );
  XOR U4084 ( .A(n3648), .B(n3647), .Z(n3766) );
  XNOR U4085 ( .A(n3765), .B(n3766), .Z(n3767) );
  XNOR U4086 ( .A(n3768), .B(n3767), .Z(n3773) );
  XOR U4087 ( .A(n3774), .B(n3773), .Z(n3640) );
  NANDN U4088 ( .A(n3622), .B(n3621), .Z(n3626) );
  NANDN U4089 ( .A(n3624), .B(n3623), .Z(n3625) );
  AND U4090 ( .A(n3626), .B(n3625), .Z(n3639) );
  XNOR U4091 ( .A(n3640), .B(n3639), .Z(n3641) );
  NANDN U4092 ( .A(n3628), .B(n3627), .Z(n3632) );
  NAND U4093 ( .A(n3630), .B(n3629), .Z(n3631) );
  NAND U4094 ( .A(n3632), .B(n3631), .Z(n3642) );
  XNOR U4095 ( .A(n3641), .B(n3642), .Z(n3633) );
  XNOR U4096 ( .A(n3634), .B(n3633), .Z(n3635) );
  XNOR U4097 ( .A(n3636), .B(n3635), .Z(n3777) );
  XNOR U4098 ( .A(sreg[68]), .B(n3777), .Z(n3778) );
  XOR U4099 ( .A(n3779), .B(n3778), .Z(c[68]) );
  NANDN U4100 ( .A(n3634), .B(n3633), .Z(n3638) );
  NANDN U4101 ( .A(n3636), .B(n3635), .Z(n3637) );
  AND U4102 ( .A(n3638), .B(n3637), .Z(n3785) );
  NANDN U4103 ( .A(n3640), .B(n3639), .Z(n3644) );
  NANDN U4104 ( .A(n3642), .B(n3641), .Z(n3643) );
  AND U4105 ( .A(n3644), .B(n3643), .Z(n3783) );
  NANDN U4106 ( .A(n3646), .B(n3645), .Z(n3650) );
  NANDN U4107 ( .A(n3648), .B(n3647), .Z(n3649) );
  AND U4108 ( .A(n3650), .B(n3649), .Z(n3921) );
  NANDN U4109 ( .A(n3652), .B(n3651), .Z(n3656) );
  NAND U4110 ( .A(n3654), .B(n3653), .Z(n3655) );
  AND U4111 ( .A(n3656), .B(n3655), .Z(n3920) );
  XNOR U4112 ( .A(n3921), .B(n3920), .Z(n3923) );
  NANDN U4113 ( .A(n3658), .B(n3657), .Z(n3662) );
  NANDN U4114 ( .A(n3660), .B(n3659), .Z(n3661) );
  AND U4115 ( .A(n3662), .B(n3661), .Z(n3868) );
  NAND U4116 ( .A(n582), .B(n3663), .Z(n3665) );
  XOR U4117 ( .A(b[27]), .B(a[11]), .Z(n3812) );
  NAND U4118 ( .A(n9770), .B(n3812), .Z(n3664) );
  AND U4119 ( .A(n3665), .B(n3664), .Z(n3875) );
  NAND U4120 ( .A(n567), .B(n3666), .Z(n3668) );
  XOR U4121 ( .A(b[5]), .B(a[33]), .Z(n3815) );
  NAND U4122 ( .A(n7235), .B(n3815), .Z(n3667) );
  AND U4123 ( .A(n3668), .B(n3667), .Z(n3873) );
  NAND U4124 ( .A(n9046), .B(n3669), .Z(n3671) );
  XOR U4125 ( .A(b[19]), .B(a[19]), .Z(n3818) );
  NAND U4126 ( .A(n575), .B(n3818), .Z(n3670) );
  NAND U4127 ( .A(n3671), .B(n3670), .Z(n3872) );
  XNOR U4128 ( .A(n3873), .B(n3872), .Z(n3874) );
  XNOR U4129 ( .A(n3875), .B(n3874), .Z(n3866) );
  NAND U4130 ( .A(n9764), .B(n3672), .Z(n3674) );
  XOR U4131 ( .A(b[31]), .B(a[7]), .Z(n3821) );
  NAND U4132 ( .A(n584), .B(n3821), .Z(n3673) );
  AND U4133 ( .A(n3674), .B(n3673), .Z(n3833) );
  NAND U4134 ( .A(n568), .B(n3675), .Z(n3677) );
  XOR U4135 ( .A(b[3]), .B(a[35]), .Z(n3824) );
  NAND U4136 ( .A(n7245), .B(n3824), .Z(n3676) );
  AND U4137 ( .A(n3677), .B(n3676), .Z(n3831) );
  NAND U4138 ( .A(n576), .B(n3678), .Z(n3680) );
  XOR U4139 ( .A(b[17]), .B(a[21]), .Z(n3827) );
  NAND U4140 ( .A(n9141), .B(n3827), .Z(n3679) );
  NAND U4141 ( .A(n3680), .B(n3679), .Z(n3830) );
  XNOR U4142 ( .A(n3831), .B(n3830), .Z(n3832) );
  XOR U4143 ( .A(n3833), .B(n3832), .Z(n3867) );
  XOR U4144 ( .A(n3866), .B(n3867), .Z(n3869) );
  XOR U4145 ( .A(n3868), .B(n3869), .Z(n3801) );
  NANDN U4146 ( .A(n3682), .B(n3681), .Z(n3686) );
  NANDN U4147 ( .A(n3684), .B(n3683), .Z(n3685) );
  AND U4148 ( .A(n3686), .B(n3685), .Z(n3854) );
  NANDN U4149 ( .A(n3688), .B(n3687), .Z(n3692) );
  NANDN U4150 ( .A(n3690), .B(n3689), .Z(n3691) );
  NAND U4151 ( .A(n3692), .B(n3691), .Z(n3855) );
  XNOR U4152 ( .A(n3854), .B(n3855), .Z(n3856) );
  NANDN U4153 ( .A(n3694), .B(n3693), .Z(n3698) );
  NANDN U4154 ( .A(n3696), .B(n3695), .Z(n3697) );
  NAND U4155 ( .A(n3698), .B(n3697), .Z(n3857) );
  XNOR U4156 ( .A(n3856), .B(n3857), .Z(n3800) );
  XNOR U4157 ( .A(n3801), .B(n3800), .Z(n3803) );
  NANDN U4158 ( .A(n3700), .B(n3699), .Z(n3704) );
  NANDN U4159 ( .A(n3702), .B(n3701), .Z(n3703) );
  AND U4160 ( .A(n3704), .B(n3703), .Z(n3802) );
  XOR U4161 ( .A(n3803), .B(n3802), .Z(n3917) );
  NANDN U4162 ( .A(n3706), .B(n3705), .Z(n3710) );
  NANDN U4163 ( .A(n3708), .B(n3707), .Z(n3709) );
  AND U4164 ( .A(n3710), .B(n3709), .Z(n3914) );
  NANDN U4165 ( .A(n3712), .B(n3711), .Z(n3716) );
  NANDN U4166 ( .A(n3714), .B(n3713), .Z(n3715) );
  AND U4167 ( .A(n3716), .B(n3715), .Z(n3797) );
  NANDN U4168 ( .A(n3718), .B(n3717), .Z(n3722) );
  OR U4169 ( .A(n3720), .B(n3719), .Z(n3721) );
  AND U4170 ( .A(n3722), .B(n3721), .Z(n3795) );
  NANDN U4171 ( .A(n3724), .B(n3723), .Z(n3728) );
  NANDN U4172 ( .A(n3726), .B(n3725), .Z(n3727) );
  AND U4173 ( .A(n3728), .B(n3727), .Z(n3861) );
  NANDN U4174 ( .A(n3730), .B(n3729), .Z(n3734) );
  NANDN U4175 ( .A(n3732), .B(n3731), .Z(n3733) );
  NAND U4176 ( .A(n3734), .B(n3733), .Z(n3860) );
  XNOR U4177 ( .A(n3861), .B(n3860), .Z(n3862) );
  NAND U4178 ( .A(n583), .B(n3735), .Z(n3737) );
  XOR U4179 ( .A(b[29]), .B(a[9]), .Z(n3887) );
  NAND U4180 ( .A(n581), .B(n3887), .Z(n3736) );
  AND U4181 ( .A(n3737), .B(n3736), .Z(n3807) );
  AND U4182 ( .A(b[31]), .B(a[5]), .Z(n3806) );
  XNOR U4183 ( .A(n3807), .B(n3806), .Z(n3808) );
  NAND U4184 ( .A(b[0]), .B(a[37]), .Z(n3738) );
  XNOR U4185 ( .A(b[1]), .B(n3738), .Z(n3740) );
  NANDN U4186 ( .A(b[0]), .B(a[36]), .Z(n3739) );
  NAND U4187 ( .A(n3740), .B(n3739), .Z(n3809) );
  XNOR U4188 ( .A(n3808), .B(n3809), .Z(n3848) );
  NAND U4189 ( .A(n578), .B(n3741), .Z(n3743) );
  XOR U4190 ( .A(b[23]), .B(a[15]), .Z(n3890) );
  NAND U4191 ( .A(n9268), .B(n3890), .Z(n3742) );
  AND U4192 ( .A(n3743), .B(n3742), .Z(n3881) );
  NAND U4193 ( .A(n569), .B(n3744), .Z(n3746) );
  XOR U4194 ( .A(b[7]), .B(a[31]), .Z(n3893) );
  NAND U4195 ( .A(n7819), .B(n3893), .Z(n3745) );
  AND U4196 ( .A(n3746), .B(n3745), .Z(n3879) );
  NAND U4197 ( .A(n579), .B(n3747), .Z(n3749) );
  XOR U4198 ( .A(b[25]), .B(a[13]), .Z(n3896) );
  NAND U4199 ( .A(n9364), .B(n3896), .Z(n3748) );
  NAND U4200 ( .A(n3749), .B(n3748), .Z(n3878) );
  XNOR U4201 ( .A(n3879), .B(n3878), .Z(n3880) );
  XOR U4202 ( .A(n3881), .B(n3880), .Z(n3849) );
  XNOR U4203 ( .A(n3848), .B(n3849), .Z(n3850) );
  NAND U4204 ( .A(n572), .B(n3750), .Z(n3752) );
  XOR U4205 ( .A(b[13]), .B(a[25]), .Z(n3899) );
  NAND U4206 ( .A(n8585), .B(n3899), .Z(n3751) );
  AND U4207 ( .A(n3752), .B(n3751), .Z(n3843) );
  NAND U4208 ( .A(n571), .B(n3753), .Z(n3755) );
  XOR U4209 ( .A(b[11]), .B(a[27]), .Z(n3902) );
  NAND U4210 ( .A(n8135), .B(n3902), .Z(n3754) );
  NAND U4211 ( .A(n3755), .B(n3754), .Z(n3842) );
  XNOR U4212 ( .A(n3843), .B(n3842), .Z(n3844) );
  NAND U4213 ( .A(n573), .B(n3756), .Z(n3758) );
  XOR U4214 ( .A(b[15]), .B(a[23]), .Z(n3905) );
  NAND U4215 ( .A(n8694), .B(n3905), .Z(n3757) );
  AND U4216 ( .A(n3758), .B(n3757), .Z(n3839) );
  NAND U4217 ( .A(n577), .B(n3759), .Z(n3761) );
  XOR U4218 ( .A(b[21]), .B(a[17]), .Z(n3908) );
  NAND U4219 ( .A(n9216), .B(n3908), .Z(n3760) );
  AND U4220 ( .A(n3761), .B(n3760), .Z(n3837) );
  NAND U4221 ( .A(n570), .B(n3762), .Z(n3764) );
  XOR U4222 ( .A(b[9]), .B(a[29]), .Z(n3911) );
  NAND U4223 ( .A(n8037), .B(n3911), .Z(n3763) );
  NAND U4224 ( .A(n3764), .B(n3763), .Z(n3836) );
  XNOR U4225 ( .A(n3837), .B(n3836), .Z(n3838) );
  XOR U4226 ( .A(n3839), .B(n3838), .Z(n3845) );
  XOR U4227 ( .A(n3844), .B(n3845), .Z(n3851) );
  XOR U4228 ( .A(n3850), .B(n3851), .Z(n3863) );
  XNOR U4229 ( .A(n3862), .B(n3863), .Z(n3794) );
  XNOR U4230 ( .A(n3795), .B(n3794), .Z(n3796) );
  XOR U4231 ( .A(n3797), .B(n3796), .Z(n3915) );
  XNOR U4232 ( .A(n3914), .B(n3915), .Z(n3916) );
  XNOR U4233 ( .A(n3917), .B(n3916), .Z(n3922) );
  XOR U4234 ( .A(n3923), .B(n3922), .Z(n3789) );
  NANDN U4235 ( .A(n3766), .B(n3765), .Z(n3770) );
  NANDN U4236 ( .A(n3768), .B(n3767), .Z(n3769) );
  AND U4237 ( .A(n3770), .B(n3769), .Z(n3788) );
  XNOR U4238 ( .A(n3789), .B(n3788), .Z(n3790) );
  NANDN U4239 ( .A(n3772), .B(n3771), .Z(n3776) );
  NAND U4240 ( .A(n3774), .B(n3773), .Z(n3775) );
  NAND U4241 ( .A(n3776), .B(n3775), .Z(n3791) );
  XNOR U4242 ( .A(n3790), .B(n3791), .Z(n3782) );
  XNOR U4243 ( .A(n3783), .B(n3782), .Z(n3784) );
  XNOR U4244 ( .A(n3785), .B(n3784), .Z(n3926) );
  XNOR U4245 ( .A(sreg[69]), .B(n3926), .Z(n3928) );
  NANDN U4246 ( .A(sreg[68]), .B(n3777), .Z(n3781) );
  NANDN U4247 ( .A(n3779), .B(n3778), .Z(n3780) );
  NAND U4248 ( .A(n3781), .B(n3780), .Z(n3927) );
  XNOR U4249 ( .A(n3928), .B(n3927), .Z(c[69]) );
  NANDN U4250 ( .A(n3783), .B(n3782), .Z(n3787) );
  NANDN U4251 ( .A(n3785), .B(n3784), .Z(n3786) );
  AND U4252 ( .A(n3787), .B(n3786), .Z(n3934) );
  NANDN U4253 ( .A(n3789), .B(n3788), .Z(n3793) );
  NANDN U4254 ( .A(n3791), .B(n3790), .Z(n3792) );
  AND U4255 ( .A(n3793), .B(n3792), .Z(n3932) );
  NANDN U4256 ( .A(n3795), .B(n3794), .Z(n3799) );
  NANDN U4257 ( .A(n3797), .B(n3796), .Z(n3798) );
  AND U4258 ( .A(n3799), .B(n3798), .Z(n3944) );
  NANDN U4259 ( .A(n3801), .B(n3800), .Z(n3805) );
  NAND U4260 ( .A(n3803), .B(n3802), .Z(n3804) );
  AND U4261 ( .A(n3805), .B(n3804), .Z(n3943) );
  XNOR U4262 ( .A(n3944), .B(n3943), .Z(n3946) );
  NANDN U4263 ( .A(n3807), .B(n3806), .Z(n3811) );
  NANDN U4264 ( .A(n3809), .B(n3808), .Z(n3810) );
  AND U4265 ( .A(n3811), .B(n3810), .Z(n4021) );
  NAND U4266 ( .A(n582), .B(n3812), .Z(n3814) );
  XOR U4267 ( .A(b[27]), .B(a[12]), .Z(n3967) );
  NAND U4268 ( .A(n9770), .B(n3967), .Z(n3813) );
  AND U4269 ( .A(n3814), .B(n3813), .Z(n4028) );
  NAND U4270 ( .A(n567), .B(n3815), .Z(n3817) );
  XOR U4271 ( .A(b[5]), .B(a[34]), .Z(n3970) );
  NAND U4272 ( .A(n7235), .B(n3970), .Z(n3816) );
  AND U4273 ( .A(n3817), .B(n3816), .Z(n4026) );
  NAND U4274 ( .A(n9046), .B(n3818), .Z(n3820) );
  XOR U4275 ( .A(b[19]), .B(a[20]), .Z(n3973) );
  NAND U4276 ( .A(n575), .B(n3973), .Z(n3819) );
  NAND U4277 ( .A(n3820), .B(n3819), .Z(n4025) );
  XNOR U4278 ( .A(n4026), .B(n4025), .Z(n4027) );
  XNOR U4279 ( .A(n4028), .B(n4027), .Z(n4019) );
  NAND U4280 ( .A(n9764), .B(n3821), .Z(n3823) );
  XOR U4281 ( .A(b[31]), .B(a[8]), .Z(n3976) );
  NAND U4282 ( .A(n584), .B(n3976), .Z(n3822) );
  AND U4283 ( .A(n3823), .B(n3822), .Z(n3988) );
  NAND U4284 ( .A(n568), .B(n3824), .Z(n3826) );
  XOR U4285 ( .A(b[3]), .B(a[36]), .Z(n3979) );
  NAND U4286 ( .A(n7245), .B(n3979), .Z(n3825) );
  AND U4287 ( .A(n3826), .B(n3825), .Z(n3986) );
  NAND U4288 ( .A(n576), .B(n3827), .Z(n3829) );
  XOR U4289 ( .A(b[17]), .B(a[22]), .Z(n3982) );
  NAND U4290 ( .A(n9141), .B(n3982), .Z(n3828) );
  NAND U4291 ( .A(n3829), .B(n3828), .Z(n3985) );
  XNOR U4292 ( .A(n3986), .B(n3985), .Z(n3987) );
  XOR U4293 ( .A(n3988), .B(n3987), .Z(n4020) );
  XOR U4294 ( .A(n4019), .B(n4020), .Z(n4022) );
  XOR U4295 ( .A(n4021), .B(n4022), .Z(n3956) );
  NANDN U4296 ( .A(n3831), .B(n3830), .Z(n3835) );
  NANDN U4297 ( .A(n3833), .B(n3832), .Z(n3834) );
  AND U4298 ( .A(n3835), .B(n3834), .Z(n4009) );
  NANDN U4299 ( .A(n3837), .B(n3836), .Z(n3841) );
  NANDN U4300 ( .A(n3839), .B(n3838), .Z(n3840) );
  NAND U4301 ( .A(n3841), .B(n3840), .Z(n4010) );
  XNOR U4302 ( .A(n4009), .B(n4010), .Z(n4011) );
  NANDN U4303 ( .A(n3843), .B(n3842), .Z(n3847) );
  NANDN U4304 ( .A(n3845), .B(n3844), .Z(n3846) );
  NAND U4305 ( .A(n3847), .B(n3846), .Z(n4012) );
  XNOR U4306 ( .A(n4011), .B(n4012), .Z(n3955) );
  XNOR U4307 ( .A(n3956), .B(n3955), .Z(n3958) );
  NANDN U4308 ( .A(n3849), .B(n3848), .Z(n3853) );
  NANDN U4309 ( .A(n3851), .B(n3850), .Z(n3852) );
  AND U4310 ( .A(n3853), .B(n3852), .Z(n3957) );
  XOR U4311 ( .A(n3958), .B(n3957), .Z(n4070) );
  NANDN U4312 ( .A(n3855), .B(n3854), .Z(n3859) );
  NANDN U4313 ( .A(n3857), .B(n3856), .Z(n3858) );
  AND U4314 ( .A(n3859), .B(n3858), .Z(n4067) );
  NANDN U4315 ( .A(n3861), .B(n3860), .Z(n3865) );
  NANDN U4316 ( .A(n3863), .B(n3862), .Z(n3864) );
  AND U4317 ( .A(n3865), .B(n3864), .Z(n3952) );
  NANDN U4318 ( .A(n3867), .B(n3866), .Z(n3871) );
  OR U4319 ( .A(n3869), .B(n3868), .Z(n3870) );
  AND U4320 ( .A(n3871), .B(n3870), .Z(n3950) );
  NANDN U4321 ( .A(n3873), .B(n3872), .Z(n3877) );
  NANDN U4322 ( .A(n3875), .B(n3874), .Z(n3876) );
  AND U4323 ( .A(n3877), .B(n3876), .Z(n4016) );
  NANDN U4324 ( .A(n3879), .B(n3878), .Z(n3883) );
  NANDN U4325 ( .A(n3881), .B(n3880), .Z(n3882) );
  NAND U4326 ( .A(n3883), .B(n3882), .Z(n4015) );
  XNOR U4327 ( .A(n4016), .B(n4015), .Z(n4018) );
  NAND U4328 ( .A(b[0]), .B(a[38]), .Z(n3884) );
  XNOR U4329 ( .A(b[1]), .B(n3884), .Z(n3886) );
  NANDN U4330 ( .A(b[0]), .B(a[37]), .Z(n3885) );
  NAND U4331 ( .A(n3886), .B(n3885), .Z(n3964) );
  NAND U4332 ( .A(n583), .B(n3887), .Z(n3889) );
  XOR U4333 ( .A(b[29]), .B(a[10]), .Z(n4037) );
  NAND U4334 ( .A(n581), .B(n4037), .Z(n3888) );
  AND U4335 ( .A(n3889), .B(n3888), .Z(n3962) );
  AND U4336 ( .A(b[31]), .B(a[6]), .Z(n3961) );
  XNOR U4337 ( .A(n3962), .B(n3961), .Z(n3963) );
  XNOR U4338 ( .A(n3964), .B(n3963), .Z(n4004) );
  NAND U4339 ( .A(n578), .B(n3890), .Z(n3892) );
  XOR U4340 ( .A(b[23]), .B(a[16]), .Z(n4043) );
  NAND U4341 ( .A(n9268), .B(n4043), .Z(n3891) );
  AND U4342 ( .A(n3892), .B(n3891), .Z(n4033) );
  NAND U4343 ( .A(n569), .B(n3893), .Z(n3895) );
  XOR U4344 ( .A(b[7]), .B(a[32]), .Z(n4046) );
  NAND U4345 ( .A(n7819), .B(n4046), .Z(n3894) );
  AND U4346 ( .A(n3895), .B(n3894), .Z(n4032) );
  NAND U4347 ( .A(n579), .B(n3896), .Z(n3898) );
  XOR U4348 ( .A(b[25]), .B(a[14]), .Z(n4049) );
  NAND U4349 ( .A(n9364), .B(n4049), .Z(n3897) );
  NAND U4350 ( .A(n3898), .B(n3897), .Z(n4031) );
  XOR U4351 ( .A(n4032), .B(n4031), .Z(n4034) );
  XOR U4352 ( .A(n4033), .B(n4034), .Z(n4003) );
  XOR U4353 ( .A(n4004), .B(n4003), .Z(n4006) );
  NAND U4354 ( .A(n572), .B(n3899), .Z(n3901) );
  XOR U4355 ( .A(b[13]), .B(a[26]), .Z(n4052) );
  NAND U4356 ( .A(n8585), .B(n4052), .Z(n3900) );
  AND U4357 ( .A(n3901), .B(n3900), .Z(n3998) );
  NAND U4358 ( .A(n571), .B(n3902), .Z(n3904) );
  XOR U4359 ( .A(b[11]), .B(a[28]), .Z(n4055) );
  NAND U4360 ( .A(n8135), .B(n4055), .Z(n3903) );
  NAND U4361 ( .A(n3904), .B(n3903), .Z(n3997) );
  XNOR U4362 ( .A(n3998), .B(n3997), .Z(n4000) );
  NAND U4363 ( .A(n573), .B(n3905), .Z(n3907) );
  XOR U4364 ( .A(b[15]), .B(a[24]), .Z(n4058) );
  NAND U4365 ( .A(n8694), .B(n4058), .Z(n3906) );
  AND U4366 ( .A(n3907), .B(n3906), .Z(n3994) );
  NAND U4367 ( .A(n577), .B(n3908), .Z(n3910) );
  XOR U4368 ( .A(b[21]), .B(a[18]), .Z(n4061) );
  NAND U4369 ( .A(n9216), .B(n4061), .Z(n3909) );
  AND U4370 ( .A(n3910), .B(n3909), .Z(n3992) );
  NAND U4371 ( .A(n570), .B(n3911), .Z(n3913) );
  XOR U4372 ( .A(b[9]), .B(a[30]), .Z(n4064) );
  NAND U4373 ( .A(n8037), .B(n4064), .Z(n3912) );
  NAND U4374 ( .A(n3913), .B(n3912), .Z(n3991) );
  XNOR U4375 ( .A(n3992), .B(n3991), .Z(n3993) );
  XNOR U4376 ( .A(n3994), .B(n3993), .Z(n3999) );
  XOR U4377 ( .A(n4000), .B(n3999), .Z(n4005) );
  XNOR U4378 ( .A(n4006), .B(n4005), .Z(n4017) );
  XNOR U4379 ( .A(n4018), .B(n4017), .Z(n3949) );
  XNOR U4380 ( .A(n3950), .B(n3949), .Z(n3951) );
  XOR U4381 ( .A(n3952), .B(n3951), .Z(n4068) );
  XNOR U4382 ( .A(n4067), .B(n4068), .Z(n4069) );
  XNOR U4383 ( .A(n4070), .B(n4069), .Z(n3945) );
  XOR U4384 ( .A(n3946), .B(n3945), .Z(n3938) );
  NANDN U4385 ( .A(n3915), .B(n3914), .Z(n3919) );
  NANDN U4386 ( .A(n3917), .B(n3916), .Z(n3918) );
  AND U4387 ( .A(n3919), .B(n3918), .Z(n3937) );
  XNOR U4388 ( .A(n3938), .B(n3937), .Z(n3939) );
  NANDN U4389 ( .A(n3921), .B(n3920), .Z(n3925) );
  NAND U4390 ( .A(n3923), .B(n3922), .Z(n3924) );
  NAND U4391 ( .A(n3925), .B(n3924), .Z(n3940) );
  XNOR U4392 ( .A(n3939), .B(n3940), .Z(n3931) );
  XNOR U4393 ( .A(n3932), .B(n3931), .Z(n3933) );
  XNOR U4394 ( .A(n3934), .B(n3933), .Z(n4073) );
  XNOR U4395 ( .A(sreg[70]), .B(n4073), .Z(n4075) );
  NANDN U4396 ( .A(sreg[69]), .B(n3926), .Z(n3930) );
  NAND U4397 ( .A(n3928), .B(n3927), .Z(n3929) );
  NAND U4398 ( .A(n3930), .B(n3929), .Z(n4074) );
  XNOR U4399 ( .A(n4075), .B(n4074), .Z(c[70]) );
  NANDN U4400 ( .A(n3932), .B(n3931), .Z(n3936) );
  NANDN U4401 ( .A(n3934), .B(n3933), .Z(n3935) );
  AND U4402 ( .A(n3936), .B(n3935), .Z(n4081) );
  NANDN U4403 ( .A(n3938), .B(n3937), .Z(n3942) );
  NANDN U4404 ( .A(n3940), .B(n3939), .Z(n3941) );
  AND U4405 ( .A(n3942), .B(n3941), .Z(n4079) );
  NANDN U4406 ( .A(n3944), .B(n3943), .Z(n3948) );
  NAND U4407 ( .A(n3946), .B(n3945), .Z(n3947) );
  AND U4408 ( .A(n3948), .B(n3947), .Z(n4086) );
  NANDN U4409 ( .A(n3950), .B(n3949), .Z(n3954) );
  NANDN U4410 ( .A(n3952), .B(n3951), .Z(n3953) );
  AND U4411 ( .A(n3954), .B(n3953), .Z(n4217) );
  NANDN U4412 ( .A(n3956), .B(n3955), .Z(n3960) );
  NAND U4413 ( .A(n3958), .B(n3957), .Z(n3959) );
  AND U4414 ( .A(n3960), .B(n3959), .Z(n4216) );
  XNOR U4415 ( .A(n4217), .B(n4216), .Z(n4219) );
  NANDN U4416 ( .A(n3962), .B(n3961), .Z(n3966) );
  NANDN U4417 ( .A(n3964), .B(n3963), .Z(n3965) );
  AND U4418 ( .A(n3966), .B(n3965), .Z(n4152) );
  NAND U4419 ( .A(n582), .B(n3967), .Z(n3969) );
  XOR U4420 ( .A(b[27]), .B(a[13]), .Z(n4096) );
  NAND U4421 ( .A(n9770), .B(n4096), .Z(n3968) );
  AND U4422 ( .A(n3969), .B(n3968), .Z(n4159) );
  NAND U4423 ( .A(n567), .B(n3970), .Z(n3972) );
  XOR U4424 ( .A(b[5]), .B(a[35]), .Z(n4099) );
  NAND U4425 ( .A(n7235), .B(n4099), .Z(n3971) );
  AND U4426 ( .A(n3972), .B(n3971), .Z(n4157) );
  NAND U4427 ( .A(n9046), .B(n3973), .Z(n3975) );
  XOR U4428 ( .A(b[19]), .B(a[21]), .Z(n4102) );
  NAND U4429 ( .A(n575), .B(n4102), .Z(n3974) );
  NAND U4430 ( .A(n3975), .B(n3974), .Z(n4156) );
  XNOR U4431 ( .A(n4157), .B(n4156), .Z(n4158) );
  XNOR U4432 ( .A(n4159), .B(n4158), .Z(n4150) );
  NAND U4433 ( .A(n9764), .B(n3976), .Z(n3978) );
  XOR U4434 ( .A(b[31]), .B(a[9]), .Z(n4105) );
  NAND U4435 ( .A(n584), .B(n4105), .Z(n3977) );
  AND U4436 ( .A(n3978), .B(n3977), .Z(n4117) );
  NAND U4437 ( .A(n568), .B(n3979), .Z(n3981) );
  XOR U4438 ( .A(a[37]), .B(b[3]), .Z(n4108) );
  NAND U4439 ( .A(n7245), .B(n4108), .Z(n3980) );
  AND U4440 ( .A(n3981), .B(n3980), .Z(n4115) );
  NAND U4441 ( .A(n576), .B(n3982), .Z(n3984) );
  XOR U4442 ( .A(b[17]), .B(a[23]), .Z(n4111) );
  NAND U4443 ( .A(n9141), .B(n4111), .Z(n3983) );
  NAND U4444 ( .A(n3984), .B(n3983), .Z(n4114) );
  XNOR U4445 ( .A(n4115), .B(n4114), .Z(n4116) );
  XOR U4446 ( .A(n4117), .B(n4116), .Z(n4151) );
  XOR U4447 ( .A(n4150), .B(n4151), .Z(n4153) );
  XOR U4448 ( .A(n4152), .B(n4153), .Z(n4199) );
  NANDN U4449 ( .A(n3986), .B(n3985), .Z(n3990) );
  NANDN U4450 ( .A(n3988), .B(n3987), .Z(n3989) );
  AND U4451 ( .A(n3990), .B(n3989), .Z(n4138) );
  NANDN U4452 ( .A(n3992), .B(n3991), .Z(n3996) );
  NANDN U4453 ( .A(n3994), .B(n3993), .Z(n3995) );
  NAND U4454 ( .A(n3996), .B(n3995), .Z(n4139) );
  XNOR U4455 ( .A(n4138), .B(n4139), .Z(n4140) );
  NANDN U4456 ( .A(n3998), .B(n3997), .Z(n4002) );
  NAND U4457 ( .A(n4000), .B(n3999), .Z(n4001) );
  NAND U4458 ( .A(n4002), .B(n4001), .Z(n4141) );
  XNOR U4459 ( .A(n4140), .B(n4141), .Z(n4198) );
  XNOR U4460 ( .A(n4199), .B(n4198), .Z(n4201) );
  NAND U4461 ( .A(n4004), .B(n4003), .Z(n4008) );
  NAND U4462 ( .A(n4006), .B(n4005), .Z(n4007) );
  AND U4463 ( .A(n4008), .B(n4007), .Z(n4200) );
  XOR U4464 ( .A(n4201), .B(n4200), .Z(n4213) );
  NANDN U4465 ( .A(n4010), .B(n4009), .Z(n4014) );
  NANDN U4466 ( .A(n4012), .B(n4011), .Z(n4013) );
  AND U4467 ( .A(n4014), .B(n4013), .Z(n4210) );
  NANDN U4468 ( .A(n4020), .B(n4019), .Z(n4024) );
  OR U4469 ( .A(n4022), .B(n4021), .Z(n4023) );
  AND U4470 ( .A(n4024), .B(n4023), .Z(n4205) );
  NANDN U4471 ( .A(n4026), .B(n4025), .Z(n4030) );
  NANDN U4472 ( .A(n4028), .B(n4027), .Z(n4029) );
  AND U4473 ( .A(n4030), .B(n4029), .Z(n4145) );
  NANDN U4474 ( .A(n4032), .B(n4031), .Z(n4036) );
  OR U4475 ( .A(n4034), .B(n4033), .Z(n4035) );
  NAND U4476 ( .A(n4036), .B(n4035), .Z(n4144) );
  XNOR U4477 ( .A(n4145), .B(n4144), .Z(n4146) );
  NAND U4478 ( .A(n583), .B(n4037), .Z(n4039) );
  XOR U4479 ( .A(b[29]), .B(a[11]), .Z(n4171) );
  NAND U4480 ( .A(n581), .B(n4171), .Z(n4038) );
  AND U4481 ( .A(n4039), .B(n4038), .Z(n4091) );
  AND U4482 ( .A(b[31]), .B(a[7]), .Z(n4090) );
  XNOR U4483 ( .A(n4091), .B(n4090), .Z(n4092) );
  NAND U4484 ( .A(b[0]), .B(a[39]), .Z(n4040) );
  XNOR U4485 ( .A(b[1]), .B(n4040), .Z(n4042) );
  NANDN U4486 ( .A(b[0]), .B(a[38]), .Z(n4041) );
  NAND U4487 ( .A(n4042), .B(n4041), .Z(n4093) );
  XNOR U4488 ( .A(n4092), .B(n4093), .Z(n4132) );
  NAND U4489 ( .A(n578), .B(n4043), .Z(n4045) );
  XOR U4490 ( .A(b[23]), .B(a[17]), .Z(n4174) );
  NAND U4491 ( .A(n9268), .B(n4174), .Z(n4044) );
  AND U4492 ( .A(n4045), .B(n4044), .Z(n4165) );
  NAND U4493 ( .A(n569), .B(n4046), .Z(n4048) );
  XOR U4494 ( .A(b[7]), .B(a[33]), .Z(n4177) );
  NAND U4495 ( .A(n7819), .B(n4177), .Z(n4047) );
  AND U4496 ( .A(n4048), .B(n4047), .Z(n4163) );
  NAND U4497 ( .A(n579), .B(n4049), .Z(n4051) );
  XOR U4498 ( .A(b[25]), .B(a[15]), .Z(n4180) );
  NAND U4499 ( .A(n9364), .B(n4180), .Z(n4050) );
  NAND U4500 ( .A(n4051), .B(n4050), .Z(n4162) );
  XNOR U4501 ( .A(n4163), .B(n4162), .Z(n4164) );
  XOR U4502 ( .A(n4165), .B(n4164), .Z(n4133) );
  XNOR U4503 ( .A(n4132), .B(n4133), .Z(n4134) );
  NAND U4504 ( .A(n572), .B(n4052), .Z(n4054) );
  XOR U4505 ( .A(b[13]), .B(a[27]), .Z(n4183) );
  NAND U4506 ( .A(n8585), .B(n4183), .Z(n4053) );
  AND U4507 ( .A(n4054), .B(n4053), .Z(n4127) );
  NAND U4508 ( .A(n571), .B(n4055), .Z(n4057) );
  XOR U4509 ( .A(b[11]), .B(a[29]), .Z(n4186) );
  NAND U4510 ( .A(n8135), .B(n4186), .Z(n4056) );
  NAND U4511 ( .A(n4057), .B(n4056), .Z(n4126) );
  XNOR U4512 ( .A(n4127), .B(n4126), .Z(n4128) );
  NAND U4513 ( .A(n573), .B(n4058), .Z(n4060) );
  XOR U4514 ( .A(b[15]), .B(a[25]), .Z(n4189) );
  NAND U4515 ( .A(n8694), .B(n4189), .Z(n4059) );
  AND U4516 ( .A(n4060), .B(n4059), .Z(n4123) );
  NAND U4517 ( .A(n577), .B(n4061), .Z(n4063) );
  XOR U4518 ( .A(b[21]), .B(a[19]), .Z(n4192) );
  NAND U4519 ( .A(n9216), .B(n4192), .Z(n4062) );
  AND U4520 ( .A(n4063), .B(n4062), .Z(n4121) );
  NAND U4521 ( .A(n570), .B(n4064), .Z(n4066) );
  XOR U4522 ( .A(b[9]), .B(a[31]), .Z(n4195) );
  NAND U4523 ( .A(n8037), .B(n4195), .Z(n4065) );
  NAND U4524 ( .A(n4066), .B(n4065), .Z(n4120) );
  XNOR U4525 ( .A(n4121), .B(n4120), .Z(n4122) );
  XOR U4526 ( .A(n4123), .B(n4122), .Z(n4129) );
  XOR U4527 ( .A(n4128), .B(n4129), .Z(n4135) );
  XOR U4528 ( .A(n4134), .B(n4135), .Z(n4147) );
  XNOR U4529 ( .A(n4146), .B(n4147), .Z(n4204) );
  XNOR U4530 ( .A(n4205), .B(n4204), .Z(n4206) );
  XOR U4531 ( .A(n4207), .B(n4206), .Z(n4211) );
  XNOR U4532 ( .A(n4210), .B(n4211), .Z(n4212) );
  XNOR U4533 ( .A(n4213), .B(n4212), .Z(n4218) );
  XOR U4534 ( .A(n4219), .B(n4218), .Z(n4085) );
  NANDN U4535 ( .A(n4068), .B(n4067), .Z(n4072) );
  NANDN U4536 ( .A(n4070), .B(n4069), .Z(n4071) );
  AND U4537 ( .A(n4072), .B(n4071), .Z(n4084) );
  XOR U4538 ( .A(n4085), .B(n4084), .Z(n4087) );
  XNOR U4539 ( .A(n4086), .B(n4087), .Z(n4078) );
  XNOR U4540 ( .A(n4079), .B(n4078), .Z(n4080) );
  XNOR U4541 ( .A(n4081), .B(n4080), .Z(n4222) );
  XNOR U4542 ( .A(sreg[71]), .B(n4222), .Z(n4224) );
  NANDN U4543 ( .A(sreg[70]), .B(n4073), .Z(n4077) );
  NAND U4544 ( .A(n4075), .B(n4074), .Z(n4076) );
  NAND U4545 ( .A(n4077), .B(n4076), .Z(n4223) );
  XNOR U4546 ( .A(n4224), .B(n4223), .Z(c[71]) );
  NANDN U4547 ( .A(n4079), .B(n4078), .Z(n4083) );
  NANDN U4548 ( .A(n4081), .B(n4080), .Z(n4082) );
  AND U4549 ( .A(n4083), .B(n4082), .Z(n4230) );
  NANDN U4550 ( .A(n4085), .B(n4084), .Z(n4089) );
  NANDN U4551 ( .A(n4087), .B(n4086), .Z(n4088) );
  AND U4552 ( .A(n4089), .B(n4088), .Z(n4228) );
  NANDN U4553 ( .A(n4091), .B(n4090), .Z(n4095) );
  NANDN U4554 ( .A(n4093), .B(n4092), .Z(n4094) );
  AND U4555 ( .A(n4095), .B(n4094), .Z(n4319) );
  NAND U4556 ( .A(n582), .B(n4096), .Z(n4098) );
  XOR U4557 ( .A(b[27]), .B(a[14]), .Z(n4263) );
  NAND U4558 ( .A(n9770), .B(n4263), .Z(n4097) );
  AND U4559 ( .A(n4098), .B(n4097), .Z(n4326) );
  NAND U4560 ( .A(n567), .B(n4099), .Z(n4101) );
  XOR U4561 ( .A(b[5]), .B(a[36]), .Z(n4266) );
  NAND U4562 ( .A(n7235), .B(n4266), .Z(n4100) );
  AND U4563 ( .A(n4101), .B(n4100), .Z(n4324) );
  NAND U4564 ( .A(n9046), .B(n4102), .Z(n4104) );
  XOR U4565 ( .A(b[19]), .B(a[22]), .Z(n4269) );
  NAND U4566 ( .A(n575), .B(n4269), .Z(n4103) );
  NAND U4567 ( .A(n4104), .B(n4103), .Z(n4323) );
  XNOR U4568 ( .A(n4324), .B(n4323), .Z(n4325) );
  XNOR U4569 ( .A(n4326), .B(n4325), .Z(n4317) );
  NAND U4570 ( .A(n9764), .B(n4105), .Z(n4107) );
  XOR U4571 ( .A(b[31]), .B(a[10]), .Z(n4272) );
  NAND U4572 ( .A(n584), .B(n4272), .Z(n4106) );
  AND U4573 ( .A(n4107), .B(n4106), .Z(n4284) );
  NAND U4574 ( .A(n568), .B(n4108), .Z(n4110) );
  XOR U4575 ( .A(a[38]), .B(b[3]), .Z(n4275) );
  NAND U4576 ( .A(n7245), .B(n4275), .Z(n4109) );
  AND U4577 ( .A(n4110), .B(n4109), .Z(n4282) );
  NAND U4578 ( .A(n576), .B(n4111), .Z(n4113) );
  XOR U4579 ( .A(b[17]), .B(a[24]), .Z(n4278) );
  NAND U4580 ( .A(n9141), .B(n4278), .Z(n4112) );
  NAND U4581 ( .A(n4113), .B(n4112), .Z(n4281) );
  XNOR U4582 ( .A(n4282), .B(n4281), .Z(n4283) );
  XOR U4583 ( .A(n4284), .B(n4283), .Z(n4318) );
  XOR U4584 ( .A(n4317), .B(n4318), .Z(n4320) );
  XOR U4585 ( .A(n4319), .B(n4320), .Z(n4252) );
  NANDN U4586 ( .A(n4115), .B(n4114), .Z(n4119) );
  NANDN U4587 ( .A(n4117), .B(n4116), .Z(n4118) );
  AND U4588 ( .A(n4119), .B(n4118), .Z(n4305) );
  NANDN U4589 ( .A(n4121), .B(n4120), .Z(n4125) );
  NANDN U4590 ( .A(n4123), .B(n4122), .Z(n4124) );
  NAND U4591 ( .A(n4125), .B(n4124), .Z(n4306) );
  XNOR U4592 ( .A(n4305), .B(n4306), .Z(n4307) );
  NANDN U4593 ( .A(n4127), .B(n4126), .Z(n4131) );
  NANDN U4594 ( .A(n4129), .B(n4128), .Z(n4130) );
  NAND U4595 ( .A(n4131), .B(n4130), .Z(n4308) );
  XNOR U4596 ( .A(n4307), .B(n4308), .Z(n4251) );
  XNOR U4597 ( .A(n4252), .B(n4251), .Z(n4254) );
  NANDN U4598 ( .A(n4133), .B(n4132), .Z(n4137) );
  NANDN U4599 ( .A(n4135), .B(n4134), .Z(n4136) );
  AND U4600 ( .A(n4137), .B(n4136), .Z(n4253) );
  XOR U4601 ( .A(n4254), .B(n4253), .Z(n4367) );
  NANDN U4602 ( .A(n4139), .B(n4138), .Z(n4143) );
  NANDN U4603 ( .A(n4141), .B(n4140), .Z(n4142) );
  AND U4604 ( .A(n4143), .B(n4142), .Z(n4365) );
  NANDN U4605 ( .A(n4145), .B(n4144), .Z(n4149) );
  NANDN U4606 ( .A(n4147), .B(n4146), .Z(n4148) );
  AND U4607 ( .A(n4149), .B(n4148), .Z(n4248) );
  NANDN U4608 ( .A(n4151), .B(n4150), .Z(n4155) );
  OR U4609 ( .A(n4153), .B(n4152), .Z(n4154) );
  AND U4610 ( .A(n4155), .B(n4154), .Z(n4246) );
  NANDN U4611 ( .A(n4157), .B(n4156), .Z(n4161) );
  NANDN U4612 ( .A(n4159), .B(n4158), .Z(n4160) );
  AND U4613 ( .A(n4161), .B(n4160), .Z(n4312) );
  NANDN U4614 ( .A(n4163), .B(n4162), .Z(n4167) );
  NANDN U4615 ( .A(n4165), .B(n4164), .Z(n4166) );
  NAND U4616 ( .A(n4167), .B(n4166), .Z(n4311) );
  XNOR U4617 ( .A(n4312), .B(n4311), .Z(n4313) );
  NAND U4618 ( .A(b[0]), .B(a[40]), .Z(n4168) );
  XNOR U4619 ( .A(b[1]), .B(n4168), .Z(n4170) );
  NANDN U4620 ( .A(b[0]), .B(a[39]), .Z(n4169) );
  NAND U4621 ( .A(n4170), .B(n4169), .Z(n4260) );
  NAND U4622 ( .A(n583), .B(n4171), .Z(n4173) );
  XOR U4623 ( .A(b[29]), .B(a[12]), .Z(n4338) );
  NAND U4624 ( .A(n581), .B(n4338), .Z(n4172) );
  AND U4625 ( .A(n4173), .B(n4172), .Z(n4258) );
  AND U4626 ( .A(b[31]), .B(a[8]), .Z(n4257) );
  XNOR U4627 ( .A(n4258), .B(n4257), .Z(n4259) );
  XNOR U4628 ( .A(n4260), .B(n4259), .Z(n4299) );
  NAND U4629 ( .A(n578), .B(n4174), .Z(n4176) );
  XOR U4630 ( .A(b[23]), .B(a[18]), .Z(n4341) );
  NAND U4631 ( .A(n9268), .B(n4341), .Z(n4175) );
  AND U4632 ( .A(n4176), .B(n4175), .Z(n4332) );
  NAND U4633 ( .A(n569), .B(n4177), .Z(n4179) );
  XOR U4634 ( .A(b[7]), .B(a[34]), .Z(n4344) );
  NAND U4635 ( .A(n7819), .B(n4344), .Z(n4178) );
  AND U4636 ( .A(n4179), .B(n4178), .Z(n4330) );
  NAND U4637 ( .A(n579), .B(n4180), .Z(n4182) );
  XOR U4638 ( .A(b[25]), .B(a[16]), .Z(n4347) );
  NAND U4639 ( .A(n9364), .B(n4347), .Z(n4181) );
  NAND U4640 ( .A(n4182), .B(n4181), .Z(n4329) );
  XNOR U4641 ( .A(n4330), .B(n4329), .Z(n4331) );
  XOR U4642 ( .A(n4332), .B(n4331), .Z(n4300) );
  XNOR U4643 ( .A(n4299), .B(n4300), .Z(n4301) );
  NAND U4644 ( .A(n572), .B(n4183), .Z(n4185) );
  XOR U4645 ( .A(b[13]), .B(a[28]), .Z(n4350) );
  NAND U4646 ( .A(n8585), .B(n4350), .Z(n4184) );
  AND U4647 ( .A(n4185), .B(n4184), .Z(n4294) );
  NAND U4648 ( .A(n571), .B(n4186), .Z(n4188) );
  XOR U4649 ( .A(b[11]), .B(a[30]), .Z(n4353) );
  NAND U4650 ( .A(n8135), .B(n4353), .Z(n4187) );
  NAND U4651 ( .A(n4188), .B(n4187), .Z(n4293) );
  XNOR U4652 ( .A(n4294), .B(n4293), .Z(n4295) );
  NAND U4653 ( .A(n573), .B(n4189), .Z(n4191) );
  XOR U4654 ( .A(b[15]), .B(a[26]), .Z(n4356) );
  NAND U4655 ( .A(n8694), .B(n4356), .Z(n4190) );
  AND U4656 ( .A(n4191), .B(n4190), .Z(n4290) );
  NAND U4657 ( .A(n577), .B(n4192), .Z(n4194) );
  XOR U4658 ( .A(b[21]), .B(a[20]), .Z(n4359) );
  NAND U4659 ( .A(n9216), .B(n4359), .Z(n4193) );
  AND U4660 ( .A(n4194), .B(n4193), .Z(n4288) );
  NAND U4661 ( .A(n570), .B(n4195), .Z(n4197) );
  XOR U4662 ( .A(b[9]), .B(a[32]), .Z(n4362) );
  NAND U4663 ( .A(n8037), .B(n4362), .Z(n4196) );
  NAND U4664 ( .A(n4197), .B(n4196), .Z(n4287) );
  XNOR U4665 ( .A(n4288), .B(n4287), .Z(n4289) );
  XOR U4666 ( .A(n4290), .B(n4289), .Z(n4296) );
  XOR U4667 ( .A(n4295), .B(n4296), .Z(n4302) );
  XOR U4668 ( .A(n4301), .B(n4302), .Z(n4314) );
  XNOR U4669 ( .A(n4313), .B(n4314), .Z(n4245) );
  XNOR U4670 ( .A(n4246), .B(n4245), .Z(n4247) );
  XOR U4671 ( .A(n4248), .B(n4247), .Z(n4366) );
  XOR U4672 ( .A(n4365), .B(n4366), .Z(n4368) );
  XOR U4673 ( .A(n4367), .B(n4368), .Z(n4242) );
  NANDN U4674 ( .A(n4199), .B(n4198), .Z(n4203) );
  NAND U4675 ( .A(n4201), .B(n4200), .Z(n4202) );
  AND U4676 ( .A(n4203), .B(n4202), .Z(n4240) );
  NANDN U4677 ( .A(n4205), .B(n4204), .Z(n4209) );
  NANDN U4678 ( .A(n4207), .B(n4206), .Z(n4208) );
  AND U4679 ( .A(n4209), .B(n4208), .Z(n4239) );
  XNOR U4680 ( .A(n4240), .B(n4239), .Z(n4241) );
  XNOR U4681 ( .A(n4242), .B(n4241), .Z(n4233) );
  NANDN U4682 ( .A(n4211), .B(n4210), .Z(n4215) );
  NANDN U4683 ( .A(n4213), .B(n4212), .Z(n4214) );
  NAND U4684 ( .A(n4215), .B(n4214), .Z(n4234) );
  XNOR U4685 ( .A(n4233), .B(n4234), .Z(n4235) );
  NANDN U4686 ( .A(n4217), .B(n4216), .Z(n4221) );
  NAND U4687 ( .A(n4219), .B(n4218), .Z(n4220) );
  NAND U4688 ( .A(n4221), .B(n4220), .Z(n4236) );
  XNOR U4689 ( .A(n4235), .B(n4236), .Z(n4227) );
  XNOR U4690 ( .A(n4228), .B(n4227), .Z(n4229) );
  XNOR U4691 ( .A(n4230), .B(n4229), .Z(n4371) );
  XNOR U4692 ( .A(sreg[72]), .B(n4371), .Z(n4373) );
  NANDN U4693 ( .A(sreg[71]), .B(n4222), .Z(n4226) );
  NAND U4694 ( .A(n4224), .B(n4223), .Z(n4225) );
  NAND U4695 ( .A(n4226), .B(n4225), .Z(n4372) );
  XNOR U4696 ( .A(n4373), .B(n4372), .Z(c[72]) );
  NANDN U4697 ( .A(n4228), .B(n4227), .Z(n4232) );
  NANDN U4698 ( .A(n4230), .B(n4229), .Z(n4231) );
  AND U4699 ( .A(n4232), .B(n4231), .Z(n4379) );
  NANDN U4700 ( .A(n4234), .B(n4233), .Z(n4238) );
  NANDN U4701 ( .A(n4236), .B(n4235), .Z(n4237) );
  AND U4702 ( .A(n4238), .B(n4237), .Z(n4377) );
  NANDN U4703 ( .A(n4240), .B(n4239), .Z(n4244) );
  NANDN U4704 ( .A(n4242), .B(n4241), .Z(n4243) );
  AND U4705 ( .A(n4244), .B(n4243), .Z(n4385) );
  NANDN U4706 ( .A(n4246), .B(n4245), .Z(n4250) );
  NANDN U4707 ( .A(n4248), .B(n4247), .Z(n4249) );
  AND U4708 ( .A(n4250), .B(n4249), .Z(n4389) );
  NANDN U4709 ( .A(n4252), .B(n4251), .Z(n4256) );
  NAND U4710 ( .A(n4254), .B(n4253), .Z(n4255) );
  AND U4711 ( .A(n4256), .B(n4255), .Z(n4388) );
  XNOR U4712 ( .A(n4389), .B(n4388), .Z(n4391) );
  NANDN U4713 ( .A(n4258), .B(n4257), .Z(n4262) );
  NANDN U4714 ( .A(n4260), .B(n4259), .Z(n4261) );
  AND U4715 ( .A(n4262), .B(n4261), .Z(n4468) );
  NAND U4716 ( .A(n582), .B(n4263), .Z(n4265) );
  XOR U4717 ( .A(b[27]), .B(a[15]), .Z(n4412) );
  NAND U4718 ( .A(n9770), .B(n4412), .Z(n4264) );
  AND U4719 ( .A(n4265), .B(n4264), .Z(n4475) );
  NAND U4720 ( .A(n567), .B(n4266), .Z(n4268) );
  XOR U4721 ( .A(b[5]), .B(a[37]), .Z(n4415) );
  NAND U4722 ( .A(n7235), .B(n4415), .Z(n4267) );
  AND U4723 ( .A(n4268), .B(n4267), .Z(n4473) );
  NAND U4724 ( .A(n9046), .B(n4269), .Z(n4271) );
  XOR U4725 ( .A(b[19]), .B(a[23]), .Z(n4418) );
  NAND U4726 ( .A(n575), .B(n4418), .Z(n4270) );
  NAND U4727 ( .A(n4271), .B(n4270), .Z(n4472) );
  XNOR U4728 ( .A(n4473), .B(n4472), .Z(n4474) );
  XNOR U4729 ( .A(n4475), .B(n4474), .Z(n4466) );
  NAND U4730 ( .A(n9764), .B(n4272), .Z(n4274) );
  XOR U4731 ( .A(b[31]), .B(a[11]), .Z(n4421) );
  NAND U4732 ( .A(n584), .B(n4421), .Z(n4273) );
  AND U4733 ( .A(n4274), .B(n4273), .Z(n4433) );
  NAND U4734 ( .A(n568), .B(n4275), .Z(n4277) );
  XOR U4735 ( .A(a[39]), .B(b[3]), .Z(n4424) );
  NAND U4736 ( .A(n7245), .B(n4424), .Z(n4276) );
  AND U4737 ( .A(n4277), .B(n4276), .Z(n4431) );
  NAND U4738 ( .A(n576), .B(n4278), .Z(n4280) );
  XOR U4739 ( .A(b[17]), .B(a[25]), .Z(n4427) );
  NAND U4740 ( .A(n9141), .B(n4427), .Z(n4279) );
  NAND U4741 ( .A(n4280), .B(n4279), .Z(n4430) );
  XNOR U4742 ( .A(n4431), .B(n4430), .Z(n4432) );
  XOR U4743 ( .A(n4433), .B(n4432), .Z(n4467) );
  XOR U4744 ( .A(n4466), .B(n4467), .Z(n4469) );
  XOR U4745 ( .A(n4468), .B(n4469), .Z(n4401) );
  NANDN U4746 ( .A(n4282), .B(n4281), .Z(n4286) );
  NANDN U4747 ( .A(n4284), .B(n4283), .Z(n4285) );
  AND U4748 ( .A(n4286), .B(n4285), .Z(n4454) );
  NANDN U4749 ( .A(n4288), .B(n4287), .Z(n4292) );
  NANDN U4750 ( .A(n4290), .B(n4289), .Z(n4291) );
  NAND U4751 ( .A(n4292), .B(n4291), .Z(n4455) );
  XNOR U4752 ( .A(n4454), .B(n4455), .Z(n4456) );
  NANDN U4753 ( .A(n4294), .B(n4293), .Z(n4298) );
  NANDN U4754 ( .A(n4296), .B(n4295), .Z(n4297) );
  NAND U4755 ( .A(n4298), .B(n4297), .Z(n4457) );
  XNOR U4756 ( .A(n4456), .B(n4457), .Z(n4400) );
  XNOR U4757 ( .A(n4401), .B(n4400), .Z(n4403) );
  NANDN U4758 ( .A(n4300), .B(n4299), .Z(n4304) );
  NANDN U4759 ( .A(n4302), .B(n4301), .Z(n4303) );
  AND U4760 ( .A(n4304), .B(n4303), .Z(n4402) );
  XOR U4761 ( .A(n4403), .B(n4402), .Z(n4517) );
  NANDN U4762 ( .A(n4306), .B(n4305), .Z(n4310) );
  NANDN U4763 ( .A(n4308), .B(n4307), .Z(n4309) );
  AND U4764 ( .A(n4310), .B(n4309), .Z(n4514) );
  NANDN U4765 ( .A(n4312), .B(n4311), .Z(n4316) );
  NANDN U4766 ( .A(n4314), .B(n4313), .Z(n4315) );
  AND U4767 ( .A(n4316), .B(n4315), .Z(n4397) );
  NANDN U4768 ( .A(n4318), .B(n4317), .Z(n4322) );
  OR U4769 ( .A(n4320), .B(n4319), .Z(n4321) );
  AND U4770 ( .A(n4322), .B(n4321), .Z(n4395) );
  NANDN U4771 ( .A(n4324), .B(n4323), .Z(n4328) );
  NANDN U4772 ( .A(n4326), .B(n4325), .Z(n4327) );
  AND U4773 ( .A(n4328), .B(n4327), .Z(n4461) );
  NANDN U4774 ( .A(n4330), .B(n4329), .Z(n4334) );
  NANDN U4775 ( .A(n4332), .B(n4331), .Z(n4333) );
  NAND U4776 ( .A(n4334), .B(n4333), .Z(n4460) );
  XNOR U4777 ( .A(n4461), .B(n4460), .Z(n4462) );
  NAND U4778 ( .A(b[0]), .B(a[41]), .Z(n4335) );
  XNOR U4779 ( .A(b[1]), .B(n4335), .Z(n4337) );
  NANDN U4780 ( .A(b[0]), .B(a[40]), .Z(n4336) );
  NAND U4781 ( .A(n4337), .B(n4336), .Z(n4409) );
  NAND U4782 ( .A(n583), .B(n4338), .Z(n4340) );
  XOR U4783 ( .A(b[29]), .B(a[13]), .Z(n4487) );
  NAND U4784 ( .A(n581), .B(n4487), .Z(n4339) );
  AND U4785 ( .A(n4340), .B(n4339), .Z(n4407) );
  AND U4786 ( .A(b[31]), .B(a[9]), .Z(n4406) );
  XNOR U4787 ( .A(n4407), .B(n4406), .Z(n4408) );
  XNOR U4788 ( .A(n4409), .B(n4408), .Z(n4448) );
  NAND U4789 ( .A(n578), .B(n4341), .Z(n4343) );
  XOR U4790 ( .A(b[23]), .B(a[19]), .Z(n4490) );
  NAND U4791 ( .A(n9268), .B(n4490), .Z(n4342) );
  AND U4792 ( .A(n4343), .B(n4342), .Z(n4481) );
  NAND U4793 ( .A(n569), .B(n4344), .Z(n4346) );
  XOR U4794 ( .A(b[7]), .B(a[35]), .Z(n4493) );
  NAND U4795 ( .A(n7819), .B(n4493), .Z(n4345) );
  AND U4796 ( .A(n4346), .B(n4345), .Z(n4479) );
  NAND U4797 ( .A(n579), .B(n4347), .Z(n4349) );
  XOR U4798 ( .A(b[25]), .B(a[17]), .Z(n4496) );
  NAND U4799 ( .A(n9364), .B(n4496), .Z(n4348) );
  NAND U4800 ( .A(n4349), .B(n4348), .Z(n4478) );
  XNOR U4801 ( .A(n4479), .B(n4478), .Z(n4480) );
  XOR U4802 ( .A(n4481), .B(n4480), .Z(n4449) );
  XNOR U4803 ( .A(n4448), .B(n4449), .Z(n4450) );
  NAND U4804 ( .A(n572), .B(n4350), .Z(n4352) );
  XOR U4805 ( .A(b[13]), .B(a[29]), .Z(n4499) );
  NAND U4806 ( .A(n8585), .B(n4499), .Z(n4351) );
  AND U4807 ( .A(n4352), .B(n4351), .Z(n4443) );
  NAND U4808 ( .A(n571), .B(n4353), .Z(n4355) );
  XOR U4809 ( .A(b[11]), .B(a[31]), .Z(n4502) );
  NAND U4810 ( .A(n8135), .B(n4502), .Z(n4354) );
  NAND U4811 ( .A(n4355), .B(n4354), .Z(n4442) );
  XNOR U4812 ( .A(n4443), .B(n4442), .Z(n4444) );
  NAND U4813 ( .A(n573), .B(n4356), .Z(n4358) );
  XOR U4814 ( .A(b[15]), .B(a[27]), .Z(n4505) );
  NAND U4815 ( .A(n8694), .B(n4505), .Z(n4357) );
  AND U4816 ( .A(n4358), .B(n4357), .Z(n4439) );
  NAND U4817 ( .A(n577), .B(n4359), .Z(n4361) );
  XOR U4818 ( .A(b[21]), .B(a[21]), .Z(n4508) );
  NAND U4819 ( .A(n9216), .B(n4508), .Z(n4360) );
  AND U4820 ( .A(n4361), .B(n4360), .Z(n4437) );
  NAND U4821 ( .A(n570), .B(n4362), .Z(n4364) );
  XOR U4822 ( .A(b[9]), .B(a[33]), .Z(n4511) );
  NAND U4823 ( .A(n8037), .B(n4511), .Z(n4363) );
  NAND U4824 ( .A(n4364), .B(n4363), .Z(n4436) );
  XNOR U4825 ( .A(n4437), .B(n4436), .Z(n4438) );
  XOR U4826 ( .A(n4439), .B(n4438), .Z(n4445) );
  XOR U4827 ( .A(n4444), .B(n4445), .Z(n4451) );
  XOR U4828 ( .A(n4450), .B(n4451), .Z(n4463) );
  XNOR U4829 ( .A(n4462), .B(n4463), .Z(n4394) );
  XNOR U4830 ( .A(n4395), .B(n4394), .Z(n4396) );
  XOR U4831 ( .A(n4397), .B(n4396), .Z(n4515) );
  XNOR U4832 ( .A(n4514), .B(n4515), .Z(n4516) );
  XNOR U4833 ( .A(n4517), .B(n4516), .Z(n4390) );
  XOR U4834 ( .A(n4391), .B(n4390), .Z(n4383) );
  NANDN U4835 ( .A(n4366), .B(n4365), .Z(n4370) );
  OR U4836 ( .A(n4368), .B(n4367), .Z(n4369) );
  AND U4837 ( .A(n4370), .B(n4369), .Z(n4382) );
  XNOR U4838 ( .A(n4383), .B(n4382), .Z(n4384) );
  XNOR U4839 ( .A(n4385), .B(n4384), .Z(n4376) );
  XNOR U4840 ( .A(n4377), .B(n4376), .Z(n4378) );
  XNOR U4841 ( .A(n4379), .B(n4378), .Z(n4520) );
  XNOR U4842 ( .A(sreg[73]), .B(n4520), .Z(n4522) );
  NANDN U4843 ( .A(sreg[72]), .B(n4371), .Z(n4375) );
  NAND U4844 ( .A(n4373), .B(n4372), .Z(n4374) );
  NAND U4845 ( .A(n4375), .B(n4374), .Z(n4521) );
  XNOR U4846 ( .A(n4522), .B(n4521), .Z(c[73]) );
  NANDN U4847 ( .A(n4377), .B(n4376), .Z(n4381) );
  NANDN U4848 ( .A(n4379), .B(n4378), .Z(n4380) );
  AND U4849 ( .A(n4381), .B(n4380), .Z(n4528) );
  NANDN U4850 ( .A(n4383), .B(n4382), .Z(n4387) );
  NANDN U4851 ( .A(n4385), .B(n4384), .Z(n4386) );
  AND U4852 ( .A(n4387), .B(n4386), .Z(n4526) );
  NANDN U4853 ( .A(n4389), .B(n4388), .Z(n4393) );
  NAND U4854 ( .A(n4391), .B(n4390), .Z(n4392) );
  AND U4855 ( .A(n4393), .B(n4392), .Z(n4533) );
  NANDN U4856 ( .A(n4395), .B(n4394), .Z(n4399) );
  NANDN U4857 ( .A(n4397), .B(n4396), .Z(n4398) );
  AND U4858 ( .A(n4399), .B(n4398), .Z(n4538) );
  NANDN U4859 ( .A(n4401), .B(n4400), .Z(n4405) );
  NAND U4860 ( .A(n4403), .B(n4402), .Z(n4404) );
  AND U4861 ( .A(n4405), .B(n4404), .Z(n4537) );
  XNOR U4862 ( .A(n4538), .B(n4537), .Z(n4540) );
  NANDN U4863 ( .A(n4407), .B(n4406), .Z(n4411) );
  NANDN U4864 ( .A(n4409), .B(n4408), .Z(n4410) );
  AND U4865 ( .A(n4411), .B(n4410), .Z(n4617) );
  NAND U4866 ( .A(n582), .B(n4412), .Z(n4414) );
  XOR U4867 ( .A(b[27]), .B(a[16]), .Z(n4561) );
  NAND U4868 ( .A(n9770), .B(n4561), .Z(n4413) );
  AND U4869 ( .A(n4414), .B(n4413), .Z(n4624) );
  NAND U4870 ( .A(n567), .B(n4415), .Z(n4417) );
  XOR U4871 ( .A(b[5]), .B(a[38]), .Z(n4564) );
  NAND U4872 ( .A(n7235), .B(n4564), .Z(n4416) );
  AND U4873 ( .A(n4417), .B(n4416), .Z(n4622) );
  NAND U4874 ( .A(n9046), .B(n4418), .Z(n4420) );
  XOR U4875 ( .A(b[19]), .B(a[24]), .Z(n4567) );
  NAND U4876 ( .A(n575), .B(n4567), .Z(n4419) );
  NAND U4877 ( .A(n4420), .B(n4419), .Z(n4621) );
  XNOR U4878 ( .A(n4622), .B(n4621), .Z(n4623) );
  XNOR U4879 ( .A(n4624), .B(n4623), .Z(n4615) );
  NAND U4880 ( .A(n9764), .B(n4421), .Z(n4423) );
  XOR U4881 ( .A(b[31]), .B(a[12]), .Z(n4570) );
  NAND U4882 ( .A(n584), .B(n4570), .Z(n4422) );
  AND U4883 ( .A(n4423), .B(n4422), .Z(n4582) );
  NAND U4884 ( .A(n568), .B(n4424), .Z(n4426) );
  XOR U4885 ( .A(a[40]), .B(b[3]), .Z(n4573) );
  NAND U4886 ( .A(n7245), .B(n4573), .Z(n4425) );
  AND U4887 ( .A(n4426), .B(n4425), .Z(n4580) );
  NAND U4888 ( .A(n576), .B(n4427), .Z(n4429) );
  XOR U4889 ( .A(b[17]), .B(a[26]), .Z(n4576) );
  NAND U4890 ( .A(n9141), .B(n4576), .Z(n4428) );
  NAND U4891 ( .A(n4429), .B(n4428), .Z(n4579) );
  XNOR U4892 ( .A(n4580), .B(n4579), .Z(n4581) );
  XOR U4893 ( .A(n4582), .B(n4581), .Z(n4616) );
  XOR U4894 ( .A(n4615), .B(n4616), .Z(n4618) );
  XOR U4895 ( .A(n4617), .B(n4618), .Z(n4550) );
  NANDN U4896 ( .A(n4431), .B(n4430), .Z(n4435) );
  NANDN U4897 ( .A(n4433), .B(n4432), .Z(n4434) );
  AND U4898 ( .A(n4435), .B(n4434), .Z(n4603) );
  NANDN U4899 ( .A(n4437), .B(n4436), .Z(n4441) );
  NANDN U4900 ( .A(n4439), .B(n4438), .Z(n4440) );
  NAND U4901 ( .A(n4441), .B(n4440), .Z(n4604) );
  XNOR U4902 ( .A(n4603), .B(n4604), .Z(n4605) );
  NANDN U4903 ( .A(n4443), .B(n4442), .Z(n4447) );
  NANDN U4904 ( .A(n4445), .B(n4444), .Z(n4446) );
  NAND U4905 ( .A(n4447), .B(n4446), .Z(n4606) );
  XNOR U4906 ( .A(n4605), .B(n4606), .Z(n4549) );
  XNOR U4907 ( .A(n4550), .B(n4549), .Z(n4552) );
  NANDN U4908 ( .A(n4449), .B(n4448), .Z(n4453) );
  NANDN U4909 ( .A(n4451), .B(n4450), .Z(n4452) );
  AND U4910 ( .A(n4453), .B(n4452), .Z(n4551) );
  XOR U4911 ( .A(n4552), .B(n4551), .Z(n4666) );
  NANDN U4912 ( .A(n4455), .B(n4454), .Z(n4459) );
  NANDN U4913 ( .A(n4457), .B(n4456), .Z(n4458) );
  AND U4914 ( .A(n4459), .B(n4458), .Z(n4663) );
  NANDN U4915 ( .A(n4461), .B(n4460), .Z(n4465) );
  NANDN U4916 ( .A(n4463), .B(n4462), .Z(n4464) );
  AND U4917 ( .A(n4465), .B(n4464), .Z(n4546) );
  NANDN U4918 ( .A(n4467), .B(n4466), .Z(n4471) );
  OR U4919 ( .A(n4469), .B(n4468), .Z(n4470) );
  AND U4920 ( .A(n4471), .B(n4470), .Z(n4544) );
  NANDN U4921 ( .A(n4473), .B(n4472), .Z(n4477) );
  NANDN U4922 ( .A(n4475), .B(n4474), .Z(n4476) );
  AND U4923 ( .A(n4477), .B(n4476), .Z(n4610) );
  NANDN U4924 ( .A(n4479), .B(n4478), .Z(n4483) );
  NANDN U4925 ( .A(n4481), .B(n4480), .Z(n4482) );
  NAND U4926 ( .A(n4483), .B(n4482), .Z(n4609) );
  XNOR U4927 ( .A(n4610), .B(n4609), .Z(n4611) );
  NAND U4928 ( .A(b[0]), .B(a[42]), .Z(n4484) );
  XNOR U4929 ( .A(b[1]), .B(n4484), .Z(n4486) );
  NANDN U4930 ( .A(b[0]), .B(a[41]), .Z(n4485) );
  NAND U4931 ( .A(n4486), .B(n4485), .Z(n4558) );
  NAND U4932 ( .A(n583), .B(n4487), .Z(n4489) );
  XOR U4933 ( .A(b[29]), .B(a[14]), .Z(n4633) );
  NAND U4934 ( .A(n581), .B(n4633), .Z(n4488) );
  AND U4935 ( .A(n4489), .B(n4488), .Z(n4556) );
  AND U4936 ( .A(b[31]), .B(a[10]), .Z(n4555) );
  XNOR U4937 ( .A(n4556), .B(n4555), .Z(n4557) );
  XNOR U4938 ( .A(n4558), .B(n4557), .Z(n4597) );
  NAND U4939 ( .A(n578), .B(n4490), .Z(n4492) );
  XOR U4940 ( .A(b[23]), .B(a[20]), .Z(n4639) );
  NAND U4941 ( .A(n9268), .B(n4639), .Z(n4491) );
  AND U4942 ( .A(n4492), .B(n4491), .Z(n4630) );
  NAND U4943 ( .A(n569), .B(n4493), .Z(n4495) );
  XOR U4944 ( .A(b[7]), .B(a[36]), .Z(n4642) );
  NAND U4945 ( .A(n7819), .B(n4642), .Z(n4494) );
  AND U4946 ( .A(n4495), .B(n4494), .Z(n4628) );
  NAND U4947 ( .A(n579), .B(n4496), .Z(n4498) );
  XOR U4948 ( .A(b[25]), .B(a[18]), .Z(n4645) );
  NAND U4949 ( .A(n9364), .B(n4645), .Z(n4497) );
  NAND U4950 ( .A(n4498), .B(n4497), .Z(n4627) );
  XNOR U4951 ( .A(n4628), .B(n4627), .Z(n4629) );
  XOR U4952 ( .A(n4630), .B(n4629), .Z(n4598) );
  XNOR U4953 ( .A(n4597), .B(n4598), .Z(n4599) );
  NAND U4954 ( .A(n572), .B(n4499), .Z(n4501) );
  XOR U4955 ( .A(b[13]), .B(a[30]), .Z(n4648) );
  NAND U4956 ( .A(n8585), .B(n4648), .Z(n4500) );
  AND U4957 ( .A(n4501), .B(n4500), .Z(n4592) );
  NAND U4958 ( .A(n571), .B(n4502), .Z(n4504) );
  XOR U4959 ( .A(b[11]), .B(a[32]), .Z(n4651) );
  NAND U4960 ( .A(n8135), .B(n4651), .Z(n4503) );
  NAND U4961 ( .A(n4504), .B(n4503), .Z(n4591) );
  XNOR U4962 ( .A(n4592), .B(n4591), .Z(n4593) );
  NAND U4963 ( .A(n573), .B(n4505), .Z(n4507) );
  XOR U4964 ( .A(b[15]), .B(a[28]), .Z(n4654) );
  NAND U4965 ( .A(n8694), .B(n4654), .Z(n4506) );
  AND U4966 ( .A(n4507), .B(n4506), .Z(n4588) );
  NAND U4967 ( .A(n577), .B(n4508), .Z(n4510) );
  XOR U4968 ( .A(b[21]), .B(a[22]), .Z(n4657) );
  NAND U4969 ( .A(n9216), .B(n4657), .Z(n4509) );
  AND U4970 ( .A(n4510), .B(n4509), .Z(n4586) );
  NAND U4971 ( .A(n570), .B(n4511), .Z(n4513) );
  XOR U4972 ( .A(b[9]), .B(a[34]), .Z(n4660) );
  NAND U4973 ( .A(n8037), .B(n4660), .Z(n4512) );
  NAND U4974 ( .A(n4513), .B(n4512), .Z(n4585) );
  XNOR U4975 ( .A(n4586), .B(n4585), .Z(n4587) );
  XOR U4976 ( .A(n4588), .B(n4587), .Z(n4594) );
  XOR U4977 ( .A(n4593), .B(n4594), .Z(n4600) );
  XOR U4978 ( .A(n4599), .B(n4600), .Z(n4612) );
  XNOR U4979 ( .A(n4611), .B(n4612), .Z(n4543) );
  XNOR U4980 ( .A(n4544), .B(n4543), .Z(n4545) );
  XOR U4981 ( .A(n4546), .B(n4545), .Z(n4664) );
  XNOR U4982 ( .A(n4663), .B(n4664), .Z(n4665) );
  XNOR U4983 ( .A(n4666), .B(n4665), .Z(n4539) );
  XOR U4984 ( .A(n4540), .B(n4539), .Z(n4532) );
  NANDN U4985 ( .A(n4515), .B(n4514), .Z(n4519) );
  NANDN U4986 ( .A(n4517), .B(n4516), .Z(n4518) );
  AND U4987 ( .A(n4519), .B(n4518), .Z(n4531) );
  XOR U4988 ( .A(n4532), .B(n4531), .Z(n4534) );
  XNOR U4989 ( .A(n4533), .B(n4534), .Z(n4525) );
  XNOR U4990 ( .A(n4526), .B(n4525), .Z(n4527) );
  XNOR U4991 ( .A(n4528), .B(n4527), .Z(n4669) );
  XNOR U4992 ( .A(sreg[74]), .B(n4669), .Z(n4671) );
  NANDN U4993 ( .A(sreg[73]), .B(n4520), .Z(n4524) );
  NAND U4994 ( .A(n4522), .B(n4521), .Z(n4523) );
  NAND U4995 ( .A(n4524), .B(n4523), .Z(n4670) );
  XNOR U4996 ( .A(n4671), .B(n4670), .Z(c[74]) );
  NANDN U4997 ( .A(n4526), .B(n4525), .Z(n4530) );
  NANDN U4998 ( .A(n4528), .B(n4527), .Z(n4529) );
  AND U4999 ( .A(n4530), .B(n4529), .Z(n4677) );
  NANDN U5000 ( .A(n4532), .B(n4531), .Z(n4536) );
  NANDN U5001 ( .A(n4534), .B(n4533), .Z(n4535) );
  AND U5002 ( .A(n4536), .B(n4535), .Z(n4675) );
  NANDN U5003 ( .A(n4538), .B(n4537), .Z(n4542) );
  NAND U5004 ( .A(n4540), .B(n4539), .Z(n4541) );
  AND U5005 ( .A(n4542), .B(n4541), .Z(n4682) );
  NANDN U5006 ( .A(n4544), .B(n4543), .Z(n4548) );
  NANDN U5007 ( .A(n4546), .B(n4545), .Z(n4547) );
  AND U5008 ( .A(n4548), .B(n4547), .Z(n4687) );
  NANDN U5009 ( .A(n4550), .B(n4549), .Z(n4554) );
  NAND U5010 ( .A(n4552), .B(n4551), .Z(n4553) );
  AND U5011 ( .A(n4554), .B(n4553), .Z(n4686) );
  XNOR U5012 ( .A(n4687), .B(n4686), .Z(n4689) );
  NANDN U5013 ( .A(n4556), .B(n4555), .Z(n4560) );
  NANDN U5014 ( .A(n4558), .B(n4557), .Z(n4559) );
  AND U5015 ( .A(n4560), .B(n4559), .Z(n4766) );
  NAND U5016 ( .A(n582), .B(n4561), .Z(n4563) );
  XOR U5017 ( .A(b[27]), .B(a[17]), .Z(n4710) );
  NAND U5018 ( .A(n9770), .B(n4710), .Z(n4562) );
  AND U5019 ( .A(n4563), .B(n4562), .Z(n4773) );
  NAND U5020 ( .A(n567), .B(n4564), .Z(n4566) );
  XOR U5021 ( .A(a[39]), .B(b[5]), .Z(n4713) );
  NAND U5022 ( .A(n7235), .B(n4713), .Z(n4565) );
  AND U5023 ( .A(n4566), .B(n4565), .Z(n4771) );
  NAND U5024 ( .A(n9046), .B(n4567), .Z(n4569) );
  XOR U5025 ( .A(b[19]), .B(a[25]), .Z(n4716) );
  NAND U5026 ( .A(n575), .B(n4716), .Z(n4568) );
  NAND U5027 ( .A(n4569), .B(n4568), .Z(n4770) );
  XNOR U5028 ( .A(n4771), .B(n4770), .Z(n4772) );
  XNOR U5029 ( .A(n4773), .B(n4772), .Z(n4764) );
  NAND U5030 ( .A(n9764), .B(n4570), .Z(n4572) );
  XOR U5031 ( .A(b[31]), .B(a[13]), .Z(n4719) );
  NAND U5032 ( .A(n584), .B(n4719), .Z(n4571) );
  AND U5033 ( .A(n4572), .B(n4571), .Z(n4731) );
  NAND U5034 ( .A(n568), .B(n4573), .Z(n4575) );
  XOR U5035 ( .A(a[41]), .B(b[3]), .Z(n4722) );
  NAND U5036 ( .A(n7245), .B(n4722), .Z(n4574) );
  AND U5037 ( .A(n4575), .B(n4574), .Z(n4729) );
  NAND U5038 ( .A(n576), .B(n4576), .Z(n4578) );
  XOR U5039 ( .A(b[17]), .B(a[27]), .Z(n4725) );
  NAND U5040 ( .A(n9141), .B(n4725), .Z(n4577) );
  NAND U5041 ( .A(n4578), .B(n4577), .Z(n4728) );
  XNOR U5042 ( .A(n4729), .B(n4728), .Z(n4730) );
  XOR U5043 ( .A(n4731), .B(n4730), .Z(n4765) );
  XOR U5044 ( .A(n4764), .B(n4765), .Z(n4767) );
  XOR U5045 ( .A(n4766), .B(n4767), .Z(n4699) );
  NANDN U5046 ( .A(n4580), .B(n4579), .Z(n4584) );
  NANDN U5047 ( .A(n4582), .B(n4581), .Z(n4583) );
  AND U5048 ( .A(n4584), .B(n4583), .Z(n4752) );
  NANDN U5049 ( .A(n4586), .B(n4585), .Z(n4590) );
  NANDN U5050 ( .A(n4588), .B(n4587), .Z(n4589) );
  NAND U5051 ( .A(n4590), .B(n4589), .Z(n4753) );
  XNOR U5052 ( .A(n4752), .B(n4753), .Z(n4754) );
  NANDN U5053 ( .A(n4592), .B(n4591), .Z(n4596) );
  NANDN U5054 ( .A(n4594), .B(n4593), .Z(n4595) );
  NAND U5055 ( .A(n4596), .B(n4595), .Z(n4755) );
  XNOR U5056 ( .A(n4754), .B(n4755), .Z(n4698) );
  XNOR U5057 ( .A(n4699), .B(n4698), .Z(n4701) );
  NANDN U5058 ( .A(n4598), .B(n4597), .Z(n4602) );
  NANDN U5059 ( .A(n4600), .B(n4599), .Z(n4601) );
  AND U5060 ( .A(n4602), .B(n4601), .Z(n4700) );
  XOR U5061 ( .A(n4701), .B(n4700), .Z(n4815) );
  NANDN U5062 ( .A(n4604), .B(n4603), .Z(n4608) );
  NANDN U5063 ( .A(n4606), .B(n4605), .Z(n4607) );
  AND U5064 ( .A(n4608), .B(n4607), .Z(n4812) );
  NANDN U5065 ( .A(n4610), .B(n4609), .Z(n4614) );
  NANDN U5066 ( .A(n4612), .B(n4611), .Z(n4613) );
  AND U5067 ( .A(n4614), .B(n4613), .Z(n4695) );
  NANDN U5068 ( .A(n4616), .B(n4615), .Z(n4620) );
  OR U5069 ( .A(n4618), .B(n4617), .Z(n4619) );
  AND U5070 ( .A(n4620), .B(n4619), .Z(n4693) );
  NANDN U5071 ( .A(n4622), .B(n4621), .Z(n4626) );
  NANDN U5072 ( .A(n4624), .B(n4623), .Z(n4625) );
  AND U5073 ( .A(n4626), .B(n4625), .Z(n4759) );
  NANDN U5074 ( .A(n4628), .B(n4627), .Z(n4632) );
  NANDN U5075 ( .A(n4630), .B(n4629), .Z(n4631) );
  NAND U5076 ( .A(n4632), .B(n4631), .Z(n4758) );
  XNOR U5077 ( .A(n4759), .B(n4758), .Z(n4760) );
  NAND U5078 ( .A(n583), .B(n4633), .Z(n4635) );
  XOR U5079 ( .A(b[29]), .B(a[15]), .Z(n4785) );
  NAND U5080 ( .A(n581), .B(n4785), .Z(n4634) );
  AND U5081 ( .A(n4635), .B(n4634), .Z(n4705) );
  AND U5082 ( .A(b[31]), .B(a[11]), .Z(n4704) );
  XNOR U5083 ( .A(n4705), .B(n4704), .Z(n4706) );
  NAND U5084 ( .A(b[0]), .B(a[43]), .Z(n4636) );
  XNOR U5085 ( .A(b[1]), .B(n4636), .Z(n4638) );
  NANDN U5086 ( .A(b[0]), .B(a[42]), .Z(n4637) );
  NAND U5087 ( .A(n4638), .B(n4637), .Z(n4707) );
  XNOR U5088 ( .A(n4706), .B(n4707), .Z(n4746) );
  NAND U5089 ( .A(n578), .B(n4639), .Z(n4641) );
  XOR U5090 ( .A(b[23]), .B(a[21]), .Z(n4788) );
  NAND U5091 ( .A(n9268), .B(n4788), .Z(n4640) );
  AND U5092 ( .A(n4641), .B(n4640), .Z(n4779) );
  NAND U5093 ( .A(n569), .B(n4642), .Z(n4644) );
  XOR U5094 ( .A(b[7]), .B(a[37]), .Z(n4791) );
  NAND U5095 ( .A(n7819), .B(n4791), .Z(n4643) );
  AND U5096 ( .A(n4644), .B(n4643), .Z(n4777) );
  NAND U5097 ( .A(n579), .B(n4645), .Z(n4647) );
  XOR U5098 ( .A(b[25]), .B(a[19]), .Z(n4794) );
  NAND U5099 ( .A(n9364), .B(n4794), .Z(n4646) );
  NAND U5100 ( .A(n4647), .B(n4646), .Z(n4776) );
  XNOR U5101 ( .A(n4777), .B(n4776), .Z(n4778) );
  XOR U5102 ( .A(n4779), .B(n4778), .Z(n4747) );
  XNOR U5103 ( .A(n4746), .B(n4747), .Z(n4748) );
  NAND U5104 ( .A(n572), .B(n4648), .Z(n4650) );
  XOR U5105 ( .A(b[13]), .B(a[31]), .Z(n4797) );
  NAND U5106 ( .A(n8585), .B(n4797), .Z(n4649) );
  AND U5107 ( .A(n4650), .B(n4649), .Z(n4741) );
  NAND U5108 ( .A(n571), .B(n4651), .Z(n4653) );
  XOR U5109 ( .A(b[11]), .B(a[33]), .Z(n4800) );
  NAND U5110 ( .A(n8135), .B(n4800), .Z(n4652) );
  NAND U5111 ( .A(n4653), .B(n4652), .Z(n4740) );
  XNOR U5112 ( .A(n4741), .B(n4740), .Z(n4742) );
  NAND U5113 ( .A(n573), .B(n4654), .Z(n4656) );
  XOR U5114 ( .A(b[15]), .B(a[29]), .Z(n4803) );
  NAND U5115 ( .A(n8694), .B(n4803), .Z(n4655) );
  AND U5116 ( .A(n4656), .B(n4655), .Z(n4737) );
  NAND U5117 ( .A(n577), .B(n4657), .Z(n4659) );
  XOR U5118 ( .A(b[21]), .B(a[23]), .Z(n4806) );
  NAND U5119 ( .A(n9216), .B(n4806), .Z(n4658) );
  AND U5120 ( .A(n4659), .B(n4658), .Z(n4735) );
  NAND U5121 ( .A(n570), .B(n4660), .Z(n4662) );
  XOR U5122 ( .A(b[9]), .B(a[35]), .Z(n4809) );
  NAND U5123 ( .A(n8037), .B(n4809), .Z(n4661) );
  NAND U5124 ( .A(n4662), .B(n4661), .Z(n4734) );
  XNOR U5125 ( .A(n4735), .B(n4734), .Z(n4736) );
  XOR U5126 ( .A(n4737), .B(n4736), .Z(n4743) );
  XOR U5127 ( .A(n4742), .B(n4743), .Z(n4749) );
  XOR U5128 ( .A(n4748), .B(n4749), .Z(n4761) );
  XNOR U5129 ( .A(n4760), .B(n4761), .Z(n4692) );
  XNOR U5130 ( .A(n4693), .B(n4692), .Z(n4694) );
  XOR U5131 ( .A(n4695), .B(n4694), .Z(n4813) );
  XNOR U5132 ( .A(n4812), .B(n4813), .Z(n4814) );
  XNOR U5133 ( .A(n4815), .B(n4814), .Z(n4688) );
  XOR U5134 ( .A(n4689), .B(n4688), .Z(n4681) );
  NANDN U5135 ( .A(n4664), .B(n4663), .Z(n4668) );
  NANDN U5136 ( .A(n4666), .B(n4665), .Z(n4667) );
  AND U5137 ( .A(n4668), .B(n4667), .Z(n4680) );
  XOR U5138 ( .A(n4681), .B(n4680), .Z(n4683) );
  XNOR U5139 ( .A(n4682), .B(n4683), .Z(n4674) );
  XNOR U5140 ( .A(n4675), .B(n4674), .Z(n4676) );
  XNOR U5141 ( .A(n4677), .B(n4676), .Z(n4818) );
  XNOR U5142 ( .A(sreg[75]), .B(n4818), .Z(n4820) );
  NANDN U5143 ( .A(sreg[74]), .B(n4669), .Z(n4673) );
  NAND U5144 ( .A(n4671), .B(n4670), .Z(n4672) );
  NAND U5145 ( .A(n4673), .B(n4672), .Z(n4819) );
  XNOR U5146 ( .A(n4820), .B(n4819), .Z(c[75]) );
  NANDN U5147 ( .A(n4675), .B(n4674), .Z(n4679) );
  NANDN U5148 ( .A(n4677), .B(n4676), .Z(n4678) );
  AND U5149 ( .A(n4679), .B(n4678), .Z(n4826) );
  NANDN U5150 ( .A(n4681), .B(n4680), .Z(n4685) );
  NANDN U5151 ( .A(n4683), .B(n4682), .Z(n4684) );
  AND U5152 ( .A(n4685), .B(n4684), .Z(n4824) );
  NANDN U5153 ( .A(n4687), .B(n4686), .Z(n4691) );
  NAND U5154 ( .A(n4689), .B(n4688), .Z(n4690) );
  AND U5155 ( .A(n4691), .B(n4690), .Z(n4831) );
  NANDN U5156 ( .A(n4693), .B(n4692), .Z(n4697) );
  NANDN U5157 ( .A(n4695), .B(n4694), .Z(n4696) );
  AND U5158 ( .A(n4697), .B(n4696), .Z(n4962) );
  NANDN U5159 ( .A(n4699), .B(n4698), .Z(n4703) );
  NAND U5160 ( .A(n4701), .B(n4700), .Z(n4702) );
  AND U5161 ( .A(n4703), .B(n4702), .Z(n4961) );
  XNOR U5162 ( .A(n4962), .B(n4961), .Z(n4964) );
  NANDN U5163 ( .A(n4705), .B(n4704), .Z(n4709) );
  NANDN U5164 ( .A(n4707), .B(n4706), .Z(n4708) );
  AND U5165 ( .A(n4709), .B(n4708), .Z(n4909) );
  NAND U5166 ( .A(n582), .B(n4710), .Z(n4712) );
  XOR U5167 ( .A(b[27]), .B(a[18]), .Z(n4853) );
  NAND U5168 ( .A(n9770), .B(n4853), .Z(n4711) );
  AND U5169 ( .A(n4712), .B(n4711), .Z(n4916) );
  NAND U5170 ( .A(n567), .B(n4713), .Z(n4715) );
  XOR U5171 ( .A(a[40]), .B(b[5]), .Z(n4856) );
  NAND U5172 ( .A(n7235), .B(n4856), .Z(n4714) );
  AND U5173 ( .A(n4715), .B(n4714), .Z(n4914) );
  NAND U5174 ( .A(n9046), .B(n4716), .Z(n4718) );
  XOR U5175 ( .A(b[19]), .B(a[26]), .Z(n4859) );
  NAND U5176 ( .A(n575), .B(n4859), .Z(n4717) );
  NAND U5177 ( .A(n4718), .B(n4717), .Z(n4913) );
  XNOR U5178 ( .A(n4914), .B(n4913), .Z(n4915) );
  XNOR U5179 ( .A(n4916), .B(n4915), .Z(n4907) );
  NAND U5180 ( .A(n9764), .B(n4719), .Z(n4721) );
  XOR U5181 ( .A(b[31]), .B(a[14]), .Z(n4862) );
  NAND U5182 ( .A(n584), .B(n4862), .Z(n4720) );
  AND U5183 ( .A(n4721), .B(n4720), .Z(n4874) );
  NAND U5184 ( .A(n568), .B(n4722), .Z(n4724) );
  XOR U5185 ( .A(a[42]), .B(b[3]), .Z(n4865) );
  NAND U5186 ( .A(n7245), .B(n4865), .Z(n4723) );
  AND U5187 ( .A(n4724), .B(n4723), .Z(n4872) );
  NAND U5188 ( .A(n576), .B(n4725), .Z(n4727) );
  XOR U5189 ( .A(b[17]), .B(a[28]), .Z(n4868) );
  NAND U5190 ( .A(n9141), .B(n4868), .Z(n4726) );
  NAND U5191 ( .A(n4727), .B(n4726), .Z(n4871) );
  XNOR U5192 ( .A(n4872), .B(n4871), .Z(n4873) );
  XOR U5193 ( .A(n4874), .B(n4873), .Z(n4908) );
  XOR U5194 ( .A(n4907), .B(n4908), .Z(n4910) );
  XOR U5195 ( .A(n4909), .B(n4910), .Z(n4842) );
  NANDN U5196 ( .A(n4729), .B(n4728), .Z(n4733) );
  NANDN U5197 ( .A(n4731), .B(n4730), .Z(n4732) );
  AND U5198 ( .A(n4733), .B(n4732), .Z(n4895) );
  NANDN U5199 ( .A(n4735), .B(n4734), .Z(n4739) );
  NANDN U5200 ( .A(n4737), .B(n4736), .Z(n4738) );
  NAND U5201 ( .A(n4739), .B(n4738), .Z(n4896) );
  XNOR U5202 ( .A(n4895), .B(n4896), .Z(n4897) );
  NANDN U5203 ( .A(n4741), .B(n4740), .Z(n4745) );
  NANDN U5204 ( .A(n4743), .B(n4742), .Z(n4744) );
  NAND U5205 ( .A(n4745), .B(n4744), .Z(n4898) );
  XNOR U5206 ( .A(n4897), .B(n4898), .Z(n4841) );
  XNOR U5207 ( .A(n4842), .B(n4841), .Z(n4844) );
  NANDN U5208 ( .A(n4747), .B(n4746), .Z(n4751) );
  NANDN U5209 ( .A(n4749), .B(n4748), .Z(n4750) );
  AND U5210 ( .A(n4751), .B(n4750), .Z(n4843) );
  XOR U5211 ( .A(n4844), .B(n4843), .Z(n4958) );
  NANDN U5212 ( .A(n4753), .B(n4752), .Z(n4757) );
  NANDN U5213 ( .A(n4755), .B(n4754), .Z(n4756) );
  AND U5214 ( .A(n4757), .B(n4756), .Z(n4955) );
  NANDN U5215 ( .A(n4759), .B(n4758), .Z(n4763) );
  NANDN U5216 ( .A(n4761), .B(n4760), .Z(n4762) );
  AND U5217 ( .A(n4763), .B(n4762), .Z(n4838) );
  NANDN U5218 ( .A(n4765), .B(n4764), .Z(n4769) );
  OR U5219 ( .A(n4767), .B(n4766), .Z(n4768) );
  AND U5220 ( .A(n4769), .B(n4768), .Z(n4836) );
  NANDN U5221 ( .A(n4771), .B(n4770), .Z(n4775) );
  NANDN U5222 ( .A(n4773), .B(n4772), .Z(n4774) );
  AND U5223 ( .A(n4775), .B(n4774), .Z(n4902) );
  NANDN U5224 ( .A(n4777), .B(n4776), .Z(n4781) );
  NANDN U5225 ( .A(n4779), .B(n4778), .Z(n4780) );
  NAND U5226 ( .A(n4781), .B(n4780), .Z(n4901) );
  XNOR U5227 ( .A(n4902), .B(n4901), .Z(n4903) );
  NAND U5228 ( .A(b[0]), .B(a[44]), .Z(n4782) );
  XNOR U5229 ( .A(b[1]), .B(n4782), .Z(n4784) );
  NANDN U5230 ( .A(b[0]), .B(a[43]), .Z(n4783) );
  NAND U5231 ( .A(n4784), .B(n4783), .Z(n4850) );
  NAND U5232 ( .A(n583), .B(n4785), .Z(n4787) );
  XOR U5233 ( .A(b[29]), .B(a[16]), .Z(n4928) );
  NAND U5234 ( .A(n581), .B(n4928), .Z(n4786) );
  AND U5235 ( .A(n4787), .B(n4786), .Z(n4848) );
  AND U5236 ( .A(b[31]), .B(a[12]), .Z(n4847) );
  XNOR U5237 ( .A(n4848), .B(n4847), .Z(n4849) );
  XNOR U5238 ( .A(n4850), .B(n4849), .Z(n4889) );
  NAND U5239 ( .A(n578), .B(n4788), .Z(n4790) );
  XOR U5240 ( .A(b[23]), .B(a[22]), .Z(n4931) );
  NAND U5241 ( .A(n9268), .B(n4931), .Z(n4789) );
  AND U5242 ( .A(n4790), .B(n4789), .Z(n4922) );
  NAND U5243 ( .A(n569), .B(n4791), .Z(n4793) );
  XOR U5244 ( .A(b[7]), .B(a[38]), .Z(n4934) );
  NAND U5245 ( .A(n7819), .B(n4934), .Z(n4792) );
  AND U5246 ( .A(n4793), .B(n4792), .Z(n4920) );
  NAND U5247 ( .A(n579), .B(n4794), .Z(n4796) );
  XOR U5248 ( .A(b[25]), .B(a[20]), .Z(n4937) );
  NAND U5249 ( .A(n9364), .B(n4937), .Z(n4795) );
  NAND U5250 ( .A(n4796), .B(n4795), .Z(n4919) );
  XNOR U5251 ( .A(n4920), .B(n4919), .Z(n4921) );
  XOR U5252 ( .A(n4922), .B(n4921), .Z(n4890) );
  XNOR U5253 ( .A(n4889), .B(n4890), .Z(n4891) );
  NAND U5254 ( .A(n572), .B(n4797), .Z(n4799) );
  XOR U5255 ( .A(b[13]), .B(a[32]), .Z(n4940) );
  NAND U5256 ( .A(n8585), .B(n4940), .Z(n4798) );
  AND U5257 ( .A(n4799), .B(n4798), .Z(n4884) );
  NAND U5258 ( .A(n571), .B(n4800), .Z(n4802) );
  XOR U5259 ( .A(b[11]), .B(a[34]), .Z(n4943) );
  NAND U5260 ( .A(n8135), .B(n4943), .Z(n4801) );
  NAND U5261 ( .A(n4802), .B(n4801), .Z(n4883) );
  XNOR U5262 ( .A(n4884), .B(n4883), .Z(n4885) );
  NAND U5263 ( .A(n573), .B(n4803), .Z(n4805) );
  XOR U5264 ( .A(b[15]), .B(a[30]), .Z(n4946) );
  NAND U5265 ( .A(n8694), .B(n4946), .Z(n4804) );
  AND U5266 ( .A(n4805), .B(n4804), .Z(n4880) );
  NAND U5267 ( .A(n577), .B(n4806), .Z(n4808) );
  XOR U5268 ( .A(b[21]), .B(a[24]), .Z(n4949) );
  NAND U5269 ( .A(n9216), .B(n4949), .Z(n4807) );
  AND U5270 ( .A(n4808), .B(n4807), .Z(n4878) );
  NAND U5271 ( .A(n570), .B(n4809), .Z(n4811) );
  XOR U5272 ( .A(b[9]), .B(a[36]), .Z(n4952) );
  NAND U5273 ( .A(n8037), .B(n4952), .Z(n4810) );
  NAND U5274 ( .A(n4811), .B(n4810), .Z(n4877) );
  XNOR U5275 ( .A(n4878), .B(n4877), .Z(n4879) );
  XOR U5276 ( .A(n4880), .B(n4879), .Z(n4886) );
  XOR U5277 ( .A(n4885), .B(n4886), .Z(n4892) );
  XOR U5278 ( .A(n4891), .B(n4892), .Z(n4904) );
  XNOR U5279 ( .A(n4903), .B(n4904), .Z(n4835) );
  XNOR U5280 ( .A(n4836), .B(n4835), .Z(n4837) );
  XOR U5281 ( .A(n4838), .B(n4837), .Z(n4956) );
  XNOR U5282 ( .A(n4955), .B(n4956), .Z(n4957) );
  XNOR U5283 ( .A(n4958), .B(n4957), .Z(n4963) );
  XOR U5284 ( .A(n4964), .B(n4963), .Z(n4830) );
  NANDN U5285 ( .A(n4813), .B(n4812), .Z(n4817) );
  NANDN U5286 ( .A(n4815), .B(n4814), .Z(n4816) );
  AND U5287 ( .A(n4817), .B(n4816), .Z(n4829) );
  XOR U5288 ( .A(n4830), .B(n4829), .Z(n4832) );
  XNOR U5289 ( .A(n4831), .B(n4832), .Z(n4823) );
  XNOR U5290 ( .A(n4824), .B(n4823), .Z(n4825) );
  XNOR U5291 ( .A(n4826), .B(n4825), .Z(n4967) );
  XNOR U5292 ( .A(sreg[76]), .B(n4967), .Z(n4969) );
  NANDN U5293 ( .A(sreg[75]), .B(n4818), .Z(n4822) );
  NAND U5294 ( .A(n4820), .B(n4819), .Z(n4821) );
  NAND U5295 ( .A(n4822), .B(n4821), .Z(n4968) );
  XNOR U5296 ( .A(n4969), .B(n4968), .Z(c[76]) );
  NANDN U5297 ( .A(n4824), .B(n4823), .Z(n4828) );
  NANDN U5298 ( .A(n4826), .B(n4825), .Z(n4827) );
  AND U5299 ( .A(n4828), .B(n4827), .Z(n4975) );
  NANDN U5300 ( .A(n4830), .B(n4829), .Z(n4834) );
  NANDN U5301 ( .A(n4832), .B(n4831), .Z(n4833) );
  AND U5302 ( .A(n4834), .B(n4833), .Z(n4973) );
  NANDN U5303 ( .A(n4836), .B(n4835), .Z(n4840) );
  NANDN U5304 ( .A(n4838), .B(n4837), .Z(n4839) );
  AND U5305 ( .A(n4840), .B(n4839), .Z(n4985) );
  NANDN U5306 ( .A(n4842), .B(n4841), .Z(n4846) );
  NAND U5307 ( .A(n4844), .B(n4843), .Z(n4845) );
  AND U5308 ( .A(n4846), .B(n4845), .Z(n4984) );
  XNOR U5309 ( .A(n4985), .B(n4984), .Z(n4987) );
  NANDN U5310 ( .A(n4848), .B(n4847), .Z(n4852) );
  NANDN U5311 ( .A(n4850), .B(n4849), .Z(n4851) );
  AND U5312 ( .A(n4852), .B(n4851), .Z(n5062) );
  NAND U5313 ( .A(n582), .B(n4853), .Z(n4855) );
  XOR U5314 ( .A(b[27]), .B(a[19]), .Z(n5008) );
  NAND U5315 ( .A(n9770), .B(n5008), .Z(n4854) );
  AND U5316 ( .A(n4855), .B(n4854), .Z(n5069) );
  NAND U5317 ( .A(n567), .B(n4856), .Z(n4858) );
  XOR U5318 ( .A(a[41]), .B(b[5]), .Z(n5011) );
  NAND U5319 ( .A(n7235), .B(n5011), .Z(n4857) );
  AND U5320 ( .A(n4858), .B(n4857), .Z(n5067) );
  NAND U5321 ( .A(n9046), .B(n4859), .Z(n4861) );
  XOR U5322 ( .A(b[19]), .B(a[27]), .Z(n5014) );
  NAND U5323 ( .A(n575), .B(n5014), .Z(n4860) );
  NAND U5324 ( .A(n4861), .B(n4860), .Z(n5066) );
  XNOR U5325 ( .A(n5067), .B(n5066), .Z(n5068) );
  XNOR U5326 ( .A(n5069), .B(n5068), .Z(n5060) );
  NAND U5327 ( .A(n9764), .B(n4862), .Z(n4864) );
  XOR U5328 ( .A(b[31]), .B(a[15]), .Z(n5017) );
  NAND U5329 ( .A(n584), .B(n5017), .Z(n4863) );
  AND U5330 ( .A(n4864), .B(n4863), .Z(n5029) );
  NAND U5331 ( .A(n568), .B(n4865), .Z(n4867) );
  XOR U5332 ( .A(a[43]), .B(b[3]), .Z(n5020) );
  NAND U5333 ( .A(n7245), .B(n5020), .Z(n4866) );
  AND U5334 ( .A(n4867), .B(n4866), .Z(n5027) );
  NAND U5335 ( .A(n576), .B(n4868), .Z(n4870) );
  XOR U5336 ( .A(b[17]), .B(a[29]), .Z(n5023) );
  NAND U5337 ( .A(n9141), .B(n5023), .Z(n4869) );
  NAND U5338 ( .A(n4870), .B(n4869), .Z(n5026) );
  XNOR U5339 ( .A(n5027), .B(n5026), .Z(n5028) );
  XOR U5340 ( .A(n5029), .B(n5028), .Z(n5061) );
  XOR U5341 ( .A(n5060), .B(n5061), .Z(n5063) );
  XOR U5342 ( .A(n5062), .B(n5063), .Z(n4997) );
  NANDN U5343 ( .A(n4872), .B(n4871), .Z(n4876) );
  NANDN U5344 ( .A(n4874), .B(n4873), .Z(n4875) );
  AND U5345 ( .A(n4876), .B(n4875), .Z(n5050) );
  NANDN U5346 ( .A(n4878), .B(n4877), .Z(n4882) );
  NANDN U5347 ( .A(n4880), .B(n4879), .Z(n4881) );
  NAND U5348 ( .A(n4882), .B(n4881), .Z(n5051) );
  XNOR U5349 ( .A(n5050), .B(n5051), .Z(n5052) );
  NANDN U5350 ( .A(n4884), .B(n4883), .Z(n4888) );
  NANDN U5351 ( .A(n4886), .B(n4885), .Z(n4887) );
  NAND U5352 ( .A(n4888), .B(n4887), .Z(n5053) );
  XNOR U5353 ( .A(n5052), .B(n5053), .Z(n4996) );
  XNOR U5354 ( .A(n4997), .B(n4996), .Z(n4999) );
  NANDN U5355 ( .A(n4890), .B(n4889), .Z(n4894) );
  NANDN U5356 ( .A(n4892), .B(n4891), .Z(n4893) );
  AND U5357 ( .A(n4894), .B(n4893), .Z(n4998) );
  XOR U5358 ( .A(n4999), .B(n4998), .Z(n5111) );
  NANDN U5359 ( .A(n4896), .B(n4895), .Z(n4900) );
  NANDN U5360 ( .A(n4898), .B(n4897), .Z(n4899) );
  AND U5361 ( .A(n4900), .B(n4899), .Z(n5108) );
  NANDN U5362 ( .A(n4902), .B(n4901), .Z(n4906) );
  NANDN U5363 ( .A(n4904), .B(n4903), .Z(n4905) );
  AND U5364 ( .A(n4906), .B(n4905), .Z(n4993) );
  NANDN U5365 ( .A(n4908), .B(n4907), .Z(n4912) );
  OR U5366 ( .A(n4910), .B(n4909), .Z(n4911) );
  AND U5367 ( .A(n4912), .B(n4911), .Z(n4991) );
  NANDN U5368 ( .A(n4914), .B(n4913), .Z(n4918) );
  NANDN U5369 ( .A(n4916), .B(n4915), .Z(n4917) );
  AND U5370 ( .A(n4918), .B(n4917), .Z(n5057) );
  NANDN U5371 ( .A(n4920), .B(n4919), .Z(n4924) );
  NANDN U5372 ( .A(n4922), .B(n4921), .Z(n4923) );
  NAND U5373 ( .A(n4924), .B(n4923), .Z(n5056) );
  XNOR U5374 ( .A(n5057), .B(n5056), .Z(n5059) );
  NAND U5375 ( .A(b[0]), .B(a[45]), .Z(n4925) );
  XNOR U5376 ( .A(b[1]), .B(n4925), .Z(n4927) );
  NANDN U5377 ( .A(b[0]), .B(a[44]), .Z(n4926) );
  NAND U5378 ( .A(n4927), .B(n4926), .Z(n5005) );
  NAND U5379 ( .A(n583), .B(n4928), .Z(n4930) );
  XOR U5380 ( .A(b[29]), .B(a[17]), .Z(n5078) );
  NAND U5381 ( .A(n581), .B(n5078), .Z(n4929) );
  AND U5382 ( .A(n4930), .B(n4929), .Z(n5003) );
  AND U5383 ( .A(b[31]), .B(a[13]), .Z(n5002) );
  XNOR U5384 ( .A(n5003), .B(n5002), .Z(n5004) );
  XNOR U5385 ( .A(n5005), .B(n5004), .Z(n5045) );
  NAND U5386 ( .A(n578), .B(n4931), .Z(n4933) );
  XOR U5387 ( .A(b[23]), .B(a[23]), .Z(n5084) );
  NAND U5388 ( .A(n9268), .B(n5084), .Z(n4932) );
  AND U5389 ( .A(n4933), .B(n4932), .Z(n5074) );
  NAND U5390 ( .A(n569), .B(n4934), .Z(n4936) );
  XOR U5391 ( .A(b[7]), .B(a[39]), .Z(n5087) );
  NAND U5392 ( .A(n7819), .B(n5087), .Z(n4935) );
  AND U5393 ( .A(n4936), .B(n4935), .Z(n5073) );
  NAND U5394 ( .A(n579), .B(n4937), .Z(n4939) );
  XOR U5395 ( .A(b[25]), .B(a[21]), .Z(n5090) );
  NAND U5396 ( .A(n9364), .B(n5090), .Z(n4938) );
  NAND U5397 ( .A(n4939), .B(n4938), .Z(n5072) );
  XOR U5398 ( .A(n5073), .B(n5072), .Z(n5075) );
  XOR U5399 ( .A(n5074), .B(n5075), .Z(n5044) );
  XOR U5400 ( .A(n5045), .B(n5044), .Z(n5047) );
  NAND U5401 ( .A(n572), .B(n4940), .Z(n4942) );
  XOR U5402 ( .A(b[13]), .B(a[33]), .Z(n5093) );
  NAND U5403 ( .A(n8585), .B(n5093), .Z(n4941) );
  AND U5404 ( .A(n4942), .B(n4941), .Z(n5039) );
  NAND U5405 ( .A(n571), .B(n4943), .Z(n4945) );
  XOR U5406 ( .A(b[11]), .B(a[35]), .Z(n5096) );
  NAND U5407 ( .A(n8135), .B(n5096), .Z(n4944) );
  NAND U5408 ( .A(n4945), .B(n4944), .Z(n5038) );
  XNOR U5409 ( .A(n5039), .B(n5038), .Z(n5041) );
  NAND U5410 ( .A(n573), .B(n4946), .Z(n4948) );
  XOR U5411 ( .A(b[15]), .B(a[31]), .Z(n5099) );
  NAND U5412 ( .A(n8694), .B(n5099), .Z(n4947) );
  AND U5413 ( .A(n4948), .B(n4947), .Z(n5035) );
  NAND U5414 ( .A(n577), .B(n4949), .Z(n4951) );
  XOR U5415 ( .A(b[21]), .B(a[25]), .Z(n5102) );
  NAND U5416 ( .A(n9216), .B(n5102), .Z(n4950) );
  AND U5417 ( .A(n4951), .B(n4950), .Z(n5033) );
  NAND U5418 ( .A(n570), .B(n4952), .Z(n4954) );
  XOR U5419 ( .A(b[9]), .B(a[37]), .Z(n5105) );
  NAND U5420 ( .A(n8037), .B(n5105), .Z(n4953) );
  NAND U5421 ( .A(n4954), .B(n4953), .Z(n5032) );
  XNOR U5422 ( .A(n5033), .B(n5032), .Z(n5034) );
  XNOR U5423 ( .A(n5035), .B(n5034), .Z(n5040) );
  XOR U5424 ( .A(n5041), .B(n5040), .Z(n5046) );
  XNOR U5425 ( .A(n5047), .B(n5046), .Z(n5058) );
  XNOR U5426 ( .A(n5059), .B(n5058), .Z(n4990) );
  XNOR U5427 ( .A(n4991), .B(n4990), .Z(n4992) );
  XOR U5428 ( .A(n4993), .B(n4992), .Z(n5109) );
  XNOR U5429 ( .A(n5108), .B(n5109), .Z(n5110) );
  XNOR U5430 ( .A(n5111), .B(n5110), .Z(n4986) );
  XOR U5431 ( .A(n4987), .B(n4986), .Z(n4979) );
  NANDN U5432 ( .A(n4956), .B(n4955), .Z(n4960) );
  NANDN U5433 ( .A(n4958), .B(n4957), .Z(n4959) );
  AND U5434 ( .A(n4960), .B(n4959), .Z(n4978) );
  XNOR U5435 ( .A(n4979), .B(n4978), .Z(n4980) );
  NANDN U5436 ( .A(n4962), .B(n4961), .Z(n4966) );
  NAND U5437 ( .A(n4964), .B(n4963), .Z(n4965) );
  NAND U5438 ( .A(n4966), .B(n4965), .Z(n4981) );
  XNOR U5439 ( .A(n4980), .B(n4981), .Z(n4972) );
  XNOR U5440 ( .A(n4973), .B(n4972), .Z(n4974) );
  XNOR U5441 ( .A(n4975), .B(n4974), .Z(n5114) );
  XNOR U5442 ( .A(sreg[77]), .B(n5114), .Z(n5116) );
  NANDN U5443 ( .A(sreg[76]), .B(n4967), .Z(n4971) );
  NAND U5444 ( .A(n4969), .B(n4968), .Z(n4970) );
  NAND U5445 ( .A(n4971), .B(n4970), .Z(n5115) );
  XNOR U5446 ( .A(n5116), .B(n5115), .Z(c[77]) );
  NANDN U5447 ( .A(n4973), .B(n4972), .Z(n4977) );
  NANDN U5448 ( .A(n4975), .B(n4974), .Z(n4976) );
  AND U5449 ( .A(n4977), .B(n4976), .Z(n5122) );
  NANDN U5450 ( .A(n4979), .B(n4978), .Z(n4983) );
  NANDN U5451 ( .A(n4981), .B(n4980), .Z(n4982) );
  AND U5452 ( .A(n4983), .B(n4982), .Z(n5120) );
  NANDN U5453 ( .A(n4985), .B(n4984), .Z(n4989) );
  NAND U5454 ( .A(n4987), .B(n4986), .Z(n4988) );
  AND U5455 ( .A(n4989), .B(n4988), .Z(n5127) );
  NANDN U5456 ( .A(n4991), .B(n4990), .Z(n4995) );
  NANDN U5457 ( .A(n4993), .B(n4992), .Z(n4994) );
  AND U5458 ( .A(n4995), .B(n4994), .Z(n5132) );
  NANDN U5459 ( .A(n4997), .B(n4996), .Z(n5001) );
  NAND U5460 ( .A(n4999), .B(n4998), .Z(n5000) );
  AND U5461 ( .A(n5001), .B(n5000), .Z(n5131) );
  XNOR U5462 ( .A(n5132), .B(n5131), .Z(n5134) );
  NANDN U5463 ( .A(n5003), .B(n5002), .Z(n5007) );
  NANDN U5464 ( .A(n5005), .B(n5004), .Z(n5006) );
  AND U5465 ( .A(n5007), .B(n5006), .Z(n5197) );
  NAND U5466 ( .A(n582), .B(n5008), .Z(n5010) );
  XOR U5467 ( .A(b[27]), .B(a[20]), .Z(n5143) );
  NAND U5468 ( .A(n9770), .B(n5143), .Z(n5009) );
  AND U5469 ( .A(n5010), .B(n5009), .Z(n5204) );
  NAND U5470 ( .A(n567), .B(n5011), .Z(n5013) );
  XOR U5471 ( .A(a[42]), .B(b[5]), .Z(n5146) );
  NAND U5472 ( .A(n7235), .B(n5146), .Z(n5012) );
  AND U5473 ( .A(n5013), .B(n5012), .Z(n5202) );
  NAND U5474 ( .A(n9046), .B(n5014), .Z(n5016) );
  XOR U5475 ( .A(b[19]), .B(a[28]), .Z(n5149) );
  NAND U5476 ( .A(n575), .B(n5149), .Z(n5015) );
  NAND U5477 ( .A(n5016), .B(n5015), .Z(n5201) );
  XNOR U5478 ( .A(n5202), .B(n5201), .Z(n5203) );
  XNOR U5479 ( .A(n5204), .B(n5203), .Z(n5195) );
  NAND U5480 ( .A(n9764), .B(n5017), .Z(n5019) );
  XOR U5481 ( .A(b[31]), .B(a[16]), .Z(n5152) );
  NAND U5482 ( .A(n584), .B(n5152), .Z(n5018) );
  AND U5483 ( .A(n5019), .B(n5018), .Z(n5164) );
  NAND U5484 ( .A(n568), .B(n5020), .Z(n5022) );
  XOR U5485 ( .A(a[44]), .B(b[3]), .Z(n5155) );
  NAND U5486 ( .A(n7245), .B(n5155), .Z(n5021) );
  AND U5487 ( .A(n5022), .B(n5021), .Z(n5162) );
  NAND U5488 ( .A(n576), .B(n5023), .Z(n5025) );
  XOR U5489 ( .A(b[17]), .B(a[30]), .Z(n5158) );
  NAND U5490 ( .A(n9141), .B(n5158), .Z(n5024) );
  NAND U5491 ( .A(n5025), .B(n5024), .Z(n5161) );
  XNOR U5492 ( .A(n5162), .B(n5161), .Z(n5163) );
  XOR U5493 ( .A(n5164), .B(n5163), .Z(n5196) );
  XOR U5494 ( .A(n5195), .B(n5196), .Z(n5198) );
  XOR U5495 ( .A(n5197), .B(n5198), .Z(n5244) );
  NANDN U5496 ( .A(n5027), .B(n5026), .Z(n5031) );
  NANDN U5497 ( .A(n5029), .B(n5028), .Z(n5030) );
  AND U5498 ( .A(n5031), .B(n5030), .Z(n5185) );
  NANDN U5499 ( .A(n5033), .B(n5032), .Z(n5037) );
  NANDN U5500 ( .A(n5035), .B(n5034), .Z(n5036) );
  NAND U5501 ( .A(n5037), .B(n5036), .Z(n5186) );
  XNOR U5502 ( .A(n5185), .B(n5186), .Z(n5187) );
  NANDN U5503 ( .A(n5039), .B(n5038), .Z(n5043) );
  NAND U5504 ( .A(n5041), .B(n5040), .Z(n5042) );
  NAND U5505 ( .A(n5043), .B(n5042), .Z(n5188) );
  XNOR U5506 ( .A(n5187), .B(n5188), .Z(n5243) );
  XNOR U5507 ( .A(n5244), .B(n5243), .Z(n5246) );
  NAND U5508 ( .A(n5045), .B(n5044), .Z(n5049) );
  NAND U5509 ( .A(n5047), .B(n5046), .Z(n5048) );
  AND U5510 ( .A(n5049), .B(n5048), .Z(n5245) );
  XOR U5511 ( .A(n5246), .B(n5245), .Z(n5258) );
  NANDN U5512 ( .A(n5051), .B(n5050), .Z(n5055) );
  NANDN U5513 ( .A(n5053), .B(n5052), .Z(n5054) );
  AND U5514 ( .A(n5055), .B(n5054), .Z(n5255) );
  NANDN U5515 ( .A(n5061), .B(n5060), .Z(n5065) );
  OR U5516 ( .A(n5063), .B(n5062), .Z(n5064) );
  AND U5517 ( .A(n5065), .B(n5064), .Z(n5250) );
  NANDN U5518 ( .A(n5067), .B(n5066), .Z(n5071) );
  NANDN U5519 ( .A(n5069), .B(n5068), .Z(n5070) );
  AND U5520 ( .A(n5071), .B(n5070), .Z(n5192) );
  NANDN U5521 ( .A(n5073), .B(n5072), .Z(n5077) );
  OR U5522 ( .A(n5075), .B(n5074), .Z(n5076) );
  NAND U5523 ( .A(n5077), .B(n5076), .Z(n5191) );
  XNOR U5524 ( .A(n5192), .B(n5191), .Z(n5194) );
  NAND U5525 ( .A(n583), .B(n5078), .Z(n5080) );
  XOR U5526 ( .A(b[29]), .B(a[18]), .Z(n5216) );
  NAND U5527 ( .A(n581), .B(n5216), .Z(n5079) );
  AND U5528 ( .A(n5080), .B(n5079), .Z(n5138) );
  AND U5529 ( .A(b[31]), .B(a[14]), .Z(n5137) );
  XNOR U5530 ( .A(n5138), .B(n5137), .Z(n5139) );
  NAND U5531 ( .A(b[0]), .B(a[46]), .Z(n5081) );
  XNOR U5532 ( .A(b[1]), .B(n5081), .Z(n5083) );
  NANDN U5533 ( .A(b[0]), .B(a[45]), .Z(n5082) );
  NAND U5534 ( .A(n5083), .B(n5082), .Z(n5140) );
  XNOR U5535 ( .A(n5139), .B(n5140), .Z(n5180) );
  NAND U5536 ( .A(n578), .B(n5084), .Z(n5086) );
  XOR U5537 ( .A(b[23]), .B(a[24]), .Z(n5219) );
  NAND U5538 ( .A(n9268), .B(n5219), .Z(n5085) );
  AND U5539 ( .A(n5086), .B(n5085), .Z(n5209) );
  NAND U5540 ( .A(n569), .B(n5087), .Z(n5089) );
  XOR U5541 ( .A(b[7]), .B(a[40]), .Z(n5222) );
  NAND U5542 ( .A(n7819), .B(n5222), .Z(n5088) );
  AND U5543 ( .A(n5089), .B(n5088), .Z(n5208) );
  NAND U5544 ( .A(n579), .B(n5090), .Z(n5092) );
  XOR U5545 ( .A(b[25]), .B(a[22]), .Z(n5225) );
  NAND U5546 ( .A(n9364), .B(n5225), .Z(n5091) );
  NAND U5547 ( .A(n5092), .B(n5091), .Z(n5207) );
  XOR U5548 ( .A(n5208), .B(n5207), .Z(n5210) );
  XOR U5549 ( .A(n5209), .B(n5210), .Z(n5179) );
  XOR U5550 ( .A(n5180), .B(n5179), .Z(n5182) );
  NAND U5551 ( .A(n572), .B(n5093), .Z(n5095) );
  XOR U5552 ( .A(b[13]), .B(a[34]), .Z(n5228) );
  NAND U5553 ( .A(n8585), .B(n5228), .Z(n5094) );
  AND U5554 ( .A(n5095), .B(n5094), .Z(n5174) );
  NAND U5555 ( .A(n571), .B(n5096), .Z(n5098) );
  XOR U5556 ( .A(b[11]), .B(a[36]), .Z(n5231) );
  NAND U5557 ( .A(n8135), .B(n5231), .Z(n5097) );
  NAND U5558 ( .A(n5098), .B(n5097), .Z(n5173) );
  XNOR U5559 ( .A(n5174), .B(n5173), .Z(n5176) );
  NAND U5560 ( .A(n573), .B(n5099), .Z(n5101) );
  XOR U5561 ( .A(b[15]), .B(a[32]), .Z(n5234) );
  NAND U5562 ( .A(n8694), .B(n5234), .Z(n5100) );
  AND U5563 ( .A(n5101), .B(n5100), .Z(n5170) );
  NAND U5564 ( .A(n577), .B(n5102), .Z(n5104) );
  XOR U5565 ( .A(b[21]), .B(a[26]), .Z(n5237) );
  NAND U5566 ( .A(n9216), .B(n5237), .Z(n5103) );
  AND U5567 ( .A(n5104), .B(n5103), .Z(n5168) );
  NAND U5568 ( .A(n570), .B(n5105), .Z(n5107) );
  XOR U5569 ( .A(b[9]), .B(a[38]), .Z(n5240) );
  NAND U5570 ( .A(n8037), .B(n5240), .Z(n5106) );
  NAND U5571 ( .A(n5107), .B(n5106), .Z(n5167) );
  XNOR U5572 ( .A(n5168), .B(n5167), .Z(n5169) );
  XNOR U5573 ( .A(n5170), .B(n5169), .Z(n5175) );
  XOR U5574 ( .A(n5176), .B(n5175), .Z(n5181) );
  XNOR U5575 ( .A(n5182), .B(n5181), .Z(n5193) );
  XNOR U5576 ( .A(n5194), .B(n5193), .Z(n5249) );
  XNOR U5577 ( .A(n5250), .B(n5249), .Z(n5251) );
  XOR U5578 ( .A(n5252), .B(n5251), .Z(n5256) );
  XNOR U5579 ( .A(n5255), .B(n5256), .Z(n5257) );
  XNOR U5580 ( .A(n5258), .B(n5257), .Z(n5133) );
  XOR U5581 ( .A(n5134), .B(n5133), .Z(n5126) );
  NANDN U5582 ( .A(n5109), .B(n5108), .Z(n5113) );
  NANDN U5583 ( .A(n5111), .B(n5110), .Z(n5112) );
  AND U5584 ( .A(n5113), .B(n5112), .Z(n5125) );
  XOR U5585 ( .A(n5126), .B(n5125), .Z(n5128) );
  XNOR U5586 ( .A(n5127), .B(n5128), .Z(n5119) );
  XNOR U5587 ( .A(n5120), .B(n5119), .Z(n5121) );
  XNOR U5588 ( .A(n5122), .B(n5121), .Z(n5261) );
  XNOR U5589 ( .A(sreg[78]), .B(n5261), .Z(n5263) );
  NANDN U5590 ( .A(sreg[77]), .B(n5114), .Z(n5118) );
  NAND U5591 ( .A(n5116), .B(n5115), .Z(n5117) );
  NAND U5592 ( .A(n5118), .B(n5117), .Z(n5262) );
  XNOR U5593 ( .A(n5263), .B(n5262), .Z(c[78]) );
  NANDN U5594 ( .A(n5120), .B(n5119), .Z(n5124) );
  NANDN U5595 ( .A(n5122), .B(n5121), .Z(n5123) );
  AND U5596 ( .A(n5124), .B(n5123), .Z(n5269) );
  NANDN U5597 ( .A(n5126), .B(n5125), .Z(n5130) );
  NANDN U5598 ( .A(n5128), .B(n5127), .Z(n5129) );
  AND U5599 ( .A(n5130), .B(n5129), .Z(n5267) );
  NANDN U5600 ( .A(n5132), .B(n5131), .Z(n5136) );
  NAND U5601 ( .A(n5134), .B(n5133), .Z(n5135) );
  AND U5602 ( .A(n5136), .B(n5135), .Z(n5274) );
  NANDN U5603 ( .A(n5138), .B(n5137), .Z(n5142) );
  NANDN U5604 ( .A(n5140), .B(n5139), .Z(n5141) );
  AND U5605 ( .A(n5142), .B(n5141), .Z(n5344) );
  NAND U5606 ( .A(n582), .B(n5143), .Z(n5145) );
  XOR U5607 ( .A(b[27]), .B(a[21]), .Z(n5290) );
  NAND U5608 ( .A(n9770), .B(n5290), .Z(n5144) );
  AND U5609 ( .A(n5145), .B(n5144), .Z(n5351) );
  NAND U5610 ( .A(n567), .B(n5146), .Z(n5148) );
  XOR U5611 ( .A(a[43]), .B(b[5]), .Z(n5293) );
  NAND U5612 ( .A(n7235), .B(n5293), .Z(n5147) );
  AND U5613 ( .A(n5148), .B(n5147), .Z(n5349) );
  NAND U5614 ( .A(n9046), .B(n5149), .Z(n5151) );
  XOR U5615 ( .A(b[19]), .B(a[29]), .Z(n5296) );
  NAND U5616 ( .A(n575), .B(n5296), .Z(n5150) );
  NAND U5617 ( .A(n5151), .B(n5150), .Z(n5348) );
  XNOR U5618 ( .A(n5349), .B(n5348), .Z(n5350) );
  XNOR U5619 ( .A(n5351), .B(n5350), .Z(n5342) );
  NAND U5620 ( .A(n9764), .B(n5152), .Z(n5154) );
  XOR U5621 ( .A(b[31]), .B(a[17]), .Z(n5299) );
  NAND U5622 ( .A(n584), .B(n5299), .Z(n5153) );
  AND U5623 ( .A(n5154), .B(n5153), .Z(n5311) );
  NAND U5624 ( .A(n568), .B(n5155), .Z(n5157) );
  XOR U5625 ( .A(a[45]), .B(b[3]), .Z(n5302) );
  NAND U5626 ( .A(n7245), .B(n5302), .Z(n5156) );
  AND U5627 ( .A(n5157), .B(n5156), .Z(n5309) );
  NAND U5628 ( .A(n576), .B(n5158), .Z(n5160) );
  XOR U5629 ( .A(b[17]), .B(a[31]), .Z(n5305) );
  NAND U5630 ( .A(n9141), .B(n5305), .Z(n5159) );
  NAND U5631 ( .A(n5160), .B(n5159), .Z(n5308) );
  XNOR U5632 ( .A(n5309), .B(n5308), .Z(n5310) );
  XOR U5633 ( .A(n5311), .B(n5310), .Z(n5343) );
  XOR U5634 ( .A(n5342), .B(n5343), .Z(n5345) );
  XOR U5635 ( .A(n5344), .B(n5345), .Z(n5391) );
  NANDN U5636 ( .A(n5162), .B(n5161), .Z(n5166) );
  NANDN U5637 ( .A(n5164), .B(n5163), .Z(n5165) );
  AND U5638 ( .A(n5166), .B(n5165), .Z(n5332) );
  NANDN U5639 ( .A(n5168), .B(n5167), .Z(n5172) );
  NANDN U5640 ( .A(n5170), .B(n5169), .Z(n5171) );
  NAND U5641 ( .A(n5172), .B(n5171), .Z(n5333) );
  XNOR U5642 ( .A(n5332), .B(n5333), .Z(n5334) );
  NANDN U5643 ( .A(n5174), .B(n5173), .Z(n5178) );
  NAND U5644 ( .A(n5176), .B(n5175), .Z(n5177) );
  NAND U5645 ( .A(n5178), .B(n5177), .Z(n5335) );
  XNOR U5646 ( .A(n5334), .B(n5335), .Z(n5390) );
  XNOR U5647 ( .A(n5391), .B(n5390), .Z(n5393) );
  NAND U5648 ( .A(n5180), .B(n5179), .Z(n5184) );
  NAND U5649 ( .A(n5182), .B(n5181), .Z(n5183) );
  AND U5650 ( .A(n5184), .B(n5183), .Z(n5392) );
  XOR U5651 ( .A(n5393), .B(n5392), .Z(n5404) );
  NANDN U5652 ( .A(n5186), .B(n5185), .Z(n5190) );
  NANDN U5653 ( .A(n5188), .B(n5187), .Z(n5189) );
  AND U5654 ( .A(n5190), .B(n5189), .Z(n5402) );
  NANDN U5655 ( .A(n5196), .B(n5195), .Z(n5200) );
  OR U5656 ( .A(n5198), .B(n5197), .Z(n5199) );
  AND U5657 ( .A(n5200), .B(n5199), .Z(n5397) );
  NANDN U5658 ( .A(n5202), .B(n5201), .Z(n5206) );
  NANDN U5659 ( .A(n5204), .B(n5203), .Z(n5205) );
  AND U5660 ( .A(n5206), .B(n5205), .Z(n5339) );
  NANDN U5661 ( .A(n5208), .B(n5207), .Z(n5212) );
  OR U5662 ( .A(n5210), .B(n5209), .Z(n5211) );
  NAND U5663 ( .A(n5212), .B(n5211), .Z(n5338) );
  XNOR U5664 ( .A(n5339), .B(n5338), .Z(n5341) );
  NAND U5665 ( .A(b[0]), .B(a[47]), .Z(n5213) );
  XNOR U5666 ( .A(b[1]), .B(n5213), .Z(n5215) );
  NANDN U5667 ( .A(b[0]), .B(a[46]), .Z(n5214) );
  NAND U5668 ( .A(n5215), .B(n5214), .Z(n5287) );
  NAND U5669 ( .A(n583), .B(n5216), .Z(n5218) );
  XOR U5670 ( .A(b[29]), .B(a[19]), .Z(n5360) );
  NAND U5671 ( .A(n581), .B(n5360), .Z(n5217) );
  AND U5672 ( .A(n5218), .B(n5217), .Z(n5285) );
  AND U5673 ( .A(b[31]), .B(a[15]), .Z(n5284) );
  XNOR U5674 ( .A(n5285), .B(n5284), .Z(n5286) );
  XNOR U5675 ( .A(n5287), .B(n5286), .Z(n5327) );
  NAND U5676 ( .A(n578), .B(n5219), .Z(n5221) );
  XOR U5677 ( .A(b[23]), .B(a[25]), .Z(n5366) );
  NAND U5678 ( .A(n9268), .B(n5366), .Z(n5220) );
  AND U5679 ( .A(n5221), .B(n5220), .Z(n5356) );
  NAND U5680 ( .A(n569), .B(n5222), .Z(n5224) );
  XOR U5681 ( .A(b[7]), .B(a[41]), .Z(n5369) );
  NAND U5682 ( .A(n7819), .B(n5369), .Z(n5223) );
  AND U5683 ( .A(n5224), .B(n5223), .Z(n5355) );
  NAND U5684 ( .A(n579), .B(n5225), .Z(n5227) );
  XOR U5685 ( .A(b[25]), .B(a[23]), .Z(n5372) );
  NAND U5686 ( .A(n9364), .B(n5372), .Z(n5226) );
  NAND U5687 ( .A(n5227), .B(n5226), .Z(n5354) );
  XOR U5688 ( .A(n5355), .B(n5354), .Z(n5357) );
  XOR U5689 ( .A(n5356), .B(n5357), .Z(n5326) );
  XOR U5690 ( .A(n5327), .B(n5326), .Z(n5329) );
  NAND U5691 ( .A(n572), .B(n5228), .Z(n5230) );
  XOR U5692 ( .A(b[13]), .B(a[35]), .Z(n5375) );
  NAND U5693 ( .A(n8585), .B(n5375), .Z(n5229) );
  AND U5694 ( .A(n5230), .B(n5229), .Z(n5321) );
  NAND U5695 ( .A(n571), .B(n5231), .Z(n5233) );
  XOR U5696 ( .A(b[11]), .B(a[37]), .Z(n5378) );
  NAND U5697 ( .A(n8135), .B(n5378), .Z(n5232) );
  NAND U5698 ( .A(n5233), .B(n5232), .Z(n5320) );
  XNOR U5699 ( .A(n5321), .B(n5320), .Z(n5323) );
  NAND U5700 ( .A(n573), .B(n5234), .Z(n5236) );
  XOR U5701 ( .A(b[15]), .B(a[33]), .Z(n5381) );
  NAND U5702 ( .A(n8694), .B(n5381), .Z(n5235) );
  AND U5703 ( .A(n5236), .B(n5235), .Z(n5317) );
  NAND U5704 ( .A(n577), .B(n5237), .Z(n5239) );
  XOR U5705 ( .A(b[21]), .B(a[27]), .Z(n5384) );
  NAND U5706 ( .A(n9216), .B(n5384), .Z(n5238) );
  AND U5707 ( .A(n5239), .B(n5238), .Z(n5315) );
  NAND U5708 ( .A(n570), .B(n5240), .Z(n5242) );
  XOR U5709 ( .A(b[9]), .B(a[39]), .Z(n5387) );
  NAND U5710 ( .A(n8037), .B(n5387), .Z(n5241) );
  NAND U5711 ( .A(n5242), .B(n5241), .Z(n5314) );
  XNOR U5712 ( .A(n5315), .B(n5314), .Z(n5316) );
  XNOR U5713 ( .A(n5317), .B(n5316), .Z(n5322) );
  XOR U5714 ( .A(n5323), .B(n5322), .Z(n5328) );
  XNOR U5715 ( .A(n5329), .B(n5328), .Z(n5340) );
  XNOR U5716 ( .A(n5341), .B(n5340), .Z(n5396) );
  XNOR U5717 ( .A(n5397), .B(n5396), .Z(n5398) );
  XOR U5718 ( .A(n5399), .B(n5398), .Z(n5403) );
  XOR U5719 ( .A(n5402), .B(n5403), .Z(n5405) );
  XOR U5720 ( .A(n5404), .B(n5405), .Z(n5281) );
  NANDN U5721 ( .A(n5244), .B(n5243), .Z(n5248) );
  NAND U5722 ( .A(n5246), .B(n5245), .Z(n5247) );
  AND U5723 ( .A(n5248), .B(n5247), .Z(n5279) );
  NANDN U5724 ( .A(n5250), .B(n5249), .Z(n5254) );
  NANDN U5725 ( .A(n5252), .B(n5251), .Z(n5253) );
  AND U5726 ( .A(n5254), .B(n5253), .Z(n5278) );
  XNOR U5727 ( .A(n5279), .B(n5278), .Z(n5280) );
  XNOR U5728 ( .A(n5281), .B(n5280), .Z(n5272) );
  NANDN U5729 ( .A(n5256), .B(n5255), .Z(n5260) );
  NANDN U5730 ( .A(n5258), .B(n5257), .Z(n5259) );
  NAND U5731 ( .A(n5260), .B(n5259), .Z(n5273) );
  XOR U5732 ( .A(n5272), .B(n5273), .Z(n5275) );
  XNOR U5733 ( .A(n5274), .B(n5275), .Z(n5266) );
  XNOR U5734 ( .A(n5267), .B(n5266), .Z(n5268) );
  XNOR U5735 ( .A(n5269), .B(n5268), .Z(n5408) );
  XNOR U5736 ( .A(sreg[79]), .B(n5408), .Z(n5410) );
  NANDN U5737 ( .A(sreg[78]), .B(n5261), .Z(n5265) );
  NAND U5738 ( .A(n5263), .B(n5262), .Z(n5264) );
  NAND U5739 ( .A(n5265), .B(n5264), .Z(n5409) );
  XNOR U5740 ( .A(n5410), .B(n5409), .Z(c[79]) );
  NANDN U5741 ( .A(n5267), .B(n5266), .Z(n5271) );
  NANDN U5742 ( .A(n5269), .B(n5268), .Z(n5270) );
  AND U5743 ( .A(n5271), .B(n5270), .Z(n5416) );
  NANDN U5744 ( .A(n5273), .B(n5272), .Z(n5277) );
  NANDN U5745 ( .A(n5275), .B(n5274), .Z(n5276) );
  AND U5746 ( .A(n5277), .B(n5276), .Z(n5414) );
  NANDN U5747 ( .A(n5279), .B(n5278), .Z(n5283) );
  NANDN U5748 ( .A(n5281), .B(n5280), .Z(n5282) );
  AND U5749 ( .A(n5283), .B(n5282), .Z(n5422) );
  NANDN U5750 ( .A(n5285), .B(n5284), .Z(n5289) );
  NANDN U5751 ( .A(n5287), .B(n5286), .Z(n5288) );
  AND U5752 ( .A(n5289), .B(n5288), .Z(n5493) );
  NAND U5753 ( .A(n582), .B(n5290), .Z(n5292) );
  XOR U5754 ( .A(b[27]), .B(a[22]), .Z(n5437) );
  NAND U5755 ( .A(n9770), .B(n5437), .Z(n5291) );
  AND U5756 ( .A(n5292), .B(n5291), .Z(n5500) );
  NAND U5757 ( .A(n567), .B(n5293), .Z(n5295) );
  XOR U5758 ( .A(a[44]), .B(b[5]), .Z(n5440) );
  NAND U5759 ( .A(n7235), .B(n5440), .Z(n5294) );
  AND U5760 ( .A(n5295), .B(n5294), .Z(n5498) );
  NAND U5761 ( .A(n9046), .B(n5296), .Z(n5298) );
  XOR U5762 ( .A(b[19]), .B(a[30]), .Z(n5443) );
  NAND U5763 ( .A(n575), .B(n5443), .Z(n5297) );
  NAND U5764 ( .A(n5298), .B(n5297), .Z(n5497) );
  XNOR U5765 ( .A(n5498), .B(n5497), .Z(n5499) );
  XNOR U5766 ( .A(n5500), .B(n5499), .Z(n5491) );
  NAND U5767 ( .A(n9764), .B(n5299), .Z(n5301) );
  XOR U5768 ( .A(b[31]), .B(a[18]), .Z(n5446) );
  NAND U5769 ( .A(n584), .B(n5446), .Z(n5300) );
  AND U5770 ( .A(n5301), .B(n5300), .Z(n5458) );
  NAND U5771 ( .A(n568), .B(n5302), .Z(n5304) );
  XOR U5772 ( .A(a[46]), .B(b[3]), .Z(n5449) );
  NAND U5773 ( .A(n7245), .B(n5449), .Z(n5303) );
  AND U5774 ( .A(n5304), .B(n5303), .Z(n5456) );
  NAND U5775 ( .A(n576), .B(n5305), .Z(n5307) );
  XOR U5776 ( .A(b[17]), .B(a[32]), .Z(n5452) );
  NAND U5777 ( .A(n9141), .B(n5452), .Z(n5306) );
  NAND U5778 ( .A(n5307), .B(n5306), .Z(n5455) );
  XNOR U5779 ( .A(n5456), .B(n5455), .Z(n5457) );
  XOR U5780 ( .A(n5458), .B(n5457), .Z(n5492) );
  XOR U5781 ( .A(n5491), .B(n5492), .Z(n5494) );
  XOR U5782 ( .A(n5493), .B(n5494), .Z(n5540) );
  NANDN U5783 ( .A(n5309), .B(n5308), .Z(n5313) );
  NANDN U5784 ( .A(n5311), .B(n5310), .Z(n5312) );
  AND U5785 ( .A(n5313), .B(n5312), .Z(n5479) );
  NANDN U5786 ( .A(n5315), .B(n5314), .Z(n5319) );
  NANDN U5787 ( .A(n5317), .B(n5316), .Z(n5318) );
  NAND U5788 ( .A(n5319), .B(n5318), .Z(n5480) );
  XNOR U5789 ( .A(n5479), .B(n5480), .Z(n5481) );
  NANDN U5790 ( .A(n5321), .B(n5320), .Z(n5325) );
  NAND U5791 ( .A(n5323), .B(n5322), .Z(n5324) );
  NAND U5792 ( .A(n5325), .B(n5324), .Z(n5482) );
  XNOR U5793 ( .A(n5481), .B(n5482), .Z(n5539) );
  XNOR U5794 ( .A(n5540), .B(n5539), .Z(n5542) );
  NAND U5795 ( .A(n5327), .B(n5326), .Z(n5331) );
  NAND U5796 ( .A(n5329), .B(n5328), .Z(n5330) );
  AND U5797 ( .A(n5331), .B(n5330), .Z(n5541) );
  XOR U5798 ( .A(n5542), .B(n5541), .Z(n5553) );
  NANDN U5799 ( .A(n5333), .B(n5332), .Z(n5337) );
  NANDN U5800 ( .A(n5335), .B(n5334), .Z(n5336) );
  AND U5801 ( .A(n5337), .B(n5336), .Z(n5551) );
  NANDN U5802 ( .A(n5343), .B(n5342), .Z(n5347) );
  OR U5803 ( .A(n5345), .B(n5344), .Z(n5346) );
  AND U5804 ( .A(n5347), .B(n5346), .Z(n5546) );
  NANDN U5805 ( .A(n5349), .B(n5348), .Z(n5353) );
  NANDN U5806 ( .A(n5351), .B(n5350), .Z(n5352) );
  AND U5807 ( .A(n5353), .B(n5352), .Z(n5486) );
  NANDN U5808 ( .A(n5355), .B(n5354), .Z(n5359) );
  OR U5809 ( .A(n5357), .B(n5356), .Z(n5358) );
  NAND U5810 ( .A(n5359), .B(n5358), .Z(n5485) );
  XNOR U5811 ( .A(n5486), .B(n5485), .Z(n5487) );
  NAND U5812 ( .A(n583), .B(n5360), .Z(n5362) );
  XOR U5813 ( .A(b[29]), .B(a[20]), .Z(n5512) );
  NAND U5814 ( .A(n581), .B(n5512), .Z(n5361) );
  AND U5815 ( .A(n5362), .B(n5361), .Z(n5432) );
  AND U5816 ( .A(b[31]), .B(a[16]), .Z(n5431) );
  XNOR U5817 ( .A(n5432), .B(n5431), .Z(n5433) );
  NAND U5818 ( .A(b[0]), .B(a[48]), .Z(n5363) );
  XNOR U5819 ( .A(b[1]), .B(n5363), .Z(n5365) );
  NANDN U5820 ( .A(b[0]), .B(a[47]), .Z(n5364) );
  NAND U5821 ( .A(n5365), .B(n5364), .Z(n5434) );
  XNOR U5822 ( .A(n5433), .B(n5434), .Z(n5473) );
  NAND U5823 ( .A(n578), .B(n5366), .Z(n5368) );
  XOR U5824 ( .A(b[23]), .B(a[26]), .Z(n5515) );
  NAND U5825 ( .A(n9268), .B(n5515), .Z(n5367) );
  AND U5826 ( .A(n5368), .B(n5367), .Z(n5506) );
  NAND U5827 ( .A(n569), .B(n5369), .Z(n5371) );
  XOR U5828 ( .A(a[42]), .B(b[7]), .Z(n5518) );
  NAND U5829 ( .A(n7819), .B(n5518), .Z(n5370) );
  AND U5830 ( .A(n5371), .B(n5370), .Z(n5504) );
  NAND U5831 ( .A(n579), .B(n5372), .Z(n5374) );
  XOR U5832 ( .A(b[25]), .B(a[24]), .Z(n5521) );
  NAND U5833 ( .A(n9364), .B(n5521), .Z(n5373) );
  NAND U5834 ( .A(n5374), .B(n5373), .Z(n5503) );
  XNOR U5835 ( .A(n5504), .B(n5503), .Z(n5505) );
  XOR U5836 ( .A(n5506), .B(n5505), .Z(n5474) );
  XNOR U5837 ( .A(n5473), .B(n5474), .Z(n5475) );
  NAND U5838 ( .A(n572), .B(n5375), .Z(n5377) );
  XOR U5839 ( .A(b[13]), .B(a[36]), .Z(n5524) );
  NAND U5840 ( .A(n8585), .B(n5524), .Z(n5376) );
  AND U5841 ( .A(n5377), .B(n5376), .Z(n5468) );
  NAND U5842 ( .A(n571), .B(n5378), .Z(n5380) );
  XOR U5843 ( .A(b[11]), .B(a[38]), .Z(n5527) );
  NAND U5844 ( .A(n8135), .B(n5527), .Z(n5379) );
  NAND U5845 ( .A(n5380), .B(n5379), .Z(n5467) );
  XNOR U5846 ( .A(n5468), .B(n5467), .Z(n5469) );
  NAND U5847 ( .A(n573), .B(n5381), .Z(n5383) );
  XOR U5848 ( .A(b[15]), .B(a[34]), .Z(n5530) );
  NAND U5849 ( .A(n8694), .B(n5530), .Z(n5382) );
  AND U5850 ( .A(n5383), .B(n5382), .Z(n5464) );
  NAND U5851 ( .A(n577), .B(n5384), .Z(n5386) );
  XOR U5852 ( .A(b[21]), .B(a[28]), .Z(n5533) );
  NAND U5853 ( .A(n9216), .B(n5533), .Z(n5385) );
  AND U5854 ( .A(n5386), .B(n5385), .Z(n5462) );
  NAND U5855 ( .A(n570), .B(n5387), .Z(n5389) );
  XOR U5856 ( .A(b[9]), .B(a[40]), .Z(n5536) );
  NAND U5857 ( .A(n8037), .B(n5536), .Z(n5388) );
  NAND U5858 ( .A(n5389), .B(n5388), .Z(n5461) );
  XNOR U5859 ( .A(n5462), .B(n5461), .Z(n5463) );
  XOR U5860 ( .A(n5464), .B(n5463), .Z(n5470) );
  XOR U5861 ( .A(n5469), .B(n5470), .Z(n5476) );
  XOR U5862 ( .A(n5475), .B(n5476), .Z(n5488) );
  XNOR U5863 ( .A(n5487), .B(n5488), .Z(n5545) );
  XNOR U5864 ( .A(n5546), .B(n5545), .Z(n5547) );
  XOR U5865 ( .A(n5548), .B(n5547), .Z(n5552) );
  XOR U5866 ( .A(n5551), .B(n5552), .Z(n5554) );
  XOR U5867 ( .A(n5553), .B(n5554), .Z(n5428) );
  NANDN U5868 ( .A(n5391), .B(n5390), .Z(n5395) );
  NAND U5869 ( .A(n5393), .B(n5392), .Z(n5394) );
  AND U5870 ( .A(n5395), .B(n5394), .Z(n5426) );
  NANDN U5871 ( .A(n5397), .B(n5396), .Z(n5401) );
  NANDN U5872 ( .A(n5399), .B(n5398), .Z(n5400) );
  AND U5873 ( .A(n5401), .B(n5400), .Z(n5425) );
  XNOR U5874 ( .A(n5426), .B(n5425), .Z(n5427) );
  XNOR U5875 ( .A(n5428), .B(n5427), .Z(n5419) );
  NANDN U5876 ( .A(n5403), .B(n5402), .Z(n5407) );
  OR U5877 ( .A(n5405), .B(n5404), .Z(n5406) );
  NAND U5878 ( .A(n5407), .B(n5406), .Z(n5420) );
  XNOR U5879 ( .A(n5419), .B(n5420), .Z(n5421) );
  XNOR U5880 ( .A(n5422), .B(n5421), .Z(n5413) );
  XNOR U5881 ( .A(n5414), .B(n5413), .Z(n5415) );
  XNOR U5882 ( .A(n5416), .B(n5415), .Z(n5557) );
  XNOR U5883 ( .A(sreg[80]), .B(n5557), .Z(n5559) );
  NANDN U5884 ( .A(sreg[79]), .B(n5408), .Z(n5412) );
  NAND U5885 ( .A(n5410), .B(n5409), .Z(n5411) );
  NAND U5886 ( .A(n5412), .B(n5411), .Z(n5558) );
  XNOR U5887 ( .A(n5559), .B(n5558), .Z(c[80]) );
  NANDN U5888 ( .A(n5414), .B(n5413), .Z(n5418) );
  NANDN U5889 ( .A(n5416), .B(n5415), .Z(n5417) );
  AND U5890 ( .A(n5418), .B(n5417), .Z(n5565) );
  NANDN U5891 ( .A(n5420), .B(n5419), .Z(n5424) );
  NANDN U5892 ( .A(n5422), .B(n5421), .Z(n5423) );
  AND U5893 ( .A(n5424), .B(n5423), .Z(n5563) );
  NANDN U5894 ( .A(n5426), .B(n5425), .Z(n5430) );
  NANDN U5895 ( .A(n5428), .B(n5427), .Z(n5429) );
  AND U5896 ( .A(n5430), .B(n5429), .Z(n5571) );
  NANDN U5897 ( .A(n5432), .B(n5431), .Z(n5436) );
  NANDN U5898 ( .A(n5434), .B(n5433), .Z(n5435) );
  AND U5899 ( .A(n5436), .B(n5435), .Z(n5654) );
  NAND U5900 ( .A(n582), .B(n5437), .Z(n5439) );
  XOR U5901 ( .A(b[27]), .B(a[23]), .Z(n5598) );
  NAND U5902 ( .A(n9770), .B(n5598), .Z(n5438) );
  AND U5903 ( .A(n5439), .B(n5438), .Z(n5661) );
  NAND U5904 ( .A(n567), .B(n5440), .Z(n5442) );
  XOR U5905 ( .A(a[45]), .B(b[5]), .Z(n5601) );
  NAND U5906 ( .A(n7235), .B(n5601), .Z(n5441) );
  AND U5907 ( .A(n5442), .B(n5441), .Z(n5659) );
  NAND U5908 ( .A(n9046), .B(n5443), .Z(n5445) );
  XOR U5909 ( .A(b[19]), .B(a[31]), .Z(n5604) );
  NAND U5910 ( .A(n575), .B(n5604), .Z(n5444) );
  NAND U5911 ( .A(n5445), .B(n5444), .Z(n5658) );
  XNOR U5912 ( .A(n5659), .B(n5658), .Z(n5660) );
  XNOR U5913 ( .A(n5661), .B(n5660), .Z(n5652) );
  NAND U5914 ( .A(n9764), .B(n5446), .Z(n5448) );
  XOR U5915 ( .A(b[31]), .B(a[19]), .Z(n5607) );
  NAND U5916 ( .A(n584), .B(n5607), .Z(n5447) );
  AND U5917 ( .A(n5448), .B(n5447), .Z(n5619) );
  NAND U5918 ( .A(n568), .B(n5449), .Z(n5451) );
  XOR U5919 ( .A(a[47]), .B(b[3]), .Z(n5610) );
  NAND U5920 ( .A(n7245), .B(n5610), .Z(n5450) );
  AND U5921 ( .A(n5451), .B(n5450), .Z(n5617) );
  NAND U5922 ( .A(n576), .B(n5452), .Z(n5454) );
  XOR U5923 ( .A(b[17]), .B(a[33]), .Z(n5613) );
  NAND U5924 ( .A(n9141), .B(n5613), .Z(n5453) );
  NAND U5925 ( .A(n5454), .B(n5453), .Z(n5616) );
  XNOR U5926 ( .A(n5617), .B(n5616), .Z(n5618) );
  XOR U5927 ( .A(n5619), .B(n5618), .Z(n5653) );
  XOR U5928 ( .A(n5652), .B(n5653), .Z(n5655) );
  XOR U5929 ( .A(n5654), .B(n5655), .Z(n5587) );
  NANDN U5930 ( .A(n5456), .B(n5455), .Z(n5460) );
  NANDN U5931 ( .A(n5458), .B(n5457), .Z(n5459) );
  AND U5932 ( .A(n5460), .B(n5459), .Z(n5640) );
  NANDN U5933 ( .A(n5462), .B(n5461), .Z(n5466) );
  NANDN U5934 ( .A(n5464), .B(n5463), .Z(n5465) );
  NAND U5935 ( .A(n5466), .B(n5465), .Z(n5641) );
  XNOR U5936 ( .A(n5640), .B(n5641), .Z(n5642) );
  NANDN U5937 ( .A(n5468), .B(n5467), .Z(n5472) );
  NANDN U5938 ( .A(n5470), .B(n5469), .Z(n5471) );
  NAND U5939 ( .A(n5472), .B(n5471), .Z(n5643) );
  XNOR U5940 ( .A(n5642), .B(n5643), .Z(n5586) );
  XNOR U5941 ( .A(n5587), .B(n5586), .Z(n5589) );
  NANDN U5942 ( .A(n5474), .B(n5473), .Z(n5478) );
  NANDN U5943 ( .A(n5476), .B(n5475), .Z(n5477) );
  AND U5944 ( .A(n5478), .B(n5477), .Z(n5588) );
  XOR U5945 ( .A(n5589), .B(n5588), .Z(n5702) );
  NANDN U5946 ( .A(n5480), .B(n5479), .Z(n5484) );
  NANDN U5947 ( .A(n5482), .B(n5481), .Z(n5483) );
  AND U5948 ( .A(n5484), .B(n5483), .Z(n5700) );
  NANDN U5949 ( .A(n5486), .B(n5485), .Z(n5490) );
  NANDN U5950 ( .A(n5488), .B(n5487), .Z(n5489) );
  AND U5951 ( .A(n5490), .B(n5489), .Z(n5583) );
  NANDN U5952 ( .A(n5492), .B(n5491), .Z(n5496) );
  OR U5953 ( .A(n5494), .B(n5493), .Z(n5495) );
  AND U5954 ( .A(n5496), .B(n5495), .Z(n5581) );
  NANDN U5955 ( .A(n5498), .B(n5497), .Z(n5502) );
  NANDN U5956 ( .A(n5500), .B(n5499), .Z(n5501) );
  AND U5957 ( .A(n5502), .B(n5501), .Z(n5647) );
  NANDN U5958 ( .A(n5504), .B(n5503), .Z(n5508) );
  NANDN U5959 ( .A(n5506), .B(n5505), .Z(n5507) );
  NAND U5960 ( .A(n5508), .B(n5507), .Z(n5646) );
  XNOR U5961 ( .A(n5647), .B(n5646), .Z(n5648) );
  NAND U5962 ( .A(b[0]), .B(a[49]), .Z(n5509) );
  XNOR U5963 ( .A(b[1]), .B(n5509), .Z(n5511) );
  NANDN U5964 ( .A(b[0]), .B(a[48]), .Z(n5510) );
  NAND U5965 ( .A(n5511), .B(n5510), .Z(n5595) );
  NAND U5966 ( .A(n583), .B(n5512), .Z(n5514) );
  XOR U5967 ( .A(b[29]), .B(a[21]), .Z(n5673) );
  NAND U5968 ( .A(n581), .B(n5673), .Z(n5513) );
  AND U5969 ( .A(n5514), .B(n5513), .Z(n5593) );
  AND U5970 ( .A(b[31]), .B(a[17]), .Z(n5592) );
  XNOR U5971 ( .A(n5593), .B(n5592), .Z(n5594) );
  XNOR U5972 ( .A(n5595), .B(n5594), .Z(n5634) );
  NAND U5973 ( .A(n578), .B(n5515), .Z(n5517) );
  XOR U5974 ( .A(b[23]), .B(a[27]), .Z(n5676) );
  NAND U5975 ( .A(n9268), .B(n5676), .Z(n5516) );
  AND U5976 ( .A(n5517), .B(n5516), .Z(n5667) );
  NAND U5977 ( .A(n569), .B(n5518), .Z(n5520) );
  XOR U5978 ( .A(a[43]), .B(b[7]), .Z(n5679) );
  NAND U5979 ( .A(n7819), .B(n5679), .Z(n5519) );
  AND U5980 ( .A(n5520), .B(n5519), .Z(n5665) );
  NAND U5981 ( .A(n579), .B(n5521), .Z(n5523) );
  XOR U5982 ( .A(b[25]), .B(a[25]), .Z(n5682) );
  NAND U5983 ( .A(n9364), .B(n5682), .Z(n5522) );
  NAND U5984 ( .A(n5523), .B(n5522), .Z(n5664) );
  XNOR U5985 ( .A(n5665), .B(n5664), .Z(n5666) );
  XOR U5986 ( .A(n5667), .B(n5666), .Z(n5635) );
  XNOR U5987 ( .A(n5634), .B(n5635), .Z(n5636) );
  NAND U5988 ( .A(n572), .B(n5524), .Z(n5526) );
  XOR U5989 ( .A(b[13]), .B(a[37]), .Z(n5685) );
  NAND U5990 ( .A(n8585), .B(n5685), .Z(n5525) );
  AND U5991 ( .A(n5526), .B(n5525), .Z(n5629) );
  NAND U5992 ( .A(n571), .B(n5527), .Z(n5529) );
  XOR U5993 ( .A(b[11]), .B(a[39]), .Z(n5688) );
  NAND U5994 ( .A(n8135), .B(n5688), .Z(n5528) );
  NAND U5995 ( .A(n5529), .B(n5528), .Z(n5628) );
  XNOR U5996 ( .A(n5629), .B(n5628), .Z(n5630) );
  NAND U5997 ( .A(n573), .B(n5530), .Z(n5532) );
  XOR U5998 ( .A(b[15]), .B(a[35]), .Z(n5691) );
  NAND U5999 ( .A(n8694), .B(n5691), .Z(n5531) );
  AND U6000 ( .A(n5532), .B(n5531), .Z(n5625) );
  NAND U6001 ( .A(n577), .B(n5533), .Z(n5535) );
  XOR U6002 ( .A(b[21]), .B(a[29]), .Z(n5694) );
  NAND U6003 ( .A(n9216), .B(n5694), .Z(n5534) );
  AND U6004 ( .A(n5535), .B(n5534), .Z(n5623) );
  NAND U6005 ( .A(n570), .B(n5536), .Z(n5538) );
  XOR U6006 ( .A(b[9]), .B(a[41]), .Z(n5697) );
  NAND U6007 ( .A(n8037), .B(n5697), .Z(n5537) );
  NAND U6008 ( .A(n5538), .B(n5537), .Z(n5622) );
  XNOR U6009 ( .A(n5623), .B(n5622), .Z(n5624) );
  XOR U6010 ( .A(n5625), .B(n5624), .Z(n5631) );
  XOR U6011 ( .A(n5630), .B(n5631), .Z(n5637) );
  XOR U6012 ( .A(n5636), .B(n5637), .Z(n5649) );
  XNOR U6013 ( .A(n5648), .B(n5649), .Z(n5580) );
  XNOR U6014 ( .A(n5581), .B(n5580), .Z(n5582) );
  XOR U6015 ( .A(n5583), .B(n5582), .Z(n5701) );
  XOR U6016 ( .A(n5700), .B(n5701), .Z(n5703) );
  XOR U6017 ( .A(n5702), .B(n5703), .Z(n5577) );
  NANDN U6018 ( .A(n5540), .B(n5539), .Z(n5544) );
  NAND U6019 ( .A(n5542), .B(n5541), .Z(n5543) );
  AND U6020 ( .A(n5544), .B(n5543), .Z(n5575) );
  NANDN U6021 ( .A(n5546), .B(n5545), .Z(n5550) );
  NANDN U6022 ( .A(n5548), .B(n5547), .Z(n5549) );
  AND U6023 ( .A(n5550), .B(n5549), .Z(n5574) );
  XNOR U6024 ( .A(n5575), .B(n5574), .Z(n5576) );
  XNOR U6025 ( .A(n5577), .B(n5576), .Z(n5568) );
  NANDN U6026 ( .A(n5552), .B(n5551), .Z(n5556) );
  OR U6027 ( .A(n5554), .B(n5553), .Z(n5555) );
  NAND U6028 ( .A(n5556), .B(n5555), .Z(n5569) );
  XNOR U6029 ( .A(n5568), .B(n5569), .Z(n5570) );
  XNOR U6030 ( .A(n5571), .B(n5570), .Z(n5562) );
  XNOR U6031 ( .A(n5563), .B(n5562), .Z(n5564) );
  XNOR U6032 ( .A(n5565), .B(n5564), .Z(n5706) );
  XNOR U6033 ( .A(sreg[81]), .B(n5706), .Z(n5708) );
  NANDN U6034 ( .A(sreg[80]), .B(n5557), .Z(n5561) );
  NAND U6035 ( .A(n5559), .B(n5558), .Z(n5560) );
  NAND U6036 ( .A(n5561), .B(n5560), .Z(n5707) );
  XNOR U6037 ( .A(n5708), .B(n5707), .Z(c[81]) );
  NANDN U6038 ( .A(n5563), .B(n5562), .Z(n5567) );
  NANDN U6039 ( .A(n5565), .B(n5564), .Z(n5566) );
  AND U6040 ( .A(n5567), .B(n5566), .Z(n5714) );
  NANDN U6041 ( .A(n5569), .B(n5568), .Z(n5573) );
  NANDN U6042 ( .A(n5571), .B(n5570), .Z(n5572) );
  AND U6043 ( .A(n5573), .B(n5572), .Z(n5712) );
  NANDN U6044 ( .A(n5575), .B(n5574), .Z(n5579) );
  NANDN U6045 ( .A(n5577), .B(n5576), .Z(n5578) );
  AND U6046 ( .A(n5579), .B(n5578), .Z(n5720) );
  NANDN U6047 ( .A(n5581), .B(n5580), .Z(n5585) );
  NANDN U6048 ( .A(n5583), .B(n5582), .Z(n5584) );
  AND U6049 ( .A(n5585), .B(n5584), .Z(n5724) );
  NANDN U6050 ( .A(n5587), .B(n5586), .Z(n5591) );
  NAND U6051 ( .A(n5589), .B(n5588), .Z(n5590) );
  AND U6052 ( .A(n5591), .B(n5590), .Z(n5723) );
  XNOR U6053 ( .A(n5724), .B(n5723), .Z(n5726) );
  NANDN U6054 ( .A(n5593), .B(n5592), .Z(n5597) );
  NANDN U6055 ( .A(n5595), .B(n5594), .Z(n5596) );
  AND U6056 ( .A(n5597), .B(n5596), .Z(n5803) );
  NAND U6057 ( .A(n582), .B(n5598), .Z(n5600) );
  XOR U6058 ( .A(b[27]), .B(a[24]), .Z(n5747) );
  NAND U6059 ( .A(n9770), .B(n5747), .Z(n5599) );
  AND U6060 ( .A(n5600), .B(n5599), .Z(n5810) );
  NAND U6061 ( .A(n567), .B(n5601), .Z(n5603) );
  XOR U6062 ( .A(a[46]), .B(b[5]), .Z(n5750) );
  NAND U6063 ( .A(n7235), .B(n5750), .Z(n5602) );
  AND U6064 ( .A(n5603), .B(n5602), .Z(n5808) );
  NAND U6065 ( .A(n9046), .B(n5604), .Z(n5606) );
  XOR U6066 ( .A(b[19]), .B(a[32]), .Z(n5753) );
  NAND U6067 ( .A(n575), .B(n5753), .Z(n5605) );
  NAND U6068 ( .A(n5606), .B(n5605), .Z(n5807) );
  XNOR U6069 ( .A(n5808), .B(n5807), .Z(n5809) );
  XNOR U6070 ( .A(n5810), .B(n5809), .Z(n5801) );
  NAND U6071 ( .A(n9764), .B(n5607), .Z(n5609) );
  XOR U6072 ( .A(b[31]), .B(a[20]), .Z(n5756) );
  NAND U6073 ( .A(n584), .B(n5756), .Z(n5608) );
  AND U6074 ( .A(n5609), .B(n5608), .Z(n5768) );
  NAND U6075 ( .A(n568), .B(n5610), .Z(n5612) );
  XOR U6076 ( .A(a[48]), .B(b[3]), .Z(n5759) );
  NAND U6077 ( .A(n7245), .B(n5759), .Z(n5611) );
  AND U6078 ( .A(n5612), .B(n5611), .Z(n5766) );
  NAND U6079 ( .A(n576), .B(n5613), .Z(n5615) );
  XOR U6080 ( .A(b[17]), .B(a[34]), .Z(n5762) );
  NAND U6081 ( .A(n9141), .B(n5762), .Z(n5614) );
  NAND U6082 ( .A(n5615), .B(n5614), .Z(n5765) );
  XNOR U6083 ( .A(n5766), .B(n5765), .Z(n5767) );
  XOR U6084 ( .A(n5768), .B(n5767), .Z(n5802) );
  XOR U6085 ( .A(n5801), .B(n5802), .Z(n5804) );
  XOR U6086 ( .A(n5803), .B(n5804), .Z(n5736) );
  NANDN U6087 ( .A(n5617), .B(n5616), .Z(n5621) );
  NANDN U6088 ( .A(n5619), .B(n5618), .Z(n5620) );
  AND U6089 ( .A(n5621), .B(n5620), .Z(n5789) );
  NANDN U6090 ( .A(n5623), .B(n5622), .Z(n5627) );
  NANDN U6091 ( .A(n5625), .B(n5624), .Z(n5626) );
  NAND U6092 ( .A(n5627), .B(n5626), .Z(n5790) );
  XNOR U6093 ( .A(n5789), .B(n5790), .Z(n5791) );
  NANDN U6094 ( .A(n5629), .B(n5628), .Z(n5633) );
  NANDN U6095 ( .A(n5631), .B(n5630), .Z(n5632) );
  NAND U6096 ( .A(n5633), .B(n5632), .Z(n5792) );
  XNOR U6097 ( .A(n5791), .B(n5792), .Z(n5735) );
  XNOR U6098 ( .A(n5736), .B(n5735), .Z(n5738) );
  NANDN U6099 ( .A(n5635), .B(n5634), .Z(n5639) );
  NANDN U6100 ( .A(n5637), .B(n5636), .Z(n5638) );
  AND U6101 ( .A(n5639), .B(n5638), .Z(n5737) );
  XOR U6102 ( .A(n5738), .B(n5737), .Z(n5852) );
  NANDN U6103 ( .A(n5641), .B(n5640), .Z(n5645) );
  NANDN U6104 ( .A(n5643), .B(n5642), .Z(n5644) );
  AND U6105 ( .A(n5645), .B(n5644), .Z(n5849) );
  NANDN U6106 ( .A(n5647), .B(n5646), .Z(n5651) );
  NANDN U6107 ( .A(n5649), .B(n5648), .Z(n5650) );
  AND U6108 ( .A(n5651), .B(n5650), .Z(n5732) );
  NANDN U6109 ( .A(n5653), .B(n5652), .Z(n5657) );
  OR U6110 ( .A(n5655), .B(n5654), .Z(n5656) );
  AND U6111 ( .A(n5657), .B(n5656), .Z(n5730) );
  NANDN U6112 ( .A(n5659), .B(n5658), .Z(n5663) );
  NANDN U6113 ( .A(n5661), .B(n5660), .Z(n5662) );
  AND U6114 ( .A(n5663), .B(n5662), .Z(n5796) );
  NANDN U6115 ( .A(n5665), .B(n5664), .Z(n5669) );
  NANDN U6116 ( .A(n5667), .B(n5666), .Z(n5668) );
  NAND U6117 ( .A(n5669), .B(n5668), .Z(n5795) );
  XNOR U6118 ( .A(n5796), .B(n5795), .Z(n5797) );
  NAND U6119 ( .A(b[0]), .B(a[50]), .Z(n5670) );
  XNOR U6120 ( .A(b[1]), .B(n5670), .Z(n5672) );
  NANDN U6121 ( .A(b[0]), .B(a[49]), .Z(n5671) );
  NAND U6122 ( .A(n5672), .B(n5671), .Z(n5744) );
  NAND U6123 ( .A(n583), .B(n5673), .Z(n5675) );
  XOR U6124 ( .A(b[29]), .B(a[22]), .Z(n5819) );
  NAND U6125 ( .A(n581), .B(n5819), .Z(n5674) );
  AND U6126 ( .A(n5675), .B(n5674), .Z(n5742) );
  AND U6127 ( .A(b[31]), .B(a[18]), .Z(n5741) );
  XNOR U6128 ( .A(n5742), .B(n5741), .Z(n5743) );
  XNOR U6129 ( .A(n5744), .B(n5743), .Z(n5783) );
  NAND U6130 ( .A(n578), .B(n5676), .Z(n5678) );
  XOR U6131 ( .A(b[23]), .B(a[28]), .Z(n5825) );
  NAND U6132 ( .A(n9268), .B(n5825), .Z(n5677) );
  AND U6133 ( .A(n5678), .B(n5677), .Z(n5816) );
  NAND U6134 ( .A(n569), .B(n5679), .Z(n5681) );
  XOR U6135 ( .A(a[44]), .B(b[7]), .Z(n5828) );
  NAND U6136 ( .A(n7819), .B(n5828), .Z(n5680) );
  AND U6137 ( .A(n5681), .B(n5680), .Z(n5814) );
  NAND U6138 ( .A(n579), .B(n5682), .Z(n5684) );
  XOR U6139 ( .A(b[25]), .B(a[26]), .Z(n5831) );
  NAND U6140 ( .A(n9364), .B(n5831), .Z(n5683) );
  NAND U6141 ( .A(n5684), .B(n5683), .Z(n5813) );
  XNOR U6142 ( .A(n5814), .B(n5813), .Z(n5815) );
  XOR U6143 ( .A(n5816), .B(n5815), .Z(n5784) );
  XNOR U6144 ( .A(n5783), .B(n5784), .Z(n5785) );
  NAND U6145 ( .A(n572), .B(n5685), .Z(n5687) );
  XOR U6146 ( .A(b[13]), .B(a[38]), .Z(n5834) );
  NAND U6147 ( .A(n8585), .B(n5834), .Z(n5686) );
  AND U6148 ( .A(n5687), .B(n5686), .Z(n5778) );
  NAND U6149 ( .A(n571), .B(n5688), .Z(n5690) );
  XOR U6150 ( .A(b[11]), .B(a[40]), .Z(n5837) );
  NAND U6151 ( .A(n8135), .B(n5837), .Z(n5689) );
  NAND U6152 ( .A(n5690), .B(n5689), .Z(n5777) );
  XNOR U6153 ( .A(n5778), .B(n5777), .Z(n5779) );
  NAND U6154 ( .A(n573), .B(n5691), .Z(n5693) );
  XOR U6155 ( .A(b[15]), .B(a[36]), .Z(n5840) );
  NAND U6156 ( .A(n8694), .B(n5840), .Z(n5692) );
  AND U6157 ( .A(n5693), .B(n5692), .Z(n5774) );
  NAND U6158 ( .A(n577), .B(n5694), .Z(n5696) );
  XOR U6159 ( .A(b[21]), .B(a[30]), .Z(n5843) );
  NAND U6160 ( .A(n9216), .B(n5843), .Z(n5695) );
  AND U6161 ( .A(n5696), .B(n5695), .Z(n5772) );
  NAND U6162 ( .A(n570), .B(n5697), .Z(n5699) );
  XOR U6163 ( .A(b[9]), .B(a[42]), .Z(n5846) );
  NAND U6164 ( .A(n8037), .B(n5846), .Z(n5698) );
  NAND U6165 ( .A(n5699), .B(n5698), .Z(n5771) );
  XNOR U6166 ( .A(n5772), .B(n5771), .Z(n5773) );
  XOR U6167 ( .A(n5774), .B(n5773), .Z(n5780) );
  XOR U6168 ( .A(n5779), .B(n5780), .Z(n5786) );
  XOR U6169 ( .A(n5785), .B(n5786), .Z(n5798) );
  XNOR U6170 ( .A(n5797), .B(n5798), .Z(n5729) );
  XNOR U6171 ( .A(n5730), .B(n5729), .Z(n5731) );
  XOR U6172 ( .A(n5732), .B(n5731), .Z(n5850) );
  XNOR U6173 ( .A(n5849), .B(n5850), .Z(n5851) );
  XNOR U6174 ( .A(n5852), .B(n5851), .Z(n5725) );
  XOR U6175 ( .A(n5726), .B(n5725), .Z(n5718) );
  NANDN U6176 ( .A(n5701), .B(n5700), .Z(n5705) );
  OR U6177 ( .A(n5703), .B(n5702), .Z(n5704) );
  AND U6178 ( .A(n5705), .B(n5704), .Z(n5717) );
  XNOR U6179 ( .A(n5718), .B(n5717), .Z(n5719) );
  XNOR U6180 ( .A(n5720), .B(n5719), .Z(n5711) );
  XNOR U6181 ( .A(n5712), .B(n5711), .Z(n5713) );
  XNOR U6182 ( .A(n5714), .B(n5713), .Z(n5855) );
  XNOR U6183 ( .A(sreg[82]), .B(n5855), .Z(n5857) );
  NANDN U6184 ( .A(sreg[81]), .B(n5706), .Z(n5710) );
  NAND U6185 ( .A(n5708), .B(n5707), .Z(n5709) );
  NAND U6186 ( .A(n5710), .B(n5709), .Z(n5856) );
  XNOR U6187 ( .A(n5857), .B(n5856), .Z(c[82]) );
  NANDN U6188 ( .A(n5712), .B(n5711), .Z(n5716) );
  NANDN U6189 ( .A(n5714), .B(n5713), .Z(n5715) );
  AND U6190 ( .A(n5716), .B(n5715), .Z(n5863) );
  NANDN U6191 ( .A(n5718), .B(n5717), .Z(n5722) );
  NANDN U6192 ( .A(n5720), .B(n5719), .Z(n5721) );
  AND U6193 ( .A(n5722), .B(n5721), .Z(n5861) );
  NANDN U6194 ( .A(n5724), .B(n5723), .Z(n5728) );
  NAND U6195 ( .A(n5726), .B(n5725), .Z(n5727) );
  AND U6196 ( .A(n5728), .B(n5727), .Z(n5868) );
  NANDN U6197 ( .A(n5730), .B(n5729), .Z(n5734) );
  NANDN U6198 ( .A(n5732), .B(n5731), .Z(n5733) );
  AND U6199 ( .A(n5734), .B(n5733), .Z(n5873) );
  NANDN U6200 ( .A(n5736), .B(n5735), .Z(n5740) );
  NAND U6201 ( .A(n5738), .B(n5737), .Z(n5739) );
  AND U6202 ( .A(n5740), .B(n5739), .Z(n5872) );
  XNOR U6203 ( .A(n5873), .B(n5872), .Z(n5875) );
  NANDN U6204 ( .A(n5742), .B(n5741), .Z(n5746) );
  NANDN U6205 ( .A(n5744), .B(n5743), .Z(n5745) );
  AND U6206 ( .A(n5746), .B(n5745), .Z(n5950) );
  NAND U6207 ( .A(n582), .B(n5747), .Z(n5749) );
  XOR U6208 ( .A(b[27]), .B(a[25]), .Z(n5896) );
  NAND U6209 ( .A(n9770), .B(n5896), .Z(n5748) );
  AND U6210 ( .A(n5749), .B(n5748), .Z(n5957) );
  NAND U6211 ( .A(n567), .B(n5750), .Z(n5752) );
  XOR U6212 ( .A(a[47]), .B(b[5]), .Z(n5899) );
  NAND U6213 ( .A(n7235), .B(n5899), .Z(n5751) );
  AND U6214 ( .A(n5752), .B(n5751), .Z(n5955) );
  NAND U6215 ( .A(n9046), .B(n5753), .Z(n5755) );
  XOR U6216 ( .A(b[19]), .B(a[33]), .Z(n5902) );
  NAND U6217 ( .A(n575), .B(n5902), .Z(n5754) );
  NAND U6218 ( .A(n5755), .B(n5754), .Z(n5954) );
  XNOR U6219 ( .A(n5955), .B(n5954), .Z(n5956) );
  XNOR U6220 ( .A(n5957), .B(n5956), .Z(n5948) );
  NAND U6221 ( .A(n9764), .B(n5756), .Z(n5758) );
  XOR U6222 ( .A(b[31]), .B(a[21]), .Z(n5905) );
  NAND U6223 ( .A(n584), .B(n5905), .Z(n5757) );
  AND U6224 ( .A(n5758), .B(n5757), .Z(n5917) );
  NAND U6225 ( .A(n568), .B(n5759), .Z(n5761) );
  XOR U6226 ( .A(a[49]), .B(b[3]), .Z(n5908) );
  NAND U6227 ( .A(n7245), .B(n5908), .Z(n5760) );
  AND U6228 ( .A(n5761), .B(n5760), .Z(n5915) );
  NAND U6229 ( .A(n576), .B(n5762), .Z(n5764) );
  XOR U6230 ( .A(b[17]), .B(a[35]), .Z(n5911) );
  NAND U6231 ( .A(n9141), .B(n5911), .Z(n5763) );
  NAND U6232 ( .A(n5764), .B(n5763), .Z(n5914) );
  XNOR U6233 ( .A(n5915), .B(n5914), .Z(n5916) );
  XOR U6234 ( .A(n5917), .B(n5916), .Z(n5949) );
  XOR U6235 ( .A(n5948), .B(n5949), .Z(n5951) );
  XOR U6236 ( .A(n5950), .B(n5951), .Z(n5885) );
  NANDN U6237 ( .A(n5766), .B(n5765), .Z(n5770) );
  NANDN U6238 ( .A(n5768), .B(n5767), .Z(n5769) );
  AND U6239 ( .A(n5770), .B(n5769), .Z(n5938) );
  NANDN U6240 ( .A(n5772), .B(n5771), .Z(n5776) );
  NANDN U6241 ( .A(n5774), .B(n5773), .Z(n5775) );
  NAND U6242 ( .A(n5776), .B(n5775), .Z(n5939) );
  XNOR U6243 ( .A(n5938), .B(n5939), .Z(n5940) );
  NANDN U6244 ( .A(n5778), .B(n5777), .Z(n5782) );
  NANDN U6245 ( .A(n5780), .B(n5779), .Z(n5781) );
  NAND U6246 ( .A(n5782), .B(n5781), .Z(n5941) );
  XNOR U6247 ( .A(n5940), .B(n5941), .Z(n5884) );
  XNOR U6248 ( .A(n5885), .B(n5884), .Z(n5887) );
  NANDN U6249 ( .A(n5784), .B(n5783), .Z(n5788) );
  NANDN U6250 ( .A(n5786), .B(n5785), .Z(n5787) );
  AND U6251 ( .A(n5788), .B(n5787), .Z(n5886) );
  XOR U6252 ( .A(n5887), .B(n5886), .Z(n5999) );
  NANDN U6253 ( .A(n5790), .B(n5789), .Z(n5794) );
  NANDN U6254 ( .A(n5792), .B(n5791), .Z(n5793) );
  AND U6255 ( .A(n5794), .B(n5793), .Z(n5996) );
  NANDN U6256 ( .A(n5796), .B(n5795), .Z(n5800) );
  NANDN U6257 ( .A(n5798), .B(n5797), .Z(n5799) );
  AND U6258 ( .A(n5800), .B(n5799), .Z(n5881) );
  NANDN U6259 ( .A(n5802), .B(n5801), .Z(n5806) );
  OR U6260 ( .A(n5804), .B(n5803), .Z(n5805) );
  AND U6261 ( .A(n5806), .B(n5805), .Z(n5879) );
  NANDN U6262 ( .A(n5808), .B(n5807), .Z(n5812) );
  NANDN U6263 ( .A(n5810), .B(n5809), .Z(n5811) );
  AND U6264 ( .A(n5812), .B(n5811), .Z(n5945) );
  NANDN U6265 ( .A(n5814), .B(n5813), .Z(n5818) );
  NANDN U6266 ( .A(n5816), .B(n5815), .Z(n5817) );
  NAND U6267 ( .A(n5818), .B(n5817), .Z(n5944) );
  XNOR U6268 ( .A(n5945), .B(n5944), .Z(n5947) );
  NAND U6269 ( .A(n583), .B(n5819), .Z(n5821) );
  XOR U6270 ( .A(b[29]), .B(a[23]), .Z(n5969) );
  NAND U6271 ( .A(n581), .B(n5969), .Z(n5820) );
  AND U6272 ( .A(n5821), .B(n5820), .Z(n5891) );
  AND U6273 ( .A(b[31]), .B(a[19]), .Z(n5890) );
  XNOR U6274 ( .A(n5891), .B(n5890), .Z(n5892) );
  NAND U6275 ( .A(b[0]), .B(a[51]), .Z(n5822) );
  XNOR U6276 ( .A(b[1]), .B(n5822), .Z(n5824) );
  NANDN U6277 ( .A(b[0]), .B(a[50]), .Z(n5823) );
  NAND U6278 ( .A(n5824), .B(n5823), .Z(n5893) );
  XNOR U6279 ( .A(n5892), .B(n5893), .Z(n5933) );
  NAND U6280 ( .A(n578), .B(n5825), .Z(n5827) );
  XOR U6281 ( .A(b[23]), .B(a[29]), .Z(n5972) );
  NAND U6282 ( .A(n9268), .B(n5972), .Z(n5826) );
  AND U6283 ( .A(n5827), .B(n5826), .Z(n5962) );
  NAND U6284 ( .A(n569), .B(n5828), .Z(n5830) );
  XOR U6285 ( .A(a[45]), .B(b[7]), .Z(n5975) );
  NAND U6286 ( .A(n7819), .B(n5975), .Z(n5829) );
  AND U6287 ( .A(n5830), .B(n5829), .Z(n5961) );
  NAND U6288 ( .A(n579), .B(n5831), .Z(n5833) );
  XOR U6289 ( .A(b[25]), .B(a[27]), .Z(n5978) );
  NAND U6290 ( .A(n9364), .B(n5978), .Z(n5832) );
  NAND U6291 ( .A(n5833), .B(n5832), .Z(n5960) );
  XOR U6292 ( .A(n5961), .B(n5960), .Z(n5963) );
  XOR U6293 ( .A(n5962), .B(n5963), .Z(n5932) );
  XOR U6294 ( .A(n5933), .B(n5932), .Z(n5935) );
  NAND U6295 ( .A(n572), .B(n5834), .Z(n5836) );
  XOR U6296 ( .A(b[13]), .B(a[39]), .Z(n5981) );
  NAND U6297 ( .A(n8585), .B(n5981), .Z(n5835) );
  AND U6298 ( .A(n5836), .B(n5835), .Z(n5927) );
  NAND U6299 ( .A(n571), .B(n5837), .Z(n5839) );
  XOR U6300 ( .A(b[11]), .B(a[41]), .Z(n5984) );
  NAND U6301 ( .A(n8135), .B(n5984), .Z(n5838) );
  NAND U6302 ( .A(n5839), .B(n5838), .Z(n5926) );
  XNOR U6303 ( .A(n5927), .B(n5926), .Z(n5929) );
  NAND U6304 ( .A(n573), .B(n5840), .Z(n5842) );
  XOR U6305 ( .A(b[15]), .B(a[37]), .Z(n5987) );
  NAND U6306 ( .A(n8694), .B(n5987), .Z(n5841) );
  AND U6307 ( .A(n5842), .B(n5841), .Z(n5923) );
  NAND U6308 ( .A(n577), .B(n5843), .Z(n5845) );
  XOR U6309 ( .A(b[21]), .B(a[31]), .Z(n5990) );
  NAND U6310 ( .A(n9216), .B(n5990), .Z(n5844) );
  AND U6311 ( .A(n5845), .B(n5844), .Z(n5921) );
  NAND U6312 ( .A(n570), .B(n5846), .Z(n5848) );
  XOR U6313 ( .A(a[43]), .B(b[9]), .Z(n5993) );
  NAND U6314 ( .A(n8037), .B(n5993), .Z(n5847) );
  NAND U6315 ( .A(n5848), .B(n5847), .Z(n5920) );
  XNOR U6316 ( .A(n5921), .B(n5920), .Z(n5922) );
  XNOR U6317 ( .A(n5923), .B(n5922), .Z(n5928) );
  XOR U6318 ( .A(n5929), .B(n5928), .Z(n5934) );
  XNOR U6319 ( .A(n5935), .B(n5934), .Z(n5946) );
  XNOR U6320 ( .A(n5947), .B(n5946), .Z(n5878) );
  XNOR U6321 ( .A(n5879), .B(n5878), .Z(n5880) );
  XOR U6322 ( .A(n5881), .B(n5880), .Z(n5997) );
  XNOR U6323 ( .A(n5996), .B(n5997), .Z(n5998) );
  XNOR U6324 ( .A(n5999), .B(n5998), .Z(n5874) );
  XOR U6325 ( .A(n5875), .B(n5874), .Z(n5867) );
  NANDN U6326 ( .A(n5850), .B(n5849), .Z(n5854) );
  NANDN U6327 ( .A(n5852), .B(n5851), .Z(n5853) );
  AND U6328 ( .A(n5854), .B(n5853), .Z(n5866) );
  XOR U6329 ( .A(n5867), .B(n5866), .Z(n5869) );
  XNOR U6330 ( .A(n5868), .B(n5869), .Z(n5860) );
  XNOR U6331 ( .A(n5861), .B(n5860), .Z(n5862) );
  XNOR U6332 ( .A(n5863), .B(n5862), .Z(n6002) );
  XNOR U6333 ( .A(sreg[83]), .B(n6002), .Z(n6004) );
  NANDN U6334 ( .A(sreg[82]), .B(n5855), .Z(n5859) );
  NAND U6335 ( .A(n5857), .B(n5856), .Z(n5858) );
  NAND U6336 ( .A(n5859), .B(n5858), .Z(n6003) );
  XNOR U6337 ( .A(n6004), .B(n6003), .Z(c[83]) );
  NANDN U6338 ( .A(n5861), .B(n5860), .Z(n5865) );
  NANDN U6339 ( .A(n5863), .B(n5862), .Z(n5864) );
  AND U6340 ( .A(n5865), .B(n5864), .Z(n6010) );
  NANDN U6341 ( .A(n5867), .B(n5866), .Z(n5871) );
  NANDN U6342 ( .A(n5869), .B(n5868), .Z(n5870) );
  AND U6343 ( .A(n5871), .B(n5870), .Z(n6008) );
  NANDN U6344 ( .A(n5873), .B(n5872), .Z(n5877) );
  NAND U6345 ( .A(n5875), .B(n5874), .Z(n5876) );
  AND U6346 ( .A(n5877), .B(n5876), .Z(n6015) );
  NANDN U6347 ( .A(n5879), .B(n5878), .Z(n5883) );
  NANDN U6348 ( .A(n5881), .B(n5880), .Z(n5882) );
  AND U6349 ( .A(n5883), .B(n5882), .Z(n6144) );
  NANDN U6350 ( .A(n5885), .B(n5884), .Z(n5889) );
  NAND U6351 ( .A(n5887), .B(n5886), .Z(n5888) );
  AND U6352 ( .A(n5889), .B(n5888), .Z(n6143) );
  XNOR U6353 ( .A(n6144), .B(n6143), .Z(n6146) );
  NANDN U6354 ( .A(n5891), .B(n5890), .Z(n5895) );
  NANDN U6355 ( .A(n5893), .B(n5892), .Z(n5894) );
  AND U6356 ( .A(n5895), .B(n5894), .Z(n6079) );
  NAND U6357 ( .A(n582), .B(n5896), .Z(n5898) );
  XOR U6358 ( .A(b[27]), .B(a[26]), .Z(n6025) );
  NAND U6359 ( .A(n9770), .B(n6025), .Z(n5897) );
  AND U6360 ( .A(n5898), .B(n5897), .Z(n6086) );
  NAND U6361 ( .A(n567), .B(n5899), .Z(n5901) );
  XOR U6362 ( .A(a[48]), .B(b[5]), .Z(n6028) );
  NAND U6363 ( .A(n7235), .B(n6028), .Z(n5900) );
  AND U6364 ( .A(n5901), .B(n5900), .Z(n6084) );
  NAND U6365 ( .A(n9046), .B(n5902), .Z(n5904) );
  XOR U6366 ( .A(b[19]), .B(a[34]), .Z(n6031) );
  NAND U6367 ( .A(n575), .B(n6031), .Z(n5903) );
  NAND U6368 ( .A(n5904), .B(n5903), .Z(n6083) );
  XNOR U6369 ( .A(n6084), .B(n6083), .Z(n6085) );
  XNOR U6370 ( .A(n6086), .B(n6085), .Z(n6077) );
  NAND U6371 ( .A(n9764), .B(n5905), .Z(n5907) );
  XOR U6372 ( .A(b[31]), .B(a[22]), .Z(n6034) );
  NAND U6373 ( .A(n584), .B(n6034), .Z(n5906) );
  AND U6374 ( .A(n5907), .B(n5906), .Z(n6046) );
  NAND U6375 ( .A(n568), .B(n5908), .Z(n5910) );
  XOR U6376 ( .A(a[50]), .B(b[3]), .Z(n6037) );
  NAND U6377 ( .A(n7245), .B(n6037), .Z(n5909) );
  AND U6378 ( .A(n5910), .B(n5909), .Z(n6044) );
  NAND U6379 ( .A(n576), .B(n5911), .Z(n5913) );
  XOR U6380 ( .A(b[17]), .B(a[36]), .Z(n6040) );
  NAND U6381 ( .A(n9141), .B(n6040), .Z(n5912) );
  NAND U6382 ( .A(n5913), .B(n5912), .Z(n6043) );
  XNOR U6383 ( .A(n6044), .B(n6043), .Z(n6045) );
  XOR U6384 ( .A(n6046), .B(n6045), .Z(n6078) );
  XOR U6385 ( .A(n6077), .B(n6078), .Z(n6080) );
  XOR U6386 ( .A(n6079), .B(n6080), .Z(n6126) );
  NANDN U6387 ( .A(n5915), .B(n5914), .Z(n5919) );
  NANDN U6388 ( .A(n5917), .B(n5916), .Z(n5918) );
  AND U6389 ( .A(n5919), .B(n5918), .Z(n6067) );
  NANDN U6390 ( .A(n5921), .B(n5920), .Z(n5925) );
  NANDN U6391 ( .A(n5923), .B(n5922), .Z(n5924) );
  NAND U6392 ( .A(n5925), .B(n5924), .Z(n6068) );
  XNOR U6393 ( .A(n6067), .B(n6068), .Z(n6069) );
  NANDN U6394 ( .A(n5927), .B(n5926), .Z(n5931) );
  NAND U6395 ( .A(n5929), .B(n5928), .Z(n5930) );
  NAND U6396 ( .A(n5931), .B(n5930), .Z(n6070) );
  XNOR U6397 ( .A(n6069), .B(n6070), .Z(n6125) );
  XNOR U6398 ( .A(n6126), .B(n6125), .Z(n6128) );
  NAND U6399 ( .A(n5933), .B(n5932), .Z(n5937) );
  NAND U6400 ( .A(n5935), .B(n5934), .Z(n5936) );
  AND U6401 ( .A(n5937), .B(n5936), .Z(n6127) );
  XOR U6402 ( .A(n6128), .B(n6127), .Z(n6140) );
  NANDN U6403 ( .A(n5939), .B(n5938), .Z(n5943) );
  NANDN U6404 ( .A(n5941), .B(n5940), .Z(n5942) );
  AND U6405 ( .A(n5943), .B(n5942), .Z(n6137) );
  NANDN U6406 ( .A(n5949), .B(n5948), .Z(n5953) );
  OR U6407 ( .A(n5951), .B(n5950), .Z(n5952) );
  AND U6408 ( .A(n5953), .B(n5952), .Z(n6132) );
  NANDN U6409 ( .A(n5955), .B(n5954), .Z(n5959) );
  NANDN U6410 ( .A(n5957), .B(n5956), .Z(n5958) );
  AND U6411 ( .A(n5959), .B(n5958), .Z(n6074) );
  NANDN U6412 ( .A(n5961), .B(n5960), .Z(n5965) );
  OR U6413 ( .A(n5963), .B(n5962), .Z(n5964) );
  NAND U6414 ( .A(n5965), .B(n5964), .Z(n6073) );
  XNOR U6415 ( .A(n6074), .B(n6073), .Z(n6076) );
  NAND U6416 ( .A(b[0]), .B(a[52]), .Z(n5966) );
  XNOR U6417 ( .A(b[1]), .B(n5966), .Z(n5968) );
  NANDN U6418 ( .A(b[0]), .B(a[51]), .Z(n5967) );
  NAND U6419 ( .A(n5968), .B(n5967), .Z(n6022) );
  NAND U6420 ( .A(n583), .B(n5969), .Z(n5971) );
  XOR U6421 ( .A(b[29]), .B(a[24]), .Z(n6098) );
  NAND U6422 ( .A(n581), .B(n6098), .Z(n5970) );
  AND U6423 ( .A(n5971), .B(n5970), .Z(n6020) );
  AND U6424 ( .A(b[31]), .B(a[20]), .Z(n6019) );
  XNOR U6425 ( .A(n6020), .B(n6019), .Z(n6021) );
  XNOR U6426 ( .A(n6022), .B(n6021), .Z(n6062) );
  NAND U6427 ( .A(n578), .B(n5972), .Z(n5974) );
  XOR U6428 ( .A(b[23]), .B(a[30]), .Z(n6101) );
  NAND U6429 ( .A(n9268), .B(n6101), .Z(n5973) );
  AND U6430 ( .A(n5974), .B(n5973), .Z(n6091) );
  NAND U6431 ( .A(n569), .B(n5975), .Z(n5977) );
  XOR U6432 ( .A(a[46]), .B(b[7]), .Z(n6104) );
  NAND U6433 ( .A(n7819), .B(n6104), .Z(n5976) );
  AND U6434 ( .A(n5977), .B(n5976), .Z(n6090) );
  NAND U6435 ( .A(n579), .B(n5978), .Z(n5980) );
  XOR U6436 ( .A(b[25]), .B(a[28]), .Z(n6107) );
  NAND U6437 ( .A(n9364), .B(n6107), .Z(n5979) );
  NAND U6438 ( .A(n5980), .B(n5979), .Z(n6089) );
  XOR U6439 ( .A(n6090), .B(n6089), .Z(n6092) );
  XOR U6440 ( .A(n6091), .B(n6092), .Z(n6061) );
  XOR U6441 ( .A(n6062), .B(n6061), .Z(n6064) );
  NAND U6442 ( .A(n572), .B(n5981), .Z(n5983) );
  XOR U6443 ( .A(b[13]), .B(a[40]), .Z(n6110) );
  NAND U6444 ( .A(n8585), .B(n6110), .Z(n5982) );
  AND U6445 ( .A(n5983), .B(n5982), .Z(n6056) );
  NAND U6446 ( .A(n571), .B(n5984), .Z(n5986) );
  XOR U6447 ( .A(b[11]), .B(a[42]), .Z(n6113) );
  NAND U6448 ( .A(n8135), .B(n6113), .Z(n5985) );
  NAND U6449 ( .A(n5986), .B(n5985), .Z(n6055) );
  XNOR U6450 ( .A(n6056), .B(n6055), .Z(n6058) );
  NAND U6451 ( .A(n573), .B(n5987), .Z(n5989) );
  XOR U6452 ( .A(b[15]), .B(a[38]), .Z(n6116) );
  NAND U6453 ( .A(n8694), .B(n6116), .Z(n5988) );
  AND U6454 ( .A(n5989), .B(n5988), .Z(n6052) );
  NAND U6455 ( .A(n577), .B(n5990), .Z(n5992) );
  XOR U6456 ( .A(b[21]), .B(a[32]), .Z(n6119) );
  NAND U6457 ( .A(n9216), .B(n6119), .Z(n5991) );
  AND U6458 ( .A(n5992), .B(n5991), .Z(n6050) );
  NAND U6459 ( .A(n570), .B(n5993), .Z(n5995) );
  XOR U6460 ( .A(a[44]), .B(b[9]), .Z(n6122) );
  NAND U6461 ( .A(n8037), .B(n6122), .Z(n5994) );
  NAND U6462 ( .A(n5995), .B(n5994), .Z(n6049) );
  XNOR U6463 ( .A(n6050), .B(n6049), .Z(n6051) );
  XNOR U6464 ( .A(n6052), .B(n6051), .Z(n6057) );
  XOR U6465 ( .A(n6058), .B(n6057), .Z(n6063) );
  XNOR U6466 ( .A(n6064), .B(n6063), .Z(n6075) );
  XNOR U6467 ( .A(n6076), .B(n6075), .Z(n6131) );
  XNOR U6468 ( .A(n6132), .B(n6131), .Z(n6133) );
  XOR U6469 ( .A(n6134), .B(n6133), .Z(n6138) );
  XNOR U6470 ( .A(n6137), .B(n6138), .Z(n6139) );
  XNOR U6471 ( .A(n6140), .B(n6139), .Z(n6145) );
  XOR U6472 ( .A(n6146), .B(n6145), .Z(n6014) );
  NANDN U6473 ( .A(n5997), .B(n5996), .Z(n6001) );
  NANDN U6474 ( .A(n5999), .B(n5998), .Z(n6000) );
  AND U6475 ( .A(n6001), .B(n6000), .Z(n6013) );
  XOR U6476 ( .A(n6014), .B(n6013), .Z(n6016) );
  XNOR U6477 ( .A(n6015), .B(n6016), .Z(n6007) );
  XNOR U6478 ( .A(n6008), .B(n6007), .Z(n6009) );
  XNOR U6479 ( .A(n6010), .B(n6009), .Z(n6149) );
  XNOR U6480 ( .A(sreg[84]), .B(n6149), .Z(n6151) );
  NANDN U6481 ( .A(sreg[83]), .B(n6002), .Z(n6006) );
  NAND U6482 ( .A(n6004), .B(n6003), .Z(n6005) );
  NAND U6483 ( .A(n6006), .B(n6005), .Z(n6150) );
  XNOR U6484 ( .A(n6151), .B(n6150), .Z(c[84]) );
  NANDN U6485 ( .A(n6008), .B(n6007), .Z(n6012) );
  NANDN U6486 ( .A(n6010), .B(n6009), .Z(n6011) );
  AND U6487 ( .A(n6012), .B(n6011), .Z(n6157) );
  NANDN U6488 ( .A(n6014), .B(n6013), .Z(n6018) );
  NANDN U6489 ( .A(n6016), .B(n6015), .Z(n6017) );
  AND U6490 ( .A(n6018), .B(n6017), .Z(n6155) );
  NANDN U6491 ( .A(n6020), .B(n6019), .Z(n6024) );
  NANDN U6492 ( .A(n6022), .B(n6021), .Z(n6023) );
  AND U6493 ( .A(n6024), .B(n6023), .Z(n6234) );
  NAND U6494 ( .A(n582), .B(n6025), .Z(n6027) );
  XOR U6495 ( .A(b[27]), .B(a[27]), .Z(n6178) );
  NAND U6496 ( .A(n9770), .B(n6178), .Z(n6026) );
  AND U6497 ( .A(n6027), .B(n6026), .Z(n6241) );
  NAND U6498 ( .A(n567), .B(n6028), .Z(n6030) );
  XOR U6499 ( .A(a[49]), .B(b[5]), .Z(n6181) );
  NAND U6500 ( .A(n7235), .B(n6181), .Z(n6029) );
  AND U6501 ( .A(n6030), .B(n6029), .Z(n6239) );
  NAND U6502 ( .A(n9046), .B(n6031), .Z(n6033) );
  XOR U6503 ( .A(b[19]), .B(a[35]), .Z(n6184) );
  NAND U6504 ( .A(n575), .B(n6184), .Z(n6032) );
  NAND U6505 ( .A(n6033), .B(n6032), .Z(n6238) );
  XNOR U6506 ( .A(n6239), .B(n6238), .Z(n6240) );
  XNOR U6507 ( .A(n6241), .B(n6240), .Z(n6232) );
  NAND U6508 ( .A(n9764), .B(n6034), .Z(n6036) );
  XOR U6509 ( .A(b[31]), .B(a[23]), .Z(n6187) );
  NAND U6510 ( .A(n584), .B(n6187), .Z(n6035) );
  AND U6511 ( .A(n6036), .B(n6035), .Z(n6199) );
  NAND U6512 ( .A(n568), .B(n6037), .Z(n6039) );
  XOR U6513 ( .A(a[51]), .B(b[3]), .Z(n6190) );
  NAND U6514 ( .A(n7245), .B(n6190), .Z(n6038) );
  AND U6515 ( .A(n6039), .B(n6038), .Z(n6197) );
  NAND U6516 ( .A(n576), .B(n6040), .Z(n6042) );
  XOR U6517 ( .A(b[17]), .B(a[37]), .Z(n6193) );
  NAND U6518 ( .A(n9141), .B(n6193), .Z(n6041) );
  NAND U6519 ( .A(n6042), .B(n6041), .Z(n6196) );
  XNOR U6520 ( .A(n6197), .B(n6196), .Z(n6198) );
  XOR U6521 ( .A(n6199), .B(n6198), .Z(n6233) );
  XOR U6522 ( .A(n6232), .B(n6233), .Z(n6235) );
  XOR U6523 ( .A(n6234), .B(n6235), .Z(n6281) );
  NANDN U6524 ( .A(n6044), .B(n6043), .Z(n6048) );
  NANDN U6525 ( .A(n6046), .B(n6045), .Z(n6047) );
  AND U6526 ( .A(n6048), .B(n6047), .Z(n6220) );
  NANDN U6527 ( .A(n6050), .B(n6049), .Z(n6054) );
  NANDN U6528 ( .A(n6052), .B(n6051), .Z(n6053) );
  NAND U6529 ( .A(n6054), .B(n6053), .Z(n6221) );
  XNOR U6530 ( .A(n6220), .B(n6221), .Z(n6222) );
  NANDN U6531 ( .A(n6056), .B(n6055), .Z(n6060) );
  NAND U6532 ( .A(n6058), .B(n6057), .Z(n6059) );
  NAND U6533 ( .A(n6060), .B(n6059), .Z(n6223) );
  XNOR U6534 ( .A(n6222), .B(n6223), .Z(n6280) );
  XNOR U6535 ( .A(n6281), .B(n6280), .Z(n6283) );
  NAND U6536 ( .A(n6062), .B(n6061), .Z(n6066) );
  NAND U6537 ( .A(n6064), .B(n6063), .Z(n6065) );
  AND U6538 ( .A(n6066), .B(n6065), .Z(n6282) );
  XOR U6539 ( .A(n6283), .B(n6282), .Z(n6294) );
  NANDN U6540 ( .A(n6068), .B(n6067), .Z(n6072) );
  NANDN U6541 ( .A(n6070), .B(n6069), .Z(n6071) );
  AND U6542 ( .A(n6072), .B(n6071), .Z(n6292) );
  NANDN U6543 ( .A(n6078), .B(n6077), .Z(n6082) );
  OR U6544 ( .A(n6080), .B(n6079), .Z(n6081) );
  AND U6545 ( .A(n6082), .B(n6081), .Z(n6287) );
  NANDN U6546 ( .A(n6084), .B(n6083), .Z(n6088) );
  NANDN U6547 ( .A(n6086), .B(n6085), .Z(n6087) );
  AND U6548 ( .A(n6088), .B(n6087), .Z(n6227) );
  NANDN U6549 ( .A(n6090), .B(n6089), .Z(n6094) );
  OR U6550 ( .A(n6092), .B(n6091), .Z(n6093) );
  NAND U6551 ( .A(n6094), .B(n6093), .Z(n6226) );
  XNOR U6552 ( .A(n6227), .B(n6226), .Z(n6228) );
  NAND U6553 ( .A(b[0]), .B(a[53]), .Z(n6095) );
  XNOR U6554 ( .A(b[1]), .B(n6095), .Z(n6097) );
  NANDN U6555 ( .A(b[0]), .B(a[52]), .Z(n6096) );
  NAND U6556 ( .A(n6097), .B(n6096), .Z(n6175) );
  NAND U6557 ( .A(n583), .B(n6098), .Z(n6100) );
  XOR U6558 ( .A(b[29]), .B(a[25]), .Z(n6250) );
  NAND U6559 ( .A(n581), .B(n6250), .Z(n6099) );
  AND U6560 ( .A(n6100), .B(n6099), .Z(n6173) );
  AND U6561 ( .A(b[31]), .B(a[21]), .Z(n6172) );
  XNOR U6562 ( .A(n6173), .B(n6172), .Z(n6174) );
  XNOR U6563 ( .A(n6175), .B(n6174), .Z(n6214) );
  NAND U6564 ( .A(n578), .B(n6101), .Z(n6103) );
  XOR U6565 ( .A(b[23]), .B(a[31]), .Z(n6256) );
  NAND U6566 ( .A(n9268), .B(n6256), .Z(n6102) );
  AND U6567 ( .A(n6103), .B(n6102), .Z(n6247) );
  NAND U6568 ( .A(n569), .B(n6104), .Z(n6106) );
  XOR U6569 ( .A(a[47]), .B(b[7]), .Z(n6259) );
  NAND U6570 ( .A(n7819), .B(n6259), .Z(n6105) );
  AND U6571 ( .A(n6106), .B(n6105), .Z(n6245) );
  NAND U6572 ( .A(n579), .B(n6107), .Z(n6109) );
  XOR U6573 ( .A(b[25]), .B(a[29]), .Z(n6262) );
  NAND U6574 ( .A(n9364), .B(n6262), .Z(n6108) );
  NAND U6575 ( .A(n6109), .B(n6108), .Z(n6244) );
  XNOR U6576 ( .A(n6245), .B(n6244), .Z(n6246) );
  XOR U6577 ( .A(n6247), .B(n6246), .Z(n6215) );
  XNOR U6578 ( .A(n6214), .B(n6215), .Z(n6216) );
  NAND U6579 ( .A(n572), .B(n6110), .Z(n6112) );
  XOR U6580 ( .A(b[13]), .B(a[41]), .Z(n6265) );
  NAND U6581 ( .A(n8585), .B(n6265), .Z(n6111) );
  AND U6582 ( .A(n6112), .B(n6111), .Z(n6209) );
  NAND U6583 ( .A(n571), .B(n6113), .Z(n6115) );
  XOR U6584 ( .A(b[11]), .B(a[43]), .Z(n6268) );
  NAND U6585 ( .A(n8135), .B(n6268), .Z(n6114) );
  NAND U6586 ( .A(n6115), .B(n6114), .Z(n6208) );
  XNOR U6587 ( .A(n6209), .B(n6208), .Z(n6210) );
  NAND U6588 ( .A(n573), .B(n6116), .Z(n6118) );
  XOR U6589 ( .A(b[15]), .B(a[39]), .Z(n6271) );
  NAND U6590 ( .A(n8694), .B(n6271), .Z(n6117) );
  AND U6591 ( .A(n6118), .B(n6117), .Z(n6205) );
  NAND U6592 ( .A(n577), .B(n6119), .Z(n6121) );
  XOR U6593 ( .A(b[21]), .B(a[33]), .Z(n6274) );
  NAND U6594 ( .A(n9216), .B(n6274), .Z(n6120) );
  AND U6595 ( .A(n6121), .B(n6120), .Z(n6203) );
  NAND U6596 ( .A(n570), .B(n6122), .Z(n6124) );
  XOR U6597 ( .A(a[45]), .B(b[9]), .Z(n6277) );
  NAND U6598 ( .A(n8037), .B(n6277), .Z(n6123) );
  NAND U6599 ( .A(n6124), .B(n6123), .Z(n6202) );
  XNOR U6600 ( .A(n6203), .B(n6202), .Z(n6204) );
  XOR U6601 ( .A(n6205), .B(n6204), .Z(n6211) );
  XOR U6602 ( .A(n6210), .B(n6211), .Z(n6217) );
  XOR U6603 ( .A(n6216), .B(n6217), .Z(n6229) );
  XNOR U6604 ( .A(n6228), .B(n6229), .Z(n6286) );
  XNOR U6605 ( .A(n6287), .B(n6286), .Z(n6288) );
  XOR U6606 ( .A(n6289), .B(n6288), .Z(n6293) );
  XOR U6607 ( .A(n6292), .B(n6293), .Z(n6295) );
  XOR U6608 ( .A(n6294), .B(n6295), .Z(n6169) );
  NANDN U6609 ( .A(n6126), .B(n6125), .Z(n6130) );
  NAND U6610 ( .A(n6128), .B(n6127), .Z(n6129) );
  AND U6611 ( .A(n6130), .B(n6129), .Z(n6167) );
  NANDN U6612 ( .A(n6132), .B(n6131), .Z(n6136) );
  NANDN U6613 ( .A(n6134), .B(n6133), .Z(n6135) );
  AND U6614 ( .A(n6136), .B(n6135), .Z(n6166) );
  XNOR U6615 ( .A(n6167), .B(n6166), .Z(n6168) );
  XNOR U6616 ( .A(n6169), .B(n6168), .Z(n6160) );
  NANDN U6617 ( .A(n6138), .B(n6137), .Z(n6142) );
  NANDN U6618 ( .A(n6140), .B(n6139), .Z(n6141) );
  NAND U6619 ( .A(n6142), .B(n6141), .Z(n6161) );
  XNOR U6620 ( .A(n6160), .B(n6161), .Z(n6162) );
  NANDN U6621 ( .A(n6144), .B(n6143), .Z(n6148) );
  NAND U6622 ( .A(n6146), .B(n6145), .Z(n6147) );
  NAND U6623 ( .A(n6148), .B(n6147), .Z(n6163) );
  XNOR U6624 ( .A(n6162), .B(n6163), .Z(n6154) );
  XNOR U6625 ( .A(n6155), .B(n6154), .Z(n6156) );
  XNOR U6626 ( .A(n6157), .B(n6156), .Z(n6298) );
  XNOR U6627 ( .A(sreg[85]), .B(n6298), .Z(n6300) );
  NANDN U6628 ( .A(sreg[84]), .B(n6149), .Z(n6153) );
  NAND U6629 ( .A(n6151), .B(n6150), .Z(n6152) );
  NAND U6630 ( .A(n6153), .B(n6152), .Z(n6299) );
  XNOR U6631 ( .A(n6300), .B(n6299), .Z(c[85]) );
  NANDN U6632 ( .A(n6155), .B(n6154), .Z(n6159) );
  NANDN U6633 ( .A(n6157), .B(n6156), .Z(n6158) );
  AND U6634 ( .A(n6159), .B(n6158), .Z(n6306) );
  NANDN U6635 ( .A(n6161), .B(n6160), .Z(n6165) );
  NANDN U6636 ( .A(n6163), .B(n6162), .Z(n6164) );
  AND U6637 ( .A(n6165), .B(n6164), .Z(n6304) );
  NANDN U6638 ( .A(n6167), .B(n6166), .Z(n6171) );
  NANDN U6639 ( .A(n6169), .B(n6168), .Z(n6170) );
  AND U6640 ( .A(n6171), .B(n6170), .Z(n6312) );
  NANDN U6641 ( .A(n6173), .B(n6172), .Z(n6177) );
  NANDN U6642 ( .A(n6175), .B(n6174), .Z(n6176) );
  AND U6643 ( .A(n6177), .B(n6176), .Z(n6393) );
  NAND U6644 ( .A(n582), .B(n6178), .Z(n6180) );
  XOR U6645 ( .A(b[27]), .B(a[28]), .Z(n6339) );
  NAND U6646 ( .A(n9770), .B(n6339), .Z(n6179) );
  AND U6647 ( .A(n6180), .B(n6179), .Z(n6400) );
  NAND U6648 ( .A(n567), .B(n6181), .Z(n6183) );
  XOR U6649 ( .A(a[50]), .B(b[5]), .Z(n6342) );
  NAND U6650 ( .A(n7235), .B(n6342), .Z(n6182) );
  AND U6651 ( .A(n6183), .B(n6182), .Z(n6398) );
  NAND U6652 ( .A(n9046), .B(n6184), .Z(n6186) );
  XOR U6653 ( .A(b[19]), .B(a[36]), .Z(n6345) );
  NAND U6654 ( .A(n575), .B(n6345), .Z(n6185) );
  NAND U6655 ( .A(n6186), .B(n6185), .Z(n6397) );
  XNOR U6656 ( .A(n6398), .B(n6397), .Z(n6399) );
  XNOR U6657 ( .A(n6400), .B(n6399), .Z(n6391) );
  NAND U6658 ( .A(n9764), .B(n6187), .Z(n6189) );
  XOR U6659 ( .A(b[31]), .B(a[24]), .Z(n6348) );
  NAND U6660 ( .A(n584), .B(n6348), .Z(n6188) );
  AND U6661 ( .A(n6189), .B(n6188), .Z(n6360) );
  NAND U6662 ( .A(n568), .B(n6190), .Z(n6192) );
  XOR U6663 ( .A(a[52]), .B(b[3]), .Z(n6351) );
  NAND U6664 ( .A(n7245), .B(n6351), .Z(n6191) );
  AND U6665 ( .A(n6192), .B(n6191), .Z(n6358) );
  NAND U6666 ( .A(n576), .B(n6193), .Z(n6195) );
  XOR U6667 ( .A(b[17]), .B(a[38]), .Z(n6354) );
  NAND U6668 ( .A(n9141), .B(n6354), .Z(n6194) );
  NAND U6669 ( .A(n6195), .B(n6194), .Z(n6357) );
  XNOR U6670 ( .A(n6358), .B(n6357), .Z(n6359) );
  XOR U6671 ( .A(n6360), .B(n6359), .Z(n6392) );
  XOR U6672 ( .A(n6391), .B(n6392), .Z(n6394) );
  XOR U6673 ( .A(n6393), .B(n6394), .Z(n6328) );
  NANDN U6674 ( .A(n6197), .B(n6196), .Z(n6201) );
  NANDN U6675 ( .A(n6199), .B(n6198), .Z(n6200) );
  AND U6676 ( .A(n6201), .B(n6200), .Z(n6381) );
  NANDN U6677 ( .A(n6203), .B(n6202), .Z(n6207) );
  NANDN U6678 ( .A(n6205), .B(n6204), .Z(n6206) );
  NAND U6679 ( .A(n6207), .B(n6206), .Z(n6382) );
  XNOR U6680 ( .A(n6381), .B(n6382), .Z(n6383) );
  NANDN U6681 ( .A(n6209), .B(n6208), .Z(n6213) );
  NANDN U6682 ( .A(n6211), .B(n6210), .Z(n6212) );
  NAND U6683 ( .A(n6213), .B(n6212), .Z(n6384) );
  XNOR U6684 ( .A(n6383), .B(n6384), .Z(n6327) );
  XNOR U6685 ( .A(n6328), .B(n6327), .Z(n6330) );
  NANDN U6686 ( .A(n6215), .B(n6214), .Z(n6219) );
  NANDN U6687 ( .A(n6217), .B(n6216), .Z(n6218) );
  AND U6688 ( .A(n6219), .B(n6218), .Z(n6329) );
  XOR U6689 ( .A(n6330), .B(n6329), .Z(n6441) );
  NANDN U6690 ( .A(n6221), .B(n6220), .Z(n6225) );
  NANDN U6691 ( .A(n6223), .B(n6222), .Z(n6224) );
  AND U6692 ( .A(n6225), .B(n6224), .Z(n6439) );
  NANDN U6693 ( .A(n6227), .B(n6226), .Z(n6231) );
  NANDN U6694 ( .A(n6229), .B(n6228), .Z(n6230) );
  AND U6695 ( .A(n6231), .B(n6230), .Z(n6324) );
  NANDN U6696 ( .A(n6233), .B(n6232), .Z(n6237) );
  OR U6697 ( .A(n6235), .B(n6234), .Z(n6236) );
  AND U6698 ( .A(n6237), .B(n6236), .Z(n6322) );
  NANDN U6699 ( .A(n6239), .B(n6238), .Z(n6243) );
  NANDN U6700 ( .A(n6241), .B(n6240), .Z(n6242) );
  AND U6701 ( .A(n6243), .B(n6242), .Z(n6388) );
  NANDN U6702 ( .A(n6245), .B(n6244), .Z(n6249) );
  NANDN U6703 ( .A(n6247), .B(n6246), .Z(n6248) );
  NAND U6704 ( .A(n6249), .B(n6248), .Z(n6387) );
  XNOR U6705 ( .A(n6388), .B(n6387), .Z(n6390) );
  NAND U6706 ( .A(n583), .B(n6250), .Z(n6252) );
  XOR U6707 ( .A(b[29]), .B(a[26]), .Z(n6409) );
  NAND U6708 ( .A(n581), .B(n6409), .Z(n6251) );
  AND U6709 ( .A(n6252), .B(n6251), .Z(n6334) );
  AND U6710 ( .A(b[31]), .B(a[22]), .Z(n6333) );
  XNOR U6711 ( .A(n6334), .B(n6333), .Z(n6335) );
  NAND U6712 ( .A(b[0]), .B(a[54]), .Z(n6253) );
  XNOR U6713 ( .A(b[1]), .B(n6253), .Z(n6255) );
  NANDN U6714 ( .A(b[0]), .B(a[53]), .Z(n6254) );
  NAND U6715 ( .A(n6255), .B(n6254), .Z(n6336) );
  XNOR U6716 ( .A(n6335), .B(n6336), .Z(n6376) );
  NAND U6717 ( .A(n578), .B(n6256), .Z(n6258) );
  XOR U6718 ( .A(b[23]), .B(a[32]), .Z(n6415) );
  NAND U6719 ( .A(n9268), .B(n6415), .Z(n6257) );
  AND U6720 ( .A(n6258), .B(n6257), .Z(n6405) );
  NAND U6721 ( .A(n569), .B(n6259), .Z(n6261) );
  XOR U6722 ( .A(a[48]), .B(b[7]), .Z(n6418) );
  NAND U6723 ( .A(n7819), .B(n6418), .Z(n6260) );
  AND U6724 ( .A(n6261), .B(n6260), .Z(n6404) );
  NAND U6725 ( .A(n579), .B(n6262), .Z(n6264) );
  XOR U6726 ( .A(b[25]), .B(a[30]), .Z(n6421) );
  NAND U6727 ( .A(n9364), .B(n6421), .Z(n6263) );
  NAND U6728 ( .A(n6264), .B(n6263), .Z(n6403) );
  XOR U6729 ( .A(n6404), .B(n6403), .Z(n6406) );
  XOR U6730 ( .A(n6405), .B(n6406), .Z(n6375) );
  XOR U6731 ( .A(n6376), .B(n6375), .Z(n6378) );
  NAND U6732 ( .A(n572), .B(n6265), .Z(n6267) );
  XOR U6733 ( .A(b[13]), .B(a[42]), .Z(n6424) );
  NAND U6734 ( .A(n8585), .B(n6424), .Z(n6266) );
  AND U6735 ( .A(n6267), .B(n6266), .Z(n6370) );
  NAND U6736 ( .A(n571), .B(n6268), .Z(n6270) );
  XOR U6737 ( .A(b[11]), .B(a[44]), .Z(n6427) );
  NAND U6738 ( .A(n8135), .B(n6427), .Z(n6269) );
  NAND U6739 ( .A(n6270), .B(n6269), .Z(n6369) );
  XNOR U6740 ( .A(n6370), .B(n6369), .Z(n6372) );
  NAND U6741 ( .A(n573), .B(n6271), .Z(n6273) );
  XOR U6742 ( .A(b[15]), .B(a[40]), .Z(n6430) );
  NAND U6743 ( .A(n8694), .B(n6430), .Z(n6272) );
  AND U6744 ( .A(n6273), .B(n6272), .Z(n6366) );
  NAND U6745 ( .A(n577), .B(n6274), .Z(n6276) );
  XOR U6746 ( .A(b[21]), .B(a[34]), .Z(n6433) );
  NAND U6747 ( .A(n9216), .B(n6433), .Z(n6275) );
  AND U6748 ( .A(n6276), .B(n6275), .Z(n6364) );
  NAND U6749 ( .A(n570), .B(n6277), .Z(n6279) );
  XOR U6750 ( .A(a[46]), .B(b[9]), .Z(n6436) );
  NAND U6751 ( .A(n8037), .B(n6436), .Z(n6278) );
  NAND U6752 ( .A(n6279), .B(n6278), .Z(n6363) );
  XNOR U6753 ( .A(n6364), .B(n6363), .Z(n6365) );
  XNOR U6754 ( .A(n6366), .B(n6365), .Z(n6371) );
  XOR U6755 ( .A(n6372), .B(n6371), .Z(n6377) );
  XNOR U6756 ( .A(n6378), .B(n6377), .Z(n6389) );
  XNOR U6757 ( .A(n6390), .B(n6389), .Z(n6321) );
  XNOR U6758 ( .A(n6322), .B(n6321), .Z(n6323) );
  XOR U6759 ( .A(n6324), .B(n6323), .Z(n6440) );
  XOR U6760 ( .A(n6439), .B(n6440), .Z(n6442) );
  XOR U6761 ( .A(n6441), .B(n6442), .Z(n6318) );
  NANDN U6762 ( .A(n6281), .B(n6280), .Z(n6285) );
  NAND U6763 ( .A(n6283), .B(n6282), .Z(n6284) );
  AND U6764 ( .A(n6285), .B(n6284), .Z(n6316) );
  NANDN U6765 ( .A(n6287), .B(n6286), .Z(n6291) );
  NANDN U6766 ( .A(n6289), .B(n6288), .Z(n6290) );
  AND U6767 ( .A(n6291), .B(n6290), .Z(n6315) );
  XNOR U6768 ( .A(n6316), .B(n6315), .Z(n6317) );
  XNOR U6769 ( .A(n6318), .B(n6317), .Z(n6309) );
  NANDN U6770 ( .A(n6293), .B(n6292), .Z(n6297) );
  OR U6771 ( .A(n6295), .B(n6294), .Z(n6296) );
  NAND U6772 ( .A(n6297), .B(n6296), .Z(n6310) );
  XNOR U6773 ( .A(n6309), .B(n6310), .Z(n6311) );
  XNOR U6774 ( .A(n6312), .B(n6311), .Z(n6303) );
  XNOR U6775 ( .A(n6304), .B(n6303), .Z(n6305) );
  XNOR U6776 ( .A(n6306), .B(n6305), .Z(n6445) );
  XNOR U6777 ( .A(sreg[86]), .B(n6445), .Z(n6447) );
  NANDN U6778 ( .A(sreg[85]), .B(n6298), .Z(n6302) );
  NAND U6779 ( .A(n6300), .B(n6299), .Z(n6301) );
  NAND U6780 ( .A(n6302), .B(n6301), .Z(n6446) );
  XNOR U6781 ( .A(n6447), .B(n6446), .Z(c[86]) );
  NANDN U6782 ( .A(n6304), .B(n6303), .Z(n6308) );
  NANDN U6783 ( .A(n6306), .B(n6305), .Z(n6307) );
  AND U6784 ( .A(n6308), .B(n6307), .Z(n6453) );
  NANDN U6785 ( .A(n6310), .B(n6309), .Z(n6314) );
  NANDN U6786 ( .A(n6312), .B(n6311), .Z(n6313) );
  AND U6787 ( .A(n6314), .B(n6313), .Z(n6451) );
  NANDN U6788 ( .A(n6316), .B(n6315), .Z(n6320) );
  NANDN U6789 ( .A(n6318), .B(n6317), .Z(n6319) );
  AND U6790 ( .A(n6320), .B(n6319), .Z(n6459) );
  NANDN U6791 ( .A(n6322), .B(n6321), .Z(n6326) );
  NANDN U6792 ( .A(n6324), .B(n6323), .Z(n6325) );
  AND U6793 ( .A(n6326), .B(n6325), .Z(n6463) );
  NANDN U6794 ( .A(n6328), .B(n6327), .Z(n6332) );
  NAND U6795 ( .A(n6330), .B(n6329), .Z(n6331) );
  AND U6796 ( .A(n6332), .B(n6331), .Z(n6462) );
  XNOR U6797 ( .A(n6463), .B(n6462), .Z(n6465) );
  NANDN U6798 ( .A(n6334), .B(n6333), .Z(n6338) );
  NANDN U6799 ( .A(n6336), .B(n6335), .Z(n6337) );
  AND U6800 ( .A(n6338), .B(n6337), .Z(n6530) );
  NAND U6801 ( .A(n582), .B(n6339), .Z(n6341) );
  XOR U6802 ( .A(b[27]), .B(a[29]), .Z(n6474) );
  NAND U6803 ( .A(n9770), .B(n6474), .Z(n6340) );
  AND U6804 ( .A(n6341), .B(n6340), .Z(n6537) );
  NAND U6805 ( .A(n567), .B(n6342), .Z(n6344) );
  XOR U6806 ( .A(a[51]), .B(b[5]), .Z(n6477) );
  NAND U6807 ( .A(n7235), .B(n6477), .Z(n6343) );
  AND U6808 ( .A(n6344), .B(n6343), .Z(n6535) );
  NAND U6809 ( .A(n9046), .B(n6345), .Z(n6347) );
  XOR U6810 ( .A(b[19]), .B(a[37]), .Z(n6480) );
  NAND U6811 ( .A(n575), .B(n6480), .Z(n6346) );
  NAND U6812 ( .A(n6347), .B(n6346), .Z(n6534) );
  XNOR U6813 ( .A(n6535), .B(n6534), .Z(n6536) );
  XNOR U6814 ( .A(n6537), .B(n6536), .Z(n6528) );
  NAND U6815 ( .A(n9764), .B(n6348), .Z(n6350) );
  XOR U6816 ( .A(b[31]), .B(a[25]), .Z(n6483) );
  NAND U6817 ( .A(n584), .B(n6483), .Z(n6349) );
  AND U6818 ( .A(n6350), .B(n6349), .Z(n6495) );
  NAND U6819 ( .A(n568), .B(n6351), .Z(n6353) );
  XOR U6820 ( .A(a[53]), .B(b[3]), .Z(n6486) );
  NAND U6821 ( .A(n7245), .B(n6486), .Z(n6352) );
  AND U6822 ( .A(n6353), .B(n6352), .Z(n6493) );
  NAND U6823 ( .A(n576), .B(n6354), .Z(n6356) );
  XOR U6824 ( .A(b[17]), .B(a[39]), .Z(n6489) );
  NAND U6825 ( .A(n9141), .B(n6489), .Z(n6355) );
  NAND U6826 ( .A(n6356), .B(n6355), .Z(n6492) );
  XNOR U6827 ( .A(n6493), .B(n6492), .Z(n6494) );
  XOR U6828 ( .A(n6495), .B(n6494), .Z(n6529) );
  XOR U6829 ( .A(n6528), .B(n6529), .Z(n6531) );
  XOR U6830 ( .A(n6530), .B(n6531), .Z(n6577) );
  NANDN U6831 ( .A(n6358), .B(n6357), .Z(n6362) );
  NANDN U6832 ( .A(n6360), .B(n6359), .Z(n6361) );
  AND U6833 ( .A(n6362), .B(n6361), .Z(n6516) );
  NANDN U6834 ( .A(n6364), .B(n6363), .Z(n6368) );
  NANDN U6835 ( .A(n6366), .B(n6365), .Z(n6367) );
  NAND U6836 ( .A(n6368), .B(n6367), .Z(n6517) );
  XNOR U6837 ( .A(n6516), .B(n6517), .Z(n6518) );
  NANDN U6838 ( .A(n6370), .B(n6369), .Z(n6374) );
  NAND U6839 ( .A(n6372), .B(n6371), .Z(n6373) );
  NAND U6840 ( .A(n6374), .B(n6373), .Z(n6519) );
  XNOR U6841 ( .A(n6518), .B(n6519), .Z(n6576) );
  XNOR U6842 ( .A(n6577), .B(n6576), .Z(n6579) );
  NAND U6843 ( .A(n6376), .B(n6375), .Z(n6380) );
  NAND U6844 ( .A(n6378), .B(n6377), .Z(n6379) );
  AND U6845 ( .A(n6380), .B(n6379), .Z(n6578) );
  XOR U6846 ( .A(n6579), .B(n6578), .Z(n6591) );
  NANDN U6847 ( .A(n6382), .B(n6381), .Z(n6386) );
  NANDN U6848 ( .A(n6384), .B(n6383), .Z(n6385) );
  AND U6849 ( .A(n6386), .B(n6385), .Z(n6588) );
  NANDN U6850 ( .A(n6392), .B(n6391), .Z(n6396) );
  OR U6851 ( .A(n6394), .B(n6393), .Z(n6395) );
  AND U6852 ( .A(n6396), .B(n6395), .Z(n6583) );
  NANDN U6853 ( .A(n6398), .B(n6397), .Z(n6402) );
  NANDN U6854 ( .A(n6400), .B(n6399), .Z(n6401) );
  AND U6855 ( .A(n6402), .B(n6401), .Z(n6523) );
  NANDN U6856 ( .A(n6404), .B(n6403), .Z(n6408) );
  OR U6857 ( .A(n6406), .B(n6405), .Z(n6407) );
  NAND U6858 ( .A(n6408), .B(n6407), .Z(n6522) );
  XNOR U6859 ( .A(n6523), .B(n6522), .Z(n6524) );
  NAND U6860 ( .A(n583), .B(n6409), .Z(n6411) );
  XOR U6861 ( .A(b[29]), .B(a[27]), .Z(n6549) );
  NAND U6862 ( .A(n581), .B(n6549), .Z(n6410) );
  AND U6863 ( .A(n6411), .B(n6410), .Z(n6469) );
  AND U6864 ( .A(b[31]), .B(a[23]), .Z(n6468) );
  XNOR U6865 ( .A(n6469), .B(n6468), .Z(n6470) );
  NAND U6866 ( .A(b[0]), .B(a[55]), .Z(n6412) );
  XNOR U6867 ( .A(b[1]), .B(n6412), .Z(n6414) );
  NANDN U6868 ( .A(b[0]), .B(a[54]), .Z(n6413) );
  NAND U6869 ( .A(n6414), .B(n6413), .Z(n6471) );
  XNOR U6870 ( .A(n6470), .B(n6471), .Z(n6510) );
  NAND U6871 ( .A(n578), .B(n6415), .Z(n6417) );
  XOR U6872 ( .A(b[23]), .B(a[33]), .Z(n6552) );
  NAND U6873 ( .A(n9268), .B(n6552), .Z(n6416) );
  AND U6874 ( .A(n6417), .B(n6416), .Z(n6543) );
  NAND U6875 ( .A(n569), .B(n6418), .Z(n6420) );
  XOR U6876 ( .A(a[49]), .B(b[7]), .Z(n6555) );
  NAND U6877 ( .A(n7819), .B(n6555), .Z(n6419) );
  AND U6878 ( .A(n6420), .B(n6419), .Z(n6541) );
  NAND U6879 ( .A(n579), .B(n6421), .Z(n6423) );
  XOR U6880 ( .A(b[25]), .B(a[31]), .Z(n6558) );
  NAND U6881 ( .A(n9364), .B(n6558), .Z(n6422) );
  NAND U6882 ( .A(n6423), .B(n6422), .Z(n6540) );
  XNOR U6883 ( .A(n6541), .B(n6540), .Z(n6542) );
  XOR U6884 ( .A(n6543), .B(n6542), .Z(n6511) );
  XNOR U6885 ( .A(n6510), .B(n6511), .Z(n6512) );
  NAND U6886 ( .A(n572), .B(n6424), .Z(n6426) );
  XOR U6887 ( .A(b[13]), .B(a[43]), .Z(n6561) );
  NAND U6888 ( .A(n8585), .B(n6561), .Z(n6425) );
  AND U6889 ( .A(n6426), .B(n6425), .Z(n6505) );
  NAND U6890 ( .A(n571), .B(n6427), .Z(n6429) );
  XOR U6891 ( .A(a[45]), .B(b[11]), .Z(n6564) );
  NAND U6892 ( .A(n8135), .B(n6564), .Z(n6428) );
  NAND U6893 ( .A(n6429), .B(n6428), .Z(n6504) );
  XNOR U6894 ( .A(n6505), .B(n6504), .Z(n6506) );
  NAND U6895 ( .A(n573), .B(n6430), .Z(n6432) );
  XOR U6896 ( .A(b[15]), .B(a[41]), .Z(n6567) );
  NAND U6897 ( .A(n8694), .B(n6567), .Z(n6431) );
  AND U6898 ( .A(n6432), .B(n6431), .Z(n6501) );
  NAND U6899 ( .A(n577), .B(n6433), .Z(n6435) );
  XOR U6900 ( .A(b[21]), .B(a[35]), .Z(n6570) );
  NAND U6901 ( .A(n9216), .B(n6570), .Z(n6434) );
  AND U6902 ( .A(n6435), .B(n6434), .Z(n6499) );
  NAND U6903 ( .A(n570), .B(n6436), .Z(n6438) );
  XOR U6904 ( .A(a[47]), .B(b[9]), .Z(n6573) );
  NAND U6905 ( .A(n8037), .B(n6573), .Z(n6437) );
  NAND U6906 ( .A(n6438), .B(n6437), .Z(n6498) );
  XNOR U6907 ( .A(n6499), .B(n6498), .Z(n6500) );
  XOR U6908 ( .A(n6501), .B(n6500), .Z(n6507) );
  XOR U6909 ( .A(n6506), .B(n6507), .Z(n6513) );
  XOR U6910 ( .A(n6512), .B(n6513), .Z(n6525) );
  XNOR U6911 ( .A(n6524), .B(n6525), .Z(n6582) );
  XNOR U6912 ( .A(n6583), .B(n6582), .Z(n6584) );
  XOR U6913 ( .A(n6585), .B(n6584), .Z(n6589) );
  XNOR U6914 ( .A(n6588), .B(n6589), .Z(n6590) );
  XNOR U6915 ( .A(n6591), .B(n6590), .Z(n6464) );
  XOR U6916 ( .A(n6465), .B(n6464), .Z(n6457) );
  NANDN U6917 ( .A(n6440), .B(n6439), .Z(n6444) );
  OR U6918 ( .A(n6442), .B(n6441), .Z(n6443) );
  AND U6919 ( .A(n6444), .B(n6443), .Z(n6456) );
  XNOR U6920 ( .A(n6457), .B(n6456), .Z(n6458) );
  XNOR U6921 ( .A(n6459), .B(n6458), .Z(n6450) );
  XNOR U6922 ( .A(n6451), .B(n6450), .Z(n6452) );
  XNOR U6923 ( .A(n6453), .B(n6452), .Z(n6594) );
  XNOR U6924 ( .A(sreg[87]), .B(n6594), .Z(n6596) );
  NANDN U6925 ( .A(sreg[86]), .B(n6445), .Z(n6449) );
  NAND U6926 ( .A(n6447), .B(n6446), .Z(n6448) );
  NAND U6927 ( .A(n6449), .B(n6448), .Z(n6595) );
  XNOR U6928 ( .A(n6596), .B(n6595), .Z(c[87]) );
  NANDN U6929 ( .A(n6451), .B(n6450), .Z(n6455) );
  NANDN U6930 ( .A(n6453), .B(n6452), .Z(n6454) );
  AND U6931 ( .A(n6455), .B(n6454), .Z(n6602) );
  NANDN U6932 ( .A(n6457), .B(n6456), .Z(n6461) );
  NANDN U6933 ( .A(n6459), .B(n6458), .Z(n6460) );
  AND U6934 ( .A(n6461), .B(n6460), .Z(n6600) );
  NANDN U6935 ( .A(n6463), .B(n6462), .Z(n6467) );
  NAND U6936 ( .A(n6465), .B(n6464), .Z(n6466) );
  AND U6937 ( .A(n6467), .B(n6466), .Z(n6607) );
  NANDN U6938 ( .A(n6469), .B(n6468), .Z(n6473) );
  NANDN U6939 ( .A(n6471), .B(n6470), .Z(n6472) );
  AND U6940 ( .A(n6473), .B(n6472), .Z(n6691) );
  NAND U6941 ( .A(n582), .B(n6474), .Z(n6476) );
  XOR U6942 ( .A(b[27]), .B(a[30]), .Z(n6635) );
  NAND U6943 ( .A(n9770), .B(n6635), .Z(n6475) );
  AND U6944 ( .A(n6476), .B(n6475), .Z(n6698) );
  NAND U6945 ( .A(n567), .B(n6477), .Z(n6479) );
  XOR U6946 ( .A(a[52]), .B(b[5]), .Z(n6638) );
  NAND U6947 ( .A(n7235), .B(n6638), .Z(n6478) );
  AND U6948 ( .A(n6479), .B(n6478), .Z(n6696) );
  NAND U6949 ( .A(n9046), .B(n6480), .Z(n6482) );
  XOR U6950 ( .A(b[19]), .B(a[38]), .Z(n6641) );
  NAND U6951 ( .A(n575), .B(n6641), .Z(n6481) );
  NAND U6952 ( .A(n6482), .B(n6481), .Z(n6695) );
  XNOR U6953 ( .A(n6696), .B(n6695), .Z(n6697) );
  XNOR U6954 ( .A(n6698), .B(n6697), .Z(n6689) );
  NAND U6955 ( .A(n9764), .B(n6483), .Z(n6485) );
  XOR U6956 ( .A(b[31]), .B(a[26]), .Z(n6644) );
  NAND U6957 ( .A(n584), .B(n6644), .Z(n6484) );
  AND U6958 ( .A(n6485), .B(n6484), .Z(n6656) );
  NAND U6959 ( .A(n568), .B(n6486), .Z(n6488) );
  XOR U6960 ( .A(a[54]), .B(b[3]), .Z(n6647) );
  NAND U6961 ( .A(n7245), .B(n6647), .Z(n6487) );
  AND U6962 ( .A(n6488), .B(n6487), .Z(n6654) );
  NAND U6963 ( .A(n576), .B(n6489), .Z(n6491) );
  XOR U6964 ( .A(b[17]), .B(a[40]), .Z(n6650) );
  NAND U6965 ( .A(n9141), .B(n6650), .Z(n6490) );
  NAND U6966 ( .A(n6491), .B(n6490), .Z(n6653) );
  XNOR U6967 ( .A(n6654), .B(n6653), .Z(n6655) );
  XOR U6968 ( .A(n6656), .B(n6655), .Z(n6690) );
  XOR U6969 ( .A(n6689), .B(n6690), .Z(n6692) );
  XOR U6970 ( .A(n6691), .B(n6692), .Z(n6624) );
  NANDN U6971 ( .A(n6493), .B(n6492), .Z(n6497) );
  NANDN U6972 ( .A(n6495), .B(n6494), .Z(n6496) );
  AND U6973 ( .A(n6497), .B(n6496), .Z(n6677) );
  NANDN U6974 ( .A(n6499), .B(n6498), .Z(n6503) );
  NANDN U6975 ( .A(n6501), .B(n6500), .Z(n6502) );
  NAND U6976 ( .A(n6503), .B(n6502), .Z(n6678) );
  XNOR U6977 ( .A(n6677), .B(n6678), .Z(n6679) );
  NANDN U6978 ( .A(n6505), .B(n6504), .Z(n6509) );
  NANDN U6979 ( .A(n6507), .B(n6506), .Z(n6508) );
  NAND U6980 ( .A(n6509), .B(n6508), .Z(n6680) );
  XNOR U6981 ( .A(n6679), .B(n6680), .Z(n6623) );
  XNOR U6982 ( .A(n6624), .B(n6623), .Z(n6626) );
  NANDN U6983 ( .A(n6511), .B(n6510), .Z(n6515) );
  NANDN U6984 ( .A(n6513), .B(n6512), .Z(n6514) );
  AND U6985 ( .A(n6515), .B(n6514), .Z(n6625) );
  XOR U6986 ( .A(n6626), .B(n6625), .Z(n6739) );
  NANDN U6987 ( .A(n6517), .B(n6516), .Z(n6521) );
  NANDN U6988 ( .A(n6519), .B(n6518), .Z(n6520) );
  AND U6989 ( .A(n6521), .B(n6520), .Z(n6737) );
  NANDN U6990 ( .A(n6523), .B(n6522), .Z(n6527) );
  NANDN U6991 ( .A(n6525), .B(n6524), .Z(n6526) );
  AND U6992 ( .A(n6527), .B(n6526), .Z(n6620) );
  NANDN U6993 ( .A(n6529), .B(n6528), .Z(n6533) );
  OR U6994 ( .A(n6531), .B(n6530), .Z(n6532) );
  AND U6995 ( .A(n6533), .B(n6532), .Z(n6618) );
  NANDN U6996 ( .A(n6535), .B(n6534), .Z(n6539) );
  NANDN U6997 ( .A(n6537), .B(n6536), .Z(n6538) );
  AND U6998 ( .A(n6539), .B(n6538), .Z(n6684) );
  NANDN U6999 ( .A(n6541), .B(n6540), .Z(n6545) );
  NANDN U7000 ( .A(n6543), .B(n6542), .Z(n6544) );
  NAND U7001 ( .A(n6545), .B(n6544), .Z(n6683) );
  XNOR U7002 ( .A(n6684), .B(n6683), .Z(n6685) );
  NAND U7003 ( .A(b[0]), .B(a[56]), .Z(n6546) );
  XNOR U7004 ( .A(b[1]), .B(n6546), .Z(n6548) );
  NANDN U7005 ( .A(b[0]), .B(a[55]), .Z(n6547) );
  NAND U7006 ( .A(n6548), .B(n6547), .Z(n6632) );
  NAND U7007 ( .A(n583), .B(n6549), .Z(n6551) );
  XOR U7008 ( .A(b[29]), .B(a[28]), .Z(n6710) );
  NAND U7009 ( .A(n581), .B(n6710), .Z(n6550) );
  AND U7010 ( .A(n6551), .B(n6550), .Z(n6630) );
  AND U7011 ( .A(b[31]), .B(a[24]), .Z(n6629) );
  XNOR U7012 ( .A(n6630), .B(n6629), .Z(n6631) );
  XNOR U7013 ( .A(n6632), .B(n6631), .Z(n6671) );
  NAND U7014 ( .A(n578), .B(n6552), .Z(n6554) );
  XOR U7015 ( .A(b[23]), .B(a[34]), .Z(n6713) );
  NAND U7016 ( .A(n9268), .B(n6713), .Z(n6553) );
  AND U7017 ( .A(n6554), .B(n6553), .Z(n6704) );
  NAND U7018 ( .A(n569), .B(n6555), .Z(n6557) );
  XOR U7019 ( .A(a[50]), .B(b[7]), .Z(n6716) );
  NAND U7020 ( .A(n7819), .B(n6716), .Z(n6556) );
  AND U7021 ( .A(n6557), .B(n6556), .Z(n6702) );
  NAND U7022 ( .A(n579), .B(n6558), .Z(n6560) );
  XOR U7023 ( .A(b[25]), .B(a[32]), .Z(n6719) );
  NAND U7024 ( .A(n9364), .B(n6719), .Z(n6559) );
  NAND U7025 ( .A(n6560), .B(n6559), .Z(n6701) );
  XNOR U7026 ( .A(n6702), .B(n6701), .Z(n6703) );
  XOR U7027 ( .A(n6704), .B(n6703), .Z(n6672) );
  XNOR U7028 ( .A(n6671), .B(n6672), .Z(n6673) );
  NAND U7029 ( .A(n572), .B(n6561), .Z(n6563) );
  XOR U7030 ( .A(b[13]), .B(a[44]), .Z(n6722) );
  NAND U7031 ( .A(n8585), .B(n6722), .Z(n6562) );
  AND U7032 ( .A(n6563), .B(n6562), .Z(n6666) );
  NAND U7033 ( .A(n571), .B(n6564), .Z(n6566) );
  XOR U7034 ( .A(a[46]), .B(b[11]), .Z(n6725) );
  NAND U7035 ( .A(n8135), .B(n6725), .Z(n6565) );
  NAND U7036 ( .A(n6566), .B(n6565), .Z(n6665) );
  XNOR U7037 ( .A(n6666), .B(n6665), .Z(n6667) );
  NAND U7038 ( .A(n573), .B(n6567), .Z(n6569) );
  XOR U7039 ( .A(b[15]), .B(a[42]), .Z(n6728) );
  NAND U7040 ( .A(n8694), .B(n6728), .Z(n6568) );
  AND U7041 ( .A(n6569), .B(n6568), .Z(n6662) );
  NAND U7042 ( .A(n577), .B(n6570), .Z(n6572) );
  XOR U7043 ( .A(b[21]), .B(a[36]), .Z(n6731) );
  NAND U7044 ( .A(n9216), .B(n6731), .Z(n6571) );
  AND U7045 ( .A(n6572), .B(n6571), .Z(n6660) );
  NAND U7046 ( .A(n570), .B(n6573), .Z(n6575) );
  XOR U7047 ( .A(a[48]), .B(b[9]), .Z(n6734) );
  NAND U7048 ( .A(n8037), .B(n6734), .Z(n6574) );
  NAND U7049 ( .A(n6575), .B(n6574), .Z(n6659) );
  XNOR U7050 ( .A(n6660), .B(n6659), .Z(n6661) );
  XOR U7051 ( .A(n6662), .B(n6661), .Z(n6668) );
  XOR U7052 ( .A(n6667), .B(n6668), .Z(n6674) );
  XOR U7053 ( .A(n6673), .B(n6674), .Z(n6686) );
  XNOR U7054 ( .A(n6685), .B(n6686), .Z(n6617) );
  XNOR U7055 ( .A(n6618), .B(n6617), .Z(n6619) );
  XOR U7056 ( .A(n6620), .B(n6619), .Z(n6738) );
  XOR U7057 ( .A(n6737), .B(n6738), .Z(n6740) );
  XOR U7058 ( .A(n6739), .B(n6740), .Z(n6614) );
  NANDN U7059 ( .A(n6577), .B(n6576), .Z(n6581) );
  NAND U7060 ( .A(n6579), .B(n6578), .Z(n6580) );
  AND U7061 ( .A(n6581), .B(n6580), .Z(n6612) );
  NANDN U7062 ( .A(n6583), .B(n6582), .Z(n6587) );
  NANDN U7063 ( .A(n6585), .B(n6584), .Z(n6586) );
  AND U7064 ( .A(n6587), .B(n6586), .Z(n6611) );
  XNOR U7065 ( .A(n6612), .B(n6611), .Z(n6613) );
  XNOR U7066 ( .A(n6614), .B(n6613), .Z(n6605) );
  NANDN U7067 ( .A(n6589), .B(n6588), .Z(n6593) );
  NANDN U7068 ( .A(n6591), .B(n6590), .Z(n6592) );
  NAND U7069 ( .A(n6593), .B(n6592), .Z(n6606) );
  XOR U7070 ( .A(n6605), .B(n6606), .Z(n6608) );
  XNOR U7071 ( .A(n6607), .B(n6608), .Z(n6599) );
  XNOR U7072 ( .A(n6600), .B(n6599), .Z(n6601) );
  XNOR U7073 ( .A(n6602), .B(n6601), .Z(n6743) );
  XNOR U7074 ( .A(sreg[88]), .B(n6743), .Z(n6745) );
  NANDN U7075 ( .A(sreg[87]), .B(n6594), .Z(n6598) );
  NAND U7076 ( .A(n6596), .B(n6595), .Z(n6597) );
  NAND U7077 ( .A(n6598), .B(n6597), .Z(n6744) );
  XNOR U7078 ( .A(n6745), .B(n6744), .Z(c[88]) );
  NANDN U7079 ( .A(n6600), .B(n6599), .Z(n6604) );
  NANDN U7080 ( .A(n6602), .B(n6601), .Z(n6603) );
  AND U7081 ( .A(n6604), .B(n6603), .Z(n6751) );
  NANDN U7082 ( .A(n6606), .B(n6605), .Z(n6610) );
  NANDN U7083 ( .A(n6608), .B(n6607), .Z(n6609) );
  AND U7084 ( .A(n6610), .B(n6609), .Z(n6749) );
  NANDN U7085 ( .A(n6612), .B(n6611), .Z(n6616) );
  NANDN U7086 ( .A(n6614), .B(n6613), .Z(n6615) );
  AND U7087 ( .A(n6616), .B(n6615), .Z(n6757) );
  NANDN U7088 ( .A(n6618), .B(n6617), .Z(n6622) );
  NANDN U7089 ( .A(n6620), .B(n6619), .Z(n6621) );
  AND U7090 ( .A(n6622), .B(n6621), .Z(n6761) );
  NANDN U7091 ( .A(n6624), .B(n6623), .Z(n6628) );
  NAND U7092 ( .A(n6626), .B(n6625), .Z(n6627) );
  AND U7093 ( .A(n6628), .B(n6627), .Z(n6760) );
  XNOR U7094 ( .A(n6761), .B(n6760), .Z(n6763) );
  NANDN U7095 ( .A(n6630), .B(n6629), .Z(n6634) );
  NANDN U7096 ( .A(n6632), .B(n6631), .Z(n6633) );
  AND U7097 ( .A(n6634), .B(n6633), .Z(n6840) );
  NAND U7098 ( .A(n582), .B(n6635), .Z(n6637) );
  XOR U7099 ( .A(b[27]), .B(a[31]), .Z(n6784) );
  NAND U7100 ( .A(n9770), .B(n6784), .Z(n6636) );
  AND U7101 ( .A(n6637), .B(n6636), .Z(n6847) );
  NAND U7102 ( .A(n567), .B(n6638), .Z(n6640) );
  XOR U7103 ( .A(a[53]), .B(b[5]), .Z(n6787) );
  NAND U7104 ( .A(n7235), .B(n6787), .Z(n6639) );
  AND U7105 ( .A(n6640), .B(n6639), .Z(n6845) );
  NAND U7106 ( .A(n9046), .B(n6641), .Z(n6643) );
  XOR U7107 ( .A(b[19]), .B(a[39]), .Z(n6790) );
  NAND U7108 ( .A(n575), .B(n6790), .Z(n6642) );
  NAND U7109 ( .A(n6643), .B(n6642), .Z(n6844) );
  XNOR U7110 ( .A(n6845), .B(n6844), .Z(n6846) );
  XNOR U7111 ( .A(n6847), .B(n6846), .Z(n6838) );
  NAND U7112 ( .A(n9764), .B(n6644), .Z(n6646) );
  XOR U7113 ( .A(b[31]), .B(a[27]), .Z(n6793) );
  NAND U7114 ( .A(n584), .B(n6793), .Z(n6645) );
  AND U7115 ( .A(n6646), .B(n6645), .Z(n6805) );
  NAND U7116 ( .A(n568), .B(n6647), .Z(n6649) );
  XOR U7117 ( .A(a[55]), .B(b[3]), .Z(n6796) );
  NAND U7118 ( .A(n7245), .B(n6796), .Z(n6648) );
  AND U7119 ( .A(n6649), .B(n6648), .Z(n6803) );
  NAND U7120 ( .A(n576), .B(n6650), .Z(n6652) );
  XOR U7121 ( .A(b[17]), .B(a[41]), .Z(n6799) );
  NAND U7122 ( .A(n9141), .B(n6799), .Z(n6651) );
  NAND U7123 ( .A(n6652), .B(n6651), .Z(n6802) );
  XNOR U7124 ( .A(n6803), .B(n6802), .Z(n6804) );
  XOR U7125 ( .A(n6805), .B(n6804), .Z(n6839) );
  XOR U7126 ( .A(n6838), .B(n6839), .Z(n6841) );
  XOR U7127 ( .A(n6840), .B(n6841), .Z(n6773) );
  NANDN U7128 ( .A(n6654), .B(n6653), .Z(n6658) );
  NANDN U7129 ( .A(n6656), .B(n6655), .Z(n6657) );
  AND U7130 ( .A(n6658), .B(n6657), .Z(n6826) );
  NANDN U7131 ( .A(n6660), .B(n6659), .Z(n6664) );
  NANDN U7132 ( .A(n6662), .B(n6661), .Z(n6663) );
  NAND U7133 ( .A(n6664), .B(n6663), .Z(n6827) );
  XNOR U7134 ( .A(n6826), .B(n6827), .Z(n6828) );
  NANDN U7135 ( .A(n6666), .B(n6665), .Z(n6670) );
  NANDN U7136 ( .A(n6668), .B(n6667), .Z(n6669) );
  NAND U7137 ( .A(n6670), .B(n6669), .Z(n6829) );
  XNOR U7138 ( .A(n6828), .B(n6829), .Z(n6772) );
  XNOR U7139 ( .A(n6773), .B(n6772), .Z(n6775) );
  NANDN U7140 ( .A(n6672), .B(n6671), .Z(n6676) );
  NANDN U7141 ( .A(n6674), .B(n6673), .Z(n6675) );
  AND U7142 ( .A(n6676), .B(n6675), .Z(n6774) );
  XOR U7143 ( .A(n6775), .B(n6774), .Z(n6889) );
  NANDN U7144 ( .A(n6678), .B(n6677), .Z(n6682) );
  NANDN U7145 ( .A(n6680), .B(n6679), .Z(n6681) );
  AND U7146 ( .A(n6682), .B(n6681), .Z(n6886) );
  NANDN U7147 ( .A(n6684), .B(n6683), .Z(n6688) );
  NANDN U7148 ( .A(n6686), .B(n6685), .Z(n6687) );
  AND U7149 ( .A(n6688), .B(n6687), .Z(n6769) );
  NANDN U7150 ( .A(n6690), .B(n6689), .Z(n6694) );
  OR U7151 ( .A(n6692), .B(n6691), .Z(n6693) );
  AND U7152 ( .A(n6694), .B(n6693), .Z(n6767) );
  NANDN U7153 ( .A(n6696), .B(n6695), .Z(n6700) );
  NANDN U7154 ( .A(n6698), .B(n6697), .Z(n6699) );
  AND U7155 ( .A(n6700), .B(n6699), .Z(n6833) );
  NANDN U7156 ( .A(n6702), .B(n6701), .Z(n6706) );
  NANDN U7157 ( .A(n6704), .B(n6703), .Z(n6705) );
  NAND U7158 ( .A(n6706), .B(n6705), .Z(n6832) );
  XNOR U7159 ( .A(n6833), .B(n6832), .Z(n6834) );
  NAND U7160 ( .A(b[0]), .B(a[57]), .Z(n6707) );
  XNOR U7161 ( .A(b[1]), .B(n6707), .Z(n6709) );
  NANDN U7162 ( .A(b[0]), .B(a[56]), .Z(n6708) );
  NAND U7163 ( .A(n6709), .B(n6708), .Z(n6781) );
  NAND U7164 ( .A(n583), .B(n6710), .Z(n6712) );
  XOR U7165 ( .A(b[29]), .B(a[29]), .Z(n6856) );
  NAND U7166 ( .A(n581), .B(n6856), .Z(n6711) );
  AND U7167 ( .A(n6712), .B(n6711), .Z(n6779) );
  AND U7168 ( .A(b[31]), .B(a[25]), .Z(n6778) );
  XNOR U7169 ( .A(n6779), .B(n6778), .Z(n6780) );
  XNOR U7170 ( .A(n6781), .B(n6780), .Z(n6820) );
  NAND U7171 ( .A(n578), .B(n6713), .Z(n6715) );
  XOR U7172 ( .A(b[23]), .B(a[35]), .Z(n6862) );
  NAND U7173 ( .A(n9268), .B(n6862), .Z(n6714) );
  AND U7174 ( .A(n6715), .B(n6714), .Z(n6853) );
  NAND U7175 ( .A(n569), .B(n6716), .Z(n6718) );
  XOR U7176 ( .A(a[51]), .B(b[7]), .Z(n6865) );
  NAND U7177 ( .A(n7819), .B(n6865), .Z(n6717) );
  AND U7178 ( .A(n6718), .B(n6717), .Z(n6851) );
  NAND U7179 ( .A(n579), .B(n6719), .Z(n6721) );
  XOR U7180 ( .A(b[25]), .B(a[33]), .Z(n6868) );
  NAND U7181 ( .A(n9364), .B(n6868), .Z(n6720) );
  NAND U7182 ( .A(n6721), .B(n6720), .Z(n6850) );
  XNOR U7183 ( .A(n6851), .B(n6850), .Z(n6852) );
  XOR U7184 ( .A(n6853), .B(n6852), .Z(n6821) );
  XNOR U7185 ( .A(n6820), .B(n6821), .Z(n6822) );
  NAND U7186 ( .A(n572), .B(n6722), .Z(n6724) );
  XOR U7187 ( .A(b[13]), .B(a[45]), .Z(n6871) );
  NAND U7188 ( .A(n8585), .B(n6871), .Z(n6723) );
  AND U7189 ( .A(n6724), .B(n6723), .Z(n6815) );
  NAND U7190 ( .A(n571), .B(n6725), .Z(n6727) );
  XOR U7191 ( .A(a[47]), .B(b[11]), .Z(n6874) );
  NAND U7192 ( .A(n8135), .B(n6874), .Z(n6726) );
  NAND U7193 ( .A(n6727), .B(n6726), .Z(n6814) );
  XNOR U7194 ( .A(n6815), .B(n6814), .Z(n6816) );
  NAND U7195 ( .A(n573), .B(n6728), .Z(n6730) );
  XOR U7196 ( .A(b[15]), .B(a[43]), .Z(n6877) );
  NAND U7197 ( .A(n8694), .B(n6877), .Z(n6729) );
  AND U7198 ( .A(n6730), .B(n6729), .Z(n6811) );
  NAND U7199 ( .A(n577), .B(n6731), .Z(n6733) );
  XOR U7200 ( .A(b[21]), .B(a[37]), .Z(n6880) );
  NAND U7201 ( .A(n9216), .B(n6880), .Z(n6732) );
  AND U7202 ( .A(n6733), .B(n6732), .Z(n6809) );
  NAND U7203 ( .A(n570), .B(n6734), .Z(n6736) );
  XOR U7204 ( .A(a[49]), .B(b[9]), .Z(n6883) );
  NAND U7205 ( .A(n8037), .B(n6883), .Z(n6735) );
  NAND U7206 ( .A(n6736), .B(n6735), .Z(n6808) );
  XNOR U7207 ( .A(n6809), .B(n6808), .Z(n6810) );
  XOR U7208 ( .A(n6811), .B(n6810), .Z(n6817) );
  XOR U7209 ( .A(n6816), .B(n6817), .Z(n6823) );
  XOR U7210 ( .A(n6822), .B(n6823), .Z(n6835) );
  XNOR U7211 ( .A(n6834), .B(n6835), .Z(n6766) );
  XNOR U7212 ( .A(n6767), .B(n6766), .Z(n6768) );
  XOR U7213 ( .A(n6769), .B(n6768), .Z(n6887) );
  XNOR U7214 ( .A(n6886), .B(n6887), .Z(n6888) );
  XNOR U7215 ( .A(n6889), .B(n6888), .Z(n6762) );
  XOR U7216 ( .A(n6763), .B(n6762), .Z(n6755) );
  NANDN U7217 ( .A(n6738), .B(n6737), .Z(n6742) );
  OR U7218 ( .A(n6740), .B(n6739), .Z(n6741) );
  AND U7219 ( .A(n6742), .B(n6741), .Z(n6754) );
  XNOR U7220 ( .A(n6755), .B(n6754), .Z(n6756) );
  XNOR U7221 ( .A(n6757), .B(n6756), .Z(n6748) );
  XNOR U7222 ( .A(n6749), .B(n6748), .Z(n6750) );
  XNOR U7223 ( .A(n6751), .B(n6750), .Z(n6892) );
  XNOR U7224 ( .A(sreg[89]), .B(n6892), .Z(n6894) );
  NANDN U7225 ( .A(sreg[88]), .B(n6743), .Z(n6747) );
  NAND U7226 ( .A(n6745), .B(n6744), .Z(n6746) );
  NAND U7227 ( .A(n6747), .B(n6746), .Z(n6893) );
  XNOR U7228 ( .A(n6894), .B(n6893), .Z(c[89]) );
  NANDN U7229 ( .A(n6749), .B(n6748), .Z(n6753) );
  NANDN U7230 ( .A(n6751), .B(n6750), .Z(n6752) );
  AND U7231 ( .A(n6753), .B(n6752), .Z(n6900) );
  NANDN U7232 ( .A(n6755), .B(n6754), .Z(n6759) );
  NANDN U7233 ( .A(n6757), .B(n6756), .Z(n6758) );
  AND U7234 ( .A(n6759), .B(n6758), .Z(n6898) );
  NANDN U7235 ( .A(n6761), .B(n6760), .Z(n6765) );
  NAND U7236 ( .A(n6763), .B(n6762), .Z(n6764) );
  AND U7237 ( .A(n6765), .B(n6764), .Z(n6905) );
  NANDN U7238 ( .A(n6767), .B(n6766), .Z(n6771) );
  NANDN U7239 ( .A(n6769), .B(n6768), .Z(n6770) );
  AND U7240 ( .A(n6771), .B(n6770), .Z(n6910) );
  NANDN U7241 ( .A(n6773), .B(n6772), .Z(n6777) );
  NAND U7242 ( .A(n6775), .B(n6774), .Z(n6776) );
  AND U7243 ( .A(n6777), .B(n6776), .Z(n6909) );
  XNOR U7244 ( .A(n6910), .B(n6909), .Z(n6912) );
  NANDN U7245 ( .A(n6779), .B(n6778), .Z(n6783) );
  NANDN U7246 ( .A(n6781), .B(n6780), .Z(n6782) );
  AND U7247 ( .A(n6783), .B(n6782), .Z(n6989) );
  NAND U7248 ( .A(n582), .B(n6784), .Z(n6786) );
  XOR U7249 ( .A(b[27]), .B(a[32]), .Z(n6933) );
  NAND U7250 ( .A(n9770), .B(n6933), .Z(n6785) );
  AND U7251 ( .A(n6786), .B(n6785), .Z(n6996) );
  NAND U7252 ( .A(n567), .B(n6787), .Z(n6789) );
  XOR U7253 ( .A(a[54]), .B(b[5]), .Z(n6936) );
  NAND U7254 ( .A(n7235), .B(n6936), .Z(n6788) );
  AND U7255 ( .A(n6789), .B(n6788), .Z(n6994) );
  NAND U7256 ( .A(n9046), .B(n6790), .Z(n6792) );
  XOR U7257 ( .A(b[19]), .B(a[40]), .Z(n6939) );
  NAND U7258 ( .A(n575), .B(n6939), .Z(n6791) );
  NAND U7259 ( .A(n6792), .B(n6791), .Z(n6993) );
  XNOR U7260 ( .A(n6994), .B(n6993), .Z(n6995) );
  XNOR U7261 ( .A(n6996), .B(n6995), .Z(n6987) );
  NAND U7262 ( .A(n9764), .B(n6793), .Z(n6795) );
  XOR U7263 ( .A(b[31]), .B(a[28]), .Z(n6942) );
  NAND U7264 ( .A(n584), .B(n6942), .Z(n6794) );
  AND U7265 ( .A(n6795), .B(n6794), .Z(n6954) );
  NAND U7266 ( .A(n568), .B(n6796), .Z(n6798) );
  XOR U7267 ( .A(a[56]), .B(b[3]), .Z(n6945) );
  NAND U7268 ( .A(n7245), .B(n6945), .Z(n6797) );
  AND U7269 ( .A(n6798), .B(n6797), .Z(n6952) );
  NAND U7270 ( .A(n576), .B(n6799), .Z(n6801) );
  XOR U7271 ( .A(b[17]), .B(a[42]), .Z(n6948) );
  NAND U7272 ( .A(n9141), .B(n6948), .Z(n6800) );
  NAND U7273 ( .A(n6801), .B(n6800), .Z(n6951) );
  XNOR U7274 ( .A(n6952), .B(n6951), .Z(n6953) );
  XOR U7275 ( .A(n6954), .B(n6953), .Z(n6988) );
  XOR U7276 ( .A(n6987), .B(n6988), .Z(n6990) );
  XOR U7277 ( .A(n6989), .B(n6990), .Z(n6922) );
  NANDN U7278 ( .A(n6803), .B(n6802), .Z(n6807) );
  NANDN U7279 ( .A(n6805), .B(n6804), .Z(n6806) );
  AND U7280 ( .A(n6807), .B(n6806), .Z(n6975) );
  NANDN U7281 ( .A(n6809), .B(n6808), .Z(n6813) );
  NANDN U7282 ( .A(n6811), .B(n6810), .Z(n6812) );
  NAND U7283 ( .A(n6813), .B(n6812), .Z(n6976) );
  XNOR U7284 ( .A(n6975), .B(n6976), .Z(n6977) );
  NANDN U7285 ( .A(n6815), .B(n6814), .Z(n6819) );
  NANDN U7286 ( .A(n6817), .B(n6816), .Z(n6818) );
  NAND U7287 ( .A(n6819), .B(n6818), .Z(n6978) );
  XNOR U7288 ( .A(n6977), .B(n6978), .Z(n6921) );
  XNOR U7289 ( .A(n6922), .B(n6921), .Z(n6924) );
  NANDN U7290 ( .A(n6821), .B(n6820), .Z(n6825) );
  NANDN U7291 ( .A(n6823), .B(n6822), .Z(n6824) );
  AND U7292 ( .A(n6825), .B(n6824), .Z(n6923) );
  XOR U7293 ( .A(n6924), .B(n6923), .Z(n7038) );
  NANDN U7294 ( .A(n6827), .B(n6826), .Z(n6831) );
  NANDN U7295 ( .A(n6829), .B(n6828), .Z(n6830) );
  AND U7296 ( .A(n6831), .B(n6830), .Z(n7035) );
  NANDN U7297 ( .A(n6833), .B(n6832), .Z(n6837) );
  NANDN U7298 ( .A(n6835), .B(n6834), .Z(n6836) );
  AND U7299 ( .A(n6837), .B(n6836), .Z(n6918) );
  NANDN U7300 ( .A(n6839), .B(n6838), .Z(n6843) );
  OR U7301 ( .A(n6841), .B(n6840), .Z(n6842) );
  AND U7302 ( .A(n6843), .B(n6842), .Z(n6916) );
  NANDN U7303 ( .A(n6845), .B(n6844), .Z(n6849) );
  NANDN U7304 ( .A(n6847), .B(n6846), .Z(n6848) );
  AND U7305 ( .A(n6849), .B(n6848), .Z(n6982) );
  NANDN U7306 ( .A(n6851), .B(n6850), .Z(n6855) );
  NANDN U7307 ( .A(n6853), .B(n6852), .Z(n6854) );
  NAND U7308 ( .A(n6855), .B(n6854), .Z(n6981) );
  XNOR U7309 ( .A(n6982), .B(n6981), .Z(n6983) );
  NAND U7310 ( .A(n583), .B(n6856), .Z(n6858) );
  XOR U7311 ( .A(b[29]), .B(a[30]), .Z(n7005) );
  NAND U7312 ( .A(n581), .B(n7005), .Z(n6857) );
  AND U7313 ( .A(n6858), .B(n6857), .Z(n6928) );
  AND U7314 ( .A(b[31]), .B(a[26]), .Z(n6927) );
  XNOR U7315 ( .A(n6928), .B(n6927), .Z(n6929) );
  NAND U7316 ( .A(b[0]), .B(a[58]), .Z(n6859) );
  XNOR U7317 ( .A(b[1]), .B(n6859), .Z(n6861) );
  NANDN U7318 ( .A(b[0]), .B(a[57]), .Z(n6860) );
  NAND U7319 ( .A(n6861), .B(n6860), .Z(n6930) );
  XNOR U7320 ( .A(n6929), .B(n6930), .Z(n6969) );
  NAND U7321 ( .A(n578), .B(n6862), .Z(n6864) );
  XOR U7322 ( .A(b[23]), .B(a[36]), .Z(n7011) );
  NAND U7323 ( .A(n9268), .B(n7011), .Z(n6863) );
  AND U7324 ( .A(n6864), .B(n6863), .Z(n7002) );
  NAND U7325 ( .A(n569), .B(n6865), .Z(n6867) );
  XOR U7326 ( .A(a[52]), .B(b[7]), .Z(n7014) );
  NAND U7327 ( .A(n7819), .B(n7014), .Z(n6866) );
  AND U7328 ( .A(n6867), .B(n6866), .Z(n7000) );
  NAND U7329 ( .A(n579), .B(n6868), .Z(n6870) );
  XOR U7330 ( .A(b[25]), .B(a[34]), .Z(n7017) );
  NAND U7331 ( .A(n9364), .B(n7017), .Z(n6869) );
  NAND U7332 ( .A(n6870), .B(n6869), .Z(n6999) );
  XNOR U7333 ( .A(n7000), .B(n6999), .Z(n7001) );
  XOR U7334 ( .A(n7002), .B(n7001), .Z(n6970) );
  XNOR U7335 ( .A(n6969), .B(n6970), .Z(n6971) );
  NAND U7336 ( .A(n572), .B(n6871), .Z(n6873) );
  XOR U7337 ( .A(b[13]), .B(a[46]), .Z(n7020) );
  NAND U7338 ( .A(n8585), .B(n7020), .Z(n6872) );
  AND U7339 ( .A(n6873), .B(n6872), .Z(n6964) );
  NAND U7340 ( .A(n571), .B(n6874), .Z(n6876) );
  XOR U7341 ( .A(a[48]), .B(b[11]), .Z(n7023) );
  NAND U7342 ( .A(n8135), .B(n7023), .Z(n6875) );
  NAND U7343 ( .A(n6876), .B(n6875), .Z(n6963) );
  XNOR U7344 ( .A(n6964), .B(n6963), .Z(n6965) );
  NAND U7345 ( .A(n573), .B(n6877), .Z(n6879) );
  XOR U7346 ( .A(b[15]), .B(a[44]), .Z(n7026) );
  NAND U7347 ( .A(n8694), .B(n7026), .Z(n6878) );
  AND U7348 ( .A(n6879), .B(n6878), .Z(n6960) );
  NAND U7349 ( .A(n577), .B(n6880), .Z(n6882) );
  XOR U7350 ( .A(b[21]), .B(a[38]), .Z(n7029) );
  NAND U7351 ( .A(n9216), .B(n7029), .Z(n6881) );
  AND U7352 ( .A(n6882), .B(n6881), .Z(n6958) );
  NAND U7353 ( .A(n570), .B(n6883), .Z(n6885) );
  XOR U7354 ( .A(a[50]), .B(b[9]), .Z(n7032) );
  NAND U7355 ( .A(n8037), .B(n7032), .Z(n6884) );
  NAND U7356 ( .A(n6885), .B(n6884), .Z(n6957) );
  XNOR U7357 ( .A(n6958), .B(n6957), .Z(n6959) );
  XOR U7358 ( .A(n6960), .B(n6959), .Z(n6966) );
  XOR U7359 ( .A(n6965), .B(n6966), .Z(n6972) );
  XOR U7360 ( .A(n6971), .B(n6972), .Z(n6984) );
  XNOR U7361 ( .A(n6983), .B(n6984), .Z(n6915) );
  XNOR U7362 ( .A(n6916), .B(n6915), .Z(n6917) );
  XOR U7363 ( .A(n6918), .B(n6917), .Z(n7036) );
  XNOR U7364 ( .A(n7035), .B(n7036), .Z(n7037) );
  XNOR U7365 ( .A(n7038), .B(n7037), .Z(n6911) );
  XOR U7366 ( .A(n6912), .B(n6911), .Z(n6904) );
  NANDN U7367 ( .A(n6887), .B(n6886), .Z(n6891) );
  NANDN U7368 ( .A(n6889), .B(n6888), .Z(n6890) );
  AND U7369 ( .A(n6891), .B(n6890), .Z(n6903) );
  XOR U7370 ( .A(n6904), .B(n6903), .Z(n6906) );
  XNOR U7371 ( .A(n6905), .B(n6906), .Z(n6897) );
  XNOR U7372 ( .A(n6898), .B(n6897), .Z(n6899) );
  XNOR U7373 ( .A(n6900), .B(n6899), .Z(n7041) );
  XNOR U7374 ( .A(sreg[90]), .B(n7041), .Z(n7043) );
  NANDN U7375 ( .A(sreg[89]), .B(n6892), .Z(n6896) );
  NAND U7376 ( .A(n6894), .B(n6893), .Z(n6895) );
  NAND U7377 ( .A(n6896), .B(n6895), .Z(n7042) );
  XNOR U7378 ( .A(n7043), .B(n7042), .Z(c[90]) );
  NANDN U7379 ( .A(n6898), .B(n6897), .Z(n6902) );
  NANDN U7380 ( .A(n6900), .B(n6899), .Z(n6901) );
  AND U7381 ( .A(n6902), .B(n6901), .Z(n7049) );
  NANDN U7382 ( .A(n6904), .B(n6903), .Z(n6908) );
  NANDN U7383 ( .A(n6906), .B(n6905), .Z(n6907) );
  AND U7384 ( .A(n6908), .B(n6907), .Z(n7047) );
  NANDN U7385 ( .A(n6910), .B(n6909), .Z(n6914) );
  NAND U7386 ( .A(n6912), .B(n6911), .Z(n6913) );
  AND U7387 ( .A(n6914), .B(n6913), .Z(n7054) );
  NANDN U7388 ( .A(n6916), .B(n6915), .Z(n6920) );
  NANDN U7389 ( .A(n6918), .B(n6917), .Z(n6919) );
  AND U7390 ( .A(n6920), .B(n6919), .Z(n7059) );
  NANDN U7391 ( .A(n6922), .B(n6921), .Z(n6926) );
  NAND U7392 ( .A(n6924), .B(n6923), .Z(n6925) );
  AND U7393 ( .A(n6926), .B(n6925), .Z(n7058) );
  XNOR U7394 ( .A(n7059), .B(n7058), .Z(n7061) );
  NANDN U7395 ( .A(n6928), .B(n6927), .Z(n6932) );
  NANDN U7396 ( .A(n6930), .B(n6929), .Z(n6931) );
  AND U7397 ( .A(n6932), .B(n6931), .Z(n7138) );
  NAND U7398 ( .A(n582), .B(n6933), .Z(n6935) );
  XOR U7399 ( .A(b[27]), .B(a[33]), .Z(n7082) );
  NAND U7400 ( .A(n9770), .B(n7082), .Z(n6934) );
  AND U7401 ( .A(n6935), .B(n6934), .Z(n7145) );
  NAND U7402 ( .A(n567), .B(n6936), .Z(n6938) );
  XOR U7403 ( .A(a[55]), .B(b[5]), .Z(n7085) );
  NAND U7404 ( .A(n7235), .B(n7085), .Z(n6937) );
  AND U7405 ( .A(n6938), .B(n6937), .Z(n7143) );
  NAND U7406 ( .A(n9046), .B(n6939), .Z(n6941) );
  XOR U7407 ( .A(b[19]), .B(a[41]), .Z(n7088) );
  NAND U7408 ( .A(n575), .B(n7088), .Z(n6940) );
  NAND U7409 ( .A(n6941), .B(n6940), .Z(n7142) );
  XNOR U7410 ( .A(n7143), .B(n7142), .Z(n7144) );
  XNOR U7411 ( .A(n7145), .B(n7144), .Z(n7136) );
  NAND U7412 ( .A(n9764), .B(n6942), .Z(n6944) );
  XOR U7413 ( .A(b[31]), .B(a[29]), .Z(n7091) );
  NAND U7414 ( .A(n584), .B(n7091), .Z(n6943) );
  AND U7415 ( .A(n6944), .B(n6943), .Z(n7103) );
  NAND U7416 ( .A(n568), .B(n6945), .Z(n6947) );
  XOR U7417 ( .A(a[57]), .B(b[3]), .Z(n7094) );
  NAND U7418 ( .A(n7245), .B(n7094), .Z(n6946) );
  AND U7419 ( .A(n6947), .B(n6946), .Z(n7101) );
  NAND U7420 ( .A(n576), .B(n6948), .Z(n6950) );
  XOR U7421 ( .A(b[17]), .B(a[43]), .Z(n7097) );
  NAND U7422 ( .A(n9141), .B(n7097), .Z(n6949) );
  NAND U7423 ( .A(n6950), .B(n6949), .Z(n7100) );
  XNOR U7424 ( .A(n7101), .B(n7100), .Z(n7102) );
  XOR U7425 ( .A(n7103), .B(n7102), .Z(n7137) );
  XOR U7426 ( .A(n7136), .B(n7137), .Z(n7139) );
  XOR U7427 ( .A(n7138), .B(n7139), .Z(n7071) );
  NANDN U7428 ( .A(n6952), .B(n6951), .Z(n6956) );
  NANDN U7429 ( .A(n6954), .B(n6953), .Z(n6955) );
  AND U7430 ( .A(n6956), .B(n6955), .Z(n7124) );
  NANDN U7431 ( .A(n6958), .B(n6957), .Z(n6962) );
  NANDN U7432 ( .A(n6960), .B(n6959), .Z(n6961) );
  NAND U7433 ( .A(n6962), .B(n6961), .Z(n7125) );
  XNOR U7434 ( .A(n7124), .B(n7125), .Z(n7126) );
  NANDN U7435 ( .A(n6964), .B(n6963), .Z(n6968) );
  NANDN U7436 ( .A(n6966), .B(n6965), .Z(n6967) );
  NAND U7437 ( .A(n6968), .B(n6967), .Z(n7127) );
  XNOR U7438 ( .A(n7126), .B(n7127), .Z(n7070) );
  XNOR U7439 ( .A(n7071), .B(n7070), .Z(n7073) );
  NANDN U7440 ( .A(n6970), .B(n6969), .Z(n6974) );
  NANDN U7441 ( .A(n6972), .B(n6971), .Z(n6973) );
  AND U7442 ( .A(n6974), .B(n6973), .Z(n7072) );
  XOR U7443 ( .A(n7073), .B(n7072), .Z(n7187) );
  NANDN U7444 ( .A(n6976), .B(n6975), .Z(n6980) );
  NANDN U7445 ( .A(n6978), .B(n6977), .Z(n6979) );
  AND U7446 ( .A(n6980), .B(n6979), .Z(n7184) );
  NANDN U7447 ( .A(n6982), .B(n6981), .Z(n6986) );
  NANDN U7448 ( .A(n6984), .B(n6983), .Z(n6985) );
  AND U7449 ( .A(n6986), .B(n6985), .Z(n7067) );
  NANDN U7450 ( .A(n6988), .B(n6987), .Z(n6992) );
  OR U7451 ( .A(n6990), .B(n6989), .Z(n6991) );
  AND U7452 ( .A(n6992), .B(n6991), .Z(n7065) );
  NANDN U7453 ( .A(n6994), .B(n6993), .Z(n6998) );
  NANDN U7454 ( .A(n6996), .B(n6995), .Z(n6997) );
  AND U7455 ( .A(n6998), .B(n6997), .Z(n7131) );
  NANDN U7456 ( .A(n7000), .B(n6999), .Z(n7004) );
  NANDN U7457 ( .A(n7002), .B(n7001), .Z(n7003) );
  NAND U7458 ( .A(n7004), .B(n7003), .Z(n7130) );
  XNOR U7459 ( .A(n7131), .B(n7130), .Z(n7132) );
  NAND U7460 ( .A(n583), .B(n7005), .Z(n7007) );
  XOR U7461 ( .A(b[29]), .B(a[31]), .Z(n7157) );
  NAND U7462 ( .A(n581), .B(n7157), .Z(n7006) );
  AND U7463 ( .A(n7007), .B(n7006), .Z(n7077) );
  AND U7464 ( .A(b[31]), .B(a[27]), .Z(n7076) );
  XNOR U7465 ( .A(n7077), .B(n7076), .Z(n7078) );
  NAND U7466 ( .A(b[0]), .B(a[59]), .Z(n7008) );
  XNOR U7467 ( .A(b[1]), .B(n7008), .Z(n7010) );
  NANDN U7468 ( .A(b[0]), .B(a[58]), .Z(n7009) );
  NAND U7469 ( .A(n7010), .B(n7009), .Z(n7079) );
  XNOR U7470 ( .A(n7078), .B(n7079), .Z(n7118) );
  NAND U7471 ( .A(n578), .B(n7011), .Z(n7013) );
  XOR U7472 ( .A(b[23]), .B(a[37]), .Z(n7160) );
  NAND U7473 ( .A(n9268), .B(n7160), .Z(n7012) );
  AND U7474 ( .A(n7013), .B(n7012), .Z(n7151) );
  NAND U7475 ( .A(n569), .B(n7014), .Z(n7016) );
  XOR U7476 ( .A(a[53]), .B(b[7]), .Z(n7163) );
  NAND U7477 ( .A(n7819), .B(n7163), .Z(n7015) );
  AND U7478 ( .A(n7016), .B(n7015), .Z(n7149) );
  NAND U7479 ( .A(n579), .B(n7017), .Z(n7019) );
  XOR U7480 ( .A(b[25]), .B(a[35]), .Z(n7166) );
  NAND U7481 ( .A(n9364), .B(n7166), .Z(n7018) );
  NAND U7482 ( .A(n7019), .B(n7018), .Z(n7148) );
  XNOR U7483 ( .A(n7149), .B(n7148), .Z(n7150) );
  XOR U7484 ( .A(n7151), .B(n7150), .Z(n7119) );
  XNOR U7485 ( .A(n7118), .B(n7119), .Z(n7120) );
  NAND U7486 ( .A(n572), .B(n7020), .Z(n7022) );
  XOR U7487 ( .A(a[47]), .B(b[13]), .Z(n7169) );
  NAND U7488 ( .A(n8585), .B(n7169), .Z(n7021) );
  AND U7489 ( .A(n7022), .B(n7021), .Z(n7113) );
  NAND U7490 ( .A(n571), .B(n7023), .Z(n7025) );
  XOR U7491 ( .A(a[49]), .B(b[11]), .Z(n7172) );
  NAND U7492 ( .A(n8135), .B(n7172), .Z(n7024) );
  NAND U7493 ( .A(n7025), .B(n7024), .Z(n7112) );
  XNOR U7494 ( .A(n7113), .B(n7112), .Z(n7114) );
  NAND U7495 ( .A(n573), .B(n7026), .Z(n7028) );
  XOR U7496 ( .A(b[15]), .B(a[45]), .Z(n7175) );
  NAND U7497 ( .A(n8694), .B(n7175), .Z(n7027) );
  AND U7498 ( .A(n7028), .B(n7027), .Z(n7109) );
  NAND U7499 ( .A(n577), .B(n7029), .Z(n7031) );
  XOR U7500 ( .A(b[21]), .B(a[39]), .Z(n7178) );
  NAND U7501 ( .A(n9216), .B(n7178), .Z(n7030) );
  AND U7502 ( .A(n7031), .B(n7030), .Z(n7107) );
  NAND U7503 ( .A(n570), .B(n7032), .Z(n7034) );
  XOR U7504 ( .A(a[51]), .B(b[9]), .Z(n7181) );
  NAND U7505 ( .A(n8037), .B(n7181), .Z(n7033) );
  NAND U7506 ( .A(n7034), .B(n7033), .Z(n7106) );
  XNOR U7507 ( .A(n7107), .B(n7106), .Z(n7108) );
  XOR U7508 ( .A(n7109), .B(n7108), .Z(n7115) );
  XOR U7509 ( .A(n7114), .B(n7115), .Z(n7121) );
  XOR U7510 ( .A(n7120), .B(n7121), .Z(n7133) );
  XNOR U7511 ( .A(n7132), .B(n7133), .Z(n7064) );
  XNOR U7512 ( .A(n7065), .B(n7064), .Z(n7066) );
  XOR U7513 ( .A(n7067), .B(n7066), .Z(n7185) );
  XNOR U7514 ( .A(n7184), .B(n7185), .Z(n7186) );
  XNOR U7515 ( .A(n7187), .B(n7186), .Z(n7060) );
  XOR U7516 ( .A(n7061), .B(n7060), .Z(n7053) );
  NANDN U7517 ( .A(n7036), .B(n7035), .Z(n7040) );
  NANDN U7518 ( .A(n7038), .B(n7037), .Z(n7039) );
  AND U7519 ( .A(n7040), .B(n7039), .Z(n7052) );
  XOR U7520 ( .A(n7053), .B(n7052), .Z(n7055) );
  XNOR U7521 ( .A(n7054), .B(n7055), .Z(n7046) );
  XNOR U7522 ( .A(n7047), .B(n7046), .Z(n7048) );
  XNOR U7523 ( .A(n7049), .B(n7048), .Z(n7190) );
  XNOR U7524 ( .A(sreg[91]), .B(n7190), .Z(n7192) );
  NANDN U7525 ( .A(sreg[90]), .B(n7041), .Z(n7045) );
  NAND U7526 ( .A(n7043), .B(n7042), .Z(n7044) );
  NAND U7527 ( .A(n7045), .B(n7044), .Z(n7191) );
  XNOR U7528 ( .A(n7192), .B(n7191), .Z(c[91]) );
  NANDN U7529 ( .A(n7047), .B(n7046), .Z(n7051) );
  NANDN U7530 ( .A(n7049), .B(n7048), .Z(n7050) );
  AND U7531 ( .A(n7051), .B(n7050), .Z(n7198) );
  NANDN U7532 ( .A(n7053), .B(n7052), .Z(n7057) );
  NANDN U7533 ( .A(n7055), .B(n7054), .Z(n7056) );
  AND U7534 ( .A(n7057), .B(n7056), .Z(n7196) );
  NANDN U7535 ( .A(n7059), .B(n7058), .Z(n7063) );
  NAND U7536 ( .A(n7061), .B(n7060), .Z(n7062) );
  AND U7537 ( .A(n7063), .B(n7062), .Z(n7335) );
  NANDN U7538 ( .A(n7065), .B(n7064), .Z(n7069) );
  NANDN U7539 ( .A(n7067), .B(n7066), .Z(n7068) );
  AND U7540 ( .A(n7069), .B(n7068), .Z(n7202) );
  NANDN U7541 ( .A(n7071), .B(n7070), .Z(n7075) );
  NAND U7542 ( .A(n7073), .B(n7072), .Z(n7074) );
  AND U7543 ( .A(n7075), .B(n7074), .Z(n7201) );
  XNOR U7544 ( .A(n7202), .B(n7201), .Z(n7204) );
  NANDN U7545 ( .A(n7077), .B(n7076), .Z(n7081) );
  NANDN U7546 ( .A(n7079), .B(n7078), .Z(n7080) );
  AND U7547 ( .A(n7081), .B(n7080), .Z(n7287) );
  NAND U7548 ( .A(n582), .B(n7082), .Z(n7084) );
  XOR U7549 ( .A(b[27]), .B(a[34]), .Z(n7231) );
  NAND U7550 ( .A(n9770), .B(n7231), .Z(n7083) );
  AND U7551 ( .A(n7084), .B(n7083), .Z(n7330) );
  NAND U7552 ( .A(n567), .B(n7085), .Z(n7087) );
  XOR U7553 ( .A(a[56]), .B(b[5]), .Z(n7234) );
  NAND U7554 ( .A(n7235), .B(n7234), .Z(n7086) );
  AND U7555 ( .A(n7087), .B(n7086), .Z(n7328) );
  NAND U7556 ( .A(n9046), .B(n7088), .Z(n7090) );
  XOR U7557 ( .A(b[19]), .B(a[42]), .Z(n7238) );
  NAND U7558 ( .A(n575), .B(n7238), .Z(n7089) );
  NAND U7559 ( .A(n7090), .B(n7089), .Z(n7327) );
  XNOR U7560 ( .A(n7328), .B(n7327), .Z(n7329) );
  XNOR U7561 ( .A(n7330), .B(n7329), .Z(n7285) );
  NAND U7562 ( .A(n9764), .B(n7091), .Z(n7093) );
  XOR U7563 ( .A(b[31]), .B(a[30]), .Z(n7241) );
  NAND U7564 ( .A(n584), .B(n7241), .Z(n7092) );
  AND U7565 ( .A(n7093), .B(n7092), .Z(n7254) );
  NAND U7566 ( .A(n568), .B(n7094), .Z(n7096) );
  XOR U7567 ( .A(a[58]), .B(b[3]), .Z(n7244) );
  NAND U7568 ( .A(n7245), .B(n7244), .Z(n7095) );
  AND U7569 ( .A(n7096), .B(n7095), .Z(n7252) );
  NAND U7570 ( .A(n576), .B(n7097), .Z(n7099) );
  XOR U7571 ( .A(b[17]), .B(a[44]), .Z(n7248) );
  NAND U7572 ( .A(n9141), .B(n7248), .Z(n7098) );
  NAND U7573 ( .A(n7099), .B(n7098), .Z(n7251) );
  XNOR U7574 ( .A(n7252), .B(n7251), .Z(n7253) );
  XOR U7575 ( .A(n7254), .B(n7253), .Z(n7286) );
  XOR U7576 ( .A(n7285), .B(n7286), .Z(n7288) );
  XOR U7577 ( .A(n7287), .B(n7288), .Z(n7220) );
  NANDN U7578 ( .A(n7101), .B(n7100), .Z(n7105) );
  NANDN U7579 ( .A(n7103), .B(n7102), .Z(n7104) );
  AND U7580 ( .A(n7105), .B(n7104), .Z(n7275) );
  NANDN U7581 ( .A(n7107), .B(n7106), .Z(n7111) );
  NANDN U7582 ( .A(n7109), .B(n7108), .Z(n7110) );
  NAND U7583 ( .A(n7111), .B(n7110), .Z(n7276) );
  XNOR U7584 ( .A(n7275), .B(n7276), .Z(n7277) );
  NANDN U7585 ( .A(n7113), .B(n7112), .Z(n7117) );
  NANDN U7586 ( .A(n7115), .B(n7114), .Z(n7116) );
  NAND U7587 ( .A(n7117), .B(n7116), .Z(n7278) );
  XNOR U7588 ( .A(n7277), .B(n7278), .Z(n7219) );
  XNOR U7589 ( .A(n7220), .B(n7219), .Z(n7222) );
  NANDN U7590 ( .A(n7119), .B(n7118), .Z(n7123) );
  NANDN U7591 ( .A(n7121), .B(n7120), .Z(n7122) );
  AND U7592 ( .A(n7123), .B(n7122), .Z(n7221) );
  XOR U7593 ( .A(n7222), .B(n7221), .Z(n7210) );
  NANDN U7594 ( .A(n7125), .B(n7124), .Z(n7129) );
  NANDN U7595 ( .A(n7127), .B(n7126), .Z(n7128) );
  AND U7596 ( .A(n7129), .B(n7128), .Z(n7207) );
  NANDN U7597 ( .A(n7131), .B(n7130), .Z(n7135) );
  NANDN U7598 ( .A(n7133), .B(n7132), .Z(n7134) );
  AND U7599 ( .A(n7135), .B(n7134), .Z(n7216) );
  NANDN U7600 ( .A(n7137), .B(n7136), .Z(n7141) );
  OR U7601 ( .A(n7139), .B(n7138), .Z(n7140) );
  AND U7602 ( .A(n7141), .B(n7140), .Z(n7214) );
  NANDN U7603 ( .A(n7143), .B(n7142), .Z(n7147) );
  NANDN U7604 ( .A(n7145), .B(n7144), .Z(n7146) );
  AND U7605 ( .A(n7147), .B(n7146), .Z(n7282) );
  NANDN U7606 ( .A(n7149), .B(n7148), .Z(n7153) );
  NANDN U7607 ( .A(n7151), .B(n7150), .Z(n7152) );
  NAND U7608 ( .A(n7153), .B(n7152), .Z(n7281) );
  XNOR U7609 ( .A(n7282), .B(n7281), .Z(n7284) );
  NAND U7610 ( .A(b[0]), .B(a[60]), .Z(n7154) );
  XNOR U7611 ( .A(b[1]), .B(n7154), .Z(n7156) );
  NANDN U7612 ( .A(b[0]), .B(a[59]), .Z(n7155) );
  NAND U7613 ( .A(n7156), .B(n7155), .Z(n7228) );
  NAND U7614 ( .A(n583), .B(n7157), .Z(n7159) );
  XOR U7615 ( .A(b[29]), .B(a[32]), .Z(n7303) );
  NAND U7616 ( .A(n581), .B(n7303), .Z(n7158) );
  AND U7617 ( .A(n7159), .B(n7158), .Z(n7226) );
  AND U7618 ( .A(b[31]), .B(a[28]), .Z(n7225) );
  XNOR U7619 ( .A(n7226), .B(n7225), .Z(n7227) );
  XNOR U7620 ( .A(n7228), .B(n7227), .Z(n7269) );
  NAND U7621 ( .A(n578), .B(n7160), .Z(n7162) );
  XOR U7622 ( .A(b[23]), .B(a[38]), .Z(n7291) );
  NAND U7623 ( .A(n9268), .B(n7291), .Z(n7161) );
  AND U7624 ( .A(n7162), .B(n7161), .Z(n7324) );
  NAND U7625 ( .A(n569), .B(n7163), .Z(n7165) );
  XOR U7626 ( .A(a[54]), .B(b[7]), .Z(n7294) );
  NAND U7627 ( .A(n7819), .B(n7294), .Z(n7164) );
  AND U7628 ( .A(n7165), .B(n7164), .Z(n7322) );
  NAND U7629 ( .A(n579), .B(n7166), .Z(n7168) );
  XOR U7630 ( .A(b[25]), .B(a[36]), .Z(n7297) );
  NAND U7631 ( .A(n9364), .B(n7297), .Z(n7167) );
  NAND U7632 ( .A(n7168), .B(n7167), .Z(n7321) );
  XNOR U7633 ( .A(n7322), .B(n7321), .Z(n7323) );
  XOR U7634 ( .A(n7324), .B(n7323), .Z(n7270) );
  XNOR U7635 ( .A(n7269), .B(n7270), .Z(n7271) );
  NAND U7636 ( .A(n572), .B(n7169), .Z(n7171) );
  XOR U7637 ( .A(a[48]), .B(b[13]), .Z(n7306) );
  NAND U7638 ( .A(n8585), .B(n7306), .Z(n7170) );
  AND U7639 ( .A(n7171), .B(n7170), .Z(n7264) );
  NAND U7640 ( .A(n571), .B(n7172), .Z(n7174) );
  XOR U7641 ( .A(a[50]), .B(b[11]), .Z(n7309) );
  NAND U7642 ( .A(n8135), .B(n7309), .Z(n7173) );
  NAND U7643 ( .A(n7174), .B(n7173), .Z(n7263) );
  XNOR U7644 ( .A(n7264), .B(n7263), .Z(n7265) );
  NAND U7645 ( .A(n573), .B(n7175), .Z(n7177) );
  XOR U7646 ( .A(b[15]), .B(a[46]), .Z(n7312) );
  NAND U7647 ( .A(n8694), .B(n7312), .Z(n7176) );
  AND U7648 ( .A(n7177), .B(n7176), .Z(n7260) );
  NAND U7649 ( .A(n577), .B(n7178), .Z(n7180) );
  XOR U7650 ( .A(b[21]), .B(a[40]), .Z(n7315) );
  NAND U7651 ( .A(n9216), .B(n7315), .Z(n7179) );
  AND U7652 ( .A(n7180), .B(n7179), .Z(n7258) );
  NAND U7653 ( .A(n570), .B(n7181), .Z(n7183) );
  XOR U7654 ( .A(a[52]), .B(b[9]), .Z(n7318) );
  NAND U7655 ( .A(n8037), .B(n7318), .Z(n7182) );
  NAND U7656 ( .A(n7183), .B(n7182), .Z(n7257) );
  XNOR U7657 ( .A(n7258), .B(n7257), .Z(n7259) );
  XOR U7658 ( .A(n7260), .B(n7259), .Z(n7266) );
  XOR U7659 ( .A(n7265), .B(n7266), .Z(n7272) );
  XOR U7660 ( .A(n7271), .B(n7272), .Z(n7283) );
  XNOR U7661 ( .A(n7284), .B(n7283), .Z(n7213) );
  XNOR U7662 ( .A(n7214), .B(n7213), .Z(n7215) );
  XOR U7663 ( .A(n7216), .B(n7215), .Z(n7208) );
  XNOR U7664 ( .A(n7207), .B(n7208), .Z(n7209) );
  XNOR U7665 ( .A(n7210), .B(n7209), .Z(n7203) );
  XOR U7666 ( .A(n7204), .B(n7203), .Z(n7334) );
  NANDN U7667 ( .A(n7185), .B(n7184), .Z(n7189) );
  NANDN U7668 ( .A(n7187), .B(n7186), .Z(n7188) );
  AND U7669 ( .A(n7189), .B(n7188), .Z(n7333) );
  XOR U7670 ( .A(n7334), .B(n7333), .Z(n7336) );
  XNOR U7671 ( .A(n7335), .B(n7336), .Z(n7195) );
  XNOR U7672 ( .A(n7196), .B(n7195), .Z(n7197) );
  XNOR U7673 ( .A(n7198), .B(n7197), .Z(n7339) );
  XNOR U7674 ( .A(sreg[92]), .B(n7339), .Z(n7341) );
  NANDN U7675 ( .A(sreg[91]), .B(n7190), .Z(n7194) );
  NAND U7676 ( .A(n7192), .B(n7191), .Z(n7193) );
  NAND U7677 ( .A(n7194), .B(n7193), .Z(n7340) );
  XNOR U7678 ( .A(n7341), .B(n7340), .Z(c[92]) );
  NANDN U7679 ( .A(n7196), .B(n7195), .Z(n7200) );
  NANDN U7680 ( .A(n7198), .B(n7197), .Z(n7199) );
  AND U7681 ( .A(n7200), .B(n7199), .Z(n7347) );
  NANDN U7682 ( .A(n7202), .B(n7201), .Z(n7206) );
  NAND U7683 ( .A(n7204), .B(n7203), .Z(n7205) );
  AND U7684 ( .A(n7206), .B(n7205), .Z(n7478) );
  NANDN U7685 ( .A(n7208), .B(n7207), .Z(n7212) );
  NANDN U7686 ( .A(n7210), .B(n7209), .Z(n7211) );
  AND U7687 ( .A(n7212), .B(n7211), .Z(n7477) );
  NANDN U7688 ( .A(n7214), .B(n7213), .Z(n7218) );
  NANDN U7689 ( .A(n7216), .B(n7215), .Z(n7217) );
  AND U7690 ( .A(n7218), .B(n7217), .Z(n7471) );
  NANDN U7691 ( .A(n7220), .B(n7219), .Z(n7224) );
  NAND U7692 ( .A(n7222), .B(n7221), .Z(n7223) );
  AND U7693 ( .A(n7224), .B(n7223), .Z(n7470) );
  XNOR U7694 ( .A(n7471), .B(n7470), .Z(n7472) );
  NANDN U7695 ( .A(n7226), .B(n7225), .Z(n7230) );
  NANDN U7696 ( .A(n7228), .B(n7227), .Z(n7229) );
  AND U7697 ( .A(n7230), .B(n7229), .Z(n7442) );
  NAND U7698 ( .A(n582), .B(n7231), .Z(n7233) );
  XOR U7699 ( .A(b[27]), .B(a[35]), .Z(n7360) );
  NAND U7700 ( .A(n9770), .B(n7360), .Z(n7232) );
  AND U7701 ( .A(n7233), .B(n7232), .Z(n7433) );
  NAND U7702 ( .A(n567), .B(n7234), .Z(n7237) );
  XOR U7703 ( .A(a[57]), .B(b[5]), .Z(n7363) );
  NAND U7704 ( .A(n7235), .B(n7363), .Z(n7236) );
  AND U7705 ( .A(n7237), .B(n7236), .Z(n7431) );
  NAND U7706 ( .A(n9046), .B(n7238), .Z(n7240) );
  XOR U7707 ( .A(b[19]), .B(a[43]), .Z(n7366) );
  NAND U7708 ( .A(n575), .B(n7366), .Z(n7239) );
  NAND U7709 ( .A(n7240), .B(n7239), .Z(n7430) );
  XNOR U7710 ( .A(n7431), .B(n7430), .Z(n7432) );
  XNOR U7711 ( .A(n7433), .B(n7432), .Z(n7440) );
  NAND U7712 ( .A(n9764), .B(n7241), .Z(n7243) );
  XOR U7713 ( .A(b[31]), .B(a[31]), .Z(n7369) );
  NAND U7714 ( .A(n584), .B(n7369), .Z(n7242) );
  AND U7715 ( .A(n7243), .B(n7242), .Z(n7385) );
  NAND U7716 ( .A(n568), .B(n7244), .Z(n7247) );
  XOR U7717 ( .A(a[59]), .B(b[3]), .Z(n7372) );
  NAND U7718 ( .A(n7245), .B(n7372), .Z(n7246) );
  AND U7719 ( .A(n7247), .B(n7246), .Z(n7383) );
  NAND U7720 ( .A(n576), .B(n7248), .Z(n7250) );
  XOR U7721 ( .A(b[17]), .B(a[45]), .Z(n7375) );
  NAND U7722 ( .A(n9141), .B(n7375), .Z(n7249) );
  NAND U7723 ( .A(n7250), .B(n7249), .Z(n7382) );
  XNOR U7724 ( .A(n7383), .B(n7382), .Z(n7384) );
  XOR U7725 ( .A(n7385), .B(n7384), .Z(n7441) );
  XOR U7726 ( .A(n7440), .B(n7441), .Z(n7443) );
  XOR U7727 ( .A(n7442), .B(n7443), .Z(n7453) );
  NANDN U7728 ( .A(n7252), .B(n7251), .Z(n7256) );
  NANDN U7729 ( .A(n7254), .B(n7253), .Z(n7255) );
  AND U7730 ( .A(n7256), .B(n7255), .Z(n7446) );
  NANDN U7731 ( .A(n7258), .B(n7257), .Z(n7262) );
  NANDN U7732 ( .A(n7260), .B(n7259), .Z(n7261) );
  NAND U7733 ( .A(n7262), .B(n7261), .Z(n7447) );
  XNOR U7734 ( .A(n7446), .B(n7447), .Z(n7448) );
  NANDN U7735 ( .A(n7264), .B(n7263), .Z(n7268) );
  NANDN U7736 ( .A(n7266), .B(n7265), .Z(n7267) );
  NAND U7737 ( .A(n7268), .B(n7267), .Z(n7449) );
  XNOR U7738 ( .A(n7448), .B(n7449), .Z(n7452) );
  XNOR U7739 ( .A(n7453), .B(n7452), .Z(n7455) );
  NANDN U7740 ( .A(n7270), .B(n7269), .Z(n7274) );
  NANDN U7741 ( .A(n7272), .B(n7271), .Z(n7273) );
  AND U7742 ( .A(n7274), .B(n7273), .Z(n7454) );
  XOR U7743 ( .A(n7455), .B(n7454), .Z(n7467) );
  NANDN U7744 ( .A(n7276), .B(n7275), .Z(n7280) );
  NANDN U7745 ( .A(n7278), .B(n7277), .Z(n7279) );
  AND U7746 ( .A(n7280), .B(n7279), .Z(n7464) );
  NANDN U7747 ( .A(n7286), .B(n7285), .Z(n7290) );
  OR U7748 ( .A(n7288), .B(n7287), .Z(n7289) );
  AND U7749 ( .A(n7290), .B(n7289), .Z(n7459) );
  NANDN U7750 ( .A(n563), .B(n7291), .Z(n7293) );
  XNOR U7751 ( .A(b[23]), .B(a[39]), .Z(n7415) );
  OR U7752 ( .A(n7415), .B(n9605), .Z(n7292) );
  NAND U7753 ( .A(n7293), .B(n7292), .Z(n7438) );
  NANDN U7754 ( .A(n558), .B(n7294), .Z(n7296) );
  XNOR U7755 ( .A(a[55]), .B(b[7]), .Z(n7418) );
  OR U7756 ( .A(n7418), .B(n8290), .Z(n7295) );
  AND U7757 ( .A(n7296), .B(n7295), .Z(n7436) );
  NANDN U7758 ( .A(n566), .B(n7297), .Z(n7299) );
  XOR U7759 ( .A(b[25]), .B(a[37]), .Z(n7421) );
  NANDN U7760 ( .A(n9684), .B(n7421), .Z(n7298) );
  NAND U7761 ( .A(n7299), .B(n7298), .Z(n7437) );
  XOR U7762 ( .A(n7436), .B(n7437), .Z(n7439) );
  XOR U7763 ( .A(n7438), .B(n7439), .Z(n7351) );
  NAND U7764 ( .A(b[0]), .B(a[61]), .Z(n7300) );
  XNOR U7765 ( .A(b[1]), .B(n7300), .Z(n7302) );
  NANDN U7766 ( .A(b[0]), .B(a[60]), .Z(n7301) );
  NAND U7767 ( .A(n7302), .B(n7301), .Z(n7359) );
  NANDN U7768 ( .A(n559), .B(n7303), .Z(n7305) );
  XNOR U7769 ( .A(b[29]), .B(a[33]), .Z(n7427) );
  OR U7770 ( .A(n7427), .B(n9796), .Z(n7304) );
  NAND U7771 ( .A(n7305), .B(n7304), .Z(n7357) );
  NAND U7772 ( .A(b[31]), .B(a[29]), .Z(n7356) );
  XOR U7773 ( .A(n7357), .B(n7356), .Z(n7358) );
  XNOR U7774 ( .A(n7359), .B(n7358), .Z(n7350) );
  XOR U7775 ( .A(n7351), .B(n7350), .Z(n7353) );
  NANDN U7776 ( .A(n553), .B(n7306), .Z(n7308) );
  XNOR U7777 ( .A(a[49]), .B(b[13]), .Z(n7400) );
  OR U7778 ( .A(n7400), .B(n8853), .Z(n7307) );
  NAND U7779 ( .A(n7308), .B(n7307), .Z(n7390) );
  NANDN U7780 ( .A(n562), .B(n7309), .Z(n7311) );
  XNOR U7781 ( .A(a[51]), .B(b[11]), .Z(n7403) );
  OR U7782 ( .A(n7403), .B(n8701), .Z(n7310) );
  NAND U7783 ( .A(n7311), .B(n7310), .Z(n7388) );
  NANDN U7784 ( .A(n557), .B(n7312), .Z(n7314) );
  XNOR U7785 ( .A(b[15]), .B(a[47]), .Z(n7406) );
  OR U7786 ( .A(n7406), .B(n9067), .Z(n7313) );
  NAND U7787 ( .A(n7314), .B(n7313), .Z(n7380) );
  NANDN U7788 ( .A(n556), .B(n7315), .Z(n7317) );
  XNOR U7789 ( .A(b[21]), .B(a[41]), .Z(n7409) );
  OR U7790 ( .A(n7409), .B(n9480), .Z(n7316) );
  AND U7791 ( .A(n7317), .B(n7316), .Z(n7378) );
  NANDN U7792 ( .A(n564), .B(n7318), .Z(n7320) );
  XOR U7793 ( .A(a[53]), .B(b[9]), .Z(n7412) );
  NANDN U7794 ( .A(n8485), .B(n7412), .Z(n7319) );
  NAND U7795 ( .A(n7320), .B(n7319), .Z(n7379) );
  XOR U7796 ( .A(n7378), .B(n7379), .Z(n7381) );
  XOR U7797 ( .A(n7380), .B(n7381), .Z(n7389) );
  XOR U7798 ( .A(n7388), .B(n7389), .Z(n7391) );
  XOR U7799 ( .A(n7390), .B(n7391), .Z(n7352) );
  XOR U7800 ( .A(n7353), .B(n7352), .Z(n7397) );
  NANDN U7801 ( .A(n7322), .B(n7321), .Z(n7326) );
  NANDN U7802 ( .A(n7324), .B(n7323), .Z(n7325) );
  AND U7803 ( .A(n7326), .B(n7325), .Z(n7395) );
  NANDN U7804 ( .A(n7328), .B(n7327), .Z(n7332) );
  NANDN U7805 ( .A(n7330), .B(n7329), .Z(n7331) );
  NAND U7806 ( .A(n7332), .B(n7331), .Z(n7394) );
  XNOR U7807 ( .A(n7395), .B(n7394), .Z(n7396) );
  XNOR U7808 ( .A(n7397), .B(n7396), .Z(n7458) );
  XNOR U7809 ( .A(n7459), .B(n7458), .Z(n7460) );
  XOR U7810 ( .A(n7461), .B(n7460), .Z(n7465) );
  XNOR U7811 ( .A(n7464), .B(n7465), .Z(n7466) );
  XOR U7812 ( .A(n7467), .B(n7466), .Z(n7473) );
  XNOR U7813 ( .A(n7472), .B(n7473), .Z(n7476) );
  XOR U7814 ( .A(n7477), .B(n7476), .Z(n7479) );
  XOR U7815 ( .A(n7478), .B(n7479), .Z(n7345) );
  NANDN U7816 ( .A(n7334), .B(n7333), .Z(n7338) );
  NANDN U7817 ( .A(n7336), .B(n7335), .Z(n7337) );
  NAND U7818 ( .A(n7338), .B(n7337), .Z(n7344) );
  XNOR U7819 ( .A(n7345), .B(n7344), .Z(n7346) );
  XNOR U7820 ( .A(n7347), .B(n7346), .Z(n7482) );
  XNOR U7821 ( .A(sreg[93]), .B(n7482), .Z(n7484) );
  NANDN U7822 ( .A(sreg[92]), .B(n7339), .Z(n7343) );
  NAND U7823 ( .A(n7341), .B(n7340), .Z(n7342) );
  NAND U7824 ( .A(n7343), .B(n7342), .Z(n7483) );
  XNOR U7825 ( .A(n7484), .B(n7483), .Z(c[93]) );
  NANDN U7826 ( .A(n7345), .B(n7344), .Z(n7349) );
  NANDN U7827 ( .A(n7347), .B(n7346), .Z(n7348) );
  AND U7828 ( .A(n7349), .B(n7348), .Z(n7490) );
  NAND U7829 ( .A(n7351), .B(n7350), .Z(n7355) );
  NAND U7830 ( .A(n7353), .B(n7352), .Z(n7354) );
  AND U7831 ( .A(n7355), .B(n7354), .Z(n7507) );
  NANDN U7832 ( .A(n565), .B(n7360), .Z(n7362) );
  XNOR U7833 ( .A(b[27]), .B(a[36]), .Z(n7534) );
  OR U7834 ( .A(n7534), .B(n9692), .Z(n7361) );
  AND U7835 ( .A(n7362), .B(n7361), .Z(n7596) );
  NANDN U7836 ( .A(n561), .B(n7363), .Z(n7365) );
  XNOR U7837 ( .A(a[58]), .B(b[5]), .Z(n7537) );
  OR U7838 ( .A(n7537), .B(n8041), .Z(n7364) );
  AND U7839 ( .A(n7365), .B(n7364), .Z(n7594) );
  NAND U7840 ( .A(n9046), .B(n7366), .Z(n7368) );
  XOR U7841 ( .A(b[19]), .B(a[44]), .Z(n7540) );
  NAND U7842 ( .A(n575), .B(n7540), .Z(n7367) );
  NAND U7843 ( .A(n7368), .B(n7367), .Z(n7595) );
  XNOR U7844 ( .A(n7594), .B(n7595), .Z(n7597) );
  XNOR U7845 ( .A(n7596), .B(n7597), .Z(n7556) );
  NANDN U7846 ( .A(n580), .B(n7369), .Z(n7371) );
  XNOR U7847 ( .A(b[31]), .B(a[32]), .Z(n7543) );
  OR U7848 ( .A(n7543), .B(n9904), .Z(n7370) );
  NAND U7849 ( .A(n7371), .B(n7370), .Z(n7522) );
  NANDN U7850 ( .A(n560), .B(n7372), .Z(n7374) );
  XNOR U7851 ( .A(a[60]), .B(b[3]), .Z(n7546) );
  OR U7852 ( .A(n7546), .B(n7784), .Z(n7373) );
  AND U7853 ( .A(n7374), .B(n7373), .Z(n7519) );
  NANDN U7854 ( .A(n554), .B(n7375), .Z(n7377) );
  XOR U7855 ( .A(b[17]), .B(a[46]), .Z(n7549) );
  NANDN U7856 ( .A(n9195), .B(n7549), .Z(n7376) );
  NAND U7857 ( .A(n7377), .B(n7376), .Z(n7520) );
  XOR U7858 ( .A(n7519), .B(n7520), .Z(n7523) );
  XOR U7859 ( .A(n7522), .B(n7523), .Z(n7557) );
  XNOR U7860 ( .A(n7556), .B(n7557), .Z(n7559) );
  XNOR U7861 ( .A(n7558), .B(n7559), .Z(n7506) );
  NANDN U7862 ( .A(n7383), .B(n7382), .Z(n7387) );
  NANDN U7863 ( .A(n7385), .B(n7384), .Z(n7386) );
  NAND U7864 ( .A(n7387), .B(n7386), .Z(n7598) );
  XNOR U7865 ( .A(n7599), .B(n7598), .Z(n7601) );
  NANDN U7866 ( .A(n7389), .B(n7388), .Z(n7393) );
  NANDN U7867 ( .A(n7391), .B(n7390), .Z(n7392) );
  NAND U7868 ( .A(n7393), .B(n7392), .Z(n7600) );
  XNOR U7869 ( .A(n7601), .B(n7600), .Z(n7505) );
  XNOR U7870 ( .A(n7506), .B(n7505), .Z(n7508) );
  XNOR U7871 ( .A(n7507), .B(n7508), .Z(n7500) );
  NANDN U7872 ( .A(n7395), .B(n7394), .Z(n7399) );
  NANDN U7873 ( .A(n7397), .B(n7396), .Z(n7398) );
  AND U7874 ( .A(n7399), .B(n7398), .Z(n7503) );
  OR U7875 ( .A(n7400), .B(n553), .Z(n7402) );
  XNOR U7876 ( .A(a[50]), .B(b[13]), .Z(n7560) );
  OR U7877 ( .A(n7560), .B(n8853), .Z(n7401) );
  AND U7878 ( .A(n7402), .B(n7401), .Z(n7528) );
  OR U7879 ( .A(n7403), .B(n562), .Z(n7405) );
  XNOR U7880 ( .A(a[52]), .B(b[11]), .Z(n7563) );
  OR U7881 ( .A(n7563), .B(n8701), .Z(n7404) );
  AND U7882 ( .A(n7405), .B(n7404), .Z(n7526) );
  OR U7883 ( .A(n7406), .B(n557), .Z(n7408) );
  XNOR U7884 ( .A(b[15]), .B(a[48]), .Z(n7566) );
  OR U7885 ( .A(n7566), .B(n9067), .Z(n7407) );
  AND U7886 ( .A(n7408), .B(n7407), .Z(n7517) );
  OR U7887 ( .A(n7409), .B(n556), .Z(n7411) );
  XNOR U7888 ( .A(b[21]), .B(a[42]), .Z(n7569) );
  OR U7889 ( .A(n7569), .B(n9480), .Z(n7410) );
  AND U7890 ( .A(n7411), .B(n7410), .Z(n7515) );
  NAND U7891 ( .A(n570), .B(n7412), .Z(n7414) );
  XOR U7892 ( .A(a[54]), .B(b[9]), .Z(n7572) );
  NAND U7893 ( .A(n8037), .B(n7572), .Z(n7413) );
  NAND U7894 ( .A(n7414), .B(n7413), .Z(n7516) );
  XNOR U7895 ( .A(n7515), .B(n7516), .Z(n7518) );
  XNOR U7896 ( .A(n7517), .B(n7518), .Z(n7527) );
  XNOR U7897 ( .A(n7526), .B(n7527), .Z(n7529) );
  XNOR U7898 ( .A(n7528), .B(n7529), .Z(n7512) );
  OR U7899 ( .A(n7415), .B(n563), .Z(n7417) );
  XNOR U7900 ( .A(b[23]), .B(a[40]), .Z(n7575) );
  OR U7901 ( .A(n7575), .B(n9605), .Z(n7416) );
  AND U7902 ( .A(n7417), .B(n7416), .Z(n7592) );
  OR U7903 ( .A(n7418), .B(n558), .Z(n7420) );
  XNOR U7904 ( .A(a[56]), .B(b[7]), .Z(n7578) );
  OR U7905 ( .A(n7578), .B(n8290), .Z(n7419) );
  AND U7906 ( .A(n7420), .B(n7419), .Z(n7590) );
  NAND U7907 ( .A(n579), .B(n7421), .Z(n7423) );
  XOR U7908 ( .A(b[25]), .B(a[38]), .Z(n7581) );
  NAND U7909 ( .A(n9364), .B(n7581), .Z(n7422) );
  NAND U7910 ( .A(n7423), .B(n7422), .Z(n7591) );
  XNOR U7911 ( .A(n7590), .B(n7591), .Z(n7593) );
  XNOR U7912 ( .A(n7592), .B(n7593), .Z(n7510) );
  NAND U7913 ( .A(b[0]), .B(a[62]), .Z(n7424) );
  XNOR U7914 ( .A(b[1]), .B(n7424), .Z(n7426) );
  NANDN U7915 ( .A(b[0]), .B(a[61]), .Z(n7425) );
  NAND U7916 ( .A(n7426), .B(n7425), .Z(n7533) );
  OR U7917 ( .A(n7427), .B(n559), .Z(n7429) );
  XNOR U7918 ( .A(b[29]), .B(a[34]), .Z(n7587) );
  OR U7919 ( .A(n7587), .B(n9796), .Z(n7428) );
  NAND U7920 ( .A(n7429), .B(n7428), .Z(n7531) );
  NAND U7921 ( .A(b[31]), .B(a[30]), .Z(n7530) );
  XOR U7922 ( .A(n7531), .B(n7530), .Z(n7532) );
  XNOR U7923 ( .A(n7533), .B(n7532), .Z(n7509) );
  XNOR U7924 ( .A(n7510), .B(n7509), .Z(n7511) );
  XNOR U7925 ( .A(n7512), .B(n7511), .Z(n7555) );
  NANDN U7926 ( .A(n7431), .B(n7430), .Z(n7435) );
  NANDN U7927 ( .A(n7433), .B(n7432), .Z(n7434) );
  AND U7928 ( .A(n7435), .B(n7434), .Z(n7552) );
  XNOR U7929 ( .A(n7552), .B(n7553), .Z(n7554) );
  XOR U7930 ( .A(n7555), .B(n7554), .Z(n7502) );
  NANDN U7931 ( .A(n7441), .B(n7440), .Z(n7445) );
  OR U7932 ( .A(n7443), .B(n7442), .Z(n7444) );
  NAND U7933 ( .A(n7445), .B(n7444), .Z(n7501) );
  XOR U7934 ( .A(n7502), .B(n7501), .Z(n7504) );
  XNOR U7935 ( .A(n7503), .B(n7504), .Z(n7497) );
  NANDN U7936 ( .A(n7447), .B(n7446), .Z(n7451) );
  NANDN U7937 ( .A(n7449), .B(n7448), .Z(n7450) );
  AND U7938 ( .A(n7451), .B(n7450), .Z(n7498) );
  XNOR U7939 ( .A(n7497), .B(n7498), .Z(n7499) );
  XNOR U7940 ( .A(n7500), .B(n7499), .Z(n7495) );
  NANDN U7941 ( .A(n7453), .B(n7452), .Z(n7457) );
  NAND U7942 ( .A(n7455), .B(n7454), .Z(n7456) );
  AND U7943 ( .A(n7457), .B(n7456), .Z(n7493) );
  NANDN U7944 ( .A(n7459), .B(n7458), .Z(n7463) );
  NANDN U7945 ( .A(n7461), .B(n7460), .Z(n7462) );
  AND U7946 ( .A(n7463), .B(n7462), .Z(n7494) );
  XNOR U7947 ( .A(n7493), .B(n7494), .Z(n7496) );
  XNOR U7948 ( .A(n7495), .B(n7496), .Z(n7603) );
  NANDN U7949 ( .A(n7465), .B(n7464), .Z(n7469) );
  NANDN U7950 ( .A(n7467), .B(n7466), .Z(n7468) );
  NAND U7951 ( .A(n7469), .B(n7468), .Z(n7602) );
  XNOR U7952 ( .A(n7603), .B(n7602), .Z(n7605) );
  NANDN U7953 ( .A(n7471), .B(n7470), .Z(n7475) );
  NANDN U7954 ( .A(n7473), .B(n7472), .Z(n7474) );
  NAND U7955 ( .A(n7475), .B(n7474), .Z(n7604) );
  XNOR U7956 ( .A(n7605), .B(n7604), .Z(n7487) );
  NANDN U7957 ( .A(n7477), .B(n7476), .Z(n7481) );
  OR U7958 ( .A(n7479), .B(n7478), .Z(n7480) );
  NAND U7959 ( .A(n7481), .B(n7480), .Z(n7488) );
  XNOR U7960 ( .A(n7487), .B(n7488), .Z(n7489) );
  XNOR U7961 ( .A(n7490), .B(n7489), .Z(n7606) );
  XNOR U7962 ( .A(sreg[94]), .B(n7606), .Z(n7608) );
  NANDN U7963 ( .A(sreg[93]), .B(n7482), .Z(n7486) );
  NAND U7964 ( .A(n7484), .B(n7483), .Z(n7485) );
  NAND U7965 ( .A(n7486), .B(n7485), .Z(n7607) );
  XNOR U7966 ( .A(n7608), .B(n7607), .Z(c[94]) );
  NANDN U7967 ( .A(n7488), .B(n7487), .Z(n7492) );
  NANDN U7968 ( .A(n7490), .B(n7489), .Z(n7491) );
  AND U7969 ( .A(n7492), .B(n7491), .Z(n7618) );
  XNOR U7970 ( .A(n7620), .B(n7621), .Z(n7623) );
  NANDN U7971 ( .A(n7510), .B(n7509), .Z(n7514) );
  NANDN U7972 ( .A(n7512), .B(n7511), .Z(n7513) );
  AND U7973 ( .A(n7514), .B(n7513), .Z(n7729) );
  IV U7974 ( .A(n7519), .Z(n7521) );
  NAND U7975 ( .A(n7521), .B(n7520), .Z(n7525) );
  NANDN U7976 ( .A(n7523), .B(n7522), .Z(n7524) );
  NAND U7977 ( .A(n7525), .B(n7524), .Z(n7718) );
  XNOR U7978 ( .A(n7719), .B(n7718), .Z(n7721) );
  XNOR U7979 ( .A(n7721), .B(n7720), .Z(n7726) );
  OR U7980 ( .A(n7534), .B(n565), .Z(n7536) );
  XNOR U7981 ( .A(b[27]), .B(a[37]), .Z(n7634) );
  OR U7982 ( .A(n7634), .B(n9692), .Z(n7535) );
  AND U7983 ( .A(n7536), .B(n7535), .Z(n7713) );
  OR U7984 ( .A(n7537), .B(n561), .Z(n7539) );
  XNOR U7985 ( .A(a[59]), .B(b[5]), .Z(n7637) );
  OR U7986 ( .A(n7637), .B(n8041), .Z(n7538) );
  AND U7987 ( .A(n7539), .B(n7538), .Z(n7710) );
  NAND U7988 ( .A(n9046), .B(n7540), .Z(n7542) );
  XOR U7989 ( .A(b[19]), .B(a[45]), .Z(n7640) );
  NAND U7990 ( .A(n575), .B(n7640), .Z(n7541) );
  NAND U7991 ( .A(n7542), .B(n7541), .Z(n7711) );
  XNOR U7992 ( .A(n7710), .B(n7711), .Z(n7714) );
  XNOR U7993 ( .A(n7713), .B(n7714), .Z(n7673) );
  OR U7994 ( .A(n7543), .B(n580), .Z(n7545) );
  XNOR U7995 ( .A(b[31]), .B(a[33]), .Z(n7643) );
  OR U7996 ( .A(n7643), .B(n9904), .Z(n7544) );
  AND U7997 ( .A(n7545), .B(n7544), .Z(n7659) );
  OR U7998 ( .A(n7546), .B(n560), .Z(n7548) );
  XNOR U7999 ( .A(a[61]), .B(b[3]), .Z(n7646) );
  OR U8000 ( .A(n7646), .B(n7784), .Z(n7547) );
  AND U8001 ( .A(n7548), .B(n7547), .Z(n7656) );
  NAND U8002 ( .A(n576), .B(n7549), .Z(n7551) );
  XOR U8003 ( .A(b[17]), .B(a[47]), .Z(n7649) );
  NAND U8004 ( .A(n9141), .B(n7649), .Z(n7550) );
  NAND U8005 ( .A(n7551), .B(n7550), .Z(n7657) );
  XNOR U8006 ( .A(n7656), .B(n7657), .Z(n7660) );
  XNOR U8007 ( .A(n7659), .B(n7660), .Z(n7672) );
  XNOR U8008 ( .A(n7673), .B(n7672), .Z(n7674) );
  XOR U8009 ( .A(n7675), .B(n7674), .Z(n7727) );
  XNOR U8010 ( .A(n7726), .B(n7727), .Z(n7728) );
  XNOR U8011 ( .A(n7729), .B(n7728), .Z(n7732) );
  OR U8012 ( .A(n7560), .B(n553), .Z(n7562) );
  XNOR U8013 ( .A(a[51]), .B(b[13]), .Z(n7682) );
  OR U8014 ( .A(n7682), .B(n8853), .Z(n7561) );
  AND U8015 ( .A(n7562), .B(n7561), .Z(n7666) );
  OR U8016 ( .A(n7563), .B(n562), .Z(n7565) );
  XNOR U8017 ( .A(a[53]), .B(b[11]), .Z(n7679) );
  OR U8018 ( .A(n7679), .B(n8701), .Z(n7564) );
  AND U8019 ( .A(n7565), .B(n7564), .Z(n7664) );
  OR U8020 ( .A(n7566), .B(n557), .Z(n7568) );
  XNOR U8021 ( .A(a[49]), .B(b[15]), .Z(n7685) );
  OR U8022 ( .A(n7685), .B(n9067), .Z(n7567) );
  AND U8023 ( .A(n7568), .B(n7567), .Z(n7654) );
  OR U8024 ( .A(n7569), .B(n556), .Z(n7571) );
  XNOR U8025 ( .A(b[21]), .B(a[43]), .Z(n7688) );
  OR U8026 ( .A(n7688), .B(n9480), .Z(n7570) );
  AND U8027 ( .A(n7571), .B(n7570), .Z(n7652) );
  NAND U8028 ( .A(n570), .B(n7572), .Z(n7574) );
  XOR U8029 ( .A(a[55]), .B(b[9]), .Z(n7691) );
  NAND U8030 ( .A(n8037), .B(n7691), .Z(n7573) );
  NAND U8031 ( .A(n7574), .B(n7573), .Z(n7653) );
  XNOR U8032 ( .A(n7652), .B(n7653), .Z(n7655) );
  XNOR U8033 ( .A(n7654), .B(n7655), .Z(n7665) );
  XNOR U8034 ( .A(n7664), .B(n7665), .Z(n7667) );
  XNOR U8035 ( .A(n7666), .B(n7667), .Z(n7627) );
  OR U8036 ( .A(n7575), .B(n563), .Z(n7577) );
  XNOR U8037 ( .A(b[23]), .B(a[41]), .Z(n7694) );
  OR U8038 ( .A(n7694), .B(n9605), .Z(n7576) );
  AND U8039 ( .A(n7577), .B(n7576), .Z(n7708) );
  OR U8040 ( .A(n7578), .B(n558), .Z(n7580) );
  XNOR U8041 ( .A(a[57]), .B(b[7]), .Z(n7697) );
  OR U8042 ( .A(n7697), .B(n8290), .Z(n7579) );
  AND U8043 ( .A(n7580), .B(n7579), .Z(n7706) );
  NAND U8044 ( .A(n579), .B(n7581), .Z(n7583) );
  XOR U8045 ( .A(b[25]), .B(a[39]), .Z(n7700) );
  NAND U8046 ( .A(n9364), .B(n7700), .Z(n7582) );
  NAND U8047 ( .A(n7583), .B(n7582), .Z(n7707) );
  XNOR U8048 ( .A(n7706), .B(n7707), .Z(n7709) );
  XNOR U8049 ( .A(n7708), .B(n7709), .Z(n7625) );
  NAND U8050 ( .A(b[0]), .B(a[63]), .Z(n7584) );
  XNOR U8051 ( .A(b[1]), .B(n7584), .Z(n7586) );
  NANDN U8052 ( .A(b[0]), .B(a[62]), .Z(n7585) );
  NAND U8053 ( .A(n7586), .B(n7585), .Z(n7633) );
  OR U8054 ( .A(n7587), .B(n559), .Z(n7589) );
  XNOR U8055 ( .A(b[29]), .B(a[35]), .Z(n7703) );
  OR U8056 ( .A(n7703), .B(n9796), .Z(n7588) );
  NAND U8057 ( .A(n7589), .B(n7588), .Z(n7631) );
  NAND U8058 ( .A(b[31]), .B(a[31]), .Z(n7630) );
  XOR U8059 ( .A(n7631), .B(n7630), .Z(n7632) );
  XNOR U8060 ( .A(n7633), .B(n7632), .Z(n7624) );
  XNOR U8061 ( .A(n7625), .B(n7624), .Z(n7626) );
  XNOR U8062 ( .A(n7627), .B(n7626), .Z(n7670) );
  XNOR U8063 ( .A(n7668), .B(n7669), .Z(n7671) );
  XNOR U8064 ( .A(n7670), .B(n7671), .Z(n7723) );
  XNOR U8065 ( .A(n7722), .B(n7723), .Z(n7725) );
  XNOR U8066 ( .A(n7724), .B(n7725), .Z(n7731) );
  XOR U8067 ( .A(n7731), .B(n7730), .Z(n7733) );
  XNOR U8068 ( .A(n7732), .B(n7733), .Z(n7622) );
  XNOR U8069 ( .A(n7623), .B(n7622), .Z(n7737) );
  XOR U8070 ( .A(n7736), .B(n7737), .Z(n7739) );
  XNOR U8071 ( .A(n7738), .B(n7739), .Z(n7616) );
  XNOR U8072 ( .A(n7616), .B(n7617), .Z(n7619) );
  XNOR U8073 ( .A(n7618), .B(n7619), .Z(n7611) );
  XNOR U8074 ( .A(sreg[95]), .B(n7611), .Z(n7613) );
  NANDN U8075 ( .A(sreg[94]), .B(n7606), .Z(n7610) );
  NAND U8076 ( .A(n7608), .B(n7607), .Z(n7609) );
  NAND U8077 ( .A(n7610), .B(n7609), .Z(n7612) );
  XNOR U8078 ( .A(n7613), .B(n7612), .Z(c[95]) );
  NANDN U8079 ( .A(sreg[95]), .B(n7611), .Z(n7615) );
  NAND U8080 ( .A(n7613), .B(n7612), .Z(n7614) );
  AND U8081 ( .A(n7615), .B(n7614), .Z(n7743) );
  NANDN U8082 ( .A(n7625), .B(n7624), .Z(n7629) );
  NANDN U8083 ( .A(n7627), .B(n7626), .Z(n7628) );
  AND U8084 ( .A(n7629), .B(n7628), .Z(n7762) );
  OR U8085 ( .A(n7634), .B(n565), .Z(n7636) );
  XNOR U8086 ( .A(b[27]), .B(a[38]), .Z(n7774) );
  OR U8087 ( .A(n7774), .B(n9692), .Z(n7635) );
  AND U8088 ( .A(n7636), .B(n7635), .Z(n7843) );
  OR U8089 ( .A(n7637), .B(n561), .Z(n7639) );
  XNOR U8090 ( .A(a[60]), .B(b[5]), .Z(n7825) );
  OR U8091 ( .A(n7825), .B(n8041), .Z(n7638) );
  AND U8092 ( .A(n7639), .B(n7638), .Z(n7841) );
  NAND U8093 ( .A(n9046), .B(n7640), .Z(n7642) );
  XOR U8094 ( .A(b[19]), .B(a[46]), .Z(n7815) );
  NAND U8095 ( .A(n575), .B(n7815), .Z(n7641) );
  NAND U8096 ( .A(n7642), .B(n7641), .Z(n7842) );
  XNOR U8097 ( .A(n7841), .B(n7842), .Z(n7844) );
  XNOR U8098 ( .A(n7843), .B(n7844), .Z(n7845) );
  OR U8099 ( .A(n7643), .B(n580), .Z(n7645) );
  XNOR U8100 ( .A(b[31]), .B(a[34]), .Z(n7831) );
  OR U8101 ( .A(n7831), .B(n9904), .Z(n7644) );
  NAND U8102 ( .A(n7645), .B(n7644), .Z(n7796) );
  OR U8103 ( .A(n7646), .B(n560), .Z(n7648) );
  XNOR U8104 ( .A(a[62]), .B(b[3]), .Z(n7783) );
  OR U8105 ( .A(n7783), .B(n7784), .Z(n7647) );
  AND U8106 ( .A(n7648), .B(n7647), .Z(n7794) );
  NANDN U8107 ( .A(n554), .B(n7649), .Z(n7651) );
  XOR U8108 ( .A(b[17]), .B(a[48]), .Z(n7787) );
  NANDN U8109 ( .A(n9195), .B(n7787), .Z(n7650) );
  NAND U8110 ( .A(n7651), .B(n7650), .Z(n7795) );
  XOR U8111 ( .A(n7794), .B(n7795), .Z(n7797) );
  XOR U8112 ( .A(n7796), .B(n7797), .Z(n7846) );
  XNOR U8113 ( .A(n7845), .B(n7846), .Z(n7848) );
  XNOR U8114 ( .A(n7847), .B(n7848), .Z(n7761) );
  IV U8115 ( .A(n7656), .Z(n7658) );
  NAND U8116 ( .A(n7658), .B(n7657), .Z(n7663) );
  IV U8117 ( .A(n7659), .Z(n7661) );
  NAND U8118 ( .A(n7661), .B(n7660), .Z(n7662) );
  NAND U8119 ( .A(n7663), .B(n7662), .Z(n7849) );
  XNOR U8120 ( .A(n7850), .B(n7849), .Z(n7852) );
  XNOR U8121 ( .A(n7852), .B(n7851), .Z(n7760) );
  XNOR U8122 ( .A(n7761), .B(n7760), .Z(n7763) );
  XNOR U8123 ( .A(n7762), .B(n7763), .Z(n7755) );
  NAND U8124 ( .A(n7673), .B(n7672), .Z(n7678) );
  IV U8125 ( .A(n7674), .Z(n7676) );
  NAND U8126 ( .A(n7676), .B(n7675), .Z(n7677) );
  AND U8127 ( .A(n7678), .B(n7677), .Z(n7756) );
  OR U8128 ( .A(n7679), .B(n562), .Z(n7681) );
  XNOR U8129 ( .A(a[54]), .B(b[11]), .Z(n7809) );
  OR U8130 ( .A(n7809), .B(n8701), .Z(n7680) );
  AND U8131 ( .A(n7681), .B(n7680), .Z(n7800) );
  OR U8132 ( .A(n7682), .B(n553), .Z(n7684) );
  XNOR U8133 ( .A(a[52]), .B(b[13]), .Z(n7812) );
  OR U8134 ( .A(n7812), .B(n8853), .Z(n7683) );
  AND U8135 ( .A(n7684), .B(n7683), .Z(n7798) );
  OR U8136 ( .A(n7685), .B(n557), .Z(n7687) );
  XOR U8137 ( .A(a[50]), .B(b[15]), .Z(n7777) );
  NANDN U8138 ( .A(n9067), .B(n7777), .Z(n7686) );
  AND U8139 ( .A(n7687), .B(n7686), .Z(n7792) );
  OR U8140 ( .A(n7688), .B(n556), .Z(n7690) );
  XNOR U8141 ( .A(b[21]), .B(a[44]), .Z(n7822) );
  OR U8142 ( .A(n7822), .B(n9480), .Z(n7689) );
  AND U8143 ( .A(n7690), .B(n7689), .Z(n7790) );
  NAND U8144 ( .A(n570), .B(n7691), .Z(n7693) );
  XOR U8145 ( .A(a[56]), .B(b[9]), .Z(n7806) );
  NAND U8146 ( .A(n8037), .B(n7806), .Z(n7692) );
  NAND U8147 ( .A(n7693), .B(n7692), .Z(n7791) );
  XNOR U8148 ( .A(n7790), .B(n7791), .Z(n7793) );
  XNOR U8149 ( .A(n7792), .B(n7793), .Z(n7799) );
  XNOR U8150 ( .A(n7798), .B(n7799), .Z(n7801) );
  XOR U8151 ( .A(n7800), .B(n7801), .Z(n7767) );
  OR U8152 ( .A(n7694), .B(n563), .Z(n7696) );
  XOR U8153 ( .A(b[23]), .B(a[42]), .Z(n7828) );
  NANDN U8154 ( .A(n9605), .B(n7828), .Z(n7695) );
  AND U8155 ( .A(n7696), .B(n7695), .Z(n7839) );
  OR U8156 ( .A(n7697), .B(n558), .Z(n7699) );
  XOR U8157 ( .A(a[58]), .B(b[7]), .Z(n7818) );
  NANDN U8158 ( .A(n8290), .B(n7818), .Z(n7698) );
  AND U8159 ( .A(n7699), .B(n7698), .Z(n7837) );
  NAND U8160 ( .A(n579), .B(n7700), .Z(n7702) );
  XOR U8161 ( .A(b[25]), .B(a[40]), .Z(n7780) );
  NAND U8162 ( .A(n9364), .B(n7780), .Z(n7701) );
  NAND U8163 ( .A(n7702), .B(n7701), .Z(n7838) );
  XNOR U8164 ( .A(n7837), .B(n7838), .Z(n7840) );
  XOR U8165 ( .A(n7839), .B(n7840), .Z(n7765) );
  OR U8166 ( .A(n7703), .B(n559), .Z(n7705) );
  XNOR U8167 ( .A(b[29]), .B(a[36]), .Z(n7834) );
  OR U8168 ( .A(n7834), .B(n9796), .Z(n7704) );
  NAND U8169 ( .A(n7705), .B(n7704), .Z(n7771) );
  NAND U8170 ( .A(b[31]), .B(a[32]), .Z(n7770) );
  XOR U8171 ( .A(n7771), .B(n7770), .Z(n7773) );
  XOR U8172 ( .A(n7772), .B(n7773), .Z(n7764) );
  IV U8173 ( .A(n7710), .Z(n7712) );
  NAND U8174 ( .A(n7712), .B(n7711), .Z(n7717) );
  IV U8175 ( .A(n7713), .Z(n7715) );
  NAND U8176 ( .A(n7715), .B(n7714), .Z(n7716) );
  NAND U8177 ( .A(n7717), .B(n7716), .Z(n7803) );
  XNOR U8178 ( .A(n7802), .B(n7803), .Z(n7804) );
  XNOR U8179 ( .A(n7805), .B(n7804), .Z(n7757) );
  XNOR U8180 ( .A(n7756), .B(n7757), .Z(n7759) );
  XNOR U8181 ( .A(n7758), .B(n7759), .Z(n7753) );
  XNOR U8182 ( .A(n7753), .B(n7752), .Z(n7754) );
  XNOR U8183 ( .A(n7755), .B(n7754), .Z(n7750) );
  XNOR U8184 ( .A(n7749), .B(n7748), .Z(n7751) );
  XNOR U8185 ( .A(n7750), .B(n7751), .Z(n7854) );
  NANDN U8186 ( .A(n7731), .B(n7730), .Z(n7735) );
  OR U8187 ( .A(n7733), .B(n7732), .Z(n7734) );
  AND U8188 ( .A(n7735), .B(n7734), .Z(n7853) );
  XOR U8189 ( .A(n7854), .B(n7853), .Z(n7856) );
  XOR U8190 ( .A(n7855), .B(n7856), .Z(n7745) );
  NANDN U8191 ( .A(n7737), .B(n7736), .Z(n7741) );
  NANDN U8192 ( .A(n7739), .B(n7738), .Z(n7740) );
  NAND U8193 ( .A(n7741), .B(n7740), .Z(n7744) );
  XOR U8194 ( .A(n7745), .B(n7744), .Z(n7747) );
  XOR U8195 ( .A(n7746), .B(n7747), .Z(n7742) );
  XOR U8196 ( .A(n7743), .B(n7742), .Z(c[96]) );
  AND U8197 ( .A(n7743), .B(n7742), .Z(n7860) );
  XNOR U8198 ( .A(n7865), .B(n7866), .Z(n7868) );
  NAND U8199 ( .A(n7765), .B(n7764), .Z(n7769) );
  NAND U8200 ( .A(n7767), .B(n7766), .Z(n7768) );
  AND U8201 ( .A(n7769), .B(n7768), .Z(n7964) );
  OR U8202 ( .A(n7774), .B(n565), .Z(n7776) );
  XNOR U8203 ( .A(b[27]), .B(a[39]), .Z(n7937) );
  OR U8204 ( .A(n7937), .B(n9692), .Z(n7775) );
  AND U8205 ( .A(n7776), .B(n7775), .Z(n7932) );
  NAND U8206 ( .A(n573), .B(n7777), .Z(n7779) );
  XOR U8207 ( .A(a[51]), .B(b[15]), .Z(n7877) );
  NAND U8208 ( .A(n8694), .B(n7877), .Z(n7778) );
  NAND U8209 ( .A(n7779), .B(n7778), .Z(n7931) );
  XNOR U8210 ( .A(b[1]), .B(n7931), .Z(n7933) );
  XNOR U8211 ( .A(n7932), .B(n7933), .Z(n7959) );
  NANDN U8212 ( .A(n566), .B(n7780), .Z(n7782) );
  XNOR U8213 ( .A(b[25]), .B(a[41]), .Z(n7916) );
  OR U8214 ( .A(n7916), .B(n9684), .Z(n7781) );
  AND U8215 ( .A(n7782), .B(n7781), .Z(n7925) );
  OR U8216 ( .A(n7783), .B(n560), .Z(n7786) );
  XNOR U8217 ( .A(a[63]), .B(b[3]), .Z(n7949) );
  OR U8218 ( .A(n7949), .B(n7784), .Z(n7785) );
  AND U8219 ( .A(n7786), .B(n7785), .Z(n7923) );
  NAND U8220 ( .A(n576), .B(n7787), .Z(n7789) );
  XOR U8221 ( .A(b[17]), .B(a[49]), .Z(n7940) );
  NAND U8222 ( .A(n9141), .B(n7940), .Z(n7788) );
  NAND U8223 ( .A(n7789), .B(n7788), .Z(n7924) );
  XNOR U8224 ( .A(n7923), .B(n7924), .Z(n7926) );
  XNOR U8225 ( .A(n7925), .B(n7926), .Z(n7958) );
  XNOR U8226 ( .A(n7959), .B(n7958), .Z(n7960) );
  XNOR U8227 ( .A(n7961), .B(n7960), .Z(n7963) );
  XNOR U8228 ( .A(n7874), .B(n7873), .Z(n7876) );
  XNOR U8229 ( .A(n7876), .B(n7875), .Z(n7962) );
  XNOR U8230 ( .A(n7963), .B(n7962), .Z(n7965) );
  XNOR U8231 ( .A(n7964), .B(n7965), .Z(n7969) );
  NANDN U8232 ( .A(n564), .B(n7806), .Z(n7808) );
  XNOR U8233 ( .A(a[57]), .B(b[9]), .Z(n7901) );
  OR U8234 ( .A(n7901), .B(n8485), .Z(n7807) );
  AND U8235 ( .A(n7808), .B(n7807), .Z(n7929) );
  OR U8236 ( .A(n7809), .B(n562), .Z(n7811) );
  XNOR U8237 ( .A(a[55]), .B(b[11]), .Z(n7913) );
  OR U8238 ( .A(n7913), .B(n8701), .Z(n7810) );
  AND U8239 ( .A(n7811), .B(n7810), .Z(n7927) );
  OR U8240 ( .A(n7812), .B(n553), .Z(n7814) );
  XNOR U8241 ( .A(a[53]), .B(b[13]), .Z(n7910) );
  OR U8242 ( .A(n7910), .B(n8853), .Z(n7813) );
  AND U8243 ( .A(n7814), .B(n7813), .Z(n7921) );
  NANDN U8244 ( .A(n574), .B(n7815), .Z(n7817) );
  XOR U8245 ( .A(b[19]), .B(a[47]), .Z(n7946) );
  NANDN U8246 ( .A(n555), .B(n7946), .Z(n7816) );
  AND U8247 ( .A(n7817), .B(n7816), .Z(n7919) );
  NAND U8248 ( .A(n569), .B(n7818), .Z(n7821) );
  XOR U8249 ( .A(a[59]), .B(b[7]), .Z(n7904) );
  NAND U8250 ( .A(n7819), .B(n7904), .Z(n7820) );
  NAND U8251 ( .A(n7821), .B(n7820), .Z(n7920) );
  XNOR U8252 ( .A(n7919), .B(n7920), .Z(n7922) );
  XNOR U8253 ( .A(n7921), .B(n7922), .Z(n7928) );
  XNOR U8254 ( .A(n7927), .B(n7928), .Z(n7930) );
  XNOR U8255 ( .A(n7929), .B(n7930), .Z(n7955) );
  OR U8256 ( .A(n7822), .B(n556), .Z(n7824) );
  XOR U8257 ( .A(b[21]), .B(a[45]), .Z(n7907) );
  NANDN U8258 ( .A(n9480), .B(n7907), .Z(n7823) );
  AND U8259 ( .A(n7824), .B(n7823), .Z(n7893) );
  OR U8260 ( .A(n7825), .B(n561), .Z(n7827) );
  XNOR U8261 ( .A(a[61]), .B(b[5]), .Z(n7943) );
  OR U8262 ( .A(n7943), .B(n8041), .Z(n7826) );
  AND U8263 ( .A(n7827), .B(n7826), .Z(n7891) );
  NAND U8264 ( .A(n578), .B(n7828), .Z(n7830) );
  XOR U8265 ( .A(b[23]), .B(a[43]), .Z(n7934) );
  NAND U8266 ( .A(n9268), .B(n7934), .Z(n7829) );
  NAND U8267 ( .A(n7830), .B(n7829), .Z(n7892) );
  XNOR U8268 ( .A(n7891), .B(n7892), .Z(n7894) );
  XNOR U8269 ( .A(n7893), .B(n7894), .Z(n7953) );
  OR U8270 ( .A(n7831), .B(n580), .Z(n7833) );
  XOR U8271 ( .A(b[31]), .B(a[35]), .Z(n7883) );
  NANDN U8272 ( .A(n9904), .B(n7883), .Z(n7832) );
  NAND U8273 ( .A(n7833), .B(n7832), .Z(n7887) );
  AND U8274 ( .A(b[31]), .B(a[33]), .Z(n8047) );
  OR U8275 ( .A(n7834), .B(n559), .Z(n7836) );
  XNOR U8276 ( .A(b[29]), .B(a[37]), .Z(n7880) );
  OR U8277 ( .A(n7880), .B(n9796), .Z(n7835) );
  NAND U8278 ( .A(n7836), .B(n7835), .Z(n7886) );
  XOR U8279 ( .A(n8047), .B(n7886), .Z(n7888) );
  XOR U8280 ( .A(n7887), .B(n7888), .Z(n7952) );
  XNOR U8281 ( .A(n7953), .B(n7952), .Z(n7954) );
  XNOR U8282 ( .A(n7955), .B(n7954), .Z(n7871) );
  XNOR U8283 ( .A(n7869), .B(n7870), .Z(n7872) );
  XNOR U8284 ( .A(n7871), .B(n7872), .Z(n7896) );
  XOR U8285 ( .A(n7896), .B(n7895), .Z(n7898) );
  XNOR U8286 ( .A(n7897), .B(n7898), .Z(n7966) );
  XNOR U8287 ( .A(n7966), .B(n7967), .Z(n7968) );
  XNOR U8288 ( .A(n7969), .B(n7968), .Z(n7867) );
  XNOR U8289 ( .A(n7868), .B(n7867), .Z(n7970) );
  XOR U8290 ( .A(n7971), .B(n7970), .Z(n7973) );
  XOR U8291 ( .A(n7972), .B(n7973), .Z(n7862) );
  NANDN U8292 ( .A(n7854), .B(n7853), .Z(n7858) );
  NANDN U8293 ( .A(n7856), .B(n7855), .Z(n7857) );
  NAND U8294 ( .A(n7858), .B(n7857), .Z(n7861) );
  XOR U8295 ( .A(n7862), .B(n7861), .Z(n7864) );
  XOR U8296 ( .A(n7863), .B(n7864), .Z(n7859) );
  XOR U8297 ( .A(n7860), .B(n7859), .Z(c[97]) );
  AND U8298 ( .A(n7860), .B(n7859), .Z(n7975) );
  NANDN U8299 ( .A(n557), .B(n7877), .Z(n7879) );
  XNOR U8300 ( .A(a[52]), .B(b[15]), .Z(n7996) );
  OR U8301 ( .A(n7996), .B(n9067), .Z(n7878) );
  AND U8302 ( .A(n7879), .B(n7878), .Z(n8072) );
  OR U8303 ( .A(n7880), .B(n559), .Z(n7882) );
  XNOR U8304 ( .A(b[29]), .B(a[38]), .Z(n8033) );
  OR U8305 ( .A(n8033), .B(n9796), .Z(n7881) );
  AND U8306 ( .A(n7882), .B(n7881), .Z(n8070) );
  NAND U8307 ( .A(n9764), .B(n7883), .Z(n7885) );
  XOR U8308 ( .A(b[31]), .B(a[36]), .Z(n8064) );
  NAND U8309 ( .A(n584), .B(n8064), .Z(n7884) );
  NAND U8310 ( .A(n7885), .B(n7884), .Z(n8071) );
  XNOR U8311 ( .A(n8070), .B(n8071), .Z(n8073) );
  XNOR U8312 ( .A(n8072), .B(n8073), .Z(n7991) );
  IV U8313 ( .A(n8047), .Z(n8181) );
  NAND U8314 ( .A(n8181), .B(n7886), .Z(n7890) );
  NANDN U8315 ( .A(n7888), .B(n7887), .Z(n7889) );
  AND U8316 ( .A(n7890), .B(n7889), .Z(n7990) );
  XNOR U8317 ( .A(n7991), .B(n7990), .Z(n7993) );
  XNOR U8318 ( .A(n7993), .B(n7992), .Z(n7982) );
  XOR U8319 ( .A(n7983), .B(n7982), .Z(n7985) );
  XNOR U8320 ( .A(n7984), .B(n7985), .Z(n8084) );
  NANDN U8321 ( .A(n7896), .B(n7895), .Z(n7900) );
  NANDN U8322 ( .A(n7898), .B(n7897), .Z(n7899) );
  AND U8323 ( .A(n7900), .B(n7899), .Z(n8085) );
  XNOR U8324 ( .A(n8084), .B(n8085), .Z(n8087) );
  OR U8325 ( .A(n7901), .B(n564), .Z(n7903) );
  XOR U8326 ( .A(a[58]), .B(b[9]), .Z(n8036) );
  NANDN U8327 ( .A(n8485), .B(n8036), .Z(n7902) );
  AND U8328 ( .A(n7903), .B(n7902), .Z(n8017) );
  NANDN U8329 ( .A(n558), .B(n7904), .Z(n7906) );
  XNOR U8330 ( .A(a[60]), .B(b[7]), .Z(n8061) );
  OR U8331 ( .A(n8061), .B(n8290), .Z(n7905) );
  AND U8332 ( .A(n7906), .B(n7905), .Z(n8015) );
  NAND U8333 ( .A(n577), .B(n7907), .Z(n7909) );
  XOR U8334 ( .A(b[21]), .B(a[46]), .Z(n8067) );
  NAND U8335 ( .A(n9216), .B(n8067), .Z(n7908) );
  NAND U8336 ( .A(n7909), .B(n7908), .Z(n8016) );
  XNOR U8337 ( .A(n8015), .B(n8016), .Z(n8018) );
  XNOR U8338 ( .A(n8017), .B(n8018), .Z(n8027) );
  OR U8339 ( .A(n7910), .B(n553), .Z(n7912) );
  XOR U8340 ( .A(a[54]), .B(b[13]), .Z(n8002) );
  NANDN U8341 ( .A(n8853), .B(n8002), .Z(n7911) );
  NAND U8342 ( .A(n7912), .B(n7911), .Z(n8050) );
  OR U8343 ( .A(n7913), .B(n562), .Z(n7915) );
  XOR U8344 ( .A(a[56]), .B(b[11]), .Z(n8058) );
  NANDN U8345 ( .A(n8701), .B(n8058), .Z(n7914) );
  AND U8346 ( .A(n7915), .B(n7914), .Z(n8048) );
  OR U8347 ( .A(n7916), .B(n566), .Z(n7918) );
  XNOR U8348 ( .A(b[25]), .B(a[42]), .Z(n8052) );
  OR U8349 ( .A(n8052), .B(n9684), .Z(n7917) );
  NAND U8350 ( .A(n7918), .B(n7917), .Z(n8049) );
  XOR U8351 ( .A(n8048), .B(n8049), .Z(n8051) );
  XOR U8352 ( .A(n8050), .B(n8051), .Z(n8026) );
  XNOR U8353 ( .A(n8027), .B(n8026), .Z(n8029) );
  XNOR U8354 ( .A(n8029), .B(n8028), .Z(n8081) );
  XNOR U8355 ( .A(n8081), .B(n8080), .Z(n8083) );
  XOR U8356 ( .A(n8083), .B(n8082), .Z(n8089) );
  NANDN U8357 ( .A(n563), .B(n7934), .Z(n7936) );
  XNOR U8358 ( .A(b[23]), .B(a[44]), .Z(n8030) );
  OR U8359 ( .A(n8030), .B(n9605), .Z(n7935) );
  AND U8360 ( .A(n7936), .B(n7935), .Z(n8013) );
  OR U8361 ( .A(n7937), .B(n565), .Z(n7939) );
  XNOR U8362 ( .A(b[27]), .B(a[40]), .Z(n8055) );
  OR U8363 ( .A(n8055), .B(n9692), .Z(n7938) );
  AND U8364 ( .A(n7939), .B(n7938), .Z(n8011) );
  NAND U8365 ( .A(n576), .B(n7940), .Z(n7942) );
  XOR U8366 ( .A(b[17]), .B(a[50]), .Z(n7999) );
  NAND U8367 ( .A(n9141), .B(n7999), .Z(n7941) );
  NAND U8368 ( .A(n7942), .B(n7941), .Z(n8012) );
  XNOR U8369 ( .A(n8011), .B(n8012), .Z(n8014) );
  XNOR U8370 ( .A(n8013), .B(n8014), .Z(n8075) );
  OR U8371 ( .A(n7943), .B(n561), .Z(n7945) );
  XNOR U8372 ( .A(a[62]), .B(b[5]), .Z(n8040) );
  OR U8373 ( .A(n8040), .B(n8041), .Z(n7944) );
  AND U8374 ( .A(n7945), .B(n7944), .Z(n8019) );
  NAND U8375 ( .A(n9046), .B(n7946), .Z(n7948) );
  XOR U8376 ( .A(b[19]), .B(a[48]), .Z(n8044) );
  NAND U8377 ( .A(n575), .B(n8044), .Z(n7947) );
  NAND U8378 ( .A(n7948), .B(n7947), .Z(n8020) );
  XNOR U8379 ( .A(n8019), .B(n8020), .Z(n8022) );
  OR U8380 ( .A(n7949), .B(n560), .Z(n7950) );
  AND U8381 ( .A(n7951), .B(n7950), .Z(n8007) );
  NAND U8382 ( .A(b[31]), .B(a[34]), .Z(n8005) );
  XNOR U8383 ( .A(n8007), .B(n8005), .Z(n8008) );
  XNOR U8384 ( .A(n8047), .B(n8008), .Z(n8023) );
  XOR U8385 ( .A(n8022), .B(n8023), .Z(n8074) );
  XOR U8386 ( .A(n8075), .B(n8074), .Z(n8077) );
  XNOR U8387 ( .A(n8076), .B(n8077), .Z(n7986) );
  NANDN U8388 ( .A(n7953), .B(n7952), .Z(n7957) );
  NANDN U8389 ( .A(n7955), .B(n7954), .Z(n7956) );
  AND U8390 ( .A(n7957), .B(n7956), .Z(n7987) );
  XNOR U8391 ( .A(n7986), .B(n7987), .Z(n7989) );
  XNOR U8392 ( .A(n7989), .B(n7988), .Z(n8088) );
  XNOR U8393 ( .A(n8091), .B(n8090), .Z(n8086) );
  XNOR U8394 ( .A(n8087), .B(n8086), .Z(n8095) );
  XOR U8395 ( .A(n8095), .B(n8094), .Z(n8097) );
  XNOR U8396 ( .A(n8096), .B(n8097), .Z(n7977) );
  XNOR U8397 ( .A(n7977), .B(n7976), .Z(n7979) );
  XOR U8398 ( .A(n7978), .B(n7979), .Z(n7974) );
  XOR U8399 ( .A(n7975), .B(n7974), .Z(c[98]) );
  AND U8400 ( .A(n7975), .B(n7974), .Z(n8101) );
  NAND U8401 ( .A(n7977), .B(n7976), .Z(n7981) );
  NANDN U8402 ( .A(n7979), .B(n7978), .Z(n7980) );
  NAND U8403 ( .A(n7981), .B(n7980), .Z(n8104) );
  XNOR U8404 ( .A(n8110), .B(n8111), .Z(n8113) );
  NANDN U8405 ( .A(n7991), .B(n7990), .Z(n7995) );
  NAND U8406 ( .A(n7993), .B(n7992), .Z(n7994) );
  AND U8407 ( .A(n7995), .B(n7994), .Z(n8199) );
  OR U8408 ( .A(n7996), .B(n557), .Z(n7998) );
  XNOR U8409 ( .A(a[53]), .B(b[15]), .Z(n8170) );
  OR U8410 ( .A(n8170), .B(n9067), .Z(n7997) );
  AND U8411 ( .A(n7998), .B(n7997), .Z(n8187) );
  NANDN U8412 ( .A(n554), .B(n7999), .Z(n8001) );
  XNOR U8413 ( .A(a[51]), .B(b[17]), .Z(n8173) );
  OR U8414 ( .A(n8173), .B(n9195), .Z(n8000) );
  AND U8415 ( .A(n8001), .B(n8000), .Z(n8185) );
  NAND U8416 ( .A(n572), .B(n8002), .Z(n8004) );
  XOR U8417 ( .A(a[55]), .B(b[13]), .Z(n8176) );
  NAND U8418 ( .A(n8585), .B(n8176), .Z(n8003) );
  NAND U8419 ( .A(n8004), .B(n8003), .Z(n8186) );
  XNOR U8420 ( .A(n8185), .B(n8186), .Z(n8188) );
  XNOR U8421 ( .A(n8187), .B(n8188), .Z(n8125) );
  IV U8422 ( .A(n8005), .Z(n8006) );
  NANDN U8423 ( .A(n8007), .B(n8006), .Z(n8010) );
  OR U8424 ( .A(n8008), .B(n8047), .Z(n8009) );
  AND U8425 ( .A(n8010), .B(n8009), .Z(n8124) );
  XNOR U8426 ( .A(n8125), .B(n8124), .Z(n8127) );
  XNOR U8427 ( .A(n8127), .B(n8126), .Z(n8204) );
  IV U8428 ( .A(n8019), .Z(n8021) );
  NAND U8429 ( .A(n8021), .B(n8020), .Z(n8025) );
  NANDN U8430 ( .A(n8023), .B(n8022), .Z(n8024) );
  NAND U8431 ( .A(n8025), .B(n8024), .Z(n8202) );
  XNOR U8432 ( .A(n8201), .B(n8202), .Z(n8203) );
  XNOR U8433 ( .A(n8204), .B(n8203), .Z(n8197) );
  XNOR U8434 ( .A(n8197), .B(n8198), .Z(n8200) );
  XNOR U8435 ( .A(n8199), .B(n8200), .Z(n8117) );
  OR U8436 ( .A(n8030), .B(n563), .Z(n8032) );
  XNOR U8437 ( .A(b[23]), .B(a[45]), .Z(n8128) );
  OR U8438 ( .A(n8128), .B(n9605), .Z(n8031) );
  AND U8439 ( .A(n8032), .B(n8031), .Z(n8168) );
  OR U8440 ( .A(n8033), .B(n559), .Z(n8035) );
  XNOR U8441 ( .A(b[29]), .B(a[39]), .Z(n8141) );
  OR U8442 ( .A(n8141), .B(n9796), .Z(n8034) );
  AND U8443 ( .A(n8035), .B(n8034), .Z(n8166) );
  NAND U8444 ( .A(n570), .B(n8036), .Z(n8039) );
  XOR U8445 ( .A(a[59]), .B(b[9]), .Z(n8154) );
  NAND U8446 ( .A(n8037), .B(n8154), .Z(n8038) );
  NAND U8447 ( .A(n8039), .B(n8038), .Z(n8167) );
  XNOR U8448 ( .A(n8166), .B(n8167), .Z(n8169) );
  XNOR U8449 ( .A(n8168), .B(n8169), .Z(n8206) );
  OR U8450 ( .A(n8040), .B(n561), .Z(n8043) );
  XNOR U8451 ( .A(a[63]), .B(b[5]), .Z(n8163) );
  OR U8452 ( .A(n8163), .B(n8041), .Z(n8042) );
  AND U8453 ( .A(n8043), .B(n8042), .Z(n8193) );
  NAND U8454 ( .A(n9046), .B(n8044), .Z(n8046) );
  XOR U8455 ( .A(b[19]), .B(a[49]), .Z(n8144) );
  NAND U8456 ( .A(n575), .B(n8144), .Z(n8045) );
  NAND U8457 ( .A(n8046), .B(n8045), .Z(n8194) );
  XNOR U8458 ( .A(n8193), .B(n8194), .Z(n8196) );
  AND U8459 ( .A(b[31]), .B(a[35]), .Z(n8179) );
  XNOR U8460 ( .A(n8180), .B(n8179), .Z(n8182) );
  XNOR U8461 ( .A(n8047), .B(n8182), .Z(n8195) );
  XNOR U8462 ( .A(n8196), .B(n8195), .Z(n8205) );
  XNOR U8463 ( .A(n8206), .B(n8205), .Z(n8208) );
  XNOR U8464 ( .A(n8208), .B(n8207), .Z(n8121) );
  OR U8465 ( .A(n8052), .B(n566), .Z(n8054) );
  XNOR U8466 ( .A(b[25]), .B(a[43]), .Z(n8131) );
  OR U8467 ( .A(n8131), .B(n9684), .Z(n8053) );
  AND U8468 ( .A(n8054), .B(n8053), .Z(n8149) );
  OR U8469 ( .A(n8055), .B(n565), .Z(n8057) );
  XNOR U8470 ( .A(b[27]), .B(a[41]), .Z(n8151) );
  OR U8471 ( .A(n8151), .B(n9692), .Z(n8056) );
  AND U8472 ( .A(n8057), .B(n8056), .Z(n8147) );
  NAND U8473 ( .A(n571), .B(n8058), .Z(n8060) );
  XOR U8474 ( .A(a[57]), .B(b[11]), .Z(n8134) );
  NAND U8475 ( .A(n8135), .B(n8134), .Z(n8059) );
  NAND U8476 ( .A(n8060), .B(n8059), .Z(n8148) );
  XNOR U8477 ( .A(n8147), .B(n8148), .Z(n8150) );
  XNOR U8478 ( .A(n8149), .B(n8150), .Z(n8210) );
  OR U8479 ( .A(n8061), .B(n558), .Z(n8063) );
  XNOR U8480 ( .A(a[61]), .B(b[7]), .Z(n8138) );
  OR U8481 ( .A(n8138), .B(n8290), .Z(n8062) );
  NAND U8482 ( .A(n8063), .B(n8062), .Z(n8191) );
  NANDN U8483 ( .A(n580), .B(n8064), .Z(n8066) );
  XNOR U8484 ( .A(b[31]), .B(a[37]), .Z(n8160) );
  OR U8485 ( .A(n8160), .B(n9904), .Z(n8065) );
  AND U8486 ( .A(n8066), .B(n8065), .Z(n8189) );
  NANDN U8487 ( .A(n556), .B(n8067), .Z(n8069) );
  XOR U8488 ( .A(b[21]), .B(a[47]), .Z(n8157) );
  NANDN U8489 ( .A(n9480), .B(n8157), .Z(n8068) );
  NAND U8490 ( .A(n8069), .B(n8068), .Z(n8190) );
  XOR U8491 ( .A(n8189), .B(n8190), .Z(n8192) );
  XOR U8492 ( .A(n8191), .B(n8192), .Z(n8209) );
  XNOR U8493 ( .A(n8210), .B(n8209), .Z(n8212) );
  XNOR U8494 ( .A(n8212), .B(n8211), .Z(n8120) );
  XNOR U8495 ( .A(n8121), .B(n8120), .Z(n8123) );
  NANDN U8496 ( .A(n8075), .B(n8074), .Z(n8079) );
  NANDN U8497 ( .A(n8077), .B(n8076), .Z(n8078) );
  NAND U8498 ( .A(n8079), .B(n8078), .Z(n8122) );
  XNOR U8499 ( .A(n8123), .B(n8122), .Z(n8115) );
  XNOR U8500 ( .A(n8115), .B(n8114), .Z(n8116) );
  XNOR U8501 ( .A(n8117), .B(n8116), .Z(n8112) );
  XNOR U8502 ( .A(n8113), .B(n8112), .Z(n8109) );
  NAND U8503 ( .A(n8089), .B(n8088), .Z(n8093) );
  NAND U8504 ( .A(n8091), .B(n8090), .Z(n8092) );
  NAND U8505 ( .A(n8093), .B(n8092), .Z(n8107) );
  XNOR U8506 ( .A(n8106), .B(n8107), .Z(n8108) );
  XNOR U8507 ( .A(n8109), .B(n8108), .Z(n8102) );
  NANDN U8508 ( .A(n8095), .B(n8094), .Z(n8099) );
  NANDN U8509 ( .A(n8097), .B(n8096), .Z(n8098) );
  NAND U8510 ( .A(n8099), .B(n8098), .Z(n8103) );
  XOR U8511 ( .A(n8102), .B(n8103), .Z(n8105) );
  XOR U8512 ( .A(n8104), .B(n8105), .Z(n8100) );
  XOR U8513 ( .A(n8101), .B(n8100), .Z(c[99]) );
  AND U8514 ( .A(n8101), .B(n8100), .Z(n8216) );
  NANDN U8515 ( .A(n8115), .B(n8114), .Z(n8119) );
  NAND U8516 ( .A(n8117), .B(n8116), .Z(n8118) );
  AND U8517 ( .A(n8119), .B(n8118), .Z(n8223) );
  OR U8518 ( .A(n8128), .B(n563), .Z(n8130) );
  XNOR U8519 ( .A(b[23]), .B(a[46]), .Z(n8261) );
  OR U8520 ( .A(n8261), .B(n9605), .Z(n8129) );
  AND U8521 ( .A(n8130), .B(n8129), .Z(n8313) );
  OR U8522 ( .A(n8131), .B(n566), .Z(n8133) );
  XNOR U8523 ( .A(b[25]), .B(a[44]), .Z(n8305) );
  OR U8524 ( .A(n8305), .B(n9684), .Z(n8132) );
  AND U8525 ( .A(n8133), .B(n8132), .Z(n8311) );
  NAND U8526 ( .A(n571), .B(n8134), .Z(n8137) );
  XOR U8527 ( .A(a[58]), .B(b[11]), .Z(n8308) );
  NAND U8528 ( .A(n8135), .B(n8308), .Z(n8136) );
  NAND U8529 ( .A(n8137), .B(n8136), .Z(n8312) );
  XNOR U8530 ( .A(n8311), .B(n8312), .Z(n8314) );
  XNOR U8531 ( .A(n8313), .B(n8314), .Z(n8236) );
  OR U8532 ( .A(n8138), .B(n558), .Z(n8140) );
  XNOR U8533 ( .A(a[62]), .B(b[7]), .Z(n8289) );
  OR U8534 ( .A(n8289), .B(n8290), .Z(n8139) );
  NAND U8535 ( .A(n8140), .B(n8139), .Z(n8284) );
  OR U8536 ( .A(n8141), .B(n559), .Z(n8143) );
  XNOR U8537 ( .A(b[29]), .B(a[40]), .Z(n8286) );
  OR U8538 ( .A(n8286), .B(n9796), .Z(n8142) );
  AND U8539 ( .A(n8143), .B(n8142), .Z(n8282) );
  NANDN U8540 ( .A(n574), .B(n8144), .Z(n8146) );
  XOR U8541 ( .A(b[19]), .B(a[50]), .Z(n8273) );
  NANDN U8542 ( .A(n555), .B(n8273), .Z(n8145) );
  NAND U8543 ( .A(n8146), .B(n8145), .Z(n8283) );
  XOR U8544 ( .A(n8282), .B(n8283), .Z(n8285) );
  XOR U8545 ( .A(n8284), .B(n8285), .Z(n8235) );
  XNOR U8546 ( .A(n8236), .B(n8235), .Z(n8238) );
  XNOR U8547 ( .A(n8238), .B(n8237), .Z(n8250) );
  OR U8548 ( .A(n8151), .B(n565), .Z(n8153) );
  XOR U8549 ( .A(b[27]), .B(a[42]), .Z(n8267) );
  NANDN U8550 ( .A(n9692), .B(n8267), .Z(n8152) );
  AND U8551 ( .A(n8153), .B(n8152), .Z(n8255) );
  NANDN U8552 ( .A(n564), .B(n8154), .Z(n8156) );
  XNOR U8553 ( .A(a[60]), .B(b[9]), .Z(n8264) );
  OR U8554 ( .A(n8264), .B(n8485), .Z(n8155) );
  AND U8555 ( .A(n8156), .B(n8155), .Z(n8253) );
  NAND U8556 ( .A(n577), .B(n8157), .Z(n8159) );
  XOR U8557 ( .A(b[21]), .B(a[48]), .Z(n8293) );
  NAND U8558 ( .A(n9216), .B(n8293), .Z(n8158) );
  NAND U8559 ( .A(n8159), .B(n8158), .Z(n8254) );
  XNOR U8560 ( .A(n8253), .B(n8254), .Z(n8256) );
  XNOR U8561 ( .A(n8255), .B(n8256), .Z(n8240) );
  OR U8562 ( .A(n8160), .B(n580), .Z(n8162) );
  XNOR U8563 ( .A(b[31]), .B(a[38]), .Z(n8270) );
  OR U8564 ( .A(n8270), .B(n9904), .Z(n8161) );
  NAND U8565 ( .A(n8162), .B(n8161), .Z(n8278) );
  AND U8566 ( .A(b[31]), .B(a[36]), .Z(n8276) );
  OR U8567 ( .A(n8163), .B(n561), .Z(n8164) );
  AND U8568 ( .A(n8165), .B(n8164), .Z(n8277) );
  XNOR U8569 ( .A(n8276), .B(n8277), .Z(n8279) );
  XOR U8570 ( .A(n8278), .B(n8279), .Z(n8239) );
  XNOR U8571 ( .A(n8240), .B(n8239), .Z(n8242) );
  XNOR U8572 ( .A(n8242), .B(n8241), .Z(n8249) );
  XNOR U8573 ( .A(n8250), .B(n8249), .Z(n8252) );
  XNOR U8574 ( .A(n8251), .B(n8252), .Z(n8228) );
  OR U8575 ( .A(n8170), .B(n557), .Z(n8172) );
  XNOR U8576 ( .A(a[54]), .B(b[15]), .Z(n8296) );
  OR U8577 ( .A(n8296), .B(n9067), .Z(n8171) );
  AND U8578 ( .A(n8172), .B(n8171), .Z(n8259) );
  OR U8579 ( .A(n8173), .B(n554), .Z(n8175) );
  XNOR U8580 ( .A(a[52]), .B(b[17]), .Z(n8302) );
  OR U8581 ( .A(n8302), .B(n9195), .Z(n8174) );
  AND U8582 ( .A(n8175), .B(n8174), .Z(n8257) );
  NAND U8583 ( .A(n572), .B(n8176), .Z(n8178) );
  XOR U8584 ( .A(a[56]), .B(b[13]), .Z(n8299) );
  NAND U8585 ( .A(n8585), .B(n8299), .Z(n8177) );
  NAND U8586 ( .A(n8178), .B(n8177), .Z(n8258) );
  XNOR U8587 ( .A(n8257), .B(n8258), .Z(n8260) );
  XOR U8588 ( .A(n8259), .B(n8260), .Z(n8316) );
  NAND U8589 ( .A(n8180), .B(n8179), .Z(n8184) );
  OR U8590 ( .A(n8182), .B(n8181), .Z(n8183) );
  AND U8591 ( .A(n8184), .B(n8183), .Z(n8315) );
  XOR U8592 ( .A(n8318), .B(n8317), .Z(n8234) );
  XNOR U8593 ( .A(n8231), .B(n8232), .Z(n8233) );
  XNOR U8594 ( .A(n8234), .B(n8233), .Z(n8227) );
  XNOR U8595 ( .A(n8228), .B(n8227), .Z(n8230) );
  XNOR U8596 ( .A(n8229), .B(n8230), .Z(n8324) );
  NANDN U8597 ( .A(n8210), .B(n8209), .Z(n8214) );
  NAND U8598 ( .A(n8212), .B(n8211), .Z(n8213) );
  NAND U8599 ( .A(n8214), .B(n8213), .Z(n8246) );
  XOR U8600 ( .A(n8245), .B(n8246), .Z(n8248) );
  XNOR U8601 ( .A(n8247), .B(n8248), .Z(n8322) );
  XNOR U8602 ( .A(n8321), .B(n8322), .Z(n8323) );
  XNOR U8603 ( .A(n8324), .B(n8323), .Z(n8224) );
  XNOR U8604 ( .A(n8223), .B(n8224), .Z(n8226) );
  XNOR U8605 ( .A(n8225), .B(n8226), .Z(n8217) );
  XNOR U8606 ( .A(n8218), .B(n8217), .Z(n8220) );
  XOR U8607 ( .A(n8219), .B(n8220), .Z(n8215) );
  XOR U8608 ( .A(n8216), .B(n8215), .Z(c[100]) );
  AND U8609 ( .A(n8216), .B(n8215), .Z(n8326) );
  NAND U8610 ( .A(n8218), .B(n8217), .Z(n8222) );
  NANDN U8611 ( .A(n8220), .B(n8219), .Z(n8221) );
  NAND U8612 ( .A(n8222), .B(n8221), .Z(n8329) );
  NANDN U8613 ( .A(n8240), .B(n8239), .Z(n8244) );
  NAND U8614 ( .A(n8242), .B(n8241), .Z(n8243) );
  NAND U8615 ( .A(n8244), .B(n8243), .Z(n8338) );
  XOR U8616 ( .A(n8337), .B(n8338), .Z(n8340) );
  XNOR U8617 ( .A(n8339), .B(n8340), .Z(n8333) );
  XNOR U8618 ( .A(n8333), .B(n8334), .Z(n8336) );
  XNOR U8619 ( .A(n8335), .B(n8336), .Z(n8431) );
  XNOR U8620 ( .A(n8371), .B(n8370), .Z(n8373) );
  OR U8621 ( .A(n8261), .B(n563), .Z(n8263) );
  XNOR U8622 ( .A(b[23]), .B(a[47]), .Z(n8384) );
  OR U8623 ( .A(n8384), .B(n9605), .Z(n8262) );
  AND U8624 ( .A(n8263), .B(n8262), .Z(n8353) );
  OR U8625 ( .A(n8264), .B(n564), .Z(n8266) );
  XNOR U8626 ( .A(a[61]), .B(b[9]), .Z(n8402) );
  OR U8627 ( .A(n8402), .B(n8485), .Z(n8265) );
  AND U8628 ( .A(n8266), .B(n8265), .Z(n8351) );
  NAND U8629 ( .A(n582), .B(n8267), .Z(n8269) );
  XOR U8630 ( .A(b[27]), .B(a[43]), .Z(n8390) );
  NAND U8631 ( .A(n9770), .B(n8390), .Z(n8268) );
  NAND U8632 ( .A(n8269), .B(n8268), .Z(n8352) );
  XNOR U8633 ( .A(n8351), .B(n8352), .Z(n8354) );
  XNOR U8634 ( .A(n8353), .B(n8354), .Z(n8379) );
  OR U8635 ( .A(n8270), .B(n580), .Z(n8272) );
  XNOR U8636 ( .A(b[31]), .B(a[39]), .Z(n8408) );
  OR U8637 ( .A(n8408), .B(n9904), .Z(n8271) );
  AND U8638 ( .A(n8272), .B(n8271), .Z(n8414) );
  NAND U8639 ( .A(n9046), .B(n8273), .Z(n8275) );
  XOR U8640 ( .A(b[19]), .B(a[51]), .Z(n8387) );
  NAND U8641 ( .A(n575), .B(n8387), .Z(n8274) );
  NAND U8642 ( .A(n8275), .B(n8274), .Z(n8415) );
  XNOR U8643 ( .A(n8414), .B(n8415), .Z(n8417) );
  AND U8644 ( .A(b[31]), .B(a[37]), .Z(n8364) );
  XOR U8645 ( .A(n8364), .B(n8365), .Z(n8367) );
  XNOR U8646 ( .A(n8276), .B(n8367), .Z(n8416) );
  XNOR U8647 ( .A(n8417), .B(n8416), .Z(n8378) );
  XNOR U8648 ( .A(n8379), .B(n8378), .Z(n8381) );
  IV U8649 ( .A(n8276), .Z(n8366) );
  NANDN U8650 ( .A(n8277), .B(n8366), .Z(n8281) );
  NANDN U8651 ( .A(n8279), .B(n8278), .Z(n8280) );
  AND U8652 ( .A(n8281), .B(n8280), .Z(n8380) );
  XNOR U8653 ( .A(n8381), .B(n8380), .Z(n8372) );
  XNOR U8654 ( .A(n8373), .B(n8372), .Z(n8424) );
  OR U8655 ( .A(n8286), .B(n559), .Z(n8288) );
  XNOR U8656 ( .A(b[29]), .B(a[41]), .Z(n8393) );
  OR U8657 ( .A(n8393), .B(n9796), .Z(n8287) );
  AND U8658 ( .A(n8288), .B(n8287), .Z(n8349) );
  OR U8659 ( .A(n8289), .B(n558), .Z(n8292) );
  XNOR U8660 ( .A(a[63]), .B(b[7]), .Z(n8411) );
  OR U8661 ( .A(n8411), .B(n8290), .Z(n8291) );
  AND U8662 ( .A(n8292), .B(n8291), .Z(n8347) );
  NAND U8663 ( .A(n577), .B(n8293), .Z(n8295) );
  XOR U8664 ( .A(b[21]), .B(a[49]), .Z(n8405) );
  NAND U8665 ( .A(n9216), .B(n8405), .Z(n8294) );
  NAND U8666 ( .A(n8295), .B(n8294), .Z(n8348) );
  XNOR U8667 ( .A(n8347), .B(n8348), .Z(n8350) );
  XNOR U8668 ( .A(n8349), .B(n8350), .Z(n8375) );
  XNOR U8669 ( .A(n8374), .B(n8375), .Z(n8376) );
  OR U8670 ( .A(n8296), .B(n557), .Z(n8298) );
  XNOR U8671 ( .A(a[55]), .B(b[15]), .Z(n8355) );
  OR U8672 ( .A(n8355), .B(n9067), .Z(n8297) );
  NAND U8673 ( .A(n8298), .B(n8297), .Z(n8343) );
  NANDN U8674 ( .A(n553), .B(n8299), .Z(n8301) );
  XNOR U8675 ( .A(a[57]), .B(b[13]), .Z(n8358) );
  OR U8676 ( .A(n8358), .B(n8853), .Z(n8300) );
  NAND U8677 ( .A(n8301), .B(n8300), .Z(n8341) );
  OR U8678 ( .A(n8302), .B(n554), .Z(n8304) );
  XOR U8679 ( .A(a[53]), .B(b[17]), .Z(n8396) );
  NANDN U8680 ( .A(n9195), .B(n8396), .Z(n8303) );
  NAND U8681 ( .A(n8304), .B(n8303), .Z(n8420) );
  OR U8682 ( .A(n8305), .B(n566), .Z(n8307) );
  XOR U8683 ( .A(b[25]), .B(a[45]), .Z(n8361) );
  NANDN U8684 ( .A(n9684), .B(n8361), .Z(n8306) );
  AND U8685 ( .A(n8307), .B(n8306), .Z(n8418) );
  NANDN U8686 ( .A(n562), .B(n8308), .Z(n8310) );
  XNOR U8687 ( .A(a[59]), .B(b[11]), .Z(n8399) );
  OR U8688 ( .A(n8399), .B(n8701), .Z(n8309) );
  NAND U8689 ( .A(n8310), .B(n8309), .Z(n8419) );
  XOR U8690 ( .A(n8418), .B(n8419), .Z(n8421) );
  XOR U8691 ( .A(n8420), .B(n8421), .Z(n8342) );
  XOR U8692 ( .A(n8341), .B(n8342), .Z(n8344) );
  XOR U8693 ( .A(n8343), .B(n8344), .Z(n8377) );
  XOR U8694 ( .A(n8376), .B(n8377), .Z(n8423) );
  XOR U8695 ( .A(n8423), .B(n8422), .Z(n8425) );
  XNOR U8696 ( .A(n8424), .B(n8425), .Z(n8426) );
  NAND U8697 ( .A(n8316), .B(n8315), .Z(n8320) );
  NAND U8698 ( .A(n8318), .B(n8317), .Z(n8319) );
  AND U8699 ( .A(n8320), .B(n8319), .Z(n8427) );
  XNOR U8700 ( .A(n8426), .B(n8427), .Z(n8428) );
  XNOR U8701 ( .A(n8429), .B(n8428), .Z(n8430) );
  XNOR U8702 ( .A(n8431), .B(n8430), .Z(n8433) );
  XNOR U8703 ( .A(n8433), .B(n8432), .Z(n8328) );
  XOR U8704 ( .A(n8327), .B(n8328), .Z(n8330) );
  XOR U8705 ( .A(n8329), .B(n8330), .Z(n8325) );
  XOR U8706 ( .A(n8326), .B(n8325), .Z(c[101]) );
  AND U8707 ( .A(n8326), .B(n8325), .Z(n8435) );
  NANDN U8708 ( .A(n8328), .B(n8327), .Z(n8332) );
  NANDN U8709 ( .A(n8330), .B(n8329), .Z(n8331) );
  NAND U8710 ( .A(n8332), .B(n8331), .Z(n8438) );
  NANDN U8711 ( .A(n8342), .B(n8341), .Z(n8346) );
  NANDN U8712 ( .A(n8344), .B(n8343), .Z(n8345) );
  AND U8713 ( .A(n8346), .B(n8345), .Z(n8445) );
  OR U8714 ( .A(n8355), .B(n557), .Z(n8357) );
  XOR U8715 ( .A(a[56]), .B(b[15]), .Z(n8468) );
  NANDN U8716 ( .A(n9067), .B(n8468), .Z(n8356) );
  AND U8717 ( .A(n8357), .B(n8356), .Z(n8448) );
  OR U8718 ( .A(n8358), .B(n553), .Z(n8360) );
  XOR U8719 ( .A(a[58]), .B(b[13]), .Z(n8465) );
  NANDN U8720 ( .A(n8853), .B(n8465), .Z(n8359) );
  AND U8721 ( .A(n8360), .B(n8359), .Z(n8446) );
  NAND U8722 ( .A(n579), .B(n8361), .Z(n8363) );
  XOR U8723 ( .A(b[25]), .B(a[46]), .Z(n8456) );
  NAND U8724 ( .A(n9364), .B(n8456), .Z(n8362) );
  NAND U8725 ( .A(n8363), .B(n8362), .Z(n8447) );
  XNOR U8726 ( .A(n8446), .B(n8447), .Z(n8449) );
  XNOR U8727 ( .A(n8448), .B(n8449), .Z(n8515) );
  NANDN U8728 ( .A(n8365), .B(n8364), .Z(n8369) );
  OR U8729 ( .A(n8367), .B(n8366), .Z(n8368) );
  AND U8730 ( .A(n8369), .B(n8368), .Z(n8514) );
  XOR U8731 ( .A(n8515), .B(n8514), .Z(n8517) );
  XNOR U8732 ( .A(n8516), .B(n8517), .Z(n8442) );
  XNOR U8733 ( .A(n8443), .B(n8442), .Z(n8444) );
  XNOR U8734 ( .A(n8445), .B(n8444), .Z(n8527) );
  XNOR U8735 ( .A(n8527), .B(n8526), .Z(n8528) );
  NANDN U8736 ( .A(n8379), .B(n8378), .Z(n8383) );
  NAND U8737 ( .A(n8381), .B(n8380), .Z(n8382) );
  AND U8738 ( .A(n8383), .B(n8382), .Z(n8507) );
  OR U8739 ( .A(n8384), .B(n563), .Z(n8386) );
  XOR U8740 ( .A(b[23]), .B(a[48]), .Z(n8481) );
  NANDN U8741 ( .A(n9605), .B(n8481), .Z(n8385) );
  AND U8742 ( .A(n8386), .B(n8385), .Z(n8473) );
  NANDN U8743 ( .A(n574), .B(n8387), .Z(n8389) );
  XNOR U8744 ( .A(a[52]), .B(b[19]), .Z(n8462) );
  OR U8745 ( .A(n8462), .B(n555), .Z(n8388) );
  AND U8746 ( .A(n8389), .B(n8388), .Z(n8471) );
  NANDN U8747 ( .A(n565), .B(n8390), .Z(n8392) );
  XNOR U8748 ( .A(b[27]), .B(a[44]), .Z(n8450) );
  OR U8749 ( .A(n8450), .B(n9692), .Z(n8391) );
  AND U8750 ( .A(n8392), .B(n8391), .Z(n8504) );
  OR U8751 ( .A(n8393), .B(n559), .Z(n8395) );
  XNOR U8752 ( .A(b[29]), .B(a[42]), .Z(n8475) );
  OR U8753 ( .A(n8475), .B(n9796), .Z(n8394) );
  AND U8754 ( .A(n8395), .B(n8394), .Z(n8502) );
  NAND U8755 ( .A(n576), .B(n8396), .Z(n8398) );
  XOR U8756 ( .A(a[54]), .B(b[17]), .Z(n8459) );
  NAND U8757 ( .A(n9141), .B(n8459), .Z(n8397) );
  NAND U8758 ( .A(n8398), .B(n8397), .Z(n8503) );
  XNOR U8759 ( .A(n8502), .B(n8503), .Z(n8505) );
  XNOR U8760 ( .A(n8504), .B(n8505), .Z(n8472) );
  XNOR U8761 ( .A(n8471), .B(n8472), .Z(n8474) );
  XNOR U8762 ( .A(n8473), .B(n8474), .Z(n8523) );
  OR U8763 ( .A(n8399), .B(n562), .Z(n8401) );
  XNOR U8764 ( .A(a[60]), .B(b[11]), .Z(n8453) );
  OR U8765 ( .A(n8453), .B(n8701), .Z(n8400) );
  AND U8766 ( .A(n8401), .B(n8400), .Z(n8500) );
  OR U8767 ( .A(n8402), .B(n564), .Z(n8404) );
  XNOR U8768 ( .A(a[62]), .B(b[9]), .Z(n8484) );
  OR U8769 ( .A(n8484), .B(n8485), .Z(n8403) );
  AND U8770 ( .A(n8404), .B(n8403), .Z(n8498) );
  NAND U8771 ( .A(n577), .B(n8405), .Z(n8407) );
  XOR U8772 ( .A(b[21]), .B(a[50]), .Z(n8488) );
  NAND U8773 ( .A(n9216), .B(n8488), .Z(n8406) );
  NAND U8774 ( .A(n8407), .B(n8406), .Z(n8499) );
  XNOR U8775 ( .A(n8498), .B(n8499), .Z(n8501) );
  XNOR U8776 ( .A(n8500), .B(n8501), .Z(n8521) );
  OR U8777 ( .A(n8408), .B(n580), .Z(n8410) );
  XNOR U8778 ( .A(b[31]), .B(a[40]), .Z(n8478) );
  OR U8779 ( .A(n8478), .B(n9904), .Z(n8409) );
  NAND U8780 ( .A(n8410), .B(n8409), .Z(n8494) );
  AND U8781 ( .A(b[31]), .B(a[38]), .Z(n8492) );
  OR U8782 ( .A(n8411), .B(n558), .Z(n8412) );
  AND U8783 ( .A(n8413), .B(n8412), .Z(n8493) );
  XNOR U8784 ( .A(n8492), .B(n8493), .Z(n8495) );
  XOR U8785 ( .A(n8494), .B(n8495), .Z(n8520) );
  XNOR U8786 ( .A(n8521), .B(n8520), .Z(n8522) );
  XNOR U8787 ( .A(n8523), .B(n8522), .Z(n8512) );
  XNOR U8788 ( .A(n8510), .B(n8511), .Z(n8513) );
  XNOR U8789 ( .A(n8512), .B(n8513), .Z(n8506) );
  XNOR U8790 ( .A(n8507), .B(n8506), .Z(n8508) );
  XOR U8791 ( .A(n8509), .B(n8508), .Z(n8529) );
  XNOR U8792 ( .A(n8528), .B(n8529), .Z(n8532) );
  XNOR U8793 ( .A(n8532), .B(n8533), .Z(n8535) );
  XNOR U8794 ( .A(n8534), .B(n8535), .Z(n8537) );
  XNOR U8795 ( .A(n8537), .B(n8536), .Z(n8539) );
  XNOR U8796 ( .A(n8538), .B(n8539), .Z(n8437) );
  XOR U8797 ( .A(n8437), .B(n8436), .Z(n8439) );
  XOR U8798 ( .A(n8438), .B(n8439), .Z(n8434) );
  XOR U8799 ( .A(n8435), .B(n8434), .Z(c[102]) );
  AND U8800 ( .A(n8435), .B(n8434), .Z(n8541) );
  NANDN U8801 ( .A(n8437), .B(n8436), .Z(n8441) );
  NANDN U8802 ( .A(n8439), .B(n8438), .Z(n8440) );
  NAND U8803 ( .A(n8441), .B(n8440), .Z(n8544) );
  OR U8804 ( .A(n8450), .B(n565), .Z(n8452) );
  XNOR U8805 ( .A(b[27]), .B(a[45]), .Z(n8572) );
  OR U8806 ( .A(n8572), .B(n9692), .Z(n8451) );
  AND U8807 ( .A(n8452), .B(n8451), .Z(n8597) );
  OR U8808 ( .A(n8453), .B(n562), .Z(n8455) );
  XNOR U8809 ( .A(a[61]), .B(b[11]), .Z(n8552) );
  OR U8810 ( .A(n8552), .B(n8701), .Z(n8454) );
  AND U8811 ( .A(n8455), .B(n8454), .Z(n8595) );
  NAND U8812 ( .A(n579), .B(n8456), .Z(n8458) );
  XOR U8813 ( .A(b[25]), .B(a[47]), .Z(n8569) );
  NAND U8814 ( .A(n9364), .B(n8569), .Z(n8457) );
  NAND U8815 ( .A(n8458), .B(n8457), .Z(n8596) );
  XNOR U8816 ( .A(n8595), .B(n8596), .Z(n8598) );
  XNOR U8817 ( .A(n8597), .B(n8598), .Z(n8621) );
  NANDN U8818 ( .A(n554), .B(n8459), .Z(n8461) );
  XNOR U8819 ( .A(a[55]), .B(b[17]), .Z(n8588) );
  OR U8820 ( .A(n8588), .B(n9195), .Z(n8460) );
  AND U8821 ( .A(n8461), .B(n8460), .Z(n8567) );
  OR U8822 ( .A(n8462), .B(n574), .Z(n8464) );
  XNOR U8823 ( .A(b[19]), .B(a[53]), .Z(n8581) );
  OR U8824 ( .A(n8581), .B(n555), .Z(n8463) );
  AND U8825 ( .A(n8464), .B(n8463), .Z(n8565) );
  NAND U8826 ( .A(n572), .B(n8465), .Z(n8467) );
  XOR U8827 ( .A(a[59]), .B(b[13]), .Z(n8584) );
  NAND U8828 ( .A(n8585), .B(n8584), .Z(n8466) );
  NAND U8829 ( .A(n8467), .B(n8466), .Z(n8566) );
  XNOR U8830 ( .A(n8565), .B(n8566), .Z(n8568) );
  XNOR U8831 ( .A(n8567), .B(n8568), .Z(n8620) );
  NAND U8832 ( .A(n573), .B(n8468), .Z(n8470) );
  XOR U8833 ( .A(a[57]), .B(b[15]), .Z(n8578) );
  NAND U8834 ( .A(n8694), .B(n8578), .Z(n8469) );
  AND U8835 ( .A(n8470), .B(n8469), .Z(n8619) );
  XOR U8836 ( .A(n8620), .B(n8619), .Z(n8622) );
  XNOR U8837 ( .A(n8621), .B(n8622), .Z(n8548) );
  XNOR U8838 ( .A(n8549), .B(n8548), .Z(n8551) );
  XNOR U8839 ( .A(n8551), .B(n8550), .Z(n8630) );
  OR U8840 ( .A(n8475), .B(n559), .Z(n8477) );
  XNOR U8841 ( .A(b[29]), .B(a[43]), .Z(n8555) );
  OR U8842 ( .A(n8555), .B(n9796), .Z(n8476) );
  AND U8843 ( .A(n8477), .B(n8476), .Z(n8593) );
  OR U8844 ( .A(n8478), .B(n580), .Z(n8480) );
  XNOR U8845 ( .A(b[31]), .B(a[41]), .Z(n8599) );
  OR U8846 ( .A(n8599), .B(n9904), .Z(n8479) );
  AND U8847 ( .A(n8480), .B(n8479), .Z(n8591) );
  NAND U8848 ( .A(n578), .B(n8481), .Z(n8483) );
  XOR U8849 ( .A(b[23]), .B(a[49]), .Z(n8575) );
  NAND U8850 ( .A(n9268), .B(n8575), .Z(n8482) );
  NAND U8851 ( .A(n8483), .B(n8482), .Z(n8592) );
  XNOR U8852 ( .A(n8591), .B(n8592), .Z(n8594) );
  XNOR U8853 ( .A(n8593), .B(n8594), .Z(n8626) );
  OR U8854 ( .A(n8484), .B(n564), .Z(n8487) );
  XNOR U8855 ( .A(a[63]), .B(b[9]), .Z(n8602) );
  OR U8856 ( .A(n8602), .B(n8485), .Z(n8486) );
  AND U8857 ( .A(n8487), .B(n8486), .Z(n8561) );
  NAND U8858 ( .A(n577), .B(n8488), .Z(n8490) );
  XOR U8859 ( .A(b[21]), .B(a[51]), .Z(n8558) );
  NAND U8860 ( .A(n9216), .B(n8558), .Z(n8489) );
  NAND U8861 ( .A(n8490), .B(n8489), .Z(n8562) );
  XNOR U8862 ( .A(n8561), .B(n8562), .Z(n8564) );
  AND U8863 ( .A(b[31]), .B(a[39]), .Z(n8605) );
  IV U8864 ( .A(n8491), .Z(n8606) );
  XNOR U8865 ( .A(n8605), .B(n8606), .Z(n8608) );
  XNOR U8866 ( .A(n8492), .B(n8608), .Z(n8563) );
  XNOR U8867 ( .A(n8564), .B(n8563), .Z(n8625) );
  XNOR U8868 ( .A(n8626), .B(n8625), .Z(n8628) );
  IV U8869 ( .A(n8492), .Z(n8607) );
  NANDN U8870 ( .A(n8493), .B(n8607), .Z(n8497) );
  NANDN U8871 ( .A(n8495), .B(n8494), .Z(n8496) );
  NAND U8872 ( .A(n8497), .B(n8496), .Z(n8627) );
  XNOR U8873 ( .A(n8628), .B(n8627), .Z(n8617) );
  XOR U8874 ( .A(n8615), .B(n8616), .Z(n8618) );
  XOR U8875 ( .A(n8617), .B(n8618), .Z(n8629) );
  XOR U8876 ( .A(n8630), .B(n8629), .Z(n8632) );
  XNOR U8877 ( .A(n8631), .B(n8632), .Z(n8637) );
  NANDN U8878 ( .A(n8515), .B(n8514), .Z(n8519) );
  NANDN U8879 ( .A(n8517), .B(n8516), .Z(n8518) );
  AND U8880 ( .A(n8519), .B(n8518), .Z(n8611) );
  NANDN U8881 ( .A(n8521), .B(n8520), .Z(n8525) );
  NANDN U8882 ( .A(n8523), .B(n8522), .Z(n8524) );
  NAND U8883 ( .A(n8525), .B(n8524), .Z(n8612) );
  XNOR U8884 ( .A(n8611), .B(n8612), .Z(n8613) );
  XNOR U8885 ( .A(n8614), .B(n8613), .Z(n8635) );
  XNOR U8886 ( .A(n8636), .B(n8635), .Z(n8638) );
  XNOR U8887 ( .A(n8637), .B(n8638), .Z(n8640) );
  NANDN U8888 ( .A(n8527), .B(n8526), .Z(n8531) );
  NANDN U8889 ( .A(n8529), .B(n8528), .Z(n8530) );
  NAND U8890 ( .A(n8531), .B(n8530), .Z(n8639) );
  XNOR U8891 ( .A(n8640), .B(n8639), .Z(n8642) );
  XNOR U8892 ( .A(n8642), .B(n8641), .Z(n8543) );
  XOR U8893 ( .A(n8543), .B(n8542), .Z(n8545) );
  XOR U8894 ( .A(n8544), .B(n8545), .Z(n8540) );
  XOR U8895 ( .A(n8541), .B(n8540), .Z(c[103]) );
  AND U8896 ( .A(n8541), .B(n8540), .Z(n8644) );
  NANDN U8897 ( .A(n8543), .B(n8542), .Z(n8547) );
  NANDN U8898 ( .A(n8545), .B(n8544), .Z(n8546) );
  NAND U8899 ( .A(n8547), .B(n8546), .Z(n8647) );
  OR U8900 ( .A(n8552), .B(n562), .Z(n8554) );
  XNOR U8901 ( .A(a[62]), .B(b[11]), .Z(n8700) );
  OR U8902 ( .A(n8700), .B(n8701), .Z(n8553) );
  AND U8903 ( .A(n8554), .B(n8553), .Z(n8729) );
  OR U8904 ( .A(n8555), .B(n559), .Z(n8557) );
  XNOR U8905 ( .A(b[29]), .B(a[44]), .Z(n8687) );
  OR U8906 ( .A(n8687), .B(n9796), .Z(n8556) );
  AND U8907 ( .A(n8557), .B(n8556), .Z(n8727) );
  NAND U8908 ( .A(n577), .B(n8558), .Z(n8560) );
  XOR U8909 ( .A(b[21]), .B(a[52]), .Z(n8723) );
  NAND U8910 ( .A(n9216), .B(n8723), .Z(n8559) );
  NAND U8911 ( .A(n8560), .B(n8559), .Z(n8728) );
  XNOR U8912 ( .A(n8727), .B(n8728), .Z(n8730) );
  XNOR U8913 ( .A(n8729), .B(n8730), .Z(n8668) );
  XNOR U8914 ( .A(n8668), .B(n8667), .Z(n8670) );
  XNOR U8915 ( .A(n8670), .B(n8669), .Z(n8659) );
  NANDN U8916 ( .A(n566), .B(n8569), .Z(n8571) );
  XNOR U8917 ( .A(b[25]), .B(a[48]), .Z(n8711) );
  OR U8918 ( .A(n8711), .B(n9684), .Z(n8570) );
  AND U8919 ( .A(n8571), .B(n8570), .Z(n8736) );
  OR U8920 ( .A(n8572), .B(n565), .Z(n8574) );
  XNOR U8921 ( .A(b[27]), .B(a[46]), .Z(n8714) );
  OR U8922 ( .A(n8714), .B(n9692), .Z(n8573) );
  AND U8923 ( .A(n8574), .B(n8573), .Z(n8734) );
  NAND U8924 ( .A(n578), .B(n8575), .Z(n8577) );
  XOR U8925 ( .A(b[23]), .B(a[50]), .Z(n8704) );
  NAND U8926 ( .A(n9268), .B(n8704), .Z(n8576) );
  NAND U8927 ( .A(n8577), .B(n8576), .Z(n8735) );
  XNOR U8928 ( .A(n8734), .B(n8735), .Z(n8737) );
  XNOR U8929 ( .A(n8736), .B(n8737), .Z(n8674) );
  NANDN U8930 ( .A(n557), .B(n8578), .Z(n8580) );
  XOR U8931 ( .A(a[58]), .B(b[15]), .Z(n8693) );
  NANDN U8932 ( .A(n9067), .B(n8693), .Z(n8579) );
  AND U8933 ( .A(n8580), .B(n8579), .Z(n8709) );
  OR U8934 ( .A(n8581), .B(n574), .Z(n8583) );
  XOR U8935 ( .A(a[54]), .B(b[19]), .Z(n8717) );
  NANDN U8936 ( .A(n555), .B(n8717), .Z(n8582) );
  AND U8937 ( .A(n8583), .B(n8582), .Z(n8707) );
  NAND U8938 ( .A(n572), .B(n8584), .Z(n8587) );
  XOR U8939 ( .A(a[60]), .B(b[13]), .Z(n8697) );
  NAND U8940 ( .A(n8585), .B(n8697), .Z(n8586) );
  NAND U8941 ( .A(n8587), .B(n8586), .Z(n8708) );
  XNOR U8942 ( .A(n8707), .B(n8708), .Z(n8710) );
  XNOR U8943 ( .A(n8709), .B(n8710), .Z(n8672) );
  OR U8944 ( .A(n8588), .B(n554), .Z(n8590) );
  XNOR U8945 ( .A(a[56]), .B(b[17]), .Z(n8690) );
  OR U8946 ( .A(n8690), .B(n9195), .Z(n8589) );
  AND U8947 ( .A(n8590), .B(n8589), .Z(n8671) );
  XNOR U8948 ( .A(n8672), .B(n8671), .Z(n8673) );
  XOR U8949 ( .A(n8674), .B(n8673), .Z(n8665) );
  OR U8950 ( .A(n8599), .B(n580), .Z(n8601) );
  XNOR U8951 ( .A(b[31]), .B(a[42]), .Z(n8720) );
  OR U8952 ( .A(n8720), .B(n9904), .Z(n8600) );
  AND U8953 ( .A(n8601), .B(n8600), .Z(n8732) );
  OR U8954 ( .A(n8602), .B(n564), .Z(n8603) );
  AND U8955 ( .A(n8604), .B(n8603), .Z(n8731) );
  NAND U8956 ( .A(b[31]), .B(a[40]), .Z(n8811) );
  XNOR U8957 ( .A(n8731), .B(n8811), .Z(n8733) );
  XNOR U8958 ( .A(n8732), .B(n8733), .Z(n8682) );
  NAND U8959 ( .A(n8606), .B(n8605), .Z(n8610) );
  OR U8960 ( .A(n8608), .B(n8607), .Z(n8609) );
  AND U8961 ( .A(n8610), .B(n8609), .Z(n8681) );
  XOR U8962 ( .A(n8682), .B(n8681), .Z(n8684) );
  XOR U8963 ( .A(n8683), .B(n8684), .Z(n8664) );
  XOR U8964 ( .A(n8663), .B(n8664), .Z(n8666) );
  XOR U8965 ( .A(n8665), .B(n8666), .Z(n8660) );
  XNOR U8966 ( .A(n8659), .B(n8660), .Z(n8661) );
  XNOR U8967 ( .A(n8662), .B(n8661), .Z(n8658) );
  NANDN U8968 ( .A(n8620), .B(n8619), .Z(n8624) );
  OR U8969 ( .A(n8622), .B(n8621), .Z(n8623) );
  AND U8970 ( .A(n8624), .B(n8623), .Z(n8677) );
  XOR U8971 ( .A(n8677), .B(n8678), .Z(n8680) );
  XNOR U8972 ( .A(n8679), .B(n8680), .Z(n8656) );
  XNOR U8973 ( .A(n8655), .B(n8656), .Z(n8657) );
  XNOR U8974 ( .A(n8658), .B(n8657), .Z(n8651) );
  NANDN U8975 ( .A(n8630), .B(n8629), .Z(n8634) );
  NANDN U8976 ( .A(n8632), .B(n8631), .Z(n8633) );
  NAND U8977 ( .A(n8634), .B(n8633), .Z(n8652) );
  XNOR U8978 ( .A(n8651), .B(n8652), .Z(n8654) );
  XNOR U8979 ( .A(n8654), .B(n8653), .Z(n8646) );
  XOR U8980 ( .A(n8646), .B(n8645), .Z(n8648) );
  XOR U8981 ( .A(n8647), .B(n8648), .Z(n8643) );
  XOR U8982 ( .A(n8644), .B(n8643), .Z(c[104]) );
  AND U8983 ( .A(n8644), .B(n8643), .Z(n8739) );
  NANDN U8984 ( .A(n8646), .B(n8645), .Z(n8650) );
  NANDN U8985 ( .A(n8648), .B(n8647), .Z(n8649) );
  NAND U8986 ( .A(n8650), .B(n8649), .Z(n8742) );
  NANDN U8987 ( .A(n8672), .B(n8671), .Z(n8676) );
  NANDN U8988 ( .A(n8674), .B(n8673), .Z(n8675) );
  NAND U8989 ( .A(n8676), .B(n8675), .Z(n8823) );
  XOR U8990 ( .A(n8822), .B(n8823), .Z(n8825) );
  XNOR U8991 ( .A(n8824), .B(n8825), .Z(n8829) );
  NANDN U8992 ( .A(n8682), .B(n8681), .Z(n8686) );
  NANDN U8993 ( .A(n8684), .B(n8683), .Z(n8685) );
  AND U8994 ( .A(n8686), .B(n8685), .Z(n8752) );
  OR U8995 ( .A(n8687), .B(n559), .Z(n8689) );
  XNOR U8996 ( .A(b[29]), .B(a[45]), .Z(n8762) );
  OR U8997 ( .A(n8762), .B(n9796), .Z(n8688) );
  AND U8998 ( .A(n8689), .B(n8688), .Z(n8809) );
  OR U8999 ( .A(n8690), .B(n554), .Z(n8692) );
  XNOR U9000 ( .A(a[57]), .B(b[17]), .Z(n8765) );
  OR U9001 ( .A(n8765), .B(n9195), .Z(n8691) );
  AND U9002 ( .A(n8692), .B(n8691), .Z(n8807) );
  NAND U9003 ( .A(n573), .B(n8693), .Z(n8696) );
  XOR U9004 ( .A(a[59]), .B(b[15]), .Z(n8774) );
  NAND U9005 ( .A(n8694), .B(n8774), .Z(n8695) );
  NAND U9006 ( .A(n8696), .B(n8695), .Z(n8808) );
  XNOR U9007 ( .A(n8807), .B(n8808), .Z(n8810) );
  XNOR U9008 ( .A(n8809), .B(n8810), .Z(n8804) );
  NANDN U9009 ( .A(n553), .B(n8697), .Z(n8699) );
  XNOR U9010 ( .A(a[61]), .B(b[13]), .Z(n8777) );
  OR U9011 ( .A(n8777), .B(n8853), .Z(n8698) );
  NAND U9012 ( .A(n8699), .B(n8698), .Z(n8818) );
  OR U9013 ( .A(n8700), .B(n562), .Z(n8703) );
  XNOR U9014 ( .A(a[63]), .B(b[11]), .Z(n8796) );
  OR U9015 ( .A(n8796), .B(n8701), .Z(n8702) );
  AND U9016 ( .A(n8703), .B(n8702), .Z(n8815) );
  NANDN U9017 ( .A(n563), .B(n8704), .Z(n8706) );
  XNOR U9018 ( .A(b[23]), .B(a[51]), .Z(n8771) );
  OR U9019 ( .A(n8771), .B(n9605), .Z(n8705) );
  NAND U9020 ( .A(n8706), .B(n8705), .Z(n8816) );
  XOR U9021 ( .A(n8815), .B(n8816), .Z(n8819) );
  XOR U9022 ( .A(n8818), .B(n8819), .Z(n8803) );
  XNOR U9023 ( .A(n8804), .B(n8803), .Z(n8806) );
  XNOR U9024 ( .A(n8806), .B(n8805), .Z(n8751) );
  OR U9025 ( .A(n8711), .B(n566), .Z(n8713) );
  XNOR U9026 ( .A(b[25]), .B(a[49]), .Z(n8784) );
  OR U9027 ( .A(n8784), .B(n9684), .Z(n8712) );
  AND U9028 ( .A(n8713), .B(n8712), .Z(n8782) );
  OR U9029 ( .A(n8714), .B(n565), .Z(n8716) );
  XOR U9030 ( .A(b[27]), .B(a[47]), .Z(n8768) );
  NANDN U9031 ( .A(n9692), .B(n8768), .Z(n8715) );
  AND U9032 ( .A(n8716), .B(n8715), .Z(n8780) );
  NAND U9033 ( .A(n9046), .B(n8717), .Z(n8719) );
  XOR U9034 ( .A(a[55]), .B(b[19]), .Z(n8790) );
  NAND U9035 ( .A(n575), .B(n8790), .Z(n8718) );
  NAND U9036 ( .A(n8719), .B(n8718), .Z(n8781) );
  XNOR U9037 ( .A(n8780), .B(n8781), .Z(n8783) );
  XNOR U9038 ( .A(n8782), .B(n8783), .Z(n8759) );
  OR U9039 ( .A(n8720), .B(n580), .Z(n8722) );
  XNOR U9040 ( .A(b[31]), .B(a[43]), .Z(n8793) );
  OR U9041 ( .A(n8793), .B(n9904), .Z(n8721) );
  AND U9042 ( .A(n8722), .B(n8721), .Z(n8799) );
  NAND U9043 ( .A(n577), .B(n8723), .Z(n8725) );
  XOR U9044 ( .A(b[21]), .B(a[53]), .Z(n8787) );
  NAND U9045 ( .A(n9216), .B(n8787), .Z(n8724) );
  NAND U9046 ( .A(n8725), .B(n8724), .Z(n8800) );
  XNOR U9047 ( .A(n8799), .B(n8800), .Z(n8802) );
  IV U9048 ( .A(n8726), .Z(n8812) );
  XNOR U9049 ( .A(n8812), .B(n8811), .Z(n8814) );
  AND U9050 ( .A(b[31]), .B(a[41]), .Z(n8813) );
  XOR U9051 ( .A(n8814), .B(n8813), .Z(n8801) );
  XNOR U9052 ( .A(n8802), .B(n8801), .Z(n8758) );
  XNOR U9053 ( .A(n8759), .B(n8758), .Z(n8761) );
  XNOR U9054 ( .A(n8761), .B(n8760), .Z(n8757) );
  XNOR U9055 ( .A(n8755), .B(n8754), .Z(n8756) );
  XNOR U9056 ( .A(n8757), .B(n8756), .Z(n8750) );
  XNOR U9057 ( .A(n8751), .B(n8750), .Z(n8753) );
  XNOR U9058 ( .A(n8752), .B(n8753), .Z(n8827) );
  XNOR U9059 ( .A(n8826), .B(n8827), .Z(n8828) );
  XNOR U9060 ( .A(n8829), .B(n8828), .Z(n8746) );
  XNOR U9061 ( .A(n8747), .B(n8746), .Z(n8749) );
  XNOR U9062 ( .A(n8748), .B(n8749), .Z(n8740) );
  XNOR U9063 ( .A(n8741), .B(n8740), .Z(n8743) );
  XOR U9064 ( .A(n8742), .B(n8743), .Z(n8738) );
  XOR U9065 ( .A(n8739), .B(n8738), .Z(c[105]) );
  AND U9066 ( .A(n8739), .B(n8738), .Z(n8831) );
  NAND U9067 ( .A(n8741), .B(n8740), .Z(n8745) );
  NANDN U9068 ( .A(n8743), .B(n8742), .Z(n8744) );
  NAND U9069 ( .A(n8745), .B(n8744), .Z(n8834) );
  OR U9070 ( .A(n8762), .B(n559), .Z(n8764) );
  XNOR U9071 ( .A(b[29]), .B(a[46]), .Z(n8849) );
  OR U9072 ( .A(n8849), .B(n9796), .Z(n8763) );
  AND U9073 ( .A(n8764), .B(n8763), .Z(n8844) );
  OR U9074 ( .A(n8765), .B(n554), .Z(n8767) );
  XNOR U9075 ( .A(a[58]), .B(b[17]), .Z(n8870) );
  OR U9076 ( .A(n8870), .B(n9195), .Z(n8766) );
  AND U9077 ( .A(n8767), .B(n8766), .Z(n8842) );
  NAND U9078 ( .A(n582), .B(n8768), .Z(n8770) );
  XOR U9079 ( .A(b[27]), .B(a[48]), .Z(n8879) );
  NAND U9080 ( .A(n9770), .B(n8879), .Z(n8769) );
  NAND U9081 ( .A(n8770), .B(n8769), .Z(n8843) );
  XNOR U9082 ( .A(n8842), .B(n8843), .Z(n8845) );
  XNOR U9083 ( .A(n8844), .B(n8845), .Z(n8894) );
  OR U9084 ( .A(n8771), .B(n563), .Z(n8773) );
  XOR U9085 ( .A(b[23]), .B(a[52]), .Z(n8862) );
  NANDN U9086 ( .A(n9605), .B(n8862), .Z(n8772) );
  NAND U9087 ( .A(n8773), .B(n8772), .Z(n8868) );
  NANDN U9088 ( .A(n557), .B(n8774), .Z(n8776) );
  XNOR U9089 ( .A(a[60]), .B(b[15]), .Z(n8873) );
  OR U9090 ( .A(n8873), .B(n9067), .Z(n8775) );
  AND U9091 ( .A(n8776), .B(n8775), .Z(n8866) );
  OR U9092 ( .A(n8777), .B(n553), .Z(n8779) );
  XNOR U9093 ( .A(a[62]), .B(b[13]), .Z(n8852) );
  OR U9094 ( .A(n8852), .B(n8853), .Z(n8778) );
  NAND U9095 ( .A(n8779), .B(n8778), .Z(n8867) );
  XOR U9096 ( .A(n8866), .B(n8867), .Z(n8869) );
  XOR U9097 ( .A(n8868), .B(n8869), .Z(n8893) );
  XNOR U9098 ( .A(n8894), .B(n8893), .Z(n8896) );
  XNOR U9099 ( .A(n8896), .B(n8895), .Z(n8901) );
  OR U9100 ( .A(n8784), .B(n566), .Z(n8786) );
  XNOR U9101 ( .A(b[25]), .B(a[50]), .Z(n8876) );
  OR U9102 ( .A(n8876), .B(n9684), .Z(n8785) );
  AND U9103 ( .A(n8786), .B(n8785), .Z(n8887) );
  NANDN U9104 ( .A(n556), .B(n8787), .Z(n8789) );
  XOR U9105 ( .A(b[21]), .B(a[54]), .Z(n8856) );
  NANDN U9106 ( .A(n9480), .B(n8856), .Z(n8788) );
  AND U9107 ( .A(n8789), .B(n8788), .Z(n8885) );
  NAND U9108 ( .A(n9046), .B(n8790), .Z(n8792) );
  XOR U9109 ( .A(a[56]), .B(b[19]), .Z(n8882) );
  NAND U9110 ( .A(n575), .B(n8882), .Z(n8791) );
  NAND U9111 ( .A(n8792), .B(n8791), .Z(n8886) );
  XNOR U9112 ( .A(n8885), .B(n8886), .Z(n8888) );
  XNOR U9113 ( .A(n8887), .B(n8888), .Z(n8890) );
  OR U9114 ( .A(n8793), .B(n580), .Z(n8795) );
  XNOR U9115 ( .A(b[31]), .B(a[44]), .Z(n8859) );
  OR U9116 ( .A(n8859), .B(n9904), .Z(n8794) );
  NAND U9117 ( .A(n8795), .B(n8794), .Z(n8847) );
  AND U9118 ( .A(b[31]), .B(a[42]), .Z(n8943) );
  OR U9119 ( .A(n8796), .B(n562), .Z(n8797) );
  AND U9120 ( .A(n8798), .B(n8797), .Z(n8846) );
  XNOR U9121 ( .A(n8943), .B(n8846), .Z(n8848) );
  XOR U9122 ( .A(n8847), .B(n8848), .Z(n8889) );
  XNOR U9123 ( .A(n8890), .B(n8889), .Z(n8892) );
  XNOR U9124 ( .A(n8892), .B(n8891), .Z(n8900) );
  XNOR U9125 ( .A(n8901), .B(n8900), .Z(n8902) );
  XNOR U9126 ( .A(n8903), .B(n8902), .Z(n8841) );
  IV U9127 ( .A(n8815), .Z(n8817) );
  NAND U9128 ( .A(n8817), .B(n8816), .Z(n8821) );
  NANDN U9129 ( .A(n8819), .B(n8818), .Z(n8820) );
  AND U9130 ( .A(n8821), .B(n8820), .Z(n8904) );
  XNOR U9131 ( .A(n8905), .B(n8904), .Z(n8906) );
  XNOR U9132 ( .A(n8907), .B(n8906), .Z(n8839) );
  XNOR U9133 ( .A(n8838), .B(n8839), .Z(n8840) );
  XNOR U9134 ( .A(n8841), .B(n8840), .Z(n8909) );
  XNOR U9135 ( .A(n8908), .B(n8909), .Z(n8911) );
  XNOR U9136 ( .A(n8910), .B(n8911), .Z(n8913) );
  XNOR U9137 ( .A(n8913), .B(n8912), .Z(n8915) );
  XNOR U9138 ( .A(n8915), .B(n8914), .Z(n8833) );
  XOR U9139 ( .A(n8832), .B(n8833), .Z(n8835) );
  XOR U9140 ( .A(n8834), .B(n8835), .Z(n8830) );
  XOR U9141 ( .A(n8831), .B(n8830), .Z(c[106]) );
  AND U9142 ( .A(n8831), .B(n8830), .Z(n8917) );
  NANDN U9143 ( .A(n8833), .B(n8832), .Z(n8837) );
  NANDN U9144 ( .A(n8835), .B(n8834), .Z(n8836) );
  NAND U9145 ( .A(n8837), .B(n8836), .Z(n8920) );
  OR U9146 ( .A(n8849), .B(n559), .Z(n8851) );
  XNOR U9147 ( .A(b[29]), .B(a[47]), .Z(n8964) );
  OR U9148 ( .A(n8964), .B(n9796), .Z(n8850) );
  AND U9149 ( .A(n8851), .B(n8850), .Z(n8972) );
  OR U9150 ( .A(n8852), .B(n553), .Z(n8855) );
  XNOR U9151 ( .A(a[63]), .B(b[13]), .Z(n8980) );
  OR U9152 ( .A(n8980), .B(n8853), .Z(n8854) );
  AND U9153 ( .A(n8855), .B(n8854), .Z(n8970) );
  NAND U9154 ( .A(n577), .B(n8856), .Z(n8858) );
  XOR U9155 ( .A(a[55]), .B(b[21]), .Z(n8958) );
  NAND U9156 ( .A(n9216), .B(n8958), .Z(n8857) );
  NAND U9157 ( .A(n8858), .B(n8857), .Z(n8971) );
  XNOR U9158 ( .A(n8970), .B(n8971), .Z(n8973) );
  XNOR U9159 ( .A(n8972), .B(n8973), .Z(n8975) );
  OR U9160 ( .A(n8859), .B(n580), .Z(n8861) );
  XOR U9161 ( .A(b[31]), .B(a[45]), .Z(n8983) );
  NANDN U9162 ( .A(n9904), .B(n8983), .Z(n8860) );
  AND U9163 ( .A(n8861), .B(n8860), .Z(n8992) );
  NAND U9164 ( .A(n578), .B(n8862), .Z(n8864) );
  XOR U9165 ( .A(b[23]), .B(a[53]), .Z(n8967) );
  NAND U9166 ( .A(n9268), .B(n8967), .Z(n8863) );
  NAND U9167 ( .A(n8864), .B(n8863), .Z(n8993) );
  XNOR U9168 ( .A(n8992), .B(n8993), .Z(n8994) );
  AND U9169 ( .A(b[31]), .B(a[43]), .Z(n8940) );
  XNOR U9170 ( .A(n8940), .B(n8865), .Z(n8942) );
  XNOR U9171 ( .A(n8943), .B(n8942), .Z(n8995) );
  XOR U9172 ( .A(n8994), .B(n8995), .Z(n8974) );
  XOR U9173 ( .A(n8975), .B(n8974), .Z(n8977) );
  XNOR U9174 ( .A(n8976), .B(n8977), .Z(n9004) );
  OR U9175 ( .A(n8870), .B(n554), .Z(n8872) );
  XNOR U9176 ( .A(a[59]), .B(b[17]), .Z(n8946) );
  OR U9177 ( .A(n8946), .B(n9195), .Z(n8871) );
  AND U9178 ( .A(n8872), .B(n8871), .Z(n8938) );
  OR U9179 ( .A(n8873), .B(n557), .Z(n8875) );
  XNOR U9180 ( .A(a[61]), .B(b[15]), .Z(n8949) );
  OR U9181 ( .A(n8949), .B(n9067), .Z(n8874) );
  AND U9182 ( .A(n8875), .B(n8874), .Z(n8936) );
  OR U9183 ( .A(n8876), .B(n566), .Z(n8878) );
  XOR U9184 ( .A(b[25]), .B(a[51]), .Z(n8952) );
  NANDN U9185 ( .A(n9684), .B(n8952), .Z(n8877) );
  NAND U9186 ( .A(n8878), .B(n8877), .Z(n8988) );
  NANDN U9187 ( .A(n565), .B(n8879), .Z(n8881) );
  XNOR U9188 ( .A(b[27]), .B(a[49]), .Z(n8961) );
  OR U9189 ( .A(n8961), .B(n9692), .Z(n8880) );
  NAND U9190 ( .A(n8881), .B(n8880), .Z(n8987) );
  NAND U9191 ( .A(n9046), .B(n8882), .Z(n8884) );
  XOR U9192 ( .A(a[57]), .B(b[19]), .Z(n8955) );
  NAND U9193 ( .A(n575), .B(n8955), .Z(n8883) );
  NAND U9194 ( .A(n8884), .B(n8883), .Z(n8986) );
  XOR U9195 ( .A(n8987), .B(n8986), .Z(n8989) );
  XOR U9196 ( .A(n8988), .B(n8989), .Z(n8937) );
  XNOR U9197 ( .A(n8936), .B(n8937), .Z(n8939) );
  XNOR U9198 ( .A(n8938), .B(n8939), .Z(n9003) );
  XNOR U9199 ( .A(n9002), .B(n9003), .Z(n9005) );
  XNOR U9200 ( .A(n9004), .B(n9005), .Z(n8997) );
  XOR U9201 ( .A(n8997), .B(n8996), .Z(n8999) );
  XNOR U9202 ( .A(n8998), .B(n8999), .Z(n8934) );
  NANDN U9203 ( .A(n8894), .B(n8893), .Z(n8899) );
  IV U9204 ( .A(n8895), .Z(n8897) );
  NAND U9205 ( .A(n8897), .B(n8896), .Z(n8898) );
  NAND U9206 ( .A(n8899), .B(n8898), .Z(n8932) );
  XNOR U9207 ( .A(n8933), .B(n8932), .Z(n8935) );
  XNOR U9208 ( .A(n8934), .B(n8935), .Z(n8931) );
  XNOR U9209 ( .A(n8928), .B(n8929), .Z(n8930) );
  XNOR U9210 ( .A(n8931), .B(n8930), .Z(n8924) );
  XNOR U9211 ( .A(n8925), .B(n8924), .Z(n8927) );
  XNOR U9212 ( .A(n8927), .B(n8926), .Z(n8919) );
  XOR U9213 ( .A(n8919), .B(n8918), .Z(n8921) );
  XOR U9214 ( .A(n8920), .B(n8921), .Z(n8916) );
  XOR U9215 ( .A(n8917), .B(n8916), .Z(c[107]) );
  AND U9216 ( .A(n8917), .B(n8916), .Z(n9007) );
  NANDN U9217 ( .A(n8919), .B(n8918), .Z(n8923) );
  NANDN U9218 ( .A(n8921), .B(n8920), .Z(n8922) );
  NAND U9219 ( .A(n8923), .B(n8922), .Z(n9010) );
  NAND U9220 ( .A(n8941), .B(n8940), .Z(n8945) );
  NAND U9221 ( .A(n8943), .B(n8942), .Z(n8944) );
  AND U9222 ( .A(n8945), .B(n8944), .Z(n9062) );
  OR U9223 ( .A(n8946), .B(n554), .Z(n8948) );
  XNOR U9224 ( .A(a[60]), .B(b[17]), .Z(n9030) );
  OR U9225 ( .A(n9030), .B(n9195), .Z(n8947) );
  AND U9226 ( .A(n8948), .B(n8947), .Z(n9054) );
  OR U9227 ( .A(n8949), .B(n557), .Z(n8951) );
  XNOR U9228 ( .A(a[62]), .B(b[15]), .Z(n9066) );
  OR U9229 ( .A(n9066), .B(n9067), .Z(n8950) );
  AND U9230 ( .A(n8951), .B(n8950), .Z(n9052) );
  NAND U9231 ( .A(n579), .B(n8952), .Z(n8954) );
  XOR U9232 ( .A(b[25]), .B(a[52]), .Z(n9070) );
  NAND U9233 ( .A(n9364), .B(n9070), .Z(n8953) );
  NAND U9234 ( .A(n8954), .B(n8953), .Z(n9053) );
  XNOR U9235 ( .A(n9052), .B(n9053), .Z(n9055) );
  XNOR U9236 ( .A(n9054), .B(n9055), .Z(n9063) );
  XNOR U9237 ( .A(n9062), .B(n9063), .Z(n9064) );
  NANDN U9238 ( .A(n574), .B(n8955), .Z(n8957) );
  XOR U9239 ( .A(a[58]), .B(b[19]), .Z(n9045) );
  NANDN U9240 ( .A(n555), .B(n9045), .Z(n8956) );
  NAND U9241 ( .A(n8957), .B(n8956), .Z(n9058) );
  NANDN U9242 ( .A(n556), .B(n8958), .Z(n8960) );
  XNOR U9243 ( .A(a[56]), .B(b[21]), .Z(n9049) );
  OR U9244 ( .A(n9049), .B(n9480), .Z(n8959) );
  NAND U9245 ( .A(n8960), .B(n8959), .Z(n9056) );
  OR U9246 ( .A(n8961), .B(n565), .Z(n8963) );
  XNOR U9247 ( .A(b[27]), .B(a[50]), .Z(n9039) );
  OR U9248 ( .A(n9039), .B(n9692), .Z(n8962) );
  NAND U9249 ( .A(n8963), .B(n8962), .Z(n9076) );
  OR U9250 ( .A(n8964), .B(n559), .Z(n8966) );
  XNOR U9251 ( .A(b[29]), .B(a[48]), .Z(n9042) );
  OR U9252 ( .A(n9042), .B(n9796), .Z(n8965) );
  AND U9253 ( .A(n8966), .B(n8965), .Z(n9074) );
  NANDN U9254 ( .A(n563), .B(n8967), .Z(n8969) );
  XOR U9255 ( .A(b[23]), .B(a[54]), .Z(n9036) );
  NANDN U9256 ( .A(n9605), .B(n9036), .Z(n8968) );
  NAND U9257 ( .A(n8969), .B(n8968), .Z(n9075) );
  XOR U9258 ( .A(n9074), .B(n9075), .Z(n9077) );
  XOR U9259 ( .A(n9076), .B(n9077), .Z(n9057) );
  XOR U9260 ( .A(n9056), .B(n9057), .Z(n9059) );
  XOR U9261 ( .A(n9058), .B(n9059), .Z(n9065) );
  XOR U9262 ( .A(n9064), .B(n9065), .Z(n9023) );
  XOR U9263 ( .A(n9023), .B(n9022), .Z(n9025) );
  XNOR U9264 ( .A(n9024), .B(n9025), .Z(n9083) );
  NANDN U9265 ( .A(n8975), .B(n8974), .Z(n8979) );
  NANDN U9266 ( .A(n8977), .B(n8976), .Z(n8978) );
  NAND U9267 ( .A(n8979), .B(n8978), .Z(n9082) );
  OR U9268 ( .A(n8980), .B(n553), .Z(n8981) );
  AND U9269 ( .A(n8982), .B(n8981), .Z(n9080) );
  AND U9270 ( .A(b[31]), .B(a[44]), .Z(n9116) );
  NAND U9271 ( .A(n9764), .B(n8983), .Z(n8985) );
  XOR U9272 ( .A(b[31]), .B(a[46]), .Z(n9033) );
  NAND U9273 ( .A(n584), .B(n9033), .Z(n8984) );
  NAND U9274 ( .A(n8985), .B(n8984), .Z(n9078) );
  XNOR U9275 ( .A(n9116), .B(n9078), .Z(n9079) );
  XNOR U9276 ( .A(n9080), .B(n9079), .Z(n9026) );
  NAND U9277 ( .A(n8987), .B(n8986), .Z(n8991) );
  NAND U9278 ( .A(n8989), .B(n8988), .Z(n8990) );
  AND U9279 ( .A(n8991), .B(n8990), .Z(n9027) );
  XNOR U9280 ( .A(n9026), .B(n9027), .Z(n9029) );
  XNOR U9281 ( .A(n9029), .B(n9028), .Z(n9081) );
  XOR U9282 ( .A(n9082), .B(n9081), .Z(n9084) );
  XNOR U9283 ( .A(n9083), .B(n9084), .Z(n9020) );
  NANDN U9284 ( .A(n8997), .B(n8996), .Z(n9001) );
  NANDN U9285 ( .A(n8999), .B(n8998), .Z(n9000) );
  NAND U9286 ( .A(n9001), .B(n9000), .Z(n9019) );
  XOR U9287 ( .A(n9019), .B(n9018), .Z(n9021) );
  XNOR U9288 ( .A(n9020), .B(n9021), .Z(n9014) );
  XNOR U9289 ( .A(n9015), .B(n9014), .Z(n9016) );
  XNOR U9290 ( .A(n9017), .B(n9016), .Z(n9008) );
  XNOR U9291 ( .A(n9009), .B(n9008), .Z(n9011) );
  XOR U9292 ( .A(n9010), .B(n9011), .Z(n9006) );
  XOR U9293 ( .A(n9007), .B(n9006), .Z(c[108]) );
  AND U9294 ( .A(n9007), .B(n9006), .Z(n9086) );
  NAND U9295 ( .A(n9009), .B(n9008), .Z(n9013) );
  NANDN U9296 ( .A(n9011), .B(n9010), .Z(n9012) );
  NAND U9297 ( .A(n9013), .B(n9012), .Z(n9089) );
  XNOR U9298 ( .A(n9100), .B(n9099), .Z(n9102) );
  OR U9299 ( .A(n9030), .B(n554), .Z(n9032) );
  XOR U9300 ( .A(a[61]), .B(b[17]), .Z(n9140) );
  NANDN U9301 ( .A(n9195), .B(n9140), .Z(n9031) );
  AND U9302 ( .A(n9032), .B(n9031), .Z(n9153) );
  NANDN U9303 ( .A(n580), .B(n9033), .Z(n9035) );
  XNOR U9304 ( .A(b[31]), .B(a[47]), .Z(n9122) );
  OR U9305 ( .A(n9122), .B(n9904), .Z(n9034) );
  AND U9306 ( .A(n9035), .B(n9034), .Z(n9151) );
  NAND U9307 ( .A(n578), .B(n9036), .Z(n9038) );
  XOR U9308 ( .A(b[23]), .B(a[55]), .Z(n9137) );
  NAND U9309 ( .A(n9268), .B(n9137), .Z(n9037) );
  NAND U9310 ( .A(n9038), .B(n9037), .Z(n9152) );
  XNOR U9311 ( .A(n9151), .B(n9152), .Z(n9154) );
  XNOR U9312 ( .A(n9153), .B(n9154), .Z(n9106) );
  OR U9313 ( .A(n9039), .B(n565), .Z(n9041) );
  XNOR U9314 ( .A(b[27]), .B(a[51]), .Z(n9125) );
  OR U9315 ( .A(n9125), .B(n9692), .Z(n9040) );
  AND U9316 ( .A(n9041), .B(n9040), .Z(n9149) );
  OR U9317 ( .A(n9042), .B(n559), .Z(n9044) );
  XNOR U9318 ( .A(b[29]), .B(a[49]), .Z(n9128) );
  OR U9319 ( .A(n9128), .B(n9796), .Z(n9043) );
  AND U9320 ( .A(n9044), .B(n9043), .Z(n9147) );
  NAND U9321 ( .A(n9046), .B(n9045), .Z(n9048) );
  XOR U9322 ( .A(a[59]), .B(b[19]), .Z(n9144) );
  NAND U9323 ( .A(n575), .B(n9144), .Z(n9047) );
  NAND U9324 ( .A(n9048), .B(n9047), .Z(n9148) );
  XNOR U9325 ( .A(n9147), .B(n9148), .Z(n9150) );
  XNOR U9326 ( .A(n9149), .B(n9150), .Z(n9104) );
  OR U9327 ( .A(n9049), .B(n556), .Z(n9051) );
  XNOR U9328 ( .A(a[57]), .B(b[21]), .Z(n9134) );
  OR U9329 ( .A(n9134), .B(n9480), .Z(n9050) );
  AND U9330 ( .A(n9051), .B(n9050), .Z(n9103) );
  XNOR U9331 ( .A(n9104), .B(n9103), .Z(n9105) );
  XNOR U9332 ( .A(n9106), .B(n9105), .Z(n9160) );
  XNOR U9333 ( .A(n9160), .B(n9159), .Z(n9162) );
  NANDN U9334 ( .A(n9057), .B(n9056), .Z(n9061) );
  NANDN U9335 ( .A(n9059), .B(n9058), .Z(n9060) );
  NAND U9336 ( .A(n9061), .B(n9060), .Z(n9161) );
  XNOR U9337 ( .A(n9162), .B(n9161), .Z(n9165) );
  OR U9338 ( .A(n9066), .B(n557), .Z(n9069) );
  XNOR U9339 ( .A(a[63]), .B(b[15]), .Z(n9119) );
  OR U9340 ( .A(n9119), .B(n9067), .Z(n9068) );
  AND U9341 ( .A(n9069), .B(n9068), .Z(n9109) );
  NAND U9342 ( .A(n579), .B(n9070), .Z(n9072) );
  XOR U9343 ( .A(b[25]), .B(a[53]), .Z(n9131) );
  NAND U9344 ( .A(n9364), .B(n9131), .Z(n9071) );
  NAND U9345 ( .A(n9072), .B(n9071), .Z(n9110) );
  XNOR U9346 ( .A(n9109), .B(n9110), .Z(n9111) );
  AND U9347 ( .A(b[31]), .B(a[45]), .Z(n9113) );
  XNOR U9348 ( .A(n9113), .B(n9073), .Z(n9115) );
  XNOR U9349 ( .A(n9116), .B(n9115), .Z(n9112) );
  XNOR U9350 ( .A(n9111), .B(n9112), .Z(n9155) );
  XNOR U9351 ( .A(n9155), .B(n9156), .Z(n9158) );
  XNOR U9352 ( .A(n9158), .B(n9157), .Z(n9164) );
  XOR U9353 ( .A(n9163), .B(n9164), .Z(n9166) );
  XNOR U9354 ( .A(n9165), .B(n9166), .Z(n9101) );
  XNOR U9355 ( .A(n9102), .B(n9101), .Z(n9094) );
  XOR U9356 ( .A(n9094), .B(n9093), .Z(n9096) );
  XOR U9357 ( .A(n9095), .B(n9096), .Z(n9088) );
  XOR U9358 ( .A(n9087), .B(n9088), .Z(n9090) );
  XOR U9359 ( .A(n9089), .B(n9090), .Z(n9085) );
  XOR U9360 ( .A(n9086), .B(n9085), .Z(c[109]) );
  AND U9361 ( .A(n9086), .B(n9085), .Z(n9170) );
  NANDN U9362 ( .A(n9088), .B(n9087), .Z(n9092) );
  NANDN U9363 ( .A(n9090), .B(n9089), .Z(n9091) );
  NAND U9364 ( .A(n9092), .B(n9091), .Z(n9173) );
  NANDN U9365 ( .A(n9094), .B(n9093), .Z(n9098) );
  NANDN U9366 ( .A(n9096), .B(n9095), .Z(n9097) );
  NAND U9367 ( .A(n9098), .B(n9097), .Z(n9171) );
  NANDN U9368 ( .A(n9104), .B(n9103), .Z(n9108) );
  NANDN U9369 ( .A(n9106), .B(n9105), .Z(n9107) );
  AND U9370 ( .A(n9108), .B(n9107), .Z(n9185) );
  NAND U9371 ( .A(n9114), .B(n9113), .Z(n9118) );
  NAND U9372 ( .A(n9116), .B(n9115), .Z(n9117) );
  NAND U9373 ( .A(n9118), .B(n9117), .Z(n9238) );
  OR U9374 ( .A(n9119), .B(n557), .Z(n9120) );
  AND U9375 ( .A(n9121), .B(n9120), .Z(n9228) );
  AND U9376 ( .A(b[31]), .B(a[46]), .Z(n9225) );
  OR U9377 ( .A(n9122), .B(n580), .Z(n9124) );
  XNOR U9378 ( .A(b[31]), .B(a[48]), .Z(n9219) );
  OR U9379 ( .A(n9219), .B(n9904), .Z(n9123) );
  NAND U9380 ( .A(n9124), .B(n9123), .Z(n9226) );
  XOR U9381 ( .A(n9225), .B(n9226), .Z(n9227) );
  XNOR U9382 ( .A(n9228), .B(n9227), .Z(n9237) );
  XOR U9383 ( .A(n9238), .B(n9237), .Z(n9240) );
  XOR U9384 ( .A(n9239), .B(n9240), .Z(n9186) );
  XNOR U9385 ( .A(n9185), .B(n9186), .Z(n9187) );
  OR U9386 ( .A(n9125), .B(n565), .Z(n9127) );
  XNOR U9387 ( .A(b[27]), .B(a[52]), .Z(n9209) );
  OR U9388 ( .A(n9209), .B(n9692), .Z(n9126) );
  AND U9389 ( .A(n9127), .B(n9126), .Z(n9203) );
  OR U9390 ( .A(n9128), .B(n559), .Z(n9130) );
  XNOR U9391 ( .A(b[29]), .B(a[50]), .Z(n9212) );
  OR U9392 ( .A(n9212), .B(n9796), .Z(n9129) );
  AND U9393 ( .A(n9130), .B(n9129), .Z(n9201) );
  NAND U9394 ( .A(n579), .B(n9131), .Z(n9133) );
  XOR U9395 ( .A(b[25]), .B(a[54]), .Z(n9222) );
  NAND U9396 ( .A(n9364), .B(n9222), .Z(n9132) );
  NAND U9397 ( .A(n9133), .B(n9132), .Z(n9202) );
  XNOR U9398 ( .A(n9201), .B(n9202), .Z(n9204) );
  XNOR U9399 ( .A(n9203), .B(n9204), .Z(n9234) );
  OR U9400 ( .A(n9134), .B(n556), .Z(n9136) );
  XOR U9401 ( .A(a[58]), .B(b[21]), .Z(n9215) );
  NANDN U9402 ( .A(n9480), .B(n9215), .Z(n9135) );
  AND U9403 ( .A(n9136), .B(n9135), .Z(n9207) );
  NANDN U9404 ( .A(n563), .B(n9137), .Z(n9139) );
  XOR U9405 ( .A(b[23]), .B(a[56]), .Z(n9198) );
  NANDN U9406 ( .A(n9605), .B(n9198), .Z(n9138) );
  AND U9407 ( .A(n9139), .B(n9138), .Z(n9205) );
  NAND U9408 ( .A(n576), .B(n9140), .Z(n9143) );
  XOR U9409 ( .A(a[62]), .B(b[17]), .Z(n9194) );
  NAND U9410 ( .A(n9141), .B(n9194), .Z(n9142) );
  NAND U9411 ( .A(n9143), .B(n9142), .Z(n9206) );
  XNOR U9412 ( .A(n9205), .B(n9206), .Z(n9208) );
  XNOR U9413 ( .A(n9207), .B(n9208), .Z(n9232) );
  NANDN U9414 ( .A(n574), .B(n9144), .Z(n9146) );
  XNOR U9415 ( .A(a[60]), .B(b[19]), .Z(n9191) );
  OR U9416 ( .A(n9191), .B(n555), .Z(n9145) );
  AND U9417 ( .A(n9146), .B(n9145), .Z(n9231) );
  XNOR U9418 ( .A(n9232), .B(n9231), .Z(n9233) );
  XOR U9419 ( .A(n9234), .B(n9233), .Z(n9243) );
  XOR U9420 ( .A(n9241), .B(n9242), .Z(n9244) );
  XOR U9421 ( .A(n9243), .B(n9244), .Z(n9188) );
  XNOR U9422 ( .A(n9187), .B(n9188), .Z(n9183) );
  XNOR U9423 ( .A(n9181), .B(n9182), .Z(n9184) );
  XNOR U9424 ( .A(n9183), .B(n9184), .Z(n9178) );
  NANDN U9425 ( .A(n9164), .B(n9163), .Z(n9168) );
  OR U9426 ( .A(n9166), .B(n9165), .Z(n9167) );
  NAND U9427 ( .A(n9168), .B(n9167), .Z(n9177) );
  XNOR U9428 ( .A(n9178), .B(n9177), .Z(n9180) );
  XNOR U9429 ( .A(n9179), .B(n9180), .Z(n9172) );
  XOR U9430 ( .A(n9171), .B(n9172), .Z(n9174) );
  XOR U9431 ( .A(n9173), .B(n9174), .Z(n9169) );
  XOR U9432 ( .A(n9170), .B(n9169), .Z(c[110]) );
  AND U9433 ( .A(n9170), .B(n9169), .Z(n9246) );
  NANDN U9434 ( .A(n9172), .B(n9171), .Z(n9176) );
  NANDN U9435 ( .A(n9174), .B(n9173), .Z(n9175) );
  NAND U9436 ( .A(n9176), .B(n9175), .Z(n9249) );
  NANDN U9437 ( .A(n9186), .B(n9185), .Z(n9190) );
  NANDN U9438 ( .A(n9188), .B(n9187), .Z(n9189) );
  AND U9439 ( .A(n9190), .B(n9189), .Z(n9253) );
  OR U9440 ( .A(n9191), .B(n574), .Z(n9193) );
  XNOR U9441 ( .A(a[61]), .B(b[19]), .Z(n9288) );
  OR U9442 ( .A(n9288), .B(n555), .Z(n9192) );
  AND U9443 ( .A(n9193), .B(n9192), .Z(n9302) );
  NANDN U9444 ( .A(n554), .B(n9194), .Z(n9197) );
  XNOR U9445 ( .A(a[63]), .B(b[17]), .Z(n9297) );
  OR U9446 ( .A(n9297), .B(n9195), .Z(n9196) );
  AND U9447 ( .A(n9197), .B(n9196), .Z(n9300) );
  NAND U9448 ( .A(n578), .B(n9198), .Z(n9200) );
  XOR U9449 ( .A(a[57]), .B(b[23]), .Z(n9267) );
  NAND U9450 ( .A(n9268), .B(n9267), .Z(n9199) );
  NAND U9451 ( .A(n9200), .B(n9199), .Z(n9301) );
  XNOR U9452 ( .A(n9300), .B(n9301), .Z(n9303) );
  XNOR U9453 ( .A(n9302), .B(n9303), .Z(n9309) );
  XNOR U9454 ( .A(n9309), .B(n9308), .Z(n9311) );
  XNOR U9455 ( .A(n9311), .B(n9310), .Z(n9315) );
  OR U9456 ( .A(n9209), .B(n565), .Z(n9211) );
  XOR U9457 ( .A(b[27]), .B(a[53]), .Z(n9291) );
  NANDN U9458 ( .A(n9692), .B(n9291), .Z(n9210) );
  AND U9459 ( .A(n9211), .B(n9210), .Z(n9279) );
  OR U9460 ( .A(n9212), .B(n559), .Z(n9214) );
  XNOR U9461 ( .A(b[29]), .B(a[51]), .Z(n9264) );
  OR U9462 ( .A(n9264), .B(n9796), .Z(n9213) );
  AND U9463 ( .A(n9214), .B(n9213), .Z(n9277) );
  NAND U9464 ( .A(n577), .B(n9215), .Z(n9218) );
  XOR U9465 ( .A(a[59]), .B(b[21]), .Z(n9285) );
  NAND U9466 ( .A(n9216), .B(n9285), .Z(n9217) );
  NAND U9467 ( .A(n9218), .B(n9217), .Z(n9278) );
  XNOR U9468 ( .A(n9277), .B(n9278), .Z(n9280) );
  XNOR U9469 ( .A(n9279), .B(n9280), .Z(n9305) );
  OR U9470 ( .A(n9219), .B(n580), .Z(n9221) );
  XNOR U9471 ( .A(b[31]), .B(a[49]), .Z(n9294) );
  OR U9472 ( .A(n9294), .B(n9904), .Z(n9220) );
  AND U9473 ( .A(n9221), .B(n9220), .Z(n9281) );
  NAND U9474 ( .A(n579), .B(n9222), .Z(n9224) );
  XOR U9475 ( .A(b[25]), .B(a[55]), .Z(n9261) );
  NAND U9476 ( .A(n9364), .B(n9261), .Z(n9223) );
  NAND U9477 ( .A(n9224), .B(n9223), .Z(n9282) );
  XNOR U9478 ( .A(n9281), .B(n9282), .Z(n9284) );
  AND U9479 ( .A(b[31]), .B(a[47]), .Z(n9271) );
  XOR U9480 ( .A(n9271), .B(n9272), .Z(n9274) );
  XNOR U9481 ( .A(n9225), .B(n9274), .Z(n9283) );
  XNOR U9482 ( .A(n9284), .B(n9283), .Z(n9304) );
  XNOR U9483 ( .A(n9305), .B(n9304), .Z(n9307) );
  IV U9484 ( .A(n9225), .Z(n9273) );
  NAND U9485 ( .A(n9273), .B(n9226), .Z(n9230) );
  OR U9486 ( .A(n9228), .B(n9227), .Z(n9229) );
  NAND U9487 ( .A(n9230), .B(n9229), .Z(n9306) );
  XNOR U9488 ( .A(n9307), .B(n9306), .Z(n9313) );
  NANDN U9489 ( .A(n9232), .B(n9231), .Z(n9236) );
  NANDN U9490 ( .A(n9234), .B(n9233), .Z(n9235) );
  AND U9491 ( .A(n9236), .B(n9235), .Z(n9312) );
  XNOR U9492 ( .A(n9313), .B(n9312), .Z(n9314) );
  XOR U9493 ( .A(n9315), .B(n9314), .Z(n9260) );
  XNOR U9494 ( .A(n9258), .B(n9257), .Z(n9259) );
  XOR U9495 ( .A(n9260), .B(n9259), .Z(n9254) );
  XNOR U9496 ( .A(n9253), .B(n9254), .Z(n9256) );
  XNOR U9497 ( .A(n9255), .B(n9256), .Z(n9247) );
  XNOR U9498 ( .A(n9248), .B(n9247), .Z(n9250) );
  XOR U9499 ( .A(n9249), .B(n9250), .Z(n9245) );
  XOR U9500 ( .A(n9246), .B(n9245), .Z(c[111]) );
  AND U9501 ( .A(n9246), .B(n9245), .Z(n9319) );
  NAND U9502 ( .A(n9248), .B(n9247), .Z(n9252) );
  NANDN U9503 ( .A(n9250), .B(n9249), .Z(n9251) );
  NAND U9504 ( .A(n9252), .B(n9251), .Z(n9322) );
  NANDN U9505 ( .A(n566), .B(n9261), .Z(n9263) );
  XOR U9506 ( .A(b[25]), .B(a[56]), .Z(n9363) );
  NANDN U9507 ( .A(n9684), .B(n9363), .Z(n9262) );
  AND U9508 ( .A(n9263), .B(n9262), .Z(n9349) );
  OR U9509 ( .A(n9264), .B(n559), .Z(n9266) );
  XNOR U9510 ( .A(b[29]), .B(a[52]), .Z(n9351) );
  OR U9511 ( .A(n9351), .B(n9796), .Z(n9265) );
  AND U9512 ( .A(n9266), .B(n9265), .Z(n9347) );
  NAND U9513 ( .A(n578), .B(n9267), .Z(n9270) );
  XOR U9514 ( .A(a[58]), .B(b[23]), .Z(n9354) );
  NAND U9515 ( .A(n9268), .B(n9354), .Z(n9269) );
  NAND U9516 ( .A(n9270), .B(n9269), .Z(n9348) );
  XNOR U9517 ( .A(n9347), .B(n9348), .Z(n9350) );
  XNOR U9518 ( .A(n9349), .B(n9350), .Z(n9335) );
  NANDN U9519 ( .A(n9272), .B(n9271), .Z(n9276) );
  OR U9520 ( .A(n9274), .B(n9273), .Z(n9275) );
  AND U9521 ( .A(n9276), .B(n9275), .Z(n9334) );
  XNOR U9522 ( .A(n9335), .B(n9334), .Z(n9337) );
  XNOR U9523 ( .A(n9337), .B(n9336), .Z(n9384) );
  NANDN U9524 ( .A(n556), .B(n9285), .Z(n9287) );
  XNOR U9525 ( .A(a[60]), .B(b[21]), .Z(n9357) );
  OR U9526 ( .A(n9357), .B(n9480), .Z(n9286) );
  AND U9527 ( .A(n9287), .B(n9286), .Z(n9340) );
  OR U9528 ( .A(n9288), .B(n574), .Z(n9290) );
  XNOR U9529 ( .A(a[62]), .B(b[19]), .Z(n9367) );
  OR U9530 ( .A(n9367), .B(n555), .Z(n9289) );
  AND U9531 ( .A(n9290), .B(n9289), .Z(n9338) );
  NAND U9532 ( .A(n582), .B(n9291), .Z(n9293) );
  XOR U9533 ( .A(b[27]), .B(a[54]), .Z(n9370) );
  NAND U9534 ( .A(n9770), .B(n9370), .Z(n9292) );
  NAND U9535 ( .A(n9293), .B(n9292), .Z(n9339) );
  XNOR U9536 ( .A(n9338), .B(n9339), .Z(n9341) );
  XNOR U9537 ( .A(n9340), .B(n9341), .Z(n9376) );
  OR U9538 ( .A(n9294), .B(n580), .Z(n9296) );
  XNOR U9539 ( .A(b[31]), .B(a[50]), .Z(n9360) );
  OR U9540 ( .A(n9360), .B(n9904), .Z(n9295) );
  NAND U9541 ( .A(n9296), .B(n9295), .Z(n9343) );
  AND U9542 ( .A(b[31]), .B(a[48]), .Z(n9374) );
  OR U9543 ( .A(n9297), .B(n554), .Z(n9298) );
  AND U9544 ( .A(n9299), .B(n9298), .Z(n9342) );
  XNOR U9545 ( .A(n9374), .B(n9342), .Z(n9344) );
  XOR U9546 ( .A(n9343), .B(n9344), .Z(n9375) );
  XNOR U9547 ( .A(n9376), .B(n9375), .Z(n9378) );
  XNOR U9548 ( .A(n9378), .B(n9377), .Z(n9382) );
  XNOR U9549 ( .A(n9381), .B(n9382), .Z(n9383) );
  XNOR U9550 ( .A(n9384), .B(n9383), .Z(n9332) );
  XNOR U9551 ( .A(n9330), .B(n9331), .Z(n9333) );
  XNOR U9552 ( .A(n9332), .B(n9333), .Z(n9327) );
  NANDN U9553 ( .A(n9313), .B(n9312), .Z(n9317) );
  NANDN U9554 ( .A(n9315), .B(n9314), .Z(n9316) );
  AND U9555 ( .A(n9317), .B(n9316), .Z(n9326) );
  XNOR U9556 ( .A(n9327), .B(n9326), .Z(n9328) );
  XOR U9557 ( .A(n9329), .B(n9328), .Z(n9321) );
  XOR U9558 ( .A(n9320), .B(n9321), .Z(n9323) );
  XOR U9559 ( .A(n9322), .B(n9323), .Z(n9318) );
  XOR U9560 ( .A(n9319), .B(n9318), .Z(c[112]) );
  AND U9561 ( .A(n9319), .B(n9318), .Z(n9386) );
  NANDN U9562 ( .A(n9321), .B(n9320), .Z(n9325) );
  NANDN U9563 ( .A(n9323), .B(n9322), .Z(n9324) );
  NAND U9564 ( .A(n9325), .B(n9324), .Z(n9389) );
  IV U9565 ( .A(n9374), .Z(n9419) );
  NANDN U9566 ( .A(n9342), .B(n9419), .Z(n9346) );
  NANDN U9567 ( .A(n9344), .B(n9343), .Z(n9345) );
  NAND U9568 ( .A(n9346), .B(n9345), .Z(n9402) );
  XOR U9569 ( .A(n9401), .B(n9402), .Z(n9404) );
  XNOR U9570 ( .A(n9403), .B(n9404), .Z(n9399) );
  OR U9571 ( .A(n9351), .B(n559), .Z(n9353) );
  XNOR U9572 ( .A(b[29]), .B(a[53]), .Z(n9438) );
  OR U9573 ( .A(n9438), .B(n9796), .Z(n9352) );
  AND U9574 ( .A(n9353), .B(n9352), .Z(n9411) );
  NANDN U9575 ( .A(n563), .B(n9354), .Z(n9356) );
  XNOR U9576 ( .A(a[59]), .B(b[23]), .Z(n9429) );
  OR U9577 ( .A(n9429), .B(n9605), .Z(n9355) );
  AND U9578 ( .A(n9356), .B(n9355), .Z(n9409) );
  OR U9579 ( .A(n9357), .B(n556), .Z(n9359) );
  XNOR U9580 ( .A(a[61]), .B(b[21]), .Z(n9432) );
  OR U9581 ( .A(n9432), .B(n9480), .Z(n9358) );
  AND U9582 ( .A(n9359), .B(n9358), .Z(n9446) );
  OR U9583 ( .A(n9360), .B(n580), .Z(n9362) );
  XNOR U9584 ( .A(b[31]), .B(a[51]), .Z(n9423) );
  OR U9585 ( .A(n9423), .B(n9904), .Z(n9361) );
  AND U9586 ( .A(n9362), .B(n9361), .Z(n9444) );
  NAND U9587 ( .A(n579), .B(n9363), .Z(n9366) );
  XOR U9588 ( .A(b[25]), .B(a[57]), .Z(n9435) );
  NAND U9589 ( .A(n9364), .B(n9435), .Z(n9365) );
  NAND U9590 ( .A(n9366), .B(n9365), .Z(n9445) );
  XNOR U9591 ( .A(n9444), .B(n9445), .Z(n9447) );
  XNOR U9592 ( .A(n9446), .B(n9447), .Z(n9410) );
  XNOR U9593 ( .A(n9409), .B(n9410), .Z(n9412) );
  XNOR U9594 ( .A(n9411), .B(n9412), .Z(n9406) );
  OR U9595 ( .A(n9367), .B(n574), .Z(n9369) );
  XNOR U9596 ( .A(a[63]), .B(b[19]), .Z(n9426) );
  OR U9597 ( .A(n9426), .B(n555), .Z(n9368) );
  AND U9598 ( .A(n9369), .B(n9368), .Z(n9413) );
  NAND U9599 ( .A(n582), .B(n9370), .Z(n9372) );
  XOR U9600 ( .A(b[27]), .B(a[55]), .Z(n9441) );
  NAND U9601 ( .A(n9770), .B(n9441), .Z(n9371) );
  NAND U9602 ( .A(n9372), .B(n9371), .Z(n9414) );
  XNOR U9603 ( .A(n9413), .B(n9414), .Z(n9416) );
  AND U9604 ( .A(b[31]), .B(a[49]), .Z(n9417) );
  IV U9605 ( .A(n9373), .Z(n9418) );
  XNOR U9606 ( .A(n9417), .B(n9418), .Z(n9420) );
  XNOR U9607 ( .A(n9374), .B(n9420), .Z(n9415) );
  XNOR U9608 ( .A(n9416), .B(n9415), .Z(n9405) );
  XNOR U9609 ( .A(n9406), .B(n9405), .Z(n9408) );
  XNOR U9610 ( .A(n9407), .B(n9408), .Z(n9398) );
  NANDN U9611 ( .A(n9376), .B(n9375), .Z(n9380) );
  NAND U9612 ( .A(n9378), .B(n9377), .Z(n9379) );
  NAND U9613 ( .A(n9380), .B(n9379), .Z(n9397) );
  XNOR U9614 ( .A(n9398), .B(n9397), .Z(n9400) );
  XNOR U9615 ( .A(n9399), .B(n9400), .Z(n9392) );
  XOR U9616 ( .A(n9392), .B(n9391), .Z(n9394) );
  XOR U9617 ( .A(n9393), .B(n9394), .Z(n9388) );
  XOR U9618 ( .A(n9387), .B(n9388), .Z(n9390) );
  XOR U9619 ( .A(n9389), .B(n9390), .Z(n9385) );
  XOR U9620 ( .A(n9386), .B(n9385), .Z(c[113]) );
  AND U9621 ( .A(n9386), .B(n9385), .Z(n9449) );
  NANDN U9622 ( .A(n9392), .B(n9391), .Z(n9396) );
  NANDN U9623 ( .A(n9394), .B(n9393), .Z(n9395) );
  AND U9624 ( .A(n9396), .B(n9395), .Z(n9451) );
  NAND U9625 ( .A(n9418), .B(n9417), .Z(n9422) );
  OR U9626 ( .A(n9420), .B(n9419), .Z(n9421) );
  AND U9627 ( .A(n9422), .B(n9421), .Z(n9491) );
  OR U9628 ( .A(n9423), .B(n580), .Z(n9425) );
  XOR U9629 ( .A(b[31]), .B(a[52]), .Z(n9476) );
  NANDN U9630 ( .A(n9904), .B(n9476), .Z(n9424) );
  AND U9631 ( .A(n9425), .B(n9424), .Z(n9465) );
  OR U9632 ( .A(n9426), .B(n574), .Z(n9427) );
  AND U9633 ( .A(n9428), .B(n9427), .Z(n9464) );
  NAND U9634 ( .A(b[31]), .B(a[50]), .Z(n9486) );
  XNOR U9635 ( .A(n9464), .B(n9486), .Z(n9466) );
  XNOR U9636 ( .A(n9465), .B(n9466), .Z(n9492) );
  XNOR U9637 ( .A(n9491), .B(n9492), .Z(n9494) );
  XNOR U9638 ( .A(n9493), .B(n9494), .Z(n9497) );
  OR U9639 ( .A(n9429), .B(n563), .Z(n9431) );
  XNOR U9640 ( .A(a[60]), .B(b[23]), .Z(n9473) );
  OR U9641 ( .A(n9473), .B(n9605), .Z(n9430) );
  AND U9642 ( .A(n9431), .B(n9430), .Z(n9489) );
  OR U9643 ( .A(n9432), .B(n556), .Z(n9434) );
  XNOR U9644 ( .A(a[62]), .B(b[21]), .Z(n9479) );
  OR U9645 ( .A(n9479), .B(n9480), .Z(n9433) );
  AND U9646 ( .A(n9434), .B(n9433), .Z(n9487) );
  NANDN U9647 ( .A(n566), .B(n9435), .Z(n9437) );
  XNOR U9648 ( .A(a[58]), .B(b[25]), .Z(n9470) );
  OR U9649 ( .A(n9470), .B(n9684), .Z(n9436) );
  AND U9650 ( .A(n9437), .B(n9436), .Z(n9462) );
  OR U9651 ( .A(n9438), .B(n559), .Z(n9440) );
  XNOR U9652 ( .A(b[29]), .B(a[54]), .Z(n9467) );
  OR U9653 ( .A(n9467), .B(n9796), .Z(n9439) );
  AND U9654 ( .A(n9440), .B(n9439), .Z(n9460) );
  NAND U9655 ( .A(n582), .B(n9441), .Z(n9443) );
  XOR U9656 ( .A(b[27]), .B(a[56]), .Z(n9483) );
  NAND U9657 ( .A(n9770), .B(n9483), .Z(n9442) );
  NAND U9658 ( .A(n9443), .B(n9442), .Z(n9461) );
  XNOR U9659 ( .A(n9460), .B(n9461), .Z(n9463) );
  XNOR U9660 ( .A(n9462), .B(n9463), .Z(n9488) );
  XNOR U9661 ( .A(n9487), .B(n9488), .Z(n9490) );
  XNOR U9662 ( .A(n9489), .B(n9490), .Z(n9496) );
  XOR U9663 ( .A(n9496), .B(n9495), .Z(n9498) );
  XNOR U9664 ( .A(n9497), .B(n9498), .Z(n9501) );
  XNOR U9665 ( .A(n9502), .B(n9501), .Z(n9503) );
  XNOR U9666 ( .A(n9504), .B(n9503), .Z(n9456) );
  XNOR U9667 ( .A(n9457), .B(n9456), .Z(n9459) );
  XNOR U9668 ( .A(n9458), .B(n9459), .Z(n9450) );
  XNOR U9669 ( .A(n9451), .B(n9450), .Z(n9453) );
  XOR U9670 ( .A(n9452), .B(n9453), .Z(n9448) );
  XOR U9671 ( .A(n9449), .B(n9448), .Z(c[114]) );
  AND U9672 ( .A(n9449), .B(n9448), .Z(n9506) );
  NAND U9673 ( .A(n9451), .B(n9450), .Z(n9455) );
  NANDN U9674 ( .A(n9453), .B(n9452), .Z(n9454) );
  NAND U9675 ( .A(n9455), .B(n9454), .Z(n9509) );
  XNOR U9676 ( .A(n9558), .B(n9559), .Z(n9561) );
  OR U9677 ( .A(n9467), .B(n559), .Z(n9469) );
  XNOR U9678 ( .A(b[29]), .B(a[55]), .Z(n9551) );
  OR U9679 ( .A(n9551), .B(n9796), .Z(n9468) );
  AND U9680 ( .A(n9469), .B(n9468), .Z(n9554) );
  OR U9681 ( .A(n9470), .B(n566), .Z(n9472) );
  XNOR U9682 ( .A(a[59]), .B(b[25]), .Z(n9542) );
  OR U9683 ( .A(n9542), .B(n9684), .Z(n9471) );
  AND U9684 ( .A(n9472), .B(n9471), .Z(n9534) );
  OR U9685 ( .A(n9473), .B(n563), .Z(n9475) );
  XNOR U9686 ( .A(a[61]), .B(b[23]), .Z(n9545) );
  OR U9687 ( .A(n9545), .B(n9605), .Z(n9474) );
  AND U9688 ( .A(n9475), .B(n9474), .Z(n9532) );
  NAND U9689 ( .A(n9764), .B(n9476), .Z(n9478) );
  XOR U9690 ( .A(b[31]), .B(a[53]), .Z(n9536) );
  NAND U9691 ( .A(n584), .B(n9536), .Z(n9477) );
  NAND U9692 ( .A(n9478), .B(n9477), .Z(n9533) );
  XNOR U9693 ( .A(n9532), .B(n9533), .Z(n9535) );
  XNOR U9694 ( .A(n9534), .B(n9535), .Z(n9555) );
  XNOR U9695 ( .A(n9554), .B(n9555), .Z(n9557) );
  OR U9696 ( .A(n9479), .B(n556), .Z(n9482) );
  XNOR U9697 ( .A(a[63]), .B(b[21]), .Z(n9539) );
  OR U9698 ( .A(n9539), .B(n9480), .Z(n9481) );
  AND U9699 ( .A(n9482), .B(n9481), .Z(n9525) );
  NAND U9700 ( .A(n582), .B(n9483), .Z(n9485) );
  XOR U9701 ( .A(b[27]), .B(a[57]), .Z(n9548) );
  NAND U9702 ( .A(n9770), .B(n9548), .Z(n9484) );
  NAND U9703 ( .A(n9485), .B(n9484), .Z(n9526) );
  XNOR U9704 ( .A(n9525), .B(n9526), .Z(n9528) );
  IV U9705 ( .A(n9486), .Z(n9524) );
  AND U9706 ( .A(b[31]), .B(a[51]), .Z(n9522) );
  XNOR U9707 ( .A(n9522), .B(n9521), .Z(n9523) );
  XNOR U9708 ( .A(n9524), .B(n9523), .Z(n9529) );
  XNOR U9709 ( .A(n9528), .B(n9529), .Z(n9556) );
  XNOR U9710 ( .A(n9557), .B(n9556), .Z(n9560) );
  XNOR U9711 ( .A(n9561), .B(n9560), .Z(n9520) );
  XNOR U9712 ( .A(n9518), .B(n9517), .Z(n9519) );
  XNOR U9713 ( .A(n9520), .B(n9519), .Z(n9513) );
  NANDN U9714 ( .A(n9496), .B(n9495), .Z(n9500) );
  OR U9715 ( .A(n9498), .B(n9497), .Z(n9499) );
  AND U9716 ( .A(n9500), .B(n9499), .Z(n9514) );
  XNOR U9717 ( .A(n9513), .B(n9514), .Z(n9516) );
  XNOR U9718 ( .A(n9516), .B(n9515), .Z(n9508) );
  XOR U9719 ( .A(n9507), .B(n9508), .Z(n9510) );
  XOR U9720 ( .A(n9509), .B(n9510), .Z(n9505) );
  XOR U9721 ( .A(n9506), .B(n9505), .Z(c[115]) );
  AND U9722 ( .A(n9506), .B(n9505), .Z(n9563) );
  NANDN U9723 ( .A(n9508), .B(n9507), .Z(n9512) );
  NANDN U9724 ( .A(n9510), .B(n9509), .Z(n9511) );
  NAND U9725 ( .A(n9512), .B(n9511), .Z(n9566) );
  IV U9726 ( .A(n9525), .Z(n9527) );
  NAND U9727 ( .A(n9527), .B(n9526), .Z(n9531) );
  NANDN U9728 ( .A(n9529), .B(n9528), .Z(n9530) );
  NAND U9729 ( .A(n9531), .B(n9530), .Z(n9578) );
  XNOR U9730 ( .A(n9579), .B(n9578), .Z(n9581) );
  XNOR U9731 ( .A(n9581), .B(n9580), .Z(n9577) );
  NANDN U9732 ( .A(n580), .B(n9536), .Z(n9538) );
  XOR U9733 ( .A(b[31]), .B(a[54]), .Z(n9601) );
  NANDN U9734 ( .A(n9904), .B(n9601), .Z(n9537) );
  AND U9735 ( .A(n9538), .B(n9537), .Z(n9589) );
  OR U9736 ( .A(n9539), .B(n556), .Z(n9540) );
  AND U9737 ( .A(n9541), .B(n9540), .Z(n9588) );
  NAND U9738 ( .A(b[31]), .B(a[52]), .Z(n9611) );
  XNOR U9739 ( .A(n9588), .B(n9611), .Z(n9590) );
  XNOR U9740 ( .A(n9589), .B(n9590), .Z(n9585) );
  OR U9741 ( .A(n9542), .B(n566), .Z(n9544) );
  XNOR U9742 ( .A(a[60]), .B(b[25]), .Z(n9595) );
  OR U9743 ( .A(n9595), .B(n9684), .Z(n9543) );
  AND U9744 ( .A(n9544), .B(n9543), .Z(n9593) );
  OR U9745 ( .A(n9545), .B(n563), .Z(n9547) );
  XNOR U9746 ( .A(a[62]), .B(b[23]), .Z(n9604) );
  OR U9747 ( .A(n9604), .B(n9605), .Z(n9546) );
  AND U9748 ( .A(n9547), .B(n9546), .Z(n9591) );
  NAND U9749 ( .A(n582), .B(n9548), .Z(n9550) );
  XOR U9750 ( .A(b[27]), .B(a[58]), .Z(n9608) );
  NAND U9751 ( .A(n9770), .B(n9608), .Z(n9549) );
  NAND U9752 ( .A(n9550), .B(n9549), .Z(n9592) );
  XNOR U9753 ( .A(n9591), .B(n9592), .Z(n9594) );
  XNOR U9754 ( .A(n9593), .B(n9594), .Z(n9583) );
  OR U9755 ( .A(n9551), .B(n559), .Z(n9553) );
  XNOR U9756 ( .A(b[29]), .B(a[56]), .Z(n9598) );
  OR U9757 ( .A(n9598), .B(n9796), .Z(n9552) );
  AND U9758 ( .A(n9553), .B(n9552), .Z(n9582) );
  XNOR U9759 ( .A(n9583), .B(n9582), .Z(n9584) );
  XNOR U9760 ( .A(n9585), .B(n9584), .Z(n9574) );
  XNOR U9761 ( .A(n9574), .B(n9575), .Z(n9576) );
  XNOR U9762 ( .A(n9577), .B(n9576), .Z(n9570) );
  XNOR U9763 ( .A(n9570), .B(n9571), .Z(n9573) );
  XNOR U9764 ( .A(n9572), .B(n9573), .Z(n9564) );
  XNOR U9765 ( .A(n9565), .B(n9564), .Z(n9567) );
  XOR U9766 ( .A(n9566), .B(n9567), .Z(n9562) );
  XOR U9767 ( .A(n9563), .B(n9562), .Z(c[116]) );
  AND U9768 ( .A(n9563), .B(n9562), .Z(n9613) );
  NAND U9769 ( .A(n9565), .B(n9564), .Z(n9569) );
  NANDN U9770 ( .A(n9567), .B(n9566), .Z(n9568) );
  NAND U9771 ( .A(n9569), .B(n9568), .Z(n9616) );
  NANDN U9772 ( .A(n9583), .B(n9582), .Z(n9587) );
  NANDN U9773 ( .A(n9585), .B(n9584), .Z(n9586) );
  AND U9774 ( .A(n9587), .B(n9586), .Z(n9624) );
  OR U9775 ( .A(n9595), .B(n566), .Z(n9597) );
  XNOR U9776 ( .A(a[61]), .B(b[25]), .Z(n9635) );
  OR U9777 ( .A(n9635), .B(n9684), .Z(n9596) );
  AND U9778 ( .A(n9597), .B(n9596), .Z(n9649) );
  OR U9779 ( .A(n9598), .B(n559), .Z(n9600) );
  XOR U9780 ( .A(b[29]), .B(a[57]), .Z(n9638) );
  NANDN U9781 ( .A(n9796), .B(n9638), .Z(n9599) );
  AND U9782 ( .A(n9600), .B(n9599), .Z(n9647) );
  NAND U9783 ( .A(n9764), .B(n9601), .Z(n9603) );
  XOR U9784 ( .A(b[31]), .B(a[55]), .Z(n9641) );
  NAND U9785 ( .A(n584), .B(n9641), .Z(n9602) );
  NAND U9786 ( .A(n9603), .B(n9602), .Z(n9648) );
  XNOR U9787 ( .A(n9647), .B(n9648), .Z(n9650) );
  XNOR U9788 ( .A(n9649), .B(n9650), .Z(n9627) );
  OR U9789 ( .A(n9604), .B(n563), .Z(n9607) );
  XNOR U9790 ( .A(a[63]), .B(b[23]), .Z(n9644) );
  OR U9791 ( .A(n9644), .B(n9605), .Z(n9606) );
  AND U9792 ( .A(n9607), .B(n9606), .Z(n9655) );
  NAND U9793 ( .A(n582), .B(n9608), .Z(n9610) );
  XOR U9794 ( .A(b[27]), .B(a[59]), .Z(n9632) );
  NAND U9795 ( .A(n9770), .B(n9632), .Z(n9609) );
  NAND U9796 ( .A(n9610), .B(n9609), .Z(n9656) );
  XNOR U9797 ( .A(n9655), .B(n9656), .Z(n9658) );
  IV U9798 ( .A(n9611), .Z(n9652) );
  XNOR U9799 ( .A(n9652), .B(n9651), .Z(n9654) );
  NAND U9800 ( .A(b[31]), .B(a[53]), .Z(n9653) );
  XNOR U9801 ( .A(n9654), .B(n9653), .Z(n9657) );
  XNOR U9802 ( .A(n9658), .B(n9657), .Z(n9626) );
  XNOR U9803 ( .A(n9627), .B(n9626), .Z(n9628) );
  XNOR U9804 ( .A(n9629), .B(n9628), .Z(n9622) );
  XNOR U9805 ( .A(n9623), .B(n9622), .Z(n9625) );
  XNOR U9806 ( .A(n9624), .B(n9625), .Z(n9619) );
  XNOR U9807 ( .A(n9618), .B(n9619), .Z(n9620) );
  XNOR U9808 ( .A(n9621), .B(n9620), .Z(n9614) );
  XOR U9809 ( .A(n9615), .B(n9614), .Z(n9617) );
  XOR U9810 ( .A(n9616), .B(n9617), .Z(n9612) );
  XOR U9811 ( .A(n9613), .B(n9612), .Z(c[117]) );
  AND U9812 ( .A(n9613), .B(n9612), .Z(n9660) );
  NANDN U9813 ( .A(n9627), .B(n9626), .Z(n9631) );
  NAND U9814 ( .A(n9629), .B(n9628), .Z(n9630) );
  AND U9815 ( .A(n9631), .B(n9630), .Z(n9667) );
  NANDN U9816 ( .A(n565), .B(n9632), .Z(n9634) );
  XNOR U9817 ( .A(b[27]), .B(a[60]), .Z(n9691) );
  OR U9818 ( .A(n9691), .B(n9692), .Z(n9633) );
  AND U9819 ( .A(n9634), .B(n9633), .Z(n9681) );
  OR U9820 ( .A(n9635), .B(n566), .Z(n9637) );
  XNOR U9821 ( .A(a[62]), .B(b[25]), .Z(n9683) );
  OR U9822 ( .A(n9683), .B(n9684), .Z(n9636) );
  AND U9823 ( .A(n9637), .B(n9636), .Z(n9679) );
  NAND U9824 ( .A(n583), .B(n9638), .Z(n9640) );
  XOR U9825 ( .A(b[29]), .B(a[58]), .Z(n9687) );
  NAND U9826 ( .A(n581), .B(n9687), .Z(n9639) );
  NAND U9827 ( .A(n9640), .B(n9639), .Z(n9680) );
  XNOR U9828 ( .A(n9679), .B(n9680), .Z(n9682) );
  XNOR U9829 ( .A(n9681), .B(n9682), .Z(n9676) );
  NANDN U9830 ( .A(n580), .B(n9641), .Z(n9643) );
  XOR U9831 ( .A(b[31]), .B(a[56]), .Z(n9695) );
  NANDN U9832 ( .A(n9904), .B(n9695), .Z(n9642) );
  NAND U9833 ( .A(n9643), .B(n9642), .Z(n9699) );
  AND U9834 ( .A(b[31]), .B(a[54]), .Z(n9726) );
  OR U9835 ( .A(n9644), .B(n563), .Z(n9645) );
  AND U9836 ( .A(n9646), .B(n9645), .Z(n9698) );
  XNOR U9837 ( .A(n9726), .B(n9698), .Z(n9700) );
  XOR U9838 ( .A(n9699), .B(n9700), .Z(n9675) );
  XNOR U9839 ( .A(n9676), .B(n9675), .Z(n9678) );
  XNOR U9840 ( .A(n9678), .B(n9677), .Z(n9674) );
  XNOR U9841 ( .A(n9671), .B(n9672), .Z(n9673) );
  XOR U9842 ( .A(n9674), .B(n9673), .Z(n9668) );
  XOR U9843 ( .A(n9667), .B(n9668), .Z(n9670) );
  XOR U9844 ( .A(n9669), .B(n9670), .Z(n9662) );
  XOR U9845 ( .A(n9661), .B(n9662), .Z(n9664) );
  XOR U9846 ( .A(n9663), .B(n9664), .Z(n9659) );
  XOR U9847 ( .A(n9660), .B(n9659), .Z(c[118]) );
  AND U9848 ( .A(n9660), .B(n9659), .Z(n9702) );
  NANDN U9849 ( .A(n9662), .B(n9661), .Z(n9666) );
  NANDN U9850 ( .A(n9664), .B(n9663), .Z(n9665) );
  NAND U9851 ( .A(n9666), .B(n9665), .Z(n9705) );
  OR U9852 ( .A(n9683), .B(n566), .Z(n9686) );
  XNOR U9853 ( .A(a[63]), .B(b[25]), .Z(n9738) );
  OR U9854 ( .A(n9738), .B(n9684), .Z(n9685) );
  AND U9855 ( .A(n9686), .B(n9685), .Z(n9741) );
  NAND U9856 ( .A(n583), .B(n9687), .Z(n9689) );
  XOR U9857 ( .A(b[29]), .B(a[59]), .Z(n9729) );
  NAND U9858 ( .A(n581), .B(n9729), .Z(n9688) );
  NAND U9859 ( .A(n9689), .B(n9688), .Z(n9742) );
  XNOR U9860 ( .A(n9741), .B(n9742), .Z(n9743) );
  AND U9861 ( .A(b[31]), .B(a[55]), .Z(n9723) );
  XNOR U9862 ( .A(n9723), .B(n9690), .Z(n9725) );
  XNOR U9863 ( .A(n9726), .B(n9725), .Z(n9744) );
  XNOR U9864 ( .A(n9743), .B(n9744), .Z(n9719) );
  OR U9865 ( .A(n9691), .B(n565), .Z(n9694) );
  XOR U9866 ( .A(b[27]), .B(a[61]), .Z(n9732) );
  NANDN U9867 ( .A(n9692), .B(n9732), .Z(n9693) );
  AND U9868 ( .A(n9694), .B(n9693), .Z(n9720) );
  XNOR U9869 ( .A(n9719), .B(n9720), .Z(n9722) );
  NAND U9870 ( .A(n9764), .B(n9695), .Z(n9697) );
  XOR U9871 ( .A(b[31]), .B(a[57]), .Z(n9735) );
  NAND U9872 ( .A(n584), .B(n9735), .Z(n9696) );
  NAND U9873 ( .A(n9697), .B(n9696), .Z(n9721) );
  XNOR U9874 ( .A(n9722), .B(n9721), .Z(n9714) );
  XOR U9875 ( .A(n9714), .B(n9713), .Z(n9716) );
  XOR U9876 ( .A(n9715), .B(n9716), .Z(n9710) );
  XNOR U9877 ( .A(n9709), .B(n9710), .Z(n9712) );
  XNOR U9878 ( .A(n9711), .B(n9712), .Z(n9704) );
  XOR U9879 ( .A(n9703), .B(n9704), .Z(n9706) );
  XOR U9880 ( .A(n9705), .B(n9706), .Z(n9701) );
  XOR U9881 ( .A(n9702), .B(n9701), .Z(c[119]) );
  AND U9882 ( .A(n9702), .B(n9701), .Z(n9746) );
  NANDN U9883 ( .A(n9704), .B(n9703), .Z(n9708) );
  NANDN U9884 ( .A(n9706), .B(n9705), .Z(n9707) );
  NAND U9885 ( .A(n9708), .B(n9707), .Z(n9749) );
  NANDN U9886 ( .A(n9714), .B(n9713), .Z(n9718) );
  NANDN U9887 ( .A(n9716), .B(n9715), .Z(n9717) );
  AND U9888 ( .A(n9718), .B(n9717), .Z(n9755) );
  NAND U9889 ( .A(n9724), .B(n9723), .Z(n9728) );
  NAND U9890 ( .A(n9726), .B(n9725), .Z(n9727) );
  AND U9891 ( .A(n9728), .B(n9727), .Z(n9775) );
  NANDN U9892 ( .A(n559), .B(n9729), .Z(n9731) );
  XNOR U9893 ( .A(b[29]), .B(a[60]), .Z(n9760) );
  OR U9894 ( .A(n9760), .B(n9796), .Z(n9730) );
  AND U9895 ( .A(n9731), .B(n9730), .Z(n9773) );
  NAND U9896 ( .A(n582), .B(n9732), .Z(n9734) );
  XOR U9897 ( .A(a[62]), .B(b[27]), .Z(n9769) );
  NAND U9898 ( .A(n9770), .B(n9769), .Z(n9733) );
  NAND U9899 ( .A(n9734), .B(n9733), .Z(n9774) );
  XNOR U9900 ( .A(n9773), .B(n9774), .Z(n9776) );
  XNOR U9901 ( .A(n9775), .B(n9776), .Z(n9779) );
  NANDN U9902 ( .A(n580), .B(n9735), .Z(n9737) );
  XOR U9903 ( .A(b[31]), .B(a[58]), .Z(n9763) );
  NANDN U9904 ( .A(n9904), .B(n9763), .Z(n9736) );
  AND U9905 ( .A(n9737), .B(n9736), .Z(n9758) );
  OR U9906 ( .A(n9738), .B(n566), .Z(n9739) );
  AND U9907 ( .A(n9740), .B(n9739), .Z(n9757) );
  NAND U9908 ( .A(b[31]), .B(a[56]), .Z(n9767) );
  XNOR U9909 ( .A(n9757), .B(n9767), .Z(n9759) );
  XNOR U9910 ( .A(n9758), .B(n9759), .Z(n9778) );
  XOR U9911 ( .A(n9778), .B(n9777), .Z(n9780) );
  XNOR U9912 ( .A(n9779), .B(n9780), .Z(n9753) );
  XOR U9913 ( .A(n9754), .B(n9753), .Z(n9756) );
  XNOR U9914 ( .A(n9755), .B(n9756), .Z(n9747) );
  XNOR U9915 ( .A(n9748), .B(n9747), .Z(n9750) );
  XOR U9916 ( .A(n9749), .B(n9750), .Z(n9745) );
  XOR U9917 ( .A(n9746), .B(n9745), .Z(c[120]) );
  AND U9918 ( .A(n9746), .B(n9745), .Z(n9784) );
  NAND U9919 ( .A(n9748), .B(n9747), .Z(n9752) );
  NANDN U9920 ( .A(n9750), .B(n9749), .Z(n9751) );
  NAND U9921 ( .A(n9752), .B(n9751), .Z(n9787) );
  OR U9922 ( .A(n9760), .B(n559), .Z(n9762) );
  XNOR U9923 ( .A(b[29]), .B(a[61]), .Z(n9795) );
  OR U9924 ( .A(n9795), .B(n9796), .Z(n9761) );
  AND U9925 ( .A(n9762), .B(n9761), .Z(n9810) );
  NAND U9926 ( .A(n9764), .B(n9763), .Z(n9766) );
  XOR U9927 ( .A(b[31]), .B(a[59]), .Z(n9805) );
  NAND U9928 ( .A(n584), .B(n9805), .Z(n9765) );
  NAND U9929 ( .A(n9766), .B(n9765), .Z(n9811) );
  XNOR U9930 ( .A(n9810), .B(n9811), .Z(n9812) );
  IV U9931 ( .A(n9767), .Z(n9802) );
  AND U9932 ( .A(b[31]), .B(a[57]), .Z(n9799) );
  XNOR U9933 ( .A(n9799), .B(n9768), .Z(n9801) );
  XNOR U9934 ( .A(n9802), .B(n9801), .Z(n9813) );
  XOR U9935 ( .A(n9812), .B(n9813), .Z(n9792) );
  NAND U9936 ( .A(n582), .B(n9769), .Z(n9772) );
  XOR U9937 ( .A(a[63]), .B(b[27]), .Z(n9808) );
  NAND U9938 ( .A(n9808), .B(n9770), .Z(n9771) );
  NAND U9939 ( .A(n9772), .B(n9771), .Z(n9791) );
  XOR U9940 ( .A(n9792), .B(n9791), .Z(n9794) );
  XNOR U9941 ( .A(n9793), .B(n9794), .Z(n9814) );
  XNOR U9942 ( .A(n9814), .B(n9815), .Z(n9817) );
  NANDN U9943 ( .A(n9778), .B(n9777), .Z(n9782) );
  OR U9944 ( .A(n9780), .B(n9779), .Z(n9781) );
  NAND U9945 ( .A(n9782), .B(n9781), .Z(n9816) );
  XNOR U9946 ( .A(n9817), .B(n9816), .Z(n9786) );
  XOR U9947 ( .A(n9785), .B(n9786), .Z(n9788) );
  XOR U9948 ( .A(n9787), .B(n9788), .Z(n9783) );
  XOR U9949 ( .A(n9784), .B(n9783), .Z(c[121]) );
  AND U9950 ( .A(n9784), .B(n9783), .Z(n9819) );
  NANDN U9951 ( .A(n9786), .B(n9785), .Z(n9790) );
  NANDN U9952 ( .A(n9788), .B(n9787), .Z(n9789) );
  NAND U9953 ( .A(n9790), .B(n9789), .Z(n9822) );
  OR U9954 ( .A(n9795), .B(n559), .Z(n9798) );
  XOR U9955 ( .A(b[29]), .B(a[62]), .Z(n9836) );
  NANDN U9956 ( .A(n9796), .B(n9836), .Z(n9797) );
  AND U9957 ( .A(n9798), .B(n9797), .Z(n9826) );
  NAND U9958 ( .A(n9800), .B(n9799), .Z(n9804) );
  NAND U9959 ( .A(n9802), .B(n9801), .Z(n9803) );
  NAND U9960 ( .A(n9804), .B(n9803), .Z(n9827) );
  XNOR U9961 ( .A(n9826), .B(n9827), .Z(n9828) );
  NANDN U9962 ( .A(n580), .B(n9805), .Z(n9807) );
  XNOR U9963 ( .A(b[31]), .B(a[60]), .Z(n9833) );
  OR U9964 ( .A(n9833), .B(n9904), .Z(n9806) );
  NAND U9965 ( .A(n9807), .B(n9806), .Z(n9831) );
  AND U9966 ( .A(b[31]), .B(a[58]), .Z(n9858) );
  XNOR U9967 ( .A(n9858), .B(n9830), .Z(n9832) );
  XOR U9968 ( .A(n9831), .B(n9832), .Z(n9829) );
  XNOR U9969 ( .A(n9828), .B(n9829), .Z(n9839) );
  XNOR U9970 ( .A(n9839), .B(n9840), .Z(n9842) );
  XNOR U9971 ( .A(n9841), .B(n9842), .Z(n9821) );
  XNOR U9972 ( .A(n9821), .B(n9820), .Z(n9823) );
  XOR U9973 ( .A(n9822), .B(n9823), .Z(n9818) );
  XOR U9974 ( .A(n9819), .B(n9818), .Z(c[122]) );
  AND U9975 ( .A(n9819), .B(n9818), .Z(n9844) );
  NAND U9976 ( .A(n9821), .B(n9820), .Z(n9825) );
  NANDN U9977 ( .A(n9823), .B(n9822), .Z(n9824) );
  NAND U9978 ( .A(n9825), .B(n9824), .Z(n9847) );
  OR U9979 ( .A(n9833), .B(n580), .Z(n9835) );
  XNOR U9980 ( .A(b[31]), .B(a[61]), .Z(n9859) );
  OR U9981 ( .A(n9859), .B(n9904), .Z(n9834) );
  AND U9982 ( .A(n9835), .B(n9834), .Z(n9851) );
  XOR U9983 ( .A(a[63]), .B(b[29]), .Z(n9862) );
  NAND U9984 ( .A(n581), .B(n9862), .Z(n9838) );
  NAND U9985 ( .A(n583), .B(n9836), .Z(n9837) );
  NAND U9986 ( .A(n9838), .B(n9837), .Z(n9852) );
  XNOR U9987 ( .A(n9851), .B(n9852), .Z(n9853) );
  AND U9988 ( .A(b[31]), .B(a[59]), .Z(n9856) );
  XNOR U9989 ( .A(n9856), .B(n9855), .Z(n9857) );
  XNOR U9990 ( .A(n9858), .B(n9857), .Z(n9854) );
  XNOR U9991 ( .A(n9853), .B(n9854), .Z(n9867) );
  XNOR U9992 ( .A(n9866), .B(n9867), .Z(n9869) );
  XNOR U9993 ( .A(n9868), .B(n9869), .Z(n9846) );
  XOR U9994 ( .A(n9846), .B(n9845), .Z(n9848) );
  XOR U9995 ( .A(n9847), .B(n9848), .Z(n9843) );
  XOR U9996 ( .A(n9844), .B(n9843), .Z(c[123]) );
  AND U9997 ( .A(n9844), .B(n9843), .Z(n9871) );
  NANDN U9998 ( .A(n9846), .B(n9845), .Z(n9850) );
  NANDN U9999 ( .A(n9848), .B(n9847), .Z(n9849) );
  NAND U10000 ( .A(n9850), .B(n9849), .Z(n9874) );
  OR U10001 ( .A(n9859), .B(n580), .Z(n9861) );
  XNOR U10002 ( .A(b[31]), .B(a[62]), .Z(n9878) );
  OR U10003 ( .A(n9878), .B(n9904), .Z(n9860) );
  NAND U10004 ( .A(n9861), .B(n9860), .Z(n9883) );
  AND U10005 ( .A(b[31]), .B(a[60]), .Z(n9907) );
  AND U10006 ( .A(n9862), .B(n583), .Z(n9865) );
  XOR U10007 ( .A(b[28]), .B(b[27]), .Z(n9863) );
  NAND U10008 ( .A(b[29]), .B(n9863), .Z(n9864) );
  NANDN U10009 ( .A(n9865), .B(n9864), .Z(n9881) );
  XNOR U10010 ( .A(n9907), .B(n9881), .Z(n9884) );
  XOR U10011 ( .A(n9883), .B(n9884), .Z(n9888) );
  XNOR U10012 ( .A(n9887), .B(n9888), .Z(n9890) );
  XNOR U10013 ( .A(n9889), .B(n9890), .Z(n9873) );
  XOR U10014 ( .A(n9873), .B(n9872), .Z(n9875) );
  XOR U10015 ( .A(n9874), .B(n9875), .Z(n9870) );
  XOR U10016 ( .A(n9871), .B(n9870), .Z(c[124]) );
  AND U10017 ( .A(n9871), .B(n9870), .Z(n9914) );
  NANDN U10018 ( .A(n9873), .B(n9872), .Z(n9877) );
  NANDN U10019 ( .A(n9875), .B(n9874), .Z(n9876) );
  NAND U10020 ( .A(n9877), .B(n9876), .Z(n9893) );
  AND U10021 ( .A(b[31]), .B(a[61]), .Z(n9910) );
  XOR U10022 ( .A(n9909), .B(n9910), .Z(n9908) );
  IV U10023 ( .A(n9907), .Z(n9882) );
  XNOR U10024 ( .A(n9908), .B(n9882), .Z(n9898) );
  OR U10025 ( .A(n9878), .B(n580), .Z(n9880) );
  XNOR U10026 ( .A(a[63]), .B(b[31]), .Z(n9903) );
  OR U10027 ( .A(n9903), .B(n9904), .Z(n9879) );
  NAND U10028 ( .A(n9880), .B(n9879), .Z(n9897) );
  XOR U10029 ( .A(n9898), .B(n9897), .Z(n9900) );
  NAND U10030 ( .A(n9882), .B(n9881), .Z(n9886) );
  NAND U10031 ( .A(n9884), .B(n9883), .Z(n9885) );
  NAND U10032 ( .A(n9886), .B(n9885), .Z(n9899) );
  XOR U10033 ( .A(n9900), .B(n9899), .Z(n9892) );
  XOR U10034 ( .A(n9892), .B(n9891), .Z(n9894) );
  XOR U10035 ( .A(n9893), .B(n9894), .Z(n9913) );
  XOR U10036 ( .A(n9914), .B(n9913), .Z(c[125]) );
  NANDN U10037 ( .A(n9892), .B(n9891), .Z(n9896) );
  NANDN U10038 ( .A(n9894), .B(n9893), .Z(n9895) );
  NAND U10039 ( .A(n9896), .B(n9895), .Z(n9920) );
  IV U10040 ( .A(n9920), .Z(n9917) );
  NAND U10041 ( .A(n9898), .B(n9897), .Z(n9902) );
  NAND U10042 ( .A(n9900), .B(n9899), .Z(n9901) );
  AND U10043 ( .A(n9902), .B(n9901), .Z(n9921) );
  XOR U10044 ( .A(n9917), .B(n9921), .Z(n9916) );
  OR U10045 ( .A(n9903), .B(n580), .Z(n9906) );
  NANDN U10046 ( .A(n9904), .B(b[31]), .Z(n9905) );
  NAND U10047 ( .A(n9906), .B(n9905), .Z(n9925) );
  NAND U10048 ( .A(b[31]), .B(a[62]), .Z(n9924) );
  XOR U10049 ( .A(n9925), .B(n9924), .Z(n9923) );
  AND U10050 ( .A(n9908), .B(n9907), .Z(n9912) );
  NAND U10051 ( .A(n9910), .B(n9909), .Z(n9911) );
  NANDN U10052 ( .A(n9912), .B(n9911), .Z(n9922) );
  XNOR U10053 ( .A(n9923), .B(n9922), .Z(n9918) );
  AND U10054 ( .A(n9914), .B(n9913), .Z(n9919) );
  XNOR U10055 ( .A(n9918), .B(n9919), .Z(n9915) );
  XNOR U10056 ( .A(n9916), .B(n9915), .Z(c[126]) );
endmodule

