
module mult_N128_CC128 ( clk, rst, g_input, e_input, o );
  input [127:0] g_input;
  input [0:0] e_input;
  output [255:0] o;
  input clk, rst;
  wire   \add_42/carry[255] , \add_42/carry[254] , \add_42/carry[253] ,
         \add_42/carry[252] , \add_42/carry[251] , \add_42/carry[250] ,
         \add_42/carry[249] , \add_42/carry[248] , \add_42/carry[247] ,
         \add_42/carry[246] , \add_42/carry[245] , \add_42/carry[244] ,
         \add_42/carry[243] , \add_42/carry[242] , \add_42/carry[241] ,
         \add_42/carry[240] , \add_42/carry[239] , \add_42/carry[238] ,
         \add_42/carry[237] , \add_42/carry[236] , \add_42/carry[235] ,
         \add_42/carry[234] , \add_42/carry[233] , \add_42/carry[232] ,
         \add_42/carry[231] , \add_42/carry[230] , \add_42/carry[229] ,
         \add_42/carry[228] , \add_42/carry[227] , \add_42/carry[226] ,
         \add_42/carry[225] , \add_42/carry[224] , \add_42/carry[223] ,
         \add_42/carry[222] , \add_42/carry[221] , \add_42/carry[220] ,
         \add_42/carry[219] , \add_42/carry[218] , \add_42/carry[217] ,
         \add_42/carry[216] , \add_42/carry[215] , \add_42/carry[214] ,
         \add_42/carry[213] , \add_42/carry[212] , \add_42/carry[211] ,
         \add_42/carry[210] , \add_42/carry[209] , \add_42/carry[208] ,
         \add_42/carry[207] , \add_42/carry[206] , \add_42/carry[205] ,
         \add_42/carry[204] , \add_42/carry[203] , \add_42/carry[202] ,
         \add_42/carry[201] , \add_42/carry[200] , \add_42/carry[199] ,
         \add_42/carry[198] , \add_42/carry[197] , \add_42/carry[196] ,
         \add_42/carry[195] , \add_42/carry[194] , \add_42/carry[193] ,
         \add_42/carry[192] , \add_42/carry[191] , \add_42/carry[190] ,
         \add_42/carry[189] , \add_42/carry[188] , \add_42/carry[187] ,
         \add_42/carry[186] , \add_42/carry[185] , \add_42/carry[184] ,
         \add_42/carry[183] , \add_42/carry[182] , \add_42/carry[181] ,
         \add_42/carry[180] , \add_42/carry[179] , \add_42/carry[178] ,
         \add_42/carry[177] , \add_42/carry[176] , \add_42/carry[175] ,
         \add_42/carry[174] , \add_42/carry[173] , \add_42/carry[172] ,
         \add_42/carry[171] , \add_42/carry[170] , \add_42/carry[169] ,
         \add_42/carry[168] , \add_42/carry[167] , \add_42/carry[166] ,
         \add_42/carry[165] , \add_42/carry[164] , \add_42/carry[163] ,
         \add_42/carry[162] , \add_42/carry[161] , \add_42/carry[160] ,
         \add_42/carry[159] , \add_42/carry[158] , \add_42/carry[157] ,
         \add_42/carry[156] , \add_42/carry[155] , \add_42/carry[154] ,
         \add_42/carry[153] , \add_42/carry[152] , \add_42/carry[151] ,
         \add_42/carry[150] , \add_42/carry[149] , \add_42/carry[148] ,
         \add_42/carry[147] , \add_42/carry[146] , \add_42/carry[145] ,
         \add_42/carry[144] , \add_42/carry[143] , \add_42/carry[142] ,
         \add_42/carry[141] , \add_42/carry[140] , \add_42/carry[139] ,
         \add_42/carry[138] , \add_42/carry[137] , \add_42/carry[136] ,
         \add_42/carry[135] , \add_42/carry[134] , \add_42/carry[133] ,
         \add_42/carry[132] , \add_42/carry[131] , \add_42/carry[130] ,
         \add_42/carry[129] , \add_42/carry[128] , n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385;
  wire   [255:0] sreg;
  assign o[126] = sreg[126];
  assign o[125] = sreg[125];
  assign o[124] = sreg[124];
  assign o[123] = sreg[123];
  assign o[122] = sreg[122];
  assign o[121] = sreg[121];
  assign o[120] = sreg[120];
  assign o[119] = sreg[119];
  assign o[118] = sreg[118];
  assign o[117] = sreg[117];
  assign o[116] = sreg[116];
  assign o[115] = sreg[115];
  assign o[114] = sreg[114];
  assign o[113] = sreg[113];
  assign o[112] = sreg[112];
  assign o[111] = sreg[111];
  assign o[110] = sreg[110];
  assign o[109] = sreg[109];
  assign o[108] = sreg[108];
  assign o[107] = sreg[107];
  assign o[106] = sreg[106];
  assign o[105] = sreg[105];
  assign o[104] = sreg[104];
  assign o[103] = sreg[103];
  assign o[102] = sreg[102];
  assign o[101] = sreg[101];
  assign o[100] = sreg[100];
  assign o[99] = sreg[99];
  assign o[98] = sreg[98];
  assign o[97] = sreg[97];
  assign o[96] = sreg[96];
  assign o[95] = sreg[95];
  assign o[94] = sreg[94];
  assign o[93] = sreg[93];
  assign o[92] = sreg[92];
  assign o[91] = sreg[91];
  assign o[90] = sreg[90];
  assign o[89] = sreg[89];
  assign o[88] = sreg[88];
  assign o[87] = sreg[87];
  assign o[86] = sreg[86];
  assign o[85] = sreg[85];
  assign o[84] = sreg[84];
  assign o[83] = sreg[83];
  assign o[82] = sreg[82];
  assign o[81] = sreg[81];
  assign o[80] = sreg[80];
  assign o[79] = sreg[79];
  assign o[78] = sreg[78];
  assign o[77] = sreg[77];
  assign o[76] = sreg[76];
  assign o[75] = sreg[75];
  assign o[74] = sreg[74];
  assign o[73] = sreg[73];
  assign o[72] = sreg[72];
  assign o[71] = sreg[71];
  assign o[70] = sreg[70];
  assign o[69] = sreg[69];
  assign o[68] = sreg[68];
  assign o[67] = sreg[67];
  assign o[66] = sreg[66];
  assign o[65] = sreg[65];
  assign o[64] = sreg[64];
  assign o[63] = sreg[63];
  assign o[62] = sreg[62];
  assign o[61] = sreg[61];
  assign o[60] = sreg[60];
  assign o[59] = sreg[59];
  assign o[58] = sreg[58];
  assign o[57] = sreg[57];
  assign o[56] = sreg[56];
  assign o[55] = sreg[55];
  assign o[54] = sreg[54];
  assign o[53] = sreg[53];
  assign o[52] = sreg[52];
  assign o[51] = sreg[51];
  assign o[50] = sreg[50];
  assign o[49] = sreg[49];
  assign o[48] = sreg[48];
  assign o[47] = sreg[47];
  assign o[46] = sreg[46];
  assign o[45] = sreg[45];
  assign o[44] = sreg[44];
  assign o[43] = sreg[43];
  assign o[42] = sreg[42];
  assign o[41] = sreg[41];
  assign o[40] = sreg[40];
  assign o[39] = sreg[39];
  assign o[38] = sreg[38];
  assign o[37] = sreg[37];
  assign o[36] = sreg[36];
  assign o[35] = sreg[35];
  assign o[34] = sreg[34];
  assign o[33] = sreg[33];
  assign o[32] = sreg[32];
  assign o[31] = sreg[31];
  assign o[30] = sreg[30];
  assign o[29] = sreg[29];
  assign o[28] = sreg[28];
  assign o[27] = sreg[27];
  assign o[26] = sreg[26];
  assign o[25] = sreg[25];
  assign o[24] = sreg[24];
  assign o[23] = sreg[23];
  assign o[22] = sreg[22];
  assign o[21] = sreg[21];
  assign o[20] = sreg[20];
  assign o[19] = sreg[19];
  assign o[18] = sreg[18];
  assign o[17] = sreg[17];
  assign o[16] = sreg[16];
  assign o[15] = sreg[15];
  assign o[14] = sreg[14];
  assign o[13] = sreg[13];
  assign o[12] = sreg[12];
  assign o[11] = sreg[11];
  assign o[10] = sreg[10];
  assign o[9] = sreg[9];
  assign o[8] = sreg[8];
  assign o[7] = sreg[7];
  assign o[6] = sreg[6];
  assign o[5] = sreg[5];
  assign o[4] = sreg[4];
  assign o[3] = sreg[3];
  assign o[2] = sreg[2];
  assign o[1] = sreg[1];
  assign o[255] = \add_42/carry[255] ;

  DFF \sreg_reg[0]  ( .D(sreg[1]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[0]) );
  DFF \sreg_reg[1]  ( .D(sreg[2]), .CLK(clk), .RST(rst), .I(1'b0), .Q(sreg[1])
         );
  DFF \sreg_reg[2]  ( .D(sreg[3]), .CLK(clk), .RST(rst), .I(1'b0), .Q(sreg[2])
         );
  DFF \sreg_reg[3]  ( .D(sreg[4]), .CLK(clk), .RST(rst), .I(1'b0), .Q(sreg[3])
         );
  DFF \sreg_reg[4]  ( .D(sreg[5]), .CLK(clk), .RST(rst), .I(1'b0), .Q(sreg[4])
         );
  DFF \sreg_reg[5]  ( .D(sreg[6]), .CLK(clk), .RST(rst), .I(1'b0), .Q(sreg[5])
         );
  DFF \sreg_reg[6]  ( .D(sreg[7]), .CLK(clk), .RST(rst), .I(1'b0), .Q(sreg[6])
         );
  DFF \sreg_reg[7]  ( .D(sreg[8]), .CLK(clk), .RST(rst), .I(1'b0), .Q(sreg[7])
         );
  DFF \sreg_reg[8]  ( .D(sreg[9]), .CLK(clk), .RST(rst), .I(1'b0), .Q(sreg[8])
         );
  DFF \sreg_reg[9]  ( .D(sreg[10]), .CLK(clk), .RST(rst), .I(1'b0), .Q(sreg[9]) );
  DFF \sreg_reg[10]  ( .D(sreg[11]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[10]) );
  DFF \sreg_reg[11]  ( .D(sreg[12]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[11]) );
  DFF \sreg_reg[12]  ( .D(sreg[13]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[12]) );
  DFF \sreg_reg[13]  ( .D(sreg[14]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[13]) );
  DFF \sreg_reg[14]  ( .D(sreg[15]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[14]) );
  DFF \sreg_reg[15]  ( .D(sreg[16]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[15]) );
  DFF \sreg_reg[16]  ( .D(sreg[17]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[16]) );
  DFF \sreg_reg[17]  ( .D(sreg[18]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[17]) );
  DFF \sreg_reg[18]  ( .D(sreg[19]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[18]) );
  DFF \sreg_reg[19]  ( .D(sreg[20]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[19]) );
  DFF \sreg_reg[20]  ( .D(sreg[21]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[20]) );
  DFF \sreg_reg[21]  ( .D(sreg[22]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[21]) );
  DFF \sreg_reg[22]  ( .D(sreg[23]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[22]) );
  DFF \sreg_reg[23]  ( .D(sreg[24]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[23]) );
  DFF \sreg_reg[24]  ( .D(sreg[25]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[24]) );
  DFF \sreg_reg[25]  ( .D(sreg[26]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[25]) );
  DFF \sreg_reg[26]  ( .D(sreg[27]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[26]) );
  DFF \sreg_reg[27]  ( .D(sreg[28]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[27]) );
  DFF \sreg_reg[28]  ( .D(sreg[29]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[28]) );
  DFF \sreg_reg[29]  ( .D(sreg[30]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[29]) );
  DFF \sreg_reg[30]  ( .D(sreg[31]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[30]) );
  DFF \sreg_reg[31]  ( .D(sreg[32]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[31]) );
  DFF \sreg_reg[32]  ( .D(sreg[33]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[32]) );
  DFF \sreg_reg[33]  ( .D(sreg[34]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[33]) );
  DFF \sreg_reg[34]  ( .D(sreg[35]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[34]) );
  DFF \sreg_reg[35]  ( .D(sreg[36]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[35]) );
  DFF \sreg_reg[36]  ( .D(sreg[37]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[36]) );
  DFF \sreg_reg[37]  ( .D(sreg[38]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[37]) );
  DFF \sreg_reg[38]  ( .D(sreg[39]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[38]) );
  DFF \sreg_reg[39]  ( .D(sreg[40]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[39]) );
  DFF \sreg_reg[40]  ( .D(sreg[41]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[40]) );
  DFF \sreg_reg[41]  ( .D(sreg[42]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[41]) );
  DFF \sreg_reg[42]  ( .D(sreg[43]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[42]) );
  DFF \sreg_reg[43]  ( .D(sreg[44]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[43]) );
  DFF \sreg_reg[44]  ( .D(sreg[45]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[44]) );
  DFF \sreg_reg[45]  ( .D(sreg[46]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[45]) );
  DFF \sreg_reg[46]  ( .D(sreg[47]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[46]) );
  DFF \sreg_reg[47]  ( .D(sreg[48]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[47]) );
  DFF \sreg_reg[48]  ( .D(sreg[49]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[48]) );
  DFF \sreg_reg[49]  ( .D(sreg[50]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[49]) );
  DFF \sreg_reg[50]  ( .D(sreg[51]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[50]) );
  DFF \sreg_reg[51]  ( .D(sreg[52]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[51]) );
  DFF \sreg_reg[52]  ( .D(sreg[53]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[52]) );
  DFF \sreg_reg[53]  ( .D(sreg[54]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[53]) );
  DFF \sreg_reg[54]  ( .D(sreg[55]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[54]) );
  DFF \sreg_reg[55]  ( .D(sreg[56]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[55]) );
  DFF \sreg_reg[56]  ( .D(sreg[57]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[56]) );
  DFF \sreg_reg[57]  ( .D(sreg[58]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[57]) );
  DFF \sreg_reg[58]  ( .D(sreg[59]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[58]) );
  DFF \sreg_reg[59]  ( .D(sreg[60]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[59]) );
  DFF \sreg_reg[60]  ( .D(sreg[61]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[60]) );
  DFF \sreg_reg[61]  ( .D(sreg[62]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[61]) );
  DFF \sreg_reg[62]  ( .D(sreg[63]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[62]) );
  DFF \sreg_reg[63]  ( .D(sreg[64]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[63]) );
  DFF \sreg_reg[64]  ( .D(sreg[65]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[64]) );
  DFF \sreg_reg[65]  ( .D(sreg[66]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[65]) );
  DFF \sreg_reg[66]  ( .D(sreg[67]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[66]) );
  DFF \sreg_reg[67]  ( .D(sreg[68]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[67]) );
  DFF \sreg_reg[68]  ( .D(sreg[69]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[68]) );
  DFF \sreg_reg[69]  ( .D(sreg[70]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[69]) );
  DFF \sreg_reg[70]  ( .D(sreg[71]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[70]) );
  DFF \sreg_reg[71]  ( .D(sreg[72]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[71]) );
  DFF \sreg_reg[72]  ( .D(sreg[73]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[72]) );
  DFF \sreg_reg[73]  ( .D(sreg[74]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[73]) );
  DFF \sreg_reg[74]  ( .D(sreg[75]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[74]) );
  DFF \sreg_reg[75]  ( .D(sreg[76]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[75]) );
  DFF \sreg_reg[76]  ( .D(sreg[77]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[76]) );
  DFF \sreg_reg[77]  ( .D(sreg[78]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[77]) );
  DFF \sreg_reg[78]  ( .D(sreg[79]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[78]) );
  DFF \sreg_reg[79]  ( .D(sreg[80]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[79]) );
  DFF \sreg_reg[80]  ( .D(sreg[81]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[80]) );
  DFF \sreg_reg[81]  ( .D(sreg[82]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[81]) );
  DFF \sreg_reg[82]  ( .D(sreg[83]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[82]) );
  DFF \sreg_reg[83]  ( .D(sreg[84]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[83]) );
  DFF \sreg_reg[84]  ( .D(sreg[85]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[84]) );
  DFF \sreg_reg[85]  ( .D(sreg[86]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[85]) );
  DFF \sreg_reg[86]  ( .D(sreg[87]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[86]) );
  DFF \sreg_reg[87]  ( .D(sreg[88]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[87]) );
  DFF \sreg_reg[88]  ( .D(sreg[89]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[88]) );
  DFF \sreg_reg[89]  ( .D(sreg[90]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[89]) );
  DFF \sreg_reg[90]  ( .D(sreg[91]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[90]) );
  DFF \sreg_reg[91]  ( .D(sreg[92]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[91]) );
  DFF \sreg_reg[92]  ( .D(sreg[93]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[92]) );
  DFF \sreg_reg[93]  ( .D(sreg[94]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[93]) );
  DFF \sreg_reg[94]  ( .D(sreg[95]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[94]) );
  DFF \sreg_reg[95]  ( .D(sreg[96]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[95]) );
  DFF \sreg_reg[96]  ( .D(sreg[97]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[96]) );
  DFF \sreg_reg[97]  ( .D(sreg[98]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[97]) );
  DFF \sreg_reg[98]  ( .D(sreg[99]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[98]) );
  DFF \sreg_reg[99]  ( .D(sreg[100]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[99]) );
  DFF \sreg_reg[100]  ( .D(sreg[101]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[100]) );
  DFF \sreg_reg[101]  ( .D(sreg[102]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[101]) );
  DFF \sreg_reg[102]  ( .D(sreg[103]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[102]) );
  DFF \sreg_reg[103]  ( .D(sreg[104]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[103]) );
  DFF \sreg_reg[104]  ( .D(sreg[105]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[104]) );
  DFF \sreg_reg[105]  ( .D(sreg[106]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[105]) );
  DFF \sreg_reg[106]  ( .D(sreg[107]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[106]) );
  DFF \sreg_reg[107]  ( .D(sreg[108]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[107]) );
  DFF \sreg_reg[108]  ( .D(sreg[109]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[108]) );
  DFF \sreg_reg[109]  ( .D(sreg[110]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[109]) );
  DFF \sreg_reg[110]  ( .D(sreg[111]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[110]) );
  DFF \sreg_reg[111]  ( .D(sreg[112]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[111]) );
  DFF \sreg_reg[112]  ( .D(sreg[113]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[112]) );
  DFF \sreg_reg[113]  ( .D(sreg[114]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[113]) );
  DFF \sreg_reg[114]  ( .D(sreg[115]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[114]) );
  DFF \sreg_reg[115]  ( .D(sreg[116]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[115]) );
  DFF \sreg_reg[116]  ( .D(sreg[117]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[116]) );
  DFF \sreg_reg[117]  ( .D(sreg[118]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[117]) );
  DFF \sreg_reg[118]  ( .D(sreg[119]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[118]) );
  DFF \sreg_reg[119]  ( .D(sreg[120]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[119]) );
  DFF \sreg_reg[120]  ( .D(sreg[121]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[120]) );
  DFF \sreg_reg[121]  ( .D(sreg[122]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[121]) );
  DFF \sreg_reg[122]  ( .D(sreg[123]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[122]) );
  DFF \sreg_reg[123]  ( .D(sreg[124]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[123]) );
  DFF \sreg_reg[124]  ( .D(sreg[125]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[124]) );
  DFF \sreg_reg[125]  ( .D(sreg[126]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[125]) );
  DFF \sreg_reg[126]  ( .D(o[127]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[126]) );
  DFF \sreg_reg[127]  ( .D(o[128]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[127]) );
  DFF \sreg_reg[128]  ( .D(o[129]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[128]) );
  DFF \sreg_reg[129]  ( .D(o[130]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[129]) );
  DFF \sreg_reg[130]  ( .D(o[131]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[130]) );
  DFF \sreg_reg[131]  ( .D(o[132]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[131]) );
  DFF \sreg_reg[132]  ( .D(o[133]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[132]) );
  DFF \sreg_reg[133]  ( .D(o[134]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[133]) );
  DFF \sreg_reg[134]  ( .D(o[135]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[134]) );
  DFF \sreg_reg[135]  ( .D(o[136]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[135]) );
  DFF \sreg_reg[136]  ( .D(o[137]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[136]) );
  DFF \sreg_reg[137]  ( .D(o[138]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[137]) );
  DFF \sreg_reg[138]  ( .D(o[139]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[138]) );
  DFF \sreg_reg[139]  ( .D(o[140]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[139]) );
  DFF \sreg_reg[140]  ( .D(o[141]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[140]) );
  DFF \sreg_reg[141]  ( .D(o[142]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[141]) );
  DFF \sreg_reg[142]  ( .D(o[143]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[142]) );
  DFF \sreg_reg[143]  ( .D(o[144]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[143]) );
  DFF \sreg_reg[144]  ( .D(o[145]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[144]) );
  DFF \sreg_reg[145]  ( .D(o[146]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[145]) );
  DFF \sreg_reg[146]  ( .D(o[147]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[146]) );
  DFF \sreg_reg[147]  ( .D(o[148]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[147]) );
  DFF \sreg_reg[148]  ( .D(o[149]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[148]) );
  DFF \sreg_reg[149]  ( .D(o[150]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[149]) );
  DFF \sreg_reg[150]  ( .D(o[151]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[150]) );
  DFF \sreg_reg[151]  ( .D(o[152]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[151]) );
  DFF \sreg_reg[152]  ( .D(o[153]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[152]) );
  DFF \sreg_reg[153]  ( .D(o[154]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[153]) );
  DFF \sreg_reg[154]  ( .D(o[155]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[154]) );
  DFF \sreg_reg[155]  ( .D(o[156]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[155]) );
  DFF \sreg_reg[156]  ( .D(o[157]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[156]) );
  DFF \sreg_reg[157]  ( .D(o[158]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[157]) );
  DFF \sreg_reg[158]  ( .D(o[159]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[158]) );
  DFF \sreg_reg[159]  ( .D(o[160]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[159]) );
  DFF \sreg_reg[160]  ( .D(o[161]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[160]) );
  DFF \sreg_reg[161]  ( .D(o[162]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[161]) );
  DFF \sreg_reg[162]  ( .D(o[163]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[162]) );
  DFF \sreg_reg[163]  ( .D(o[164]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[163]) );
  DFF \sreg_reg[164]  ( .D(o[165]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[164]) );
  DFF \sreg_reg[165]  ( .D(o[166]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[165]) );
  DFF \sreg_reg[166]  ( .D(o[167]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[166]) );
  DFF \sreg_reg[167]  ( .D(o[168]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[167]) );
  DFF \sreg_reg[168]  ( .D(o[169]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[168]) );
  DFF \sreg_reg[169]  ( .D(o[170]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[169]) );
  DFF \sreg_reg[170]  ( .D(o[171]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[170]) );
  DFF \sreg_reg[171]  ( .D(o[172]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[171]) );
  DFF \sreg_reg[172]  ( .D(o[173]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[172]) );
  DFF \sreg_reg[173]  ( .D(o[174]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[173]) );
  DFF \sreg_reg[174]  ( .D(o[175]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[174]) );
  DFF \sreg_reg[175]  ( .D(o[176]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[175]) );
  DFF \sreg_reg[176]  ( .D(o[177]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[176]) );
  DFF \sreg_reg[177]  ( .D(o[178]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[177]) );
  DFF \sreg_reg[178]  ( .D(o[179]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[178]) );
  DFF \sreg_reg[179]  ( .D(o[180]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[179]) );
  DFF \sreg_reg[180]  ( .D(o[181]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[180]) );
  DFF \sreg_reg[181]  ( .D(o[182]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[181]) );
  DFF \sreg_reg[182]  ( .D(o[183]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[182]) );
  DFF \sreg_reg[183]  ( .D(o[184]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[183]) );
  DFF \sreg_reg[184]  ( .D(o[185]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[184]) );
  DFF \sreg_reg[185]  ( .D(o[186]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[185]) );
  DFF \sreg_reg[186]  ( .D(o[187]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[186]) );
  DFF \sreg_reg[187]  ( .D(o[188]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[187]) );
  DFF \sreg_reg[188]  ( .D(o[189]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[188]) );
  DFF \sreg_reg[189]  ( .D(o[190]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[189]) );
  DFF \sreg_reg[190]  ( .D(o[191]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[190]) );
  DFF \sreg_reg[191]  ( .D(o[192]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[191]) );
  DFF \sreg_reg[192]  ( .D(o[193]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[192]) );
  DFF \sreg_reg[193]  ( .D(o[194]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[193]) );
  DFF \sreg_reg[194]  ( .D(o[195]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[194]) );
  DFF \sreg_reg[195]  ( .D(o[196]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[195]) );
  DFF \sreg_reg[196]  ( .D(o[197]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[196]) );
  DFF \sreg_reg[197]  ( .D(o[198]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[197]) );
  DFF \sreg_reg[198]  ( .D(o[199]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[198]) );
  DFF \sreg_reg[199]  ( .D(o[200]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[199]) );
  DFF \sreg_reg[200]  ( .D(o[201]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[200]) );
  DFF \sreg_reg[201]  ( .D(o[202]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[201]) );
  DFF \sreg_reg[202]  ( .D(o[203]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[202]) );
  DFF \sreg_reg[203]  ( .D(o[204]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[203]) );
  DFF \sreg_reg[204]  ( .D(o[205]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[204]) );
  DFF \sreg_reg[205]  ( .D(o[206]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[205]) );
  DFF \sreg_reg[206]  ( .D(o[207]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[206]) );
  DFF \sreg_reg[207]  ( .D(o[208]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[207]) );
  DFF \sreg_reg[208]  ( .D(o[209]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[208]) );
  DFF \sreg_reg[209]  ( .D(o[210]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[209]) );
  DFF \sreg_reg[210]  ( .D(o[211]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[210]) );
  DFF \sreg_reg[211]  ( .D(o[212]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[211]) );
  DFF \sreg_reg[212]  ( .D(o[213]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[212]) );
  DFF \sreg_reg[213]  ( .D(o[214]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[213]) );
  DFF \sreg_reg[214]  ( .D(o[215]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[214]) );
  DFF \sreg_reg[215]  ( .D(o[216]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[215]) );
  DFF \sreg_reg[216]  ( .D(o[217]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[216]) );
  DFF \sreg_reg[217]  ( .D(o[218]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[217]) );
  DFF \sreg_reg[218]  ( .D(o[219]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[218]) );
  DFF \sreg_reg[219]  ( .D(o[220]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[219]) );
  DFF \sreg_reg[220]  ( .D(o[221]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[220]) );
  DFF \sreg_reg[221]  ( .D(o[222]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[221]) );
  DFF \sreg_reg[222]  ( .D(o[223]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[222]) );
  DFF \sreg_reg[223]  ( .D(o[224]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[223]) );
  DFF \sreg_reg[224]  ( .D(o[225]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[224]) );
  DFF \sreg_reg[225]  ( .D(o[226]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[225]) );
  DFF \sreg_reg[226]  ( .D(o[227]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[226]) );
  DFF \sreg_reg[227]  ( .D(o[228]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[227]) );
  DFF \sreg_reg[228]  ( .D(o[229]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[228]) );
  DFF \sreg_reg[229]  ( .D(o[230]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[229]) );
  DFF \sreg_reg[230]  ( .D(o[231]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[230]) );
  DFF \sreg_reg[231]  ( .D(o[232]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[231]) );
  DFF \sreg_reg[232]  ( .D(o[233]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[232]) );
  DFF \sreg_reg[233]  ( .D(o[234]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[233]) );
  DFF \sreg_reg[234]  ( .D(o[235]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[234]) );
  DFF \sreg_reg[235]  ( .D(o[236]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[235]) );
  DFF \sreg_reg[236]  ( .D(o[237]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[236]) );
  DFF \sreg_reg[237]  ( .D(o[238]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[237]) );
  DFF \sreg_reg[238]  ( .D(o[239]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[238]) );
  DFF \sreg_reg[239]  ( .D(o[240]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[239]) );
  DFF \sreg_reg[240]  ( .D(o[241]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[240]) );
  DFF \sreg_reg[241]  ( .D(o[242]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[241]) );
  DFF \sreg_reg[242]  ( .D(o[243]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[242]) );
  DFF \sreg_reg[243]  ( .D(o[244]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[243]) );
  DFF \sreg_reg[244]  ( .D(o[245]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[244]) );
  DFF \sreg_reg[245]  ( .D(o[246]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[245]) );
  DFF \sreg_reg[246]  ( .D(o[247]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[246]) );
  DFF \sreg_reg[247]  ( .D(o[248]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[247]) );
  DFF \sreg_reg[248]  ( .D(o[249]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[248]) );
  DFF \sreg_reg[249]  ( .D(o[250]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[249]) );
  DFF \sreg_reg[250]  ( .D(o[251]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[250]) );
  DFF \sreg_reg[251]  ( .D(o[252]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[251]) );
  DFF \sreg_reg[252]  ( .D(o[253]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[252]) );
  DFF \sreg_reg[253]  ( .D(o[254]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[253]) );
  DFF \sreg_reg[254]  ( .D(\add_42/carry[255] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(sreg[254]) );
  FADDER \add_42/U1_128  ( .CIN(sreg[128]), .IN0(n384), .IN1(
        \add_42/carry[128] ), .COUT(\add_42/carry[129] ), .SUM(o[128]) );
  FADDER \add_42/U1_129  ( .CIN(sreg[129]), .IN0(n383), .IN1(
        \add_42/carry[129] ), .COUT(\add_42/carry[130] ), .SUM(o[129]) );
  FADDER \add_42/U1_130  ( .CIN(sreg[130]), .IN0(n382), .IN1(
        \add_42/carry[130] ), .COUT(\add_42/carry[131] ), .SUM(o[130]) );
  FADDER \add_42/U1_131  ( .CIN(sreg[131]), .IN0(n381), .IN1(
        \add_42/carry[131] ), .COUT(\add_42/carry[132] ), .SUM(o[131]) );
  FADDER \add_42/U1_132  ( .CIN(sreg[132]), .IN0(n380), .IN1(
        \add_42/carry[132] ), .COUT(\add_42/carry[133] ), .SUM(o[132]) );
  FADDER \add_42/U1_133  ( .CIN(sreg[133]), .IN0(n379), .IN1(
        \add_42/carry[133] ), .COUT(\add_42/carry[134] ), .SUM(o[133]) );
  FADDER \add_42/U1_134  ( .CIN(sreg[134]), .IN0(n378), .IN1(
        \add_42/carry[134] ), .COUT(\add_42/carry[135] ), .SUM(o[134]) );
  FADDER \add_42/U1_135  ( .CIN(sreg[135]), .IN0(n377), .IN1(
        \add_42/carry[135] ), .COUT(\add_42/carry[136] ), .SUM(o[135]) );
  FADDER \add_42/U1_136  ( .CIN(sreg[136]), .IN0(n376), .IN1(
        \add_42/carry[136] ), .COUT(\add_42/carry[137] ), .SUM(o[136]) );
  FADDER \add_42/U1_137  ( .CIN(sreg[137]), .IN0(n375), .IN1(
        \add_42/carry[137] ), .COUT(\add_42/carry[138] ), .SUM(o[137]) );
  FADDER \add_42/U1_138  ( .CIN(sreg[138]), .IN0(n374), .IN1(
        \add_42/carry[138] ), .COUT(\add_42/carry[139] ), .SUM(o[138]) );
  FADDER \add_42/U1_139  ( .CIN(sreg[139]), .IN0(n373), .IN1(
        \add_42/carry[139] ), .COUT(\add_42/carry[140] ), .SUM(o[139]) );
  FADDER \add_42/U1_140  ( .CIN(sreg[140]), .IN0(n372), .IN1(
        \add_42/carry[140] ), .COUT(\add_42/carry[141] ), .SUM(o[140]) );
  FADDER \add_42/U1_141  ( .CIN(sreg[141]), .IN0(n371), .IN1(
        \add_42/carry[141] ), .COUT(\add_42/carry[142] ), .SUM(o[141]) );
  FADDER \add_42/U1_142  ( .CIN(sreg[142]), .IN0(n370), .IN1(
        \add_42/carry[142] ), .COUT(\add_42/carry[143] ), .SUM(o[142]) );
  FADDER \add_42/U1_143  ( .CIN(sreg[143]), .IN0(n369), .IN1(
        \add_42/carry[143] ), .COUT(\add_42/carry[144] ), .SUM(o[143]) );
  FADDER \add_42/U1_144  ( .CIN(sreg[144]), .IN0(n368), .IN1(
        \add_42/carry[144] ), .COUT(\add_42/carry[145] ), .SUM(o[144]) );
  FADDER \add_42/U1_145  ( .CIN(sreg[145]), .IN0(n367), .IN1(
        \add_42/carry[145] ), .COUT(\add_42/carry[146] ), .SUM(o[145]) );
  FADDER \add_42/U1_146  ( .CIN(sreg[146]), .IN0(n366), .IN1(
        \add_42/carry[146] ), .COUT(\add_42/carry[147] ), .SUM(o[146]) );
  FADDER \add_42/U1_147  ( .CIN(sreg[147]), .IN0(n365), .IN1(
        \add_42/carry[147] ), .COUT(\add_42/carry[148] ), .SUM(o[147]) );
  FADDER \add_42/U1_148  ( .CIN(sreg[148]), .IN0(n364), .IN1(
        \add_42/carry[148] ), .COUT(\add_42/carry[149] ), .SUM(o[148]) );
  FADDER \add_42/U1_149  ( .CIN(sreg[149]), .IN0(n363), .IN1(
        \add_42/carry[149] ), .COUT(\add_42/carry[150] ), .SUM(o[149]) );
  FADDER \add_42/U1_150  ( .CIN(sreg[150]), .IN0(n362), .IN1(
        \add_42/carry[150] ), .COUT(\add_42/carry[151] ), .SUM(o[150]) );
  FADDER \add_42/U1_151  ( .CIN(sreg[151]), .IN0(n361), .IN1(
        \add_42/carry[151] ), .COUT(\add_42/carry[152] ), .SUM(o[151]) );
  FADDER \add_42/U1_152  ( .CIN(sreg[152]), .IN0(n360), .IN1(
        \add_42/carry[152] ), .COUT(\add_42/carry[153] ), .SUM(o[152]) );
  FADDER \add_42/U1_153  ( .CIN(sreg[153]), .IN0(n359), .IN1(
        \add_42/carry[153] ), .COUT(\add_42/carry[154] ), .SUM(o[153]) );
  FADDER \add_42/U1_154  ( .CIN(sreg[154]), .IN0(n358), .IN1(
        \add_42/carry[154] ), .COUT(\add_42/carry[155] ), .SUM(o[154]) );
  FADDER \add_42/U1_155  ( .CIN(sreg[155]), .IN0(n357), .IN1(
        \add_42/carry[155] ), .COUT(\add_42/carry[156] ), .SUM(o[155]) );
  FADDER \add_42/U1_156  ( .CIN(sreg[156]), .IN0(n356), .IN1(
        \add_42/carry[156] ), .COUT(\add_42/carry[157] ), .SUM(o[156]) );
  FADDER \add_42/U1_157  ( .CIN(sreg[157]), .IN0(n355), .IN1(
        \add_42/carry[157] ), .COUT(\add_42/carry[158] ), .SUM(o[157]) );
  FADDER \add_42/U1_158  ( .CIN(sreg[158]), .IN0(n354), .IN1(
        \add_42/carry[158] ), .COUT(\add_42/carry[159] ), .SUM(o[158]) );
  FADDER \add_42/U1_159  ( .CIN(sreg[159]), .IN0(n353), .IN1(
        \add_42/carry[159] ), .COUT(\add_42/carry[160] ), .SUM(o[159]) );
  FADDER \add_42/U1_160  ( .CIN(sreg[160]), .IN0(n352), .IN1(
        \add_42/carry[160] ), .COUT(\add_42/carry[161] ), .SUM(o[160]) );
  FADDER \add_42/U1_161  ( .CIN(sreg[161]), .IN0(n351), .IN1(
        \add_42/carry[161] ), .COUT(\add_42/carry[162] ), .SUM(o[161]) );
  FADDER \add_42/U1_162  ( .CIN(sreg[162]), .IN0(n350), .IN1(
        \add_42/carry[162] ), .COUT(\add_42/carry[163] ), .SUM(o[162]) );
  FADDER \add_42/U1_163  ( .CIN(sreg[163]), .IN0(n349), .IN1(
        \add_42/carry[163] ), .COUT(\add_42/carry[164] ), .SUM(o[163]) );
  FADDER \add_42/U1_164  ( .CIN(sreg[164]), .IN0(n348), .IN1(
        \add_42/carry[164] ), .COUT(\add_42/carry[165] ), .SUM(o[164]) );
  FADDER \add_42/U1_165  ( .CIN(sreg[165]), .IN0(n347), .IN1(
        \add_42/carry[165] ), .COUT(\add_42/carry[166] ), .SUM(o[165]) );
  FADDER \add_42/U1_166  ( .CIN(sreg[166]), .IN0(n346), .IN1(
        \add_42/carry[166] ), .COUT(\add_42/carry[167] ), .SUM(o[166]) );
  FADDER \add_42/U1_167  ( .CIN(sreg[167]), .IN0(n345), .IN1(
        \add_42/carry[167] ), .COUT(\add_42/carry[168] ), .SUM(o[167]) );
  FADDER \add_42/U1_168  ( .CIN(sreg[168]), .IN0(n344), .IN1(
        \add_42/carry[168] ), .COUT(\add_42/carry[169] ), .SUM(o[168]) );
  FADDER \add_42/U1_169  ( .CIN(sreg[169]), .IN0(n343), .IN1(
        \add_42/carry[169] ), .COUT(\add_42/carry[170] ), .SUM(o[169]) );
  FADDER \add_42/U1_170  ( .CIN(sreg[170]), .IN0(n342), .IN1(
        \add_42/carry[170] ), .COUT(\add_42/carry[171] ), .SUM(o[170]) );
  FADDER \add_42/U1_171  ( .CIN(sreg[171]), .IN0(n341), .IN1(
        \add_42/carry[171] ), .COUT(\add_42/carry[172] ), .SUM(o[171]) );
  FADDER \add_42/U1_172  ( .CIN(sreg[172]), .IN0(n340), .IN1(
        \add_42/carry[172] ), .COUT(\add_42/carry[173] ), .SUM(o[172]) );
  FADDER \add_42/U1_173  ( .CIN(sreg[173]), .IN0(n339), .IN1(
        \add_42/carry[173] ), .COUT(\add_42/carry[174] ), .SUM(o[173]) );
  FADDER \add_42/U1_174  ( .CIN(sreg[174]), .IN0(n338), .IN1(
        \add_42/carry[174] ), .COUT(\add_42/carry[175] ), .SUM(o[174]) );
  FADDER \add_42/U1_175  ( .CIN(sreg[175]), .IN0(n337), .IN1(
        \add_42/carry[175] ), .COUT(\add_42/carry[176] ), .SUM(o[175]) );
  FADDER \add_42/U1_176  ( .CIN(sreg[176]), .IN0(n336), .IN1(
        \add_42/carry[176] ), .COUT(\add_42/carry[177] ), .SUM(o[176]) );
  FADDER \add_42/U1_177  ( .CIN(sreg[177]), .IN0(n335), .IN1(
        \add_42/carry[177] ), .COUT(\add_42/carry[178] ), .SUM(o[177]) );
  FADDER \add_42/U1_178  ( .CIN(sreg[178]), .IN0(n334), .IN1(
        \add_42/carry[178] ), .COUT(\add_42/carry[179] ), .SUM(o[178]) );
  FADDER \add_42/U1_179  ( .CIN(sreg[179]), .IN0(n333), .IN1(
        \add_42/carry[179] ), .COUT(\add_42/carry[180] ), .SUM(o[179]) );
  FADDER \add_42/U1_180  ( .CIN(sreg[180]), .IN0(n332), .IN1(
        \add_42/carry[180] ), .COUT(\add_42/carry[181] ), .SUM(o[180]) );
  FADDER \add_42/U1_181  ( .CIN(sreg[181]), .IN0(n331), .IN1(
        \add_42/carry[181] ), .COUT(\add_42/carry[182] ), .SUM(o[181]) );
  FADDER \add_42/U1_182  ( .CIN(sreg[182]), .IN0(n330), .IN1(
        \add_42/carry[182] ), .COUT(\add_42/carry[183] ), .SUM(o[182]) );
  FADDER \add_42/U1_183  ( .CIN(sreg[183]), .IN0(n329), .IN1(
        \add_42/carry[183] ), .COUT(\add_42/carry[184] ), .SUM(o[183]) );
  FADDER \add_42/U1_184  ( .CIN(sreg[184]), .IN0(n328), .IN1(
        \add_42/carry[184] ), .COUT(\add_42/carry[185] ), .SUM(o[184]) );
  FADDER \add_42/U1_185  ( .CIN(sreg[185]), .IN0(n327), .IN1(
        \add_42/carry[185] ), .COUT(\add_42/carry[186] ), .SUM(o[185]) );
  FADDER \add_42/U1_186  ( .CIN(sreg[186]), .IN0(n326), .IN1(
        \add_42/carry[186] ), .COUT(\add_42/carry[187] ), .SUM(o[186]) );
  FADDER \add_42/U1_187  ( .CIN(sreg[187]), .IN0(n325), .IN1(
        \add_42/carry[187] ), .COUT(\add_42/carry[188] ), .SUM(o[187]) );
  FADDER \add_42/U1_188  ( .CIN(sreg[188]), .IN0(n324), .IN1(
        \add_42/carry[188] ), .COUT(\add_42/carry[189] ), .SUM(o[188]) );
  FADDER \add_42/U1_189  ( .CIN(sreg[189]), .IN0(n323), .IN1(
        \add_42/carry[189] ), .COUT(\add_42/carry[190] ), .SUM(o[189]) );
  FADDER \add_42/U1_190  ( .CIN(sreg[190]), .IN0(n322), .IN1(
        \add_42/carry[190] ), .COUT(\add_42/carry[191] ), .SUM(o[190]) );
  FADDER \add_42/U1_191  ( .CIN(sreg[191]), .IN0(n321), .IN1(
        \add_42/carry[191] ), .COUT(\add_42/carry[192] ), .SUM(o[191]) );
  FADDER \add_42/U1_192  ( .CIN(sreg[192]), .IN0(n320), .IN1(
        \add_42/carry[192] ), .COUT(\add_42/carry[193] ), .SUM(o[192]) );
  FADDER \add_42/U1_193  ( .CIN(sreg[193]), .IN0(n319), .IN1(
        \add_42/carry[193] ), .COUT(\add_42/carry[194] ), .SUM(o[193]) );
  FADDER \add_42/U1_194  ( .CIN(sreg[194]), .IN0(n318), .IN1(
        \add_42/carry[194] ), .COUT(\add_42/carry[195] ), .SUM(o[194]) );
  FADDER \add_42/U1_195  ( .CIN(sreg[195]), .IN0(n317), .IN1(
        \add_42/carry[195] ), .COUT(\add_42/carry[196] ), .SUM(o[195]) );
  FADDER \add_42/U1_196  ( .CIN(sreg[196]), .IN0(n316), .IN1(
        \add_42/carry[196] ), .COUT(\add_42/carry[197] ), .SUM(o[196]) );
  FADDER \add_42/U1_197  ( .CIN(sreg[197]), .IN0(n315), .IN1(
        \add_42/carry[197] ), .COUT(\add_42/carry[198] ), .SUM(o[197]) );
  FADDER \add_42/U1_198  ( .CIN(sreg[198]), .IN0(n314), .IN1(
        \add_42/carry[198] ), .COUT(\add_42/carry[199] ), .SUM(o[198]) );
  FADDER \add_42/U1_199  ( .CIN(sreg[199]), .IN0(n313), .IN1(
        \add_42/carry[199] ), .COUT(\add_42/carry[200] ), .SUM(o[199]) );
  FADDER \add_42/U1_200  ( .CIN(sreg[200]), .IN0(n312), .IN1(
        \add_42/carry[200] ), .COUT(\add_42/carry[201] ), .SUM(o[200]) );
  FADDER \add_42/U1_201  ( .CIN(sreg[201]), .IN0(n311), .IN1(
        \add_42/carry[201] ), .COUT(\add_42/carry[202] ), .SUM(o[201]) );
  FADDER \add_42/U1_202  ( .CIN(sreg[202]), .IN0(n310), .IN1(
        \add_42/carry[202] ), .COUT(\add_42/carry[203] ), .SUM(o[202]) );
  FADDER \add_42/U1_203  ( .CIN(sreg[203]), .IN0(n309), .IN1(
        \add_42/carry[203] ), .COUT(\add_42/carry[204] ), .SUM(o[203]) );
  FADDER \add_42/U1_204  ( .CIN(sreg[204]), .IN0(n308), .IN1(
        \add_42/carry[204] ), .COUT(\add_42/carry[205] ), .SUM(o[204]) );
  FADDER \add_42/U1_205  ( .CIN(sreg[205]), .IN0(n307), .IN1(
        \add_42/carry[205] ), .COUT(\add_42/carry[206] ), .SUM(o[205]) );
  FADDER \add_42/U1_206  ( .CIN(sreg[206]), .IN0(n306), .IN1(
        \add_42/carry[206] ), .COUT(\add_42/carry[207] ), .SUM(o[206]) );
  FADDER \add_42/U1_207  ( .CIN(sreg[207]), .IN0(n305), .IN1(
        \add_42/carry[207] ), .COUT(\add_42/carry[208] ), .SUM(o[207]) );
  FADDER \add_42/U1_208  ( .CIN(sreg[208]), .IN0(n304), .IN1(
        \add_42/carry[208] ), .COUT(\add_42/carry[209] ), .SUM(o[208]) );
  FADDER \add_42/U1_209  ( .CIN(sreg[209]), .IN0(n303), .IN1(
        \add_42/carry[209] ), .COUT(\add_42/carry[210] ), .SUM(o[209]) );
  FADDER \add_42/U1_210  ( .CIN(sreg[210]), .IN0(n302), .IN1(
        \add_42/carry[210] ), .COUT(\add_42/carry[211] ), .SUM(o[210]) );
  FADDER \add_42/U1_211  ( .CIN(sreg[211]), .IN0(n301), .IN1(
        \add_42/carry[211] ), .COUT(\add_42/carry[212] ), .SUM(o[211]) );
  FADDER \add_42/U1_212  ( .CIN(sreg[212]), .IN0(n300), .IN1(
        \add_42/carry[212] ), .COUT(\add_42/carry[213] ), .SUM(o[212]) );
  FADDER \add_42/U1_213  ( .CIN(sreg[213]), .IN0(n299), .IN1(
        \add_42/carry[213] ), .COUT(\add_42/carry[214] ), .SUM(o[213]) );
  FADDER \add_42/U1_214  ( .CIN(sreg[214]), .IN0(n298), .IN1(
        \add_42/carry[214] ), .COUT(\add_42/carry[215] ), .SUM(o[214]) );
  FADDER \add_42/U1_215  ( .CIN(sreg[215]), .IN0(n297), .IN1(
        \add_42/carry[215] ), .COUT(\add_42/carry[216] ), .SUM(o[215]) );
  FADDER \add_42/U1_216  ( .CIN(sreg[216]), .IN0(n296), .IN1(
        \add_42/carry[216] ), .COUT(\add_42/carry[217] ), .SUM(o[216]) );
  FADDER \add_42/U1_217  ( .CIN(sreg[217]), .IN0(n295), .IN1(
        \add_42/carry[217] ), .COUT(\add_42/carry[218] ), .SUM(o[217]) );
  FADDER \add_42/U1_218  ( .CIN(sreg[218]), .IN0(n294), .IN1(
        \add_42/carry[218] ), .COUT(\add_42/carry[219] ), .SUM(o[218]) );
  FADDER \add_42/U1_219  ( .CIN(sreg[219]), .IN0(n293), .IN1(
        \add_42/carry[219] ), .COUT(\add_42/carry[220] ), .SUM(o[219]) );
  FADDER \add_42/U1_220  ( .CIN(sreg[220]), .IN0(n292), .IN1(
        \add_42/carry[220] ), .COUT(\add_42/carry[221] ), .SUM(o[220]) );
  FADDER \add_42/U1_221  ( .CIN(sreg[221]), .IN0(n291), .IN1(
        \add_42/carry[221] ), .COUT(\add_42/carry[222] ), .SUM(o[221]) );
  FADDER \add_42/U1_222  ( .CIN(sreg[222]), .IN0(n290), .IN1(
        \add_42/carry[222] ), .COUT(\add_42/carry[223] ), .SUM(o[222]) );
  FADDER \add_42/U1_223  ( .CIN(sreg[223]), .IN0(n289), .IN1(
        \add_42/carry[223] ), .COUT(\add_42/carry[224] ), .SUM(o[223]) );
  FADDER \add_42/U1_224  ( .CIN(sreg[224]), .IN0(n288), .IN1(
        \add_42/carry[224] ), .COUT(\add_42/carry[225] ), .SUM(o[224]) );
  FADDER \add_42/U1_225  ( .CIN(sreg[225]), .IN0(n287), .IN1(
        \add_42/carry[225] ), .COUT(\add_42/carry[226] ), .SUM(o[225]) );
  FADDER \add_42/U1_226  ( .CIN(sreg[226]), .IN0(n286), .IN1(
        \add_42/carry[226] ), .COUT(\add_42/carry[227] ), .SUM(o[226]) );
  FADDER \add_42/U1_227  ( .CIN(sreg[227]), .IN0(n285), .IN1(
        \add_42/carry[227] ), .COUT(\add_42/carry[228] ), .SUM(o[227]) );
  FADDER \add_42/U1_228  ( .CIN(sreg[228]), .IN0(n284), .IN1(
        \add_42/carry[228] ), .COUT(\add_42/carry[229] ), .SUM(o[228]) );
  FADDER \add_42/U1_229  ( .CIN(sreg[229]), .IN0(n283), .IN1(
        \add_42/carry[229] ), .COUT(\add_42/carry[230] ), .SUM(o[229]) );
  FADDER \add_42/U1_230  ( .CIN(sreg[230]), .IN0(n282), .IN1(
        \add_42/carry[230] ), .COUT(\add_42/carry[231] ), .SUM(o[230]) );
  FADDER \add_42/U1_231  ( .CIN(sreg[231]), .IN0(n281), .IN1(
        \add_42/carry[231] ), .COUT(\add_42/carry[232] ), .SUM(o[231]) );
  FADDER \add_42/U1_232  ( .CIN(sreg[232]), .IN0(n280), .IN1(
        \add_42/carry[232] ), .COUT(\add_42/carry[233] ), .SUM(o[232]) );
  FADDER \add_42/U1_233  ( .CIN(sreg[233]), .IN0(n279), .IN1(
        \add_42/carry[233] ), .COUT(\add_42/carry[234] ), .SUM(o[233]) );
  FADDER \add_42/U1_234  ( .CIN(sreg[234]), .IN0(n278), .IN1(
        \add_42/carry[234] ), .COUT(\add_42/carry[235] ), .SUM(o[234]) );
  FADDER \add_42/U1_235  ( .CIN(sreg[235]), .IN0(n277), .IN1(
        \add_42/carry[235] ), .COUT(\add_42/carry[236] ), .SUM(o[235]) );
  FADDER \add_42/U1_236  ( .CIN(sreg[236]), .IN0(n276), .IN1(
        \add_42/carry[236] ), .COUT(\add_42/carry[237] ), .SUM(o[236]) );
  FADDER \add_42/U1_237  ( .CIN(sreg[237]), .IN0(n275), .IN1(
        \add_42/carry[237] ), .COUT(\add_42/carry[238] ), .SUM(o[237]) );
  FADDER \add_42/U1_238  ( .CIN(sreg[238]), .IN0(n274), .IN1(
        \add_42/carry[238] ), .COUT(\add_42/carry[239] ), .SUM(o[238]) );
  FADDER \add_42/U1_239  ( .CIN(sreg[239]), .IN0(n273), .IN1(
        \add_42/carry[239] ), .COUT(\add_42/carry[240] ), .SUM(o[239]) );
  FADDER \add_42/U1_240  ( .CIN(sreg[240]), .IN0(n272), .IN1(
        \add_42/carry[240] ), .COUT(\add_42/carry[241] ), .SUM(o[240]) );
  FADDER \add_42/U1_241  ( .CIN(sreg[241]), .IN0(n271), .IN1(
        \add_42/carry[241] ), .COUT(\add_42/carry[242] ), .SUM(o[241]) );
  FADDER \add_42/U1_242  ( .CIN(sreg[242]), .IN0(n270), .IN1(
        \add_42/carry[242] ), .COUT(\add_42/carry[243] ), .SUM(o[242]) );
  FADDER \add_42/U1_243  ( .CIN(sreg[243]), .IN0(n269), .IN1(
        \add_42/carry[243] ), .COUT(\add_42/carry[244] ), .SUM(o[243]) );
  FADDER \add_42/U1_244  ( .CIN(sreg[244]), .IN0(n268), .IN1(
        \add_42/carry[244] ), .COUT(\add_42/carry[245] ), .SUM(o[244]) );
  FADDER \add_42/U1_245  ( .CIN(sreg[245]), .IN0(n267), .IN1(
        \add_42/carry[245] ), .COUT(\add_42/carry[246] ), .SUM(o[245]) );
  FADDER \add_42/U1_246  ( .CIN(sreg[246]), .IN0(n266), .IN1(
        \add_42/carry[246] ), .COUT(\add_42/carry[247] ), .SUM(o[246]) );
  FADDER \add_42/U1_247  ( .CIN(sreg[247]), .IN0(n265), .IN1(
        \add_42/carry[247] ), .COUT(\add_42/carry[248] ), .SUM(o[247]) );
  FADDER \add_42/U1_248  ( .CIN(sreg[248]), .IN0(n264), .IN1(
        \add_42/carry[248] ), .COUT(\add_42/carry[249] ), .SUM(o[248]) );
  FADDER \add_42/U1_249  ( .CIN(sreg[249]), .IN0(n263), .IN1(
        \add_42/carry[249] ), .COUT(\add_42/carry[250] ), .SUM(o[249]) );
  FADDER \add_42/U1_250  ( .CIN(sreg[250]), .IN0(n262), .IN1(
        \add_42/carry[250] ), .COUT(\add_42/carry[251] ), .SUM(o[250]) );
  FADDER \add_42/U1_251  ( .CIN(sreg[251]), .IN0(n261), .IN1(
        \add_42/carry[251] ), .COUT(\add_42/carry[252] ), .SUM(o[251]) );
  FADDER \add_42/U1_252  ( .CIN(sreg[252]), .IN0(n260), .IN1(
        \add_42/carry[252] ), .COUT(\add_42/carry[253] ), .SUM(o[252]) );
  FADDER \add_42/U1_253  ( .CIN(sreg[253]), .IN0(n259), .IN1(
        \add_42/carry[253] ), .COUT(\add_42/carry[254] ), .SUM(o[253]) );
  FADDER \add_42/U1_254  ( .CIN(sreg[254]), .IN0(n258), .IN1(
        \add_42/carry[254] ), .COUT(\add_42/carry[255] ), .SUM(o[254]) );
  AND U261 ( .A(sreg[127]), .B(n385), .Z(\add_42/carry[128] ) );
  XOR U262 ( .A(n385), .B(sreg[127]), .Z(o[127]) );
  AND U263 ( .A(g_input[127]), .B(e_input[0]), .Z(n258) );
  AND U264 ( .A(g_input[126]), .B(e_input[0]), .Z(n259) );
  AND U265 ( .A(g_input[125]), .B(e_input[0]), .Z(n260) );
  AND U266 ( .A(g_input[124]), .B(e_input[0]), .Z(n261) );
  AND U267 ( .A(g_input[123]), .B(e_input[0]), .Z(n262) );
  AND U268 ( .A(g_input[122]), .B(e_input[0]), .Z(n263) );
  AND U269 ( .A(g_input[121]), .B(e_input[0]), .Z(n264) );
  AND U270 ( .A(g_input[120]), .B(e_input[0]), .Z(n265) );
  AND U271 ( .A(g_input[119]), .B(e_input[0]), .Z(n266) );
  AND U272 ( .A(g_input[118]), .B(e_input[0]), .Z(n267) );
  AND U273 ( .A(g_input[117]), .B(e_input[0]), .Z(n268) );
  AND U274 ( .A(g_input[116]), .B(e_input[0]), .Z(n269) );
  AND U275 ( .A(g_input[115]), .B(e_input[0]), .Z(n270) );
  AND U276 ( .A(g_input[114]), .B(e_input[0]), .Z(n271) );
  AND U277 ( .A(g_input[113]), .B(e_input[0]), .Z(n272) );
  AND U278 ( .A(g_input[112]), .B(e_input[0]), .Z(n273) );
  AND U279 ( .A(g_input[111]), .B(e_input[0]), .Z(n274) );
  AND U280 ( .A(g_input[110]), .B(e_input[0]), .Z(n275) );
  AND U281 ( .A(g_input[109]), .B(e_input[0]), .Z(n276) );
  AND U282 ( .A(g_input[108]), .B(e_input[0]), .Z(n277) );
  AND U283 ( .A(g_input[107]), .B(e_input[0]), .Z(n278) );
  AND U284 ( .A(g_input[106]), .B(e_input[0]), .Z(n279) );
  AND U285 ( .A(g_input[105]), .B(e_input[0]), .Z(n280) );
  AND U286 ( .A(g_input[104]), .B(e_input[0]), .Z(n281) );
  AND U287 ( .A(g_input[103]), .B(e_input[0]), .Z(n282) );
  AND U288 ( .A(g_input[102]), .B(e_input[0]), .Z(n283) );
  AND U289 ( .A(g_input[101]), .B(e_input[0]), .Z(n284) );
  AND U290 ( .A(g_input[100]), .B(e_input[0]), .Z(n285) );
  AND U291 ( .A(g_input[99]), .B(e_input[0]), .Z(n286) );
  AND U292 ( .A(g_input[98]), .B(e_input[0]), .Z(n287) );
  AND U293 ( .A(g_input[97]), .B(e_input[0]), .Z(n288) );
  AND U294 ( .A(g_input[96]), .B(e_input[0]), .Z(n289) );
  AND U295 ( .A(g_input[95]), .B(e_input[0]), .Z(n290) );
  AND U296 ( .A(g_input[94]), .B(e_input[0]), .Z(n291) );
  AND U297 ( .A(g_input[93]), .B(e_input[0]), .Z(n292) );
  AND U298 ( .A(g_input[92]), .B(e_input[0]), .Z(n293) );
  AND U299 ( .A(g_input[91]), .B(e_input[0]), .Z(n294) );
  AND U300 ( .A(g_input[90]), .B(e_input[0]), .Z(n295) );
  AND U301 ( .A(g_input[89]), .B(e_input[0]), .Z(n296) );
  AND U302 ( .A(g_input[88]), .B(e_input[0]), .Z(n297) );
  AND U303 ( .A(g_input[87]), .B(e_input[0]), .Z(n298) );
  AND U304 ( .A(g_input[86]), .B(e_input[0]), .Z(n299) );
  AND U305 ( .A(g_input[85]), .B(e_input[0]), .Z(n300) );
  AND U306 ( .A(g_input[84]), .B(e_input[0]), .Z(n301) );
  AND U307 ( .A(g_input[83]), .B(e_input[0]), .Z(n302) );
  AND U308 ( .A(g_input[82]), .B(e_input[0]), .Z(n303) );
  AND U309 ( .A(g_input[81]), .B(e_input[0]), .Z(n304) );
  AND U310 ( .A(g_input[80]), .B(e_input[0]), .Z(n305) );
  AND U311 ( .A(g_input[79]), .B(e_input[0]), .Z(n306) );
  AND U312 ( .A(g_input[78]), .B(e_input[0]), .Z(n307) );
  AND U313 ( .A(g_input[77]), .B(e_input[0]), .Z(n308) );
  AND U314 ( .A(g_input[76]), .B(e_input[0]), .Z(n309) );
  AND U315 ( .A(g_input[75]), .B(e_input[0]), .Z(n310) );
  AND U316 ( .A(g_input[74]), .B(e_input[0]), .Z(n311) );
  AND U317 ( .A(g_input[73]), .B(e_input[0]), .Z(n312) );
  AND U318 ( .A(g_input[72]), .B(e_input[0]), .Z(n313) );
  AND U319 ( .A(g_input[71]), .B(e_input[0]), .Z(n314) );
  AND U320 ( .A(g_input[70]), .B(e_input[0]), .Z(n315) );
  AND U321 ( .A(g_input[69]), .B(e_input[0]), .Z(n316) );
  AND U322 ( .A(g_input[68]), .B(e_input[0]), .Z(n317) );
  AND U323 ( .A(g_input[67]), .B(e_input[0]), .Z(n318) );
  AND U324 ( .A(g_input[66]), .B(e_input[0]), .Z(n319) );
  AND U325 ( .A(g_input[65]), .B(e_input[0]), .Z(n320) );
  AND U326 ( .A(g_input[64]), .B(e_input[0]), .Z(n321) );
  AND U327 ( .A(g_input[63]), .B(e_input[0]), .Z(n322) );
  AND U328 ( .A(g_input[62]), .B(e_input[0]), .Z(n323) );
  AND U329 ( .A(g_input[61]), .B(e_input[0]), .Z(n324) );
  AND U330 ( .A(g_input[60]), .B(e_input[0]), .Z(n325) );
  AND U331 ( .A(g_input[59]), .B(e_input[0]), .Z(n326) );
  AND U332 ( .A(g_input[58]), .B(e_input[0]), .Z(n327) );
  AND U333 ( .A(g_input[57]), .B(e_input[0]), .Z(n328) );
  AND U334 ( .A(g_input[56]), .B(e_input[0]), .Z(n329) );
  AND U335 ( .A(g_input[55]), .B(e_input[0]), .Z(n330) );
  AND U336 ( .A(g_input[54]), .B(e_input[0]), .Z(n331) );
  AND U337 ( .A(g_input[53]), .B(e_input[0]), .Z(n332) );
  AND U338 ( .A(g_input[52]), .B(e_input[0]), .Z(n333) );
  AND U339 ( .A(g_input[51]), .B(e_input[0]), .Z(n334) );
  AND U340 ( .A(g_input[50]), .B(e_input[0]), .Z(n335) );
  AND U341 ( .A(g_input[49]), .B(e_input[0]), .Z(n336) );
  AND U342 ( .A(g_input[48]), .B(e_input[0]), .Z(n337) );
  AND U343 ( .A(g_input[47]), .B(e_input[0]), .Z(n338) );
  AND U344 ( .A(g_input[46]), .B(e_input[0]), .Z(n339) );
  AND U345 ( .A(g_input[45]), .B(e_input[0]), .Z(n340) );
  AND U346 ( .A(g_input[44]), .B(e_input[0]), .Z(n341) );
  AND U347 ( .A(g_input[43]), .B(e_input[0]), .Z(n342) );
  AND U348 ( .A(g_input[42]), .B(e_input[0]), .Z(n343) );
  AND U349 ( .A(g_input[41]), .B(e_input[0]), .Z(n344) );
  AND U350 ( .A(g_input[40]), .B(e_input[0]), .Z(n345) );
  AND U351 ( .A(g_input[39]), .B(e_input[0]), .Z(n346) );
  AND U352 ( .A(g_input[38]), .B(e_input[0]), .Z(n347) );
  AND U353 ( .A(g_input[37]), .B(e_input[0]), .Z(n348) );
  AND U354 ( .A(g_input[36]), .B(e_input[0]), .Z(n349) );
  AND U355 ( .A(g_input[35]), .B(e_input[0]), .Z(n350) );
  AND U356 ( .A(g_input[34]), .B(e_input[0]), .Z(n351) );
  AND U357 ( .A(g_input[33]), .B(e_input[0]), .Z(n352) );
  AND U358 ( .A(g_input[32]), .B(e_input[0]), .Z(n353) );
  AND U359 ( .A(g_input[31]), .B(e_input[0]), .Z(n354) );
  AND U360 ( .A(g_input[30]), .B(e_input[0]), .Z(n355) );
  AND U361 ( .A(g_input[29]), .B(e_input[0]), .Z(n356) );
  AND U362 ( .A(g_input[28]), .B(e_input[0]), .Z(n357) );
  AND U363 ( .A(g_input[27]), .B(e_input[0]), .Z(n358) );
  AND U364 ( .A(g_input[26]), .B(e_input[0]), .Z(n359) );
  AND U365 ( .A(g_input[25]), .B(e_input[0]), .Z(n360) );
  AND U366 ( .A(g_input[24]), .B(e_input[0]), .Z(n361) );
  AND U367 ( .A(g_input[23]), .B(e_input[0]), .Z(n362) );
  AND U368 ( .A(g_input[22]), .B(e_input[0]), .Z(n363) );
  AND U369 ( .A(g_input[21]), .B(e_input[0]), .Z(n364) );
  AND U370 ( .A(g_input[20]), .B(e_input[0]), .Z(n365) );
  AND U371 ( .A(g_input[19]), .B(e_input[0]), .Z(n366) );
  AND U372 ( .A(g_input[18]), .B(e_input[0]), .Z(n367) );
  AND U373 ( .A(g_input[17]), .B(e_input[0]), .Z(n368) );
  AND U374 ( .A(g_input[16]), .B(e_input[0]), .Z(n369) );
  AND U375 ( .A(g_input[15]), .B(e_input[0]), .Z(n370) );
  AND U376 ( .A(g_input[14]), .B(e_input[0]), .Z(n371) );
  AND U377 ( .A(g_input[13]), .B(e_input[0]), .Z(n372) );
  AND U378 ( .A(g_input[12]), .B(e_input[0]), .Z(n373) );
  AND U379 ( .A(g_input[11]), .B(e_input[0]), .Z(n374) );
  AND U380 ( .A(g_input[10]), .B(e_input[0]), .Z(n375) );
  AND U381 ( .A(g_input[9]), .B(e_input[0]), .Z(n376) );
  AND U382 ( .A(g_input[8]), .B(e_input[0]), .Z(n377) );
  AND U383 ( .A(g_input[7]), .B(e_input[0]), .Z(n378) );
  AND U384 ( .A(g_input[6]), .B(e_input[0]), .Z(n379) );
  AND U385 ( .A(g_input[5]), .B(e_input[0]), .Z(n380) );
  AND U386 ( .A(g_input[4]), .B(e_input[0]), .Z(n381) );
  AND U387 ( .A(g_input[3]), .B(e_input[0]), .Z(n382) );
  AND U388 ( .A(g_input[2]), .B(e_input[0]), .Z(n383) );
  AND U389 ( .A(g_input[1]), .B(e_input[0]), .Z(n384) );
  AND U390 ( .A(g_input[0]), .B(e_input[0]), .Z(n385) );
endmodule

