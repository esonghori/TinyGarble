
module alu ( x, y, c, o );
  input [7:0] x;
  input [7:0] y;
  input [2:0] c;
  output [15:0] o;
  wire   \C1/Z_7 , \C1/Z_6 , \C1/Z_5 , \C1/Z_4 , \C1/Z_3 , \C1/Z_2 , \C1/Z_1 ,
         \DP_OP_20_64_5734/n173 , \DP_OP_20_64_5734/n166 ,
         \DP_OP_20_64_5734/n165 , \DP_OP_20_64_5734/n164 ,
         \DP_OP_20_64_5734/n156 , \DP_OP_20_64_5734/n155 ,
         \DP_OP_20_64_5734/n142 , \DP_OP_20_64_5734/n141 ,
         \DP_OP_20_64_5734/n140 , \DP_OP_20_64_5734/n139 ,
         \DP_OP_20_64_5734/n138 , \DP_OP_20_64_5734/n137 ,
         \DP_OP_20_64_5734/n136 , \DP_OP_20_64_5734/n129 ,
         \DP_OP_20_64_5734/n128 , \DP_OP_20_64_5734/n127 ,
         \DP_OP_20_64_5734/n126 , \DP_OP_20_64_5734/n125 ,
         \DP_OP_20_64_5734/n123 , \DP_OP_20_64_5734/n111 ,
         \DP_OP_20_64_5734/n110 , \DP_OP_20_64_5734/n109 ,
         \DP_OP_20_64_5734/n107 , \DP_OP_20_64_5734/n105 ,
         \DP_OP_20_64_5734/n98 , \DP_OP_20_64_5734/n97 ,
         \DP_OP_20_64_5734/n96 , \DP_OP_20_64_5734/n94 ,
         \DP_OP_20_64_5734/n90 , \DP_OP_20_64_5734/n76 ,
         \DP_OP_20_64_5734/n75 , \DP_OP_20_64_5734/n74 ,
         \DP_OP_20_64_5734/n70 , \DP_OP_20_64_5734/n68 ,
         \DP_OP_20_64_5734/n57 , \DP_OP_20_64_5734/n56 ,
         \DP_OP_20_64_5734/n55 , \DP_OP_20_64_5734/n53 ,
         \DP_OP_20_64_5734/n49 , \DP_OP_20_64_5734/n35 ,
         \DP_OP_20_64_5734/n34 , \DP_OP_20_64_5734/n33 ,
         \DP_OP_20_64_5734/n31 , \DP_OP_20_64_5734/n29 ,
         \DP_OP_20_64_5734/n23 , \DP_OP_20_64_5734/n22 ,
         \DP_OP_20_64_5734/n21 , \DP_OP_20_64_5734/n19 ,
         \DP_OP_20_64_5734/n17 , n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766;

  XOR \DP_OP_20_64_5734/U88  ( .A(x[0]), .B(\DP_OP_20_64_5734/n173 ), .Z(
        \DP_OP_20_64_5734/n164 ) );
  XOR \DP_OP_20_64_5734/U87  ( .A(x[1]), .B(\C1/Z_1 ), .Z(
        \DP_OP_20_64_5734/n142 ) );
  XOR \DP_OP_20_64_5734/U80  ( .A(\DP_OP_20_64_5734/n156 ), .B(
        \DP_OP_20_64_5734/n142 ), .Z(\DP_OP_20_64_5734/n165 ) );
  XOR \DP_OP_20_64_5734/U79  ( .A(x[2]), .B(\C1/Z_2 ), .Z(
        \DP_OP_20_64_5734/n141 ) );
  XOR \DP_OP_20_64_5734/U78  ( .A(\DP_OP_20_64_5734/n155 ), .B(
        \DP_OP_20_64_5734/n141 ), .Z(\DP_OP_20_64_5734/n166 ) );
  XOR \DP_OP_20_64_5734/U69  ( .A(x[3]), .B(\C1/Z_3 ), .Z(
        \DP_OP_20_64_5734/n140 ) );
  XOR \DP_OP_20_64_5734/U67  ( .A(x[4]), .B(\C1/Z_4 ), .Z(
        \DP_OP_20_64_5734/n139 ) );
  XOR \DP_OP_20_64_5734/U57  ( .A(x[5]), .B(\C1/Z_5 ), .Z(
        \DP_OP_20_64_5734/n138 ) );
  XOR \DP_OP_20_64_5734/U49  ( .A(x[6]), .B(\C1/Z_6 ), .Z(
        \DP_OP_20_64_5734/n137 ) );
  XOR \DP_OP_20_64_5734/U30  ( .A(x[7]), .B(\C1/Z_7 ), .Z(
        \DP_OP_20_64_5734/n136 ) );
  IV \DP_OP_20_64_5734/U110  ( .A(\C1/Z_7 ), .Z(\DP_OP_20_64_5734/n17 ) );
  IV \DP_OP_20_64_5734/U39  ( .A(\DP_OP_20_64_5734/n136 ), .Z(
        \DP_OP_20_64_5734/n19 ) );
  NOR \DP_OP_20_64_5734/U56  ( .A(\DP_OP_20_64_5734/n17 ), .B(n671), .Z(
        \DP_OP_20_64_5734/n21 ) );
  NOR \DP_OP_20_64_5734/U66  ( .A(\DP_OP_20_64_5734/n19 ), .B(
        \DP_OP_20_64_5734/n35 ), .Z(\DP_OP_20_64_5734/n22 ) );
  NOR \DP_OP_20_64_5734/U76  ( .A(\DP_OP_20_64_5734/n21 ), .B(
        \DP_OP_20_64_5734/n22 ), .Z(\DP_OP_20_64_5734/n23 ) );
  IV \DP_OP_20_64_5734/U19  ( .A(\C1/Z_6 ), .Z(\DP_OP_20_64_5734/n29 ) );
  IV \DP_OP_20_64_5734/U38  ( .A(\DP_OP_20_64_5734/n137 ), .Z(
        \DP_OP_20_64_5734/n31 ) );
  NOR \DP_OP_20_64_5734/U55  ( .A(\DP_OP_20_64_5734/n29 ), .B(n574), .Z(
        \DP_OP_20_64_5734/n33 ) );
  NOR \DP_OP_20_64_5734/U65  ( .A(\DP_OP_20_64_5734/n31 ), .B(
        \DP_OP_20_64_5734/n57 ), .Z(\DP_OP_20_64_5734/n34 ) );
  NOR \DP_OP_20_64_5734/U75  ( .A(\DP_OP_20_64_5734/n33 ), .B(
        \DP_OP_20_64_5734/n34 ), .Z(\DP_OP_20_64_5734/n35 ) );
  IV \DP_OP_20_64_5734/U17  ( .A(\C1/Z_5 ), .Z(\DP_OP_20_64_5734/n49 ) );
  IV \DP_OP_20_64_5734/U36  ( .A(\DP_OP_20_64_5734/n138 ), .Z(
        \DP_OP_20_64_5734/n53 ) );
  NOR \DP_OP_20_64_5734/U54  ( .A(\DP_OP_20_64_5734/n49 ), .B(n543), .Z(
        \DP_OP_20_64_5734/n55 ) );
  NOR \DP_OP_20_64_5734/U64  ( .A(\DP_OP_20_64_5734/n53 ), .B(
        \DP_OP_20_64_5734/n76 ), .Z(\DP_OP_20_64_5734/n56 ) );
  NOR \DP_OP_20_64_5734/U74  ( .A(\DP_OP_20_64_5734/n55 ), .B(
        \DP_OP_20_64_5734/n56 ), .Z(\DP_OP_20_64_5734/n57 ) );
  IV \DP_OP_20_64_5734/U16  ( .A(\C1/Z_4 ), .Z(\DP_OP_20_64_5734/n68 ) );
  IV \DP_OP_20_64_5734/U35  ( .A(\DP_OP_20_64_5734/n139 ), .Z(
        \DP_OP_20_64_5734/n70 ) );
  NOR \DP_OP_20_64_5734/U53  ( .A(\DP_OP_20_64_5734/n68 ), .B(n534), .Z(
        \DP_OP_20_64_5734/n74 ) );
  NOR \DP_OP_20_64_5734/U63  ( .A(\DP_OP_20_64_5734/n70 ), .B(
        \DP_OP_20_64_5734/n98 ), .Z(\DP_OP_20_64_5734/n75 ) );
  NOR \DP_OP_20_64_5734/U73  ( .A(\DP_OP_20_64_5734/n74 ), .B(
        \DP_OP_20_64_5734/n75 ), .Z(\DP_OP_20_64_5734/n76 ) );
  IV \DP_OP_20_64_5734/U14  ( .A(\C1/Z_3 ), .Z(\DP_OP_20_64_5734/n90 ) );
  IV \DP_OP_20_64_5734/U33  ( .A(\DP_OP_20_64_5734/n140 ), .Z(
        \DP_OP_20_64_5734/n94 ) );
  NOR \DP_OP_20_64_5734/U52  ( .A(\DP_OP_20_64_5734/n90 ), .B(n515), .Z(
        \DP_OP_20_64_5734/n96 ) );
  NOR \DP_OP_20_64_5734/U62  ( .A(\DP_OP_20_64_5734/n94 ), .B(
        \DP_OP_20_64_5734/n111 ), .Z(\DP_OP_20_64_5734/n97 ) );
  NOR \DP_OP_20_64_5734/U72  ( .A(\DP_OP_20_64_5734/n96 ), .B(
        \DP_OP_20_64_5734/n97 ), .Z(\DP_OP_20_64_5734/n98 ) );
  IV \DP_OP_20_64_5734/U13  ( .A(\C1/Z_2 ), .Z(\DP_OP_20_64_5734/n105 ) );
  IV \DP_OP_20_64_5734/U32  ( .A(\DP_OP_20_64_5734/n141 ), .Z(
        \DP_OP_20_64_5734/n107 ) );
  NOR \DP_OP_20_64_5734/U51  ( .A(\DP_OP_20_64_5734/n105 ), .B(n444), .Z(
        \DP_OP_20_64_5734/n109 ) );
  NOR \DP_OP_20_64_5734/U61  ( .A(\DP_OP_20_64_5734/n107 ), .B(
        \DP_OP_20_64_5734/n129 ), .Z(\DP_OP_20_64_5734/n110 ) );
  NOR \DP_OP_20_64_5734/U71  ( .A(\DP_OP_20_64_5734/n109 ), .B(
        \DP_OP_20_64_5734/n110 ), .Z(\DP_OP_20_64_5734/n111 ) );
  IV \DP_OP_20_64_5734/U11  ( .A(\C1/Z_1 ), .Z(\DP_OP_20_64_5734/n123 ) );
  IV \DP_OP_20_64_5734/U3  ( .A(\DP_OP_20_64_5734/n142 ), .Z(
        \DP_OP_20_64_5734/n125 ) );
  IV \DP_OP_20_64_5734/U4  ( .A(\DP_OP_20_64_5734/n156 ), .Z(
        \DP_OP_20_64_5734/n126 ) );
  NOR \DP_OP_20_64_5734/U5  ( .A(\DP_OP_20_64_5734/n123 ), .B(n363), .Z(
        \DP_OP_20_64_5734/n127 ) );
  NOR \DP_OP_20_64_5734/U6  ( .A(\DP_OP_20_64_5734/n125 ), .B(
        \DP_OP_20_64_5734/n126 ), .Z(\DP_OP_20_64_5734/n128 ) );
  NOR \DP_OP_20_64_5734/U7  ( .A(\DP_OP_20_64_5734/n127 ), .B(
        \DP_OP_20_64_5734/n128 ), .Z(\DP_OP_20_64_5734/n129 ) );
  IV \DP_OP_20_64_5734/U8  ( .A(\DP_OP_20_64_5734/n129 ), .Z(
        \DP_OP_20_64_5734/n155 ) );
  NOR \DP_OP_20_64_5734/AND2i  ( .A(n307), .B(n145), .Z(
        \DP_OP_20_64_5734/n156 ) );
  XOR U53 ( .A(n515), .B(n215), .Z(n58) );
  NOR U54 ( .A(n744), .B(n58), .Z(n59) );
  XOR U55 ( .A(n212), .B(n209), .Z(n60) );
  XOR U56 ( .A(n207), .B(n60), .Z(n61) );
  NOR U57 ( .A(n747), .B(n61), .Z(n62) );
  NOR U58 ( .A(n59), .B(n62), .Z(n63) );
  IV U59 ( .A(n63), .Z(n64) );
  XOR U60 ( .A(\DP_OP_20_64_5734/n111 ), .B(\DP_OP_20_64_5734/n140 ), .Z(n65)
         );
  NOR U61 ( .A(n714), .B(n65), .Z(n66) );
  XOR U62 ( .A(n515), .B(n604), .Z(n67) );
  XOR U63 ( .A(n217), .B(n67), .Z(n68) );
  NOR U64 ( .A(n745), .B(n68), .Z(n69) );
  NOR U65 ( .A(n66), .B(n69), .Z(n70) );
  IV U66 ( .A(n70), .Z(n71) );
  NOR U67 ( .A(n64), .B(n71), .Z(n72) );
  IV U68 ( .A(n72), .Z(o[3]) );
  XOR U69 ( .A(n534), .B(n255), .Z(n73) );
  NOR U70 ( .A(n744), .B(n73), .Z(n74) );
  XOR U71 ( .A(n251), .B(n248), .Z(n75) );
  XOR U72 ( .A(n247), .B(n75), .Z(n76) );
  NOR U73 ( .A(n747), .B(n76), .Z(n77) );
  NOR U74 ( .A(n74), .B(n77), .Z(n78) );
  IV U75 ( .A(n78), .Z(n79) );
  XOR U76 ( .A(\DP_OP_20_64_5734/n98 ), .B(\DP_OP_20_64_5734/n139 ), .Z(n80)
         );
  NOR U77 ( .A(n714), .B(n80), .Z(n81) );
  XOR U78 ( .A(n534), .B(n584), .Z(n82) );
  XOR U79 ( .A(n259), .B(n82), .Z(n83) );
  NOR U80 ( .A(n745), .B(n83), .Z(n84) );
  NOR U81 ( .A(n81), .B(n84), .Z(n85) );
  IV U82 ( .A(n85), .Z(n86) );
  NOR U83 ( .A(n79), .B(n86), .Z(n87) );
  IV U84 ( .A(n87), .Z(o[4]) );
  IV U85 ( .A(n353), .Z(n88) );
  IV U86 ( .A(n354), .Z(n89) );
  NOR U87 ( .A(n353), .B(n89), .Z(n90) );
  NOR U88 ( .A(n354), .B(n88), .Z(n91) );
  NOR U89 ( .A(n352), .B(n91), .Z(n92) );
  NOR U90 ( .A(n90), .B(n92), .Z(n412) );
  XOR U91 ( .A(n543), .B(n299), .Z(n93) );
  NOR U92 ( .A(n744), .B(n93), .Z(n94) );
  XOR U93 ( .A(n295), .B(n293), .Z(n95) );
  XOR U94 ( .A(n291), .B(n95), .Z(n96) );
  NOR U95 ( .A(n747), .B(n96), .Z(n97) );
  NOR U96 ( .A(n94), .B(n97), .Z(n98) );
  IV U97 ( .A(n98), .Z(n99) );
  XOR U98 ( .A(\DP_OP_20_64_5734/n76 ), .B(\DP_OP_20_64_5734/n138 ), .Z(n100)
         );
  NOR U99 ( .A(n714), .B(n100), .Z(n101) );
  XOR U100 ( .A(n543), .B(n540), .Z(n102) );
  XOR U101 ( .A(n301), .B(n102), .Z(n103) );
  NOR U102 ( .A(n745), .B(n103), .Z(n104) );
  NOR U103 ( .A(n101), .B(n104), .Z(n105) );
  IV U104 ( .A(n105), .Z(n106) );
  NOR U105 ( .A(n99), .B(n106), .Z(n107) );
  IV U106 ( .A(n107), .Z(o[5]) );
  XOR U107 ( .A(n574), .B(n413), .Z(n108) );
  NOR U108 ( .A(n744), .B(n108), .Z(n109) );
  XOR U109 ( .A(n352), .B(n354), .Z(n110) );
  XOR U110 ( .A(n353), .B(n110), .Z(n111) );
  NOR U111 ( .A(n747), .B(n111), .Z(n112) );
  NOR U112 ( .A(n109), .B(n112), .Z(n113) );
  IV U113 ( .A(n113), .Z(n114) );
  XOR U114 ( .A(\DP_OP_20_64_5734/n57 ), .B(\DP_OP_20_64_5734/n137 ), .Z(n115)
         );
  NOR U115 ( .A(n714), .B(n115), .Z(n116) );
  XOR U116 ( .A(n574), .B(n554), .Z(n117) );
  XOR U117 ( .A(n418), .B(n117), .Z(n118) );
  NOR U118 ( .A(n745), .B(n118), .Z(n119) );
  NOR U119 ( .A(n116), .B(n119), .Z(n120) );
  IV U120 ( .A(n120), .Z(n121) );
  NOR U121 ( .A(n114), .B(n121), .Z(n122) );
  IV U122 ( .A(n122), .Z(o[6]) );
  XOR U123 ( .A(\DP_OP_20_64_5734/n35 ), .B(\DP_OP_20_64_5734/n136 ), .Z(n123)
         );
  NOR U124 ( .A(n714), .B(n123), .Z(n124) );
  XOR U125 ( .A(n671), .B(n415), .Z(n125) );
  NOR U126 ( .A(n744), .B(n125), .Z(n126) );
  XOR U127 ( .A(n412), .B(n411), .Z(n127) );
  XOR U128 ( .A(n410), .B(n127), .Z(n128) );
  NOR U129 ( .A(n747), .B(n128), .Z(n129) );
  XOR U130 ( .A(n671), .B(n669), .Z(n130) );
  XOR U131 ( .A(n423), .B(n130), .Z(n131) );
  NOR U132 ( .A(n745), .B(n131), .Z(n132) );
  NOR U133 ( .A(n126), .B(n129), .Z(n133) );
  IV U134 ( .A(n133), .Z(n134) );
  NOR U135 ( .A(n124), .B(n132), .Z(n135) );
  IV U136 ( .A(n135), .Z(n136) );
  NOR U137 ( .A(n134), .B(n136), .Z(n137) );
  IV U138 ( .A(n137), .Z(o[7]) );
  IV U139 ( .A(c[1]), .Z(n157) );
  IV U140 ( .A(c[0]), .Z(n158) );
  NOR U141 ( .A(c[1]), .B(c[0]), .Z(n138) );
  IV U142 ( .A(n138), .Z(n434) );
  NOR U143 ( .A(c[2]), .B(n434), .Z(n139) );
  IV U144 ( .A(n139), .Z(n142) );
  NOR U145 ( .A(n142), .B(n669), .Z(\C1/Z_7 ) );
  NOR U146 ( .A(n142), .B(n554), .Z(\C1/Z_6 ) );
  NOR U147 ( .A(n142), .B(n540), .Z(\C1/Z_5 ) );
  NOR U148 ( .A(n142), .B(n584), .Z(\C1/Z_4 ) );
  NOR U149 ( .A(n142), .B(n604), .Z(\C1/Z_3 ) );
  NOR U150 ( .A(n142), .B(n489), .Z(\C1/Z_2 ) );
  NOR U151 ( .A(n142), .B(n358), .Z(\C1/Z_1 ) );
  NOR U152 ( .A(c[2]), .B(n158), .Z(n140) );
  IV U153 ( .A(n140), .Z(n141) );
  NOR U154 ( .A(n157), .B(n141), .Z(n144) );
  NOR U155 ( .A(n142), .B(n306), .Z(n143) );
  NOR U156 ( .A(n144), .B(n143), .Z(n145) );
  IV U157 ( .A(n145), .Z(\DP_OP_20_64_5734/n173 ) );
  IV U158 ( .A(\DP_OP_20_64_5734/n164 ), .Z(n146) );
  NOR U159 ( .A(n714), .B(n146), .Z(n147) );
  NOR U160 ( .A(n147), .B(n720), .Z(n148) );
  IV U161 ( .A(n148), .Z(n749) );
  IV U162 ( .A(\DP_OP_20_64_5734/n165 ), .Z(n149) );
  NOR U163 ( .A(n714), .B(n149), .Z(n150) );
  NOR U164 ( .A(n150), .B(n725), .Z(n151) );
  IV U165 ( .A(n151), .Z(n754) );
  IV U166 ( .A(\DP_OP_20_64_5734/n166 ), .Z(n152) );
  NOR U167 ( .A(n714), .B(n152), .Z(n153) );
  NOR U168 ( .A(n153), .B(n730), .Z(n154) );
  IV U169 ( .A(n154), .Z(n759) );
  NOR U170 ( .A(n714), .B(\DP_OP_20_64_5734/n23 ), .Z(n155) );
  NOR U171 ( .A(n155), .B(n735), .Z(n156) );
  IV U172 ( .A(n156), .Z(n764) );
  IV U173 ( .A(n717), .Z(n740) );
  IV U174 ( .A(n710), .Z(n741) );
  IV U175 ( .A(n711), .Z(n742) );
  IV U176 ( .A(n715), .Z(n743) );
  IV U177 ( .A(n716), .Z(n744) );
  IV U178 ( .A(n719), .Z(n745) );
  IV U179 ( .A(c[2]), .Z(n746) );
  IV U180 ( .A(n718), .Z(n747) );
  IV U181 ( .A(x[0]), .Z(n307) );
  IV U182 ( .A(y[0]), .Z(n306) );
  NOR U183 ( .A(n307), .B(n306), .Z(n159) );
  IV U184 ( .A(n159), .Z(n748) );
  XOR U185 ( .A(n307), .B(y[0]), .Z(n750) );
  IV U186 ( .A(n723), .Z(n751) );
  IV U187 ( .A(n724), .Z(o[0]) );
  IV U188 ( .A(x[1]), .Z(n363) );
  NOR U189 ( .A(n363), .B(n306), .Z(n160) );
  IV U190 ( .A(n160), .Z(n178) );
  IV U191 ( .A(y[1]), .Z(n358) );
  NOR U192 ( .A(n358), .B(n307), .Z(n162) );
  XOR U193 ( .A(n178), .B(n162), .Z(n752) );
  XOR U194 ( .A(n363), .B(n307), .Z(n753) );
  NOR U195 ( .A(x[0]), .B(n306), .Z(n167) );
  IV U196 ( .A(n167), .Z(n166) );
  XOR U197 ( .A(n358), .B(n363), .Z(n161) );
  XOR U198 ( .A(n166), .B(n161), .Z(n755) );
  IV U199 ( .A(n728), .Z(n756) );
  IV U200 ( .A(n729), .Z(o[1]) );
  IV U201 ( .A(x[2]), .Z(n444) );
  IV U202 ( .A(n162), .Z(n177) );
  NOR U203 ( .A(n177), .B(n363), .Z(n163) );
  XOR U204 ( .A(n444), .B(n163), .Z(n164) );
  NOR U205 ( .A(n306), .B(n164), .Z(n181) );
  NOR U206 ( .A(n358), .B(n363), .Z(n165) );
  IV U207 ( .A(n165), .Z(n174) );
  IV U208 ( .A(y[2]), .Z(n489) );
  NOR U209 ( .A(n489), .B(n307), .Z(n172) );
  XOR U210 ( .A(n174), .B(n172), .Z(n182) );
  XOR U211 ( .A(n181), .B(n182), .Z(n757) );
  NOR U212 ( .A(x[1]), .B(x[0]), .Z(n186) );
  XOR U213 ( .A(n444), .B(n186), .Z(n758) );
  NOR U214 ( .A(x[1]), .B(n166), .Z(n170) );
  NOR U215 ( .A(n167), .B(n363), .Z(n168) );
  NOR U216 ( .A(n358), .B(n168), .Z(n169) );
  NOR U217 ( .A(n170), .B(n169), .Z(n188) );
  XOR U218 ( .A(n489), .B(n444), .Z(n171) );
  XOR U219 ( .A(n188), .B(n171), .Z(n760) );
  IV U220 ( .A(n733), .Z(n761) );
  IV U221 ( .A(n734), .Z(o[2]) );
  NOR U222 ( .A(n444), .B(n358), .Z(n198) );
  IV U223 ( .A(n172), .Z(n173) );
  NOR U224 ( .A(n174), .B(n173), .Z(n175) );
  IV U225 ( .A(n175), .Z(n200) );
  XOR U226 ( .A(n198), .B(n200), .Z(n202) );
  NOR U227 ( .A(n489), .B(n363), .Z(n194) );
  IV U228 ( .A(y[3]), .Z(n604) );
  NOR U229 ( .A(n604), .B(n307), .Z(n176) );
  IV U230 ( .A(n176), .Z(n195) );
  XOR U231 ( .A(n194), .B(n195), .Z(n201) );
  XOR U232 ( .A(n202), .B(n201), .Z(n212) );
  IV U233 ( .A(x[3]), .Z(n515) );
  NOR U234 ( .A(n515), .B(n306), .Z(n208) );
  IV U235 ( .A(n208), .Z(n209) );
  NOR U236 ( .A(n178), .B(n177), .Z(n179) );
  IV U237 ( .A(n179), .Z(n180) );
  NOR U238 ( .A(n444), .B(n180), .Z(n185) );
  IV U239 ( .A(n181), .Z(n183) );
  NOR U240 ( .A(n183), .B(n182), .Z(n184) );
  NOR U241 ( .A(n185), .B(n184), .Z(n210) );
  IV U242 ( .A(n210), .Z(n207) );
  IV U243 ( .A(n186), .Z(n187) );
  NOR U244 ( .A(x[2]), .B(n187), .Z(n215) );
  NOR U245 ( .A(x[2]), .B(n188), .Z(n192) );
  IV U246 ( .A(n188), .Z(n189) );
  NOR U247 ( .A(n444), .B(n189), .Z(n190) );
  NOR U248 ( .A(n190), .B(n489), .Z(n191) );
  NOR U249 ( .A(n192), .B(n191), .Z(n217) );
  NOR U250 ( .A(n604), .B(n363), .Z(n193) );
  IV U251 ( .A(n193), .Z(n236) );
  IV U252 ( .A(y[4]), .Z(n584) );
  NOR U253 ( .A(n584), .B(n307), .Z(n234) );
  XOR U254 ( .A(n236), .B(n234), .Z(n226) );
  IV U255 ( .A(n194), .Z(n196) );
  NOR U256 ( .A(n196), .B(n195), .Z(n225) );
  IV U257 ( .A(n225), .Z(n223) );
  NOR U258 ( .A(n489), .B(n444), .Z(n224) );
  IV U259 ( .A(n224), .Z(n222) );
  XOR U260 ( .A(n223), .B(n222), .Z(n197) );
  XOR U261 ( .A(n226), .B(n197), .Z(n242) );
  NOR U262 ( .A(n515), .B(n358), .Z(n241) );
  IV U263 ( .A(n241), .Z(n238) );
  IV U264 ( .A(n198), .Z(n199) );
  NOR U265 ( .A(n200), .B(n199), .Z(n204) );
  NOR U266 ( .A(n202), .B(n201), .Z(n203) );
  NOR U267 ( .A(n204), .B(n203), .Z(n239) );
  IV U268 ( .A(n239), .Z(n240) );
  XOR U269 ( .A(n238), .B(n240), .Z(n205) );
  XOR U270 ( .A(n242), .B(n205), .Z(n206) );
  IV U271 ( .A(n206), .Z(n251) );
  NOR U272 ( .A(n208), .B(n207), .Z(n214) );
  NOR U273 ( .A(n210), .B(n209), .Z(n211) );
  NOR U274 ( .A(n212), .B(n211), .Z(n213) );
  NOR U275 ( .A(n214), .B(n213), .Z(n250) );
  IV U276 ( .A(n250), .Z(n248) );
  IV U277 ( .A(x[4]), .Z(n534) );
  NOR U278 ( .A(n534), .B(n306), .Z(n249) );
  IV U279 ( .A(n249), .Z(n247) );
  IV U280 ( .A(n215), .Z(n216) );
  NOR U281 ( .A(x[3]), .B(n216), .Z(n255) );
  NOR U282 ( .A(x[3]), .B(n217), .Z(n221) );
  IV U283 ( .A(n217), .Z(n218) );
  NOR U284 ( .A(n515), .B(n218), .Z(n219) );
  NOR U285 ( .A(n219), .B(n604), .Z(n220) );
  NOR U286 ( .A(n221), .B(n220), .Z(n259) );
  NOR U287 ( .A(n515), .B(n489), .Z(n231) );
  NOR U288 ( .A(n223), .B(n222), .Z(n229) );
  NOR U289 ( .A(n225), .B(n224), .Z(n227) );
  NOR U290 ( .A(n227), .B(n226), .Z(n228) );
  NOR U291 ( .A(n229), .B(n228), .Z(n232) );
  IV U292 ( .A(n232), .Z(n230) );
  NOR U293 ( .A(n231), .B(n230), .Z(n278) );
  NOR U294 ( .A(n232), .B(n515), .Z(n280) );
  NOR U295 ( .A(n278), .B(n280), .Z(n237) );
  NOR U296 ( .A(n584), .B(n363), .Z(n262) );
  IV U297 ( .A(y[5]), .Z(n540) );
  NOR U298 ( .A(n540), .B(n307), .Z(n263) );
  XOR U299 ( .A(n262), .B(n263), .Z(n271) );
  NOR U300 ( .A(n604), .B(n444), .Z(n233) );
  IV U301 ( .A(n233), .Z(n269) );
  IV U302 ( .A(n234), .Z(n235) );
  NOR U303 ( .A(n236), .B(n235), .Z(n268) );
  XOR U304 ( .A(n269), .B(n268), .Z(n273) );
  XOR U305 ( .A(n271), .B(n273), .Z(n277) );
  XOR U306 ( .A(n237), .B(n277), .Z(n284) );
  NOR U307 ( .A(n239), .B(n238), .Z(n245) );
  NOR U308 ( .A(n241), .B(n240), .Z(n243) );
  NOR U309 ( .A(n243), .B(n242), .Z(n244) );
  NOR U310 ( .A(n245), .B(n244), .Z(n287) );
  NOR U311 ( .A(n534), .B(n358), .Z(n282) );
  XOR U312 ( .A(n287), .B(n282), .Z(n246) );
  XOR U313 ( .A(n284), .B(n246), .Z(n295) );
  IV U314 ( .A(x[5]), .Z(n543) );
  NOR U315 ( .A(n543), .B(n306), .Z(n292) );
  IV U316 ( .A(n292), .Z(n293) );
  NOR U317 ( .A(n248), .B(n247), .Z(n254) );
  NOR U318 ( .A(n250), .B(n249), .Z(n252) );
  NOR U319 ( .A(n252), .B(n251), .Z(n253) );
  NOR U320 ( .A(n254), .B(n253), .Z(n294) );
  IV U321 ( .A(n294), .Z(n291) );
  IV U322 ( .A(n255), .Z(n256) );
  NOR U323 ( .A(x[4]), .B(n256), .Z(n299) );
  IV U324 ( .A(n259), .Z(n257) );
  NOR U325 ( .A(n534), .B(n257), .Z(n258) );
  NOR U326 ( .A(n258), .B(n584), .Z(n261) );
  NOR U327 ( .A(x[4]), .B(n259), .Z(n260) );
  NOR U328 ( .A(n261), .B(n260), .Z(n301) );
  IV U329 ( .A(x[6]), .Z(n574) );
  NOR U330 ( .A(n574), .B(n306), .Z(n352) );
  NOR U331 ( .A(n584), .B(n444), .Z(n313) );
  IV U332 ( .A(n262), .Z(n265) );
  IV U333 ( .A(n263), .Z(n264) );
  NOR U334 ( .A(n265), .B(n264), .Z(n266) );
  IV U335 ( .A(n266), .Z(n315) );
  XOR U336 ( .A(n313), .B(n315), .Z(n317) );
  NOR U337 ( .A(n540), .B(n363), .Z(n308) );
  IV U338 ( .A(y[6]), .Z(n554) );
  NOR U339 ( .A(n554), .B(n307), .Z(n267) );
  IV U340 ( .A(n267), .Z(n309) );
  XOR U341 ( .A(n308), .B(n309), .Z(n316) );
  XOR U342 ( .A(n317), .B(n316), .Z(n326) );
  NOR U343 ( .A(n604), .B(n515), .Z(n322) );
  IV U344 ( .A(n322), .Z(n323) );
  IV U345 ( .A(n268), .Z(n270) );
  NOR U346 ( .A(n270), .B(n269), .Z(n275) );
  IV U347 ( .A(n271), .Z(n272) );
  NOR U348 ( .A(n273), .B(n272), .Z(n274) );
  NOR U349 ( .A(n275), .B(n274), .Z(n324) );
  IV U350 ( .A(n324), .Z(n321) );
  XOR U351 ( .A(n323), .B(n321), .Z(n276) );
  XOR U352 ( .A(n326), .B(n276), .Z(n332) );
  NOR U353 ( .A(n278), .B(n277), .Z(n279) );
  NOR U354 ( .A(n280), .B(n279), .Z(n336) );
  NOR U355 ( .A(n534), .B(n489), .Z(n334) );
  XOR U356 ( .A(n336), .B(n334), .Z(n281) );
  XOR U357 ( .A(n332), .B(n281), .Z(n344) );
  IV U358 ( .A(n282), .Z(n283) );
  NOR U359 ( .A(n284), .B(n283), .Z(n289) );
  IV U360 ( .A(n284), .Z(n285) );
  NOR U361 ( .A(x[4]), .B(n285), .Z(n286) );
  NOR U362 ( .A(n287), .B(n286), .Z(n288) );
  NOR U363 ( .A(n289), .B(n288), .Z(n341) );
  IV U364 ( .A(n341), .Z(n342) );
  NOR U365 ( .A(n543), .B(n358), .Z(n343) );
  IV U366 ( .A(n343), .Z(n340) );
  XOR U367 ( .A(n342), .B(n340), .Z(n290) );
  XOR U368 ( .A(n344), .B(n290), .Z(n354) );
  NOR U369 ( .A(n292), .B(n291), .Z(n298) );
  NOR U370 ( .A(n294), .B(n293), .Z(n296) );
  NOR U371 ( .A(n296), .B(n295), .Z(n297) );
  NOR U372 ( .A(n298), .B(n297), .Z(n353) );
  IV U373 ( .A(n299), .Z(n300) );
  NOR U374 ( .A(x[5]), .B(n300), .Z(n413) );
  NOR U375 ( .A(x[5]), .B(n301), .Z(n305) );
  IV U376 ( .A(n301), .Z(n302) );
  NOR U377 ( .A(n543), .B(n302), .Z(n303) );
  NOR U378 ( .A(n303), .B(n540), .Z(n304) );
  NOR U379 ( .A(n305), .B(n304), .Z(n418) );
  IV U380 ( .A(x[7]), .Z(n671) );
  NOR U381 ( .A(n671), .B(n306), .Z(n350) );
  NOR U382 ( .A(n554), .B(n363), .Z(n359) );
  IV U383 ( .A(y[7]), .Z(n669) );
  NOR U384 ( .A(n669), .B(n307), .Z(n360) );
  XOR U385 ( .A(n359), .B(n360), .Z(n367) );
  IV U386 ( .A(n367), .Z(n365) );
  IV U387 ( .A(n308), .Z(n310) );
  NOR U388 ( .A(n310), .B(n309), .Z(n368) );
  IV U389 ( .A(n368), .Z(n366) );
  NOR U390 ( .A(n540), .B(n444), .Z(n311) );
  IV U391 ( .A(n311), .Z(n369) );
  XOR U392 ( .A(n366), .B(n369), .Z(n312) );
  XOR U393 ( .A(n365), .B(n312), .Z(n378) );
  NOR U394 ( .A(n584), .B(n515), .Z(n377) );
  IV U395 ( .A(n377), .Z(n374) );
  IV U396 ( .A(n313), .Z(n314) );
  NOR U397 ( .A(n315), .B(n314), .Z(n319) );
  NOR U398 ( .A(n317), .B(n316), .Z(n318) );
  NOR U399 ( .A(n319), .B(n318), .Z(n375) );
  IV U400 ( .A(n375), .Z(n376) );
  XOR U401 ( .A(n374), .B(n376), .Z(n320) );
  XOR U402 ( .A(n378), .B(n320), .Z(n385) );
  IV U403 ( .A(n385), .Z(n383) );
  NOR U404 ( .A(n534), .B(n604), .Z(n386) );
  IV U405 ( .A(n386), .Z(n384) );
  NOR U406 ( .A(n322), .B(n321), .Z(n328) );
  NOR U407 ( .A(n324), .B(n323), .Z(n325) );
  NOR U408 ( .A(n326), .B(n325), .Z(n327) );
  NOR U409 ( .A(n328), .B(n327), .Z(n329) );
  IV U410 ( .A(n329), .Z(n387) );
  XOR U411 ( .A(n384), .B(n387), .Z(n330) );
  XOR U412 ( .A(n383), .B(n330), .Z(n396) );
  IV U413 ( .A(n334), .Z(n331) );
  NOR U414 ( .A(n331), .B(n332), .Z(n338) );
  IV U415 ( .A(n332), .Z(n333) );
  NOR U416 ( .A(n334), .B(n333), .Z(n335) );
  NOR U417 ( .A(n336), .B(n335), .Z(n337) );
  NOR U418 ( .A(n338), .B(n337), .Z(n393) );
  IV U419 ( .A(n393), .Z(n394) );
  NOR U420 ( .A(n543), .B(n489), .Z(n395) );
  IV U421 ( .A(n395), .Z(n392) );
  XOR U422 ( .A(n394), .B(n392), .Z(n339) );
  XOR U423 ( .A(n396), .B(n339), .Z(n404) );
  NOR U424 ( .A(n341), .B(n340), .Z(n348) );
  NOR U425 ( .A(n343), .B(n342), .Z(n346) );
  IV U426 ( .A(n344), .Z(n345) );
  NOR U427 ( .A(n346), .B(n345), .Z(n347) );
  NOR U428 ( .A(n348), .B(n347), .Z(n406) );
  NOR U429 ( .A(n574), .B(n358), .Z(n401) );
  XOR U430 ( .A(n406), .B(n401), .Z(n349) );
  XOR U431 ( .A(n404), .B(n349), .Z(n351) );
  IV U432 ( .A(n351), .Z(n411) );
  NOR U433 ( .A(n350), .B(n411), .Z(n357) );
  IV U434 ( .A(n350), .Z(n410) );
  NOR U435 ( .A(n351), .B(n410), .Z(n355) );
  NOR U436 ( .A(n355), .B(n412), .Z(n356) );
  NOR U437 ( .A(n357), .B(n356), .Z(n491) );
  NOR U438 ( .A(n671), .B(n358), .Z(n437) );
  IV U439 ( .A(n359), .Z(n362) );
  IV U440 ( .A(n360), .Z(n361) );
  NOR U441 ( .A(n362), .B(n361), .Z(n447) );
  NOR U442 ( .A(n669), .B(n363), .Z(n448) );
  NOR U443 ( .A(n554), .B(n444), .Z(n446) );
  XOR U444 ( .A(n448), .B(n446), .Z(n364) );
  XOR U445 ( .A(n447), .B(n364), .Z(n456) );
  NOR U446 ( .A(n366), .B(n365), .Z(n372) );
  NOR U447 ( .A(n368), .B(n367), .Z(n370) );
  NOR U448 ( .A(n370), .B(n369), .Z(n371) );
  NOR U449 ( .A(n372), .B(n371), .Z(n453) );
  IV U450 ( .A(n453), .Z(n454) );
  NOR U451 ( .A(n540), .B(n515), .Z(n455) );
  IV U452 ( .A(n455), .Z(n452) );
  XOR U453 ( .A(n454), .B(n452), .Z(n373) );
  XOR U454 ( .A(n456), .B(n373), .Z(n466) );
  NOR U455 ( .A(n584), .B(n534), .Z(n465) );
  IV U456 ( .A(n465), .Z(n462) );
  NOR U457 ( .A(n375), .B(n374), .Z(n381) );
  NOR U458 ( .A(n377), .B(n376), .Z(n379) );
  NOR U459 ( .A(n379), .B(n378), .Z(n380) );
  NOR U460 ( .A(n381), .B(n380), .Z(n463) );
  IV U461 ( .A(n463), .Z(n464) );
  XOR U462 ( .A(n462), .B(n464), .Z(n382) );
  XOR U463 ( .A(n466), .B(n382), .Z(n473) );
  NOR U464 ( .A(n543), .B(n604), .Z(n475) );
  IV U465 ( .A(n475), .Z(n471) );
  NOR U466 ( .A(n384), .B(n383), .Z(n390) );
  NOR U467 ( .A(n386), .B(n385), .Z(n388) );
  NOR U468 ( .A(n388), .B(n387), .Z(n389) );
  NOR U469 ( .A(n390), .B(n389), .Z(n472) );
  IV U470 ( .A(n472), .Z(n474) );
  XOR U471 ( .A(n471), .B(n474), .Z(n391) );
  XOR U472 ( .A(n473), .B(n391), .Z(n485) );
  NOR U473 ( .A(n393), .B(n392), .Z(n399) );
  NOR U474 ( .A(n395), .B(n394), .Z(n397) );
  NOR U475 ( .A(n397), .B(n396), .Z(n398) );
  NOR U476 ( .A(n399), .B(n398), .Z(n482) );
  IV U477 ( .A(n482), .Z(n483) );
  NOR U478 ( .A(n574), .B(n489), .Z(n484) );
  IV U479 ( .A(n484), .Z(n481) );
  XOR U480 ( .A(n483), .B(n481), .Z(n400) );
  XOR U481 ( .A(n485), .B(n400), .Z(n441) );
  IV U482 ( .A(n404), .Z(n403) );
  IV U483 ( .A(n401), .Z(n402) );
  NOR U484 ( .A(n403), .B(n402), .Z(n408) );
  NOR U485 ( .A(x[6]), .B(n404), .Z(n405) );
  NOR U486 ( .A(n406), .B(n405), .Z(n407) );
  NOR U487 ( .A(n408), .B(n407), .Z(n439) );
  XOR U488 ( .A(n441), .B(n439), .Z(n409) );
  XOR U489 ( .A(n437), .B(n409), .Z(n493) );
  XOR U490 ( .A(n491), .B(n493), .Z(n762) );
  IV U491 ( .A(n413), .Z(n414) );
  NOR U492 ( .A(x[6]), .B(n414), .Z(n415) );
  IV U493 ( .A(n415), .Z(n416) );
  NOR U494 ( .A(x[7]), .B(n416), .Z(n417) );
  IV U495 ( .A(n417), .Z(n763) );
  NOR U496 ( .A(x[6]), .B(n418), .Z(n422) );
  IV U497 ( .A(n418), .Z(n419) );
  NOR U498 ( .A(n574), .B(n419), .Z(n420) );
  NOR U499 ( .A(n420), .B(n554), .Z(n421) );
  NOR U500 ( .A(n422), .B(n421), .Z(n423) );
  NOR U501 ( .A(n423), .B(n669), .Z(n427) );
  IV U502 ( .A(n423), .Z(n424) );
  NOR U503 ( .A(y[7]), .B(n424), .Z(n425) );
  NOR U504 ( .A(x[7]), .B(n425), .Z(n426) );
  NOR U505 ( .A(n427), .B(n426), .Z(n765) );
  IV U506 ( .A(n738), .Z(n766) );
  IV U507 ( .A(n739), .Z(o[8]) );
  NOR U508 ( .A(n763), .B(c[0]), .Z(n428) );
  NOR U509 ( .A(n428), .B(n157), .Z(n431) );
  NOR U510 ( .A(n765), .B(n158), .Z(n429) );
  NOR U511 ( .A(c[1]), .B(n429), .Z(n430) );
  NOR U512 ( .A(n431), .B(n430), .Z(n432) );
  IV U513 ( .A(n432), .Z(n433) );
  NOR U514 ( .A(c[2]), .B(n433), .Z(n708) );
  NOR U515 ( .A(n746), .B(n434), .Z(n435) );
  IV U516 ( .A(n435), .Z(n706) );
  IV U517 ( .A(n439), .Z(n436) );
  NOR U518 ( .A(n437), .B(n436), .Z(n443) );
  IV U519 ( .A(n437), .Z(n438) );
  NOR U520 ( .A(n439), .B(n438), .Z(n440) );
  NOR U521 ( .A(n441), .B(n440), .Z(n442) );
  NOR U522 ( .A(n443), .B(n442), .Z(n636) );
  NOR U523 ( .A(n669), .B(n444), .Z(n445) );
  IV U524 ( .A(n445), .Z(n511) );
  NOR U525 ( .A(n554), .B(n515), .Z(n510) );
  IV U526 ( .A(n510), .Z(n508) );
  NOR U527 ( .A(n447), .B(n446), .Z(n450) );
  IV U528 ( .A(n448), .Z(n449) );
  NOR U529 ( .A(n450), .B(n449), .Z(n509) );
  IV U530 ( .A(n509), .Z(n507) );
  XOR U531 ( .A(n508), .B(n507), .Z(n451) );
  XOR U532 ( .A(n511), .B(n451), .Z(n501) );
  NOR U533 ( .A(n540), .B(n534), .Z(n500) );
  IV U534 ( .A(n500), .Z(n497) );
  NOR U535 ( .A(n453), .B(n452), .Z(n460) );
  NOR U536 ( .A(n455), .B(n454), .Z(n458) );
  IV U537 ( .A(n456), .Z(n457) );
  NOR U538 ( .A(n458), .B(n457), .Z(n459) );
  NOR U539 ( .A(n460), .B(n459), .Z(n498) );
  IV U540 ( .A(n498), .Z(n499) );
  XOR U541 ( .A(n497), .B(n499), .Z(n461) );
  XOR U542 ( .A(n501), .B(n461), .Z(n567) );
  NOR U543 ( .A(n543), .B(n584), .Z(n569) );
  IV U544 ( .A(n569), .Z(n565) );
  NOR U545 ( .A(n463), .B(n462), .Z(n469) );
  NOR U546 ( .A(n465), .B(n464), .Z(n467) );
  NOR U547 ( .A(n467), .B(n466), .Z(n468) );
  NOR U548 ( .A(n469), .B(n468), .Z(n566) );
  IV U549 ( .A(n566), .Z(n568) );
  XOR U550 ( .A(n565), .B(n568), .Z(n470) );
  XOR U551 ( .A(n567), .B(n470), .Z(n609) );
  NOR U552 ( .A(n574), .B(n604), .Z(n608) );
  IV U553 ( .A(n608), .Z(n605) );
  NOR U554 ( .A(n472), .B(n471), .Z(n479) );
  IV U555 ( .A(n473), .Z(n477) );
  NOR U556 ( .A(n475), .B(n474), .Z(n476) );
  NOR U557 ( .A(n477), .B(n476), .Z(n478) );
  NOR U558 ( .A(n479), .B(n478), .Z(n606) );
  IV U559 ( .A(n606), .Z(n607) );
  XOR U560 ( .A(n605), .B(n607), .Z(n480) );
  XOR U561 ( .A(n609), .B(n480), .Z(n631) );
  NOR U562 ( .A(n482), .B(n481), .Z(n488) );
  NOR U563 ( .A(n484), .B(n483), .Z(n486) );
  NOR U564 ( .A(n486), .B(n485), .Z(n487) );
  NOR U565 ( .A(n488), .B(n487), .Z(n630) );
  IV U566 ( .A(n630), .Z(n627) );
  NOR U567 ( .A(n671), .B(n489), .Z(n628) );
  IV U568 ( .A(n628), .Z(n629) );
  XOR U569 ( .A(n627), .B(n629), .Z(n490) );
  XOR U570 ( .A(n631), .B(n490), .Z(n638) );
  XOR U571 ( .A(n636), .B(n638), .Z(n641) );
  IV U572 ( .A(n491), .Z(n492) );
  NOR U573 ( .A(n493), .B(n492), .Z(n639) );
  XOR U574 ( .A(n641), .B(n639), .Z(n494) );
  NOR U575 ( .A(n706), .B(n494), .Z(n495) );
  NOR U576 ( .A(n708), .B(n495), .Z(n496) );
  IV U577 ( .A(n496), .Z(o[9]) );
  NOR U578 ( .A(n574), .B(n540), .Z(n521) );
  NOR U579 ( .A(n540), .B(n543), .Z(n505) );
  NOR U580 ( .A(n498), .B(n497), .Z(n504) );
  NOR U581 ( .A(n500), .B(n499), .Z(n502) );
  NOR U582 ( .A(n502), .B(n501), .Z(n503) );
  NOR U583 ( .A(n504), .B(n503), .Z(n506) );
  IV U584 ( .A(n506), .Z(n577) );
  NOR U585 ( .A(n505), .B(n577), .Z(n520) );
  IV U586 ( .A(n505), .Z(n578) );
  NOR U587 ( .A(n506), .B(n578), .Z(n518) );
  NOR U588 ( .A(n554), .B(n534), .Z(n525) );
  IV U589 ( .A(n525), .Z(n545) );
  NOR U590 ( .A(n508), .B(n507), .Z(n514) );
  NOR U591 ( .A(n510), .B(n509), .Z(n512) );
  NOR U592 ( .A(n512), .B(n511), .Z(n513) );
  NOR U593 ( .A(n514), .B(n513), .Z(n523) );
  IV U594 ( .A(n523), .Z(n524) );
  NOR U595 ( .A(n669), .B(n515), .Z(n516) );
  IV U596 ( .A(n516), .Z(n526) );
  XOR U597 ( .A(n524), .B(n526), .Z(n517) );
  XOR U598 ( .A(n545), .B(n517), .Z(n580) );
  NOR U599 ( .A(n518), .B(n580), .Z(n519) );
  NOR U600 ( .A(n520), .B(n519), .Z(n522) );
  NOR U601 ( .A(n521), .B(n522), .Z(n539) );
  IV U602 ( .A(n521), .Z(n588) );
  IV U603 ( .A(n522), .Z(n587) );
  NOR U604 ( .A(n588), .B(n587), .Z(n537) );
  NOR U605 ( .A(n523), .B(n545), .Z(n529) );
  NOR U606 ( .A(n525), .B(n524), .Z(n527) );
  NOR U607 ( .A(n527), .B(n526), .Z(n528) );
  NOR U608 ( .A(n529), .B(n528), .Z(n547) );
  NOR U609 ( .A(n547), .B(n543), .Z(n533) );
  IV U610 ( .A(n547), .Z(n531) );
  NOR U611 ( .A(n554), .B(n543), .Z(n530) );
  NOR U612 ( .A(n531), .B(n530), .Z(n532) );
  NOR U613 ( .A(n533), .B(n532), .Z(n536) );
  NOR U614 ( .A(n534), .B(n669), .Z(n535) );
  XOR U615 ( .A(n536), .B(n535), .Z(n590) );
  NOR U616 ( .A(n537), .B(n590), .Z(n538) );
  NOR U617 ( .A(n539), .B(n538), .Z(n541) );
  NOR U618 ( .A(n671), .B(n540), .Z(n542) );
  NOR U619 ( .A(n541), .B(n542), .Z(n553) );
  IV U620 ( .A(n541), .Z(n596) );
  IV U621 ( .A(n542), .Z(n595) );
  NOR U622 ( .A(n596), .B(n595), .Z(n551) );
  NOR U623 ( .A(n669), .B(n543), .Z(n544) );
  IV U624 ( .A(n544), .Z(n559) );
  NOR U625 ( .A(n545), .B(n559), .Z(n549) );
  NOR U626 ( .A(x[5]), .B(x[4]), .Z(n546) );
  NOR U627 ( .A(n547), .B(n546), .Z(n548) );
  NOR U628 ( .A(n549), .B(n548), .Z(n556) );
  IV U629 ( .A(n556), .Z(n557) );
  NOR U630 ( .A(n554), .B(n574), .Z(n558) );
  IV U631 ( .A(n558), .Z(n555) );
  XOR U632 ( .A(n557), .B(n555), .Z(n550) );
  XOR U633 ( .A(n559), .B(n550), .Z(n598) );
  NOR U634 ( .A(n551), .B(n598), .Z(n552) );
  NOR U635 ( .A(n553), .B(n552), .Z(n657) );
  IV U636 ( .A(n657), .Z(n564) );
  NOR U637 ( .A(n669), .B(n574), .Z(n664) );
  NOR U638 ( .A(n671), .B(n554), .Z(n663) );
  IV U639 ( .A(n663), .Z(n660) );
  NOR U640 ( .A(n556), .B(n555), .Z(n562) );
  NOR U641 ( .A(n558), .B(n557), .Z(n560) );
  NOR U642 ( .A(n560), .B(n559), .Z(n561) );
  NOR U643 ( .A(n562), .B(n561), .Z(n661) );
  IV U644 ( .A(n661), .Z(n662) );
  XOR U645 ( .A(n660), .B(n662), .Z(n563) );
  XOR U646 ( .A(n664), .B(n563), .Z(n656) );
  NOR U647 ( .A(n564), .B(n656), .Z(n659) );
  NOR U648 ( .A(n566), .B(n565), .Z(n573) );
  IV U649 ( .A(n567), .Z(n571) );
  NOR U650 ( .A(n569), .B(n568), .Z(n570) );
  NOR U651 ( .A(n571), .B(n570), .Z(n572) );
  NOR U652 ( .A(n573), .B(n572), .Z(n575) );
  NOR U653 ( .A(n574), .B(n584), .Z(n576) );
  IV U654 ( .A(n576), .Z(n616) );
  NOR U655 ( .A(n575), .B(n616), .Z(n583) );
  IV U656 ( .A(n575), .Z(n615) );
  NOR U657 ( .A(n576), .B(n615), .Z(n581) );
  XOR U658 ( .A(n578), .B(n577), .Z(n579) );
  XOR U659 ( .A(n580), .B(n579), .Z(n618) );
  NOR U660 ( .A(n581), .B(n618), .Z(n582) );
  NOR U661 ( .A(n583), .B(n582), .Z(n585) );
  NOR U662 ( .A(n671), .B(n584), .Z(n586) );
  IV U663 ( .A(n586), .Z(n601) );
  NOR U664 ( .A(n585), .B(n601), .Z(n594) );
  IV U665 ( .A(n585), .Z(n600) );
  NOR U666 ( .A(n586), .B(n600), .Z(n592) );
  XOR U667 ( .A(n588), .B(n587), .Z(n589) );
  XOR U668 ( .A(n590), .B(n589), .Z(n603) );
  IV U669 ( .A(n603), .Z(n591) );
  NOR U670 ( .A(n592), .B(n591), .Z(n593) );
  NOR U671 ( .A(n594), .B(n593), .Z(n653) );
  XOR U672 ( .A(n596), .B(n595), .Z(n597) );
  XOR U673 ( .A(n598), .B(n597), .Z(n652) );
  IV U674 ( .A(n652), .Z(n599) );
  NOR U675 ( .A(n653), .B(n599), .Z(n655) );
  XOR U676 ( .A(n601), .B(n600), .Z(n602) );
  XOR U677 ( .A(n603), .B(n602), .Z(n648) );
  NOR U678 ( .A(n671), .B(n604), .Z(n613) );
  NOR U679 ( .A(n606), .B(n605), .Z(n612) );
  NOR U680 ( .A(n608), .B(n607), .Z(n610) );
  NOR U681 ( .A(n610), .B(n609), .Z(n611) );
  NOR U682 ( .A(n612), .B(n611), .Z(n614) );
  IV U683 ( .A(n614), .Z(n623) );
  NOR U684 ( .A(n613), .B(n623), .Z(n621) );
  IV U685 ( .A(n613), .Z(n624) );
  NOR U686 ( .A(n614), .B(n624), .Z(n619) );
  XOR U687 ( .A(n616), .B(n615), .Z(n617) );
  XOR U688 ( .A(n618), .B(n617), .Z(n626) );
  NOR U689 ( .A(n619), .B(n626), .Z(n620) );
  NOR U690 ( .A(n621), .B(n620), .Z(n649) );
  IV U691 ( .A(n649), .Z(n622) );
  NOR U692 ( .A(n648), .B(n622), .Z(n651) );
  XOR U693 ( .A(n624), .B(n623), .Z(n625) );
  XOR U694 ( .A(n626), .B(n625), .Z(n644) );
  NOR U695 ( .A(n628), .B(n627), .Z(n634) );
  NOR U696 ( .A(n630), .B(n629), .Z(n632) );
  NOR U697 ( .A(n632), .B(n631), .Z(n633) );
  NOR U698 ( .A(n634), .B(n633), .Z(n645) );
  IV U699 ( .A(n645), .Z(n635) );
  NOR U700 ( .A(n644), .B(n635), .Z(n647) );
  IV U701 ( .A(n636), .Z(n637) );
  NOR U702 ( .A(n638), .B(n637), .Z(n643) );
  IV U703 ( .A(n639), .Z(n640) );
  NOR U704 ( .A(n641), .B(n640), .Z(n642) );
  NOR U705 ( .A(n643), .B(n642), .Z(n702) );
  XOR U706 ( .A(n645), .B(n644), .Z(n703) );
  NOR U707 ( .A(n702), .B(n703), .Z(n646) );
  NOR U708 ( .A(n647), .B(n646), .Z(n696) );
  XOR U709 ( .A(n649), .B(n648), .Z(n697) );
  NOR U710 ( .A(n696), .B(n697), .Z(n650) );
  NOR U711 ( .A(n651), .B(n650), .Z(n690) );
  XOR U712 ( .A(n653), .B(n652), .Z(n691) );
  NOR U713 ( .A(n690), .B(n691), .Z(n654) );
  NOR U714 ( .A(n655), .B(n654), .Z(n684) );
  XOR U715 ( .A(n657), .B(n656), .Z(n685) );
  NOR U716 ( .A(n684), .B(n685), .Z(n658) );
  NOR U717 ( .A(n659), .B(n658), .Z(n679) );
  NOR U718 ( .A(n661), .B(n660), .Z(n668) );
  NOR U719 ( .A(n663), .B(n662), .Z(n666) );
  IV U720 ( .A(n664), .Z(n665) );
  NOR U721 ( .A(n666), .B(n665), .Z(n667) );
  NOR U722 ( .A(n668), .B(n667), .Z(n672) );
  NOR U723 ( .A(n669), .B(n671), .Z(n670) );
  XOR U724 ( .A(n672), .B(n670), .Z(n678) );
  NOR U725 ( .A(n679), .B(n678), .Z(n674) );
  NOR U726 ( .A(n672), .B(n671), .Z(n673) );
  NOR U727 ( .A(n674), .B(n673), .Z(n675) );
  NOR U728 ( .A(n706), .B(n675), .Z(n676) );
  NOR U729 ( .A(n708), .B(n676), .Z(n677) );
  IV U730 ( .A(n677), .Z(o[15]) );
  XOR U731 ( .A(n679), .B(n678), .Z(n680) );
  IV U732 ( .A(n680), .Z(n681) );
  NOR U733 ( .A(n706), .B(n681), .Z(n682) );
  NOR U734 ( .A(n708), .B(n682), .Z(n683) );
  IV U735 ( .A(n683), .Z(o[14]) );
  IV U736 ( .A(n684), .Z(n686) );
  XOR U737 ( .A(n686), .B(n685), .Z(n687) );
  NOR U738 ( .A(n706), .B(n687), .Z(n688) );
  NOR U739 ( .A(n708), .B(n688), .Z(n689) );
  IV U740 ( .A(n689), .Z(o[13]) );
  IV U741 ( .A(n690), .Z(n692) );
  XOR U742 ( .A(n692), .B(n691), .Z(n693) );
  NOR U743 ( .A(n706), .B(n693), .Z(n694) );
  NOR U744 ( .A(n708), .B(n694), .Z(n695) );
  IV U745 ( .A(n695), .Z(o[12]) );
  IV U746 ( .A(n696), .Z(n698) );
  XOR U747 ( .A(n698), .B(n697), .Z(n699) );
  NOR U748 ( .A(n706), .B(n699), .Z(n700) );
  NOR U749 ( .A(n708), .B(n700), .Z(n701) );
  IV U750 ( .A(n701), .Z(o[11]) );
  IV U751 ( .A(n702), .Z(n704) );
  XOR U752 ( .A(n704), .B(n703), .Z(n705) );
  NOR U753 ( .A(n706), .B(n705), .Z(n707) );
  NOR U754 ( .A(n708), .B(n707), .Z(n709) );
  IV U755 ( .A(n709), .Z(o[10]) );
  NOR U756 ( .A(c[2]), .B(n157), .Z(n710) );
  NOR U757 ( .A(c[2]), .B(c[1]), .Z(n711) );
  NOR U758 ( .A(n158), .B(n741), .Z(n712) );
  NOR U759 ( .A(c[0]), .B(n742), .Z(n713) );
  NOR U760 ( .A(n712), .B(n713), .Z(n714) );
  NOR U761 ( .A(c[0]), .B(c[2]), .Z(n715) );
  NOR U762 ( .A(n157), .B(n743), .Z(n716) );
  NOR U763 ( .A(c[0]), .B(c[1]), .Z(n717) );
  NOR U764 ( .A(n746), .B(n740), .Z(n718) );
  NOR U765 ( .A(n158), .B(n742), .Z(n719) );
  NOR U766 ( .A(n744), .B(x[0]), .Z(n720) );
  NOR U767 ( .A(n747), .B(n748), .Z(n721) );
  NOR U768 ( .A(n745), .B(n750), .Z(n722) );
  NOR U769 ( .A(n721), .B(n722), .Z(n723) );
  NOR U770 ( .A(n749), .B(n751), .Z(n724) );
  NOR U771 ( .A(n744), .B(n753), .Z(n725) );
  NOR U772 ( .A(n747), .B(n752), .Z(n726) );
  NOR U773 ( .A(n745), .B(n755), .Z(n727) );
  NOR U774 ( .A(n726), .B(n727), .Z(n728) );
  NOR U775 ( .A(n754), .B(n756), .Z(n729) );
  NOR U776 ( .A(n744), .B(n758), .Z(n730) );
  NOR U777 ( .A(n747), .B(n757), .Z(n731) );
  NOR U778 ( .A(n745), .B(n760), .Z(n732) );
  NOR U779 ( .A(n731), .B(n732), .Z(n733) );
  NOR U780 ( .A(n759), .B(n761), .Z(n734) );
  NOR U781 ( .A(n744), .B(n763), .Z(n735) );
  NOR U782 ( .A(n747), .B(n762), .Z(n736) );
  NOR U783 ( .A(n745), .B(n765), .Z(n737) );
  NOR U784 ( .A(n736), .B(n737), .Z(n738) );
  NOR U785 ( .A(n764), .B(n766), .Z(n739) );
endmodule

