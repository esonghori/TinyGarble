
module MUX_N256_3 ( A, B, S, O );
  input [255:0] A;
  input [255:0] B;
  output [255:0] O;
  input S;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512;

  XOR U1 ( .A(A[9]), .B(n1), .Z(O[9]) );
  AND U2 ( .A(S), .B(n2), .Z(n1) );
  XOR U3 ( .A(B[9]), .B(A[9]), .Z(n2) );
  XOR U4 ( .A(A[99]), .B(n3), .Z(O[99]) );
  AND U5 ( .A(S), .B(n4), .Z(n3) );
  XOR U6 ( .A(B[99]), .B(A[99]), .Z(n4) );
  XOR U7 ( .A(A[98]), .B(n5), .Z(O[98]) );
  AND U8 ( .A(S), .B(n6), .Z(n5) );
  XOR U9 ( .A(B[98]), .B(A[98]), .Z(n6) );
  XOR U10 ( .A(A[97]), .B(n7), .Z(O[97]) );
  AND U11 ( .A(S), .B(n8), .Z(n7) );
  XOR U12 ( .A(B[97]), .B(A[97]), .Z(n8) );
  XOR U13 ( .A(A[96]), .B(n9), .Z(O[96]) );
  AND U14 ( .A(S), .B(n10), .Z(n9) );
  XOR U15 ( .A(B[96]), .B(A[96]), .Z(n10) );
  XOR U16 ( .A(A[95]), .B(n11), .Z(O[95]) );
  AND U17 ( .A(S), .B(n12), .Z(n11) );
  XOR U18 ( .A(B[95]), .B(A[95]), .Z(n12) );
  XOR U19 ( .A(A[94]), .B(n13), .Z(O[94]) );
  AND U20 ( .A(S), .B(n14), .Z(n13) );
  XOR U21 ( .A(B[94]), .B(A[94]), .Z(n14) );
  XOR U22 ( .A(A[93]), .B(n15), .Z(O[93]) );
  AND U23 ( .A(S), .B(n16), .Z(n15) );
  XOR U24 ( .A(B[93]), .B(A[93]), .Z(n16) );
  XOR U25 ( .A(A[92]), .B(n17), .Z(O[92]) );
  AND U26 ( .A(S), .B(n18), .Z(n17) );
  XOR U27 ( .A(B[92]), .B(A[92]), .Z(n18) );
  XOR U28 ( .A(A[91]), .B(n19), .Z(O[91]) );
  AND U29 ( .A(S), .B(n20), .Z(n19) );
  XOR U30 ( .A(B[91]), .B(A[91]), .Z(n20) );
  XOR U31 ( .A(A[90]), .B(n21), .Z(O[90]) );
  AND U32 ( .A(S), .B(n22), .Z(n21) );
  XOR U33 ( .A(B[90]), .B(A[90]), .Z(n22) );
  XOR U34 ( .A(A[8]), .B(n23), .Z(O[8]) );
  AND U35 ( .A(S), .B(n24), .Z(n23) );
  XOR U36 ( .A(B[8]), .B(A[8]), .Z(n24) );
  XOR U37 ( .A(A[89]), .B(n25), .Z(O[89]) );
  AND U38 ( .A(S), .B(n26), .Z(n25) );
  XOR U39 ( .A(B[89]), .B(A[89]), .Z(n26) );
  XOR U40 ( .A(A[88]), .B(n27), .Z(O[88]) );
  AND U41 ( .A(S), .B(n28), .Z(n27) );
  XOR U42 ( .A(B[88]), .B(A[88]), .Z(n28) );
  XOR U43 ( .A(A[87]), .B(n29), .Z(O[87]) );
  AND U44 ( .A(S), .B(n30), .Z(n29) );
  XOR U45 ( .A(B[87]), .B(A[87]), .Z(n30) );
  XOR U46 ( .A(A[86]), .B(n31), .Z(O[86]) );
  AND U47 ( .A(S), .B(n32), .Z(n31) );
  XOR U48 ( .A(B[86]), .B(A[86]), .Z(n32) );
  XOR U49 ( .A(A[85]), .B(n33), .Z(O[85]) );
  AND U50 ( .A(S), .B(n34), .Z(n33) );
  XOR U51 ( .A(B[85]), .B(A[85]), .Z(n34) );
  XOR U52 ( .A(A[84]), .B(n35), .Z(O[84]) );
  AND U53 ( .A(S), .B(n36), .Z(n35) );
  XOR U54 ( .A(B[84]), .B(A[84]), .Z(n36) );
  XOR U55 ( .A(A[83]), .B(n37), .Z(O[83]) );
  AND U56 ( .A(S), .B(n38), .Z(n37) );
  XOR U57 ( .A(B[83]), .B(A[83]), .Z(n38) );
  XOR U58 ( .A(A[82]), .B(n39), .Z(O[82]) );
  AND U59 ( .A(S), .B(n40), .Z(n39) );
  XOR U60 ( .A(B[82]), .B(A[82]), .Z(n40) );
  XOR U61 ( .A(A[81]), .B(n41), .Z(O[81]) );
  AND U62 ( .A(S), .B(n42), .Z(n41) );
  XOR U63 ( .A(B[81]), .B(A[81]), .Z(n42) );
  XOR U64 ( .A(A[80]), .B(n43), .Z(O[80]) );
  AND U65 ( .A(S), .B(n44), .Z(n43) );
  XOR U66 ( .A(B[80]), .B(A[80]), .Z(n44) );
  XOR U67 ( .A(A[7]), .B(n45), .Z(O[7]) );
  AND U68 ( .A(S), .B(n46), .Z(n45) );
  XOR U69 ( .A(B[7]), .B(A[7]), .Z(n46) );
  XOR U70 ( .A(A[79]), .B(n47), .Z(O[79]) );
  AND U71 ( .A(S), .B(n48), .Z(n47) );
  XOR U72 ( .A(B[79]), .B(A[79]), .Z(n48) );
  XOR U73 ( .A(A[78]), .B(n49), .Z(O[78]) );
  AND U74 ( .A(S), .B(n50), .Z(n49) );
  XOR U75 ( .A(B[78]), .B(A[78]), .Z(n50) );
  XOR U76 ( .A(A[77]), .B(n51), .Z(O[77]) );
  AND U77 ( .A(S), .B(n52), .Z(n51) );
  XOR U78 ( .A(B[77]), .B(A[77]), .Z(n52) );
  XOR U79 ( .A(A[76]), .B(n53), .Z(O[76]) );
  AND U80 ( .A(S), .B(n54), .Z(n53) );
  XOR U81 ( .A(B[76]), .B(A[76]), .Z(n54) );
  XOR U82 ( .A(A[75]), .B(n55), .Z(O[75]) );
  AND U83 ( .A(S), .B(n56), .Z(n55) );
  XOR U84 ( .A(B[75]), .B(A[75]), .Z(n56) );
  XOR U85 ( .A(A[74]), .B(n57), .Z(O[74]) );
  AND U86 ( .A(S), .B(n58), .Z(n57) );
  XOR U87 ( .A(B[74]), .B(A[74]), .Z(n58) );
  XOR U88 ( .A(A[73]), .B(n59), .Z(O[73]) );
  AND U89 ( .A(S), .B(n60), .Z(n59) );
  XOR U90 ( .A(B[73]), .B(A[73]), .Z(n60) );
  XOR U91 ( .A(A[72]), .B(n61), .Z(O[72]) );
  AND U92 ( .A(S), .B(n62), .Z(n61) );
  XOR U93 ( .A(B[72]), .B(A[72]), .Z(n62) );
  XOR U94 ( .A(A[71]), .B(n63), .Z(O[71]) );
  AND U95 ( .A(S), .B(n64), .Z(n63) );
  XOR U96 ( .A(B[71]), .B(A[71]), .Z(n64) );
  XOR U97 ( .A(A[70]), .B(n65), .Z(O[70]) );
  AND U98 ( .A(S), .B(n66), .Z(n65) );
  XOR U99 ( .A(B[70]), .B(A[70]), .Z(n66) );
  XOR U100 ( .A(A[6]), .B(n67), .Z(O[6]) );
  AND U101 ( .A(S), .B(n68), .Z(n67) );
  XOR U102 ( .A(B[6]), .B(A[6]), .Z(n68) );
  XOR U103 ( .A(A[69]), .B(n69), .Z(O[69]) );
  AND U104 ( .A(S), .B(n70), .Z(n69) );
  XOR U105 ( .A(B[69]), .B(A[69]), .Z(n70) );
  XOR U106 ( .A(A[68]), .B(n71), .Z(O[68]) );
  AND U107 ( .A(S), .B(n72), .Z(n71) );
  XOR U108 ( .A(B[68]), .B(A[68]), .Z(n72) );
  XOR U109 ( .A(A[67]), .B(n73), .Z(O[67]) );
  AND U110 ( .A(S), .B(n74), .Z(n73) );
  XOR U111 ( .A(B[67]), .B(A[67]), .Z(n74) );
  XOR U112 ( .A(A[66]), .B(n75), .Z(O[66]) );
  AND U113 ( .A(S), .B(n76), .Z(n75) );
  XOR U114 ( .A(B[66]), .B(A[66]), .Z(n76) );
  XOR U115 ( .A(A[65]), .B(n77), .Z(O[65]) );
  AND U116 ( .A(S), .B(n78), .Z(n77) );
  XOR U117 ( .A(B[65]), .B(A[65]), .Z(n78) );
  XOR U118 ( .A(A[64]), .B(n79), .Z(O[64]) );
  AND U119 ( .A(S), .B(n80), .Z(n79) );
  XOR U120 ( .A(B[64]), .B(A[64]), .Z(n80) );
  XOR U121 ( .A(A[63]), .B(n81), .Z(O[63]) );
  AND U122 ( .A(S), .B(n82), .Z(n81) );
  XOR U123 ( .A(B[63]), .B(A[63]), .Z(n82) );
  XOR U124 ( .A(A[62]), .B(n83), .Z(O[62]) );
  AND U125 ( .A(S), .B(n84), .Z(n83) );
  XOR U126 ( .A(B[62]), .B(A[62]), .Z(n84) );
  XOR U127 ( .A(A[61]), .B(n85), .Z(O[61]) );
  AND U128 ( .A(S), .B(n86), .Z(n85) );
  XOR U129 ( .A(B[61]), .B(A[61]), .Z(n86) );
  XOR U130 ( .A(A[60]), .B(n87), .Z(O[60]) );
  AND U131 ( .A(S), .B(n88), .Z(n87) );
  XOR U132 ( .A(B[60]), .B(A[60]), .Z(n88) );
  XOR U133 ( .A(A[5]), .B(n89), .Z(O[5]) );
  AND U134 ( .A(S), .B(n90), .Z(n89) );
  XOR U135 ( .A(B[5]), .B(A[5]), .Z(n90) );
  XOR U136 ( .A(A[59]), .B(n91), .Z(O[59]) );
  AND U137 ( .A(S), .B(n92), .Z(n91) );
  XOR U138 ( .A(B[59]), .B(A[59]), .Z(n92) );
  XOR U139 ( .A(A[58]), .B(n93), .Z(O[58]) );
  AND U140 ( .A(S), .B(n94), .Z(n93) );
  XOR U141 ( .A(B[58]), .B(A[58]), .Z(n94) );
  XOR U142 ( .A(A[57]), .B(n95), .Z(O[57]) );
  AND U143 ( .A(S), .B(n96), .Z(n95) );
  XOR U144 ( .A(B[57]), .B(A[57]), .Z(n96) );
  XOR U145 ( .A(A[56]), .B(n97), .Z(O[56]) );
  AND U146 ( .A(S), .B(n98), .Z(n97) );
  XOR U147 ( .A(B[56]), .B(A[56]), .Z(n98) );
  XOR U148 ( .A(A[55]), .B(n99), .Z(O[55]) );
  AND U149 ( .A(S), .B(n100), .Z(n99) );
  XOR U150 ( .A(B[55]), .B(A[55]), .Z(n100) );
  XOR U151 ( .A(A[54]), .B(n101), .Z(O[54]) );
  AND U152 ( .A(S), .B(n102), .Z(n101) );
  XOR U153 ( .A(B[54]), .B(A[54]), .Z(n102) );
  XOR U154 ( .A(A[53]), .B(n103), .Z(O[53]) );
  AND U155 ( .A(S), .B(n104), .Z(n103) );
  XOR U156 ( .A(B[53]), .B(A[53]), .Z(n104) );
  XOR U157 ( .A(A[52]), .B(n105), .Z(O[52]) );
  AND U158 ( .A(S), .B(n106), .Z(n105) );
  XOR U159 ( .A(B[52]), .B(A[52]), .Z(n106) );
  XOR U160 ( .A(A[51]), .B(n107), .Z(O[51]) );
  AND U161 ( .A(S), .B(n108), .Z(n107) );
  XOR U162 ( .A(B[51]), .B(A[51]), .Z(n108) );
  XOR U163 ( .A(A[50]), .B(n109), .Z(O[50]) );
  AND U164 ( .A(S), .B(n110), .Z(n109) );
  XOR U165 ( .A(B[50]), .B(A[50]), .Z(n110) );
  XOR U166 ( .A(A[4]), .B(n111), .Z(O[4]) );
  AND U167 ( .A(S), .B(n112), .Z(n111) );
  XOR U168 ( .A(B[4]), .B(A[4]), .Z(n112) );
  XOR U169 ( .A(A[49]), .B(n113), .Z(O[49]) );
  AND U170 ( .A(S), .B(n114), .Z(n113) );
  XOR U171 ( .A(B[49]), .B(A[49]), .Z(n114) );
  XOR U172 ( .A(A[48]), .B(n115), .Z(O[48]) );
  AND U173 ( .A(S), .B(n116), .Z(n115) );
  XOR U174 ( .A(B[48]), .B(A[48]), .Z(n116) );
  XOR U175 ( .A(A[47]), .B(n117), .Z(O[47]) );
  AND U176 ( .A(S), .B(n118), .Z(n117) );
  XOR U177 ( .A(B[47]), .B(A[47]), .Z(n118) );
  XOR U178 ( .A(A[46]), .B(n119), .Z(O[46]) );
  AND U179 ( .A(S), .B(n120), .Z(n119) );
  XOR U180 ( .A(B[46]), .B(A[46]), .Z(n120) );
  XOR U181 ( .A(A[45]), .B(n121), .Z(O[45]) );
  AND U182 ( .A(S), .B(n122), .Z(n121) );
  XOR U183 ( .A(B[45]), .B(A[45]), .Z(n122) );
  XOR U184 ( .A(A[44]), .B(n123), .Z(O[44]) );
  AND U185 ( .A(S), .B(n124), .Z(n123) );
  XOR U186 ( .A(B[44]), .B(A[44]), .Z(n124) );
  XOR U187 ( .A(A[43]), .B(n125), .Z(O[43]) );
  AND U188 ( .A(S), .B(n126), .Z(n125) );
  XOR U189 ( .A(B[43]), .B(A[43]), .Z(n126) );
  XOR U190 ( .A(A[42]), .B(n127), .Z(O[42]) );
  AND U191 ( .A(S), .B(n128), .Z(n127) );
  XOR U192 ( .A(B[42]), .B(A[42]), .Z(n128) );
  XOR U193 ( .A(A[41]), .B(n129), .Z(O[41]) );
  AND U194 ( .A(S), .B(n130), .Z(n129) );
  XOR U195 ( .A(B[41]), .B(A[41]), .Z(n130) );
  XOR U196 ( .A(A[40]), .B(n131), .Z(O[40]) );
  AND U197 ( .A(S), .B(n132), .Z(n131) );
  XOR U198 ( .A(B[40]), .B(A[40]), .Z(n132) );
  XOR U199 ( .A(A[3]), .B(n133), .Z(O[3]) );
  AND U200 ( .A(S), .B(n134), .Z(n133) );
  XOR U201 ( .A(B[3]), .B(A[3]), .Z(n134) );
  XOR U202 ( .A(A[39]), .B(n135), .Z(O[39]) );
  AND U203 ( .A(S), .B(n136), .Z(n135) );
  XOR U204 ( .A(B[39]), .B(A[39]), .Z(n136) );
  XOR U205 ( .A(A[38]), .B(n137), .Z(O[38]) );
  AND U206 ( .A(S), .B(n138), .Z(n137) );
  XOR U207 ( .A(B[38]), .B(A[38]), .Z(n138) );
  XOR U208 ( .A(A[37]), .B(n139), .Z(O[37]) );
  AND U209 ( .A(S), .B(n140), .Z(n139) );
  XOR U210 ( .A(B[37]), .B(A[37]), .Z(n140) );
  XOR U211 ( .A(A[36]), .B(n141), .Z(O[36]) );
  AND U212 ( .A(S), .B(n142), .Z(n141) );
  XOR U213 ( .A(B[36]), .B(A[36]), .Z(n142) );
  XOR U214 ( .A(A[35]), .B(n143), .Z(O[35]) );
  AND U215 ( .A(S), .B(n144), .Z(n143) );
  XOR U216 ( .A(B[35]), .B(A[35]), .Z(n144) );
  XOR U217 ( .A(A[34]), .B(n145), .Z(O[34]) );
  AND U218 ( .A(S), .B(n146), .Z(n145) );
  XOR U219 ( .A(B[34]), .B(A[34]), .Z(n146) );
  XOR U220 ( .A(A[33]), .B(n147), .Z(O[33]) );
  AND U221 ( .A(S), .B(n148), .Z(n147) );
  XOR U222 ( .A(B[33]), .B(A[33]), .Z(n148) );
  XOR U223 ( .A(A[32]), .B(n149), .Z(O[32]) );
  AND U224 ( .A(S), .B(n150), .Z(n149) );
  XOR U225 ( .A(B[32]), .B(A[32]), .Z(n150) );
  XOR U226 ( .A(A[31]), .B(n151), .Z(O[31]) );
  AND U227 ( .A(S), .B(n152), .Z(n151) );
  XOR U228 ( .A(B[31]), .B(A[31]), .Z(n152) );
  XOR U229 ( .A(A[30]), .B(n153), .Z(O[30]) );
  AND U230 ( .A(S), .B(n154), .Z(n153) );
  XOR U231 ( .A(B[30]), .B(A[30]), .Z(n154) );
  XOR U232 ( .A(A[2]), .B(n155), .Z(O[2]) );
  AND U233 ( .A(S), .B(n156), .Z(n155) );
  XOR U234 ( .A(B[2]), .B(A[2]), .Z(n156) );
  XOR U235 ( .A(A[29]), .B(n157), .Z(O[29]) );
  AND U236 ( .A(S), .B(n158), .Z(n157) );
  XOR U237 ( .A(B[29]), .B(A[29]), .Z(n158) );
  XOR U238 ( .A(A[28]), .B(n159), .Z(O[28]) );
  AND U239 ( .A(S), .B(n160), .Z(n159) );
  XOR U240 ( .A(B[28]), .B(A[28]), .Z(n160) );
  XOR U241 ( .A(A[27]), .B(n161), .Z(O[27]) );
  AND U242 ( .A(S), .B(n162), .Z(n161) );
  XOR U243 ( .A(B[27]), .B(A[27]), .Z(n162) );
  XOR U244 ( .A(A[26]), .B(n163), .Z(O[26]) );
  AND U245 ( .A(S), .B(n164), .Z(n163) );
  XOR U246 ( .A(B[26]), .B(A[26]), .Z(n164) );
  XOR U247 ( .A(A[25]), .B(n165), .Z(O[25]) );
  AND U248 ( .A(S), .B(n166), .Z(n165) );
  XOR U249 ( .A(B[25]), .B(A[25]), .Z(n166) );
  XOR U250 ( .A(A[255]), .B(n167), .Z(O[255]) );
  AND U251 ( .A(S), .B(n168), .Z(n167) );
  XOR U252 ( .A(B[255]), .B(A[255]), .Z(n168) );
  XOR U253 ( .A(A[254]), .B(n169), .Z(O[254]) );
  AND U254 ( .A(S), .B(n170), .Z(n169) );
  XOR U255 ( .A(B[254]), .B(A[254]), .Z(n170) );
  XOR U256 ( .A(A[253]), .B(n171), .Z(O[253]) );
  AND U257 ( .A(S), .B(n172), .Z(n171) );
  XOR U258 ( .A(B[253]), .B(A[253]), .Z(n172) );
  XOR U259 ( .A(A[252]), .B(n173), .Z(O[252]) );
  AND U260 ( .A(S), .B(n174), .Z(n173) );
  XOR U261 ( .A(B[252]), .B(A[252]), .Z(n174) );
  XOR U262 ( .A(A[251]), .B(n175), .Z(O[251]) );
  AND U263 ( .A(S), .B(n176), .Z(n175) );
  XOR U264 ( .A(B[251]), .B(A[251]), .Z(n176) );
  XOR U265 ( .A(A[250]), .B(n177), .Z(O[250]) );
  AND U266 ( .A(S), .B(n178), .Z(n177) );
  XOR U267 ( .A(B[250]), .B(A[250]), .Z(n178) );
  XOR U268 ( .A(A[24]), .B(n179), .Z(O[24]) );
  AND U269 ( .A(S), .B(n180), .Z(n179) );
  XOR U270 ( .A(B[24]), .B(A[24]), .Z(n180) );
  XOR U271 ( .A(A[249]), .B(n181), .Z(O[249]) );
  AND U272 ( .A(S), .B(n182), .Z(n181) );
  XOR U273 ( .A(B[249]), .B(A[249]), .Z(n182) );
  XOR U274 ( .A(A[248]), .B(n183), .Z(O[248]) );
  AND U275 ( .A(S), .B(n184), .Z(n183) );
  XOR U276 ( .A(B[248]), .B(A[248]), .Z(n184) );
  XOR U277 ( .A(A[247]), .B(n185), .Z(O[247]) );
  AND U278 ( .A(S), .B(n186), .Z(n185) );
  XOR U279 ( .A(B[247]), .B(A[247]), .Z(n186) );
  XOR U280 ( .A(A[246]), .B(n187), .Z(O[246]) );
  AND U281 ( .A(S), .B(n188), .Z(n187) );
  XOR U282 ( .A(B[246]), .B(A[246]), .Z(n188) );
  XOR U283 ( .A(A[245]), .B(n189), .Z(O[245]) );
  AND U284 ( .A(S), .B(n190), .Z(n189) );
  XOR U285 ( .A(B[245]), .B(A[245]), .Z(n190) );
  XOR U286 ( .A(A[244]), .B(n191), .Z(O[244]) );
  AND U287 ( .A(S), .B(n192), .Z(n191) );
  XOR U288 ( .A(B[244]), .B(A[244]), .Z(n192) );
  XOR U289 ( .A(A[243]), .B(n193), .Z(O[243]) );
  AND U290 ( .A(S), .B(n194), .Z(n193) );
  XOR U291 ( .A(B[243]), .B(A[243]), .Z(n194) );
  XOR U292 ( .A(A[242]), .B(n195), .Z(O[242]) );
  AND U293 ( .A(S), .B(n196), .Z(n195) );
  XOR U294 ( .A(B[242]), .B(A[242]), .Z(n196) );
  XOR U295 ( .A(A[241]), .B(n197), .Z(O[241]) );
  AND U296 ( .A(S), .B(n198), .Z(n197) );
  XOR U297 ( .A(B[241]), .B(A[241]), .Z(n198) );
  XOR U298 ( .A(A[240]), .B(n199), .Z(O[240]) );
  AND U299 ( .A(S), .B(n200), .Z(n199) );
  XOR U300 ( .A(B[240]), .B(A[240]), .Z(n200) );
  XOR U301 ( .A(A[23]), .B(n201), .Z(O[23]) );
  AND U302 ( .A(S), .B(n202), .Z(n201) );
  XOR U303 ( .A(B[23]), .B(A[23]), .Z(n202) );
  XOR U304 ( .A(A[239]), .B(n203), .Z(O[239]) );
  AND U305 ( .A(S), .B(n204), .Z(n203) );
  XOR U306 ( .A(B[239]), .B(A[239]), .Z(n204) );
  XOR U307 ( .A(A[238]), .B(n205), .Z(O[238]) );
  AND U308 ( .A(S), .B(n206), .Z(n205) );
  XOR U309 ( .A(B[238]), .B(A[238]), .Z(n206) );
  XOR U310 ( .A(A[237]), .B(n207), .Z(O[237]) );
  AND U311 ( .A(S), .B(n208), .Z(n207) );
  XOR U312 ( .A(B[237]), .B(A[237]), .Z(n208) );
  XOR U313 ( .A(A[236]), .B(n209), .Z(O[236]) );
  AND U314 ( .A(S), .B(n210), .Z(n209) );
  XOR U315 ( .A(B[236]), .B(A[236]), .Z(n210) );
  XOR U316 ( .A(A[235]), .B(n211), .Z(O[235]) );
  AND U317 ( .A(S), .B(n212), .Z(n211) );
  XOR U318 ( .A(B[235]), .B(A[235]), .Z(n212) );
  XOR U319 ( .A(A[234]), .B(n213), .Z(O[234]) );
  AND U320 ( .A(S), .B(n214), .Z(n213) );
  XOR U321 ( .A(B[234]), .B(A[234]), .Z(n214) );
  XOR U322 ( .A(A[233]), .B(n215), .Z(O[233]) );
  AND U323 ( .A(S), .B(n216), .Z(n215) );
  XOR U324 ( .A(B[233]), .B(A[233]), .Z(n216) );
  XOR U325 ( .A(A[232]), .B(n217), .Z(O[232]) );
  AND U326 ( .A(S), .B(n218), .Z(n217) );
  XOR U327 ( .A(B[232]), .B(A[232]), .Z(n218) );
  XOR U328 ( .A(A[231]), .B(n219), .Z(O[231]) );
  AND U329 ( .A(S), .B(n220), .Z(n219) );
  XOR U330 ( .A(B[231]), .B(A[231]), .Z(n220) );
  XOR U331 ( .A(A[230]), .B(n221), .Z(O[230]) );
  AND U332 ( .A(S), .B(n222), .Z(n221) );
  XOR U333 ( .A(B[230]), .B(A[230]), .Z(n222) );
  XOR U334 ( .A(A[22]), .B(n223), .Z(O[22]) );
  AND U335 ( .A(S), .B(n224), .Z(n223) );
  XOR U336 ( .A(B[22]), .B(A[22]), .Z(n224) );
  XOR U337 ( .A(A[229]), .B(n225), .Z(O[229]) );
  AND U338 ( .A(S), .B(n226), .Z(n225) );
  XOR U339 ( .A(B[229]), .B(A[229]), .Z(n226) );
  XOR U340 ( .A(A[228]), .B(n227), .Z(O[228]) );
  AND U341 ( .A(S), .B(n228), .Z(n227) );
  XOR U342 ( .A(B[228]), .B(A[228]), .Z(n228) );
  XOR U343 ( .A(A[227]), .B(n229), .Z(O[227]) );
  AND U344 ( .A(S), .B(n230), .Z(n229) );
  XOR U345 ( .A(B[227]), .B(A[227]), .Z(n230) );
  XOR U346 ( .A(A[226]), .B(n231), .Z(O[226]) );
  AND U347 ( .A(S), .B(n232), .Z(n231) );
  XOR U348 ( .A(B[226]), .B(A[226]), .Z(n232) );
  XOR U349 ( .A(A[225]), .B(n233), .Z(O[225]) );
  AND U350 ( .A(S), .B(n234), .Z(n233) );
  XOR U351 ( .A(B[225]), .B(A[225]), .Z(n234) );
  XOR U352 ( .A(A[224]), .B(n235), .Z(O[224]) );
  AND U353 ( .A(S), .B(n236), .Z(n235) );
  XOR U354 ( .A(B[224]), .B(A[224]), .Z(n236) );
  XOR U355 ( .A(A[223]), .B(n237), .Z(O[223]) );
  AND U356 ( .A(S), .B(n238), .Z(n237) );
  XOR U357 ( .A(B[223]), .B(A[223]), .Z(n238) );
  XOR U358 ( .A(A[222]), .B(n239), .Z(O[222]) );
  AND U359 ( .A(S), .B(n240), .Z(n239) );
  XOR U360 ( .A(B[222]), .B(A[222]), .Z(n240) );
  XOR U361 ( .A(A[221]), .B(n241), .Z(O[221]) );
  AND U362 ( .A(S), .B(n242), .Z(n241) );
  XOR U363 ( .A(B[221]), .B(A[221]), .Z(n242) );
  XOR U364 ( .A(A[220]), .B(n243), .Z(O[220]) );
  AND U365 ( .A(S), .B(n244), .Z(n243) );
  XOR U366 ( .A(B[220]), .B(A[220]), .Z(n244) );
  XOR U367 ( .A(A[21]), .B(n245), .Z(O[21]) );
  AND U368 ( .A(S), .B(n246), .Z(n245) );
  XOR U369 ( .A(B[21]), .B(A[21]), .Z(n246) );
  XOR U370 ( .A(A[219]), .B(n247), .Z(O[219]) );
  AND U371 ( .A(S), .B(n248), .Z(n247) );
  XOR U372 ( .A(B[219]), .B(A[219]), .Z(n248) );
  XOR U373 ( .A(A[218]), .B(n249), .Z(O[218]) );
  AND U374 ( .A(S), .B(n250), .Z(n249) );
  XOR U375 ( .A(B[218]), .B(A[218]), .Z(n250) );
  XOR U376 ( .A(A[217]), .B(n251), .Z(O[217]) );
  AND U377 ( .A(S), .B(n252), .Z(n251) );
  XOR U378 ( .A(B[217]), .B(A[217]), .Z(n252) );
  XOR U379 ( .A(A[216]), .B(n253), .Z(O[216]) );
  AND U380 ( .A(S), .B(n254), .Z(n253) );
  XOR U381 ( .A(B[216]), .B(A[216]), .Z(n254) );
  XOR U382 ( .A(A[215]), .B(n255), .Z(O[215]) );
  AND U383 ( .A(S), .B(n256), .Z(n255) );
  XOR U384 ( .A(B[215]), .B(A[215]), .Z(n256) );
  XOR U385 ( .A(A[214]), .B(n257), .Z(O[214]) );
  AND U386 ( .A(S), .B(n258), .Z(n257) );
  XOR U387 ( .A(B[214]), .B(A[214]), .Z(n258) );
  XOR U388 ( .A(A[213]), .B(n259), .Z(O[213]) );
  AND U389 ( .A(S), .B(n260), .Z(n259) );
  XOR U390 ( .A(B[213]), .B(A[213]), .Z(n260) );
  XOR U391 ( .A(A[212]), .B(n261), .Z(O[212]) );
  AND U392 ( .A(S), .B(n262), .Z(n261) );
  XOR U393 ( .A(B[212]), .B(A[212]), .Z(n262) );
  XOR U394 ( .A(A[211]), .B(n263), .Z(O[211]) );
  AND U395 ( .A(S), .B(n264), .Z(n263) );
  XOR U396 ( .A(B[211]), .B(A[211]), .Z(n264) );
  XOR U397 ( .A(A[210]), .B(n265), .Z(O[210]) );
  AND U398 ( .A(S), .B(n266), .Z(n265) );
  XOR U399 ( .A(B[210]), .B(A[210]), .Z(n266) );
  XOR U400 ( .A(A[20]), .B(n267), .Z(O[20]) );
  AND U401 ( .A(S), .B(n268), .Z(n267) );
  XOR U402 ( .A(B[20]), .B(A[20]), .Z(n268) );
  XOR U403 ( .A(A[209]), .B(n269), .Z(O[209]) );
  AND U404 ( .A(S), .B(n270), .Z(n269) );
  XOR U405 ( .A(B[209]), .B(A[209]), .Z(n270) );
  XOR U406 ( .A(A[208]), .B(n271), .Z(O[208]) );
  AND U407 ( .A(S), .B(n272), .Z(n271) );
  XOR U408 ( .A(B[208]), .B(A[208]), .Z(n272) );
  XOR U409 ( .A(A[207]), .B(n273), .Z(O[207]) );
  AND U410 ( .A(S), .B(n274), .Z(n273) );
  XOR U411 ( .A(B[207]), .B(A[207]), .Z(n274) );
  XOR U412 ( .A(A[206]), .B(n275), .Z(O[206]) );
  AND U413 ( .A(S), .B(n276), .Z(n275) );
  XOR U414 ( .A(B[206]), .B(A[206]), .Z(n276) );
  XOR U415 ( .A(A[205]), .B(n277), .Z(O[205]) );
  AND U416 ( .A(S), .B(n278), .Z(n277) );
  XOR U417 ( .A(B[205]), .B(A[205]), .Z(n278) );
  XOR U418 ( .A(A[204]), .B(n279), .Z(O[204]) );
  AND U419 ( .A(S), .B(n280), .Z(n279) );
  XOR U420 ( .A(B[204]), .B(A[204]), .Z(n280) );
  XOR U421 ( .A(A[203]), .B(n281), .Z(O[203]) );
  AND U422 ( .A(S), .B(n282), .Z(n281) );
  XOR U423 ( .A(B[203]), .B(A[203]), .Z(n282) );
  XOR U424 ( .A(A[202]), .B(n283), .Z(O[202]) );
  AND U425 ( .A(S), .B(n284), .Z(n283) );
  XOR U426 ( .A(B[202]), .B(A[202]), .Z(n284) );
  XOR U427 ( .A(A[201]), .B(n285), .Z(O[201]) );
  AND U428 ( .A(S), .B(n286), .Z(n285) );
  XOR U429 ( .A(B[201]), .B(A[201]), .Z(n286) );
  XOR U430 ( .A(A[200]), .B(n287), .Z(O[200]) );
  AND U431 ( .A(S), .B(n288), .Z(n287) );
  XOR U432 ( .A(B[200]), .B(A[200]), .Z(n288) );
  XOR U433 ( .A(A[1]), .B(n289), .Z(O[1]) );
  AND U434 ( .A(S), .B(n290), .Z(n289) );
  XOR U435 ( .A(B[1]), .B(A[1]), .Z(n290) );
  XOR U436 ( .A(A[19]), .B(n291), .Z(O[19]) );
  AND U437 ( .A(S), .B(n292), .Z(n291) );
  XOR U438 ( .A(B[19]), .B(A[19]), .Z(n292) );
  XOR U439 ( .A(A[199]), .B(n293), .Z(O[199]) );
  AND U440 ( .A(S), .B(n294), .Z(n293) );
  XOR U441 ( .A(B[199]), .B(A[199]), .Z(n294) );
  XOR U442 ( .A(A[198]), .B(n295), .Z(O[198]) );
  AND U443 ( .A(S), .B(n296), .Z(n295) );
  XOR U444 ( .A(B[198]), .B(A[198]), .Z(n296) );
  XOR U445 ( .A(A[197]), .B(n297), .Z(O[197]) );
  AND U446 ( .A(S), .B(n298), .Z(n297) );
  XOR U447 ( .A(B[197]), .B(A[197]), .Z(n298) );
  XOR U448 ( .A(A[196]), .B(n299), .Z(O[196]) );
  AND U449 ( .A(S), .B(n300), .Z(n299) );
  XOR U450 ( .A(B[196]), .B(A[196]), .Z(n300) );
  XOR U451 ( .A(A[195]), .B(n301), .Z(O[195]) );
  AND U452 ( .A(S), .B(n302), .Z(n301) );
  XOR U453 ( .A(B[195]), .B(A[195]), .Z(n302) );
  XOR U454 ( .A(A[194]), .B(n303), .Z(O[194]) );
  AND U455 ( .A(S), .B(n304), .Z(n303) );
  XOR U456 ( .A(B[194]), .B(A[194]), .Z(n304) );
  XOR U457 ( .A(A[193]), .B(n305), .Z(O[193]) );
  AND U458 ( .A(S), .B(n306), .Z(n305) );
  XOR U459 ( .A(B[193]), .B(A[193]), .Z(n306) );
  XOR U460 ( .A(A[192]), .B(n307), .Z(O[192]) );
  AND U461 ( .A(S), .B(n308), .Z(n307) );
  XOR U462 ( .A(B[192]), .B(A[192]), .Z(n308) );
  XOR U463 ( .A(A[191]), .B(n309), .Z(O[191]) );
  AND U464 ( .A(S), .B(n310), .Z(n309) );
  XOR U465 ( .A(B[191]), .B(A[191]), .Z(n310) );
  XOR U466 ( .A(A[190]), .B(n311), .Z(O[190]) );
  AND U467 ( .A(S), .B(n312), .Z(n311) );
  XOR U468 ( .A(B[190]), .B(A[190]), .Z(n312) );
  XOR U469 ( .A(A[18]), .B(n313), .Z(O[18]) );
  AND U470 ( .A(S), .B(n314), .Z(n313) );
  XOR U471 ( .A(B[18]), .B(A[18]), .Z(n314) );
  XOR U472 ( .A(A[189]), .B(n315), .Z(O[189]) );
  AND U473 ( .A(S), .B(n316), .Z(n315) );
  XOR U474 ( .A(B[189]), .B(A[189]), .Z(n316) );
  XOR U475 ( .A(A[188]), .B(n317), .Z(O[188]) );
  AND U476 ( .A(S), .B(n318), .Z(n317) );
  XOR U477 ( .A(B[188]), .B(A[188]), .Z(n318) );
  XOR U478 ( .A(A[187]), .B(n319), .Z(O[187]) );
  AND U479 ( .A(S), .B(n320), .Z(n319) );
  XOR U480 ( .A(B[187]), .B(A[187]), .Z(n320) );
  XOR U481 ( .A(A[186]), .B(n321), .Z(O[186]) );
  AND U482 ( .A(S), .B(n322), .Z(n321) );
  XOR U483 ( .A(B[186]), .B(A[186]), .Z(n322) );
  XOR U484 ( .A(A[185]), .B(n323), .Z(O[185]) );
  AND U485 ( .A(S), .B(n324), .Z(n323) );
  XOR U486 ( .A(B[185]), .B(A[185]), .Z(n324) );
  XOR U487 ( .A(A[184]), .B(n325), .Z(O[184]) );
  AND U488 ( .A(S), .B(n326), .Z(n325) );
  XOR U489 ( .A(B[184]), .B(A[184]), .Z(n326) );
  XOR U490 ( .A(A[183]), .B(n327), .Z(O[183]) );
  AND U491 ( .A(S), .B(n328), .Z(n327) );
  XOR U492 ( .A(B[183]), .B(A[183]), .Z(n328) );
  XOR U493 ( .A(A[182]), .B(n329), .Z(O[182]) );
  AND U494 ( .A(S), .B(n330), .Z(n329) );
  XOR U495 ( .A(B[182]), .B(A[182]), .Z(n330) );
  XOR U496 ( .A(A[181]), .B(n331), .Z(O[181]) );
  AND U497 ( .A(S), .B(n332), .Z(n331) );
  XOR U498 ( .A(B[181]), .B(A[181]), .Z(n332) );
  XOR U499 ( .A(A[180]), .B(n333), .Z(O[180]) );
  AND U500 ( .A(S), .B(n334), .Z(n333) );
  XOR U501 ( .A(B[180]), .B(A[180]), .Z(n334) );
  XOR U502 ( .A(A[17]), .B(n335), .Z(O[17]) );
  AND U503 ( .A(S), .B(n336), .Z(n335) );
  XOR U504 ( .A(B[17]), .B(A[17]), .Z(n336) );
  XOR U505 ( .A(A[179]), .B(n337), .Z(O[179]) );
  AND U506 ( .A(S), .B(n338), .Z(n337) );
  XOR U507 ( .A(B[179]), .B(A[179]), .Z(n338) );
  XOR U508 ( .A(A[178]), .B(n339), .Z(O[178]) );
  AND U509 ( .A(S), .B(n340), .Z(n339) );
  XOR U510 ( .A(B[178]), .B(A[178]), .Z(n340) );
  XOR U511 ( .A(A[177]), .B(n341), .Z(O[177]) );
  AND U512 ( .A(S), .B(n342), .Z(n341) );
  XOR U513 ( .A(B[177]), .B(A[177]), .Z(n342) );
  XOR U514 ( .A(A[176]), .B(n343), .Z(O[176]) );
  AND U515 ( .A(S), .B(n344), .Z(n343) );
  XOR U516 ( .A(B[176]), .B(A[176]), .Z(n344) );
  XOR U517 ( .A(A[175]), .B(n345), .Z(O[175]) );
  AND U518 ( .A(S), .B(n346), .Z(n345) );
  XOR U519 ( .A(B[175]), .B(A[175]), .Z(n346) );
  XOR U520 ( .A(A[174]), .B(n347), .Z(O[174]) );
  AND U521 ( .A(S), .B(n348), .Z(n347) );
  XOR U522 ( .A(B[174]), .B(A[174]), .Z(n348) );
  XOR U523 ( .A(A[173]), .B(n349), .Z(O[173]) );
  AND U524 ( .A(S), .B(n350), .Z(n349) );
  XOR U525 ( .A(B[173]), .B(A[173]), .Z(n350) );
  XOR U526 ( .A(A[172]), .B(n351), .Z(O[172]) );
  AND U527 ( .A(S), .B(n352), .Z(n351) );
  XOR U528 ( .A(B[172]), .B(A[172]), .Z(n352) );
  XOR U529 ( .A(A[171]), .B(n353), .Z(O[171]) );
  AND U530 ( .A(S), .B(n354), .Z(n353) );
  XOR U531 ( .A(B[171]), .B(A[171]), .Z(n354) );
  XOR U532 ( .A(A[170]), .B(n355), .Z(O[170]) );
  AND U533 ( .A(S), .B(n356), .Z(n355) );
  XOR U534 ( .A(B[170]), .B(A[170]), .Z(n356) );
  XOR U535 ( .A(A[16]), .B(n357), .Z(O[16]) );
  AND U536 ( .A(S), .B(n358), .Z(n357) );
  XOR U537 ( .A(B[16]), .B(A[16]), .Z(n358) );
  XOR U538 ( .A(A[169]), .B(n359), .Z(O[169]) );
  AND U539 ( .A(S), .B(n360), .Z(n359) );
  XOR U540 ( .A(B[169]), .B(A[169]), .Z(n360) );
  XOR U541 ( .A(A[168]), .B(n361), .Z(O[168]) );
  AND U542 ( .A(S), .B(n362), .Z(n361) );
  XOR U543 ( .A(B[168]), .B(A[168]), .Z(n362) );
  XOR U544 ( .A(A[167]), .B(n363), .Z(O[167]) );
  AND U545 ( .A(S), .B(n364), .Z(n363) );
  XOR U546 ( .A(B[167]), .B(A[167]), .Z(n364) );
  XOR U547 ( .A(A[166]), .B(n365), .Z(O[166]) );
  AND U548 ( .A(S), .B(n366), .Z(n365) );
  XOR U549 ( .A(B[166]), .B(A[166]), .Z(n366) );
  XOR U550 ( .A(A[165]), .B(n367), .Z(O[165]) );
  AND U551 ( .A(S), .B(n368), .Z(n367) );
  XOR U552 ( .A(B[165]), .B(A[165]), .Z(n368) );
  XOR U553 ( .A(A[164]), .B(n369), .Z(O[164]) );
  AND U554 ( .A(S), .B(n370), .Z(n369) );
  XOR U555 ( .A(B[164]), .B(A[164]), .Z(n370) );
  XOR U556 ( .A(A[163]), .B(n371), .Z(O[163]) );
  AND U557 ( .A(S), .B(n372), .Z(n371) );
  XOR U558 ( .A(B[163]), .B(A[163]), .Z(n372) );
  XOR U559 ( .A(A[162]), .B(n373), .Z(O[162]) );
  AND U560 ( .A(S), .B(n374), .Z(n373) );
  XOR U561 ( .A(B[162]), .B(A[162]), .Z(n374) );
  XOR U562 ( .A(A[161]), .B(n375), .Z(O[161]) );
  AND U563 ( .A(S), .B(n376), .Z(n375) );
  XOR U564 ( .A(B[161]), .B(A[161]), .Z(n376) );
  XOR U565 ( .A(A[160]), .B(n377), .Z(O[160]) );
  AND U566 ( .A(S), .B(n378), .Z(n377) );
  XOR U567 ( .A(B[160]), .B(A[160]), .Z(n378) );
  XOR U568 ( .A(A[15]), .B(n379), .Z(O[15]) );
  AND U569 ( .A(S), .B(n380), .Z(n379) );
  XOR U570 ( .A(B[15]), .B(A[15]), .Z(n380) );
  XOR U571 ( .A(A[159]), .B(n381), .Z(O[159]) );
  AND U572 ( .A(S), .B(n382), .Z(n381) );
  XOR U573 ( .A(B[159]), .B(A[159]), .Z(n382) );
  XOR U574 ( .A(A[158]), .B(n383), .Z(O[158]) );
  AND U575 ( .A(S), .B(n384), .Z(n383) );
  XOR U576 ( .A(B[158]), .B(A[158]), .Z(n384) );
  XOR U577 ( .A(A[157]), .B(n385), .Z(O[157]) );
  AND U578 ( .A(S), .B(n386), .Z(n385) );
  XOR U579 ( .A(B[157]), .B(A[157]), .Z(n386) );
  XOR U580 ( .A(A[156]), .B(n387), .Z(O[156]) );
  AND U581 ( .A(S), .B(n388), .Z(n387) );
  XOR U582 ( .A(B[156]), .B(A[156]), .Z(n388) );
  XOR U583 ( .A(A[155]), .B(n389), .Z(O[155]) );
  AND U584 ( .A(S), .B(n390), .Z(n389) );
  XOR U585 ( .A(B[155]), .B(A[155]), .Z(n390) );
  XOR U586 ( .A(A[154]), .B(n391), .Z(O[154]) );
  AND U587 ( .A(S), .B(n392), .Z(n391) );
  XOR U588 ( .A(B[154]), .B(A[154]), .Z(n392) );
  XOR U589 ( .A(A[153]), .B(n393), .Z(O[153]) );
  AND U590 ( .A(S), .B(n394), .Z(n393) );
  XOR U591 ( .A(B[153]), .B(A[153]), .Z(n394) );
  XOR U592 ( .A(A[152]), .B(n395), .Z(O[152]) );
  AND U593 ( .A(S), .B(n396), .Z(n395) );
  XOR U594 ( .A(B[152]), .B(A[152]), .Z(n396) );
  XOR U595 ( .A(A[151]), .B(n397), .Z(O[151]) );
  AND U596 ( .A(S), .B(n398), .Z(n397) );
  XOR U597 ( .A(B[151]), .B(A[151]), .Z(n398) );
  XOR U598 ( .A(A[150]), .B(n399), .Z(O[150]) );
  AND U599 ( .A(S), .B(n400), .Z(n399) );
  XOR U600 ( .A(B[150]), .B(A[150]), .Z(n400) );
  XOR U601 ( .A(A[14]), .B(n401), .Z(O[14]) );
  AND U602 ( .A(S), .B(n402), .Z(n401) );
  XOR U603 ( .A(B[14]), .B(A[14]), .Z(n402) );
  XOR U604 ( .A(A[149]), .B(n403), .Z(O[149]) );
  AND U605 ( .A(S), .B(n404), .Z(n403) );
  XOR U606 ( .A(B[149]), .B(A[149]), .Z(n404) );
  XOR U607 ( .A(A[148]), .B(n405), .Z(O[148]) );
  AND U608 ( .A(S), .B(n406), .Z(n405) );
  XOR U609 ( .A(B[148]), .B(A[148]), .Z(n406) );
  XOR U610 ( .A(A[147]), .B(n407), .Z(O[147]) );
  AND U611 ( .A(S), .B(n408), .Z(n407) );
  XOR U612 ( .A(B[147]), .B(A[147]), .Z(n408) );
  XOR U613 ( .A(A[146]), .B(n409), .Z(O[146]) );
  AND U614 ( .A(S), .B(n410), .Z(n409) );
  XOR U615 ( .A(B[146]), .B(A[146]), .Z(n410) );
  XOR U616 ( .A(A[145]), .B(n411), .Z(O[145]) );
  AND U617 ( .A(S), .B(n412), .Z(n411) );
  XOR U618 ( .A(B[145]), .B(A[145]), .Z(n412) );
  XOR U619 ( .A(A[144]), .B(n413), .Z(O[144]) );
  AND U620 ( .A(S), .B(n414), .Z(n413) );
  XOR U621 ( .A(B[144]), .B(A[144]), .Z(n414) );
  XOR U622 ( .A(A[143]), .B(n415), .Z(O[143]) );
  AND U623 ( .A(S), .B(n416), .Z(n415) );
  XOR U624 ( .A(B[143]), .B(A[143]), .Z(n416) );
  XOR U625 ( .A(A[142]), .B(n417), .Z(O[142]) );
  AND U626 ( .A(S), .B(n418), .Z(n417) );
  XOR U627 ( .A(B[142]), .B(A[142]), .Z(n418) );
  XOR U628 ( .A(A[141]), .B(n419), .Z(O[141]) );
  AND U629 ( .A(S), .B(n420), .Z(n419) );
  XOR U630 ( .A(B[141]), .B(A[141]), .Z(n420) );
  XOR U631 ( .A(A[140]), .B(n421), .Z(O[140]) );
  AND U632 ( .A(S), .B(n422), .Z(n421) );
  XOR U633 ( .A(B[140]), .B(A[140]), .Z(n422) );
  XOR U634 ( .A(A[13]), .B(n423), .Z(O[13]) );
  AND U635 ( .A(S), .B(n424), .Z(n423) );
  XOR U636 ( .A(B[13]), .B(A[13]), .Z(n424) );
  XOR U637 ( .A(A[139]), .B(n425), .Z(O[139]) );
  AND U638 ( .A(S), .B(n426), .Z(n425) );
  XOR U639 ( .A(B[139]), .B(A[139]), .Z(n426) );
  XOR U640 ( .A(A[138]), .B(n427), .Z(O[138]) );
  AND U641 ( .A(S), .B(n428), .Z(n427) );
  XOR U642 ( .A(B[138]), .B(A[138]), .Z(n428) );
  XOR U643 ( .A(A[137]), .B(n429), .Z(O[137]) );
  AND U644 ( .A(S), .B(n430), .Z(n429) );
  XOR U645 ( .A(B[137]), .B(A[137]), .Z(n430) );
  XOR U646 ( .A(A[136]), .B(n431), .Z(O[136]) );
  AND U647 ( .A(S), .B(n432), .Z(n431) );
  XOR U648 ( .A(B[136]), .B(A[136]), .Z(n432) );
  XOR U649 ( .A(A[135]), .B(n433), .Z(O[135]) );
  AND U650 ( .A(S), .B(n434), .Z(n433) );
  XOR U651 ( .A(B[135]), .B(A[135]), .Z(n434) );
  XOR U652 ( .A(A[134]), .B(n435), .Z(O[134]) );
  AND U653 ( .A(S), .B(n436), .Z(n435) );
  XOR U654 ( .A(B[134]), .B(A[134]), .Z(n436) );
  XOR U655 ( .A(A[133]), .B(n437), .Z(O[133]) );
  AND U656 ( .A(S), .B(n438), .Z(n437) );
  XOR U657 ( .A(B[133]), .B(A[133]), .Z(n438) );
  XOR U658 ( .A(A[132]), .B(n439), .Z(O[132]) );
  AND U659 ( .A(S), .B(n440), .Z(n439) );
  XOR U660 ( .A(B[132]), .B(A[132]), .Z(n440) );
  XOR U661 ( .A(A[131]), .B(n441), .Z(O[131]) );
  AND U662 ( .A(S), .B(n442), .Z(n441) );
  XOR U663 ( .A(B[131]), .B(A[131]), .Z(n442) );
  XOR U664 ( .A(A[130]), .B(n443), .Z(O[130]) );
  AND U665 ( .A(S), .B(n444), .Z(n443) );
  XOR U666 ( .A(B[130]), .B(A[130]), .Z(n444) );
  XOR U667 ( .A(A[12]), .B(n445), .Z(O[12]) );
  AND U668 ( .A(S), .B(n446), .Z(n445) );
  XOR U669 ( .A(B[12]), .B(A[12]), .Z(n446) );
  XOR U670 ( .A(A[129]), .B(n447), .Z(O[129]) );
  AND U671 ( .A(S), .B(n448), .Z(n447) );
  XOR U672 ( .A(B[129]), .B(A[129]), .Z(n448) );
  XOR U673 ( .A(A[128]), .B(n449), .Z(O[128]) );
  AND U674 ( .A(S), .B(n450), .Z(n449) );
  XOR U675 ( .A(B[128]), .B(A[128]), .Z(n450) );
  XOR U676 ( .A(A[127]), .B(n451), .Z(O[127]) );
  AND U677 ( .A(S), .B(n452), .Z(n451) );
  XOR U678 ( .A(B[127]), .B(A[127]), .Z(n452) );
  XOR U679 ( .A(A[126]), .B(n453), .Z(O[126]) );
  AND U680 ( .A(S), .B(n454), .Z(n453) );
  XOR U681 ( .A(B[126]), .B(A[126]), .Z(n454) );
  XOR U682 ( .A(A[125]), .B(n455), .Z(O[125]) );
  AND U683 ( .A(S), .B(n456), .Z(n455) );
  XOR U684 ( .A(B[125]), .B(A[125]), .Z(n456) );
  XOR U685 ( .A(A[124]), .B(n457), .Z(O[124]) );
  AND U686 ( .A(S), .B(n458), .Z(n457) );
  XOR U687 ( .A(B[124]), .B(A[124]), .Z(n458) );
  XOR U688 ( .A(A[123]), .B(n459), .Z(O[123]) );
  AND U689 ( .A(S), .B(n460), .Z(n459) );
  XOR U690 ( .A(B[123]), .B(A[123]), .Z(n460) );
  XOR U691 ( .A(A[122]), .B(n461), .Z(O[122]) );
  AND U692 ( .A(S), .B(n462), .Z(n461) );
  XOR U693 ( .A(B[122]), .B(A[122]), .Z(n462) );
  XOR U694 ( .A(A[121]), .B(n463), .Z(O[121]) );
  AND U695 ( .A(S), .B(n464), .Z(n463) );
  XOR U696 ( .A(B[121]), .B(A[121]), .Z(n464) );
  XOR U697 ( .A(A[120]), .B(n465), .Z(O[120]) );
  AND U698 ( .A(S), .B(n466), .Z(n465) );
  XOR U699 ( .A(B[120]), .B(A[120]), .Z(n466) );
  XOR U700 ( .A(A[11]), .B(n467), .Z(O[11]) );
  AND U701 ( .A(S), .B(n468), .Z(n467) );
  XOR U702 ( .A(B[11]), .B(A[11]), .Z(n468) );
  XOR U703 ( .A(A[119]), .B(n469), .Z(O[119]) );
  AND U704 ( .A(S), .B(n470), .Z(n469) );
  XOR U705 ( .A(B[119]), .B(A[119]), .Z(n470) );
  XOR U706 ( .A(A[118]), .B(n471), .Z(O[118]) );
  AND U707 ( .A(S), .B(n472), .Z(n471) );
  XOR U708 ( .A(B[118]), .B(A[118]), .Z(n472) );
  XOR U709 ( .A(A[117]), .B(n473), .Z(O[117]) );
  AND U710 ( .A(S), .B(n474), .Z(n473) );
  XOR U711 ( .A(B[117]), .B(A[117]), .Z(n474) );
  XOR U712 ( .A(A[116]), .B(n475), .Z(O[116]) );
  AND U713 ( .A(S), .B(n476), .Z(n475) );
  XOR U714 ( .A(B[116]), .B(A[116]), .Z(n476) );
  XOR U715 ( .A(A[115]), .B(n477), .Z(O[115]) );
  AND U716 ( .A(S), .B(n478), .Z(n477) );
  XOR U717 ( .A(B[115]), .B(A[115]), .Z(n478) );
  XOR U718 ( .A(A[114]), .B(n479), .Z(O[114]) );
  AND U719 ( .A(S), .B(n480), .Z(n479) );
  XOR U720 ( .A(B[114]), .B(A[114]), .Z(n480) );
  XOR U721 ( .A(A[113]), .B(n481), .Z(O[113]) );
  AND U722 ( .A(S), .B(n482), .Z(n481) );
  XOR U723 ( .A(B[113]), .B(A[113]), .Z(n482) );
  XOR U724 ( .A(A[112]), .B(n483), .Z(O[112]) );
  AND U725 ( .A(S), .B(n484), .Z(n483) );
  XOR U726 ( .A(B[112]), .B(A[112]), .Z(n484) );
  XOR U727 ( .A(A[111]), .B(n485), .Z(O[111]) );
  AND U728 ( .A(S), .B(n486), .Z(n485) );
  XOR U729 ( .A(B[111]), .B(A[111]), .Z(n486) );
  XOR U730 ( .A(A[110]), .B(n487), .Z(O[110]) );
  AND U731 ( .A(S), .B(n488), .Z(n487) );
  XOR U732 ( .A(B[110]), .B(A[110]), .Z(n488) );
  XOR U733 ( .A(A[10]), .B(n489), .Z(O[10]) );
  AND U734 ( .A(S), .B(n490), .Z(n489) );
  XOR U735 ( .A(B[10]), .B(A[10]), .Z(n490) );
  XOR U736 ( .A(A[109]), .B(n491), .Z(O[109]) );
  AND U737 ( .A(S), .B(n492), .Z(n491) );
  XOR U738 ( .A(B[109]), .B(A[109]), .Z(n492) );
  XOR U739 ( .A(A[108]), .B(n493), .Z(O[108]) );
  AND U740 ( .A(S), .B(n494), .Z(n493) );
  XOR U741 ( .A(B[108]), .B(A[108]), .Z(n494) );
  XOR U742 ( .A(A[107]), .B(n495), .Z(O[107]) );
  AND U743 ( .A(S), .B(n496), .Z(n495) );
  XOR U744 ( .A(B[107]), .B(A[107]), .Z(n496) );
  XOR U745 ( .A(A[106]), .B(n497), .Z(O[106]) );
  AND U746 ( .A(S), .B(n498), .Z(n497) );
  XOR U747 ( .A(B[106]), .B(A[106]), .Z(n498) );
  XOR U748 ( .A(A[105]), .B(n499), .Z(O[105]) );
  AND U749 ( .A(S), .B(n500), .Z(n499) );
  XOR U750 ( .A(B[105]), .B(A[105]), .Z(n500) );
  XOR U751 ( .A(A[104]), .B(n501), .Z(O[104]) );
  AND U752 ( .A(S), .B(n502), .Z(n501) );
  XOR U753 ( .A(B[104]), .B(A[104]), .Z(n502) );
  XOR U754 ( .A(A[103]), .B(n503), .Z(O[103]) );
  AND U755 ( .A(S), .B(n504), .Z(n503) );
  XOR U756 ( .A(B[103]), .B(A[103]), .Z(n504) );
  XOR U757 ( .A(A[102]), .B(n505), .Z(O[102]) );
  AND U758 ( .A(S), .B(n506), .Z(n505) );
  XOR U759 ( .A(B[102]), .B(A[102]), .Z(n506) );
  XOR U760 ( .A(A[101]), .B(n507), .Z(O[101]) );
  AND U761 ( .A(S), .B(n508), .Z(n507) );
  XOR U762 ( .A(B[101]), .B(A[101]), .Z(n508) );
  XOR U763 ( .A(A[100]), .B(n509), .Z(O[100]) );
  AND U764 ( .A(S), .B(n510), .Z(n509) );
  XOR U765 ( .A(B[100]), .B(A[100]), .Z(n510) );
  XOR U766 ( .A(A[0]), .B(n511), .Z(O[0]) );
  AND U767 ( .A(S), .B(n512), .Z(n511) );
  XOR U768 ( .A(B[0]), .B(A[0]), .Z(n512) );
endmodule


module MUX_N258_3 ( A, B, S, O );
  input [257:0] A;
  input [257:0] B;
  output [257:0] O;
  input S;


  ANDN U1 ( .B(A[9]), .A(S), .Z(O[9]) );
  ANDN U2 ( .B(A[99]), .A(S), .Z(O[99]) );
  ANDN U3 ( .B(A[98]), .A(S), .Z(O[98]) );
  ANDN U4 ( .B(A[97]), .A(S), .Z(O[97]) );
  ANDN U5 ( .B(A[96]), .A(S), .Z(O[96]) );
  ANDN U6 ( .B(A[95]), .A(S), .Z(O[95]) );
  ANDN U7 ( .B(A[94]), .A(S), .Z(O[94]) );
  ANDN U8 ( .B(A[93]), .A(S), .Z(O[93]) );
  ANDN U9 ( .B(A[92]), .A(S), .Z(O[92]) );
  ANDN U10 ( .B(A[91]), .A(S), .Z(O[91]) );
  ANDN U11 ( .B(A[90]), .A(S), .Z(O[90]) );
  ANDN U12 ( .B(A[8]), .A(S), .Z(O[8]) );
  ANDN U13 ( .B(A[89]), .A(S), .Z(O[89]) );
  ANDN U14 ( .B(A[88]), .A(S), .Z(O[88]) );
  ANDN U15 ( .B(A[87]), .A(S), .Z(O[87]) );
  ANDN U16 ( .B(A[86]), .A(S), .Z(O[86]) );
  ANDN U17 ( .B(A[85]), .A(S), .Z(O[85]) );
  ANDN U18 ( .B(A[84]), .A(S), .Z(O[84]) );
  ANDN U19 ( .B(A[83]), .A(S), .Z(O[83]) );
  ANDN U20 ( .B(A[82]), .A(S), .Z(O[82]) );
  ANDN U21 ( .B(A[81]), .A(S), .Z(O[81]) );
  ANDN U22 ( .B(A[80]), .A(S), .Z(O[80]) );
  ANDN U23 ( .B(A[7]), .A(S), .Z(O[7]) );
  ANDN U24 ( .B(A[79]), .A(S), .Z(O[79]) );
  ANDN U25 ( .B(A[78]), .A(S), .Z(O[78]) );
  ANDN U26 ( .B(A[77]), .A(S), .Z(O[77]) );
  ANDN U27 ( .B(A[76]), .A(S), .Z(O[76]) );
  ANDN U28 ( .B(A[75]), .A(S), .Z(O[75]) );
  ANDN U29 ( .B(A[74]), .A(S), .Z(O[74]) );
  ANDN U30 ( .B(A[73]), .A(S), .Z(O[73]) );
  ANDN U31 ( .B(A[72]), .A(S), .Z(O[72]) );
  ANDN U32 ( .B(A[71]), .A(S), .Z(O[71]) );
  ANDN U33 ( .B(A[70]), .A(S), .Z(O[70]) );
  ANDN U34 ( .B(A[6]), .A(S), .Z(O[6]) );
  ANDN U35 ( .B(A[69]), .A(S), .Z(O[69]) );
  ANDN U36 ( .B(A[68]), .A(S), .Z(O[68]) );
  ANDN U37 ( .B(A[67]), .A(S), .Z(O[67]) );
  ANDN U38 ( .B(A[66]), .A(S), .Z(O[66]) );
  ANDN U39 ( .B(A[65]), .A(S), .Z(O[65]) );
  ANDN U40 ( .B(A[64]), .A(S), .Z(O[64]) );
  ANDN U41 ( .B(A[63]), .A(S), .Z(O[63]) );
  ANDN U42 ( .B(A[62]), .A(S), .Z(O[62]) );
  ANDN U43 ( .B(A[61]), .A(S), .Z(O[61]) );
  ANDN U44 ( .B(A[60]), .A(S), .Z(O[60]) );
  ANDN U45 ( .B(A[5]), .A(S), .Z(O[5]) );
  ANDN U46 ( .B(A[59]), .A(S), .Z(O[59]) );
  ANDN U47 ( .B(A[58]), .A(S), .Z(O[58]) );
  ANDN U48 ( .B(A[57]), .A(S), .Z(O[57]) );
  ANDN U49 ( .B(A[56]), .A(S), .Z(O[56]) );
  ANDN U50 ( .B(A[55]), .A(S), .Z(O[55]) );
  ANDN U51 ( .B(A[54]), .A(S), .Z(O[54]) );
  ANDN U52 ( .B(A[53]), .A(S), .Z(O[53]) );
  ANDN U53 ( .B(A[52]), .A(S), .Z(O[52]) );
  ANDN U54 ( .B(A[51]), .A(S), .Z(O[51]) );
  ANDN U55 ( .B(A[50]), .A(S), .Z(O[50]) );
  ANDN U56 ( .B(A[4]), .A(S), .Z(O[4]) );
  ANDN U57 ( .B(A[49]), .A(S), .Z(O[49]) );
  ANDN U58 ( .B(A[48]), .A(S), .Z(O[48]) );
  ANDN U59 ( .B(A[47]), .A(S), .Z(O[47]) );
  ANDN U60 ( .B(A[46]), .A(S), .Z(O[46]) );
  ANDN U61 ( .B(A[45]), .A(S), .Z(O[45]) );
  ANDN U62 ( .B(A[44]), .A(S), .Z(O[44]) );
  ANDN U63 ( .B(A[43]), .A(S), .Z(O[43]) );
  ANDN U64 ( .B(A[42]), .A(S), .Z(O[42]) );
  ANDN U65 ( .B(A[41]), .A(S), .Z(O[41]) );
  ANDN U66 ( .B(A[40]), .A(S), .Z(O[40]) );
  ANDN U67 ( .B(A[3]), .A(S), .Z(O[3]) );
  ANDN U68 ( .B(A[39]), .A(S), .Z(O[39]) );
  ANDN U69 ( .B(A[38]), .A(S), .Z(O[38]) );
  ANDN U70 ( .B(A[37]), .A(S), .Z(O[37]) );
  ANDN U71 ( .B(A[36]), .A(S), .Z(O[36]) );
  ANDN U72 ( .B(A[35]), .A(S), .Z(O[35]) );
  ANDN U73 ( .B(A[34]), .A(S), .Z(O[34]) );
  ANDN U74 ( .B(A[33]), .A(S), .Z(O[33]) );
  ANDN U75 ( .B(A[32]), .A(S), .Z(O[32]) );
  ANDN U76 ( .B(A[31]), .A(S), .Z(O[31]) );
  ANDN U77 ( .B(A[30]), .A(S), .Z(O[30]) );
  ANDN U78 ( .B(A[2]), .A(S), .Z(O[2]) );
  ANDN U79 ( .B(A[29]), .A(S), .Z(O[29]) );
  ANDN U80 ( .B(A[28]), .A(S), .Z(O[28]) );
  ANDN U81 ( .B(A[27]), .A(S), .Z(O[27]) );
  ANDN U82 ( .B(A[26]), .A(S), .Z(O[26]) );
  ANDN U83 ( .B(A[25]), .A(S), .Z(O[25]) );
  ANDN U84 ( .B(A[255]), .A(S), .Z(O[255]) );
  ANDN U85 ( .B(A[254]), .A(S), .Z(O[254]) );
  ANDN U86 ( .B(A[253]), .A(S), .Z(O[253]) );
  ANDN U87 ( .B(A[252]), .A(S), .Z(O[252]) );
  ANDN U88 ( .B(A[251]), .A(S), .Z(O[251]) );
  ANDN U89 ( .B(A[250]), .A(S), .Z(O[250]) );
  ANDN U90 ( .B(A[24]), .A(S), .Z(O[24]) );
  ANDN U91 ( .B(A[249]), .A(S), .Z(O[249]) );
  ANDN U92 ( .B(A[248]), .A(S), .Z(O[248]) );
  ANDN U93 ( .B(A[247]), .A(S), .Z(O[247]) );
  ANDN U94 ( .B(A[246]), .A(S), .Z(O[246]) );
  ANDN U95 ( .B(A[245]), .A(S), .Z(O[245]) );
  ANDN U96 ( .B(A[244]), .A(S), .Z(O[244]) );
  ANDN U97 ( .B(A[243]), .A(S), .Z(O[243]) );
  ANDN U98 ( .B(A[242]), .A(S), .Z(O[242]) );
  ANDN U99 ( .B(A[241]), .A(S), .Z(O[241]) );
  ANDN U100 ( .B(A[240]), .A(S), .Z(O[240]) );
  ANDN U101 ( .B(A[23]), .A(S), .Z(O[23]) );
  ANDN U102 ( .B(A[239]), .A(S), .Z(O[239]) );
  ANDN U103 ( .B(A[238]), .A(S), .Z(O[238]) );
  ANDN U104 ( .B(A[237]), .A(S), .Z(O[237]) );
  ANDN U105 ( .B(A[236]), .A(S), .Z(O[236]) );
  ANDN U106 ( .B(A[235]), .A(S), .Z(O[235]) );
  ANDN U107 ( .B(A[234]), .A(S), .Z(O[234]) );
  ANDN U108 ( .B(A[233]), .A(S), .Z(O[233]) );
  ANDN U109 ( .B(A[232]), .A(S), .Z(O[232]) );
  ANDN U110 ( .B(A[231]), .A(S), .Z(O[231]) );
  ANDN U111 ( .B(A[230]), .A(S), .Z(O[230]) );
  ANDN U112 ( .B(A[22]), .A(S), .Z(O[22]) );
  ANDN U113 ( .B(A[229]), .A(S), .Z(O[229]) );
  ANDN U114 ( .B(A[228]), .A(S), .Z(O[228]) );
  ANDN U115 ( .B(A[227]), .A(S), .Z(O[227]) );
  ANDN U116 ( .B(A[226]), .A(S), .Z(O[226]) );
  ANDN U117 ( .B(A[225]), .A(S), .Z(O[225]) );
  ANDN U118 ( .B(A[224]), .A(S), .Z(O[224]) );
  ANDN U119 ( .B(A[223]), .A(S), .Z(O[223]) );
  ANDN U120 ( .B(A[222]), .A(S), .Z(O[222]) );
  ANDN U121 ( .B(A[221]), .A(S), .Z(O[221]) );
  ANDN U122 ( .B(A[220]), .A(S), .Z(O[220]) );
  ANDN U123 ( .B(A[21]), .A(S), .Z(O[21]) );
  ANDN U124 ( .B(A[219]), .A(S), .Z(O[219]) );
  ANDN U125 ( .B(A[218]), .A(S), .Z(O[218]) );
  ANDN U126 ( .B(A[217]), .A(S), .Z(O[217]) );
  ANDN U127 ( .B(A[216]), .A(S), .Z(O[216]) );
  ANDN U128 ( .B(A[215]), .A(S), .Z(O[215]) );
  ANDN U129 ( .B(A[214]), .A(S), .Z(O[214]) );
  ANDN U130 ( .B(A[213]), .A(S), .Z(O[213]) );
  ANDN U131 ( .B(A[212]), .A(S), .Z(O[212]) );
  ANDN U132 ( .B(A[211]), .A(S), .Z(O[211]) );
  ANDN U133 ( .B(A[210]), .A(S), .Z(O[210]) );
  ANDN U134 ( .B(A[20]), .A(S), .Z(O[20]) );
  ANDN U135 ( .B(A[209]), .A(S), .Z(O[209]) );
  ANDN U136 ( .B(A[208]), .A(S), .Z(O[208]) );
  ANDN U137 ( .B(A[207]), .A(S), .Z(O[207]) );
  ANDN U138 ( .B(A[206]), .A(S), .Z(O[206]) );
  ANDN U139 ( .B(A[205]), .A(S), .Z(O[205]) );
  ANDN U140 ( .B(A[204]), .A(S), .Z(O[204]) );
  ANDN U141 ( .B(A[203]), .A(S), .Z(O[203]) );
  ANDN U142 ( .B(A[202]), .A(S), .Z(O[202]) );
  ANDN U143 ( .B(A[201]), .A(S), .Z(O[201]) );
  ANDN U144 ( .B(A[200]), .A(S), .Z(O[200]) );
  ANDN U145 ( .B(A[1]), .A(S), .Z(O[1]) );
  ANDN U146 ( .B(A[19]), .A(S), .Z(O[19]) );
  ANDN U147 ( .B(A[199]), .A(S), .Z(O[199]) );
  ANDN U148 ( .B(A[198]), .A(S), .Z(O[198]) );
  ANDN U149 ( .B(A[197]), .A(S), .Z(O[197]) );
  ANDN U150 ( .B(A[196]), .A(S), .Z(O[196]) );
  ANDN U151 ( .B(A[195]), .A(S), .Z(O[195]) );
  ANDN U152 ( .B(A[194]), .A(S), .Z(O[194]) );
  ANDN U153 ( .B(A[193]), .A(S), .Z(O[193]) );
  ANDN U154 ( .B(A[192]), .A(S), .Z(O[192]) );
  ANDN U155 ( .B(A[191]), .A(S), .Z(O[191]) );
  ANDN U156 ( .B(A[190]), .A(S), .Z(O[190]) );
  ANDN U157 ( .B(A[18]), .A(S), .Z(O[18]) );
  ANDN U158 ( .B(A[189]), .A(S), .Z(O[189]) );
  ANDN U159 ( .B(A[188]), .A(S), .Z(O[188]) );
  ANDN U160 ( .B(A[187]), .A(S), .Z(O[187]) );
  ANDN U161 ( .B(A[186]), .A(S), .Z(O[186]) );
  ANDN U162 ( .B(A[185]), .A(S), .Z(O[185]) );
  ANDN U163 ( .B(A[184]), .A(S), .Z(O[184]) );
  ANDN U164 ( .B(A[183]), .A(S), .Z(O[183]) );
  ANDN U165 ( .B(A[182]), .A(S), .Z(O[182]) );
  ANDN U166 ( .B(A[181]), .A(S), .Z(O[181]) );
  ANDN U167 ( .B(A[180]), .A(S), .Z(O[180]) );
  ANDN U168 ( .B(A[17]), .A(S), .Z(O[17]) );
  ANDN U169 ( .B(A[179]), .A(S), .Z(O[179]) );
  ANDN U170 ( .B(A[178]), .A(S), .Z(O[178]) );
  ANDN U171 ( .B(A[177]), .A(S), .Z(O[177]) );
  ANDN U172 ( .B(A[176]), .A(S), .Z(O[176]) );
  ANDN U173 ( .B(A[175]), .A(S), .Z(O[175]) );
  ANDN U174 ( .B(A[174]), .A(S), .Z(O[174]) );
  ANDN U175 ( .B(A[173]), .A(S), .Z(O[173]) );
  ANDN U176 ( .B(A[172]), .A(S), .Z(O[172]) );
  ANDN U177 ( .B(A[171]), .A(S), .Z(O[171]) );
  ANDN U178 ( .B(A[170]), .A(S), .Z(O[170]) );
  ANDN U179 ( .B(A[16]), .A(S), .Z(O[16]) );
  ANDN U180 ( .B(A[169]), .A(S), .Z(O[169]) );
  ANDN U181 ( .B(A[168]), .A(S), .Z(O[168]) );
  ANDN U182 ( .B(A[167]), .A(S), .Z(O[167]) );
  ANDN U183 ( .B(A[166]), .A(S), .Z(O[166]) );
  ANDN U184 ( .B(A[165]), .A(S), .Z(O[165]) );
  ANDN U185 ( .B(A[164]), .A(S), .Z(O[164]) );
  ANDN U186 ( .B(A[163]), .A(S), .Z(O[163]) );
  ANDN U187 ( .B(A[162]), .A(S), .Z(O[162]) );
  ANDN U188 ( .B(A[161]), .A(S), .Z(O[161]) );
  ANDN U189 ( .B(A[160]), .A(S), .Z(O[160]) );
  ANDN U190 ( .B(A[15]), .A(S), .Z(O[15]) );
  ANDN U191 ( .B(A[159]), .A(S), .Z(O[159]) );
  ANDN U192 ( .B(A[158]), .A(S), .Z(O[158]) );
  ANDN U193 ( .B(A[157]), .A(S), .Z(O[157]) );
  ANDN U194 ( .B(A[156]), .A(S), .Z(O[156]) );
  ANDN U195 ( .B(A[155]), .A(S), .Z(O[155]) );
  ANDN U196 ( .B(A[154]), .A(S), .Z(O[154]) );
  ANDN U197 ( .B(A[153]), .A(S), .Z(O[153]) );
  ANDN U198 ( .B(A[152]), .A(S), .Z(O[152]) );
  ANDN U199 ( .B(A[151]), .A(S), .Z(O[151]) );
  ANDN U200 ( .B(A[150]), .A(S), .Z(O[150]) );
  ANDN U201 ( .B(A[14]), .A(S), .Z(O[14]) );
  ANDN U202 ( .B(A[149]), .A(S), .Z(O[149]) );
  ANDN U203 ( .B(A[148]), .A(S), .Z(O[148]) );
  ANDN U204 ( .B(A[147]), .A(S), .Z(O[147]) );
  ANDN U205 ( .B(A[146]), .A(S), .Z(O[146]) );
  ANDN U206 ( .B(A[145]), .A(S), .Z(O[145]) );
  ANDN U207 ( .B(A[144]), .A(S), .Z(O[144]) );
  ANDN U208 ( .B(A[143]), .A(S), .Z(O[143]) );
  ANDN U209 ( .B(A[142]), .A(S), .Z(O[142]) );
  ANDN U210 ( .B(A[141]), .A(S), .Z(O[141]) );
  ANDN U211 ( .B(A[140]), .A(S), .Z(O[140]) );
  ANDN U212 ( .B(A[13]), .A(S), .Z(O[13]) );
  ANDN U213 ( .B(A[139]), .A(S), .Z(O[139]) );
  ANDN U214 ( .B(A[138]), .A(S), .Z(O[138]) );
  ANDN U215 ( .B(A[137]), .A(S), .Z(O[137]) );
  ANDN U216 ( .B(A[136]), .A(S), .Z(O[136]) );
  ANDN U217 ( .B(A[135]), .A(S), .Z(O[135]) );
  ANDN U218 ( .B(A[134]), .A(S), .Z(O[134]) );
  ANDN U219 ( .B(A[133]), .A(S), .Z(O[133]) );
  ANDN U220 ( .B(A[132]), .A(S), .Z(O[132]) );
  ANDN U221 ( .B(A[131]), .A(S), .Z(O[131]) );
  ANDN U222 ( .B(A[130]), .A(S), .Z(O[130]) );
  ANDN U223 ( .B(A[12]), .A(S), .Z(O[12]) );
  ANDN U224 ( .B(A[129]), .A(S), .Z(O[129]) );
  ANDN U225 ( .B(A[128]), .A(S), .Z(O[128]) );
  ANDN U226 ( .B(A[127]), .A(S), .Z(O[127]) );
  ANDN U227 ( .B(A[126]), .A(S), .Z(O[126]) );
  ANDN U228 ( .B(A[125]), .A(S), .Z(O[125]) );
  ANDN U229 ( .B(A[124]), .A(S), .Z(O[124]) );
  ANDN U230 ( .B(A[123]), .A(S), .Z(O[123]) );
  ANDN U231 ( .B(A[122]), .A(S), .Z(O[122]) );
  ANDN U232 ( .B(A[121]), .A(S), .Z(O[121]) );
  ANDN U233 ( .B(A[120]), .A(S), .Z(O[120]) );
  ANDN U234 ( .B(A[11]), .A(S), .Z(O[11]) );
  ANDN U235 ( .B(A[119]), .A(S), .Z(O[119]) );
  ANDN U236 ( .B(A[118]), .A(S), .Z(O[118]) );
  ANDN U237 ( .B(A[117]), .A(S), .Z(O[117]) );
  ANDN U238 ( .B(A[116]), .A(S), .Z(O[116]) );
  ANDN U239 ( .B(A[115]), .A(S), .Z(O[115]) );
  ANDN U240 ( .B(A[114]), .A(S), .Z(O[114]) );
  ANDN U241 ( .B(A[113]), .A(S), .Z(O[113]) );
  ANDN U242 ( .B(A[112]), .A(S), .Z(O[112]) );
  ANDN U243 ( .B(A[111]), .A(S), .Z(O[111]) );
  ANDN U244 ( .B(A[110]), .A(S), .Z(O[110]) );
  ANDN U245 ( .B(A[10]), .A(S), .Z(O[10]) );
  ANDN U246 ( .B(A[109]), .A(S), .Z(O[109]) );
  ANDN U247 ( .B(A[108]), .A(S), .Z(O[108]) );
  ANDN U248 ( .B(A[107]), .A(S), .Z(O[107]) );
  ANDN U249 ( .B(A[106]), .A(S), .Z(O[106]) );
  ANDN U250 ( .B(A[105]), .A(S), .Z(O[105]) );
  ANDN U251 ( .B(A[104]), .A(S), .Z(O[104]) );
  ANDN U252 ( .B(A[103]), .A(S), .Z(O[103]) );
  ANDN U253 ( .B(A[102]), .A(S), .Z(O[102]) );
  ANDN U254 ( .B(A[101]), .A(S), .Z(O[101]) );
  ANDN U255 ( .B(A[100]), .A(S), .Z(O[100]) );
  ANDN U256 ( .B(A[0]), .A(S), .Z(O[0]) );
endmodule


module FA_1 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3612 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(CI), .B(A), .Z(S) );
endmodule


module FA_3613 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  ANDN U1 ( .B(CI), .A(S), .Z(CO) );
  XOR U2 ( .A(A), .B(CI), .Z(S) );
endmodule


module FA_3614 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3615 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3616 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3617 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3618 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3619 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3620 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3621 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3622 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3623 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3624 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3625 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3626 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3627 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3628 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3629 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3630 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3631 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3632 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3633 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3634 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3635 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3636 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3637 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3638 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3639 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3640 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3641 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3642 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3643 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3644 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3645 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3646 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3647 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3648 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3649 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3650 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3651 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3652 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3653 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3654 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3655 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3656 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3657 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3658 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3659 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3660 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3661 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3662 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3663 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3664 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3665 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3666 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3667 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3668 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3669 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3670 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3671 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3672 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3673 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3674 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3675 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3676 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3677 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3678 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3679 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3680 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3681 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3682 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3683 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3684 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3685 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3686 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3687 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3688 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3689 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3690 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3691 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3692 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3693 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3694 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3695 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3696 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3697 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3698 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3699 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3700 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3701 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3702 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3703 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3704 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3705 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3706 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3707 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3708 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3709 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3710 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3711 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3712 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3713 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3714 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3715 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3716 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3717 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3718 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3719 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3720 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3721 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3722 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3723 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3724 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3725 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3726 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3727 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3728 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3729 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3730 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3731 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3732 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3733 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3734 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3735 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3736 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3737 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3738 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3739 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3740 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3741 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3742 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3743 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3744 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3745 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3746 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3747 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3748 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3749 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3750 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3751 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3752 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3753 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3754 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3755 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3756 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3757 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3758 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3759 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3760 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3761 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3762 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3763 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3764 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3765 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3766 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3767 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3768 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3769 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3770 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3771 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3772 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3773 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3774 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3775 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3776 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3777 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3778 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3779 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3780 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3781 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3782 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3783 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3784 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3785 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3786 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3787 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3788 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3789 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3790 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3791 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3792 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3793 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3794 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3795 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3796 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3797 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3798 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3799 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3800 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3801 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3802 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3803 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3804 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3805 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3806 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3807 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3808 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3809 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3810 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3811 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3812 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3813 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3814 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3815 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3816 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3817 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3818 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3819 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3820 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3821 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3822 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3823 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3824 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3825 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3826 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3827 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3828 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3829 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3830 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3831 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3832 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3833 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3834 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3835 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3836 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3837 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3838 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3839 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3840 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3841 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3842 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3843 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3844 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3845 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3846 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3847 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3848 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3849 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3850 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3851 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3852 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3853 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3854 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3855 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3856 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3857 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3858 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3859 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3860 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3861 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3862 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3863 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3864 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3865 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3866 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3867 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3868 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module ADD_N258_1_0 ( A, B, CI, S, CO );
  input [257:0] A;
  input [257:0] B;
  output [257:0] S;
  input CI;
  output CO;

  wire   [257:1] C;

  FA_1 \FAINST[0].FA_  ( .A(1'b0), .B(B[0]), .CI(1'b0), .S(S[0]) );
  FA_3868 \FAINST[1].FA_  ( .A(A[1]), .B(B[1]), .CI(1'b0), .S(S[1]), .CO(C[2])
         );
  FA_3867 \FAINST[2].FA_  ( .A(A[2]), .B(B[2]), .CI(C[2]), .S(S[2]), .CO(C[3])
         );
  FA_3866 \FAINST[3].FA_  ( .A(A[3]), .B(B[3]), .CI(C[3]), .S(S[3]), .CO(C[4])
         );
  FA_3865 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(C[4]), .S(S[4]), .CO(C[5])
         );
  FA_3864 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_3863 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_3862 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_3861 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_3860 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_3859 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_3858 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_3857 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_3856 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_3855 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_3854 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_3853 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_3852 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_3851 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_3850 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_3849 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_3848 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_3847 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3846 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3845 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3844 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3843 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3842 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3841 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3840 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3839 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3838 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]), .CO(
        C[32]) );
  FA_3837 \FAINST[32].FA_  ( .A(A[32]), .B(B[32]), .CI(C[32]), .S(S[32]), .CO(
        C[33]) );
  FA_3836 \FAINST[33].FA_  ( .A(A[33]), .B(B[33]), .CI(C[33]), .S(S[33]), .CO(
        C[34]) );
  FA_3835 \FAINST[34].FA_  ( .A(A[34]), .B(B[34]), .CI(C[34]), .S(S[34]), .CO(
        C[35]) );
  FA_3834 \FAINST[35].FA_  ( .A(A[35]), .B(B[35]), .CI(C[35]), .S(S[35]), .CO(
        C[36]) );
  FA_3833 \FAINST[36].FA_  ( .A(A[36]), .B(B[36]), .CI(C[36]), .S(S[36]), .CO(
        C[37]) );
  FA_3832 \FAINST[37].FA_  ( .A(A[37]), .B(B[37]), .CI(C[37]), .S(S[37]), .CO(
        C[38]) );
  FA_3831 \FAINST[38].FA_  ( .A(A[38]), .B(B[38]), .CI(C[38]), .S(S[38]), .CO(
        C[39]) );
  FA_3830 \FAINST[39].FA_  ( .A(A[39]), .B(B[39]), .CI(C[39]), .S(S[39]), .CO(
        C[40]) );
  FA_3829 \FAINST[40].FA_  ( .A(A[40]), .B(B[40]), .CI(C[40]), .S(S[40]), .CO(
        C[41]) );
  FA_3828 \FAINST[41].FA_  ( .A(A[41]), .B(B[41]), .CI(C[41]), .S(S[41]), .CO(
        C[42]) );
  FA_3827 \FAINST[42].FA_  ( .A(A[42]), .B(B[42]), .CI(C[42]), .S(S[42]), .CO(
        C[43]) );
  FA_3826 \FAINST[43].FA_  ( .A(A[43]), .B(B[43]), .CI(C[43]), .S(S[43]), .CO(
        C[44]) );
  FA_3825 \FAINST[44].FA_  ( .A(A[44]), .B(B[44]), .CI(C[44]), .S(S[44]), .CO(
        C[45]) );
  FA_3824 \FAINST[45].FA_  ( .A(A[45]), .B(B[45]), .CI(C[45]), .S(S[45]), .CO(
        C[46]) );
  FA_3823 \FAINST[46].FA_  ( .A(A[46]), .B(B[46]), .CI(C[46]), .S(S[46]), .CO(
        C[47]) );
  FA_3822 \FAINST[47].FA_  ( .A(A[47]), .B(B[47]), .CI(C[47]), .S(S[47]), .CO(
        C[48]) );
  FA_3821 \FAINST[48].FA_  ( .A(A[48]), .B(B[48]), .CI(C[48]), .S(S[48]), .CO(
        C[49]) );
  FA_3820 \FAINST[49].FA_  ( .A(A[49]), .B(B[49]), .CI(C[49]), .S(S[49]), .CO(
        C[50]) );
  FA_3819 \FAINST[50].FA_  ( .A(A[50]), .B(B[50]), .CI(C[50]), .S(S[50]), .CO(
        C[51]) );
  FA_3818 \FAINST[51].FA_  ( .A(A[51]), .B(B[51]), .CI(C[51]), .S(S[51]), .CO(
        C[52]) );
  FA_3817 \FAINST[52].FA_  ( .A(A[52]), .B(B[52]), .CI(C[52]), .S(S[52]), .CO(
        C[53]) );
  FA_3816 \FAINST[53].FA_  ( .A(A[53]), .B(B[53]), .CI(C[53]), .S(S[53]), .CO(
        C[54]) );
  FA_3815 \FAINST[54].FA_  ( .A(A[54]), .B(B[54]), .CI(C[54]), .S(S[54]), .CO(
        C[55]) );
  FA_3814 \FAINST[55].FA_  ( .A(A[55]), .B(B[55]), .CI(C[55]), .S(S[55]), .CO(
        C[56]) );
  FA_3813 \FAINST[56].FA_  ( .A(A[56]), .B(B[56]), .CI(C[56]), .S(S[56]), .CO(
        C[57]) );
  FA_3812 \FAINST[57].FA_  ( .A(A[57]), .B(B[57]), .CI(C[57]), .S(S[57]), .CO(
        C[58]) );
  FA_3811 \FAINST[58].FA_  ( .A(A[58]), .B(B[58]), .CI(C[58]), .S(S[58]), .CO(
        C[59]) );
  FA_3810 \FAINST[59].FA_  ( .A(A[59]), .B(B[59]), .CI(C[59]), .S(S[59]), .CO(
        C[60]) );
  FA_3809 \FAINST[60].FA_  ( .A(A[60]), .B(B[60]), .CI(C[60]), .S(S[60]), .CO(
        C[61]) );
  FA_3808 \FAINST[61].FA_  ( .A(A[61]), .B(B[61]), .CI(C[61]), .S(S[61]), .CO(
        C[62]) );
  FA_3807 \FAINST[62].FA_  ( .A(A[62]), .B(B[62]), .CI(C[62]), .S(S[62]), .CO(
        C[63]) );
  FA_3806 \FAINST[63].FA_  ( .A(A[63]), .B(B[63]), .CI(C[63]), .S(S[63]), .CO(
        C[64]) );
  FA_3805 \FAINST[64].FA_  ( .A(A[64]), .B(B[64]), .CI(C[64]), .S(S[64]), .CO(
        C[65]) );
  FA_3804 \FAINST[65].FA_  ( .A(A[65]), .B(B[65]), .CI(C[65]), .S(S[65]), .CO(
        C[66]) );
  FA_3803 \FAINST[66].FA_  ( .A(A[66]), .B(B[66]), .CI(C[66]), .S(S[66]), .CO(
        C[67]) );
  FA_3802 \FAINST[67].FA_  ( .A(A[67]), .B(B[67]), .CI(C[67]), .S(S[67]), .CO(
        C[68]) );
  FA_3801 \FAINST[68].FA_  ( .A(A[68]), .B(B[68]), .CI(C[68]), .S(S[68]), .CO(
        C[69]) );
  FA_3800 \FAINST[69].FA_  ( .A(A[69]), .B(B[69]), .CI(C[69]), .S(S[69]), .CO(
        C[70]) );
  FA_3799 \FAINST[70].FA_  ( .A(A[70]), .B(B[70]), .CI(C[70]), .S(S[70]), .CO(
        C[71]) );
  FA_3798 \FAINST[71].FA_  ( .A(A[71]), .B(B[71]), .CI(C[71]), .S(S[71]), .CO(
        C[72]) );
  FA_3797 \FAINST[72].FA_  ( .A(A[72]), .B(B[72]), .CI(C[72]), .S(S[72]), .CO(
        C[73]) );
  FA_3796 \FAINST[73].FA_  ( .A(A[73]), .B(B[73]), .CI(C[73]), .S(S[73]), .CO(
        C[74]) );
  FA_3795 \FAINST[74].FA_  ( .A(A[74]), .B(B[74]), .CI(C[74]), .S(S[74]), .CO(
        C[75]) );
  FA_3794 \FAINST[75].FA_  ( .A(A[75]), .B(B[75]), .CI(C[75]), .S(S[75]), .CO(
        C[76]) );
  FA_3793 \FAINST[76].FA_  ( .A(A[76]), .B(B[76]), .CI(C[76]), .S(S[76]), .CO(
        C[77]) );
  FA_3792 \FAINST[77].FA_  ( .A(A[77]), .B(B[77]), .CI(C[77]), .S(S[77]), .CO(
        C[78]) );
  FA_3791 \FAINST[78].FA_  ( .A(A[78]), .B(B[78]), .CI(C[78]), .S(S[78]), .CO(
        C[79]) );
  FA_3790 \FAINST[79].FA_  ( .A(A[79]), .B(B[79]), .CI(C[79]), .S(S[79]), .CO(
        C[80]) );
  FA_3789 \FAINST[80].FA_  ( .A(A[80]), .B(B[80]), .CI(C[80]), .S(S[80]), .CO(
        C[81]) );
  FA_3788 \FAINST[81].FA_  ( .A(A[81]), .B(B[81]), .CI(C[81]), .S(S[81]), .CO(
        C[82]) );
  FA_3787 \FAINST[82].FA_  ( .A(A[82]), .B(B[82]), .CI(C[82]), .S(S[82]), .CO(
        C[83]) );
  FA_3786 \FAINST[83].FA_  ( .A(A[83]), .B(B[83]), .CI(C[83]), .S(S[83]), .CO(
        C[84]) );
  FA_3785 \FAINST[84].FA_  ( .A(A[84]), .B(B[84]), .CI(C[84]), .S(S[84]), .CO(
        C[85]) );
  FA_3784 \FAINST[85].FA_  ( .A(A[85]), .B(B[85]), .CI(C[85]), .S(S[85]), .CO(
        C[86]) );
  FA_3783 \FAINST[86].FA_  ( .A(A[86]), .B(B[86]), .CI(C[86]), .S(S[86]), .CO(
        C[87]) );
  FA_3782 \FAINST[87].FA_  ( .A(A[87]), .B(B[87]), .CI(C[87]), .S(S[87]), .CO(
        C[88]) );
  FA_3781 \FAINST[88].FA_  ( .A(A[88]), .B(B[88]), .CI(C[88]), .S(S[88]), .CO(
        C[89]) );
  FA_3780 \FAINST[89].FA_  ( .A(A[89]), .B(B[89]), .CI(C[89]), .S(S[89]), .CO(
        C[90]) );
  FA_3779 \FAINST[90].FA_  ( .A(A[90]), .B(B[90]), .CI(C[90]), .S(S[90]), .CO(
        C[91]) );
  FA_3778 \FAINST[91].FA_  ( .A(A[91]), .B(B[91]), .CI(C[91]), .S(S[91]), .CO(
        C[92]) );
  FA_3777 \FAINST[92].FA_  ( .A(A[92]), .B(B[92]), .CI(C[92]), .S(S[92]), .CO(
        C[93]) );
  FA_3776 \FAINST[93].FA_  ( .A(A[93]), .B(B[93]), .CI(C[93]), .S(S[93]), .CO(
        C[94]) );
  FA_3775 \FAINST[94].FA_  ( .A(A[94]), .B(B[94]), .CI(C[94]), .S(S[94]), .CO(
        C[95]) );
  FA_3774 \FAINST[95].FA_  ( .A(A[95]), .B(B[95]), .CI(C[95]), .S(S[95]), .CO(
        C[96]) );
  FA_3773 \FAINST[96].FA_  ( .A(A[96]), .B(B[96]), .CI(C[96]), .S(S[96]), .CO(
        C[97]) );
  FA_3772 \FAINST[97].FA_  ( .A(A[97]), .B(B[97]), .CI(C[97]), .S(S[97]), .CO(
        C[98]) );
  FA_3771 \FAINST[98].FA_  ( .A(A[98]), .B(B[98]), .CI(C[98]), .S(S[98]), .CO(
        C[99]) );
  FA_3770 \FAINST[99].FA_  ( .A(A[99]), .B(B[99]), .CI(C[99]), .S(S[99]), .CO(
        C[100]) );
  FA_3769 \FAINST[100].FA_  ( .A(A[100]), .B(B[100]), .CI(C[100]), .S(S[100]), 
        .CO(C[101]) );
  FA_3768 \FAINST[101].FA_  ( .A(A[101]), .B(B[101]), .CI(C[101]), .S(S[101]), 
        .CO(C[102]) );
  FA_3767 \FAINST[102].FA_  ( .A(A[102]), .B(B[102]), .CI(C[102]), .S(S[102]), 
        .CO(C[103]) );
  FA_3766 \FAINST[103].FA_  ( .A(A[103]), .B(B[103]), .CI(C[103]), .S(S[103]), 
        .CO(C[104]) );
  FA_3765 \FAINST[104].FA_  ( .A(A[104]), .B(B[104]), .CI(C[104]), .S(S[104]), 
        .CO(C[105]) );
  FA_3764 \FAINST[105].FA_  ( .A(A[105]), .B(B[105]), .CI(C[105]), .S(S[105]), 
        .CO(C[106]) );
  FA_3763 \FAINST[106].FA_  ( .A(A[106]), .B(B[106]), .CI(C[106]), .S(S[106]), 
        .CO(C[107]) );
  FA_3762 \FAINST[107].FA_  ( .A(A[107]), .B(B[107]), .CI(C[107]), .S(S[107]), 
        .CO(C[108]) );
  FA_3761 \FAINST[108].FA_  ( .A(A[108]), .B(B[108]), .CI(C[108]), .S(S[108]), 
        .CO(C[109]) );
  FA_3760 \FAINST[109].FA_  ( .A(A[109]), .B(B[109]), .CI(C[109]), .S(S[109]), 
        .CO(C[110]) );
  FA_3759 \FAINST[110].FA_  ( .A(A[110]), .B(B[110]), .CI(C[110]), .S(S[110]), 
        .CO(C[111]) );
  FA_3758 \FAINST[111].FA_  ( .A(A[111]), .B(B[111]), .CI(C[111]), .S(S[111]), 
        .CO(C[112]) );
  FA_3757 \FAINST[112].FA_  ( .A(A[112]), .B(B[112]), .CI(C[112]), .S(S[112]), 
        .CO(C[113]) );
  FA_3756 \FAINST[113].FA_  ( .A(A[113]), .B(B[113]), .CI(C[113]), .S(S[113]), 
        .CO(C[114]) );
  FA_3755 \FAINST[114].FA_  ( .A(A[114]), .B(B[114]), .CI(C[114]), .S(S[114]), 
        .CO(C[115]) );
  FA_3754 \FAINST[115].FA_  ( .A(A[115]), .B(B[115]), .CI(C[115]), .S(S[115]), 
        .CO(C[116]) );
  FA_3753 \FAINST[116].FA_  ( .A(A[116]), .B(B[116]), .CI(C[116]), .S(S[116]), 
        .CO(C[117]) );
  FA_3752 \FAINST[117].FA_  ( .A(A[117]), .B(B[117]), .CI(C[117]), .S(S[117]), 
        .CO(C[118]) );
  FA_3751 \FAINST[118].FA_  ( .A(A[118]), .B(B[118]), .CI(C[118]), .S(S[118]), 
        .CO(C[119]) );
  FA_3750 \FAINST[119].FA_  ( .A(A[119]), .B(B[119]), .CI(C[119]), .S(S[119]), 
        .CO(C[120]) );
  FA_3749 \FAINST[120].FA_  ( .A(A[120]), .B(B[120]), .CI(C[120]), .S(S[120]), 
        .CO(C[121]) );
  FA_3748 \FAINST[121].FA_  ( .A(A[121]), .B(B[121]), .CI(C[121]), .S(S[121]), 
        .CO(C[122]) );
  FA_3747 \FAINST[122].FA_  ( .A(A[122]), .B(B[122]), .CI(C[122]), .S(S[122]), 
        .CO(C[123]) );
  FA_3746 \FAINST[123].FA_  ( .A(A[123]), .B(B[123]), .CI(C[123]), .S(S[123]), 
        .CO(C[124]) );
  FA_3745 \FAINST[124].FA_  ( .A(A[124]), .B(B[124]), .CI(C[124]), .S(S[124]), 
        .CO(C[125]) );
  FA_3744 \FAINST[125].FA_  ( .A(A[125]), .B(B[125]), .CI(C[125]), .S(S[125]), 
        .CO(C[126]) );
  FA_3743 \FAINST[126].FA_  ( .A(A[126]), .B(B[126]), .CI(C[126]), .S(S[126]), 
        .CO(C[127]) );
  FA_3742 \FAINST[127].FA_  ( .A(A[127]), .B(B[127]), .CI(C[127]), .S(S[127]), 
        .CO(C[128]) );
  FA_3741 \FAINST[128].FA_  ( .A(A[128]), .B(B[128]), .CI(C[128]), .S(S[128]), 
        .CO(C[129]) );
  FA_3740 \FAINST[129].FA_  ( .A(A[129]), .B(B[129]), .CI(C[129]), .S(S[129]), 
        .CO(C[130]) );
  FA_3739 \FAINST[130].FA_  ( .A(A[130]), .B(B[130]), .CI(C[130]), .S(S[130]), 
        .CO(C[131]) );
  FA_3738 \FAINST[131].FA_  ( .A(A[131]), .B(B[131]), .CI(C[131]), .S(S[131]), 
        .CO(C[132]) );
  FA_3737 \FAINST[132].FA_  ( .A(A[132]), .B(B[132]), .CI(C[132]), .S(S[132]), 
        .CO(C[133]) );
  FA_3736 \FAINST[133].FA_  ( .A(A[133]), .B(B[133]), .CI(C[133]), .S(S[133]), 
        .CO(C[134]) );
  FA_3735 \FAINST[134].FA_  ( .A(A[134]), .B(B[134]), .CI(C[134]), .S(S[134]), 
        .CO(C[135]) );
  FA_3734 \FAINST[135].FA_  ( .A(A[135]), .B(B[135]), .CI(C[135]), .S(S[135]), 
        .CO(C[136]) );
  FA_3733 \FAINST[136].FA_  ( .A(A[136]), .B(B[136]), .CI(C[136]), .S(S[136]), 
        .CO(C[137]) );
  FA_3732 \FAINST[137].FA_  ( .A(A[137]), .B(B[137]), .CI(C[137]), .S(S[137]), 
        .CO(C[138]) );
  FA_3731 \FAINST[138].FA_  ( .A(A[138]), .B(B[138]), .CI(C[138]), .S(S[138]), 
        .CO(C[139]) );
  FA_3730 \FAINST[139].FA_  ( .A(A[139]), .B(B[139]), .CI(C[139]), .S(S[139]), 
        .CO(C[140]) );
  FA_3729 \FAINST[140].FA_  ( .A(A[140]), .B(B[140]), .CI(C[140]), .S(S[140]), 
        .CO(C[141]) );
  FA_3728 \FAINST[141].FA_  ( .A(A[141]), .B(B[141]), .CI(C[141]), .S(S[141]), 
        .CO(C[142]) );
  FA_3727 \FAINST[142].FA_  ( .A(A[142]), .B(B[142]), .CI(C[142]), .S(S[142]), 
        .CO(C[143]) );
  FA_3726 \FAINST[143].FA_  ( .A(A[143]), .B(B[143]), .CI(C[143]), .S(S[143]), 
        .CO(C[144]) );
  FA_3725 \FAINST[144].FA_  ( .A(A[144]), .B(B[144]), .CI(C[144]), .S(S[144]), 
        .CO(C[145]) );
  FA_3724 \FAINST[145].FA_  ( .A(A[145]), .B(B[145]), .CI(C[145]), .S(S[145]), 
        .CO(C[146]) );
  FA_3723 \FAINST[146].FA_  ( .A(A[146]), .B(B[146]), .CI(C[146]), .S(S[146]), 
        .CO(C[147]) );
  FA_3722 \FAINST[147].FA_  ( .A(A[147]), .B(B[147]), .CI(C[147]), .S(S[147]), 
        .CO(C[148]) );
  FA_3721 \FAINST[148].FA_  ( .A(A[148]), .B(B[148]), .CI(C[148]), .S(S[148]), 
        .CO(C[149]) );
  FA_3720 \FAINST[149].FA_  ( .A(A[149]), .B(B[149]), .CI(C[149]), .S(S[149]), 
        .CO(C[150]) );
  FA_3719 \FAINST[150].FA_  ( .A(A[150]), .B(B[150]), .CI(C[150]), .S(S[150]), 
        .CO(C[151]) );
  FA_3718 \FAINST[151].FA_  ( .A(A[151]), .B(B[151]), .CI(C[151]), .S(S[151]), 
        .CO(C[152]) );
  FA_3717 \FAINST[152].FA_  ( .A(A[152]), .B(B[152]), .CI(C[152]), .S(S[152]), 
        .CO(C[153]) );
  FA_3716 \FAINST[153].FA_  ( .A(A[153]), .B(B[153]), .CI(C[153]), .S(S[153]), 
        .CO(C[154]) );
  FA_3715 \FAINST[154].FA_  ( .A(A[154]), .B(B[154]), .CI(C[154]), .S(S[154]), 
        .CO(C[155]) );
  FA_3714 \FAINST[155].FA_  ( .A(A[155]), .B(B[155]), .CI(C[155]), .S(S[155]), 
        .CO(C[156]) );
  FA_3713 \FAINST[156].FA_  ( .A(A[156]), .B(B[156]), .CI(C[156]), .S(S[156]), 
        .CO(C[157]) );
  FA_3712 \FAINST[157].FA_  ( .A(A[157]), .B(B[157]), .CI(C[157]), .S(S[157]), 
        .CO(C[158]) );
  FA_3711 \FAINST[158].FA_  ( .A(A[158]), .B(B[158]), .CI(C[158]), .S(S[158]), 
        .CO(C[159]) );
  FA_3710 \FAINST[159].FA_  ( .A(A[159]), .B(B[159]), .CI(C[159]), .S(S[159]), 
        .CO(C[160]) );
  FA_3709 \FAINST[160].FA_  ( .A(A[160]), .B(B[160]), .CI(C[160]), .S(S[160]), 
        .CO(C[161]) );
  FA_3708 \FAINST[161].FA_  ( .A(A[161]), .B(B[161]), .CI(C[161]), .S(S[161]), 
        .CO(C[162]) );
  FA_3707 \FAINST[162].FA_  ( .A(A[162]), .B(B[162]), .CI(C[162]), .S(S[162]), 
        .CO(C[163]) );
  FA_3706 \FAINST[163].FA_  ( .A(A[163]), .B(B[163]), .CI(C[163]), .S(S[163]), 
        .CO(C[164]) );
  FA_3705 \FAINST[164].FA_  ( .A(A[164]), .B(B[164]), .CI(C[164]), .S(S[164]), 
        .CO(C[165]) );
  FA_3704 \FAINST[165].FA_  ( .A(A[165]), .B(B[165]), .CI(C[165]), .S(S[165]), 
        .CO(C[166]) );
  FA_3703 \FAINST[166].FA_  ( .A(A[166]), .B(B[166]), .CI(C[166]), .S(S[166]), 
        .CO(C[167]) );
  FA_3702 \FAINST[167].FA_  ( .A(A[167]), .B(B[167]), .CI(C[167]), .S(S[167]), 
        .CO(C[168]) );
  FA_3701 \FAINST[168].FA_  ( .A(A[168]), .B(B[168]), .CI(C[168]), .S(S[168]), 
        .CO(C[169]) );
  FA_3700 \FAINST[169].FA_  ( .A(A[169]), .B(B[169]), .CI(C[169]), .S(S[169]), 
        .CO(C[170]) );
  FA_3699 \FAINST[170].FA_  ( .A(A[170]), .B(B[170]), .CI(C[170]), .S(S[170]), 
        .CO(C[171]) );
  FA_3698 \FAINST[171].FA_  ( .A(A[171]), .B(B[171]), .CI(C[171]), .S(S[171]), 
        .CO(C[172]) );
  FA_3697 \FAINST[172].FA_  ( .A(A[172]), .B(B[172]), .CI(C[172]), .S(S[172]), 
        .CO(C[173]) );
  FA_3696 \FAINST[173].FA_  ( .A(A[173]), .B(B[173]), .CI(C[173]), .S(S[173]), 
        .CO(C[174]) );
  FA_3695 \FAINST[174].FA_  ( .A(A[174]), .B(B[174]), .CI(C[174]), .S(S[174]), 
        .CO(C[175]) );
  FA_3694 \FAINST[175].FA_  ( .A(A[175]), .B(B[175]), .CI(C[175]), .S(S[175]), 
        .CO(C[176]) );
  FA_3693 \FAINST[176].FA_  ( .A(A[176]), .B(B[176]), .CI(C[176]), .S(S[176]), 
        .CO(C[177]) );
  FA_3692 \FAINST[177].FA_  ( .A(A[177]), .B(B[177]), .CI(C[177]), .S(S[177]), 
        .CO(C[178]) );
  FA_3691 \FAINST[178].FA_  ( .A(A[178]), .B(B[178]), .CI(C[178]), .S(S[178]), 
        .CO(C[179]) );
  FA_3690 \FAINST[179].FA_  ( .A(A[179]), .B(B[179]), .CI(C[179]), .S(S[179]), 
        .CO(C[180]) );
  FA_3689 \FAINST[180].FA_  ( .A(A[180]), .B(B[180]), .CI(C[180]), .S(S[180]), 
        .CO(C[181]) );
  FA_3688 \FAINST[181].FA_  ( .A(A[181]), .B(B[181]), .CI(C[181]), .S(S[181]), 
        .CO(C[182]) );
  FA_3687 \FAINST[182].FA_  ( .A(A[182]), .B(B[182]), .CI(C[182]), .S(S[182]), 
        .CO(C[183]) );
  FA_3686 \FAINST[183].FA_  ( .A(A[183]), .B(B[183]), .CI(C[183]), .S(S[183]), 
        .CO(C[184]) );
  FA_3685 \FAINST[184].FA_  ( .A(A[184]), .B(B[184]), .CI(C[184]), .S(S[184]), 
        .CO(C[185]) );
  FA_3684 \FAINST[185].FA_  ( .A(A[185]), .B(B[185]), .CI(C[185]), .S(S[185]), 
        .CO(C[186]) );
  FA_3683 \FAINST[186].FA_  ( .A(A[186]), .B(B[186]), .CI(C[186]), .S(S[186]), 
        .CO(C[187]) );
  FA_3682 \FAINST[187].FA_  ( .A(A[187]), .B(B[187]), .CI(C[187]), .S(S[187]), 
        .CO(C[188]) );
  FA_3681 \FAINST[188].FA_  ( .A(A[188]), .B(B[188]), .CI(C[188]), .S(S[188]), 
        .CO(C[189]) );
  FA_3680 \FAINST[189].FA_  ( .A(A[189]), .B(B[189]), .CI(C[189]), .S(S[189]), 
        .CO(C[190]) );
  FA_3679 \FAINST[190].FA_  ( .A(A[190]), .B(B[190]), .CI(C[190]), .S(S[190]), 
        .CO(C[191]) );
  FA_3678 \FAINST[191].FA_  ( .A(A[191]), .B(B[191]), .CI(C[191]), .S(S[191]), 
        .CO(C[192]) );
  FA_3677 \FAINST[192].FA_  ( .A(A[192]), .B(B[192]), .CI(C[192]), .S(S[192]), 
        .CO(C[193]) );
  FA_3676 \FAINST[193].FA_  ( .A(A[193]), .B(B[193]), .CI(C[193]), .S(S[193]), 
        .CO(C[194]) );
  FA_3675 \FAINST[194].FA_  ( .A(A[194]), .B(B[194]), .CI(C[194]), .S(S[194]), 
        .CO(C[195]) );
  FA_3674 \FAINST[195].FA_  ( .A(A[195]), .B(B[195]), .CI(C[195]), .S(S[195]), 
        .CO(C[196]) );
  FA_3673 \FAINST[196].FA_  ( .A(A[196]), .B(B[196]), .CI(C[196]), .S(S[196]), 
        .CO(C[197]) );
  FA_3672 \FAINST[197].FA_  ( .A(A[197]), .B(B[197]), .CI(C[197]), .S(S[197]), 
        .CO(C[198]) );
  FA_3671 \FAINST[198].FA_  ( .A(A[198]), .B(B[198]), .CI(C[198]), .S(S[198]), 
        .CO(C[199]) );
  FA_3670 \FAINST[199].FA_  ( .A(A[199]), .B(B[199]), .CI(C[199]), .S(S[199]), 
        .CO(C[200]) );
  FA_3669 \FAINST[200].FA_  ( .A(A[200]), .B(B[200]), .CI(C[200]), .S(S[200]), 
        .CO(C[201]) );
  FA_3668 \FAINST[201].FA_  ( .A(A[201]), .B(B[201]), .CI(C[201]), .S(S[201]), 
        .CO(C[202]) );
  FA_3667 \FAINST[202].FA_  ( .A(A[202]), .B(B[202]), .CI(C[202]), .S(S[202]), 
        .CO(C[203]) );
  FA_3666 \FAINST[203].FA_  ( .A(A[203]), .B(B[203]), .CI(C[203]), .S(S[203]), 
        .CO(C[204]) );
  FA_3665 \FAINST[204].FA_  ( .A(A[204]), .B(B[204]), .CI(C[204]), .S(S[204]), 
        .CO(C[205]) );
  FA_3664 \FAINST[205].FA_  ( .A(A[205]), .B(B[205]), .CI(C[205]), .S(S[205]), 
        .CO(C[206]) );
  FA_3663 \FAINST[206].FA_  ( .A(A[206]), .B(B[206]), .CI(C[206]), .S(S[206]), 
        .CO(C[207]) );
  FA_3662 \FAINST[207].FA_  ( .A(A[207]), .B(B[207]), .CI(C[207]), .S(S[207]), 
        .CO(C[208]) );
  FA_3661 \FAINST[208].FA_  ( .A(A[208]), .B(B[208]), .CI(C[208]), .S(S[208]), 
        .CO(C[209]) );
  FA_3660 \FAINST[209].FA_  ( .A(A[209]), .B(B[209]), .CI(C[209]), .S(S[209]), 
        .CO(C[210]) );
  FA_3659 \FAINST[210].FA_  ( .A(A[210]), .B(B[210]), .CI(C[210]), .S(S[210]), 
        .CO(C[211]) );
  FA_3658 \FAINST[211].FA_  ( .A(A[211]), .B(B[211]), .CI(C[211]), .S(S[211]), 
        .CO(C[212]) );
  FA_3657 \FAINST[212].FA_  ( .A(A[212]), .B(B[212]), .CI(C[212]), .S(S[212]), 
        .CO(C[213]) );
  FA_3656 \FAINST[213].FA_  ( .A(A[213]), .B(B[213]), .CI(C[213]), .S(S[213]), 
        .CO(C[214]) );
  FA_3655 \FAINST[214].FA_  ( .A(A[214]), .B(B[214]), .CI(C[214]), .S(S[214]), 
        .CO(C[215]) );
  FA_3654 \FAINST[215].FA_  ( .A(A[215]), .B(B[215]), .CI(C[215]), .S(S[215]), 
        .CO(C[216]) );
  FA_3653 \FAINST[216].FA_  ( .A(A[216]), .B(B[216]), .CI(C[216]), .S(S[216]), 
        .CO(C[217]) );
  FA_3652 \FAINST[217].FA_  ( .A(A[217]), .B(B[217]), .CI(C[217]), .S(S[217]), 
        .CO(C[218]) );
  FA_3651 \FAINST[218].FA_  ( .A(A[218]), .B(B[218]), .CI(C[218]), .S(S[218]), 
        .CO(C[219]) );
  FA_3650 \FAINST[219].FA_  ( .A(A[219]), .B(B[219]), .CI(C[219]), .S(S[219]), 
        .CO(C[220]) );
  FA_3649 \FAINST[220].FA_  ( .A(A[220]), .B(B[220]), .CI(C[220]), .S(S[220]), 
        .CO(C[221]) );
  FA_3648 \FAINST[221].FA_  ( .A(A[221]), .B(B[221]), .CI(C[221]), .S(S[221]), 
        .CO(C[222]) );
  FA_3647 \FAINST[222].FA_  ( .A(A[222]), .B(B[222]), .CI(C[222]), .S(S[222]), 
        .CO(C[223]) );
  FA_3646 \FAINST[223].FA_  ( .A(A[223]), .B(B[223]), .CI(C[223]), .S(S[223]), 
        .CO(C[224]) );
  FA_3645 \FAINST[224].FA_  ( .A(A[224]), .B(B[224]), .CI(C[224]), .S(S[224]), 
        .CO(C[225]) );
  FA_3644 \FAINST[225].FA_  ( .A(A[225]), .B(B[225]), .CI(C[225]), .S(S[225]), 
        .CO(C[226]) );
  FA_3643 \FAINST[226].FA_  ( .A(A[226]), .B(B[226]), .CI(C[226]), .S(S[226]), 
        .CO(C[227]) );
  FA_3642 \FAINST[227].FA_  ( .A(A[227]), .B(B[227]), .CI(C[227]), .S(S[227]), 
        .CO(C[228]) );
  FA_3641 \FAINST[228].FA_  ( .A(A[228]), .B(B[228]), .CI(C[228]), .S(S[228]), 
        .CO(C[229]) );
  FA_3640 \FAINST[229].FA_  ( .A(A[229]), .B(B[229]), .CI(C[229]), .S(S[229]), 
        .CO(C[230]) );
  FA_3639 \FAINST[230].FA_  ( .A(A[230]), .B(B[230]), .CI(C[230]), .S(S[230]), 
        .CO(C[231]) );
  FA_3638 \FAINST[231].FA_  ( .A(A[231]), .B(B[231]), .CI(C[231]), .S(S[231]), 
        .CO(C[232]) );
  FA_3637 \FAINST[232].FA_  ( .A(A[232]), .B(B[232]), .CI(C[232]), .S(S[232]), 
        .CO(C[233]) );
  FA_3636 \FAINST[233].FA_  ( .A(A[233]), .B(B[233]), .CI(C[233]), .S(S[233]), 
        .CO(C[234]) );
  FA_3635 \FAINST[234].FA_  ( .A(A[234]), .B(B[234]), .CI(C[234]), .S(S[234]), 
        .CO(C[235]) );
  FA_3634 \FAINST[235].FA_  ( .A(A[235]), .B(B[235]), .CI(C[235]), .S(S[235]), 
        .CO(C[236]) );
  FA_3633 \FAINST[236].FA_  ( .A(A[236]), .B(B[236]), .CI(C[236]), .S(S[236]), 
        .CO(C[237]) );
  FA_3632 \FAINST[237].FA_  ( .A(A[237]), .B(B[237]), .CI(C[237]), .S(S[237]), 
        .CO(C[238]) );
  FA_3631 \FAINST[238].FA_  ( .A(A[238]), .B(B[238]), .CI(C[238]), .S(S[238]), 
        .CO(C[239]) );
  FA_3630 \FAINST[239].FA_  ( .A(A[239]), .B(B[239]), .CI(C[239]), .S(S[239]), 
        .CO(C[240]) );
  FA_3629 \FAINST[240].FA_  ( .A(A[240]), .B(B[240]), .CI(C[240]), .S(S[240]), 
        .CO(C[241]) );
  FA_3628 \FAINST[241].FA_  ( .A(A[241]), .B(B[241]), .CI(C[241]), .S(S[241]), 
        .CO(C[242]) );
  FA_3627 \FAINST[242].FA_  ( .A(A[242]), .B(B[242]), .CI(C[242]), .S(S[242]), 
        .CO(C[243]) );
  FA_3626 \FAINST[243].FA_  ( .A(A[243]), .B(B[243]), .CI(C[243]), .S(S[243]), 
        .CO(C[244]) );
  FA_3625 \FAINST[244].FA_  ( .A(A[244]), .B(B[244]), .CI(C[244]), .S(S[244]), 
        .CO(C[245]) );
  FA_3624 \FAINST[245].FA_  ( .A(A[245]), .B(B[245]), .CI(C[245]), .S(S[245]), 
        .CO(C[246]) );
  FA_3623 \FAINST[246].FA_  ( .A(A[246]), .B(B[246]), .CI(C[246]), .S(S[246]), 
        .CO(C[247]) );
  FA_3622 \FAINST[247].FA_  ( .A(A[247]), .B(B[247]), .CI(C[247]), .S(S[247]), 
        .CO(C[248]) );
  FA_3621 \FAINST[248].FA_  ( .A(A[248]), .B(B[248]), .CI(C[248]), .S(S[248]), 
        .CO(C[249]) );
  FA_3620 \FAINST[249].FA_  ( .A(A[249]), .B(B[249]), .CI(C[249]), .S(S[249]), 
        .CO(C[250]) );
  FA_3619 \FAINST[250].FA_  ( .A(A[250]), .B(B[250]), .CI(C[250]), .S(S[250]), 
        .CO(C[251]) );
  FA_3618 \FAINST[251].FA_  ( .A(A[251]), .B(B[251]), .CI(C[251]), .S(S[251]), 
        .CO(C[252]) );
  FA_3617 \FAINST[252].FA_  ( .A(A[252]), .B(B[252]), .CI(C[252]), .S(S[252]), 
        .CO(C[253]) );
  FA_3616 \FAINST[253].FA_  ( .A(A[253]), .B(B[253]), .CI(C[253]), .S(S[253]), 
        .CO(C[254]) );
  FA_3615 \FAINST[254].FA_  ( .A(A[254]), .B(B[254]), .CI(C[254]), .S(S[254]), 
        .CO(C[255]) );
  FA_3614 \FAINST[255].FA_  ( .A(A[255]), .B(B[255]), .CI(C[255]), .S(S[255]), 
        .CO(C[256]) );
  FA_3613 \FAINST[256].FA_  ( .A(A[256]), .B(1'b0), .CI(C[256]), .S(S[256]), 
        .CO(C[257]) );
  FA_3612 \FAINST[257].FA_  ( .A(A[257]), .B(1'b0), .CI(C[257]), .S(S[257]) );
endmodule


module FA_3354 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  OR U1 ( .A(CI), .B(A), .Z(CO) );
endmodule


module FA_3355 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  OR U1 ( .A(CI), .B(A), .Z(CO) );
endmodule


module FA_3356 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3357 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3358 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3359 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3360 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3361 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3362 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3363 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3364 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3365 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3366 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3367 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3368 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3369 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3370 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3371 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3372 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3373 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3374 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3375 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3376 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3377 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3378 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3379 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3380 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3381 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3382 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3383 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3384 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3385 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3386 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3387 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3388 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3389 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3390 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3391 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3392 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3393 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3394 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3395 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3396 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3397 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3398 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3399 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3400 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3401 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3402 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3403 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3404 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3405 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3406 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3407 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3408 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3409 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3410 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3411 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3412 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3413 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3414 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3415 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3416 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3417 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3418 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3419 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3420 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3421 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3422 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3423 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3424 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3425 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3426 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3427 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3428 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3429 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3430 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3431 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3432 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3433 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3434 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3435 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3436 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3437 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3438 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3439 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3440 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3441 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3442 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3443 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3444 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3445 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3446 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3447 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3448 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3449 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3450 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3451 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3452 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3453 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3454 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3455 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3456 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3457 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3458 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3459 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3460 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3461 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3462 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3463 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3464 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3465 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3466 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3467 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3468 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3469 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3470 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3471 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3472 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3473 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3474 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3475 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3476 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3477 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3478 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3479 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3480 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3481 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3482 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3483 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3484 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3485 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3486 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3487 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3488 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3489 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3490 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3491 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3492 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3493 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3494 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3495 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3496 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3497 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3498 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3499 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3500 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3501 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3502 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3503 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3504 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3505 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3506 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3507 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3508 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3509 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3510 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3511 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3512 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3513 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3514 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3515 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3516 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3517 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3518 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3519 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3520 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3521 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3522 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3523 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3524 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3525 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3526 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3527 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3528 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3529 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3530 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3531 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3532 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3533 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3534 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3535 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3536 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3537 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3538 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3539 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3540 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3541 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3542 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3543 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3544 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3545 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3546 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3547 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3548 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3549 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3550 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3551 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3552 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3553 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3554 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3555 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3556 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3557 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3558 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3559 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3560 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3561 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3562 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3563 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3564 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3565 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3566 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3567 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3568 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3569 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3570 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3571 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3572 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3573 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3574 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3575 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3576 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3577 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3578 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3579 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3580 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3581 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3582 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3583 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3584 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3585 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3586 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3587 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3588 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3589 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3590 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3591 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3592 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3593 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3594 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3595 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3596 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3597 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3598 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3599 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3600 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3601 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3602 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3603 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3604 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3605 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3606 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3607 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3608 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3609 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3610 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3611 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  OR U1 ( .A(B), .B(A), .Z(CO) );
endmodule


module COMP_N258_2 ( A, B, O );
  input [257:0] A;
  input [257:0] B;
  output O;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258;
  wire   [257:1] C;

  FA_3611 \FAINST[0].FA_  ( .A(A[0]), .B(n258), .CI(1'b1), .CO(C[1]) );
  FA_3610 \FAINST[1].FA_  ( .A(A[1]), .B(n257), .CI(C[1]), .CO(C[2]) );
  FA_3609 \FAINST[2].FA_  ( .A(A[2]), .B(n256), .CI(C[2]), .CO(C[3]) );
  FA_3608 \FAINST[3].FA_  ( .A(A[3]), .B(n255), .CI(C[3]), .CO(C[4]) );
  FA_3607 \FAINST[4].FA_  ( .A(A[4]), .B(n254), .CI(C[4]), .CO(C[5]) );
  FA_3606 \FAINST[5].FA_  ( .A(A[5]), .B(n253), .CI(C[5]), .CO(C[6]) );
  FA_3605 \FAINST[6].FA_  ( .A(A[6]), .B(n252), .CI(C[6]), .CO(C[7]) );
  FA_3604 \FAINST[7].FA_  ( .A(A[7]), .B(n251), .CI(C[7]), .CO(C[8]) );
  FA_3603 \FAINST[8].FA_  ( .A(A[8]), .B(n250), .CI(C[8]), .CO(C[9]) );
  FA_3602 \FAINST[9].FA_  ( .A(A[9]), .B(n249), .CI(C[9]), .CO(C[10]) );
  FA_3601 \FAINST[10].FA_  ( .A(A[10]), .B(n248), .CI(C[10]), .CO(C[11]) );
  FA_3600 \FAINST[11].FA_  ( .A(A[11]), .B(n247), .CI(C[11]), .CO(C[12]) );
  FA_3599 \FAINST[12].FA_  ( .A(A[12]), .B(n246), .CI(C[12]), .CO(C[13]) );
  FA_3598 \FAINST[13].FA_  ( .A(A[13]), .B(n245), .CI(C[13]), .CO(C[14]) );
  FA_3597 \FAINST[14].FA_  ( .A(A[14]), .B(n244), .CI(C[14]), .CO(C[15]) );
  FA_3596 \FAINST[15].FA_  ( .A(A[15]), .B(n243), .CI(C[15]), .CO(C[16]) );
  FA_3595 \FAINST[16].FA_  ( .A(A[16]), .B(n242), .CI(C[16]), .CO(C[17]) );
  FA_3594 \FAINST[17].FA_  ( .A(A[17]), .B(n241), .CI(C[17]), .CO(C[18]) );
  FA_3593 \FAINST[18].FA_  ( .A(A[18]), .B(n240), .CI(C[18]), .CO(C[19]) );
  FA_3592 \FAINST[19].FA_  ( .A(A[19]), .B(n239), .CI(C[19]), .CO(C[20]) );
  FA_3591 \FAINST[20].FA_  ( .A(A[20]), .B(n238), .CI(C[20]), .CO(C[21]) );
  FA_3590 \FAINST[21].FA_  ( .A(A[21]), .B(n237), .CI(C[21]), .CO(C[22]) );
  FA_3589 \FAINST[22].FA_  ( .A(A[22]), .B(n236), .CI(C[22]), .CO(C[23]) );
  FA_3588 \FAINST[23].FA_  ( .A(A[23]), .B(n235), .CI(C[23]), .CO(C[24]) );
  FA_3587 \FAINST[24].FA_  ( .A(A[24]), .B(n234), .CI(C[24]), .CO(C[25]) );
  FA_3586 \FAINST[25].FA_  ( .A(A[25]), .B(n233), .CI(C[25]), .CO(C[26]) );
  FA_3585 \FAINST[26].FA_  ( .A(A[26]), .B(n232), .CI(C[26]), .CO(C[27]) );
  FA_3584 \FAINST[27].FA_  ( .A(A[27]), .B(n231), .CI(C[27]), .CO(C[28]) );
  FA_3583 \FAINST[28].FA_  ( .A(A[28]), .B(n230), .CI(C[28]), .CO(C[29]) );
  FA_3582 \FAINST[29].FA_  ( .A(A[29]), .B(n229), .CI(C[29]), .CO(C[30]) );
  FA_3581 \FAINST[30].FA_  ( .A(A[30]), .B(n228), .CI(C[30]), .CO(C[31]) );
  FA_3580 \FAINST[31].FA_  ( .A(A[31]), .B(n227), .CI(C[31]), .CO(C[32]) );
  FA_3579 \FAINST[32].FA_  ( .A(A[32]), .B(n226), .CI(C[32]), .CO(C[33]) );
  FA_3578 \FAINST[33].FA_  ( .A(A[33]), .B(n225), .CI(C[33]), .CO(C[34]) );
  FA_3577 \FAINST[34].FA_  ( .A(A[34]), .B(n224), .CI(C[34]), .CO(C[35]) );
  FA_3576 \FAINST[35].FA_  ( .A(A[35]), .B(n223), .CI(C[35]), .CO(C[36]) );
  FA_3575 \FAINST[36].FA_  ( .A(A[36]), .B(n222), .CI(C[36]), .CO(C[37]) );
  FA_3574 \FAINST[37].FA_  ( .A(A[37]), .B(n221), .CI(C[37]), .CO(C[38]) );
  FA_3573 \FAINST[38].FA_  ( .A(A[38]), .B(n220), .CI(C[38]), .CO(C[39]) );
  FA_3572 \FAINST[39].FA_  ( .A(A[39]), .B(n219), .CI(C[39]), .CO(C[40]) );
  FA_3571 \FAINST[40].FA_  ( .A(A[40]), .B(n218), .CI(C[40]), .CO(C[41]) );
  FA_3570 \FAINST[41].FA_  ( .A(A[41]), .B(n217), .CI(C[41]), .CO(C[42]) );
  FA_3569 \FAINST[42].FA_  ( .A(A[42]), .B(n216), .CI(C[42]), .CO(C[43]) );
  FA_3568 \FAINST[43].FA_  ( .A(A[43]), .B(n215), .CI(C[43]), .CO(C[44]) );
  FA_3567 \FAINST[44].FA_  ( .A(A[44]), .B(n214), .CI(C[44]), .CO(C[45]) );
  FA_3566 \FAINST[45].FA_  ( .A(A[45]), .B(n213), .CI(C[45]), .CO(C[46]) );
  FA_3565 \FAINST[46].FA_  ( .A(A[46]), .B(n212), .CI(C[46]), .CO(C[47]) );
  FA_3564 \FAINST[47].FA_  ( .A(A[47]), .B(n211), .CI(C[47]), .CO(C[48]) );
  FA_3563 \FAINST[48].FA_  ( .A(A[48]), .B(n210), .CI(C[48]), .CO(C[49]) );
  FA_3562 \FAINST[49].FA_  ( .A(A[49]), .B(n209), .CI(C[49]), .CO(C[50]) );
  FA_3561 \FAINST[50].FA_  ( .A(A[50]), .B(n208), .CI(C[50]), .CO(C[51]) );
  FA_3560 \FAINST[51].FA_  ( .A(A[51]), .B(n207), .CI(C[51]), .CO(C[52]) );
  FA_3559 \FAINST[52].FA_  ( .A(A[52]), .B(n206), .CI(C[52]), .CO(C[53]) );
  FA_3558 \FAINST[53].FA_  ( .A(A[53]), .B(n205), .CI(C[53]), .CO(C[54]) );
  FA_3557 \FAINST[54].FA_  ( .A(A[54]), .B(n204), .CI(C[54]), .CO(C[55]) );
  FA_3556 \FAINST[55].FA_  ( .A(A[55]), .B(n203), .CI(C[55]), .CO(C[56]) );
  FA_3555 \FAINST[56].FA_  ( .A(A[56]), .B(n202), .CI(C[56]), .CO(C[57]) );
  FA_3554 \FAINST[57].FA_  ( .A(A[57]), .B(n201), .CI(C[57]), .CO(C[58]) );
  FA_3553 \FAINST[58].FA_  ( .A(A[58]), .B(n200), .CI(C[58]), .CO(C[59]) );
  FA_3552 \FAINST[59].FA_  ( .A(A[59]), .B(n199), .CI(C[59]), .CO(C[60]) );
  FA_3551 \FAINST[60].FA_  ( .A(A[60]), .B(n198), .CI(C[60]), .CO(C[61]) );
  FA_3550 \FAINST[61].FA_  ( .A(A[61]), .B(n197), .CI(C[61]), .CO(C[62]) );
  FA_3549 \FAINST[62].FA_  ( .A(A[62]), .B(n196), .CI(C[62]), .CO(C[63]) );
  FA_3548 \FAINST[63].FA_  ( .A(A[63]), .B(n195), .CI(C[63]), .CO(C[64]) );
  FA_3547 \FAINST[64].FA_  ( .A(A[64]), .B(n194), .CI(C[64]), .CO(C[65]) );
  FA_3546 \FAINST[65].FA_  ( .A(A[65]), .B(n193), .CI(C[65]), .CO(C[66]) );
  FA_3545 \FAINST[66].FA_  ( .A(A[66]), .B(n192), .CI(C[66]), .CO(C[67]) );
  FA_3544 \FAINST[67].FA_  ( .A(A[67]), .B(n191), .CI(C[67]), .CO(C[68]) );
  FA_3543 \FAINST[68].FA_  ( .A(A[68]), .B(n190), .CI(C[68]), .CO(C[69]) );
  FA_3542 \FAINST[69].FA_  ( .A(A[69]), .B(n189), .CI(C[69]), .CO(C[70]) );
  FA_3541 \FAINST[70].FA_  ( .A(A[70]), .B(n188), .CI(C[70]), .CO(C[71]) );
  FA_3540 \FAINST[71].FA_  ( .A(A[71]), .B(n187), .CI(C[71]), .CO(C[72]) );
  FA_3539 \FAINST[72].FA_  ( .A(A[72]), .B(n186), .CI(C[72]), .CO(C[73]) );
  FA_3538 \FAINST[73].FA_  ( .A(A[73]), .B(n185), .CI(C[73]), .CO(C[74]) );
  FA_3537 \FAINST[74].FA_  ( .A(A[74]), .B(n184), .CI(C[74]), .CO(C[75]) );
  FA_3536 \FAINST[75].FA_  ( .A(A[75]), .B(n183), .CI(C[75]), .CO(C[76]) );
  FA_3535 \FAINST[76].FA_  ( .A(A[76]), .B(n182), .CI(C[76]), .CO(C[77]) );
  FA_3534 \FAINST[77].FA_  ( .A(A[77]), .B(n181), .CI(C[77]), .CO(C[78]) );
  FA_3533 \FAINST[78].FA_  ( .A(A[78]), .B(n180), .CI(C[78]), .CO(C[79]) );
  FA_3532 \FAINST[79].FA_  ( .A(A[79]), .B(n179), .CI(C[79]), .CO(C[80]) );
  FA_3531 \FAINST[80].FA_  ( .A(A[80]), .B(n178), .CI(C[80]), .CO(C[81]) );
  FA_3530 \FAINST[81].FA_  ( .A(A[81]), .B(n177), .CI(C[81]), .CO(C[82]) );
  FA_3529 \FAINST[82].FA_  ( .A(A[82]), .B(n176), .CI(C[82]), .CO(C[83]) );
  FA_3528 \FAINST[83].FA_  ( .A(A[83]), .B(n175), .CI(C[83]), .CO(C[84]) );
  FA_3527 \FAINST[84].FA_  ( .A(A[84]), .B(n174), .CI(C[84]), .CO(C[85]) );
  FA_3526 \FAINST[85].FA_  ( .A(A[85]), .B(n173), .CI(C[85]), .CO(C[86]) );
  FA_3525 \FAINST[86].FA_  ( .A(A[86]), .B(n172), .CI(C[86]), .CO(C[87]) );
  FA_3524 \FAINST[87].FA_  ( .A(A[87]), .B(n171), .CI(C[87]), .CO(C[88]) );
  FA_3523 \FAINST[88].FA_  ( .A(A[88]), .B(n170), .CI(C[88]), .CO(C[89]) );
  FA_3522 \FAINST[89].FA_  ( .A(A[89]), .B(n169), .CI(C[89]), .CO(C[90]) );
  FA_3521 \FAINST[90].FA_  ( .A(A[90]), .B(n168), .CI(C[90]), .CO(C[91]) );
  FA_3520 \FAINST[91].FA_  ( .A(A[91]), .B(n167), .CI(C[91]), .CO(C[92]) );
  FA_3519 \FAINST[92].FA_  ( .A(A[92]), .B(n166), .CI(C[92]), .CO(C[93]) );
  FA_3518 \FAINST[93].FA_  ( .A(A[93]), .B(n165), .CI(C[93]), .CO(C[94]) );
  FA_3517 \FAINST[94].FA_  ( .A(A[94]), .B(n164), .CI(C[94]), .CO(C[95]) );
  FA_3516 \FAINST[95].FA_  ( .A(A[95]), .B(n163), .CI(C[95]), .CO(C[96]) );
  FA_3515 \FAINST[96].FA_  ( .A(A[96]), .B(n162), .CI(C[96]), .CO(C[97]) );
  FA_3514 \FAINST[97].FA_  ( .A(A[97]), .B(n161), .CI(C[97]), .CO(C[98]) );
  FA_3513 \FAINST[98].FA_  ( .A(A[98]), .B(n160), .CI(C[98]), .CO(C[99]) );
  FA_3512 \FAINST[99].FA_  ( .A(A[99]), .B(n159), .CI(C[99]), .CO(C[100]) );
  FA_3511 \FAINST[100].FA_  ( .A(A[100]), .B(n158), .CI(C[100]), .CO(C[101])
         );
  FA_3510 \FAINST[101].FA_  ( .A(A[101]), .B(n157), .CI(C[101]), .CO(C[102])
         );
  FA_3509 \FAINST[102].FA_  ( .A(A[102]), .B(n156), .CI(C[102]), .CO(C[103])
         );
  FA_3508 \FAINST[103].FA_  ( .A(A[103]), .B(n155), .CI(C[103]), .CO(C[104])
         );
  FA_3507 \FAINST[104].FA_  ( .A(A[104]), .B(n154), .CI(C[104]), .CO(C[105])
         );
  FA_3506 \FAINST[105].FA_  ( .A(A[105]), .B(n153), .CI(C[105]), .CO(C[106])
         );
  FA_3505 \FAINST[106].FA_  ( .A(A[106]), .B(n152), .CI(C[106]), .CO(C[107])
         );
  FA_3504 \FAINST[107].FA_  ( .A(A[107]), .B(n151), .CI(C[107]), .CO(C[108])
         );
  FA_3503 \FAINST[108].FA_  ( .A(A[108]), .B(n150), .CI(C[108]), .CO(C[109])
         );
  FA_3502 \FAINST[109].FA_  ( .A(A[109]), .B(n149), .CI(C[109]), .CO(C[110])
         );
  FA_3501 \FAINST[110].FA_  ( .A(A[110]), .B(n148), .CI(C[110]), .CO(C[111])
         );
  FA_3500 \FAINST[111].FA_  ( .A(A[111]), .B(n147), .CI(C[111]), .CO(C[112])
         );
  FA_3499 \FAINST[112].FA_  ( .A(A[112]), .B(n146), .CI(C[112]), .CO(C[113])
         );
  FA_3498 \FAINST[113].FA_  ( .A(A[113]), .B(n145), .CI(C[113]), .CO(C[114])
         );
  FA_3497 \FAINST[114].FA_  ( .A(A[114]), .B(n144), .CI(C[114]), .CO(C[115])
         );
  FA_3496 \FAINST[115].FA_  ( .A(A[115]), .B(n143), .CI(C[115]), .CO(C[116])
         );
  FA_3495 \FAINST[116].FA_  ( .A(A[116]), .B(n142), .CI(C[116]), .CO(C[117])
         );
  FA_3494 \FAINST[117].FA_  ( .A(A[117]), .B(n141), .CI(C[117]), .CO(C[118])
         );
  FA_3493 \FAINST[118].FA_  ( .A(A[118]), .B(n140), .CI(C[118]), .CO(C[119])
         );
  FA_3492 \FAINST[119].FA_  ( .A(A[119]), .B(n139), .CI(C[119]), .CO(C[120])
         );
  FA_3491 \FAINST[120].FA_  ( .A(A[120]), .B(n138), .CI(C[120]), .CO(C[121])
         );
  FA_3490 \FAINST[121].FA_  ( .A(A[121]), .B(n137), .CI(C[121]), .CO(C[122])
         );
  FA_3489 \FAINST[122].FA_  ( .A(A[122]), .B(n136), .CI(C[122]), .CO(C[123])
         );
  FA_3488 \FAINST[123].FA_  ( .A(A[123]), .B(n135), .CI(C[123]), .CO(C[124])
         );
  FA_3487 \FAINST[124].FA_  ( .A(A[124]), .B(n134), .CI(C[124]), .CO(C[125])
         );
  FA_3486 \FAINST[125].FA_  ( .A(A[125]), .B(n133), .CI(C[125]), .CO(C[126])
         );
  FA_3485 \FAINST[126].FA_  ( .A(A[126]), .B(n132), .CI(C[126]), .CO(C[127])
         );
  FA_3484 \FAINST[127].FA_  ( .A(A[127]), .B(n131), .CI(C[127]), .CO(C[128])
         );
  FA_3483 \FAINST[128].FA_  ( .A(A[128]), .B(n130), .CI(C[128]), .CO(C[129])
         );
  FA_3482 \FAINST[129].FA_  ( .A(A[129]), .B(n129), .CI(C[129]), .CO(C[130])
         );
  FA_3481 \FAINST[130].FA_  ( .A(A[130]), .B(n128), .CI(C[130]), .CO(C[131])
         );
  FA_3480 \FAINST[131].FA_  ( .A(A[131]), .B(n127), .CI(C[131]), .CO(C[132])
         );
  FA_3479 \FAINST[132].FA_  ( .A(A[132]), .B(n126), .CI(C[132]), .CO(C[133])
         );
  FA_3478 \FAINST[133].FA_  ( .A(A[133]), .B(n125), .CI(C[133]), .CO(C[134])
         );
  FA_3477 \FAINST[134].FA_  ( .A(A[134]), .B(n124), .CI(C[134]), .CO(C[135])
         );
  FA_3476 \FAINST[135].FA_  ( .A(A[135]), .B(n123), .CI(C[135]), .CO(C[136])
         );
  FA_3475 \FAINST[136].FA_  ( .A(A[136]), .B(n122), .CI(C[136]), .CO(C[137])
         );
  FA_3474 \FAINST[137].FA_  ( .A(A[137]), .B(n121), .CI(C[137]), .CO(C[138])
         );
  FA_3473 \FAINST[138].FA_  ( .A(A[138]), .B(n120), .CI(C[138]), .CO(C[139])
         );
  FA_3472 \FAINST[139].FA_  ( .A(A[139]), .B(n119), .CI(C[139]), .CO(C[140])
         );
  FA_3471 \FAINST[140].FA_  ( .A(A[140]), .B(n118), .CI(C[140]), .CO(C[141])
         );
  FA_3470 \FAINST[141].FA_  ( .A(A[141]), .B(n117), .CI(C[141]), .CO(C[142])
         );
  FA_3469 \FAINST[142].FA_  ( .A(A[142]), .B(n116), .CI(C[142]), .CO(C[143])
         );
  FA_3468 \FAINST[143].FA_  ( .A(A[143]), .B(n115), .CI(C[143]), .CO(C[144])
         );
  FA_3467 \FAINST[144].FA_  ( .A(A[144]), .B(n114), .CI(C[144]), .CO(C[145])
         );
  FA_3466 \FAINST[145].FA_  ( .A(A[145]), .B(n113), .CI(C[145]), .CO(C[146])
         );
  FA_3465 \FAINST[146].FA_  ( .A(A[146]), .B(n112), .CI(C[146]), .CO(C[147])
         );
  FA_3464 \FAINST[147].FA_  ( .A(A[147]), .B(n111), .CI(C[147]), .CO(C[148])
         );
  FA_3463 \FAINST[148].FA_  ( .A(A[148]), .B(n110), .CI(C[148]), .CO(C[149])
         );
  FA_3462 \FAINST[149].FA_  ( .A(A[149]), .B(n109), .CI(C[149]), .CO(C[150])
         );
  FA_3461 \FAINST[150].FA_  ( .A(A[150]), .B(n108), .CI(C[150]), .CO(C[151])
         );
  FA_3460 \FAINST[151].FA_  ( .A(A[151]), .B(n107), .CI(C[151]), .CO(C[152])
         );
  FA_3459 \FAINST[152].FA_  ( .A(A[152]), .B(n106), .CI(C[152]), .CO(C[153])
         );
  FA_3458 \FAINST[153].FA_  ( .A(A[153]), .B(n105), .CI(C[153]), .CO(C[154])
         );
  FA_3457 \FAINST[154].FA_  ( .A(A[154]), .B(n104), .CI(C[154]), .CO(C[155])
         );
  FA_3456 \FAINST[155].FA_  ( .A(A[155]), .B(n103), .CI(C[155]), .CO(C[156])
         );
  FA_3455 \FAINST[156].FA_  ( .A(A[156]), .B(n102), .CI(C[156]), .CO(C[157])
         );
  FA_3454 \FAINST[157].FA_  ( .A(A[157]), .B(n101), .CI(C[157]), .CO(C[158])
         );
  FA_3453 \FAINST[158].FA_  ( .A(A[158]), .B(n100), .CI(C[158]), .CO(C[159])
         );
  FA_3452 \FAINST[159].FA_  ( .A(A[159]), .B(n99), .CI(C[159]), .CO(C[160]) );
  FA_3451 \FAINST[160].FA_  ( .A(A[160]), .B(n98), .CI(C[160]), .CO(C[161]) );
  FA_3450 \FAINST[161].FA_  ( .A(A[161]), .B(n97), .CI(C[161]), .CO(C[162]) );
  FA_3449 \FAINST[162].FA_  ( .A(A[162]), .B(n96), .CI(C[162]), .CO(C[163]) );
  FA_3448 \FAINST[163].FA_  ( .A(A[163]), .B(n95), .CI(C[163]), .CO(C[164]) );
  FA_3447 \FAINST[164].FA_  ( .A(A[164]), .B(n94), .CI(C[164]), .CO(C[165]) );
  FA_3446 \FAINST[165].FA_  ( .A(A[165]), .B(n93), .CI(C[165]), .CO(C[166]) );
  FA_3445 \FAINST[166].FA_  ( .A(A[166]), .B(n92), .CI(C[166]), .CO(C[167]) );
  FA_3444 \FAINST[167].FA_  ( .A(A[167]), .B(n91), .CI(C[167]), .CO(C[168]) );
  FA_3443 \FAINST[168].FA_  ( .A(A[168]), .B(n90), .CI(C[168]), .CO(C[169]) );
  FA_3442 \FAINST[169].FA_  ( .A(A[169]), .B(n89), .CI(C[169]), .CO(C[170]) );
  FA_3441 \FAINST[170].FA_  ( .A(A[170]), .B(n88), .CI(C[170]), .CO(C[171]) );
  FA_3440 \FAINST[171].FA_  ( .A(A[171]), .B(n87), .CI(C[171]), .CO(C[172]) );
  FA_3439 \FAINST[172].FA_  ( .A(A[172]), .B(n86), .CI(C[172]), .CO(C[173]) );
  FA_3438 \FAINST[173].FA_  ( .A(A[173]), .B(n85), .CI(C[173]), .CO(C[174]) );
  FA_3437 \FAINST[174].FA_  ( .A(A[174]), .B(n84), .CI(C[174]), .CO(C[175]) );
  FA_3436 \FAINST[175].FA_  ( .A(A[175]), .B(n83), .CI(C[175]), .CO(C[176]) );
  FA_3435 \FAINST[176].FA_  ( .A(A[176]), .B(n82), .CI(C[176]), .CO(C[177]) );
  FA_3434 \FAINST[177].FA_  ( .A(A[177]), .B(n81), .CI(C[177]), .CO(C[178]) );
  FA_3433 \FAINST[178].FA_  ( .A(A[178]), .B(n80), .CI(C[178]), .CO(C[179]) );
  FA_3432 \FAINST[179].FA_  ( .A(A[179]), .B(n79), .CI(C[179]), .CO(C[180]) );
  FA_3431 \FAINST[180].FA_  ( .A(A[180]), .B(n78), .CI(C[180]), .CO(C[181]) );
  FA_3430 \FAINST[181].FA_  ( .A(A[181]), .B(n77), .CI(C[181]), .CO(C[182]) );
  FA_3429 \FAINST[182].FA_  ( .A(A[182]), .B(n76), .CI(C[182]), .CO(C[183]) );
  FA_3428 \FAINST[183].FA_  ( .A(A[183]), .B(n75), .CI(C[183]), .CO(C[184]) );
  FA_3427 \FAINST[184].FA_  ( .A(A[184]), .B(n74), .CI(C[184]), .CO(C[185]) );
  FA_3426 \FAINST[185].FA_  ( .A(A[185]), .B(n73), .CI(C[185]), .CO(C[186]) );
  FA_3425 \FAINST[186].FA_  ( .A(A[186]), .B(n72), .CI(C[186]), .CO(C[187]) );
  FA_3424 \FAINST[187].FA_  ( .A(A[187]), .B(n71), .CI(C[187]), .CO(C[188]) );
  FA_3423 \FAINST[188].FA_  ( .A(A[188]), .B(n70), .CI(C[188]), .CO(C[189]) );
  FA_3422 \FAINST[189].FA_  ( .A(A[189]), .B(n69), .CI(C[189]), .CO(C[190]) );
  FA_3421 \FAINST[190].FA_  ( .A(A[190]), .B(n68), .CI(C[190]), .CO(C[191]) );
  FA_3420 \FAINST[191].FA_  ( .A(A[191]), .B(n67), .CI(C[191]), .CO(C[192]) );
  FA_3419 \FAINST[192].FA_  ( .A(A[192]), .B(n66), .CI(C[192]), .CO(C[193]) );
  FA_3418 \FAINST[193].FA_  ( .A(A[193]), .B(n65), .CI(C[193]), .CO(C[194]) );
  FA_3417 \FAINST[194].FA_  ( .A(A[194]), .B(n64), .CI(C[194]), .CO(C[195]) );
  FA_3416 \FAINST[195].FA_  ( .A(A[195]), .B(n63), .CI(C[195]), .CO(C[196]) );
  FA_3415 \FAINST[196].FA_  ( .A(A[196]), .B(n62), .CI(C[196]), .CO(C[197]) );
  FA_3414 \FAINST[197].FA_  ( .A(A[197]), .B(n61), .CI(C[197]), .CO(C[198]) );
  FA_3413 \FAINST[198].FA_  ( .A(A[198]), .B(n60), .CI(C[198]), .CO(C[199]) );
  FA_3412 \FAINST[199].FA_  ( .A(A[199]), .B(n59), .CI(C[199]), .CO(C[200]) );
  FA_3411 \FAINST[200].FA_  ( .A(A[200]), .B(n58), .CI(C[200]), .CO(C[201]) );
  FA_3410 \FAINST[201].FA_  ( .A(A[201]), .B(n57), .CI(C[201]), .CO(C[202]) );
  FA_3409 \FAINST[202].FA_  ( .A(A[202]), .B(n56), .CI(C[202]), .CO(C[203]) );
  FA_3408 \FAINST[203].FA_  ( .A(A[203]), .B(n55), .CI(C[203]), .CO(C[204]) );
  FA_3407 \FAINST[204].FA_  ( .A(A[204]), .B(n54), .CI(C[204]), .CO(C[205]) );
  FA_3406 \FAINST[205].FA_  ( .A(A[205]), .B(n53), .CI(C[205]), .CO(C[206]) );
  FA_3405 \FAINST[206].FA_  ( .A(A[206]), .B(n52), .CI(C[206]), .CO(C[207]) );
  FA_3404 \FAINST[207].FA_  ( .A(A[207]), .B(n51), .CI(C[207]), .CO(C[208]) );
  FA_3403 \FAINST[208].FA_  ( .A(A[208]), .B(n50), .CI(C[208]), .CO(C[209]) );
  FA_3402 \FAINST[209].FA_  ( .A(A[209]), .B(n49), .CI(C[209]), .CO(C[210]) );
  FA_3401 \FAINST[210].FA_  ( .A(A[210]), .B(n48), .CI(C[210]), .CO(C[211]) );
  FA_3400 \FAINST[211].FA_  ( .A(A[211]), .B(n47), .CI(C[211]), .CO(C[212]) );
  FA_3399 \FAINST[212].FA_  ( .A(A[212]), .B(n46), .CI(C[212]), .CO(C[213]) );
  FA_3398 \FAINST[213].FA_  ( .A(A[213]), .B(n45), .CI(C[213]), .CO(C[214]) );
  FA_3397 \FAINST[214].FA_  ( .A(A[214]), .B(n44), .CI(C[214]), .CO(C[215]) );
  FA_3396 \FAINST[215].FA_  ( .A(A[215]), .B(n43), .CI(C[215]), .CO(C[216]) );
  FA_3395 \FAINST[216].FA_  ( .A(A[216]), .B(n42), .CI(C[216]), .CO(C[217]) );
  FA_3394 \FAINST[217].FA_  ( .A(A[217]), .B(n41), .CI(C[217]), .CO(C[218]) );
  FA_3393 \FAINST[218].FA_  ( .A(A[218]), .B(n40), .CI(C[218]), .CO(C[219]) );
  FA_3392 \FAINST[219].FA_  ( .A(A[219]), .B(n39), .CI(C[219]), .CO(C[220]) );
  FA_3391 \FAINST[220].FA_  ( .A(A[220]), .B(n38), .CI(C[220]), .CO(C[221]) );
  FA_3390 \FAINST[221].FA_  ( .A(A[221]), .B(n37), .CI(C[221]), .CO(C[222]) );
  FA_3389 \FAINST[222].FA_  ( .A(A[222]), .B(n36), .CI(C[222]), .CO(C[223]) );
  FA_3388 \FAINST[223].FA_  ( .A(A[223]), .B(n35), .CI(C[223]), .CO(C[224]) );
  FA_3387 \FAINST[224].FA_  ( .A(A[224]), .B(n34), .CI(C[224]), .CO(C[225]) );
  FA_3386 \FAINST[225].FA_  ( .A(A[225]), .B(n33), .CI(C[225]), .CO(C[226]) );
  FA_3385 \FAINST[226].FA_  ( .A(A[226]), .B(n32), .CI(C[226]), .CO(C[227]) );
  FA_3384 \FAINST[227].FA_  ( .A(A[227]), .B(n31), .CI(C[227]), .CO(C[228]) );
  FA_3383 \FAINST[228].FA_  ( .A(A[228]), .B(n30), .CI(C[228]), .CO(C[229]) );
  FA_3382 \FAINST[229].FA_  ( .A(A[229]), .B(n29), .CI(C[229]), .CO(C[230]) );
  FA_3381 \FAINST[230].FA_  ( .A(A[230]), .B(n28), .CI(C[230]), .CO(C[231]) );
  FA_3380 \FAINST[231].FA_  ( .A(A[231]), .B(n27), .CI(C[231]), .CO(C[232]) );
  FA_3379 \FAINST[232].FA_  ( .A(A[232]), .B(n26), .CI(C[232]), .CO(C[233]) );
  FA_3378 \FAINST[233].FA_  ( .A(A[233]), .B(n25), .CI(C[233]), .CO(C[234]) );
  FA_3377 \FAINST[234].FA_  ( .A(A[234]), .B(n24), .CI(C[234]), .CO(C[235]) );
  FA_3376 \FAINST[235].FA_  ( .A(A[235]), .B(n23), .CI(C[235]), .CO(C[236]) );
  FA_3375 \FAINST[236].FA_  ( .A(A[236]), .B(n22), .CI(C[236]), .CO(C[237]) );
  FA_3374 \FAINST[237].FA_  ( .A(A[237]), .B(n21), .CI(C[237]), .CO(C[238]) );
  FA_3373 \FAINST[238].FA_  ( .A(A[238]), .B(n20), .CI(C[238]), .CO(C[239]) );
  FA_3372 \FAINST[239].FA_  ( .A(A[239]), .B(n19), .CI(C[239]), .CO(C[240]) );
  FA_3371 \FAINST[240].FA_  ( .A(A[240]), .B(n18), .CI(C[240]), .CO(C[241]) );
  FA_3370 \FAINST[241].FA_  ( .A(A[241]), .B(n17), .CI(C[241]), .CO(C[242]) );
  FA_3369 \FAINST[242].FA_  ( .A(A[242]), .B(n16), .CI(C[242]), .CO(C[243]) );
  FA_3368 \FAINST[243].FA_  ( .A(A[243]), .B(n15), .CI(C[243]), .CO(C[244]) );
  FA_3367 \FAINST[244].FA_  ( .A(A[244]), .B(n14), .CI(C[244]), .CO(C[245]) );
  FA_3366 \FAINST[245].FA_  ( .A(A[245]), .B(n13), .CI(C[245]), .CO(C[246]) );
  FA_3365 \FAINST[246].FA_  ( .A(A[246]), .B(n12), .CI(C[246]), .CO(C[247]) );
  FA_3364 \FAINST[247].FA_  ( .A(A[247]), .B(n11), .CI(C[247]), .CO(C[248]) );
  FA_3363 \FAINST[248].FA_  ( .A(A[248]), .B(n10), .CI(C[248]), .CO(C[249]) );
  FA_3362 \FAINST[249].FA_  ( .A(A[249]), .B(n9), .CI(C[249]), .CO(C[250]) );
  FA_3361 \FAINST[250].FA_  ( .A(A[250]), .B(n8), .CI(C[250]), .CO(C[251]) );
  FA_3360 \FAINST[251].FA_  ( .A(A[251]), .B(n7), .CI(C[251]), .CO(C[252]) );
  FA_3359 \FAINST[252].FA_  ( .A(A[252]), .B(n6), .CI(C[252]), .CO(C[253]) );
  FA_3358 \FAINST[253].FA_  ( .A(A[253]), .B(n5), .CI(C[253]), .CO(C[254]) );
  FA_3357 \FAINST[254].FA_  ( .A(A[254]), .B(n4), .CI(C[254]), .CO(C[255]) );
  FA_3356 \FAINST[255].FA_  ( .A(A[255]), .B(n3), .CI(C[255]), .CO(C[256]) );
  FA_3355 \FAINST[256].FA_  ( .A(A[256]), .B(1'b1), .CI(C[256]), .CO(C[257])
         );
  FA_3354 \FAINST[257].FA_  ( .A(A[257]), .B(1'b1), .CI(C[257]), .CO(O) );
  IV U2 ( .A(B[159]), .Z(n99) );
  IV U3 ( .A(B[160]), .Z(n98) );
  IV U4 ( .A(B[161]), .Z(n97) );
  IV U5 ( .A(B[162]), .Z(n96) );
  IV U6 ( .A(B[163]), .Z(n95) );
  IV U7 ( .A(B[164]), .Z(n94) );
  IV U8 ( .A(B[165]), .Z(n93) );
  IV U9 ( .A(B[166]), .Z(n92) );
  IV U10 ( .A(B[167]), .Z(n91) );
  IV U11 ( .A(B[168]), .Z(n90) );
  IV U12 ( .A(B[249]), .Z(n9) );
  IV U13 ( .A(B[169]), .Z(n89) );
  IV U14 ( .A(B[170]), .Z(n88) );
  IV U15 ( .A(B[171]), .Z(n87) );
  IV U16 ( .A(B[172]), .Z(n86) );
  IV U17 ( .A(B[173]), .Z(n85) );
  IV U18 ( .A(B[174]), .Z(n84) );
  IV U19 ( .A(B[175]), .Z(n83) );
  IV U20 ( .A(B[176]), .Z(n82) );
  IV U21 ( .A(B[177]), .Z(n81) );
  IV U22 ( .A(B[178]), .Z(n80) );
  IV U23 ( .A(B[250]), .Z(n8) );
  IV U24 ( .A(B[179]), .Z(n79) );
  IV U25 ( .A(B[180]), .Z(n78) );
  IV U26 ( .A(B[181]), .Z(n77) );
  IV U27 ( .A(B[182]), .Z(n76) );
  IV U28 ( .A(B[183]), .Z(n75) );
  IV U29 ( .A(B[184]), .Z(n74) );
  IV U30 ( .A(B[185]), .Z(n73) );
  IV U31 ( .A(B[186]), .Z(n72) );
  IV U32 ( .A(B[187]), .Z(n71) );
  IV U33 ( .A(B[188]), .Z(n70) );
  IV U34 ( .A(B[251]), .Z(n7) );
  IV U35 ( .A(B[189]), .Z(n69) );
  IV U36 ( .A(B[190]), .Z(n68) );
  IV U37 ( .A(B[191]), .Z(n67) );
  IV U38 ( .A(B[192]), .Z(n66) );
  IV U39 ( .A(B[193]), .Z(n65) );
  IV U40 ( .A(B[194]), .Z(n64) );
  IV U41 ( .A(B[195]), .Z(n63) );
  IV U42 ( .A(B[196]), .Z(n62) );
  IV U43 ( .A(B[197]), .Z(n61) );
  IV U44 ( .A(B[198]), .Z(n60) );
  IV U45 ( .A(B[252]), .Z(n6) );
  IV U46 ( .A(B[199]), .Z(n59) );
  IV U47 ( .A(B[200]), .Z(n58) );
  IV U48 ( .A(B[201]), .Z(n57) );
  IV U49 ( .A(B[202]), .Z(n56) );
  IV U50 ( .A(B[203]), .Z(n55) );
  IV U51 ( .A(B[204]), .Z(n54) );
  IV U52 ( .A(B[205]), .Z(n53) );
  IV U53 ( .A(B[206]), .Z(n52) );
  IV U54 ( .A(B[207]), .Z(n51) );
  IV U55 ( .A(B[208]), .Z(n50) );
  IV U56 ( .A(B[253]), .Z(n5) );
  IV U57 ( .A(B[209]), .Z(n49) );
  IV U58 ( .A(B[210]), .Z(n48) );
  IV U59 ( .A(B[211]), .Z(n47) );
  IV U60 ( .A(B[212]), .Z(n46) );
  IV U61 ( .A(B[213]), .Z(n45) );
  IV U62 ( .A(B[214]), .Z(n44) );
  IV U63 ( .A(B[215]), .Z(n43) );
  IV U64 ( .A(B[216]), .Z(n42) );
  IV U65 ( .A(B[217]), .Z(n41) );
  IV U66 ( .A(B[218]), .Z(n40) );
  IV U67 ( .A(B[254]), .Z(n4) );
  IV U68 ( .A(B[219]), .Z(n39) );
  IV U69 ( .A(B[220]), .Z(n38) );
  IV U70 ( .A(B[221]), .Z(n37) );
  IV U71 ( .A(B[222]), .Z(n36) );
  IV U72 ( .A(B[223]), .Z(n35) );
  IV U73 ( .A(B[224]), .Z(n34) );
  IV U74 ( .A(B[225]), .Z(n33) );
  IV U75 ( .A(B[226]), .Z(n32) );
  IV U76 ( .A(B[227]), .Z(n31) );
  IV U77 ( .A(B[228]), .Z(n30) );
  IV U78 ( .A(B[255]), .Z(n3) );
  IV U79 ( .A(B[229]), .Z(n29) );
  IV U80 ( .A(B[230]), .Z(n28) );
  IV U81 ( .A(B[231]), .Z(n27) );
  IV U82 ( .A(B[232]), .Z(n26) );
  IV U83 ( .A(B[0]), .Z(n258) );
  IV U84 ( .A(B[1]), .Z(n257) );
  IV U85 ( .A(B[2]), .Z(n256) );
  IV U86 ( .A(B[3]), .Z(n255) );
  IV U87 ( .A(B[4]), .Z(n254) );
  IV U88 ( .A(B[5]), .Z(n253) );
  IV U89 ( .A(B[6]), .Z(n252) );
  IV U90 ( .A(B[7]), .Z(n251) );
  IV U91 ( .A(B[8]), .Z(n250) );
  IV U92 ( .A(B[233]), .Z(n25) );
  IV U93 ( .A(B[9]), .Z(n249) );
  IV U94 ( .A(B[10]), .Z(n248) );
  IV U95 ( .A(B[11]), .Z(n247) );
  IV U96 ( .A(B[12]), .Z(n246) );
  IV U97 ( .A(B[13]), .Z(n245) );
  IV U98 ( .A(B[14]), .Z(n244) );
  IV U99 ( .A(B[15]), .Z(n243) );
  IV U100 ( .A(B[16]), .Z(n242) );
  IV U101 ( .A(B[17]), .Z(n241) );
  IV U102 ( .A(B[18]), .Z(n240) );
  IV U103 ( .A(B[234]), .Z(n24) );
  IV U104 ( .A(B[19]), .Z(n239) );
  IV U105 ( .A(B[20]), .Z(n238) );
  IV U106 ( .A(B[21]), .Z(n237) );
  IV U107 ( .A(B[22]), .Z(n236) );
  IV U108 ( .A(B[23]), .Z(n235) );
  IV U109 ( .A(B[24]), .Z(n234) );
  IV U110 ( .A(B[25]), .Z(n233) );
  IV U111 ( .A(B[26]), .Z(n232) );
  IV U112 ( .A(B[27]), .Z(n231) );
  IV U113 ( .A(B[28]), .Z(n230) );
  IV U114 ( .A(B[235]), .Z(n23) );
  IV U115 ( .A(B[29]), .Z(n229) );
  IV U116 ( .A(B[30]), .Z(n228) );
  IV U117 ( .A(B[31]), .Z(n227) );
  IV U118 ( .A(B[32]), .Z(n226) );
  IV U119 ( .A(B[33]), .Z(n225) );
  IV U120 ( .A(B[34]), .Z(n224) );
  IV U121 ( .A(B[35]), .Z(n223) );
  IV U122 ( .A(B[36]), .Z(n222) );
  IV U123 ( .A(B[37]), .Z(n221) );
  IV U124 ( .A(B[38]), .Z(n220) );
  IV U125 ( .A(B[236]), .Z(n22) );
  IV U126 ( .A(B[39]), .Z(n219) );
  IV U127 ( .A(B[40]), .Z(n218) );
  IV U128 ( .A(B[41]), .Z(n217) );
  IV U129 ( .A(B[42]), .Z(n216) );
  IV U130 ( .A(B[43]), .Z(n215) );
  IV U131 ( .A(B[44]), .Z(n214) );
  IV U132 ( .A(B[45]), .Z(n213) );
  IV U133 ( .A(B[46]), .Z(n212) );
  IV U134 ( .A(B[47]), .Z(n211) );
  IV U135 ( .A(B[48]), .Z(n210) );
  IV U136 ( .A(B[237]), .Z(n21) );
  IV U137 ( .A(B[49]), .Z(n209) );
  IV U138 ( .A(B[50]), .Z(n208) );
  IV U139 ( .A(B[51]), .Z(n207) );
  IV U140 ( .A(B[52]), .Z(n206) );
  IV U141 ( .A(B[53]), .Z(n205) );
  IV U142 ( .A(B[54]), .Z(n204) );
  IV U143 ( .A(B[55]), .Z(n203) );
  IV U144 ( .A(B[56]), .Z(n202) );
  IV U145 ( .A(B[57]), .Z(n201) );
  IV U146 ( .A(B[58]), .Z(n200) );
  IV U147 ( .A(B[238]), .Z(n20) );
  IV U148 ( .A(B[59]), .Z(n199) );
  IV U149 ( .A(B[60]), .Z(n198) );
  IV U150 ( .A(B[61]), .Z(n197) );
  IV U151 ( .A(B[62]), .Z(n196) );
  IV U152 ( .A(B[63]), .Z(n195) );
  IV U153 ( .A(B[64]), .Z(n194) );
  IV U154 ( .A(B[65]), .Z(n193) );
  IV U155 ( .A(B[66]), .Z(n192) );
  IV U156 ( .A(B[67]), .Z(n191) );
  IV U157 ( .A(B[68]), .Z(n190) );
  IV U158 ( .A(B[239]), .Z(n19) );
  IV U159 ( .A(B[69]), .Z(n189) );
  IV U160 ( .A(B[70]), .Z(n188) );
  IV U161 ( .A(B[71]), .Z(n187) );
  IV U162 ( .A(B[72]), .Z(n186) );
  IV U163 ( .A(B[73]), .Z(n185) );
  IV U164 ( .A(B[74]), .Z(n184) );
  IV U165 ( .A(B[75]), .Z(n183) );
  IV U166 ( .A(B[76]), .Z(n182) );
  IV U167 ( .A(B[77]), .Z(n181) );
  IV U168 ( .A(B[78]), .Z(n180) );
  IV U169 ( .A(B[240]), .Z(n18) );
  IV U170 ( .A(B[79]), .Z(n179) );
  IV U171 ( .A(B[80]), .Z(n178) );
  IV U172 ( .A(B[81]), .Z(n177) );
  IV U173 ( .A(B[82]), .Z(n176) );
  IV U174 ( .A(B[83]), .Z(n175) );
  IV U175 ( .A(B[84]), .Z(n174) );
  IV U176 ( .A(B[85]), .Z(n173) );
  IV U177 ( .A(B[86]), .Z(n172) );
  IV U178 ( .A(B[87]), .Z(n171) );
  IV U179 ( .A(B[88]), .Z(n170) );
  IV U180 ( .A(B[241]), .Z(n17) );
  IV U181 ( .A(B[89]), .Z(n169) );
  IV U182 ( .A(B[90]), .Z(n168) );
  IV U183 ( .A(B[91]), .Z(n167) );
  IV U184 ( .A(B[92]), .Z(n166) );
  IV U185 ( .A(B[93]), .Z(n165) );
  IV U186 ( .A(B[94]), .Z(n164) );
  IV U187 ( .A(B[95]), .Z(n163) );
  IV U188 ( .A(B[96]), .Z(n162) );
  IV U189 ( .A(B[97]), .Z(n161) );
  IV U190 ( .A(B[98]), .Z(n160) );
  IV U191 ( .A(B[242]), .Z(n16) );
  IV U192 ( .A(B[99]), .Z(n159) );
  IV U193 ( .A(B[100]), .Z(n158) );
  IV U194 ( .A(B[101]), .Z(n157) );
  IV U195 ( .A(B[102]), .Z(n156) );
  IV U196 ( .A(B[103]), .Z(n155) );
  IV U197 ( .A(B[104]), .Z(n154) );
  IV U198 ( .A(B[105]), .Z(n153) );
  IV U199 ( .A(B[106]), .Z(n152) );
  IV U200 ( .A(B[107]), .Z(n151) );
  IV U201 ( .A(B[108]), .Z(n150) );
  IV U202 ( .A(B[243]), .Z(n15) );
  IV U203 ( .A(B[109]), .Z(n149) );
  IV U204 ( .A(B[110]), .Z(n148) );
  IV U205 ( .A(B[111]), .Z(n147) );
  IV U206 ( .A(B[112]), .Z(n146) );
  IV U207 ( .A(B[113]), .Z(n145) );
  IV U208 ( .A(B[114]), .Z(n144) );
  IV U209 ( .A(B[115]), .Z(n143) );
  IV U210 ( .A(B[116]), .Z(n142) );
  IV U211 ( .A(B[117]), .Z(n141) );
  IV U212 ( .A(B[118]), .Z(n140) );
  IV U213 ( .A(B[244]), .Z(n14) );
  IV U214 ( .A(B[119]), .Z(n139) );
  IV U215 ( .A(B[120]), .Z(n138) );
  IV U216 ( .A(B[121]), .Z(n137) );
  IV U217 ( .A(B[122]), .Z(n136) );
  IV U218 ( .A(B[123]), .Z(n135) );
  IV U219 ( .A(B[124]), .Z(n134) );
  IV U220 ( .A(B[125]), .Z(n133) );
  IV U221 ( .A(B[126]), .Z(n132) );
  IV U222 ( .A(B[127]), .Z(n131) );
  IV U223 ( .A(B[128]), .Z(n130) );
  IV U224 ( .A(B[245]), .Z(n13) );
  IV U225 ( .A(B[129]), .Z(n129) );
  IV U226 ( .A(B[130]), .Z(n128) );
  IV U227 ( .A(B[131]), .Z(n127) );
  IV U228 ( .A(B[132]), .Z(n126) );
  IV U229 ( .A(B[133]), .Z(n125) );
  IV U230 ( .A(B[134]), .Z(n124) );
  IV U231 ( .A(B[135]), .Z(n123) );
  IV U232 ( .A(B[136]), .Z(n122) );
  IV U233 ( .A(B[137]), .Z(n121) );
  IV U234 ( .A(B[138]), .Z(n120) );
  IV U235 ( .A(B[246]), .Z(n12) );
  IV U236 ( .A(B[139]), .Z(n119) );
  IV U237 ( .A(B[140]), .Z(n118) );
  IV U238 ( .A(B[141]), .Z(n117) );
  IV U239 ( .A(B[142]), .Z(n116) );
  IV U240 ( .A(B[143]), .Z(n115) );
  IV U241 ( .A(B[144]), .Z(n114) );
  IV U242 ( .A(B[145]), .Z(n113) );
  IV U243 ( .A(B[146]), .Z(n112) );
  IV U244 ( .A(B[147]), .Z(n111) );
  IV U245 ( .A(B[148]), .Z(n110) );
  IV U246 ( .A(B[247]), .Z(n11) );
  IV U247 ( .A(B[149]), .Z(n109) );
  IV U248 ( .A(B[150]), .Z(n108) );
  IV U249 ( .A(B[151]), .Z(n107) );
  IV U250 ( .A(B[152]), .Z(n106) );
  IV U251 ( .A(B[153]), .Z(n105) );
  IV U252 ( .A(B[154]), .Z(n104) );
  IV U253 ( .A(B[155]), .Z(n103) );
  IV U254 ( .A(B[156]), .Z(n102) );
  IV U255 ( .A(B[157]), .Z(n101) );
  IV U256 ( .A(B[158]), .Z(n100) );
  IV U257 ( .A(B[248]), .Z(n10) );
endmodule


module FA_3096 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XNOR U1 ( .A(CI), .B(A), .Z(S) );
endmodule


module FA_3097 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  NANDN U1 ( .A(CI), .B(S), .Z(CO) );
  XNOR U2 ( .A(A), .B(CI), .Z(S) );
endmodule


module FA_3098 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3099 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3100 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3101 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3102 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3103 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3104 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3105 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3106 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3107 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3108 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3109 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3110 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3111 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3112 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3113 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3114 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3115 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3116 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3117 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3118 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3119 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3120 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3121 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3122 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3123 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3124 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3125 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3126 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3127 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3128 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3129 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3130 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3131 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3132 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3133 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3134 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3135 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3136 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3137 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3138 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3139 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3140 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3141 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3142 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3143 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3144 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3145 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3146 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3147 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3148 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3149 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3150 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3151 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3152 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3153 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3154 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3155 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3156 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3157 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3158 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3159 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3160 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3161 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3162 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3163 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3164 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3165 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3166 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3167 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3168 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3169 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3170 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3171 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3172 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3173 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3174 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3175 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3176 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3177 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3178 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3179 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3180 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3181 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3182 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3183 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3184 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3185 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3186 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3187 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3188 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3189 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3190 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3191 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3192 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3193 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3194 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3195 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3196 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3197 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3198 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3199 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3200 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3201 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3202 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3203 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3204 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3205 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3206 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3207 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3208 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3209 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3210 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3211 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3212 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3213 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3214 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3215 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3216 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3217 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3218 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3219 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3220 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3221 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3222 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3223 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3224 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3225 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3226 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3227 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3228 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3229 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3230 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3231 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3232 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3233 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3234 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3235 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3236 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3237 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3238 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3239 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3240 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3241 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3242 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3243 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3244 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3245 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3246 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3247 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3248 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3249 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3250 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3251 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3252 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3253 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3254 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3255 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3256 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3257 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3258 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3259 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3260 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3261 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3262 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3263 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3264 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3265 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3266 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3267 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3268 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3269 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3270 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3271 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3272 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3273 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3274 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3275 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3276 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3277 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3278 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3279 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3280 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3281 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3282 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3283 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3284 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3285 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3286 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3287 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3288 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3289 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3290 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3291 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3292 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3293 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3294 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3295 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3296 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3297 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3298 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3299 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3300 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3301 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3302 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3303 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3304 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3305 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3306 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3307 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3308 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3309 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3310 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3311 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3312 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3313 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3314 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3315 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3316 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3317 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3318 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3319 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3320 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3321 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3322 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3323 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3324 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3325 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3326 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3327 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3328 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3329 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3330 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3331 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3332 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3333 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3334 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3335 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3336 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3337 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3338 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3339 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3340 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3341 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3342 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3343 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3344 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3345 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3346 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3347 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3348 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3349 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3350 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3351 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3352 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3353 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XNOR U1 ( .A(B), .B(A), .Z(S) );
  OR U2 ( .A(B), .B(A), .Z(CO) );
endmodule


module SUB_N258_2 ( A, B, S, CO );
  input [257:0] A;
  input [257:0] B;
  output [257:0] S;
  output CO;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258;
  wire   [257:1] C;

  FA_3353 \FAINST[0].FA_  ( .A(A[0]), .B(n258), .CI(1'b1), .S(S[0]), .CO(C[1])
         );
  FA_3352 \FAINST[1].FA_  ( .A(A[1]), .B(n257), .CI(C[1]), .S(S[1]), .CO(C[2])
         );
  FA_3351 \FAINST[2].FA_  ( .A(A[2]), .B(n256), .CI(C[2]), .S(S[2]), .CO(C[3])
         );
  FA_3350 \FAINST[3].FA_  ( .A(A[3]), .B(n255), .CI(C[3]), .S(S[3]), .CO(C[4])
         );
  FA_3349 \FAINST[4].FA_  ( .A(A[4]), .B(n254), .CI(C[4]), .S(S[4]), .CO(C[5])
         );
  FA_3348 \FAINST[5].FA_  ( .A(A[5]), .B(n253), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_3347 \FAINST[6].FA_  ( .A(A[6]), .B(n252), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_3346 \FAINST[7].FA_  ( .A(A[7]), .B(n251), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_3345 \FAINST[8].FA_  ( .A(A[8]), .B(n250), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_3344 \FAINST[9].FA_  ( .A(A[9]), .B(n249), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_3343 \FAINST[10].FA_  ( .A(A[10]), .B(n248), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_3342 \FAINST[11].FA_  ( .A(A[11]), .B(n247), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_3341 \FAINST[12].FA_  ( .A(A[12]), .B(n246), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_3340 \FAINST[13].FA_  ( .A(A[13]), .B(n245), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_3339 \FAINST[14].FA_  ( .A(A[14]), .B(n244), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_3338 \FAINST[15].FA_  ( .A(A[15]), .B(n243), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_3337 \FAINST[16].FA_  ( .A(A[16]), .B(n242), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_3336 \FAINST[17].FA_  ( .A(A[17]), .B(n241), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_3335 \FAINST[18].FA_  ( .A(A[18]), .B(n240), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_3334 \FAINST[19].FA_  ( .A(A[19]), .B(n239), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_3333 \FAINST[20].FA_  ( .A(A[20]), .B(n238), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_3332 \FAINST[21].FA_  ( .A(A[21]), .B(n237), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_3331 \FAINST[22].FA_  ( .A(A[22]), .B(n236), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3330 \FAINST[23].FA_  ( .A(A[23]), .B(n235), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3329 \FAINST[24].FA_  ( .A(A[24]), .B(n234), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3328 \FAINST[25].FA_  ( .A(A[25]), .B(n233), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3327 \FAINST[26].FA_  ( .A(A[26]), .B(n232), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3326 \FAINST[27].FA_  ( .A(A[27]), .B(n231), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3325 \FAINST[28].FA_  ( .A(A[28]), .B(n230), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3324 \FAINST[29].FA_  ( .A(A[29]), .B(n229), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3323 \FAINST[30].FA_  ( .A(A[30]), .B(n228), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3322 \FAINST[31].FA_  ( .A(A[31]), .B(n227), .CI(C[31]), .S(S[31]), .CO(
        C[32]) );
  FA_3321 \FAINST[32].FA_  ( .A(A[32]), .B(n226), .CI(C[32]), .S(S[32]), .CO(
        C[33]) );
  FA_3320 \FAINST[33].FA_  ( .A(A[33]), .B(n225), .CI(C[33]), .S(S[33]), .CO(
        C[34]) );
  FA_3319 \FAINST[34].FA_  ( .A(A[34]), .B(n224), .CI(C[34]), .S(S[34]), .CO(
        C[35]) );
  FA_3318 \FAINST[35].FA_  ( .A(A[35]), .B(n223), .CI(C[35]), .S(S[35]), .CO(
        C[36]) );
  FA_3317 \FAINST[36].FA_  ( .A(A[36]), .B(n222), .CI(C[36]), .S(S[36]), .CO(
        C[37]) );
  FA_3316 \FAINST[37].FA_  ( .A(A[37]), .B(n221), .CI(C[37]), .S(S[37]), .CO(
        C[38]) );
  FA_3315 \FAINST[38].FA_  ( .A(A[38]), .B(n220), .CI(C[38]), .S(S[38]), .CO(
        C[39]) );
  FA_3314 \FAINST[39].FA_  ( .A(A[39]), .B(n219), .CI(C[39]), .S(S[39]), .CO(
        C[40]) );
  FA_3313 \FAINST[40].FA_  ( .A(A[40]), .B(n218), .CI(C[40]), .S(S[40]), .CO(
        C[41]) );
  FA_3312 \FAINST[41].FA_  ( .A(A[41]), .B(n217), .CI(C[41]), .S(S[41]), .CO(
        C[42]) );
  FA_3311 \FAINST[42].FA_  ( .A(A[42]), .B(n216), .CI(C[42]), .S(S[42]), .CO(
        C[43]) );
  FA_3310 \FAINST[43].FA_  ( .A(A[43]), .B(n215), .CI(C[43]), .S(S[43]), .CO(
        C[44]) );
  FA_3309 \FAINST[44].FA_  ( .A(A[44]), .B(n214), .CI(C[44]), .S(S[44]), .CO(
        C[45]) );
  FA_3308 \FAINST[45].FA_  ( .A(A[45]), .B(n213), .CI(C[45]), .S(S[45]), .CO(
        C[46]) );
  FA_3307 \FAINST[46].FA_  ( .A(A[46]), .B(n212), .CI(C[46]), .S(S[46]), .CO(
        C[47]) );
  FA_3306 \FAINST[47].FA_  ( .A(A[47]), .B(n211), .CI(C[47]), .S(S[47]), .CO(
        C[48]) );
  FA_3305 \FAINST[48].FA_  ( .A(A[48]), .B(n210), .CI(C[48]), .S(S[48]), .CO(
        C[49]) );
  FA_3304 \FAINST[49].FA_  ( .A(A[49]), .B(n209), .CI(C[49]), .S(S[49]), .CO(
        C[50]) );
  FA_3303 \FAINST[50].FA_  ( .A(A[50]), .B(n208), .CI(C[50]), .S(S[50]), .CO(
        C[51]) );
  FA_3302 \FAINST[51].FA_  ( .A(A[51]), .B(n207), .CI(C[51]), .S(S[51]), .CO(
        C[52]) );
  FA_3301 \FAINST[52].FA_  ( .A(A[52]), .B(n206), .CI(C[52]), .S(S[52]), .CO(
        C[53]) );
  FA_3300 \FAINST[53].FA_  ( .A(A[53]), .B(n205), .CI(C[53]), .S(S[53]), .CO(
        C[54]) );
  FA_3299 \FAINST[54].FA_  ( .A(A[54]), .B(n204), .CI(C[54]), .S(S[54]), .CO(
        C[55]) );
  FA_3298 \FAINST[55].FA_  ( .A(A[55]), .B(n203), .CI(C[55]), .S(S[55]), .CO(
        C[56]) );
  FA_3297 \FAINST[56].FA_  ( .A(A[56]), .B(n202), .CI(C[56]), .S(S[56]), .CO(
        C[57]) );
  FA_3296 \FAINST[57].FA_  ( .A(A[57]), .B(n201), .CI(C[57]), .S(S[57]), .CO(
        C[58]) );
  FA_3295 \FAINST[58].FA_  ( .A(A[58]), .B(n200), .CI(C[58]), .S(S[58]), .CO(
        C[59]) );
  FA_3294 \FAINST[59].FA_  ( .A(A[59]), .B(n199), .CI(C[59]), .S(S[59]), .CO(
        C[60]) );
  FA_3293 \FAINST[60].FA_  ( .A(A[60]), .B(n198), .CI(C[60]), .S(S[60]), .CO(
        C[61]) );
  FA_3292 \FAINST[61].FA_  ( .A(A[61]), .B(n197), .CI(C[61]), .S(S[61]), .CO(
        C[62]) );
  FA_3291 \FAINST[62].FA_  ( .A(A[62]), .B(n196), .CI(C[62]), .S(S[62]), .CO(
        C[63]) );
  FA_3290 \FAINST[63].FA_  ( .A(A[63]), .B(n195), .CI(C[63]), .S(S[63]), .CO(
        C[64]) );
  FA_3289 \FAINST[64].FA_  ( .A(A[64]), .B(n194), .CI(C[64]), .S(S[64]), .CO(
        C[65]) );
  FA_3288 \FAINST[65].FA_  ( .A(A[65]), .B(n193), .CI(C[65]), .S(S[65]), .CO(
        C[66]) );
  FA_3287 \FAINST[66].FA_  ( .A(A[66]), .B(n192), .CI(C[66]), .S(S[66]), .CO(
        C[67]) );
  FA_3286 \FAINST[67].FA_  ( .A(A[67]), .B(n191), .CI(C[67]), .S(S[67]), .CO(
        C[68]) );
  FA_3285 \FAINST[68].FA_  ( .A(A[68]), .B(n190), .CI(C[68]), .S(S[68]), .CO(
        C[69]) );
  FA_3284 \FAINST[69].FA_  ( .A(A[69]), .B(n189), .CI(C[69]), .S(S[69]), .CO(
        C[70]) );
  FA_3283 \FAINST[70].FA_  ( .A(A[70]), .B(n188), .CI(C[70]), .S(S[70]), .CO(
        C[71]) );
  FA_3282 \FAINST[71].FA_  ( .A(A[71]), .B(n187), .CI(C[71]), .S(S[71]), .CO(
        C[72]) );
  FA_3281 \FAINST[72].FA_  ( .A(A[72]), .B(n186), .CI(C[72]), .S(S[72]), .CO(
        C[73]) );
  FA_3280 \FAINST[73].FA_  ( .A(A[73]), .B(n185), .CI(C[73]), .S(S[73]), .CO(
        C[74]) );
  FA_3279 \FAINST[74].FA_  ( .A(A[74]), .B(n184), .CI(C[74]), .S(S[74]), .CO(
        C[75]) );
  FA_3278 \FAINST[75].FA_  ( .A(A[75]), .B(n183), .CI(C[75]), .S(S[75]), .CO(
        C[76]) );
  FA_3277 \FAINST[76].FA_  ( .A(A[76]), .B(n182), .CI(C[76]), .S(S[76]), .CO(
        C[77]) );
  FA_3276 \FAINST[77].FA_  ( .A(A[77]), .B(n181), .CI(C[77]), .S(S[77]), .CO(
        C[78]) );
  FA_3275 \FAINST[78].FA_  ( .A(A[78]), .B(n180), .CI(C[78]), .S(S[78]), .CO(
        C[79]) );
  FA_3274 \FAINST[79].FA_  ( .A(A[79]), .B(n179), .CI(C[79]), .S(S[79]), .CO(
        C[80]) );
  FA_3273 \FAINST[80].FA_  ( .A(A[80]), .B(n178), .CI(C[80]), .S(S[80]), .CO(
        C[81]) );
  FA_3272 \FAINST[81].FA_  ( .A(A[81]), .B(n177), .CI(C[81]), .S(S[81]), .CO(
        C[82]) );
  FA_3271 \FAINST[82].FA_  ( .A(A[82]), .B(n176), .CI(C[82]), .S(S[82]), .CO(
        C[83]) );
  FA_3270 \FAINST[83].FA_  ( .A(A[83]), .B(n175), .CI(C[83]), .S(S[83]), .CO(
        C[84]) );
  FA_3269 \FAINST[84].FA_  ( .A(A[84]), .B(n174), .CI(C[84]), .S(S[84]), .CO(
        C[85]) );
  FA_3268 \FAINST[85].FA_  ( .A(A[85]), .B(n173), .CI(C[85]), .S(S[85]), .CO(
        C[86]) );
  FA_3267 \FAINST[86].FA_  ( .A(A[86]), .B(n172), .CI(C[86]), .S(S[86]), .CO(
        C[87]) );
  FA_3266 \FAINST[87].FA_  ( .A(A[87]), .B(n171), .CI(C[87]), .S(S[87]), .CO(
        C[88]) );
  FA_3265 \FAINST[88].FA_  ( .A(A[88]), .B(n170), .CI(C[88]), .S(S[88]), .CO(
        C[89]) );
  FA_3264 \FAINST[89].FA_  ( .A(A[89]), .B(n169), .CI(C[89]), .S(S[89]), .CO(
        C[90]) );
  FA_3263 \FAINST[90].FA_  ( .A(A[90]), .B(n168), .CI(C[90]), .S(S[90]), .CO(
        C[91]) );
  FA_3262 \FAINST[91].FA_  ( .A(A[91]), .B(n167), .CI(C[91]), .S(S[91]), .CO(
        C[92]) );
  FA_3261 \FAINST[92].FA_  ( .A(A[92]), .B(n166), .CI(C[92]), .S(S[92]), .CO(
        C[93]) );
  FA_3260 \FAINST[93].FA_  ( .A(A[93]), .B(n165), .CI(C[93]), .S(S[93]), .CO(
        C[94]) );
  FA_3259 \FAINST[94].FA_  ( .A(A[94]), .B(n164), .CI(C[94]), .S(S[94]), .CO(
        C[95]) );
  FA_3258 \FAINST[95].FA_  ( .A(A[95]), .B(n163), .CI(C[95]), .S(S[95]), .CO(
        C[96]) );
  FA_3257 \FAINST[96].FA_  ( .A(A[96]), .B(n162), .CI(C[96]), .S(S[96]), .CO(
        C[97]) );
  FA_3256 \FAINST[97].FA_  ( .A(A[97]), .B(n161), .CI(C[97]), .S(S[97]), .CO(
        C[98]) );
  FA_3255 \FAINST[98].FA_  ( .A(A[98]), .B(n160), .CI(C[98]), .S(S[98]), .CO(
        C[99]) );
  FA_3254 \FAINST[99].FA_  ( .A(A[99]), .B(n159), .CI(C[99]), .S(S[99]), .CO(
        C[100]) );
  FA_3253 \FAINST[100].FA_  ( .A(A[100]), .B(n158), .CI(C[100]), .S(S[100]), 
        .CO(C[101]) );
  FA_3252 \FAINST[101].FA_  ( .A(A[101]), .B(n157), .CI(C[101]), .S(S[101]), 
        .CO(C[102]) );
  FA_3251 \FAINST[102].FA_  ( .A(A[102]), .B(n156), .CI(C[102]), .S(S[102]), 
        .CO(C[103]) );
  FA_3250 \FAINST[103].FA_  ( .A(A[103]), .B(n155), .CI(C[103]), .S(S[103]), 
        .CO(C[104]) );
  FA_3249 \FAINST[104].FA_  ( .A(A[104]), .B(n154), .CI(C[104]), .S(S[104]), 
        .CO(C[105]) );
  FA_3248 \FAINST[105].FA_  ( .A(A[105]), .B(n153), .CI(C[105]), .S(S[105]), 
        .CO(C[106]) );
  FA_3247 \FAINST[106].FA_  ( .A(A[106]), .B(n152), .CI(C[106]), .S(S[106]), 
        .CO(C[107]) );
  FA_3246 \FAINST[107].FA_  ( .A(A[107]), .B(n151), .CI(C[107]), .S(S[107]), 
        .CO(C[108]) );
  FA_3245 \FAINST[108].FA_  ( .A(A[108]), .B(n150), .CI(C[108]), .S(S[108]), 
        .CO(C[109]) );
  FA_3244 \FAINST[109].FA_  ( .A(A[109]), .B(n149), .CI(C[109]), .S(S[109]), 
        .CO(C[110]) );
  FA_3243 \FAINST[110].FA_  ( .A(A[110]), .B(n148), .CI(C[110]), .S(S[110]), 
        .CO(C[111]) );
  FA_3242 \FAINST[111].FA_  ( .A(A[111]), .B(n147), .CI(C[111]), .S(S[111]), 
        .CO(C[112]) );
  FA_3241 \FAINST[112].FA_  ( .A(A[112]), .B(n146), .CI(C[112]), .S(S[112]), 
        .CO(C[113]) );
  FA_3240 \FAINST[113].FA_  ( .A(A[113]), .B(n145), .CI(C[113]), .S(S[113]), 
        .CO(C[114]) );
  FA_3239 \FAINST[114].FA_  ( .A(A[114]), .B(n144), .CI(C[114]), .S(S[114]), 
        .CO(C[115]) );
  FA_3238 \FAINST[115].FA_  ( .A(A[115]), .B(n143), .CI(C[115]), .S(S[115]), 
        .CO(C[116]) );
  FA_3237 \FAINST[116].FA_  ( .A(A[116]), .B(n142), .CI(C[116]), .S(S[116]), 
        .CO(C[117]) );
  FA_3236 \FAINST[117].FA_  ( .A(A[117]), .B(n141), .CI(C[117]), .S(S[117]), 
        .CO(C[118]) );
  FA_3235 \FAINST[118].FA_  ( .A(A[118]), .B(n140), .CI(C[118]), .S(S[118]), 
        .CO(C[119]) );
  FA_3234 \FAINST[119].FA_  ( .A(A[119]), .B(n139), .CI(C[119]), .S(S[119]), 
        .CO(C[120]) );
  FA_3233 \FAINST[120].FA_  ( .A(A[120]), .B(n138), .CI(C[120]), .S(S[120]), 
        .CO(C[121]) );
  FA_3232 \FAINST[121].FA_  ( .A(A[121]), .B(n137), .CI(C[121]), .S(S[121]), 
        .CO(C[122]) );
  FA_3231 \FAINST[122].FA_  ( .A(A[122]), .B(n136), .CI(C[122]), .S(S[122]), 
        .CO(C[123]) );
  FA_3230 \FAINST[123].FA_  ( .A(A[123]), .B(n135), .CI(C[123]), .S(S[123]), 
        .CO(C[124]) );
  FA_3229 \FAINST[124].FA_  ( .A(A[124]), .B(n134), .CI(C[124]), .S(S[124]), 
        .CO(C[125]) );
  FA_3228 \FAINST[125].FA_  ( .A(A[125]), .B(n133), .CI(C[125]), .S(S[125]), 
        .CO(C[126]) );
  FA_3227 \FAINST[126].FA_  ( .A(A[126]), .B(n132), .CI(C[126]), .S(S[126]), 
        .CO(C[127]) );
  FA_3226 \FAINST[127].FA_  ( .A(A[127]), .B(n131), .CI(C[127]), .S(S[127]), 
        .CO(C[128]) );
  FA_3225 \FAINST[128].FA_  ( .A(A[128]), .B(n130), .CI(C[128]), .S(S[128]), 
        .CO(C[129]) );
  FA_3224 \FAINST[129].FA_  ( .A(A[129]), .B(n129), .CI(C[129]), .S(S[129]), 
        .CO(C[130]) );
  FA_3223 \FAINST[130].FA_  ( .A(A[130]), .B(n128), .CI(C[130]), .S(S[130]), 
        .CO(C[131]) );
  FA_3222 \FAINST[131].FA_  ( .A(A[131]), .B(n127), .CI(C[131]), .S(S[131]), 
        .CO(C[132]) );
  FA_3221 \FAINST[132].FA_  ( .A(A[132]), .B(n126), .CI(C[132]), .S(S[132]), 
        .CO(C[133]) );
  FA_3220 \FAINST[133].FA_  ( .A(A[133]), .B(n125), .CI(C[133]), .S(S[133]), 
        .CO(C[134]) );
  FA_3219 \FAINST[134].FA_  ( .A(A[134]), .B(n124), .CI(C[134]), .S(S[134]), 
        .CO(C[135]) );
  FA_3218 \FAINST[135].FA_  ( .A(A[135]), .B(n123), .CI(C[135]), .S(S[135]), 
        .CO(C[136]) );
  FA_3217 \FAINST[136].FA_  ( .A(A[136]), .B(n122), .CI(C[136]), .S(S[136]), 
        .CO(C[137]) );
  FA_3216 \FAINST[137].FA_  ( .A(A[137]), .B(n121), .CI(C[137]), .S(S[137]), 
        .CO(C[138]) );
  FA_3215 \FAINST[138].FA_  ( .A(A[138]), .B(n120), .CI(C[138]), .S(S[138]), 
        .CO(C[139]) );
  FA_3214 \FAINST[139].FA_  ( .A(A[139]), .B(n119), .CI(C[139]), .S(S[139]), 
        .CO(C[140]) );
  FA_3213 \FAINST[140].FA_  ( .A(A[140]), .B(n118), .CI(C[140]), .S(S[140]), 
        .CO(C[141]) );
  FA_3212 \FAINST[141].FA_  ( .A(A[141]), .B(n117), .CI(C[141]), .S(S[141]), 
        .CO(C[142]) );
  FA_3211 \FAINST[142].FA_  ( .A(A[142]), .B(n116), .CI(C[142]), .S(S[142]), 
        .CO(C[143]) );
  FA_3210 \FAINST[143].FA_  ( .A(A[143]), .B(n115), .CI(C[143]), .S(S[143]), 
        .CO(C[144]) );
  FA_3209 \FAINST[144].FA_  ( .A(A[144]), .B(n114), .CI(C[144]), .S(S[144]), 
        .CO(C[145]) );
  FA_3208 \FAINST[145].FA_  ( .A(A[145]), .B(n113), .CI(C[145]), .S(S[145]), 
        .CO(C[146]) );
  FA_3207 \FAINST[146].FA_  ( .A(A[146]), .B(n112), .CI(C[146]), .S(S[146]), 
        .CO(C[147]) );
  FA_3206 \FAINST[147].FA_  ( .A(A[147]), .B(n111), .CI(C[147]), .S(S[147]), 
        .CO(C[148]) );
  FA_3205 \FAINST[148].FA_  ( .A(A[148]), .B(n110), .CI(C[148]), .S(S[148]), 
        .CO(C[149]) );
  FA_3204 \FAINST[149].FA_  ( .A(A[149]), .B(n109), .CI(C[149]), .S(S[149]), 
        .CO(C[150]) );
  FA_3203 \FAINST[150].FA_  ( .A(A[150]), .B(n108), .CI(C[150]), .S(S[150]), 
        .CO(C[151]) );
  FA_3202 \FAINST[151].FA_  ( .A(A[151]), .B(n107), .CI(C[151]), .S(S[151]), 
        .CO(C[152]) );
  FA_3201 \FAINST[152].FA_  ( .A(A[152]), .B(n106), .CI(C[152]), .S(S[152]), 
        .CO(C[153]) );
  FA_3200 \FAINST[153].FA_  ( .A(A[153]), .B(n105), .CI(C[153]), .S(S[153]), 
        .CO(C[154]) );
  FA_3199 \FAINST[154].FA_  ( .A(A[154]), .B(n104), .CI(C[154]), .S(S[154]), 
        .CO(C[155]) );
  FA_3198 \FAINST[155].FA_  ( .A(A[155]), .B(n103), .CI(C[155]), .S(S[155]), 
        .CO(C[156]) );
  FA_3197 \FAINST[156].FA_  ( .A(A[156]), .B(n102), .CI(C[156]), .S(S[156]), 
        .CO(C[157]) );
  FA_3196 \FAINST[157].FA_  ( .A(A[157]), .B(n101), .CI(C[157]), .S(S[157]), 
        .CO(C[158]) );
  FA_3195 \FAINST[158].FA_  ( .A(A[158]), .B(n100), .CI(C[158]), .S(S[158]), 
        .CO(C[159]) );
  FA_3194 \FAINST[159].FA_  ( .A(A[159]), .B(n99), .CI(C[159]), .S(S[159]), 
        .CO(C[160]) );
  FA_3193 \FAINST[160].FA_  ( .A(A[160]), .B(n98), .CI(C[160]), .S(S[160]), 
        .CO(C[161]) );
  FA_3192 \FAINST[161].FA_  ( .A(A[161]), .B(n97), .CI(C[161]), .S(S[161]), 
        .CO(C[162]) );
  FA_3191 \FAINST[162].FA_  ( .A(A[162]), .B(n96), .CI(C[162]), .S(S[162]), 
        .CO(C[163]) );
  FA_3190 \FAINST[163].FA_  ( .A(A[163]), .B(n95), .CI(C[163]), .S(S[163]), 
        .CO(C[164]) );
  FA_3189 \FAINST[164].FA_  ( .A(A[164]), .B(n94), .CI(C[164]), .S(S[164]), 
        .CO(C[165]) );
  FA_3188 \FAINST[165].FA_  ( .A(A[165]), .B(n93), .CI(C[165]), .S(S[165]), 
        .CO(C[166]) );
  FA_3187 \FAINST[166].FA_  ( .A(A[166]), .B(n92), .CI(C[166]), .S(S[166]), 
        .CO(C[167]) );
  FA_3186 \FAINST[167].FA_  ( .A(A[167]), .B(n91), .CI(C[167]), .S(S[167]), 
        .CO(C[168]) );
  FA_3185 \FAINST[168].FA_  ( .A(A[168]), .B(n90), .CI(C[168]), .S(S[168]), 
        .CO(C[169]) );
  FA_3184 \FAINST[169].FA_  ( .A(A[169]), .B(n89), .CI(C[169]), .S(S[169]), 
        .CO(C[170]) );
  FA_3183 \FAINST[170].FA_  ( .A(A[170]), .B(n88), .CI(C[170]), .S(S[170]), 
        .CO(C[171]) );
  FA_3182 \FAINST[171].FA_  ( .A(A[171]), .B(n87), .CI(C[171]), .S(S[171]), 
        .CO(C[172]) );
  FA_3181 \FAINST[172].FA_  ( .A(A[172]), .B(n86), .CI(C[172]), .S(S[172]), 
        .CO(C[173]) );
  FA_3180 \FAINST[173].FA_  ( .A(A[173]), .B(n85), .CI(C[173]), .S(S[173]), 
        .CO(C[174]) );
  FA_3179 \FAINST[174].FA_  ( .A(A[174]), .B(n84), .CI(C[174]), .S(S[174]), 
        .CO(C[175]) );
  FA_3178 \FAINST[175].FA_  ( .A(A[175]), .B(n83), .CI(C[175]), .S(S[175]), 
        .CO(C[176]) );
  FA_3177 \FAINST[176].FA_  ( .A(A[176]), .B(n82), .CI(C[176]), .S(S[176]), 
        .CO(C[177]) );
  FA_3176 \FAINST[177].FA_  ( .A(A[177]), .B(n81), .CI(C[177]), .S(S[177]), 
        .CO(C[178]) );
  FA_3175 \FAINST[178].FA_  ( .A(A[178]), .B(n80), .CI(C[178]), .S(S[178]), 
        .CO(C[179]) );
  FA_3174 \FAINST[179].FA_  ( .A(A[179]), .B(n79), .CI(C[179]), .S(S[179]), 
        .CO(C[180]) );
  FA_3173 \FAINST[180].FA_  ( .A(A[180]), .B(n78), .CI(C[180]), .S(S[180]), 
        .CO(C[181]) );
  FA_3172 \FAINST[181].FA_  ( .A(A[181]), .B(n77), .CI(C[181]), .S(S[181]), 
        .CO(C[182]) );
  FA_3171 \FAINST[182].FA_  ( .A(A[182]), .B(n76), .CI(C[182]), .S(S[182]), 
        .CO(C[183]) );
  FA_3170 \FAINST[183].FA_  ( .A(A[183]), .B(n75), .CI(C[183]), .S(S[183]), 
        .CO(C[184]) );
  FA_3169 \FAINST[184].FA_  ( .A(A[184]), .B(n74), .CI(C[184]), .S(S[184]), 
        .CO(C[185]) );
  FA_3168 \FAINST[185].FA_  ( .A(A[185]), .B(n73), .CI(C[185]), .S(S[185]), 
        .CO(C[186]) );
  FA_3167 \FAINST[186].FA_  ( .A(A[186]), .B(n72), .CI(C[186]), .S(S[186]), 
        .CO(C[187]) );
  FA_3166 \FAINST[187].FA_  ( .A(A[187]), .B(n71), .CI(C[187]), .S(S[187]), 
        .CO(C[188]) );
  FA_3165 \FAINST[188].FA_  ( .A(A[188]), .B(n70), .CI(C[188]), .S(S[188]), 
        .CO(C[189]) );
  FA_3164 \FAINST[189].FA_  ( .A(A[189]), .B(n69), .CI(C[189]), .S(S[189]), 
        .CO(C[190]) );
  FA_3163 \FAINST[190].FA_  ( .A(A[190]), .B(n68), .CI(C[190]), .S(S[190]), 
        .CO(C[191]) );
  FA_3162 \FAINST[191].FA_  ( .A(A[191]), .B(n67), .CI(C[191]), .S(S[191]), 
        .CO(C[192]) );
  FA_3161 \FAINST[192].FA_  ( .A(A[192]), .B(n66), .CI(C[192]), .S(S[192]), 
        .CO(C[193]) );
  FA_3160 \FAINST[193].FA_  ( .A(A[193]), .B(n65), .CI(C[193]), .S(S[193]), 
        .CO(C[194]) );
  FA_3159 \FAINST[194].FA_  ( .A(A[194]), .B(n64), .CI(C[194]), .S(S[194]), 
        .CO(C[195]) );
  FA_3158 \FAINST[195].FA_  ( .A(A[195]), .B(n63), .CI(C[195]), .S(S[195]), 
        .CO(C[196]) );
  FA_3157 \FAINST[196].FA_  ( .A(A[196]), .B(n62), .CI(C[196]), .S(S[196]), 
        .CO(C[197]) );
  FA_3156 \FAINST[197].FA_  ( .A(A[197]), .B(n61), .CI(C[197]), .S(S[197]), 
        .CO(C[198]) );
  FA_3155 \FAINST[198].FA_  ( .A(A[198]), .B(n60), .CI(C[198]), .S(S[198]), 
        .CO(C[199]) );
  FA_3154 \FAINST[199].FA_  ( .A(A[199]), .B(n59), .CI(C[199]), .S(S[199]), 
        .CO(C[200]) );
  FA_3153 \FAINST[200].FA_  ( .A(A[200]), .B(n58), .CI(C[200]), .S(S[200]), 
        .CO(C[201]) );
  FA_3152 \FAINST[201].FA_  ( .A(A[201]), .B(n57), .CI(C[201]), .S(S[201]), 
        .CO(C[202]) );
  FA_3151 \FAINST[202].FA_  ( .A(A[202]), .B(n56), .CI(C[202]), .S(S[202]), 
        .CO(C[203]) );
  FA_3150 \FAINST[203].FA_  ( .A(A[203]), .B(n55), .CI(C[203]), .S(S[203]), 
        .CO(C[204]) );
  FA_3149 \FAINST[204].FA_  ( .A(A[204]), .B(n54), .CI(C[204]), .S(S[204]), 
        .CO(C[205]) );
  FA_3148 \FAINST[205].FA_  ( .A(A[205]), .B(n53), .CI(C[205]), .S(S[205]), 
        .CO(C[206]) );
  FA_3147 \FAINST[206].FA_  ( .A(A[206]), .B(n52), .CI(C[206]), .S(S[206]), 
        .CO(C[207]) );
  FA_3146 \FAINST[207].FA_  ( .A(A[207]), .B(n51), .CI(C[207]), .S(S[207]), 
        .CO(C[208]) );
  FA_3145 \FAINST[208].FA_  ( .A(A[208]), .B(n50), .CI(C[208]), .S(S[208]), 
        .CO(C[209]) );
  FA_3144 \FAINST[209].FA_  ( .A(A[209]), .B(n49), .CI(C[209]), .S(S[209]), 
        .CO(C[210]) );
  FA_3143 \FAINST[210].FA_  ( .A(A[210]), .B(n48), .CI(C[210]), .S(S[210]), 
        .CO(C[211]) );
  FA_3142 \FAINST[211].FA_  ( .A(A[211]), .B(n47), .CI(C[211]), .S(S[211]), 
        .CO(C[212]) );
  FA_3141 \FAINST[212].FA_  ( .A(A[212]), .B(n46), .CI(C[212]), .S(S[212]), 
        .CO(C[213]) );
  FA_3140 \FAINST[213].FA_  ( .A(A[213]), .B(n45), .CI(C[213]), .S(S[213]), 
        .CO(C[214]) );
  FA_3139 \FAINST[214].FA_  ( .A(A[214]), .B(n44), .CI(C[214]), .S(S[214]), 
        .CO(C[215]) );
  FA_3138 \FAINST[215].FA_  ( .A(A[215]), .B(n43), .CI(C[215]), .S(S[215]), 
        .CO(C[216]) );
  FA_3137 \FAINST[216].FA_  ( .A(A[216]), .B(n42), .CI(C[216]), .S(S[216]), 
        .CO(C[217]) );
  FA_3136 \FAINST[217].FA_  ( .A(A[217]), .B(n41), .CI(C[217]), .S(S[217]), 
        .CO(C[218]) );
  FA_3135 \FAINST[218].FA_  ( .A(A[218]), .B(n40), .CI(C[218]), .S(S[218]), 
        .CO(C[219]) );
  FA_3134 \FAINST[219].FA_  ( .A(A[219]), .B(n39), .CI(C[219]), .S(S[219]), 
        .CO(C[220]) );
  FA_3133 \FAINST[220].FA_  ( .A(A[220]), .B(n38), .CI(C[220]), .S(S[220]), 
        .CO(C[221]) );
  FA_3132 \FAINST[221].FA_  ( .A(A[221]), .B(n37), .CI(C[221]), .S(S[221]), 
        .CO(C[222]) );
  FA_3131 \FAINST[222].FA_  ( .A(A[222]), .B(n36), .CI(C[222]), .S(S[222]), 
        .CO(C[223]) );
  FA_3130 \FAINST[223].FA_  ( .A(A[223]), .B(n35), .CI(C[223]), .S(S[223]), 
        .CO(C[224]) );
  FA_3129 \FAINST[224].FA_  ( .A(A[224]), .B(n34), .CI(C[224]), .S(S[224]), 
        .CO(C[225]) );
  FA_3128 \FAINST[225].FA_  ( .A(A[225]), .B(n33), .CI(C[225]), .S(S[225]), 
        .CO(C[226]) );
  FA_3127 \FAINST[226].FA_  ( .A(A[226]), .B(n32), .CI(C[226]), .S(S[226]), 
        .CO(C[227]) );
  FA_3126 \FAINST[227].FA_  ( .A(A[227]), .B(n31), .CI(C[227]), .S(S[227]), 
        .CO(C[228]) );
  FA_3125 \FAINST[228].FA_  ( .A(A[228]), .B(n30), .CI(C[228]), .S(S[228]), 
        .CO(C[229]) );
  FA_3124 \FAINST[229].FA_  ( .A(A[229]), .B(n29), .CI(C[229]), .S(S[229]), 
        .CO(C[230]) );
  FA_3123 \FAINST[230].FA_  ( .A(A[230]), .B(n28), .CI(C[230]), .S(S[230]), 
        .CO(C[231]) );
  FA_3122 \FAINST[231].FA_  ( .A(A[231]), .B(n27), .CI(C[231]), .S(S[231]), 
        .CO(C[232]) );
  FA_3121 \FAINST[232].FA_  ( .A(A[232]), .B(n26), .CI(C[232]), .S(S[232]), 
        .CO(C[233]) );
  FA_3120 \FAINST[233].FA_  ( .A(A[233]), .B(n25), .CI(C[233]), .S(S[233]), 
        .CO(C[234]) );
  FA_3119 \FAINST[234].FA_  ( .A(A[234]), .B(n24), .CI(C[234]), .S(S[234]), 
        .CO(C[235]) );
  FA_3118 \FAINST[235].FA_  ( .A(A[235]), .B(n23), .CI(C[235]), .S(S[235]), 
        .CO(C[236]) );
  FA_3117 \FAINST[236].FA_  ( .A(A[236]), .B(n22), .CI(C[236]), .S(S[236]), 
        .CO(C[237]) );
  FA_3116 \FAINST[237].FA_  ( .A(A[237]), .B(n21), .CI(C[237]), .S(S[237]), 
        .CO(C[238]) );
  FA_3115 \FAINST[238].FA_  ( .A(A[238]), .B(n20), .CI(C[238]), .S(S[238]), 
        .CO(C[239]) );
  FA_3114 \FAINST[239].FA_  ( .A(A[239]), .B(n19), .CI(C[239]), .S(S[239]), 
        .CO(C[240]) );
  FA_3113 \FAINST[240].FA_  ( .A(A[240]), .B(n18), .CI(C[240]), .S(S[240]), 
        .CO(C[241]) );
  FA_3112 \FAINST[241].FA_  ( .A(A[241]), .B(n17), .CI(C[241]), .S(S[241]), 
        .CO(C[242]) );
  FA_3111 \FAINST[242].FA_  ( .A(A[242]), .B(n16), .CI(C[242]), .S(S[242]), 
        .CO(C[243]) );
  FA_3110 \FAINST[243].FA_  ( .A(A[243]), .B(n15), .CI(C[243]), .S(S[243]), 
        .CO(C[244]) );
  FA_3109 \FAINST[244].FA_  ( .A(A[244]), .B(n14), .CI(C[244]), .S(S[244]), 
        .CO(C[245]) );
  FA_3108 \FAINST[245].FA_  ( .A(A[245]), .B(n13), .CI(C[245]), .S(S[245]), 
        .CO(C[246]) );
  FA_3107 \FAINST[246].FA_  ( .A(A[246]), .B(n12), .CI(C[246]), .S(S[246]), 
        .CO(C[247]) );
  FA_3106 \FAINST[247].FA_  ( .A(A[247]), .B(n11), .CI(C[247]), .S(S[247]), 
        .CO(C[248]) );
  FA_3105 \FAINST[248].FA_  ( .A(A[248]), .B(n10), .CI(C[248]), .S(S[248]), 
        .CO(C[249]) );
  FA_3104 \FAINST[249].FA_  ( .A(A[249]), .B(n9), .CI(C[249]), .S(S[249]), 
        .CO(C[250]) );
  FA_3103 \FAINST[250].FA_  ( .A(A[250]), .B(n8), .CI(C[250]), .S(S[250]), 
        .CO(C[251]) );
  FA_3102 \FAINST[251].FA_  ( .A(A[251]), .B(n7), .CI(C[251]), .S(S[251]), 
        .CO(C[252]) );
  FA_3101 \FAINST[252].FA_  ( .A(A[252]), .B(n6), .CI(C[252]), .S(S[252]), 
        .CO(C[253]) );
  FA_3100 \FAINST[253].FA_  ( .A(A[253]), .B(n5), .CI(C[253]), .S(S[253]), 
        .CO(C[254]) );
  FA_3099 \FAINST[254].FA_  ( .A(A[254]), .B(n4), .CI(C[254]), .S(S[254]), 
        .CO(C[255]) );
  FA_3098 \FAINST[255].FA_  ( .A(A[255]), .B(n3), .CI(C[255]), .S(S[255]), 
        .CO(C[256]) );
  FA_3097 \FAINST[256].FA_  ( .A(A[256]), .B(1'b1), .CI(C[256]), .S(S[256]), 
        .CO(C[257]) );
  FA_3096 \FAINST[257].FA_  ( .A(A[257]), .B(1'b1), .CI(C[257]), .S(S[257]) );
  IV U2 ( .A(B[159]), .Z(n99) );
  IV U3 ( .A(B[160]), .Z(n98) );
  IV U4 ( .A(B[161]), .Z(n97) );
  IV U5 ( .A(B[162]), .Z(n96) );
  IV U6 ( .A(B[163]), .Z(n95) );
  IV U7 ( .A(B[164]), .Z(n94) );
  IV U8 ( .A(B[165]), .Z(n93) );
  IV U9 ( .A(B[166]), .Z(n92) );
  IV U10 ( .A(B[167]), .Z(n91) );
  IV U11 ( .A(B[168]), .Z(n90) );
  IV U12 ( .A(B[249]), .Z(n9) );
  IV U13 ( .A(B[169]), .Z(n89) );
  IV U14 ( .A(B[170]), .Z(n88) );
  IV U15 ( .A(B[171]), .Z(n87) );
  IV U16 ( .A(B[172]), .Z(n86) );
  IV U17 ( .A(B[173]), .Z(n85) );
  IV U18 ( .A(B[174]), .Z(n84) );
  IV U19 ( .A(B[175]), .Z(n83) );
  IV U20 ( .A(B[176]), .Z(n82) );
  IV U21 ( .A(B[177]), .Z(n81) );
  IV U22 ( .A(B[178]), .Z(n80) );
  IV U23 ( .A(B[250]), .Z(n8) );
  IV U24 ( .A(B[179]), .Z(n79) );
  IV U25 ( .A(B[180]), .Z(n78) );
  IV U26 ( .A(B[181]), .Z(n77) );
  IV U27 ( .A(B[182]), .Z(n76) );
  IV U28 ( .A(B[183]), .Z(n75) );
  IV U29 ( .A(B[184]), .Z(n74) );
  IV U30 ( .A(B[185]), .Z(n73) );
  IV U31 ( .A(B[186]), .Z(n72) );
  IV U32 ( .A(B[187]), .Z(n71) );
  IV U33 ( .A(B[188]), .Z(n70) );
  IV U34 ( .A(B[251]), .Z(n7) );
  IV U35 ( .A(B[189]), .Z(n69) );
  IV U36 ( .A(B[190]), .Z(n68) );
  IV U37 ( .A(B[191]), .Z(n67) );
  IV U38 ( .A(B[192]), .Z(n66) );
  IV U39 ( .A(B[193]), .Z(n65) );
  IV U40 ( .A(B[194]), .Z(n64) );
  IV U41 ( .A(B[195]), .Z(n63) );
  IV U42 ( .A(B[196]), .Z(n62) );
  IV U43 ( .A(B[197]), .Z(n61) );
  IV U44 ( .A(B[198]), .Z(n60) );
  IV U45 ( .A(B[252]), .Z(n6) );
  IV U46 ( .A(B[199]), .Z(n59) );
  IV U47 ( .A(B[200]), .Z(n58) );
  IV U48 ( .A(B[201]), .Z(n57) );
  IV U49 ( .A(B[202]), .Z(n56) );
  IV U50 ( .A(B[203]), .Z(n55) );
  IV U51 ( .A(B[204]), .Z(n54) );
  IV U52 ( .A(B[205]), .Z(n53) );
  IV U53 ( .A(B[206]), .Z(n52) );
  IV U54 ( .A(B[207]), .Z(n51) );
  IV U55 ( .A(B[208]), .Z(n50) );
  IV U56 ( .A(B[253]), .Z(n5) );
  IV U57 ( .A(B[209]), .Z(n49) );
  IV U58 ( .A(B[210]), .Z(n48) );
  IV U59 ( .A(B[211]), .Z(n47) );
  IV U60 ( .A(B[212]), .Z(n46) );
  IV U61 ( .A(B[213]), .Z(n45) );
  IV U62 ( .A(B[214]), .Z(n44) );
  IV U63 ( .A(B[215]), .Z(n43) );
  IV U64 ( .A(B[216]), .Z(n42) );
  IV U65 ( .A(B[217]), .Z(n41) );
  IV U66 ( .A(B[218]), .Z(n40) );
  IV U67 ( .A(B[254]), .Z(n4) );
  IV U68 ( .A(B[219]), .Z(n39) );
  IV U69 ( .A(B[220]), .Z(n38) );
  IV U70 ( .A(B[221]), .Z(n37) );
  IV U71 ( .A(B[222]), .Z(n36) );
  IV U72 ( .A(B[223]), .Z(n35) );
  IV U73 ( .A(B[224]), .Z(n34) );
  IV U74 ( .A(B[225]), .Z(n33) );
  IV U75 ( .A(B[226]), .Z(n32) );
  IV U76 ( .A(B[227]), .Z(n31) );
  IV U77 ( .A(B[228]), .Z(n30) );
  IV U78 ( .A(B[255]), .Z(n3) );
  IV U79 ( .A(B[229]), .Z(n29) );
  IV U80 ( .A(B[230]), .Z(n28) );
  IV U81 ( .A(B[231]), .Z(n27) );
  IV U82 ( .A(B[232]), .Z(n26) );
  IV U83 ( .A(B[0]), .Z(n258) );
  IV U84 ( .A(B[1]), .Z(n257) );
  IV U85 ( .A(B[2]), .Z(n256) );
  IV U86 ( .A(B[3]), .Z(n255) );
  IV U87 ( .A(B[4]), .Z(n254) );
  IV U88 ( .A(B[5]), .Z(n253) );
  IV U89 ( .A(B[6]), .Z(n252) );
  IV U90 ( .A(B[7]), .Z(n251) );
  IV U91 ( .A(B[8]), .Z(n250) );
  IV U92 ( .A(B[233]), .Z(n25) );
  IV U93 ( .A(B[9]), .Z(n249) );
  IV U94 ( .A(B[10]), .Z(n248) );
  IV U95 ( .A(B[11]), .Z(n247) );
  IV U96 ( .A(B[12]), .Z(n246) );
  IV U97 ( .A(B[13]), .Z(n245) );
  IV U98 ( .A(B[14]), .Z(n244) );
  IV U99 ( .A(B[15]), .Z(n243) );
  IV U100 ( .A(B[16]), .Z(n242) );
  IV U101 ( .A(B[17]), .Z(n241) );
  IV U102 ( .A(B[18]), .Z(n240) );
  IV U103 ( .A(B[234]), .Z(n24) );
  IV U104 ( .A(B[19]), .Z(n239) );
  IV U105 ( .A(B[20]), .Z(n238) );
  IV U106 ( .A(B[21]), .Z(n237) );
  IV U107 ( .A(B[22]), .Z(n236) );
  IV U108 ( .A(B[23]), .Z(n235) );
  IV U109 ( .A(B[24]), .Z(n234) );
  IV U110 ( .A(B[25]), .Z(n233) );
  IV U111 ( .A(B[26]), .Z(n232) );
  IV U112 ( .A(B[27]), .Z(n231) );
  IV U113 ( .A(B[28]), .Z(n230) );
  IV U114 ( .A(B[235]), .Z(n23) );
  IV U115 ( .A(B[29]), .Z(n229) );
  IV U116 ( .A(B[30]), .Z(n228) );
  IV U117 ( .A(B[31]), .Z(n227) );
  IV U118 ( .A(B[32]), .Z(n226) );
  IV U119 ( .A(B[33]), .Z(n225) );
  IV U120 ( .A(B[34]), .Z(n224) );
  IV U121 ( .A(B[35]), .Z(n223) );
  IV U122 ( .A(B[36]), .Z(n222) );
  IV U123 ( .A(B[37]), .Z(n221) );
  IV U124 ( .A(B[38]), .Z(n220) );
  IV U125 ( .A(B[236]), .Z(n22) );
  IV U126 ( .A(B[39]), .Z(n219) );
  IV U127 ( .A(B[40]), .Z(n218) );
  IV U128 ( .A(B[41]), .Z(n217) );
  IV U129 ( .A(B[42]), .Z(n216) );
  IV U130 ( .A(B[43]), .Z(n215) );
  IV U131 ( .A(B[44]), .Z(n214) );
  IV U132 ( .A(B[45]), .Z(n213) );
  IV U133 ( .A(B[46]), .Z(n212) );
  IV U134 ( .A(B[47]), .Z(n211) );
  IV U135 ( .A(B[48]), .Z(n210) );
  IV U136 ( .A(B[237]), .Z(n21) );
  IV U137 ( .A(B[49]), .Z(n209) );
  IV U138 ( .A(B[50]), .Z(n208) );
  IV U139 ( .A(B[51]), .Z(n207) );
  IV U140 ( .A(B[52]), .Z(n206) );
  IV U141 ( .A(B[53]), .Z(n205) );
  IV U142 ( .A(B[54]), .Z(n204) );
  IV U143 ( .A(B[55]), .Z(n203) );
  IV U144 ( .A(B[56]), .Z(n202) );
  IV U145 ( .A(B[57]), .Z(n201) );
  IV U146 ( .A(B[58]), .Z(n200) );
  IV U147 ( .A(B[238]), .Z(n20) );
  IV U148 ( .A(B[59]), .Z(n199) );
  IV U149 ( .A(B[60]), .Z(n198) );
  IV U150 ( .A(B[61]), .Z(n197) );
  IV U151 ( .A(B[62]), .Z(n196) );
  IV U152 ( .A(B[63]), .Z(n195) );
  IV U153 ( .A(B[64]), .Z(n194) );
  IV U154 ( .A(B[65]), .Z(n193) );
  IV U155 ( .A(B[66]), .Z(n192) );
  IV U156 ( .A(B[67]), .Z(n191) );
  IV U157 ( .A(B[68]), .Z(n190) );
  IV U158 ( .A(B[239]), .Z(n19) );
  IV U159 ( .A(B[69]), .Z(n189) );
  IV U160 ( .A(B[70]), .Z(n188) );
  IV U161 ( .A(B[71]), .Z(n187) );
  IV U162 ( .A(B[72]), .Z(n186) );
  IV U163 ( .A(B[73]), .Z(n185) );
  IV U164 ( .A(B[74]), .Z(n184) );
  IV U165 ( .A(B[75]), .Z(n183) );
  IV U166 ( .A(B[76]), .Z(n182) );
  IV U167 ( .A(B[77]), .Z(n181) );
  IV U168 ( .A(B[78]), .Z(n180) );
  IV U169 ( .A(B[240]), .Z(n18) );
  IV U170 ( .A(B[79]), .Z(n179) );
  IV U171 ( .A(B[80]), .Z(n178) );
  IV U172 ( .A(B[81]), .Z(n177) );
  IV U173 ( .A(B[82]), .Z(n176) );
  IV U174 ( .A(B[83]), .Z(n175) );
  IV U175 ( .A(B[84]), .Z(n174) );
  IV U176 ( .A(B[85]), .Z(n173) );
  IV U177 ( .A(B[86]), .Z(n172) );
  IV U178 ( .A(B[87]), .Z(n171) );
  IV U179 ( .A(B[88]), .Z(n170) );
  IV U180 ( .A(B[241]), .Z(n17) );
  IV U181 ( .A(B[89]), .Z(n169) );
  IV U182 ( .A(B[90]), .Z(n168) );
  IV U183 ( .A(B[91]), .Z(n167) );
  IV U184 ( .A(B[92]), .Z(n166) );
  IV U185 ( .A(B[93]), .Z(n165) );
  IV U186 ( .A(B[94]), .Z(n164) );
  IV U187 ( .A(B[95]), .Z(n163) );
  IV U188 ( .A(B[96]), .Z(n162) );
  IV U189 ( .A(B[97]), .Z(n161) );
  IV U190 ( .A(B[98]), .Z(n160) );
  IV U191 ( .A(B[242]), .Z(n16) );
  IV U192 ( .A(B[99]), .Z(n159) );
  IV U193 ( .A(B[100]), .Z(n158) );
  IV U194 ( .A(B[101]), .Z(n157) );
  IV U195 ( .A(B[102]), .Z(n156) );
  IV U196 ( .A(B[103]), .Z(n155) );
  IV U197 ( .A(B[104]), .Z(n154) );
  IV U198 ( .A(B[105]), .Z(n153) );
  IV U199 ( .A(B[106]), .Z(n152) );
  IV U200 ( .A(B[107]), .Z(n151) );
  IV U201 ( .A(B[108]), .Z(n150) );
  IV U202 ( .A(B[243]), .Z(n15) );
  IV U203 ( .A(B[109]), .Z(n149) );
  IV U204 ( .A(B[110]), .Z(n148) );
  IV U205 ( .A(B[111]), .Z(n147) );
  IV U206 ( .A(B[112]), .Z(n146) );
  IV U207 ( .A(B[113]), .Z(n145) );
  IV U208 ( .A(B[114]), .Z(n144) );
  IV U209 ( .A(B[115]), .Z(n143) );
  IV U210 ( .A(B[116]), .Z(n142) );
  IV U211 ( .A(B[117]), .Z(n141) );
  IV U212 ( .A(B[118]), .Z(n140) );
  IV U213 ( .A(B[244]), .Z(n14) );
  IV U214 ( .A(B[119]), .Z(n139) );
  IV U215 ( .A(B[120]), .Z(n138) );
  IV U216 ( .A(B[121]), .Z(n137) );
  IV U217 ( .A(B[122]), .Z(n136) );
  IV U218 ( .A(B[123]), .Z(n135) );
  IV U219 ( .A(B[124]), .Z(n134) );
  IV U220 ( .A(B[125]), .Z(n133) );
  IV U221 ( .A(B[126]), .Z(n132) );
  IV U222 ( .A(B[127]), .Z(n131) );
  IV U223 ( .A(B[128]), .Z(n130) );
  IV U224 ( .A(B[245]), .Z(n13) );
  IV U225 ( .A(B[129]), .Z(n129) );
  IV U226 ( .A(B[130]), .Z(n128) );
  IV U227 ( .A(B[131]), .Z(n127) );
  IV U228 ( .A(B[132]), .Z(n126) );
  IV U229 ( .A(B[133]), .Z(n125) );
  IV U230 ( .A(B[134]), .Z(n124) );
  IV U231 ( .A(B[135]), .Z(n123) );
  IV U232 ( .A(B[136]), .Z(n122) );
  IV U233 ( .A(B[137]), .Z(n121) );
  IV U234 ( .A(B[138]), .Z(n120) );
  IV U235 ( .A(B[246]), .Z(n12) );
  IV U236 ( .A(B[139]), .Z(n119) );
  IV U237 ( .A(B[140]), .Z(n118) );
  IV U238 ( .A(B[141]), .Z(n117) );
  IV U239 ( .A(B[142]), .Z(n116) );
  IV U240 ( .A(B[143]), .Z(n115) );
  IV U241 ( .A(B[144]), .Z(n114) );
  IV U242 ( .A(B[145]), .Z(n113) );
  IV U243 ( .A(B[146]), .Z(n112) );
  IV U244 ( .A(B[147]), .Z(n111) );
  IV U245 ( .A(B[148]), .Z(n110) );
  IV U246 ( .A(B[247]), .Z(n11) );
  IV U247 ( .A(B[149]), .Z(n109) );
  IV U248 ( .A(B[150]), .Z(n108) );
  IV U249 ( .A(B[151]), .Z(n107) );
  IV U250 ( .A(B[152]), .Z(n106) );
  IV U251 ( .A(B[153]), .Z(n105) );
  IV U252 ( .A(B[154]), .Z(n104) );
  IV U253 ( .A(B[155]), .Z(n103) );
  IV U254 ( .A(B[156]), .Z(n102) );
  IV U255 ( .A(B[157]), .Z(n101) );
  IV U256 ( .A(B[158]), .Z(n100) );
  IV U257 ( .A(B[248]), .Z(n10) );
endmodule


module MUX_N258_7 ( A, B, S, O );
  input [257:0] A;
  input [257:0] B;
  output [257:0] O;
  input S;


  ANDN U1 ( .B(A[9]), .A(S), .Z(O[9]) );
  ANDN U2 ( .B(A[99]), .A(S), .Z(O[99]) );
  ANDN U3 ( .B(A[98]), .A(S), .Z(O[98]) );
  ANDN U4 ( .B(A[97]), .A(S), .Z(O[97]) );
  ANDN U5 ( .B(A[96]), .A(S), .Z(O[96]) );
  ANDN U6 ( .B(A[95]), .A(S), .Z(O[95]) );
  ANDN U7 ( .B(A[94]), .A(S), .Z(O[94]) );
  ANDN U8 ( .B(A[93]), .A(S), .Z(O[93]) );
  ANDN U9 ( .B(A[92]), .A(S), .Z(O[92]) );
  ANDN U10 ( .B(A[91]), .A(S), .Z(O[91]) );
  ANDN U11 ( .B(A[90]), .A(S), .Z(O[90]) );
  ANDN U12 ( .B(A[8]), .A(S), .Z(O[8]) );
  ANDN U13 ( .B(A[89]), .A(S), .Z(O[89]) );
  ANDN U14 ( .B(A[88]), .A(S), .Z(O[88]) );
  ANDN U15 ( .B(A[87]), .A(S), .Z(O[87]) );
  ANDN U16 ( .B(A[86]), .A(S), .Z(O[86]) );
  ANDN U17 ( .B(A[85]), .A(S), .Z(O[85]) );
  ANDN U18 ( .B(A[84]), .A(S), .Z(O[84]) );
  ANDN U19 ( .B(A[83]), .A(S), .Z(O[83]) );
  ANDN U20 ( .B(A[82]), .A(S), .Z(O[82]) );
  ANDN U21 ( .B(A[81]), .A(S), .Z(O[81]) );
  ANDN U22 ( .B(A[80]), .A(S), .Z(O[80]) );
  ANDN U23 ( .B(A[7]), .A(S), .Z(O[7]) );
  ANDN U24 ( .B(A[79]), .A(S), .Z(O[79]) );
  ANDN U25 ( .B(A[78]), .A(S), .Z(O[78]) );
  ANDN U26 ( .B(A[77]), .A(S), .Z(O[77]) );
  ANDN U27 ( .B(A[76]), .A(S), .Z(O[76]) );
  ANDN U28 ( .B(A[75]), .A(S), .Z(O[75]) );
  ANDN U29 ( .B(A[74]), .A(S), .Z(O[74]) );
  ANDN U30 ( .B(A[73]), .A(S), .Z(O[73]) );
  ANDN U31 ( .B(A[72]), .A(S), .Z(O[72]) );
  ANDN U32 ( .B(A[71]), .A(S), .Z(O[71]) );
  ANDN U33 ( .B(A[70]), .A(S), .Z(O[70]) );
  ANDN U34 ( .B(A[6]), .A(S), .Z(O[6]) );
  ANDN U35 ( .B(A[69]), .A(S), .Z(O[69]) );
  ANDN U36 ( .B(A[68]), .A(S), .Z(O[68]) );
  ANDN U37 ( .B(A[67]), .A(S), .Z(O[67]) );
  ANDN U38 ( .B(A[66]), .A(S), .Z(O[66]) );
  ANDN U39 ( .B(A[65]), .A(S), .Z(O[65]) );
  ANDN U40 ( .B(A[64]), .A(S), .Z(O[64]) );
  ANDN U41 ( .B(A[63]), .A(S), .Z(O[63]) );
  ANDN U42 ( .B(A[62]), .A(S), .Z(O[62]) );
  ANDN U43 ( .B(A[61]), .A(S), .Z(O[61]) );
  ANDN U44 ( .B(A[60]), .A(S), .Z(O[60]) );
  ANDN U45 ( .B(A[5]), .A(S), .Z(O[5]) );
  ANDN U46 ( .B(A[59]), .A(S), .Z(O[59]) );
  ANDN U47 ( .B(A[58]), .A(S), .Z(O[58]) );
  ANDN U48 ( .B(A[57]), .A(S), .Z(O[57]) );
  ANDN U49 ( .B(A[56]), .A(S), .Z(O[56]) );
  ANDN U50 ( .B(A[55]), .A(S), .Z(O[55]) );
  ANDN U51 ( .B(A[54]), .A(S), .Z(O[54]) );
  ANDN U52 ( .B(A[53]), .A(S), .Z(O[53]) );
  ANDN U53 ( .B(A[52]), .A(S), .Z(O[52]) );
  ANDN U54 ( .B(A[51]), .A(S), .Z(O[51]) );
  ANDN U55 ( .B(A[50]), .A(S), .Z(O[50]) );
  ANDN U56 ( .B(A[4]), .A(S), .Z(O[4]) );
  ANDN U57 ( .B(A[49]), .A(S), .Z(O[49]) );
  ANDN U58 ( .B(A[48]), .A(S), .Z(O[48]) );
  ANDN U59 ( .B(A[47]), .A(S), .Z(O[47]) );
  ANDN U60 ( .B(A[46]), .A(S), .Z(O[46]) );
  ANDN U61 ( .B(A[45]), .A(S), .Z(O[45]) );
  ANDN U62 ( .B(A[44]), .A(S), .Z(O[44]) );
  ANDN U63 ( .B(A[43]), .A(S), .Z(O[43]) );
  ANDN U64 ( .B(A[42]), .A(S), .Z(O[42]) );
  ANDN U65 ( .B(A[41]), .A(S), .Z(O[41]) );
  ANDN U66 ( .B(A[40]), .A(S), .Z(O[40]) );
  ANDN U67 ( .B(A[3]), .A(S), .Z(O[3]) );
  ANDN U68 ( .B(A[39]), .A(S), .Z(O[39]) );
  ANDN U69 ( .B(A[38]), .A(S), .Z(O[38]) );
  ANDN U70 ( .B(A[37]), .A(S), .Z(O[37]) );
  ANDN U71 ( .B(A[36]), .A(S), .Z(O[36]) );
  ANDN U72 ( .B(A[35]), .A(S), .Z(O[35]) );
  ANDN U73 ( .B(A[34]), .A(S), .Z(O[34]) );
  ANDN U74 ( .B(A[33]), .A(S), .Z(O[33]) );
  ANDN U75 ( .B(A[32]), .A(S), .Z(O[32]) );
  ANDN U76 ( .B(A[31]), .A(S), .Z(O[31]) );
  ANDN U77 ( .B(A[30]), .A(S), .Z(O[30]) );
  ANDN U78 ( .B(A[2]), .A(S), .Z(O[2]) );
  ANDN U79 ( .B(A[29]), .A(S), .Z(O[29]) );
  ANDN U80 ( .B(A[28]), .A(S), .Z(O[28]) );
  ANDN U81 ( .B(A[27]), .A(S), .Z(O[27]) );
  ANDN U82 ( .B(A[26]), .A(S), .Z(O[26]) );
  ANDN U83 ( .B(A[25]), .A(S), .Z(O[25]) );
  ANDN U84 ( .B(A[255]), .A(S), .Z(O[255]) );
  ANDN U85 ( .B(A[254]), .A(S), .Z(O[254]) );
  ANDN U86 ( .B(A[253]), .A(S), .Z(O[253]) );
  ANDN U87 ( .B(A[252]), .A(S), .Z(O[252]) );
  ANDN U88 ( .B(A[251]), .A(S), .Z(O[251]) );
  ANDN U89 ( .B(A[250]), .A(S), .Z(O[250]) );
  ANDN U90 ( .B(A[24]), .A(S), .Z(O[24]) );
  ANDN U91 ( .B(A[249]), .A(S), .Z(O[249]) );
  ANDN U92 ( .B(A[248]), .A(S), .Z(O[248]) );
  ANDN U93 ( .B(A[247]), .A(S), .Z(O[247]) );
  ANDN U94 ( .B(A[246]), .A(S), .Z(O[246]) );
  ANDN U95 ( .B(A[245]), .A(S), .Z(O[245]) );
  ANDN U96 ( .B(A[244]), .A(S), .Z(O[244]) );
  ANDN U97 ( .B(A[243]), .A(S), .Z(O[243]) );
  ANDN U98 ( .B(A[242]), .A(S), .Z(O[242]) );
  ANDN U99 ( .B(A[241]), .A(S), .Z(O[241]) );
  ANDN U100 ( .B(A[240]), .A(S), .Z(O[240]) );
  ANDN U101 ( .B(A[23]), .A(S), .Z(O[23]) );
  ANDN U102 ( .B(A[239]), .A(S), .Z(O[239]) );
  ANDN U103 ( .B(A[238]), .A(S), .Z(O[238]) );
  ANDN U104 ( .B(A[237]), .A(S), .Z(O[237]) );
  ANDN U105 ( .B(A[236]), .A(S), .Z(O[236]) );
  ANDN U106 ( .B(A[235]), .A(S), .Z(O[235]) );
  ANDN U107 ( .B(A[234]), .A(S), .Z(O[234]) );
  ANDN U108 ( .B(A[233]), .A(S), .Z(O[233]) );
  ANDN U109 ( .B(A[232]), .A(S), .Z(O[232]) );
  ANDN U110 ( .B(A[231]), .A(S), .Z(O[231]) );
  ANDN U111 ( .B(A[230]), .A(S), .Z(O[230]) );
  ANDN U112 ( .B(A[22]), .A(S), .Z(O[22]) );
  ANDN U113 ( .B(A[229]), .A(S), .Z(O[229]) );
  ANDN U114 ( .B(A[228]), .A(S), .Z(O[228]) );
  ANDN U115 ( .B(A[227]), .A(S), .Z(O[227]) );
  ANDN U116 ( .B(A[226]), .A(S), .Z(O[226]) );
  ANDN U117 ( .B(A[225]), .A(S), .Z(O[225]) );
  ANDN U118 ( .B(A[224]), .A(S), .Z(O[224]) );
  ANDN U119 ( .B(A[223]), .A(S), .Z(O[223]) );
  ANDN U120 ( .B(A[222]), .A(S), .Z(O[222]) );
  ANDN U121 ( .B(A[221]), .A(S), .Z(O[221]) );
  ANDN U122 ( .B(A[220]), .A(S), .Z(O[220]) );
  ANDN U123 ( .B(A[21]), .A(S), .Z(O[21]) );
  ANDN U124 ( .B(A[219]), .A(S), .Z(O[219]) );
  ANDN U125 ( .B(A[218]), .A(S), .Z(O[218]) );
  ANDN U126 ( .B(A[217]), .A(S), .Z(O[217]) );
  ANDN U127 ( .B(A[216]), .A(S), .Z(O[216]) );
  ANDN U128 ( .B(A[215]), .A(S), .Z(O[215]) );
  ANDN U129 ( .B(A[214]), .A(S), .Z(O[214]) );
  ANDN U130 ( .B(A[213]), .A(S), .Z(O[213]) );
  ANDN U131 ( .B(A[212]), .A(S), .Z(O[212]) );
  ANDN U132 ( .B(A[211]), .A(S), .Z(O[211]) );
  ANDN U133 ( .B(A[210]), .A(S), .Z(O[210]) );
  ANDN U134 ( .B(A[20]), .A(S), .Z(O[20]) );
  ANDN U135 ( .B(A[209]), .A(S), .Z(O[209]) );
  ANDN U136 ( .B(A[208]), .A(S), .Z(O[208]) );
  ANDN U137 ( .B(A[207]), .A(S), .Z(O[207]) );
  ANDN U138 ( .B(A[206]), .A(S), .Z(O[206]) );
  ANDN U139 ( .B(A[205]), .A(S), .Z(O[205]) );
  ANDN U140 ( .B(A[204]), .A(S), .Z(O[204]) );
  ANDN U141 ( .B(A[203]), .A(S), .Z(O[203]) );
  ANDN U142 ( .B(A[202]), .A(S), .Z(O[202]) );
  ANDN U143 ( .B(A[201]), .A(S), .Z(O[201]) );
  ANDN U144 ( .B(A[200]), .A(S), .Z(O[200]) );
  ANDN U145 ( .B(A[1]), .A(S), .Z(O[1]) );
  ANDN U146 ( .B(A[19]), .A(S), .Z(O[19]) );
  ANDN U147 ( .B(A[199]), .A(S), .Z(O[199]) );
  ANDN U148 ( .B(A[198]), .A(S), .Z(O[198]) );
  ANDN U149 ( .B(A[197]), .A(S), .Z(O[197]) );
  ANDN U150 ( .B(A[196]), .A(S), .Z(O[196]) );
  ANDN U151 ( .B(A[195]), .A(S), .Z(O[195]) );
  ANDN U152 ( .B(A[194]), .A(S), .Z(O[194]) );
  ANDN U153 ( .B(A[193]), .A(S), .Z(O[193]) );
  ANDN U154 ( .B(A[192]), .A(S), .Z(O[192]) );
  ANDN U155 ( .B(A[191]), .A(S), .Z(O[191]) );
  ANDN U156 ( .B(A[190]), .A(S), .Z(O[190]) );
  ANDN U157 ( .B(A[18]), .A(S), .Z(O[18]) );
  ANDN U158 ( .B(A[189]), .A(S), .Z(O[189]) );
  ANDN U159 ( .B(A[188]), .A(S), .Z(O[188]) );
  ANDN U160 ( .B(A[187]), .A(S), .Z(O[187]) );
  ANDN U161 ( .B(A[186]), .A(S), .Z(O[186]) );
  ANDN U162 ( .B(A[185]), .A(S), .Z(O[185]) );
  ANDN U163 ( .B(A[184]), .A(S), .Z(O[184]) );
  ANDN U164 ( .B(A[183]), .A(S), .Z(O[183]) );
  ANDN U165 ( .B(A[182]), .A(S), .Z(O[182]) );
  ANDN U166 ( .B(A[181]), .A(S), .Z(O[181]) );
  ANDN U167 ( .B(A[180]), .A(S), .Z(O[180]) );
  ANDN U168 ( .B(A[17]), .A(S), .Z(O[17]) );
  ANDN U169 ( .B(A[179]), .A(S), .Z(O[179]) );
  ANDN U170 ( .B(A[178]), .A(S), .Z(O[178]) );
  ANDN U171 ( .B(A[177]), .A(S), .Z(O[177]) );
  ANDN U172 ( .B(A[176]), .A(S), .Z(O[176]) );
  ANDN U173 ( .B(A[175]), .A(S), .Z(O[175]) );
  ANDN U174 ( .B(A[174]), .A(S), .Z(O[174]) );
  ANDN U175 ( .B(A[173]), .A(S), .Z(O[173]) );
  ANDN U176 ( .B(A[172]), .A(S), .Z(O[172]) );
  ANDN U177 ( .B(A[171]), .A(S), .Z(O[171]) );
  ANDN U178 ( .B(A[170]), .A(S), .Z(O[170]) );
  ANDN U179 ( .B(A[16]), .A(S), .Z(O[16]) );
  ANDN U180 ( .B(A[169]), .A(S), .Z(O[169]) );
  ANDN U181 ( .B(A[168]), .A(S), .Z(O[168]) );
  ANDN U182 ( .B(A[167]), .A(S), .Z(O[167]) );
  ANDN U183 ( .B(A[166]), .A(S), .Z(O[166]) );
  ANDN U184 ( .B(A[165]), .A(S), .Z(O[165]) );
  ANDN U185 ( .B(A[164]), .A(S), .Z(O[164]) );
  ANDN U186 ( .B(A[163]), .A(S), .Z(O[163]) );
  ANDN U187 ( .B(A[162]), .A(S), .Z(O[162]) );
  ANDN U188 ( .B(A[161]), .A(S), .Z(O[161]) );
  ANDN U189 ( .B(A[160]), .A(S), .Z(O[160]) );
  ANDN U190 ( .B(A[15]), .A(S), .Z(O[15]) );
  ANDN U191 ( .B(A[159]), .A(S), .Z(O[159]) );
  ANDN U192 ( .B(A[158]), .A(S), .Z(O[158]) );
  ANDN U193 ( .B(A[157]), .A(S), .Z(O[157]) );
  ANDN U194 ( .B(A[156]), .A(S), .Z(O[156]) );
  ANDN U195 ( .B(A[155]), .A(S), .Z(O[155]) );
  ANDN U196 ( .B(A[154]), .A(S), .Z(O[154]) );
  ANDN U197 ( .B(A[153]), .A(S), .Z(O[153]) );
  ANDN U198 ( .B(A[152]), .A(S), .Z(O[152]) );
  ANDN U199 ( .B(A[151]), .A(S), .Z(O[151]) );
  ANDN U200 ( .B(A[150]), .A(S), .Z(O[150]) );
  ANDN U201 ( .B(A[14]), .A(S), .Z(O[14]) );
  ANDN U202 ( .B(A[149]), .A(S), .Z(O[149]) );
  ANDN U203 ( .B(A[148]), .A(S), .Z(O[148]) );
  ANDN U204 ( .B(A[147]), .A(S), .Z(O[147]) );
  ANDN U205 ( .B(A[146]), .A(S), .Z(O[146]) );
  ANDN U206 ( .B(A[145]), .A(S), .Z(O[145]) );
  ANDN U207 ( .B(A[144]), .A(S), .Z(O[144]) );
  ANDN U208 ( .B(A[143]), .A(S), .Z(O[143]) );
  ANDN U209 ( .B(A[142]), .A(S), .Z(O[142]) );
  ANDN U210 ( .B(A[141]), .A(S), .Z(O[141]) );
  ANDN U211 ( .B(A[140]), .A(S), .Z(O[140]) );
  ANDN U212 ( .B(A[13]), .A(S), .Z(O[13]) );
  ANDN U213 ( .B(A[139]), .A(S), .Z(O[139]) );
  ANDN U214 ( .B(A[138]), .A(S), .Z(O[138]) );
  ANDN U215 ( .B(A[137]), .A(S), .Z(O[137]) );
  ANDN U216 ( .B(A[136]), .A(S), .Z(O[136]) );
  ANDN U217 ( .B(A[135]), .A(S), .Z(O[135]) );
  ANDN U218 ( .B(A[134]), .A(S), .Z(O[134]) );
  ANDN U219 ( .B(A[133]), .A(S), .Z(O[133]) );
  ANDN U220 ( .B(A[132]), .A(S), .Z(O[132]) );
  ANDN U221 ( .B(A[131]), .A(S), .Z(O[131]) );
  ANDN U222 ( .B(A[130]), .A(S), .Z(O[130]) );
  ANDN U223 ( .B(A[12]), .A(S), .Z(O[12]) );
  ANDN U224 ( .B(A[129]), .A(S), .Z(O[129]) );
  ANDN U225 ( .B(A[128]), .A(S), .Z(O[128]) );
  ANDN U226 ( .B(A[127]), .A(S), .Z(O[127]) );
  ANDN U227 ( .B(A[126]), .A(S), .Z(O[126]) );
  ANDN U228 ( .B(A[125]), .A(S), .Z(O[125]) );
  ANDN U229 ( .B(A[124]), .A(S), .Z(O[124]) );
  ANDN U230 ( .B(A[123]), .A(S), .Z(O[123]) );
  ANDN U231 ( .B(A[122]), .A(S), .Z(O[122]) );
  ANDN U232 ( .B(A[121]), .A(S), .Z(O[121]) );
  ANDN U233 ( .B(A[120]), .A(S), .Z(O[120]) );
  ANDN U234 ( .B(A[11]), .A(S), .Z(O[11]) );
  ANDN U235 ( .B(A[119]), .A(S), .Z(O[119]) );
  ANDN U236 ( .B(A[118]), .A(S), .Z(O[118]) );
  ANDN U237 ( .B(A[117]), .A(S), .Z(O[117]) );
  ANDN U238 ( .B(A[116]), .A(S), .Z(O[116]) );
  ANDN U239 ( .B(A[115]), .A(S), .Z(O[115]) );
  ANDN U240 ( .B(A[114]), .A(S), .Z(O[114]) );
  ANDN U241 ( .B(A[113]), .A(S), .Z(O[113]) );
  ANDN U242 ( .B(A[112]), .A(S), .Z(O[112]) );
  ANDN U243 ( .B(A[111]), .A(S), .Z(O[111]) );
  ANDN U244 ( .B(A[110]), .A(S), .Z(O[110]) );
  ANDN U245 ( .B(A[10]), .A(S), .Z(O[10]) );
  ANDN U246 ( .B(A[109]), .A(S), .Z(O[109]) );
  ANDN U247 ( .B(A[108]), .A(S), .Z(O[108]) );
  ANDN U248 ( .B(A[107]), .A(S), .Z(O[107]) );
  ANDN U249 ( .B(A[106]), .A(S), .Z(O[106]) );
  ANDN U250 ( .B(A[105]), .A(S), .Z(O[105]) );
  ANDN U251 ( .B(A[104]), .A(S), .Z(O[104]) );
  ANDN U252 ( .B(A[103]), .A(S), .Z(O[103]) );
  ANDN U253 ( .B(A[102]), .A(S), .Z(O[102]) );
  ANDN U254 ( .B(A[101]), .A(S), .Z(O[101]) );
  ANDN U255 ( .B(A[100]), .A(S), .Z(O[100]) );
  ANDN U256 ( .B(A[0]), .A(S), .Z(O[0]) );
endmodule


module MUX_N258_8 ( A, B, S, O );
  input [257:0] A;
  input [257:0] B;
  output [257:0] O;
  input S;


  ANDN U1 ( .B(A[9]), .A(S), .Z(O[9]) );
  ANDN U2 ( .B(A[99]), .A(S), .Z(O[99]) );
  ANDN U3 ( .B(A[98]), .A(S), .Z(O[98]) );
  ANDN U4 ( .B(A[97]), .A(S), .Z(O[97]) );
  ANDN U5 ( .B(A[96]), .A(S), .Z(O[96]) );
  ANDN U6 ( .B(A[95]), .A(S), .Z(O[95]) );
  ANDN U7 ( .B(A[94]), .A(S), .Z(O[94]) );
  ANDN U8 ( .B(A[93]), .A(S), .Z(O[93]) );
  ANDN U9 ( .B(A[92]), .A(S), .Z(O[92]) );
  ANDN U10 ( .B(A[91]), .A(S), .Z(O[91]) );
  ANDN U11 ( .B(A[90]), .A(S), .Z(O[90]) );
  ANDN U12 ( .B(A[8]), .A(S), .Z(O[8]) );
  ANDN U13 ( .B(A[89]), .A(S), .Z(O[89]) );
  ANDN U14 ( .B(A[88]), .A(S), .Z(O[88]) );
  ANDN U15 ( .B(A[87]), .A(S), .Z(O[87]) );
  ANDN U16 ( .B(A[86]), .A(S), .Z(O[86]) );
  ANDN U17 ( .B(A[85]), .A(S), .Z(O[85]) );
  ANDN U18 ( .B(A[84]), .A(S), .Z(O[84]) );
  ANDN U19 ( .B(A[83]), .A(S), .Z(O[83]) );
  ANDN U20 ( .B(A[82]), .A(S), .Z(O[82]) );
  ANDN U21 ( .B(A[81]), .A(S), .Z(O[81]) );
  ANDN U22 ( .B(A[80]), .A(S), .Z(O[80]) );
  ANDN U23 ( .B(A[7]), .A(S), .Z(O[7]) );
  ANDN U24 ( .B(A[79]), .A(S), .Z(O[79]) );
  ANDN U25 ( .B(A[78]), .A(S), .Z(O[78]) );
  ANDN U26 ( .B(A[77]), .A(S), .Z(O[77]) );
  ANDN U27 ( .B(A[76]), .A(S), .Z(O[76]) );
  ANDN U28 ( .B(A[75]), .A(S), .Z(O[75]) );
  ANDN U29 ( .B(A[74]), .A(S), .Z(O[74]) );
  ANDN U30 ( .B(A[73]), .A(S), .Z(O[73]) );
  ANDN U31 ( .B(A[72]), .A(S), .Z(O[72]) );
  ANDN U32 ( .B(A[71]), .A(S), .Z(O[71]) );
  ANDN U33 ( .B(A[70]), .A(S), .Z(O[70]) );
  ANDN U34 ( .B(A[6]), .A(S), .Z(O[6]) );
  ANDN U35 ( .B(A[69]), .A(S), .Z(O[69]) );
  ANDN U36 ( .B(A[68]), .A(S), .Z(O[68]) );
  ANDN U37 ( .B(A[67]), .A(S), .Z(O[67]) );
  ANDN U38 ( .B(A[66]), .A(S), .Z(O[66]) );
  ANDN U39 ( .B(A[65]), .A(S), .Z(O[65]) );
  ANDN U40 ( .B(A[64]), .A(S), .Z(O[64]) );
  ANDN U41 ( .B(A[63]), .A(S), .Z(O[63]) );
  ANDN U42 ( .B(A[62]), .A(S), .Z(O[62]) );
  ANDN U43 ( .B(A[61]), .A(S), .Z(O[61]) );
  ANDN U44 ( .B(A[60]), .A(S), .Z(O[60]) );
  ANDN U45 ( .B(A[5]), .A(S), .Z(O[5]) );
  ANDN U46 ( .B(A[59]), .A(S), .Z(O[59]) );
  ANDN U47 ( .B(A[58]), .A(S), .Z(O[58]) );
  ANDN U48 ( .B(A[57]), .A(S), .Z(O[57]) );
  ANDN U49 ( .B(A[56]), .A(S), .Z(O[56]) );
  ANDN U50 ( .B(A[55]), .A(S), .Z(O[55]) );
  ANDN U51 ( .B(A[54]), .A(S), .Z(O[54]) );
  ANDN U52 ( .B(A[53]), .A(S), .Z(O[53]) );
  ANDN U53 ( .B(A[52]), .A(S), .Z(O[52]) );
  ANDN U54 ( .B(A[51]), .A(S), .Z(O[51]) );
  ANDN U55 ( .B(A[50]), .A(S), .Z(O[50]) );
  ANDN U56 ( .B(A[4]), .A(S), .Z(O[4]) );
  ANDN U57 ( .B(A[49]), .A(S), .Z(O[49]) );
  ANDN U58 ( .B(A[48]), .A(S), .Z(O[48]) );
  ANDN U59 ( .B(A[47]), .A(S), .Z(O[47]) );
  ANDN U60 ( .B(A[46]), .A(S), .Z(O[46]) );
  ANDN U61 ( .B(A[45]), .A(S), .Z(O[45]) );
  ANDN U62 ( .B(A[44]), .A(S), .Z(O[44]) );
  ANDN U63 ( .B(A[43]), .A(S), .Z(O[43]) );
  ANDN U64 ( .B(A[42]), .A(S), .Z(O[42]) );
  ANDN U65 ( .B(A[41]), .A(S), .Z(O[41]) );
  ANDN U66 ( .B(A[40]), .A(S), .Z(O[40]) );
  ANDN U67 ( .B(A[3]), .A(S), .Z(O[3]) );
  ANDN U68 ( .B(A[39]), .A(S), .Z(O[39]) );
  ANDN U69 ( .B(A[38]), .A(S), .Z(O[38]) );
  ANDN U70 ( .B(A[37]), .A(S), .Z(O[37]) );
  ANDN U71 ( .B(A[36]), .A(S), .Z(O[36]) );
  ANDN U72 ( .B(A[35]), .A(S), .Z(O[35]) );
  ANDN U73 ( .B(A[34]), .A(S), .Z(O[34]) );
  ANDN U74 ( .B(A[33]), .A(S), .Z(O[33]) );
  ANDN U75 ( .B(A[32]), .A(S), .Z(O[32]) );
  ANDN U76 ( .B(A[31]), .A(S), .Z(O[31]) );
  ANDN U77 ( .B(A[30]), .A(S), .Z(O[30]) );
  ANDN U78 ( .B(A[2]), .A(S), .Z(O[2]) );
  ANDN U79 ( .B(A[29]), .A(S), .Z(O[29]) );
  ANDN U80 ( .B(A[28]), .A(S), .Z(O[28]) );
  ANDN U81 ( .B(A[27]), .A(S), .Z(O[27]) );
  ANDN U82 ( .B(A[26]), .A(S), .Z(O[26]) );
  ANDN U83 ( .B(A[25]), .A(S), .Z(O[25]) );
  ANDN U84 ( .B(A[255]), .A(S), .Z(O[255]) );
  ANDN U85 ( .B(A[254]), .A(S), .Z(O[254]) );
  ANDN U86 ( .B(A[253]), .A(S), .Z(O[253]) );
  ANDN U87 ( .B(A[252]), .A(S), .Z(O[252]) );
  ANDN U88 ( .B(A[251]), .A(S), .Z(O[251]) );
  ANDN U89 ( .B(A[250]), .A(S), .Z(O[250]) );
  ANDN U90 ( .B(A[24]), .A(S), .Z(O[24]) );
  ANDN U91 ( .B(A[249]), .A(S), .Z(O[249]) );
  ANDN U92 ( .B(A[248]), .A(S), .Z(O[248]) );
  ANDN U93 ( .B(A[247]), .A(S), .Z(O[247]) );
  ANDN U94 ( .B(A[246]), .A(S), .Z(O[246]) );
  ANDN U95 ( .B(A[245]), .A(S), .Z(O[245]) );
  ANDN U96 ( .B(A[244]), .A(S), .Z(O[244]) );
  ANDN U97 ( .B(A[243]), .A(S), .Z(O[243]) );
  ANDN U98 ( .B(A[242]), .A(S), .Z(O[242]) );
  ANDN U99 ( .B(A[241]), .A(S), .Z(O[241]) );
  ANDN U100 ( .B(A[240]), .A(S), .Z(O[240]) );
  ANDN U101 ( .B(A[23]), .A(S), .Z(O[23]) );
  ANDN U102 ( .B(A[239]), .A(S), .Z(O[239]) );
  ANDN U103 ( .B(A[238]), .A(S), .Z(O[238]) );
  ANDN U104 ( .B(A[237]), .A(S), .Z(O[237]) );
  ANDN U105 ( .B(A[236]), .A(S), .Z(O[236]) );
  ANDN U106 ( .B(A[235]), .A(S), .Z(O[235]) );
  ANDN U107 ( .B(A[234]), .A(S), .Z(O[234]) );
  ANDN U108 ( .B(A[233]), .A(S), .Z(O[233]) );
  ANDN U109 ( .B(A[232]), .A(S), .Z(O[232]) );
  ANDN U110 ( .B(A[231]), .A(S), .Z(O[231]) );
  ANDN U111 ( .B(A[230]), .A(S), .Z(O[230]) );
  ANDN U112 ( .B(A[22]), .A(S), .Z(O[22]) );
  ANDN U113 ( .B(A[229]), .A(S), .Z(O[229]) );
  ANDN U114 ( .B(A[228]), .A(S), .Z(O[228]) );
  ANDN U115 ( .B(A[227]), .A(S), .Z(O[227]) );
  ANDN U116 ( .B(A[226]), .A(S), .Z(O[226]) );
  ANDN U117 ( .B(A[225]), .A(S), .Z(O[225]) );
  ANDN U118 ( .B(A[224]), .A(S), .Z(O[224]) );
  ANDN U119 ( .B(A[223]), .A(S), .Z(O[223]) );
  ANDN U120 ( .B(A[222]), .A(S), .Z(O[222]) );
  ANDN U121 ( .B(A[221]), .A(S), .Z(O[221]) );
  ANDN U122 ( .B(A[220]), .A(S), .Z(O[220]) );
  ANDN U123 ( .B(A[21]), .A(S), .Z(O[21]) );
  ANDN U124 ( .B(A[219]), .A(S), .Z(O[219]) );
  ANDN U125 ( .B(A[218]), .A(S), .Z(O[218]) );
  ANDN U126 ( .B(A[217]), .A(S), .Z(O[217]) );
  ANDN U127 ( .B(A[216]), .A(S), .Z(O[216]) );
  ANDN U128 ( .B(A[215]), .A(S), .Z(O[215]) );
  ANDN U129 ( .B(A[214]), .A(S), .Z(O[214]) );
  ANDN U130 ( .B(A[213]), .A(S), .Z(O[213]) );
  ANDN U131 ( .B(A[212]), .A(S), .Z(O[212]) );
  ANDN U132 ( .B(A[211]), .A(S), .Z(O[211]) );
  ANDN U133 ( .B(A[210]), .A(S), .Z(O[210]) );
  ANDN U134 ( .B(A[20]), .A(S), .Z(O[20]) );
  ANDN U135 ( .B(A[209]), .A(S), .Z(O[209]) );
  ANDN U136 ( .B(A[208]), .A(S), .Z(O[208]) );
  ANDN U137 ( .B(A[207]), .A(S), .Z(O[207]) );
  ANDN U138 ( .B(A[206]), .A(S), .Z(O[206]) );
  ANDN U139 ( .B(A[205]), .A(S), .Z(O[205]) );
  ANDN U140 ( .B(A[204]), .A(S), .Z(O[204]) );
  ANDN U141 ( .B(A[203]), .A(S), .Z(O[203]) );
  ANDN U142 ( .B(A[202]), .A(S), .Z(O[202]) );
  ANDN U143 ( .B(A[201]), .A(S), .Z(O[201]) );
  ANDN U144 ( .B(A[200]), .A(S), .Z(O[200]) );
  ANDN U145 ( .B(A[1]), .A(S), .Z(O[1]) );
  ANDN U146 ( .B(A[19]), .A(S), .Z(O[19]) );
  ANDN U147 ( .B(A[199]), .A(S), .Z(O[199]) );
  ANDN U148 ( .B(A[198]), .A(S), .Z(O[198]) );
  ANDN U149 ( .B(A[197]), .A(S), .Z(O[197]) );
  ANDN U150 ( .B(A[196]), .A(S), .Z(O[196]) );
  ANDN U151 ( .B(A[195]), .A(S), .Z(O[195]) );
  ANDN U152 ( .B(A[194]), .A(S), .Z(O[194]) );
  ANDN U153 ( .B(A[193]), .A(S), .Z(O[193]) );
  ANDN U154 ( .B(A[192]), .A(S), .Z(O[192]) );
  ANDN U155 ( .B(A[191]), .A(S), .Z(O[191]) );
  ANDN U156 ( .B(A[190]), .A(S), .Z(O[190]) );
  ANDN U157 ( .B(A[18]), .A(S), .Z(O[18]) );
  ANDN U158 ( .B(A[189]), .A(S), .Z(O[189]) );
  ANDN U159 ( .B(A[188]), .A(S), .Z(O[188]) );
  ANDN U160 ( .B(A[187]), .A(S), .Z(O[187]) );
  ANDN U161 ( .B(A[186]), .A(S), .Z(O[186]) );
  ANDN U162 ( .B(A[185]), .A(S), .Z(O[185]) );
  ANDN U163 ( .B(A[184]), .A(S), .Z(O[184]) );
  ANDN U164 ( .B(A[183]), .A(S), .Z(O[183]) );
  ANDN U165 ( .B(A[182]), .A(S), .Z(O[182]) );
  ANDN U166 ( .B(A[181]), .A(S), .Z(O[181]) );
  ANDN U167 ( .B(A[180]), .A(S), .Z(O[180]) );
  ANDN U168 ( .B(A[17]), .A(S), .Z(O[17]) );
  ANDN U169 ( .B(A[179]), .A(S), .Z(O[179]) );
  ANDN U170 ( .B(A[178]), .A(S), .Z(O[178]) );
  ANDN U171 ( .B(A[177]), .A(S), .Z(O[177]) );
  ANDN U172 ( .B(A[176]), .A(S), .Z(O[176]) );
  ANDN U173 ( .B(A[175]), .A(S), .Z(O[175]) );
  ANDN U174 ( .B(A[174]), .A(S), .Z(O[174]) );
  ANDN U175 ( .B(A[173]), .A(S), .Z(O[173]) );
  ANDN U176 ( .B(A[172]), .A(S), .Z(O[172]) );
  ANDN U177 ( .B(A[171]), .A(S), .Z(O[171]) );
  ANDN U178 ( .B(A[170]), .A(S), .Z(O[170]) );
  ANDN U179 ( .B(A[16]), .A(S), .Z(O[16]) );
  ANDN U180 ( .B(A[169]), .A(S), .Z(O[169]) );
  ANDN U181 ( .B(A[168]), .A(S), .Z(O[168]) );
  ANDN U182 ( .B(A[167]), .A(S), .Z(O[167]) );
  ANDN U183 ( .B(A[166]), .A(S), .Z(O[166]) );
  ANDN U184 ( .B(A[165]), .A(S), .Z(O[165]) );
  ANDN U185 ( .B(A[164]), .A(S), .Z(O[164]) );
  ANDN U186 ( .B(A[163]), .A(S), .Z(O[163]) );
  ANDN U187 ( .B(A[162]), .A(S), .Z(O[162]) );
  ANDN U188 ( .B(A[161]), .A(S), .Z(O[161]) );
  ANDN U189 ( .B(A[160]), .A(S), .Z(O[160]) );
  ANDN U190 ( .B(A[15]), .A(S), .Z(O[15]) );
  ANDN U191 ( .B(A[159]), .A(S), .Z(O[159]) );
  ANDN U192 ( .B(A[158]), .A(S), .Z(O[158]) );
  ANDN U193 ( .B(A[157]), .A(S), .Z(O[157]) );
  ANDN U194 ( .B(A[156]), .A(S), .Z(O[156]) );
  ANDN U195 ( .B(A[155]), .A(S), .Z(O[155]) );
  ANDN U196 ( .B(A[154]), .A(S), .Z(O[154]) );
  ANDN U197 ( .B(A[153]), .A(S), .Z(O[153]) );
  ANDN U198 ( .B(A[152]), .A(S), .Z(O[152]) );
  ANDN U199 ( .B(A[151]), .A(S), .Z(O[151]) );
  ANDN U200 ( .B(A[150]), .A(S), .Z(O[150]) );
  ANDN U201 ( .B(A[14]), .A(S), .Z(O[14]) );
  ANDN U202 ( .B(A[149]), .A(S), .Z(O[149]) );
  ANDN U203 ( .B(A[148]), .A(S), .Z(O[148]) );
  ANDN U204 ( .B(A[147]), .A(S), .Z(O[147]) );
  ANDN U205 ( .B(A[146]), .A(S), .Z(O[146]) );
  ANDN U206 ( .B(A[145]), .A(S), .Z(O[145]) );
  ANDN U207 ( .B(A[144]), .A(S), .Z(O[144]) );
  ANDN U208 ( .B(A[143]), .A(S), .Z(O[143]) );
  ANDN U209 ( .B(A[142]), .A(S), .Z(O[142]) );
  ANDN U210 ( .B(A[141]), .A(S), .Z(O[141]) );
  ANDN U211 ( .B(A[140]), .A(S), .Z(O[140]) );
  ANDN U212 ( .B(A[13]), .A(S), .Z(O[13]) );
  ANDN U213 ( .B(A[139]), .A(S), .Z(O[139]) );
  ANDN U214 ( .B(A[138]), .A(S), .Z(O[138]) );
  ANDN U215 ( .B(A[137]), .A(S), .Z(O[137]) );
  ANDN U216 ( .B(A[136]), .A(S), .Z(O[136]) );
  ANDN U217 ( .B(A[135]), .A(S), .Z(O[135]) );
  ANDN U218 ( .B(A[134]), .A(S), .Z(O[134]) );
  ANDN U219 ( .B(A[133]), .A(S), .Z(O[133]) );
  ANDN U220 ( .B(A[132]), .A(S), .Z(O[132]) );
  ANDN U221 ( .B(A[131]), .A(S), .Z(O[131]) );
  ANDN U222 ( .B(A[130]), .A(S), .Z(O[130]) );
  ANDN U223 ( .B(A[12]), .A(S), .Z(O[12]) );
  ANDN U224 ( .B(A[129]), .A(S), .Z(O[129]) );
  ANDN U225 ( .B(A[128]), .A(S), .Z(O[128]) );
  ANDN U226 ( .B(A[127]), .A(S), .Z(O[127]) );
  ANDN U227 ( .B(A[126]), .A(S), .Z(O[126]) );
  ANDN U228 ( .B(A[125]), .A(S), .Z(O[125]) );
  ANDN U229 ( .B(A[124]), .A(S), .Z(O[124]) );
  ANDN U230 ( .B(A[123]), .A(S), .Z(O[123]) );
  ANDN U231 ( .B(A[122]), .A(S), .Z(O[122]) );
  ANDN U232 ( .B(A[121]), .A(S), .Z(O[121]) );
  ANDN U233 ( .B(A[120]), .A(S), .Z(O[120]) );
  ANDN U234 ( .B(A[11]), .A(S), .Z(O[11]) );
  ANDN U235 ( .B(A[119]), .A(S), .Z(O[119]) );
  ANDN U236 ( .B(A[118]), .A(S), .Z(O[118]) );
  ANDN U237 ( .B(A[117]), .A(S), .Z(O[117]) );
  ANDN U238 ( .B(A[116]), .A(S), .Z(O[116]) );
  ANDN U239 ( .B(A[115]), .A(S), .Z(O[115]) );
  ANDN U240 ( .B(A[114]), .A(S), .Z(O[114]) );
  ANDN U241 ( .B(A[113]), .A(S), .Z(O[113]) );
  ANDN U242 ( .B(A[112]), .A(S), .Z(O[112]) );
  ANDN U243 ( .B(A[111]), .A(S), .Z(O[111]) );
  ANDN U244 ( .B(A[110]), .A(S), .Z(O[110]) );
  ANDN U245 ( .B(A[10]), .A(S), .Z(O[10]) );
  ANDN U246 ( .B(A[109]), .A(S), .Z(O[109]) );
  ANDN U247 ( .B(A[108]), .A(S), .Z(O[108]) );
  ANDN U248 ( .B(A[107]), .A(S), .Z(O[107]) );
  ANDN U249 ( .B(A[106]), .A(S), .Z(O[106]) );
  ANDN U250 ( .B(A[105]), .A(S), .Z(O[105]) );
  ANDN U251 ( .B(A[104]), .A(S), .Z(O[104]) );
  ANDN U252 ( .B(A[103]), .A(S), .Z(O[103]) );
  ANDN U253 ( .B(A[102]), .A(S), .Z(O[102]) );
  ANDN U254 ( .B(A[101]), .A(S), .Z(O[101]) );
  ANDN U255 ( .B(A[100]), .A(S), .Z(O[100]) );
  ANDN U256 ( .B(A[0]), .A(S), .Z(O[0]) );
endmodule


module FA_2838 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  AND U1 ( .A(CI), .B(B), .Z(CO) );
endmodule


module FA_2839 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  AND U1 ( .A(CI), .B(B), .Z(CO) );
endmodule


module FA_2840 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2841 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2842 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2843 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2844 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2845 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2846 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2847 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2848 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2849 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2850 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2851 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2852 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2853 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2854 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2855 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2856 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2857 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2858 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2859 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2860 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2861 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2862 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2863 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2864 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2865 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2866 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2867 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2868 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2869 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2870 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2871 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2872 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2873 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2874 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2875 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2876 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2877 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2878 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2879 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2880 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2881 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2882 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2883 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2884 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2885 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2886 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2887 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2888 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2889 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2890 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2891 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2892 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2893 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2894 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2895 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2896 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2897 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2898 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2899 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2900 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2901 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2902 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2903 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2904 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2905 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2906 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2907 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2908 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2909 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2910 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2911 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2912 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2913 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2914 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2915 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2916 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2917 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2918 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2919 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2920 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2921 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2922 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2923 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2924 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2925 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2926 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2927 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2928 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2929 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2930 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2931 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2932 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2933 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2934 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2935 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2936 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2937 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2938 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2939 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2940 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2941 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2942 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2943 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2944 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2945 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2946 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2947 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2948 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2949 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2950 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2951 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2952 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2953 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2954 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2955 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2956 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2957 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2958 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2959 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2960 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2961 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2962 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2963 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2964 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2965 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2966 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2967 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2968 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2969 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2970 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2971 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2972 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2973 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2974 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2975 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2976 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2977 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2978 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2979 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2980 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2981 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2982 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2983 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2984 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2985 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2986 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2987 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2988 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2989 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2990 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2991 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2992 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2993 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2994 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2995 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2996 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2997 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2998 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2999 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3000 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3001 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3002 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3003 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3004 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3005 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3006 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3007 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3008 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3009 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3010 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3011 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3012 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3013 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3014 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3015 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3016 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3017 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3018 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3019 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3020 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3021 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3022 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3023 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3024 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3025 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3026 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3027 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3028 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3029 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3030 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3031 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3032 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3033 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3034 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3035 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3036 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3037 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3038 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3039 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3040 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3041 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3042 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3043 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3044 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3045 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3046 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3047 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3048 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3049 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3050 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3051 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3052 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3053 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3054 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3055 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3056 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3057 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3058 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3059 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3060 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3061 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3062 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3063 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3064 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3065 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3066 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3067 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3068 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3069 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3070 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3071 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3072 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3073 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3074 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3075 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3076 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3077 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3078 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3079 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3080 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3081 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3082 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3083 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3084 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3085 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3086 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3087 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3088 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3089 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3090 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3091 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3092 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3093 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3094 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_3095 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  OR U1 ( .A(B), .B(A), .Z(CO) );
endmodule


module COMP_N258_5 ( A, B, O );
  input [257:0] A;
  input [257:0] B;
  output O;
  wire   n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517;
  wire   [257:1] C;

  FA_3095 \FAINST[0].FA_  ( .A(A[0]), .B(n260), .CI(1'b1), .CO(C[1]) );
  FA_3094 \FAINST[1].FA_  ( .A(A[1]), .B(n261), .CI(C[1]), .CO(C[2]) );
  FA_3093 \FAINST[2].FA_  ( .A(A[2]), .B(n262), .CI(C[2]), .CO(C[3]) );
  FA_3092 \FAINST[3].FA_  ( .A(A[3]), .B(n263), .CI(C[3]), .CO(C[4]) );
  FA_3091 \FAINST[4].FA_  ( .A(A[4]), .B(n264), .CI(C[4]), .CO(C[5]) );
  FA_3090 \FAINST[5].FA_  ( .A(A[5]), .B(n265), .CI(C[5]), .CO(C[6]) );
  FA_3089 \FAINST[6].FA_  ( .A(A[6]), .B(n266), .CI(C[6]), .CO(C[7]) );
  FA_3088 \FAINST[7].FA_  ( .A(A[7]), .B(n267), .CI(C[7]), .CO(C[8]) );
  FA_3087 \FAINST[8].FA_  ( .A(A[8]), .B(n268), .CI(C[8]), .CO(C[9]) );
  FA_3086 \FAINST[9].FA_  ( .A(A[9]), .B(n269), .CI(C[9]), .CO(C[10]) );
  FA_3085 \FAINST[10].FA_  ( .A(A[10]), .B(n270), .CI(C[10]), .CO(C[11]) );
  FA_3084 \FAINST[11].FA_  ( .A(A[11]), .B(n271), .CI(C[11]), .CO(C[12]) );
  FA_3083 \FAINST[12].FA_  ( .A(A[12]), .B(n272), .CI(C[12]), .CO(C[13]) );
  FA_3082 \FAINST[13].FA_  ( .A(A[13]), .B(n273), .CI(C[13]), .CO(C[14]) );
  FA_3081 \FAINST[14].FA_  ( .A(A[14]), .B(n274), .CI(C[14]), .CO(C[15]) );
  FA_3080 \FAINST[15].FA_  ( .A(A[15]), .B(n275), .CI(C[15]), .CO(C[16]) );
  FA_3079 \FAINST[16].FA_  ( .A(A[16]), .B(n276), .CI(C[16]), .CO(C[17]) );
  FA_3078 \FAINST[17].FA_  ( .A(A[17]), .B(n277), .CI(C[17]), .CO(C[18]) );
  FA_3077 \FAINST[18].FA_  ( .A(A[18]), .B(n278), .CI(C[18]), .CO(C[19]) );
  FA_3076 \FAINST[19].FA_  ( .A(A[19]), .B(n279), .CI(C[19]), .CO(C[20]) );
  FA_3075 \FAINST[20].FA_  ( .A(A[20]), .B(n280), .CI(C[20]), .CO(C[21]) );
  FA_3074 \FAINST[21].FA_  ( .A(A[21]), .B(n281), .CI(C[21]), .CO(C[22]) );
  FA_3073 \FAINST[22].FA_  ( .A(A[22]), .B(n282), .CI(C[22]), .CO(C[23]) );
  FA_3072 \FAINST[23].FA_  ( .A(A[23]), .B(n283), .CI(C[23]), .CO(C[24]) );
  FA_3071 \FAINST[24].FA_  ( .A(A[24]), .B(n284), .CI(C[24]), .CO(C[25]) );
  FA_3070 \FAINST[25].FA_  ( .A(A[25]), .B(n285), .CI(C[25]), .CO(C[26]) );
  FA_3069 \FAINST[26].FA_  ( .A(A[26]), .B(n286), .CI(C[26]), .CO(C[27]) );
  FA_3068 \FAINST[27].FA_  ( .A(A[27]), .B(n287), .CI(C[27]), .CO(C[28]) );
  FA_3067 \FAINST[28].FA_  ( .A(A[28]), .B(n288), .CI(C[28]), .CO(C[29]) );
  FA_3066 \FAINST[29].FA_  ( .A(A[29]), .B(n289), .CI(C[29]), .CO(C[30]) );
  FA_3065 \FAINST[30].FA_  ( .A(A[30]), .B(n290), .CI(C[30]), .CO(C[31]) );
  FA_3064 \FAINST[31].FA_  ( .A(A[31]), .B(n291), .CI(C[31]), .CO(C[32]) );
  FA_3063 \FAINST[32].FA_  ( .A(A[32]), .B(n292), .CI(C[32]), .CO(C[33]) );
  FA_3062 \FAINST[33].FA_  ( .A(A[33]), .B(n293), .CI(C[33]), .CO(C[34]) );
  FA_3061 \FAINST[34].FA_  ( .A(A[34]), .B(n294), .CI(C[34]), .CO(C[35]) );
  FA_3060 \FAINST[35].FA_  ( .A(A[35]), .B(n295), .CI(C[35]), .CO(C[36]) );
  FA_3059 \FAINST[36].FA_  ( .A(A[36]), .B(n296), .CI(C[36]), .CO(C[37]) );
  FA_3058 \FAINST[37].FA_  ( .A(A[37]), .B(n297), .CI(C[37]), .CO(C[38]) );
  FA_3057 \FAINST[38].FA_  ( .A(A[38]), .B(n298), .CI(C[38]), .CO(C[39]) );
  FA_3056 \FAINST[39].FA_  ( .A(A[39]), .B(n299), .CI(C[39]), .CO(C[40]) );
  FA_3055 \FAINST[40].FA_  ( .A(A[40]), .B(n300), .CI(C[40]), .CO(C[41]) );
  FA_3054 \FAINST[41].FA_  ( .A(A[41]), .B(n301), .CI(C[41]), .CO(C[42]) );
  FA_3053 \FAINST[42].FA_  ( .A(A[42]), .B(n302), .CI(C[42]), .CO(C[43]) );
  FA_3052 \FAINST[43].FA_  ( .A(A[43]), .B(n303), .CI(C[43]), .CO(C[44]) );
  FA_3051 \FAINST[44].FA_  ( .A(A[44]), .B(n304), .CI(C[44]), .CO(C[45]) );
  FA_3050 \FAINST[45].FA_  ( .A(A[45]), .B(n305), .CI(C[45]), .CO(C[46]) );
  FA_3049 \FAINST[46].FA_  ( .A(A[46]), .B(n306), .CI(C[46]), .CO(C[47]) );
  FA_3048 \FAINST[47].FA_  ( .A(A[47]), .B(n307), .CI(C[47]), .CO(C[48]) );
  FA_3047 \FAINST[48].FA_  ( .A(A[48]), .B(n308), .CI(C[48]), .CO(C[49]) );
  FA_3046 \FAINST[49].FA_  ( .A(A[49]), .B(n309), .CI(C[49]), .CO(C[50]) );
  FA_3045 \FAINST[50].FA_  ( .A(A[50]), .B(n310), .CI(C[50]), .CO(C[51]) );
  FA_3044 \FAINST[51].FA_  ( .A(A[51]), .B(n311), .CI(C[51]), .CO(C[52]) );
  FA_3043 \FAINST[52].FA_  ( .A(A[52]), .B(n312), .CI(C[52]), .CO(C[53]) );
  FA_3042 \FAINST[53].FA_  ( .A(A[53]), .B(n313), .CI(C[53]), .CO(C[54]) );
  FA_3041 \FAINST[54].FA_  ( .A(A[54]), .B(n314), .CI(C[54]), .CO(C[55]) );
  FA_3040 \FAINST[55].FA_  ( .A(A[55]), .B(n315), .CI(C[55]), .CO(C[56]) );
  FA_3039 \FAINST[56].FA_  ( .A(A[56]), .B(n316), .CI(C[56]), .CO(C[57]) );
  FA_3038 \FAINST[57].FA_  ( .A(A[57]), .B(n317), .CI(C[57]), .CO(C[58]) );
  FA_3037 \FAINST[58].FA_  ( .A(A[58]), .B(n318), .CI(C[58]), .CO(C[59]) );
  FA_3036 \FAINST[59].FA_  ( .A(A[59]), .B(n319), .CI(C[59]), .CO(C[60]) );
  FA_3035 \FAINST[60].FA_  ( .A(A[60]), .B(n320), .CI(C[60]), .CO(C[61]) );
  FA_3034 \FAINST[61].FA_  ( .A(A[61]), .B(n321), .CI(C[61]), .CO(C[62]) );
  FA_3033 \FAINST[62].FA_  ( .A(A[62]), .B(n322), .CI(C[62]), .CO(C[63]) );
  FA_3032 \FAINST[63].FA_  ( .A(A[63]), .B(n323), .CI(C[63]), .CO(C[64]) );
  FA_3031 \FAINST[64].FA_  ( .A(A[64]), .B(n324), .CI(C[64]), .CO(C[65]) );
  FA_3030 \FAINST[65].FA_  ( .A(A[65]), .B(n325), .CI(C[65]), .CO(C[66]) );
  FA_3029 \FAINST[66].FA_  ( .A(A[66]), .B(n326), .CI(C[66]), .CO(C[67]) );
  FA_3028 \FAINST[67].FA_  ( .A(A[67]), .B(n327), .CI(C[67]), .CO(C[68]) );
  FA_3027 \FAINST[68].FA_  ( .A(A[68]), .B(n328), .CI(C[68]), .CO(C[69]) );
  FA_3026 \FAINST[69].FA_  ( .A(A[69]), .B(n329), .CI(C[69]), .CO(C[70]) );
  FA_3025 \FAINST[70].FA_  ( .A(A[70]), .B(n330), .CI(C[70]), .CO(C[71]) );
  FA_3024 \FAINST[71].FA_  ( .A(A[71]), .B(n331), .CI(C[71]), .CO(C[72]) );
  FA_3023 \FAINST[72].FA_  ( .A(A[72]), .B(n332), .CI(C[72]), .CO(C[73]) );
  FA_3022 \FAINST[73].FA_  ( .A(A[73]), .B(n333), .CI(C[73]), .CO(C[74]) );
  FA_3021 \FAINST[74].FA_  ( .A(A[74]), .B(n334), .CI(C[74]), .CO(C[75]) );
  FA_3020 \FAINST[75].FA_  ( .A(A[75]), .B(n335), .CI(C[75]), .CO(C[76]) );
  FA_3019 \FAINST[76].FA_  ( .A(A[76]), .B(n336), .CI(C[76]), .CO(C[77]) );
  FA_3018 \FAINST[77].FA_  ( .A(A[77]), .B(n337), .CI(C[77]), .CO(C[78]) );
  FA_3017 \FAINST[78].FA_  ( .A(A[78]), .B(n338), .CI(C[78]), .CO(C[79]) );
  FA_3016 \FAINST[79].FA_  ( .A(A[79]), .B(n339), .CI(C[79]), .CO(C[80]) );
  FA_3015 \FAINST[80].FA_  ( .A(A[80]), .B(n340), .CI(C[80]), .CO(C[81]) );
  FA_3014 \FAINST[81].FA_  ( .A(A[81]), .B(n341), .CI(C[81]), .CO(C[82]) );
  FA_3013 \FAINST[82].FA_  ( .A(A[82]), .B(n342), .CI(C[82]), .CO(C[83]) );
  FA_3012 \FAINST[83].FA_  ( .A(A[83]), .B(n343), .CI(C[83]), .CO(C[84]) );
  FA_3011 \FAINST[84].FA_  ( .A(A[84]), .B(n344), .CI(C[84]), .CO(C[85]) );
  FA_3010 \FAINST[85].FA_  ( .A(A[85]), .B(n345), .CI(C[85]), .CO(C[86]) );
  FA_3009 \FAINST[86].FA_  ( .A(A[86]), .B(n346), .CI(C[86]), .CO(C[87]) );
  FA_3008 \FAINST[87].FA_  ( .A(A[87]), .B(n347), .CI(C[87]), .CO(C[88]) );
  FA_3007 \FAINST[88].FA_  ( .A(A[88]), .B(n348), .CI(C[88]), .CO(C[89]) );
  FA_3006 \FAINST[89].FA_  ( .A(A[89]), .B(n349), .CI(C[89]), .CO(C[90]) );
  FA_3005 \FAINST[90].FA_  ( .A(A[90]), .B(n350), .CI(C[90]), .CO(C[91]) );
  FA_3004 \FAINST[91].FA_  ( .A(A[91]), .B(n351), .CI(C[91]), .CO(C[92]) );
  FA_3003 \FAINST[92].FA_  ( .A(A[92]), .B(n352), .CI(C[92]), .CO(C[93]) );
  FA_3002 \FAINST[93].FA_  ( .A(A[93]), .B(n353), .CI(C[93]), .CO(C[94]) );
  FA_3001 \FAINST[94].FA_  ( .A(A[94]), .B(n354), .CI(C[94]), .CO(C[95]) );
  FA_3000 \FAINST[95].FA_  ( .A(A[95]), .B(n355), .CI(C[95]), .CO(C[96]) );
  FA_2999 \FAINST[96].FA_  ( .A(A[96]), .B(n356), .CI(C[96]), .CO(C[97]) );
  FA_2998 \FAINST[97].FA_  ( .A(A[97]), .B(n357), .CI(C[97]), .CO(C[98]) );
  FA_2997 \FAINST[98].FA_  ( .A(A[98]), .B(n358), .CI(C[98]), .CO(C[99]) );
  FA_2996 \FAINST[99].FA_  ( .A(A[99]), .B(n359), .CI(C[99]), .CO(C[100]) );
  FA_2995 \FAINST[100].FA_  ( .A(A[100]), .B(n360), .CI(C[100]), .CO(C[101])
         );
  FA_2994 \FAINST[101].FA_  ( .A(A[101]), .B(n361), .CI(C[101]), .CO(C[102])
         );
  FA_2993 \FAINST[102].FA_  ( .A(A[102]), .B(n362), .CI(C[102]), .CO(C[103])
         );
  FA_2992 \FAINST[103].FA_  ( .A(A[103]), .B(n363), .CI(C[103]), .CO(C[104])
         );
  FA_2991 \FAINST[104].FA_  ( .A(A[104]), .B(n364), .CI(C[104]), .CO(C[105])
         );
  FA_2990 \FAINST[105].FA_  ( .A(A[105]), .B(n365), .CI(C[105]), .CO(C[106])
         );
  FA_2989 \FAINST[106].FA_  ( .A(A[106]), .B(n366), .CI(C[106]), .CO(C[107])
         );
  FA_2988 \FAINST[107].FA_  ( .A(A[107]), .B(n367), .CI(C[107]), .CO(C[108])
         );
  FA_2987 \FAINST[108].FA_  ( .A(A[108]), .B(n368), .CI(C[108]), .CO(C[109])
         );
  FA_2986 \FAINST[109].FA_  ( .A(A[109]), .B(n369), .CI(C[109]), .CO(C[110])
         );
  FA_2985 \FAINST[110].FA_  ( .A(A[110]), .B(n370), .CI(C[110]), .CO(C[111])
         );
  FA_2984 \FAINST[111].FA_  ( .A(A[111]), .B(n371), .CI(C[111]), .CO(C[112])
         );
  FA_2983 \FAINST[112].FA_  ( .A(A[112]), .B(n372), .CI(C[112]), .CO(C[113])
         );
  FA_2982 \FAINST[113].FA_  ( .A(A[113]), .B(n373), .CI(C[113]), .CO(C[114])
         );
  FA_2981 \FAINST[114].FA_  ( .A(A[114]), .B(n374), .CI(C[114]), .CO(C[115])
         );
  FA_2980 \FAINST[115].FA_  ( .A(A[115]), .B(n375), .CI(C[115]), .CO(C[116])
         );
  FA_2979 \FAINST[116].FA_  ( .A(A[116]), .B(n376), .CI(C[116]), .CO(C[117])
         );
  FA_2978 \FAINST[117].FA_  ( .A(A[117]), .B(n377), .CI(C[117]), .CO(C[118])
         );
  FA_2977 \FAINST[118].FA_  ( .A(A[118]), .B(n378), .CI(C[118]), .CO(C[119])
         );
  FA_2976 \FAINST[119].FA_  ( .A(A[119]), .B(n379), .CI(C[119]), .CO(C[120])
         );
  FA_2975 \FAINST[120].FA_  ( .A(A[120]), .B(n380), .CI(C[120]), .CO(C[121])
         );
  FA_2974 \FAINST[121].FA_  ( .A(A[121]), .B(n381), .CI(C[121]), .CO(C[122])
         );
  FA_2973 \FAINST[122].FA_  ( .A(A[122]), .B(n382), .CI(C[122]), .CO(C[123])
         );
  FA_2972 \FAINST[123].FA_  ( .A(A[123]), .B(n383), .CI(C[123]), .CO(C[124])
         );
  FA_2971 \FAINST[124].FA_  ( .A(A[124]), .B(n384), .CI(C[124]), .CO(C[125])
         );
  FA_2970 \FAINST[125].FA_  ( .A(A[125]), .B(n385), .CI(C[125]), .CO(C[126])
         );
  FA_2969 \FAINST[126].FA_  ( .A(A[126]), .B(n386), .CI(C[126]), .CO(C[127])
         );
  FA_2968 \FAINST[127].FA_  ( .A(A[127]), .B(n387), .CI(C[127]), .CO(C[128])
         );
  FA_2967 \FAINST[128].FA_  ( .A(A[128]), .B(n388), .CI(C[128]), .CO(C[129])
         );
  FA_2966 \FAINST[129].FA_  ( .A(A[129]), .B(n389), .CI(C[129]), .CO(C[130])
         );
  FA_2965 \FAINST[130].FA_  ( .A(A[130]), .B(n390), .CI(C[130]), .CO(C[131])
         );
  FA_2964 \FAINST[131].FA_  ( .A(A[131]), .B(n391), .CI(C[131]), .CO(C[132])
         );
  FA_2963 \FAINST[132].FA_  ( .A(A[132]), .B(n392), .CI(C[132]), .CO(C[133])
         );
  FA_2962 \FAINST[133].FA_  ( .A(A[133]), .B(n393), .CI(C[133]), .CO(C[134])
         );
  FA_2961 \FAINST[134].FA_  ( .A(A[134]), .B(n394), .CI(C[134]), .CO(C[135])
         );
  FA_2960 \FAINST[135].FA_  ( .A(A[135]), .B(n395), .CI(C[135]), .CO(C[136])
         );
  FA_2959 \FAINST[136].FA_  ( .A(A[136]), .B(n396), .CI(C[136]), .CO(C[137])
         );
  FA_2958 \FAINST[137].FA_  ( .A(A[137]), .B(n397), .CI(C[137]), .CO(C[138])
         );
  FA_2957 \FAINST[138].FA_  ( .A(A[138]), .B(n398), .CI(C[138]), .CO(C[139])
         );
  FA_2956 \FAINST[139].FA_  ( .A(A[139]), .B(n399), .CI(C[139]), .CO(C[140])
         );
  FA_2955 \FAINST[140].FA_  ( .A(A[140]), .B(n400), .CI(C[140]), .CO(C[141])
         );
  FA_2954 \FAINST[141].FA_  ( .A(A[141]), .B(n401), .CI(C[141]), .CO(C[142])
         );
  FA_2953 \FAINST[142].FA_  ( .A(A[142]), .B(n402), .CI(C[142]), .CO(C[143])
         );
  FA_2952 \FAINST[143].FA_  ( .A(A[143]), .B(n403), .CI(C[143]), .CO(C[144])
         );
  FA_2951 \FAINST[144].FA_  ( .A(A[144]), .B(n404), .CI(C[144]), .CO(C[145])
         );
  FA_2950 \FAINST[145].FA_  ( .A(A[145]), .B(n405), .CI(C[145]), .CO(C[146])
         );
  FA_2949 \FAINST[146].FA_  ( .A(A[146]), .B(n406), .CI(C[146]), .CO(C[147])
         );
  FA_2948 \FAINST[147].FA_  ( .A(A[147]), .B(n407), .CI(C[147]), .CO(C[148])
         );
  FA_2947 \FAINST[148].FA_  ( .A(A[148]), .B(n408), .CI(C[148]), .CO(C[149])
         );
  FA_2946 \FAINST[149].FA_  ( .A(A[149]), .B(n409), .CI(C[149]), .CO(C[150])
         );
  FA_2945 \FAINST[150].FA_  ( .A(A[150]), .B(n410), .CI(C[150]), .CO(C[151])
         );
  FA_2944 \FAINST[151].FA_  ( .A(A[151]), .B(n411), .CI(C[151]), .CO(C[152])
         );
  FA_2943 \FAINST[152].FA_  ( .A(A[152]), .B(n412), .CI(C[152]), .CO(C[153])
         );
  FA_2942 \FAINST[153].FA_  ( .A(A[153]), .B(n413), .CI(C[153]), .CO(C[154])
         );
  FA_2941 \FAINST[154].FA_  ( .A(A[154]), .B(n414), .CI(C[154]), .CO(C[155])
         );
  FA_2940 \FAINST[155].FA_  ( .A(A[155]), .B(n415), .CI(C[155]), .CO(C[156])
         );
  FA_2939 \FAINST[156].FA_  ( .A(A[156]), .B(n416), .CI(C[156]), .CO(C[157])
         );
  FA_2938 \FAINST[157].FA_  ( .A(A[157]), .B(n417), .CI(C[157]), .CO(C[158])
         );
  FA_2937 \FAINST[158].FA_  ( .A(A[158]), .B(n418), .CI(C[158]), .CO(C[159])
         );
  FA_2936 \FAINST[159].FA_  ( .A(A[159]), .B(n419), .CI(C[159]), .CO(C[160])
         );
  FA_2935 \FAINST[160].FA_  ( .A(A[160]), .B(n420), .CI(C[160]), .CO(C[161])
         );
  FA_2934 \FAINST[161].FA_  ( .A(A[161]), .B(n421), .CI(C[161]), .CO(C[162])
         );
  FA_2933 \FAINST[162].FA_  ( .A(A[162]), .B(n422), .CI(C[162]), .CO(C[163])
         );
  FA_2932 \FAINST[163].FA_  ( .A(A[163]), .B(n423), .CI(C[163]), .CO(C[164])
         );
  FA_2931 \FAINST[164].FA_  ( .A(A[164]), .B(n424), .CI(C[164]), .CO(C[165])
         );
  FA_2930 \FAINST[165].FA_  ( .A(A[165]), .B(n425), .CI(C[165]), .CO(C[166])
         );
  FA_2929 \FAINST[166].FA_  ( .A(A[166]), .B(n426), .CI(C[166]), .CO(C[167])
         );
  FA_2928 \FAINST[167].FA_  ( .A(A[167]), .B(n427), .CI(C[167]), .CO(C[168])
         );
  FA_2927 \FAINST[168].FA_  ( .A(A[168]), .B(n428), .CI(C[168]), .CO(C[169])
         );
  FA_2926 \FAINST[169].FA_  ( .A(A[169]), .B(n429), .CI(C[169]), .CO(C[170])
         );
  FA_2925 \FAINST[170].FA_  ( .A(A[170]), .B(n430), .CI(C[170]), .CO(C[171])
         );
  FA_2924 \FAINST[171].FA_  ( .A(A[171]), .B(n431), .CI(C[171]), .CO(C[172])
         );
  FA_2923 \FAINST[172].FA_  ( .A(A[172]), .B(n432), .CI(C[172]), .CO(C[173])
         );
  FA_2922 \FAINST[173].FA_  ( .A(A[173]), .B(n433), .CI(C[173]), .CO(C[174])
         );
  FA_2921 \FAINST[174].FA_  ( .A(A[174]), .B(n434), .CI(C[174]), .CO(C[175])
         );
  FA_2920 \FAINST[175].FA_  ( .A(A[175]), .B(n435), .CI(C[175]), .CO(C[176])
         );
  FA_2919 \FAINST[176].FA_  ( .A(A[176]), .B(n436), .CI(C[176]), .CO(C[177])
         );
  FA_2918 \FAINST[177].FA_  ( .A(A[177]), .B(n437), .CI(C[177]), .CO(C[178])
         );
  FA_2917 \FAINST[178].FA_  ( .A(A[178]), .B(n438), .CI(C[178]), .CO(C[179])
         );
  FA_2916 \FAINST[179].FA_  ( .A(A[179]), .B(n439), .CI(C[179]), .CO(C[180])
         );
  FA_2915 \FAINST[180].FA_  ( .A(A[180]), .B(n440), .CI(C[180]), .CO(C[181])
         );
  FA_2914 \FAINST[181].FA_  ( .A(A[181]), .B(n441), .CI(C[181]), .CO(C[182])
         );
  FA_2913 \FAINST[182].FA_  ( .A(A[182]), .B(n442), .CI(C[182]), .CO(C[183])
         );
  FA_2912 \FAINST[183].FA_  ( .A(A[183]), .B(n443), .CI(C[183]), .CO(C[184])
         );
  FA_2911 \FAINST[184].FA_  ( .A(A[184]), .B(n444), .CI(C[184]), .CO(C[185])
         );
  FA_2910 \FAINST[185].FA_  ( .A(A[185]), .B(n445), .CI(C[185]), .CO(C[186])
         );
  FA_2909 \FAINST[186].FA_  ( .A(A[186]), .B(n446), .CI(C[186]), .CO(C[187])
         );
  FA_2908 \FAINST[187].FA_  ( .A(A[187]), .B(n447), .CI(C[187]), .CO(C[188])
         );
  FA_2907 \FAINST[188].FA_  ( .A(A[188]), .B(n448), .CI(C[188]), .CO(C[189])
         );
  FA_2906 \FAINST[189].FA_  ( .A(A[189]), .B(n449), .CI(C[189]), .CO(C[190])
         );
  FA_2905 \FAINST[190].FA_  ( .A(A[190]), .B(n450), .CI(C[190]), .CO(C[191])
         );
  FA_2904 \FAINST[191].FA_  ( .A(A[191]), .B(n451), .CI(C[191]), .CO(C[192])
         );
  FA_2903 \FAINST[192].FA_  ( .A(A[192]), .B(n452), .CI(C[192]), .CO(C[193])
         );
  FA_2902 \FAINST[193].FA_  ( .A(A[193]), .B(n453), .CI(C[193]), .CO(C[194])
         );
  FA_2901 \FAINST[194].FA_  ( .A(A[194]), .B(n454), .CI(C[194]), .CO(C[195])
         );
  FA_2900 \FAINST[195].FA_  ( .A(A[195]), .B(n455), .CI(C[195]), .CO(C[196])
         );
  FA_2899 \FAINST[196].FA_  ( .A(A[196]), .B(n456), .CI(C[196]), .CO(C[197])
         );
  FA_2898 \FAINST[197].FA_  ( .A(A[197]), .B(n457), .CI(C[197]), .CO(C[198])
         );
  FA_2897 \FAINST[198].FA_  ( .A(A[198]), .B(n458), .CI(C[198]), .CO(C[199])
         );
  FA_2896 \FAINST[199].FA_  ( .A(A[199]), .B(n459), .CI(C[199]), .CO(C[200])
         );
  FA_2895 \FAINST[200].FA_  ( .A(A[200]), .B(n460), .CI(C[200]), .CO(C[201])
         );
  FA_2894 \FAINST[201].FA_  ( .A(A[201]), .B(n461), .CI(C[201]), .CO(C[202])
         );
  FA_2893 \FAINST[202].FA_  ( .A(A[202]), .B(n462), .CI(C[202]), .CO(C[203])
         );
  FA_2892 \FAINST[203].FA_  ( .A(A[203]), .B(n463), .CI(C[203]), .CO(C[204])
         );
  FA_2891 \FAINST[204].FA_  ( .A(A[204]), .B(n464), .CI(C[204]), .CO(C[205])
         );
  FA_2890 \FAINST[205].FA_  ( .A(A[205]), .B(n465), .CI(C[205]), .CO(C[206])
         );
  FA_2889 \FAINST[206].FA_  ( .A(A[206]), .B(n466), .CI(C[206]), .CO(C[207])
         );
  FA_2888 \FAINST[207].FA_  ( .A(A[207]), .B(n467), .CI(C[207]), .CO(C[208])
         );
  FA_2887 \FAINST[208].FA_  ( .A(A[208]), .B(n468), .CI(C[208]), .CO(C[209])
         );
  FA_2886 \FAINST[209].FA_  ( .A(A[209]), .B(n469), .CI(C[209]), .CO(C[210])
         );
  FA_2885 \FAINST[210].FA_  ( .A(A[210]), .B(n470), .CI(C[210]), .CO(C[211])
         );
  FA_2884 \FAINST[211].FA_  ( .A(A[211]), .B(n471), .CI(C[211]), .CO(C[212])
         );
  FA_2883 \FAINST[212].FA_  ( .A(A[212]), .B(n472), .CI(C[212]), .CO(C[213])
         );
  FA_2882 \FAINST[213].FA_  ( .A(A[213]), .B(n473), .CI(C[213]), .CO(C[214])
         );
  FA_2881 \FAINST[214].FA_  ( .A(A[214]), .B(n474), .CI(C[214]), .CO(C[215])
         );
  FA_2880 \FAINST[215].FA_  ( .A(A[215]), .B(n475), .CI(C[215]), .CO(C[216])
         );
  FA_2879 \FAINST[216].FA_  ( .A(A[216]), .B(n476), .CI(C[216]), .CO(C[217])
         );
  FA_2878 \FAINST[217].FA_  ( .A(A[217]), .B(n477), .CI(C[217]), .CO(C[218])
         );
  FA_2877 \FAINST[218].FA_  ( .A(A[218]), .B(n478), .CI(C[218]), .CO(C[219])
         );
  FA_2876 \FAINST[219].FA_  ( .A(A[219]), .B(n479), .CI(C[219]), .CO(C[220])
         );
  FA_2875 \FAINST[220].FA_  ( .A(A[220]), .B(n480), .CI(C[220]), .CO(C[221])
         );
  FA_2874 \FAINST[221].FA_  ( .A(A[221]), .B(n481), .CI(C[221]), .CO(C[222])
         );
  FA_2873 \FAINST[222].FA_  ( .A(A[222]), .B(n482), .CI(C[222]), .CO(C[223])
         );
  FA_2872 \FAINST[223].FA_  ( .A(A[223]), .B(n483), .CI(C[223]), .CO(C[224])
         );
  FA_2871 \FAINST[224].FA_  ( .A(A[224]), .B(n484), .CI(C[224]), .CO(C[225])
         );
  FA_2870 \FAINST[225].FA_  ( .A(A[225]), .B(n485), .CI(C[225]), .CO(C[226])
         );
  FA_2869 \FAINST[226].FA_  ( .A(A[226]), .B(n486), .CI(C[226]), .CO(C[227])
         );
  FA_2868 \FAINST[227].FA_  ( .A(A[227]), .B(n487), .CI(C[227]), .CO(C[228])
         );
  FA_2867 \FAINST[228].FA_  ( .A(A[228]), .B(n488), .CI(C[228]), .CO(C[229])
         );
  FA_2866 \FAINST[229].FA_  ( .A(A[229]), .B(n489), .CI(C[229]), .CO(C[230])
         );
  FA_2865 \FAINST[230].FA_  ( .A(A[230]), .B(n490), .CI(C[230]), .CO(C[231])
         );
  FA_2864 \FAINST[231].FA_  ( .A(A[231]), .B(n491), .CI(C[231]), .CO(C[232])
         );
  FA_2863 \FAINST[232].FA_  ( .A(A[232]), .B(n492), .CI(C[232]), .CO(C[233])
         );
  FA_2862 \FAINST[233].FA_  ( .A(A[233]), .B(n493), .CI(C[233]), .CO(C[234])
         );
  FA_2861 \FAINST[234].FA_  ( .A(A[234]), .B(n494), .CI(C[234]), .CO(C[235])
         );
  FA_2860 \FAINST[235].FA_  ( .A(A[235]), .B(n495), .CI(C[235]), .CO(C[236])
         );
  FA_2859 \FAINST[236].FA_  ( .A(A[236]), .B(n496), .CI(C[236]), .CO(C[237])
         );
  FA_2858 \FAINST[237].FA_  ( .A(A[237]), .B(n497), .CI(C[237]), .CO(C[238])
         );
  FA_2857 \FAINST[238].FA_  ( .A(A[238]), .B(n498), .CI(C[238]), .CO(C[239])
         );
  FA_2856 \FAINST[239].FA_  ( .A(A[239]), .B(n499), .CI(C[239]), .CO(C[240])
         );
  FA_2855 \FAINST[240].FA_  ( .A(A[240]), .B(n500), .CI(C[240]), .CO(C[241])
         );
  FA_2854 \FAINST[241].FA_  ( .A(A[241]), .B(n501), .CI(C[241]), .CO(C[242])
         );
  FA_2853 \FAINST[242].FA_  ( .A(A[242]), .B(n502), .CI(C[242]), .CO(C[243])
         );
  FA_2852 \FAINST[243].FA_  ( .A(A[243]), .B(n503), .CI(C[243]), .CO(C[244])
         );
  FA_2851 \FAINST[244].FA_  ( .A(A[244]), .B(n504), .CI(C[244]), .CO(C[245])
         );
  FA_2850 \FAINST[245].FA_  ( .A(A[245]), .B(n505), .CI(C[245]), .CO(C[246])
         );
  FA_2849 \FAINST[246].FA_  ( .A(A[246]), .B(n506), .CI(C[246]), .CO(C[247])
         );
  FA_2848 \FAINST[247].FA_  ( .A(A[247]), .B(n507), .CI(C[247]), .CO(C[248])
         );
  FA_2847 \FAINST[248].FA_  ( .A(A[248]), .B(n508), .CI(C[248]), .CO(C[249])
         );
  FA_2846 \FAINST[249].FA_  ( .A(A[249]), .B(n509), .CI(C[249]), .CO(C[250])
         );
  FA_2845 \FAINST[250].FA_  ( .A(A[250]), .B(n510), .CI(C[250]), .CO(C[251])
         );
  FA_2844 \FAINST[251].FA_  ( .A(A[251]), .B(n511), .CI(C[251]), .CO(C[252])
         );
  FA_2843 \FAINST[252].FA_  ( .A(A[252]), .B(n512), .CI(C[252]), .CO(C[253])
         );
  FA_2842 \FAINST[253].FA_  ( .A(A[253]), .B(n513), .CI(C[253]), .CO(C[254])
         );
  FA_2841 \FAINST[254].FA_  ( .A(A[254]), .B(n514), .CI(C[254]), .CO(C[255])
         );
  FA_2840 \FAINST[255].FA_  ( .A(A[255]), .B(n515), .CI(C[255]), .CO(C[256])
         );
  FA_2839 \FAINST[256].FA_  ( .A(1'b0), .B(n516), .CI(C[256]), .CO(C[257]) );
  FA_2838 \FAINST[257].FA_  ( .A(1'b0), .B(n517), .CI(C[257]), .CO(O) );
  IV U2 ( .A(B[159]), .Z(n419) );
  IV U3 ( .A(B[160]), .Z(n420) );
  IV U4 ( .A(B[161]), .Z(n421) );
  IV U5 ( .A(B[162]), .Z(n422) );
  IV U6 ( .A(B[163]), .Z(n423) );
  IV U7 ( .A(B[164]), .Z(n424) );
  IV U8 ( .A(B[165]), .Z(n425) );
  IV U9 ( .A(B[166]), .Z(n426) );
  IV U10 ( .A(B[167]), .Z(n427) );
  IV U11 ( .A(B[168]), .Z(n428) );
  IV U12 ( .A(B[249]), .Z(n509) );
  IV U13 ( .A(B[169]), .Z(n429) );
  IV U14 ( .A(B[170]), .Z(n430) );
  IV U15 ( .A(B[171]), .Z(n431) );
  IV U16 ( .A(B[172]), .Z(n432) );
  IV U17 ( .A(B[173]), .Z(n433) );
  IV U18 ( .A(B[174]), .Z(n434) );
  IV U19 ( .A(B[175]), .Z(n435) );
  IV U20 ( .A(B[176]), .Z(n436) );
  IV U21 ( .A(B[177]), .Z(n437) );
  IV U22 ( .A(B[178]), .Z(n438) );
  IV U23 ( .A(B[250]), .Z(n510) );
  IV U24 ( .A(B[179]), .Z(n439) );
  IV U25 ( .A(B[180]), .Z(n440) );
  IV U26 ( .A(B[181]), .Z(n441) );
  IV U27 ( .A(B[182]), .Z(n442) );
  IV U28 ( .A(B[183]), .Z(n443) );
  IV U29 ( .A(B[184]), .Z(n444) );
  IV U30 ( .A(B[185]), .Z(n445) );
  IV U31 ( .A(B[186]), .Z(n446) );
  IV U32 ( .A(B[187]), .Z(n447) );
  IV U33 ( .A(B[188]), .Z(n448) );
  IV U34 ( .A(B[251]), .Z(n511) );
  IV U35 ( .A(B[189]), .Z(n449) );
  IV U36 ( .A(B[190]), .Z(n450) );
  IV U37 ( .A(B[191]), .Z(n451) );
  IV U38 ( .A(B[192]), .Z(n452) );
  IV U39 ( .A(B[193]), .Z(n453) );
  IV U40 ( .A(B[194]), .Z(n454) );
  IV U41 ( .A(B[195]), .Z(n455) );
  IV U42 ( .A(B[196]), .Z(n456) );
  IV U43 ( .A(B[197]), .Z(n457) );
  IV U44 ( .A(B[198]), .Z(n458) );
  IV U45 ( .A(B[252]), .Z(n512) );
  IV U46 ( .A(B[199]), .Z(n459) );
  IV U47 ( .A(B[200]), .Z(n460) );
  IV U48 ( .A(B[201]), .Z(n461) );
  IV U49 ( .A(B[202]), .Z(n462) );
  IV U50 ( .A(B[203]), .Z(n463) );
  IV U51 ( .A(B[204]), .Z(n464) );
  IV U52 ( .A(B[205]), .Z(n465) );
  IV U53 ( .A(B[206]), .Z(n466) );
  IV U54 ( .A(B[207]), .Z(n467) );
  IV U55 ( .A(B[208]), .Z(n468) );
  IV U56 ( .A(B[253]), .Z(n513) );
  IV U57 ( .A(B[209]), .Z(n469) );
  IV U58 ( .A(B[210]), .Z(n470) );
  IV U59 ( .A(B[211]), .Z(n471) );
  IV U60 ( .A(B[212]), .Z(n472) );
  IV U61 ( .A(B[213]), .Z(n473) );
  IV U62 ( .A(B[214]), .Z(n474) );
  IV U63 ( .A(B[215]), .Z(n475) );
  IV U64 ( .A(B[216]), .Z(n476) );
  IV U65 ( .A(B[217]), .Z(n477) );
  IV U66 ( .A(B[218]), .Z(n478) );
  IV U67 ( .A(B[254]), .Z(n514) );
  IV U68 ( .A(B[219]), .Z(n479) );
  IV U69 ( .A(B[220]), .Z(n480) );
  IV U70 ( .A(B[221]), .Z(n481) );
  IV U71 ( .A(B[222]), .Z(n482) );
  IV U72 ( .A(B[223]), .Z(n483) );
  IV U73 ( .A(B[224]), .Z(n484) );
  IV U74 ( .A(B[225]), .Z(n485) );
  IV U75 ( .A(B[226]), .Z(n486) );
  IV U76 ( .A(B[227]), .Z(n487) );
  IV U77 ( .A(B[228]), .Z(n488) );
  IV U78 ( .A(B[255]), .Z(n515) );
  IV U79 ( .A(B[229]), .Z(n489) );
  IV U80 ( .A(B[230]), .Z(n490) );
  IV U81 ( .A(B[231]), .Z(n491) );
  IV U82 ( .A(B[232]), .Z(n492) );
  IV U83 ( .A(B[0]), .Z(n260) );
  IV U84 ( .A(B[1]), .Z(n261) );
  IV U85 ( .A(B[2]), .Z(n262) );
  IV U86 ( .A(B[3]), .Z(n263) );
  IV U87 ( .A(B[4]), .Z(n264) );
  IV U88 ( .A(B[5]), .Z(n265) );
  IV U89 ( .A(B[6]), .Z(n266) );
  IV U90 ( .A(B[7]), .Z(n267) );
  IV U91 ( .A(B[8]), .Z(n268) );
  IV U92 ( .A(B[233]), .Z(n493) );
  IV U93 ( .A(B[9]), .Z(n269) );
  IV U94 ( .A(B[10]), .Z(n270) );
  IV U95 ( .A(B[11]), .Z(n271) );
  IV U96 ( .A(B[12]), .Z(n272) );
  IV U97 ( .A(B[13]), .Z(n273) );
  IV U98 ( .A(B[14]), .Z(n274) );
  IV U99 ( .A(B[15]), .Z(n275) );
  IV U100 ( .A(B[16]), .Z(n276) );
  IV U101 ( .A(B[17]), .Z(n277) );
  IV U102 ( .A(B[18]), .Z(n278) );
  IV U103 ( .A(B[234]), .Z(n494) );
  IV U104 ( .A(B[19]), .Z(n279) );
  IV U105 ( .A(B[20]), .Z(n280) );
  IV U106 ( .A(B[21]), .Z(n281) );
  IV U107 ( .A(B[22]), .Z(n282) );
  IV U108 ( .A(B[23]), .Z(n283) );
  IV U109 ( .A(B[24]), .Z(n284) );
  IV U110 ( .A(B[25]), .Z(n285) );
  IV U111 ( .A(B[26]), .Z(n286) );
  IV U112 ( .A(B[27]), .Z(n287) );
  IV U113 ( .A(B[28]), .Z(n288) );
  IV U114 ( .A(B[235]), .Z(n495) );
  IV U115 ( .A(B[29]), .Z(n289) );
  IV U116 ( .A(B[30]), .Z(n290) );
  IV U117 ( .A(B[31]), .Z(n291) );
  IV U118 ( .A(B[32]), .Z(n292) );
  IV U119 ( .A(B[33]), .Z(n293) );
  IV U120 ( .A(B[34]), .Z(n294) );
  IV U121 ( .A(B[35]), .Z(n295) );
  IV U122 ( .A(B[36]), .Z(n296) );
  IV U123 ( .A(B[37]), .Z(n297) );
  IV U124 ( .A(B[38]), .Z(n298) );
  IV U125 ( .A(B[236]), .Z(n496) );
  IV U126 ( .A(B[39]), .Z(n299) );
  IV U127 ( .A(B[40]), .Z(n300) );
  IV U128 ( .A(B[41]), .Z(n301) );
  IV U129 ( .A(B[42]), .Z(n302) );
  IV U130 ( .A(B[43]), .Z(n303) );
  IV U131 ( .A(B[44]), .Z(n304) );
  IV U132 ( .A(B[45]), .Z(n305) );
  IV U133 ( .A(B[46]), .Z(n306) );
  IV U134 ( .A(B[47]), .Z(n307) );
  IV U135 ( .A(B[48]), .Z(n308) );
  IV U136 ( .A(B[237]), .Z(n497) );
  IV U137 ( .A(B[49]), .Z(n309) );
  IV U138 ( .A(B[50]), .Z(n310) );
  IV U139 ( .A(B[51]), .Z(n311) );
  IV U140 ( .A(B[52]), .Z(n312) );
  IV U141 ( .A(B[53]), .Z(n313) );
  IV U142 ( .A(B[54]), .Z(n314) );
  IV U143 ( .A(B[55]), .Z(n315) );
  IV U144 ( .A(B[56]), .Z(n316) );
  IV U145 ( .A(B[57]), .Z(n317) );
  IV U146 ( .A(B[58]), .Z(n318) );
  IV U147 ( .A(B[238]), .Z(n498) );
  IV U148 ( .A(B[256]), .Z(n516) );
  IV U149 ( .A(B[59]), .Z(n319) );
  IV U150 ( .A(B[60]), .Z(n320) );
  IV U151 ( .A(B[61]), .Z(n321) );
  IV U152 ( .A(B[62]), .Z(n322) );
  IV U153 ( .A(B[63]), .Z(n323) );
  IV U154 ( .A(B[64]), .Z(n324) );
  IV U155 ( .A(B[65]), .Z(n325) );
  IV U156 ( .A(B[66]), .Z(n326) );
  IV U157 ( .A(B[67]), .Z(n327) );
  IV U158 ( .A(B[68]), .Z(n328) );
  IV U159 ( .A(B[239]), .Z(n499) );
  IV U160 ( .A(B[69]), .Z(n329) );
  IV U161 ( .A(B[70]), .Z(n330) );
  IV U162 ( .A(B[71]), .Z(n331) );
  IV U163 ( .A(B[72]), .Z(n332) );
  IV U164 ( .A(B[73]), .Z(n333) );
  IV U165 ( .A(B[74]), .Z(n334) );
  IV U166 ( .A(B[75]), .Z(n335) );
  IV U167 ( .A(B[76]), .Z(n336) );
  IV U168 ( .A(B[77]), .Z(n337) );
  IV U169 ( .A(B[78]), .Z(n338) );
  IV U170 ( .A(B[240]), .Z(n500) );
  IV U171 ( .A(B[79]), .Z(n339) );
  IV U172 ( .A(B[80]), .Z(n340) );
  IV U173 ( .A(B[81]), .Z(n341) );
  IV U174 ( .A(B[82]), .Z(n342) );
  IV U175 ( .A(B[83]), .Z(n343) );
  IV U176 ( .A(B[84]), .Z(n344) );
  IV U177 ( .A(B[85]), .Z(n345) );
  IV U178 ( .A(B[86]), .Z(n346) );
  IV U179 ( .A(B[87]), .Z(n347) );
  IV U180 ( .A(B[88]), .Z(n348) );
  IV U181 ( .A(B[241]), .Z(n501) );
  IV U182 ( .A(B[89]), .Z(n349) );
  IV U183 ( .A(B[90]), .Z(n350) );
  IV U184 ( .A(B[91]), .Z(n351) );
  IV U185 ( .A(B[92]), .Z(n352) );
  IV U186 ( .A(B[93]), .Z(n353) );
  IV U187 ( .A(B[94]), .Z(n354) );
  IV U188 ( .A(B[95]), .Z(n355) );
  IV U189 ( .A(B[96]), .Z(n356) );
  IV U190 ( .A(B[97]), .Z(n357) );
  IV U191 ( .A(B[98]), .Z(n358) );
  IV U192 ( .A(B[242]), .Z(n502) );
  IV U193 ( .A(B[99]), .Z(n359) );
  IV U194 ( .A(B[100]), .Z(n360) );
  IV U195 ( .A(B[101]), .Z(n361) );
  IV U196 ( .A(B[102]), .Z(n362) );
  IV U197 ( .A(B[103]), .Z(n363) );
  IV U198 ( .A(B[104]), .Z(n364) );
  IV U199 ( .A(B[105]), .Z(n365) );
  IV U200 ( .A(B[106]), .Z(n366) );
  IV U201 ( .A(B[107]), .Z(n367) );
  IV U202 ( .A(B[108]), .Z(n368) );
  IV U203 ( .A(B[243]), .Z(n503) );
  IV U204 ( .A(B[109]), .Z(n369) );
  IV U205 ( .A(B[110]), .Z(n370) );
  IV U206 ( .A(B[111]), .Z(n371) );
  IV U207 ( .A(B[112]), .Z(n372) );
  IV U208 ( .A(B[113]), .Z(n373) );
  IV U209 ( .A(B[114]), .Z(n374) );
  IV U210 ( .A(B[115]), .Z(n375) );
  IV U211 ( .A(B[116]), .Z(n376) );
  IV U212 ( .A(B[117]), .Z(n377) );
  IV U213 ( .A(B[118]), .Z(n378) );
  IV U214 ( .A(B[244]), .Z(n504) );
  IV U215 ( .A(B[119]), .Z(n379) );
  IV U216 ( .A(B[120]), .Z(n380) );
  IV U217 ( .A(B[121]), .Z(n381) );
  IV U218 ( .A(B[122]), .Z(n382) );
  IV U219 ( .A(B[123]), .Z(n383) );
  IV U220 ( .A(B[124]), .Z(n384) );
  IV U221 ( .A(B[125]), .Z(n385) );
  IV U222 ( .A(B[126]), .Z(n386) );
  IV U223 ( .A(B[127]), .Z(n387) );
  IV U224 ( .A(B[128]), .Z(n388) );
  IV U225 ( .A(B[245]), .Z(n505) );
  IV U226 ( .A(B[129]), .Z(n389) );
  IV U227 ( .A(B[130]), .Z(n390) );
  IV U228 ( .A(B[131]), .Z(n391) );
  IV U229 ( .A(B[132]), .Z(n392) );
  IV U230 ( .A(B[133]), .Z(n393) );
  IV U231 ( .A(B[134]), .Z(n394) );
  IV U232 ( .A(B[135]), .Z(n395) );
  IV U233 ( .A(B[136]), .Z(n396) );
  IV U234 ( .A(B[137]), .Z(n397) );
  IV U235 ( .A(B[138]), .Z(n398) );
  IV U236 ( .A(B[246]), .Z(n506) );
  IV U237 ( .A(B[139]), .Z(n399) );
  IV U238 ( .A(B[140]), .Z(n400) );
  IV U239 ( .A(B[141]), .Z(n401) );
  IV U240 ( .A(B[142]), .Z(n402) );
  IV U241 ( .A(B[143]), .Z(n403) );
  IV U242 ( .A(B[144]), .Z(n404) );
  IV U243 ( .A(B[145]), .Z(n405) );
  IV U244 ( .A(B[146]), .Z(n406) );
  IV U245 ( .A(B[147]), .Z(n407) );
  IV U246 ( .A(B[148]), .Z(n408) );
  IV U247 ( .A(B[247]), .Z(n507) );
  IV U248 ( .A(B[149]), .Z(n409) );
  IV U249 ( .A(B[150]), .Z(n410) );
  IV U250 ( .A(B[151]), .Z(n411) );
  IV U251 ( .A(B[152]), .Z(n412) );
  IV U252 ( .A(B[153]), .Z(n413) );
  IV U253 ( .A(B[154]), .Z(n414) );
  IV U254 ( .A(B[155]), .Z(n415) );
  IV U255 ( .A(B[156]), .Z(n416) );
  IV U256 ( .A(B[157]), .Z(n417) );
  IV U257 ( .A(B[158]), .Z(n418) );
  IV U258 ( .A(B[248]), .Z(n508) );
  IV U259 ( .A(B[257]), .Z(n517) );
endmodule


module FA_2581 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XNOR U1 ( .A(CI), .B(A), .Z(S) );
endmodule


module FA_2582 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2583 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2584 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2585 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2586 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2587 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2588 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2589 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2590 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2591 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2592 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2593 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2594 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2595 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2596 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2597 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2598 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2599 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2600 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2601 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2602 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2603 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2604 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2605 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2606 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2607 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2608 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2609 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2610 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2611 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2612 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2613 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2614 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2615 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2616 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2617 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2618 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2619 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2620 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2621 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2622 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2623 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2624 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2625 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2626 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2627 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2628 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2629 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2630 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2631 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2632 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2633 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2634 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2635 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2636 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2637 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2638 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2639 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2640 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2641 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2642 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2643 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2644 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2645 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2646 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2647 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2648 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2649 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2650 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2651 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2652 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2653 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2654 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2655 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2656 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2657 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2658 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2659 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2660 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2661 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2662 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2663 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2664 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2665 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2666 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2667 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2668 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2669 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2670 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2671 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2672 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2673 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2674 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2675 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2676 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2677 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2678 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2679 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2680 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2681 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2682 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2683 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2684 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2685 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2686 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2687 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2688 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2689 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2690 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2691 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2692 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2693 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2694 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2695 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2696 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2697 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2698 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2699 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2700 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2701 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2702 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2703 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2704 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2705 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2706 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2707 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2708 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2709 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2710 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2711 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2712 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2713 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2714 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2715 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2716 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2717 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2718 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2719 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2720 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2721 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2722 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2723 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2724 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2725 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2726 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2727 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2728 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2729 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2730 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2731 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2732 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2733 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2734 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2735 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2736 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2737 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2738 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2739 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2740 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2741 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2742 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2743 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2744 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2745 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2746 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2747 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2748 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2749 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2750 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2751 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2752 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2753 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2754 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2755 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2756 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2757 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2758 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2759 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2760 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2761 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2762 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2763 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2764 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2765 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2766 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2767 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2768 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2769 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2770 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2771 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2772 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2773 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2774 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2775 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2776 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2777 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2778 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2779 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2780 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2781 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2782 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2783 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2784 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2785 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2786 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2787 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2788 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2789 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2790 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2791 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2792 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2793 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2794 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2795 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2796 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2797 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2798 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2799 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2800 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2801 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2802 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2803 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2804 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2805 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2806 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2807 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2808 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2809 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2810 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2811 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2812 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2813 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2814 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2815 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2816 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2817 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2818 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2819 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2820 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2821 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2822 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2823 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2824 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2825 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2826 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2827 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2828 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2829 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2830 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2831 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2832 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2833 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2834 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2835 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2836 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2837 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XNOR U1 ( .A(B), .B(A), .Z(S) );
  OR U2 ( .A(B), .B(A), .Z(CO) );
endmodule


module SUB_N258_5 ( A, B, S, CO );
  input [257:0] A;
  input [257:0] B;
  output [257:0] S;
  output CO;
  wire   n2, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512;
  wire   [257:1] C;

  FA_2837 \FAINST[0].FA_  ( .A(A[0]), .B(n2), .CI(1'b1), .S(S[0]), .CO(C[1])
         );
  FA_2836 \FAINST[1].FA_  ( .A(A[1]), .B(n258), .CI(C[1]), .S(S[1]), .CO(C[2])
         );
  FA_2835 \FAINST[2].FA_  ( .A(A[2]), .B(n259), .CI(C[2]), .S(S[2]), .CO(C[3])
         );
  FA_2834 \FAINST[3].FA_  ( .A(A[3]), .B(n260), .CI(C[3]), .S(S[3]), .CO(C[4])
         );
  FA_2833 \FAINST[4].FA_  ( .A(A[4]), .B(n261), .CI(C[4]), .S(S[4]), .CO(C[5])
         );
  FA_2832 \FAINST[5].FA_  ( .A(A[5]), .B(n262), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_2831 \FAINST[6].FA_  ( .A(A[6]), .B(n263), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_2830 \FAINST[7].FA_  ( .A(A[7]), .B(n264), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_2829 \FAINST[8].FA_  ( .A(A[8]), .B(n265), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_2828 \FAINST[9].FA_  ( .A(A[9]), .B(n266), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_2827 \FAINST[10].FA_  ( .A(A[10]), .B(n267), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_2826 \FAINST[11].FA_  ( .A(A[11]), .B(n268), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_2825 \FAINST[12].FA_  ( .A(A[12]), .B(n269), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_2824 \FAINST[13].FA_  ( .A(A[13]), .B(n270), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_2823 \FAINST[14].FA_  ( .A(A[14]), .B(n271), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_2822 \FAINST[15].FA_  ( .A(A[15]), .B(n272), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_2821 \FAINST[16].FA_  ( .A(A[16]), .B(n273), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_2820 \FAINST[17].FA_  ( .A(A[17]), .B(n274), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_2819 \FAINST[18].FA_  ( .A(A[18]), .B(n275), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_2818 \FAINST[19].FA_  ( .A(A[19]), .B(n276), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_2817 \FAINST[20].FA_  ( .A(A[20]), .B(n277), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_2816 \FAINST[21].FA_  ( .A(A[21]), .B(n278), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_2815 \FAINST[22].FA_  ( .A(A[22]), .B(n279), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_2814 \FAINST[23].FA_  ( .A(A[23]), .B(n280), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_2813 \FAINST[24].FA_  ( .A(A[24]), .B(n281), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_2812 \FAINST[25].FA_  ( .A(A[25]), .B(n282), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_2811 \FAINST[26].FA_  ( .A(A[26]), .B(n283), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_2810 \FAINST[27].FA_  ( .A(A[27]), .B(n284), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_2809 \FAINST[28].FA_  ( .A(A[28]), .B(n285), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_2808 \FAINST[29].FA_  ( .A(A[29]), .B(n286), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_2807 \FAINST[30].FA_  ( .A(A[30]), .B(n287), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_2806 \FAINST[31].FA_  ( .A(A[31]), .B(n288), .CI(C[31]), .S(S[31]), .CO(
        C[32]) );
  FA_2805 \FAINST[32].FA_  ( .A(A[32]), .B(n289), .CI(C[32]), .S(S[32]), .CO(
        C[33]) );
  FA_2804 \FAINST[33].FA_  ( .A(A[33]), .B(n290), .CI(C[33]), .S(S[33]), .CO(
        C[34]) );
  FA_2803 \FAINST[34].FA_  ( .A(A[34]), .B(n291), .CI(C[34]), .S(S[34]), .CO(
        C[35]) );
  FA_2802 \FAINST[35].FA_  ( .A(A[35]), .B(n292), .CI(C[35]), .S(S[35]), .CO(
        C[36]) );
  FA_2801 \FAINST[36].FA_  ( .A(A[36]), .B(n293), .CI(C[36]), .S(S[36]), .CO(
        C[37]) );
  FA_2800 \FAINST[37].FA_  ( .A(A[37]), .B(n294), .CI(C[37]), .S(S[37]), .CO(
        C[38]) );
  FA_2799 \FAINST[38].FA_  ( .A(A[38]), .B(n295), .CI(C[38]), .S(S[38]), .CO(
        C[39]) );
  FA_2798 \FAINST[39].FA_  ( .A(A[39]), .B(n296), .CI(C[39]), .S(S[39]), .CO(
        C[40]) );
  FA_2797 \FAINST[40].FA_  ( .A(A[40]), .B(n297), .CI(C[40]), .S(S[40]), .CO(
        C[41]) );
  FA_2796 \FAINST[41].FA_  ( .A(A[41]), .B(n298), .CI(C[41]), .S(S[41]), .CO(
        C[42]) );
  FA_2795 \FAINST[42].FA_  ( .A(A[42]), .B(n299), .CI(C[42]), .S(S[42]), .CO(
        C[43]) );
  FA_2794 \FAINST[43].FA_  ( .A(A[43]), .B(n300), .CI(C[43]), .S(S[43]), .CO(
        C[44]) );
  FA_2793 \FAINST[44].FA_  ( .A(A[44]), .B(n301), .CI(C[44]), .S(S[44]), .CO(
        C[45]) );
  FA_2792 \FAINST[45].FA_  ( .A(A[45]), .B(n302), .CI(C[45]), .S(S[45]), .CO(
        C[46]) );
  FA_2791 \FAINST[46].FA_  ( .A(A[46]), .B(n303), .CI(C[46]), .S(S[46]), .CO(
        C[47]) );
  FA_2790 \FAINST[47].FA_  ( .A(A[47]), .B(n304), .CI(C[47]), .S(S[47]), .CO(
        C[48]) );
  FA_2789 \FAINST[48].FA_  ( .A(A[48]), .B(n305), .CI(C[48]), .S(S[48]), .CO(
        C[49]) );
  FA_2788 \FAINST[49].FA_  ( .A(A[49]), .B(n306), .CI(C[49]), .S(S[49]), .CO(
        C[50]) );
  FA_2787 \FAINST[50].FA_  ( .A(A[50]), .B(n307), .CI(C[50]), .S(S[50]), .CO(
        C[51]) );
  FA_2786 \FAINST[51].FA_  ( .A(A[51]), .B(n308), .CI(C[51]), .S(S[51]), .CO(
        C[52]) );
  FA_2785 \FAINST[52].FA_  ( .A(A[52]), .B(n309), .CI(C[52]), .S(S[52]), .CO(
        C[53]) );
  FA_2784 \FAINST[53].FA_  ( .A(A[53]), .B(n310), .CI(C[53]), .S(S[53]), .CO(
        C[54]) );
  FA_2783 \FAINST[54].FA_  ( .A(A[54]), .B(n311), .CI(C[54]), .S(S[54]), .CO(
        C[55]) );
  FA_2782 \FAINST[55].FA_  ( .A(A[55]), .B(n312), .CI(C[55]), .S(S[55]), .CO(
        C[56]) );
  FA_2781 \FAINST[56].FA_  ( .A(A[56]), .B(n313), .CI(C[56]), .S(S[56]), .CO(
        C[57]) );
  FA_2780 \FAINST[57].FA_  ( .A(A[57]), .B(n314), .CI(C[57]), .S(S[57]), .CO(
        C[58]) );
  FA_2779 \FAINST[58].FA_  ( .A(A[58]), .B(n315), .CI(C[58]), .S(S[58]), .CO(
        C[59]) );
  FA_2778 \FAINST[59].FA_  ( .A(A[59]), .B(n316), .CI(C[59]), .S(S[59]), .CO(
        C[60]) );
  FA_2777 \FAINST[60].FA_  ( .A(A[60]), .B(n317), .CI(C[60]), .S(S[60]), .CO(
        C[61]) );
  FA_2776 \FAINST[61].FA_  ( .A(A[61]), .B(n318), .CI(C[61]), .S(S[61]), .CO(
        C[62]) );
  FA_2775 \FAINST[62].FA_  ( .A(A[62]), .B(n319), .CI(C[62]), .S(S[62]), .CO(
        C[63]) );
  FA_2774 \FAINST[63].FA_  ( .A(A[63]), .B(n320), .CI(C[63]), .S(S[63]), .CO(
        C[64]) );
  FA_2773 \FAINST[64].FA_  ( .A(A[64]), .B(n321), .CI(C[64]), .S(S[64]), .CO(
        C[65]) );
  FA_2772 \FAINST[65].FA_  ( .A(A[65]), .B(n322), .CI(C[65]), .S(S[65]), .CO(
        C[66]) );
  FA_2771 \FAINST[66].FA_  ( .A(A[66]), .B(n323), .CI(C[66]), .S(S[66]), .CO(
        C[67]) );
  FA_2770 \FAINST[67].FA_  ( .A(A[67]), .B(n324), .CI(C[67]), .S(S[67]), .CO(
        C[68]) );
  FA_2769 \FAINST[68].FA_  ( .A(A[68]), .B(n325), .CI(C[68]), .S(S[68]), .CO(
        C[69]) );
  FA_2768 \FAINST[69].FA_  ( .A(A[69]), .B(n326), .CI(C[69]), .S(S[69]), .CO(
        C[70]) );
  FA_2767 \FAINST[70].FA_  ( .A(A[70]), .B(n327), .CI(C[70]), .S(S[70]), .CO(
        C[71]) );
  FA_2766 \FAINST[71].FA_  ( .A(A[71]), .B(n328), .CI(C[71]), .S(S[71]), .CO(
        C[72]) );
  FA_2765 \FAINST[72].FA_  ( .A(A[72]), .B(n329), .CI(C[72]), .S(S[72]), .CO(
        C[73]) );
  FA_2764 \FAINST[73].FA_  ( .A(A[73]), .B(n330), .CI(C[73]), .S(S[73]), .CO(
        C[74]) );
  FA_2763 \FAINST[74].FA_  ( .A(A[74]), .B(n331), .CI(C[74]), .S(S[74]), .CO(
        C[75]) );
  FA_2762 \FAINST[75].FA_  ( .A(A[75]), .B(n332), .CI(C[75]), .S(S[75]), .CO(
        C[76]) );
  FA_2761 \FAINST[76].FA_  ( .A(A[76]), .B(n333), .CI(C[76]), .S(S[76]), .CO(
        C[77]) );
  FA_2760 \FAINST[77].FA_  ( .A(A[77]), .B(n334), .CI(C[77]), .S(S[77]), .CO(
        C[78]) );
  FA_2759 \FAINST[78].FA_  ( .A(A[78]), .B(n335), .CI(C[78]), .S(S[78]), .CO(
        C[79]) );
  FA_2758 \FAINST[79].FA_  ( .A(A[79]), .B(n336), .CI(C[79]), .S(S[79]), .CO(
        C[80]) );
  FA_2757 \FAINST[80].FA_  ( .A(A[80]), .B(n337), .CI(C[80]), .S(S[80]), .CO(
        C[81]) );
  FA_2756 \FAINST[81].FA_  ( .A(A[81]), .B(n338), .CI(C[81]), .S(S[81]), .CO(
        C[82]) );
  FA_2755 \FAINST[82].FA_  ( .A(A[82]), .B(n339), .CI(C[82]), .S(S[82]), .CO(
        C[83]) );
  FA_2754 \FAINST[83].FA_  ( .A(A[83]), .B(n340), .CI(C[83]), .S(S[83]), .CO(
        C[84]) );
  FA_2753 \FAINST[84].FA_  ( .A(A[84]), .B(n341), .CI(C[84]), .S(S[84]), .CO(
        C[85]) );
  FA_2752 \FAINST[85].FA_  ( .A(A[85]), .B(n342), .CI(C[85]), .S(S[85]), .CO(
        C[86]) );
  FA_2751 \FAINST[86].FA_  ( .A(A[86]), .B(n343), .CI(C[86]), .S(S[86]), .CO(
        C[87]) );
  FA_2750 \FAINST[87].FA_  ( .A(A[87]), .B(n344), .CI(C[87]), .S(S[87]), .CO(
        C[88]) );
  FA_2749 \FAINST[88].FA_  ( .A(A[88]), .B(n345), .CI(C[88]), .S(S[88]), .CO(
        C[89]) );
  FA_2748 \FAINST[89].FA_  ( .A(A[89]), .B(n346), .CI(C[89]), .S(S[89]), .CO(
        C[90]) );
  FA_2747 \FAINST[90].FA_  ( .A(A[90]), .B(n347), .CI(C[90]), .S(S[90]), .CO(
        C[91]) );
  FA_2746 \FAINST[91].FA_  ( .A(A[91]), .B(n348), .CI(C[91]), .S(S[91]), .CO(
        C[92]) );
  FA_2745 \FAINST[92].FA_  ( .A(A[92]), .B(n349), .CI(C[92]), .S(S[92]), .CO(
        C[93]) );
  FA_2744 \FAINST[93].FA_  ( .A(A[93]), .B(n350), .CI(C[93]), .S(S[93]), .CO(
        C[94]) );
  FA_2743 \FAINST[94].FA_  ( .A(A[94]), .B(n351), .CI(C[94]), .S(S[94]), .CO(
        C[95]) );
  FA_2742 \FAINST[95].FA_  ( .A(A[95]), .B(n352), .CI(C[95]), .S(S[95]), .CO(
        C[96]) );
  FA_2741 \FAINST[96].FA_  ( .A(A[96]), .B(n353), .CI(C[96]), .S(S[96]), .CO(
        C[97]) );
  FA_2740 \FAINST[97].FA_  ( .A(A[97]), .B(n354), .CI(C[97]), .S(S[97]), .CO(
        C[98]) );
  FA_2739 \FAINST[98].FA_  ( .A(A[98]), .B(n355), .CI(C[98]), .S(S[98]), .CO(
        C[99]) );
  FA_2738 \FAINST[99].FA_  ( .A(A[99]), .B(n356), .CI(C[99]), .S(S[99]), .CO(
        C[100]) );
  FA_2737 \FAINST[100].FA_  ( .A(A[100]), .B(n357), .CI(C[100]), .S(S[100]), 
        .CO(C[101]) );
  FA_2736 \FAINST[101].FA_  ( .A(A[101]), .B(n358), .CI(C[101]), .S(S[101]), 
        .CO(C[102]) );
  FA_2735 \FAINST[102].FA_  ( .A(A[102]), .B(n359), .CI(C[102]), .S(S[102]), 
        .CO(C[103]) );
  FA_2734 \FAINST[103].FA_  ( .A(A[103]), .B(n360), .CI(C[103]), .S(S[103]), 
        .CO(C[104]) );
  FA_2733 \FAINST[104].FA_  ( .A(A[104]), .B(n361), .CI(C[104]), .S(S[104]), 
        .CO(C[105]) );
  FA_2732 \FAINST[105].FA_  ( .A(A[105]), .B(n362), .CI(C[105]), .S(S[105]), 
        .CO(C[106]) );
  FA_2731 \FAINST[106].FA_  ( .A(A[106]), .B(n363), .CI(C[106]), .S(S[106]), 
        .CO(C[107]) );
  FA_2730 \FAINST[107].FA_  ( .A(A[107]), .B(n364), .CI(C[107]), .S(S[107]), 
        .CO(C[108]) );
  FA_2729 \FAINST[108].FA_  ( .A(A[108]), .B(n365), .CI(C[108]), .S(S[108]), 
        .CO(C[109]) );
  FA_2728 \FAINST[109].FA_  ( .A(A[109]), .B(n366), .CI(C[109]), .S(S[109]), 
        .CO(C[110]) );
  FA_2727 \FAINST[110].FA_  ( .A(A[110]), .B(n367), .CI(C[110]), .S(S[110]), 
        .CO(C[111]) );
  FA_2726 \FAINST[111].FA_  ( .A(A[111]), .B(n368), .CI(C[111]), .S(S[111]), 
        .CO(C[112]) );
  FA_2725 \FAINST[112].FA_  ( .A(A[112]), .B(n369), .CI(C[112]), .S(S[112]), 
        .CO(C[113]) );
  FA_2724 \FAINST[113].FA_  ( .A(A[113]), .B(n370), .CI(C[113]), .S(S[113]), 
        .CO(C[114]) );
  FA_2723 \FAINST[114].FA_  ( .A(A[114]), .B(n371), .CI(C[114]), .S(S[114]), 
        .CO(C[115]) );
  FA_2722 \FAINST[115].FA_  ( .A(A[115]), .B(n372), .CI(C[115]), .S(S[115]), 
        .CO(C[116]) );
  FA_2721 \FAINST[116].FA_  ( .A(A[116]), .B(n373), .CI(C[116]), .S(S[116]), 
        .CO(C[117]) );
  FA_2720 \FAINST[117].FA_  ( .A(A[117]), .B(n374), .CI(C[117]), .S(S[117]), 
        .CO(C[118]) );
  FA_2719 \FAINST[118].FA_  ( .A(A[118]), .B(n375), .CI(C[118]), .S(S[118]), 
        .CO(C[119]) );
  FA_2718 \FAINST[119].FA_  ( .A(A[119]), .B(n376), .CI(C[119]), .S(S[119]), 
        .CO(C[120]) );
  FA_2717 \FAINST[120].FA_  ( .A(A[120]), .B(n377), .CI(C[120]), .S(S[120]), 
        .CO(C[121]) );
  FA_2716 \FAINST[121].FA_  ( .A(A[121]), .B(n378), .CI(C[121]), .S(S[121]), 
        .CO(C[122]) );
  FA_2715 \FAINST[122].FA_  ( .A(A[122]), .B(n379), .CI(C[122]), .S(S[122]), 
        .CO(C[123]) );
  FA_2714 \FAINST[123].FA_  ( .A(A[123]), .B(n380), .CI(C[123]), .S(S[123]), 
        .CO(C[124]) );
  FA_2713 \FAINST[124].FA_  ( .A(A[124]), .B(n381), .CI(C[124]), .S(S[124]), 
        .CO(C[125]) );
  FA_2712 \FAINST[125].FA_  ( .A(A[125]), .B(n382), .CI(C[125]), .S(S[125]), 
        .CO(C[126]) );
  FA_2711 \FAINST[126].FA_  ( .A(A[126]), .B(n383), .CI(C[126]), .S(S[126]), 
        .CO(C[127]) );
  FA_2710 \FAINST[127].FA_  ( .A(A[127]), .B(n384), .CI(C[127]), .S(S[127]), 
        .CO(C[128]) );
  FA_2709 \FAINST[128].FA_  ( .A(A[128]), .B(n385), .CI(C[128]), .S(S[128]), 
        .CO(C[129]) );
  FA_2708 \FAINST[129].FA_  ( .A(A[129]), .B(n386), .CI(C[129]), .S(S[129]), 
        .CO(C[130]) );
  FA_2707 \FAINST[130].FA_  ( .A(A[130]), .B(n387), .CI(C[130]), .S(S[130]), 
        .CO(C[131]) );
  FA_2706 \FAINST[131].FA_  ( .A(A[131]), .B(n388), .CI(C[131]), .S(S[131]), 
        .CO(C[132]) );
  FA_2705 \FAINST[132].FA_  ( .A(A[132]), .B(n389), .CI(C[132]), .S(S[132]), 
        .CO(C[133]) );
  FA_2704 \FAINST[133].FA_  ( .A(A[133]), .B(n390), .CI(C[133]), .S(S[133]), 
        .CO(C[134]) );
  FA_2703 \FAINST[134].FA_  ( .A(A[134]), .B(n391), .CI(C[134]), .S(S[134]), 
        .CO(C[135]) );
  FA_2702 \FAINST[135].FA_  ( .A(A[135]), .B(n392), .CI(C[135]), .S(S[135]), 
        .CO(C[136]) );
  FA_2701 \FAINST[136].FA_  ( .A(A[136]), .B(n393), .CI(C[136]), .S(S[136]), 
        .CO(C[137]) );
  FA_2700 \FAINST[137].FA_  ( .A(A[137]), .B(n394), .CI(C[137]), .S(S[137]), 
        .CO(C[138]) );
  FA_2699 \FAINST[138].FA_  ( .A(A[138]), .B(n395), .CI(C[138]), .S(S[138]), 
        .CO(C[139]) );
  FA_2698 \FAINST[139].FA_  ( .A(A[139]), .B(n396), .CI(C[139]), .S(S[139]), 
        .CO(C[140]) );
  FA_2697 \FAINST[140].FA_  ( .A(A[140]), .B(n397), .CI(C[140]), .S(S[140]), 
        .CO(C[141]) );
  FA_2696 \FAINST[141].FA_  ( .A(A[141]), .B(n398), .CI(C[141]), .S(S[141]), 
        .CO(C[142]) );
  FA_2695 \FAINST[142].FA_  ( .A(A[142]), .B(n399), .CI(C[142]), .S(S[142]), 
        .CO(C[143]) );
  FA_2694 \FAINST[143].FA_  ( .A(A[143]), .B(n400), .CI(C[143]), .S(S[143]), 
        .CO(C[144]) );
  FA_2693 \FAINST[144].FA_  ( .A(A[144]), .B(n401), .CI(C[144]), .S(S[144]), 
        .CO(C[145]) );
  FA_2692 \FAINST[145].FA_  ( .A(A[145]), .B(n402), .CI(C[145]), .S(S[145]), 
        .CO(C[146]) );
  FA_2691 \FAINST[146].FA_  ( .A(A[146]), .B(n403), .CI(C[146]), .S(S[146]), 
        .CO(C[147]) );
  FA_2690 \FAINST[147].FA_  ( .A(A[147]), .B(n404), .CI(C[147]), .S(S[147]), 
        .CO(C[148]) );
  FA_2689 \FAINST[148].FA_  ( .A(A[148]), .B(n405), .CI(C[148]), .S(S[148]), 
        .CO(C[149]) );
  FA_2688 \FAINST[149].FA_  ( .A(A[149]), .B(n406), .CI(C[149]), .S(S[149]), 
        .CO(C[150]) );
  FA_2687 \FAINST[150].FA_  ( .A(A[150]), .B(n407), .CI(C[150]), .S(S[150]), 
        .CO(C[151]) );
  FA_2686 \FAINST[151].FA_  ( .A(A[151]), .B(n408), .CI(C[151]), .S(S[151]), 
        .CO(C[152]) );
  FA_2685 \FAINST[152].FA_  ( .A(A[152]), .B(n409), .CI(C[152]), .S(S[152]), 
        .CO(C[153]) );
  FA_2684 \FAINST[153].FA_  ( .A(A[153]), .B(n410), .CI(C[153]), .S(S[153]), 
        .CO(C[154]) );
  FA_2683 \FAINST[154].FA_  ( .A(A[154]), .B(n411), .CI(C[154]), .S(S[154]), 
        .CO(C[155]) );
  FA_2682 \FAINST[155].FA_  ( .A(A[155]), .B(n412), .CI(C[155]), .S(S[155]), 
        .CO(C[156]) );
  FA_2681 \FAINST[156].FA_  ( .A(A[156]), .B(n413), .CI(C[156]), .S(S[156]), 
        .CO(C[157]) );
  FA_2680 \FAINST[157].FA_  ( .A(A[157]), .B(n414), .CI(C[157]), .S(S[157]), 
        .CO(C[158]) );
  FA_2679 \FAINST[158].FA_  ( .A(A[158]), .B(n415), .CI(C[158]), .S(S[158]), 
        .CO(C[159]) );
  FA_2678 \FAINST[159].FA_  ( .A(A[159]), .B(n416), .CI(C[159]), .S(S[159]), 
        .CO(C[160]) );
  FA_2677 \FAINST[160].FA_  ( .A(A[160]), .B(n417), .CI(C[160]), .S(S[160]), 
        .CO(C[161]) );
  FA_2676 \FAINST[161].FA_  ( .A(A[161]), .B(n418), .CI(C[161]), .S(S[161]), 
        .CO(C[162]) );
  FA_2675 \FAINST[162].FA_  ( .A(A[162]), .B(n419), .CI(C[162]), .S(S[162]), 
        .CO(C[163]) );
  FA_2674 \FAINST[163].FA_  ( .A(A[163]), .B(n420), .CI(C[163]), .S(S[163]), 
        .CO(C[164]) );
  FA_2673 \FAINST[164].FA_  ( .A(A[164]), .B(n421), .CI(C[164]), .S(S[164]), 
        .CO(C[165]) );
  FA_2672 \FAINST[165].FA_  ( .A(A[165]), .B(n422), .CI(C[165]), .S(S[165]), 
        .CO(C[166]) );
  FA_2671 \FAINST[166].FA_  ( .A(A[166]), .B(n423), .CI(C[166]), .S(S[166]), 
        .CO(C[167]) );
  FA_2670 \FAINST[167].FA_  ( .A(A[167]), .B(n424), .CI(C[167]), .S(S[167]), 
        .CO(C[168]) );
  FA_2669 \FAINST[168].FA_  ( .A(A[168]), .B(n425), .CI(C[168]), .S(S[168]), 
        .CO(C[169]) );
  FA_2668 \FAINST[169].FA_  ( .A(A[169]), .B(n426), .CI(C[169]), .S(S[169]), 
        .CO(C[170]) );
  FA_2667 \FAINST[170].FA_  ( .A(A[170]), .B(n427), .CI(C[170]), .S(S[170]), 
        .CO(C[171]) );
  FA_2666 \FAINST[171].FA_  ( .A(A[171]), .B(n428), .CI(C[171]), .S(S[171]), 
        .CO(C[172]) );
  FA_2665 \FAINST[172].FA_  ( .A(A[172]), .B(n429), .CI(C[172]), .S(S[172]), 
        .CO(C[173]) );
  FA_2664 \FAINST[173].FA_  ( .A(A[173]), .B(n430), .CI(C[173]), .S(S[173]), 
        .CO(C[174]) );
  FA_2663 \FAINST[174].FA_  ( .A(A[174]), .B(n431), .CI(C[174]), .S(S[174]), 
        .CO(C[175]) );
  FA_2662 \FAINST[175].FA_  ( .A(A[175]), .B(n432), .CI(C[175]), .S(S[175]), 
        .CO(C[176]) );
  FA_2661 \FAINST[176].FA_  ( .A(A[176]), .B(n433), .CI(C[176]), .S(S[176]), 
        .CO(C[177]) );
  FA_2660 \FAINST[177].FA_  ( .A(A[177]), .B(n434), .CI(C[177]), .S(S[177]), 
        .CO(C[178]) );
  FA_2659 \FAINST[178].FA_  ( .A(A[178]), .B(n435), .CI(C[178]), .S(S[178]), 
        .CO(C[179]) );
  FA_2658 \FAINST[179].FA_  ( .A(A[179]), .B(n436), .CI(C[179]), .S(S[179]), 
        .CO(C[180]) );
  FA_2657 \FAINST[180].FA_  ( .A(A[180]), .B(n437), .CI(C[180]), .S(S[180]), 
        .CO(C[181]) );
  FA_2656 \FAINST[181].FA_  ( .A(A[181]), .B(n438), .CI(C[181]), .S(S[181]), 
        .CO(C[182]) );
  FA_2655 \FAINST[182].FA_  ( .A(A[182]), .B(n439), .CI(C[182]), .S(S[182]), 
        .CO(C[183]) );
  FA_2654 \FAINST[183].FA_  ( .A(A[183]), .B(n440), .CI(C[183]), .S(S[183]), 
        .CO(C[184]) );
  FA_2653 \FAINST[184].FA_  ( .A(A[184]), .B(n441), .CI(C[184]), .S(S[184]), 
        .CO(C[185]) );
  FA_2652 \FAINST[185].FA_  ( .A(A[185]), .B(n442), .CI(C[185]), .S(S[185]), 
        .CO(C[186]) );
  FA_2651 \FAINST[186].FA_  ( .A(A[186]), .B(n443), .CI(C[186]), .S(S[186]), 
        .CO(C[187]) );
  FA_2650 \FAINST[187].FA_  ( .A(A[187]), .B(n444), .CI(C[187]), .S(S[187]), 
        .CO(C[188]) );
  FA_2649 \FAINST[188].FA_  ( .A(A[188]), .B(n445), .CI(C[188]), .S(S[188]), 
        .CO(C[189]) );
  FA_2648 \FAINST[189].FA_  ( .A(A[189]), .B(n446), .CI(C[189]), .S(S[189]), 
        .CO(C[190]) );
  FA_2647 \FAINST[190].FA_  ( .A(A[190]), .B(n447), .CI(C[190]), .S(S[190]), 
        .CO(C[191]) );
  FA_2646 \FAINST[191].FA_  ( .A(A[191]), .B(n448), .CI(C[191]), .S(S[191]), 
        .CO(C[192]) );
  FA_2645 \FAINST[192].FA_  ( .A(A[192]), .B(n449), .CI(C[192]), .S(S[192]), 
        .CO(C[193]) );
  FA_2644 \FAINST[193].FA_  ( .A(A[193]), .B(n450), .CI(C[193]), .S(S[193]), 
        .CO(C[194]) );
  FA_2643 \FAINST[194].FA_  ( .A(A[194]), .B(n451), .CI(C[194]), .S(S[194]), 
        .CO(C[195]) );
  FA_2642 \FAINST[195].FA_  ( .A(A[195]), .B(n452), .CI(C[195]), .S(S[195]), 
        .CO(C[196]) );
  FA_2641 \FAINST[196].FA_  ( .A(A[196]), .B(n453), .CI(C[196]), .S(S[196]), 
        .CO(C[197]) );
  FA_2640 \FAINST[197].FA_  ( .A(A[197]), .B(n454), .CI(C[197]), .S(S[197]), 
        .CO(C[198]) );
  FA_2639 \FAINST[198].FA_  ( .A(A[198]), .B(n455), .CI(C[198]), .S(S[198]), 
        .CO(C[199]) );
  FA_2638 \FAINST[199].FA_  ( .A(A[199]), .B(n456), .CI(C[199]), .S(S[199]), 
        .CO(C[200]) );
  FA_2637 \FAINST[200].FA_  ( .A(A[200]), .B(n457), .CI(C[200]), .S(S[200]), 
        .CO(C[201]) );
  FA_2636 \FAINST[201].FA_  ( .A(A[201]), .B(n458), .CI(C[201]), .S(S[201]), 
        .CO(C[202]) );
  FA_2635 \FAINST[202].FA_  ( .A(A[202]), .B(n459), .CI(C[202]), .S(S[202]), 
        .CO(C[203]) );
  FA_2634 \FAINST[203].FA_  ( .A(A[203]), .B(n460), .CI(C[203]), .S(S[203]), 
        .CO(C[204]) );
  FA_2633 \FAINST[204].FA_  ( .A(A[204]), .B(n461), .CI(C[204]), .S(S[204]), 
        .CO(C[205]) );
  FA_2632 \FAINST[205].FA_  ( .A(A[205]), .B(n462), .CI(C[205]), .S(S[205]), 
        .CO(C[206]) );
  FA_2631 \FAINST[206].FA_  ( .A(A[206]), .B(n463), .CI(C[206]), .S(S[206]), 
        .CO(C[207]) );
  FA_2630 \FAINST[207].FA_  ( .A(A[207]), .B(n464), .CI(C[207]), .S(S[207]), 
        .CO(C[208]) );
  FA_2629 \FAINST[208].FA_  ( .A(A[208]), .B(n465), .CI(C[208]), .S(S[208]), 
        .CO(C[209]) );
  FA_2628 \FAINST[209].FA_  ( .A(A[209]), .B(n466), .CI(C[209]), .S(S[209]), 
        .CO(C[210]) );
  FA_2627 \FAINST[210].FA_  ( .A(A[210]), .B(n467), .CI(C[210]), .S(S[210]), 
        .CO(C[211]) );
  FA_2626 \FAINST[211].FA_  ( .A(A[211]), .B(n468), .CI(C[211]), .S(S[211]), 
        .CO(C[212]) );
  FA_2625 \FAINST[212].FA_  ( .A(A[212]), .B(n469), .CI(C[212]), .S(S[212]), 
        .CO(C[213]) );
  FA_2624 \FAINST[213].FA_  ( .A(A[213]), .B(n470), .CI(C[213]), .S(S[213]), 
        .CO(C[214]) );
  FA_2623 \FAINST[214].FA_  ( .A(A[214]), .B(n471), .CI(C[214]), .S(S[214]), 
        .CO(C[215]) );
  FA_2622 \FAINST[215].FA_  ( .A(A[215]), .B(n472), .CI(C[215]), .S(S[215]), 
        .CO(C[216]) );
  FA_2621 \FAINST[216].FA_  ( .A(A[216]), .B(n473), .CI(C[216]), .S(S[216]), 
        .CO(C[217]) );
  FA_2620 \FAINST[217].FA_  ( .A(A[217]), .B(n474), .CI(C[217]), .S(S[217]), 
        .CO(C[218]) );
  FA_2619 \FAINST[218].FA_  ( .A(A[218]), .B(n475), .CI(C[218]), .S(S[218]), 
        .CO(C[219]) );
  FA_2618 \FAINST[219].FA_  ( .A(A[219]), .B(n476), .CI(C[219]), .S(S[219]), 
        .CO(C[220]) );
  FA_2617 \FAINST[220].FA_  ( .A(A[220]), .B(n477), .CI(C[220]), .S(S[220]), 
        .CO(C[221]) );
  FA_2616 \FAINST[221].FA_  ( .A(A[221]), .B(n478), .CI(C[221]), .S(S[221]), 
        .CO(C[222]) );
  FA_2615 \FAINST[222].FA_  ( .A(A[222]), .B(n479), .CI(C[222]), .S(S[222]), 
        .CO(C[223]) );
  FA_2614 \FAINST[223].FA_  ( .A(A[223]), .B(n480), .CI(C[223]), .S(S[223]), 
        .CO(C[224]) );
  FA_2613 \FAINST[224].FA_  ( .A(A[224]), .B(n481), .CI(C[224]), .S(S[224]), 
        .CO(C[225]) );
  FA_2612 \FAINST[225].FA_  ( .A(A[225]), .B(n482), .CI(C[225]), .S(S[225]), 
        .CO(C[226]) );
  FA_2611 \FAINST[226].FA_  ( .A(A[226]), .B(n483), .CI(C[226]), .S(S[226]), 
        .CO(C[227]) );
  FA_2610 \FAINST[227].FA_  ( .A(A[227]), .B(n484), .CI(C[227]), .S(S[227]), 
        .CO(C[228]) );
  FA_2609 \FAINST[228].FA_  ( .A(A[228]), .B(n485), .CI(C[228]), .S(S[228]), 
        .CO(C[229]) );
  FA_2608 \FAINST[229].FA_  ( .A(A[229]), .B(n486), .CI(C[229]), .S(S[229]), 
        .CO(C[230]) );
  FA_2607 \FAINST[230].FA_  ( .A(A[230]), .B(n487), .CI(C[230]), .S(S[230]), 
        .CO(C[231]) );
  FA_2606 \FAINST[231].FA_  ( .A(A[231]), .B(n488), .CI(C[231]), .S(S[231]), 
        .CO(C[232]) );
  FA_2605 \FAINST[232].FA_  ( .A(A[232]), .B(n489), .CI(C[232]), .S(S[232]), 
        .CO(C[233]) );
  FA_2604 \FAINST[233].FA_  ( .A(A[233]), .B(n490), .CI(C[233]), .S(S[233]), 
        .CO(C[234]) );
  FA_2603 \FAINST[234].FA_  ( .A(A[234]), .B(n491), .CI(C[234]), .S(S[234]), 
        .CO(C[235]) );
  FA_2602 \FAINST[235].FA_  ( .A(A[235]), .B(n492), .CI(C[235]), .S(S[235]), 
        .CO(C[236]) );
  FA_2601 \FAINST[236].FA_  ( .A(A[236]), .B(n493), .CI(C[236]), .S(S[236]), 
        .CO(C[237]) );
  FA_2600 \FAINST[237].FA_  ( .A(A[237]), .B(n494), .CI(C[237]), .S(S[237]), 
        .CO(C[238]) );
  FA_2599 \FAINST[238].FA_  ( .A(A[238]), .B(n495), .CI(C[238]), .S(S[238]), 
        .CO(C[239]) );
  FA_2598 \FAINST[239].FA_  ( .A(A[239]), .B(n496), .CI(C[239]), .S(S[239]), 
        .CO(C[240]) );
  FA_2597 \FAINST[240].FA_  ( .A(A[240]), .B(n497), .CI(C[240]), .S(S[240]), 
        .CO(C[241]) );
  FA_2596 \FAINST[241].FA_  ( .A(A[241]), .B(n498), .CI(C[241]), .S(S[241]), 
        .CO(C[242]) );
  FA_2595 \FAINST[242].FA_  ( .A(A[242]), .B(n499), .CI(C[242]), .S(S[242]), 
        .CO(C[243]) );
  FA_2594 \FAINST[243].FA_  ( .A(A[243]), .B(n500), .CI(C[243]), .S(S[243]), 
        .CO(C[244]) );
  FA_2593 \FAINST[244].FA_  ( .A(A[244]), .B(n501), .CI(C[244]), .S(S[244]), 
        .CO(C[245]) );
  FA_2592 \FAINST[245].FA_  ( .A(A[245]), .B(n502), .CI(C[245]), .S(S[245]), 
        .CO(C[246]) );
  FA_2591 \FAINST[246].FA_  ( .A(A[246]), .B(n503), .CI(C[246]), .S(S[246]), 
        .CO(C[247]) );
  FA_2590 \FAINST[247].FA_  ( .A(A[247]), .B(n504), .CI(C[247]), .S(S[247]), 
        .CO(C[248]) );
  FA_2589 \FAINST[248].FA_  ( .A(A[248]), .B(n505), .CI(C[248]), .S(S[248]), 
        .CO(C[249]) );
  FA_2588 \FAINST[249].FA_  ( .A(A[249]), .B(n506), .CI(C[249]), .S(S[249]), 
        .CO(C[250]) );
  FA_2587 \FAINST[250].FA_  ( .A(A[250]), .B(n507), .CI(C[250]), .S(S[250]), 
        .CO(C[251]) );
  FA_2586 \FAINST[251].FA_  ( .A(A[251]), .B(n508), .CI(C[251]), .S(S[251]), 
        .CO(C[252]) );
  FA_2585 \FAINST[252].FA_  ( .A(A[252]), .B(n509), .CI(C[252]), .S(S[252]), 
        .CO(C[253]) );
  FA_2584 \FAINST[253].FA_  ( .A(A[253]), .B(n510), .CI(C[253]), .S(S[253]), 
        .CO(C[254]) );
  FA_2583 \FAINST[254].FA_  ( .A(A[254]), .B(n511), .CI(C[254]), .S(S[254]), 
        .CO(C[255]) );
  FA_2582 \FAINST[255].FA_  ( .A(A[255]), .B(n512), .CI(C[255]), .S(S[255]), 
        .CO(C[256]) );
  FA_2581 \FAINST[256].FA_  ( .A(A[256]), .B(1'b1), .CI(C[256]), .S(S[256]) );
  IV U2 ( .A(B[159]), .Z(n416) );
  IV U3 ( .A(B[160]), .Z(n417) );
  IV U4 ( .A(B[161]), .Z(n418) );
  IV U5 ( .A(B[162]), .Z(n419) );
  IV U6 ( .A(B[163]), .Z(n420) );
  IV U7 ( .A(B[164]), .Z(n421) );
  IV U8 ( .A(B[165]), .Z(n422) );
  IV U9 ( .A(B[166]), .Z(n423) );
  IV U10 ( .A(B[167]), .Z(n424) );
  IV U11 ( .A(B[168]), .Z(n425) );
  IV U12 ( .A(B[249]), .Z(n506) );
  IV U13 ( .A(B[169]), .Z(n426) );
  IV U14 ( .A(B[170]), .Z(n427) );
  IV U15 ( .A(B[171]), .Z(n428) );
  IV U16 ( .A(B[172]), .Z(n429) );
  IV U17 ( .A(B[173]), .Z(n430) );
  IV U18 ( .A(B[174]), .Z(n431) );
  IV U19 ( .A(B[175]), .Z(n432) );
  IV U20 ( .A(B[176]), .Z(n433) );
  IV U21 ( .A(B[177]), .Z(n434) );
  IV U22 ( .A(B[178]), .Z(n435) );
  IV U23 ( .A(B[250]), .Z(n507) );
  IV U24 ( .A(B[179]), .Z(n436) );
  IV U25 ( .A(B[180]), .Z(n437) );
  IV U26 ( .A(B[181]), .Z(n438) );
  IV U27 ( .A(B[182]), .Z(n439) );
  IV U28 ( .A(B[183]), .Z(n440) );
  IV U29 ( .A(B[184]), .Z(n441) );
  IV U30 ( .A(B[185]), .Z(n442) );
  IV U31 ( .A(B[186]), .Z(n443) );
  IV U32 ( .A(B[187]), .Z(n444) );
  IV U33 ( .A(B[188]), .Z(n445) );
  IV U34 ( .A(B[251]), .Z(n508) );
  IV U35 ( .A(B[189]), .Z(n446) );
  IV U36 ( .A(B[190]), .Z(n447) );
  IV U37 ( .A(B[191]), .Z(n448) );
  IV U38 ( .A(B[192]), .Z(n449) );
  IV U39 ( .A(B[193]), .Z(n450) );
  IV U40 ( .A(B[194]), .Z(n451) );
  IV U41 ( .A(B[195]), .Z(n452) );
  IV U42 ( .A(B[196]), .Z(n453) );
  IV U43 ( .A(B[197]), .Z(n454) );
  IV U44 ( .A(B[198]), .Z(n455) );
  IV U45 ( .A(B[252]), .Z(n509) );
  IV U46 ( .A(B[199]), .Z(n456) );
  IV U47 ( .A(B[200]), .Z(n457) );
  IV U48 ( .A(B[201]), .Z(n458) );
  IV U49 ( .A(B[202]), .Z(n459) );
  IV U50 ( .A(B[203]), .Z(n460) );
  IV U51 ( .A(B[204]), .Z(n461) );
  IV U52 ( .A(B[205]), .Z(n462) );
  IV U53 ( .A(B[206]), .Z(n463) );
  IV U54 ( .A(B[207]), .Z(n464) );
  IV U55 ( .A(B[208]), .Z(n465) );
  IV U56 ( .A(B[253]), .Z(n510) );
  IV U57 ( .A(B[209]), .Z(n466) );
  IV U58 ( .A(B[210]), .Z(n467) );
  IV U59 ( .A(B[211]), .Z(n468) );
  IV U60 ( .A(B[212]), .Z(n469) );
  IV U61 ( .A(B[213]), .Z(n470) );
  IV U62 ( .A(B[214]), .Z(n471) );
  IV U63 ( .A(B[215]), .Z(n472) );
  IV U64 ( .A(B[216]), .Z(n473) );
  IV U65 ( .A(B[217]), .Z(n474) );
  IV U66 ( .A(B[218]), .Z(n475) );
  IV U67 ( .A(B[254]), .Z(n511) );
  IV U68 ( .A(B[219]), .Z(n476) );
  IV U69 ( .A(B[220]), .Z(n477) );
  IV U70 ( .A(B[221]), .Z(n478) );
  IV U71 ( .A(B[222]), .Z(n479) );
  IV U72 ( .A(B[223]), .Z(n480) );
  IV U73 ( .A(B[224]), .Z(n481) );
  IV U74 ( .A(B[225]), .Z(n482) );
  IV U75 ( .A(B[226]), .Z(n483) );
  IV U76 ( .A(B[227]), .Z(n484) );
  IV U77 ( .A(B[228]), .Z(n485) );
  IV U78 ( .A(B[255]), .Z(n512) );
  IV U79 ( .A(B[229]), .Z(n486) );
  IV U80 ( .A(B[230]), .Z(n487) );
  IV U81 ( .A(B[231]), .Z(n488) );
  IV U82 ( .A(B[232]), .Z(n489) );
  IV U83 ( .A(B[0]), .Z(n2) );
  IV U84 ( .A(B[1]), .Z(n258) );
  IV U85 ( .A(B[2]), .Z(n259) );
  IV U86 ( .A(B[3]), .Z(n260) );
  IV U87 ( .A(B[4]), .Z(n261) );
  IV U88 ( .A(B[5]), .Z(n262) );
  IV U89 ( .A(B[6]), .Z(n263) );
  IV U90 ( .A(B[7]), .Z(n264) );
  IV U91 ( .A(B[8]), .Z(n265) );
  IV U92 ( .A(B[233]), .Z(n490) );
  IV U93 ( .A(B[9]), .Z(n266) );
  IV U94 ( .A(B[10]), .Z(n267) );
  IV U95 ( .A(B[11]), .Z(n268) );
  IV U96 ( .A(B[12]), .Z(n269) );
  IV U97 ( .A(B[13]), .Z(n270) );
  IV U98 ( .A(B[14]), .Z(n271) );
  IV U99 ( .A(B[15]), .Z(n272) );
  IV U100 ( .A(B[16]), .Z(n273) );
  IV U101 ( .A(B[17]), .Z(n274) );
  IV U102 ( .A(B[18]), .Z(n275) );
  IV U103 ( .A(B[234]), .Z(n491) );
  IV U104 ( .A(B[19]), .Z(n276) );
  IV U105 ( .A(B[20]), .Z(n277) );
  IV U106 ( .A(B[21]), .Z(n278) );
  IV U107 ( .A(B[22]), .Z(n279) );
  IV U108 ( .A(B[23]), .Z(n280) );
  IV U109 ( .A(B[24]), .Z(n281) );
  IV U110 ( .A(B[25]), .Z(n282) );
  IV U111 ( .A(B[26]), .Z(n283) );
  IV U112 ( .A(B[27]), .Z(n284) );
  IV U113 ( .A(B[28]), .Z(n285) );
  IV U114 ( .A(B[235]), .Z(n492) );
  IV U115 ( .A(B[29]), .Z(n286) );
  IV U116 ( .A(B[30]), .Z(n287) );
  IV U117 ( .A(B[31]), .Z(n288) );
  IV U118 ( .A(B[32]), .Z(n289) );
  IV U119 ( .A(B[33]), .Z(n290) );
  IV U120 ( .A(B[34]), .Z(n291) );
  IV U121 ( .A(B[35]), .Z(n292) );
  IV U122 ( .A(B[36]), .Z(n293) );
  IV U123 ( .A(B[37]), .Z(n294) );
  IV U124 ( .A(B[38]), .Z(n295) );
  IV U125 ( .A(B[236]), .Z(n493) );
  IV U126 ( .A(B[39]), .Z(n296) );
  IV U127 ( .A(B[40]), .Z(n297) );
  IV U128 ( .A(B[41]), .Z(n298) );
  IV U129 ( .A(B[42]), .Z(n299) );
  IV U130 ( .A(B[43]), .Z(n300) );
  IV U131 ( .A(B[44]), .Z(n301) );
  IV U132 ( .A(B[45]), .Z(n302) );
  IV U133 ( .A(B[46]), .Z(n303) );
  IV U134 ( .A(B[47]), .Z(n304) );
  IV U135 ( .A(B[48]), .Z(n305) );
  IV U136 ( .A(B[237]), .Z(n494) );
  IV U137 ( .A(B[49]), .Z(n306) );
  IV U138 ( .A(B[50]), .Z(n307) );
  IV U139 ( .A(B[51]), .Z(n308) );
  IV U140 ( .A(B[52]), .Z(n309) );
  IV U141 ( .A(B[53]), .Z(n310) );
  IV U142 ( .A(B[54]), .Z(n311) );
  IV U143 ( .A(B[55]), .Z(n312) );
  IV U144 ( .A(B[56]), .Z(n313) );
  IV U145 ( .A(B[57]), .Z(n314) );
  IV U146 ( .A(B[58]), .Z(n315) );
  IV U147 ( .A(B[238]), .Z(n495) );
  IV U148 ( .A(B[59]), .Z(n316) );
  IV U149 ( .A(B[60]), .Z(n317) );
  IV U150 ( .A(B[61]), .Z(n318) );
  IV U151 ( .A(B[62]), .Z(n319) );
  IV U152 ( .A(B[63]), .Z(n320) );
  IV U153 ( .A(B[64]), .Z(n321) );
  IV U154 ( .A(B[65]), .Z(n322) );
  IV U155 ( .A(B[66]), .Z(n323) );
  IV U156 ( .A(B[67]), .Z(n324) );
  IV U157 ( .A(B[68]), .Z(n325) );
  IV U158 ( .A(B[239]), .Z(n496) );
  IV U159 ( .A(B[69]), .Z(n326) );
  IV U160 ( .A(B[70]), .Z(n327) );
  IV U161 ( .A(B[71]), .Z(n328) );
  IV U162 ( .A(B[72]), .Z(n329) );
  IV U163 ( .A(B[73]), .Z(n330) );
  IV U164 ( .A(B[74]), .Z(n331) );
  IV U165 ( .A(B[75]), .Z(n332) );
  IV U166 ( .A(B[76]), .Z(n333) );
  IV U167 ( .A(B[77]), .Z(n334) );
  IV U168 ( .A(B[78]), .Z(n335) );
  IV U169 ( .A(B[240]), .Z(n497) );
  IV U170 ( .A(B[79]), .Z(n336) );
  IV U171 ( .A(B[80]), .Z(n337) );
  IV U172 ( .A(B[81]), .Z(n338) );
  IV U173 ( .A(B[82]), .Z(n339) );
  IV U174 ( .A(B[83]), .Z(n340) );
  IV U175 ( .A(B[84]), .Z(n341) );
  IV U176 ( .A(B[85]), .Z(n342) );
  IV U177 ( .A(B[86]), .Z(n343) );
  IV U178 ( .A(B[87]), .Z(n344) );
  IV U179 ( .A(B[88]), .Z(n345) );
  IV U180 ( .A(B[241]), .Z(n498) );
  IV U181 ( .A(B[89]), .Z(n346) );
  IV U182 ( .A(B[90]), .Z(n347) );
  IV U183 ( .A(B[91]), .Z(n348) );
  IV U184 ( .A(B[92]), .Z(n349) );
  IV U185 ( .A(B[93]), .Z(n350) );
  IV U186 ( .A(B[94]), .Z(n351) );
  IV U187 ( .A(B[95]), .Z(n352) );
  IV U188 ( .A(B[96]), .Z(n353) );
  IV U189 ( .A(B[97]), .Z(n354) );
  IV U190 ( .A(B[98]), .Z(n355) );
  IV U191 ( .A(B[242]), .Z(n499) );
  IV U192 ( .A(B[99]), .Z(n356) );
  IV U193 ( .A(B[100]), .Z(n357) );
  IV U194 ( .A(B[101]), .Z(n358) );
  IV U195 ( .A(B[102]), .Z(n359) );
  IV U196 ( .A(B[103]), .Z(n360) );
  IV U197 ( .A(B[104]), .Z(n361) );
  IV U198 ( .A(B[105]), .Z(n362) );
  IV U199 ( .A(B[106]), .Z(n363) );
  IV U200 ( .A(B[107]), .Z(n364) );
  IV U201 ( .A(B[108]), .Z(n365) );
  IV U202 ( .A(B[243]), .Z(n500) );
  IV U203 ( .A(B[109]), .Z(n366) );
  IV U204 ( .A(B[110]), .Z(n367) );
  IV U205 ( .A(B[111]), .Z(n368) );
  IV U206 ( .A(B[112]), .Z(n369) );
  IV U207 ( .A(B[113]), .Z(n370) );
  IV U208 ( .A(B[114]), .Z(n371) );
  IV U209 ( .A(B[115]), .Z(n372) );
  IV U210 ( .A(B[116]), .Z(n373) );
  IV U211 ( .A(B[117]), .Z(n374) );
  IV U212 ( .A(B[118]), .Z(n375) );
  IV U213 ( .A(B[244]), .Z(n501) );
  IV U214 ( .A(B[119]), .Z(n376) );
  IV U215 ( .A(B[120]), .Z(n377) );
  IV U216 ( .A(B[121]), .Z(n378) );
  IV U217 ( .A(B[122]), .Z(n379) );
  IV U218 ( .A(B[123]), .Z(n380) );
  IV U219 ( .A(B[124]), .Z(n381) );
  IV U220 ( .A(B[125]), .Z(n382) );
  IV U221 ( .A(B[126]), .Z(n383) );
  IV U222 ( .A(B[127]), .Z(n384) );
  IV U223 ( .A(B[128]), .Z(n385) );
  IV U224 ( .A(B[245]), .Z(n502) );
  IV U225 ( .A(B[129]), .Z(n386) );
  IV U226 ( .A(B[130]), .Z(n387) );
  IV U227 ( .A(B[131]), .Z(n388) );
  IV U228 ( .A(B[132]), .Z(n389) );
  IV U229 ( .A(B[133]), .Z(n390) );
  IV U230 ( .A(B[134]), .Z(n391) );
  IV U231 ( .A(B[135]), .Z(n392) );
  IV U232 ( .A(B[136]), .Z(n393) );
  IV U233 ( .A(B[137]), .Z(n394) );
  IV U234 ( .A(B[138]), .Z(n395) );
  IV U235 ( .A(B[246]), .Z(n503) );
  IV U236 ( .A(B[139]), .Z(n396) );
  IV U237 ( .A(B[140]), .Z(n397) );
  IV U238 ( .A(B[141]), .Z(n398) );
  IV U239 ( .A(B[142]), .Z(n399) );
  IV U240 ( .A(B[143]), .Z(n400) );
  IV U241 ( .A(B[144]), .Z(n401) );
  IV U242 ( .A(B[145]), .Z(n402) );
  IV U243 ( .A(B[146]), .Z(n403) );
  IV U244 ( .A(B[147]), .Z(n404) );
  IV U245 ( .A(B[148]), .Z(n405) );
  IV U246 ( .A(B[247]), .Z(n504) );
  IV U247 ( .A(B[149]), .Z(n406) );
  IV U248 ( .A(B[150]), .Z(n407) );
  IV U249 ( .A(B[151]), .Z(n408) );
  IV U250 ( .A(B[152]), .Z(n409) );
  IV U251 ( .A(B[153]), .Z(n410) );
  IV U252 ( .A(B[154]), .Z(n411) );
  IV U253 ( .A(B[155]), .Z(n412) );
  IV U254 ( .A(B[156]), .Z(n413) );
  IV U255 ( .A(B[157]), .Z(n414) );
  IV U256 ( .A(B[158]), .Z(n415) );
  IV U257 ( .A(B[248]), .Z(n505) );
endmodule


module modmult_step_N256_1_0 ( xregN_1, y, n, zin, zout );
  input [255:0] y;
  input [255:0] n;
  input [257:0] zin;
  output [257:0] zout;
  input xregN_1;
  wire   c1, c2, n1;
  wire   [257:0] w1;
  wire   [257:0] w2;
  wire   [257:0] w3;
  wire   [257:0] z2;
  wire   [257:0] z3;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6;

  MUX_N258_3 MUX_1 ( .A({1'b0, 1'b0, y}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .S(xregN_1), .O({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, w1[255:0]}) );
  MUX_N258_8 MUX_2 ( .A({1'b0, 1'b0, n}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .S(c1), .O({SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        w2[255:0]}) );
  MUX_N258_7 MUX_3 ( .A({1'b0, 1'b0, n}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .S(n1), .O({SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        w3[255:0]}) );
  ADD_N258_1_0 ADD_1 ( .A({zin[256:0], 1'b0}), .B({1'b0, 1'b0, w1[255:0]}), 
        .CI(1'b0), .S(z2) );
  COMP_N258_2 COMP_1 ( .A(z2), .B({1'b0, 1'b0, n}), .O(c1) );
  SUB_N258_2 SUB_1 ( .A(z2), .B({1'b0, 1'b0, w2[255:0]}), .S(z3) );
  COMP_N258_5 COMP_2 ( .A({1'b0, 1'b0, n}), .B(z3), .O(c2) );
  SUB_N258_5 SUB_2 ( .A({1'b0, z3[256:0]}), .B({1'b0, 1'b0, w3[255:0]}), .S({
        SYNOPSYS_UNCONNECTED__6, zout[256:0]}) );
  IV U2 ( .A(c2), .Z(n1) );
endmodule


module MUX_N258_4 ( A, B, S, O );
  input [257:0] A;
  input [257:0] B;
  output [257:0] O;
  input S;


  ANDN U1 ( .B(A[9]), .A(S), .Z(O[9]) );
  ANDN U2 ( .B(A[99]), .A(S), .Z(O[99]) );
  ANDN U3 ( .B(A[98]), .A(S), .Z(O[98]) );
  ANDN U4 ( .B(A[97]), .A(S), .Z(O[97]) );
  ANDN U5 ( .B(A[96]), .A(S), .Z(O[96]) );
  ANDN U6 ( .B(A[95]), .A(S), .Z(O[95]) );
  ANDN U7 ( .B(A[94]), .A(S), .Z(O[94]) );
  ANDN U8 ( .B(A[93]), .A(S), .Z(O[93]) );
  ANDN U9 ( .B(A[92]), .A(S), .Z(O[92]) );
  ANDN U10 ( .B(A[91]), .A(S), .Z(O[91]) );
  ANDN U11 ( .B(A[90]), .A(S), .Z(O[90]) );
  ANDN U12 ( .B(A[8]), .A(S), .Z(O[8]) );
  ANDN U13 ( .B(A[89]), .A(S), .Z(O[89]) );
  ANDN U14 ( .B(A[88]), .A(S), .Z(O[88]) );
  ANDN U15 ( .B(A[87]), .A(S), .Z(O[87]) );
  ANDN U16 ( .B(A[86]), .A(S), .Z(O[86]) );
  ANDN U17 ( .B(A[85]), .A(S), .Z(O[85]) );
  ANDN U18 ( .B(A[84]), .A(S), .Z(O[84]) );
  ANDN U19 ( .B(A[83]), .A(S), .Z(O[83]) );
  ANDN U20 ( .B(A[82]), .A(S), .Z(O[82]) );
  ANDN U21 ( .B(A[81]), .A(S), .Z(O[81]) );
  ANDN U22 ( .B(A[80]), .A(S), .Z(O[80]) );
  ANDN U23 ( .B(A[7]), .A(S), .Z(O[7]) );
  ANDN U24 ( .B(A[79]), .A(S), .Z(O[79]) );
  ANDN U25 ( .B(A[78]), .A(S), .Z(O[78]) );
  ANDN U26 ( .B(A[77]), .A(S), .Z(O[77]) );
  ANDN U27 ( .B(A[76]), .A(S), .Z(O[76]) );
  ANDN U28 ( .B(A[75]), .A(S), .Z(O[75]) );
  ANDN U29 ( .B(A[74]), .A(S), .Z(O[74]) );
  ANDN U30 ( .B(A[73]), .A(S), .Z(O[73]) );
  ANDN U31 ( .B(A[72]), .A(S), .Z(O[72]) );
  ANDN U32 ( .B(A[71]), .A(S), .Z(O[71]) );
  ANDN U33 ( .B(A[70]), .A(S), .Z(O[70]) );
  ANDN U34 ( .B(A[6]), .A(S), .Z(O[6]) );
  ANDN U35 ( .B(A[69]), .A(S), .Z(O[69]) );
  ANDN U36 ( .B(A[68]), .A(S), .Z(O[68]) );
  ANDN U37 ( .B(A[67]), .A(S), .Z(O[67]) );
  ANDN U38 ( .B(A[66]), .A(S), .Z(O[66]) );
  ANDN U39 ( .B(A[65]), .A(S), .Z(O[65]) );
  ANDN U40 ( .B(A[64]), .A(S), .Z(O[64]) );
  ANDN U41 ( .B(A[63]), .A(S), .Z(O[63]) );
  ANDN U42 ( .B(A[62]), .A(S), .Z(O[62]) );
  ANDN U43 ( .B(A[61]), .A(S), .Z(O[61]) );
  ANDN U44 ( .B(A[60]), .A(S), .Z(O[60]) );
  ANDN U45 ( .B(A[5]), .A(S), .Z(O[5]) );
  ANDN U46 ( .B(A[59]), .A(S), .Z(O[59]) );
  ANDN U47 ( .B(A[58]), .A(S), .Z(O[58]) );
  ANDN U48 ( .B(A[57]), .A(S), .Z(O[57]) );
  ANDN U49 ( .B(A[56]), .A(S), .Z(O[56]) );
  ANDN U50 ( .B(A[55]), .A(S), .Z(O[55]) );
  ANDN U51 ( .B(A[54]), .A(S), .Z(O[54]) );
  ANDN U52 ( .B(A[53]), .A(S), .Z(O[53]) );
  ANDN U53 ( .B(A[52]), .A(S), .Z(O[52]) );
  ANDN U54 ( .B(A[51]), .A(S), .Z(O[51]) );
  ANDN U55 ( .B(A[50]), .A(S), .Z(O[50]) );
  ANDN U56 ( .B(A[4]), .A(S), .Z(O[4]) );
  ANDN U57 ( .B(A[49]), .A(S), .Z(O[49]) );
  ANDN U58 ( .B(A[48]), .A(S), .Z(O[48]) );
  ANDN U59 ( .B(A[47]), .A(S), .Z(O[47]) );
  ANDN U60 ( .B(A[46]), .A(S), .Z(O[46]) );
  ANDN U61 ( .B(A[45]), .A(S), .Z(O[45]) );
  ANDN U62 ( .B(A[44]), .A(S), .Z(O[44]) );
  ANDN U63 ( .B(A[43]), .A(S), .Z(O[43]) );
  ANDN U64 ( .B(A[42]), .A(S), .Z(O[42]) );
  ANDN U65 ( .B(A[41]), .A(S), .Z(O[41]) );
  ANDN U66 ( .B(A[40]), .A(S), .Z(O[40]) );
  ANDN U67 ( .B(A[3]), .A(S), .Z(O[3]) );
  ANDN U68 ( .B(A[39]), .A(S), .Z(O[39]) );
  ANDN U69 ( .B(A[38]), .A(S), .Z(O[38]) );
  ANDN U70 ( .B(A[37]), .A(S), .Z(O[37]) );
  ANDN U71 ( .B(A[36]), .A(S), .Z(O[36]) );
  ANDN U72 ( .B(A[35]), .A(S), .Z(O[35]) );
  ANDN U73 ( .B(A[34]), .A(S), .Z(O[34]) );
  ANDN U74 ( .B(A[33]), .A(S), .Z(O[33]) );
  ANDN U75 ( .B(A[32]), .A(S), .Z(O[32]) );
  ANDN U76 ( .B(A[31]), .A(S), .Z(O[31]) );
  ANDN U77 ( .B(A[30]), .A(S), .Z(O[30]) );
  ANDN U78 ( .B(A[2]), .A(S), .Z(O[2]) );
  ANDN U79 ( .B(A[29]), .A(S), .Z(O[29]) );
  ANDN U80 ( .B(A[28]), .A(S), .Z(O[28]) );
  ANDN U81 ( .B(A[27]), .A(S), .Z(O[27]) );
  ANDN U82 ( .B(A[26]), .A(S), .Z(O[26]) );
  ANDN U83 ( .B(A[25]), .A(S), .Z(O[25]) );
  ANDN U84 ( .B(A[255]), .A(S), .Z(O[255]) );
  ANDN U85 ( .B(A[254]), .A(S), .Z(O[254]) );
  ANDN U86 ( .B(A[253]), .A(S), .Z(O[253]) );
  ANDN U87 ( .B(A[252]), .A(S), .Z(O[252]) );
  ANDN U88 ( .B(A[251]), .A(S), .Z(O[251]) );
  ANDN U89 ( .B(A[250]), .A(S), .Z(O[250]) );
  ANDN U90 ( .B(A[24]), .A(S), .Z(O[24]) );
  ANDN U91 ( .B(A[249]), .A(S), .Z(O[249]) );
  ANDN U92 ( .B(A[248]), .A(S), .Z(O[248]) );
  ANDN U93 ( .B(A[247]), .A(S), .Z(O[247]) );
  ANDN U94 ( .B(A[246]), .A(S), .Z(O[246]) );
  ANDN U95 ( .B(A[245]), .A(S), .Z(O[245]) );
  ANDN U96 ( .B(A[244]), .A(S), .Z(O[244]) );
  ANDN U97 ( .B(A[243]), .A(S), .Z(O[243]) );
  ANDN U98 ( .B(A[242]), .A(S), .Z(O[242]) );
  ANDN U99 ( .B(A[241]), .A(S), .Z(O[241]) );
  ANDN U100 ( .B(A[240]), .A(S), .Z(O[240]) );
  ANDN U101 ( .B(A[23]), .A(S), .Z(O[23]) );
  ANDN U102 ( .B(A[239]), .A(S), .Z(O[239]) );
  ANDN U103 ( .B(A[238]), .A(S), .Z(O[238]) );
  ANDN U104 ( .B(A[237]), .A(S), .Z(O[237]) );
  ANDN U105 ( .B(A[236]), .A(S), .Z(O[236]) );
  ANDN U106 ( .B(A[235]), .A(S), .Z(O[235]) );
  ANDN U107 ( .B(A[234]), .A(S), .Z(O[234]) );
  ANDN U108 ( .B(A[233]), .A(S), .Z(O[233]) );
  ANDN U109 ( .B(A[232]), .A(S), .Z(O[232]) );
  ANDN U110 ( .B(A[231]), .A(S), .Z(O[231]) );
  ANDN U111 ( .B(A[230]), .A(S), .Z(O[230]) );
  ANDN U112 ( .B(A[22]), .A(S), .Z(O[22]) );
  ANDN U113 ( .B(A[229]), .A(S), .Z(O[229]) );
  ANDN U114 ( .B(A[228]), .A(S), .Z(O[228]) );
  ANDN U115 ( .B(A[227]), .A(S), .Z(O[227]) );
  ANDN U116 ( .B(A[226]), .A(S), .Z(O[226]) );
  ANDN U117 ( .B(A[225]), .A(S), .Z(O[225]) );
  ANDN U118 ( .B(A[224]), .A(S), .Z(O[224]) );
  ANDN U119 ( .B(A[223]), .A(S), .Z(O[223]) );
  ANDN U120 ( .B(A[222]), .A(S), .Z(O[222]) );
  ANDN U121 ( .B(A[221]), .A(S), .Z(O[221]) );
  ANDN U122 ( .B(A[220]), .A(S), .Z(O[220]) );
  ANDN U123 ( .B(A[21]), .A(S), .Z(O[21]) );
  ANDN U124 ( .B(A[219]), .A(S), .Z(O[219]) );
  ANDN U125 ( .B(A[218]), .A(S), .Z(O[218]) );
  ANDN U126 ( .B(A[217]), .A(S), .Z(O[217]) );
  ANDN U127 ( .B(A[216]), .A(S), .Z(O[216]) );
  ANDN U128 ( .B(A[215]), .A(S), .Z(O[215]) );
  ANDN U129 ( .B(A[214]), .A(S), .Z(O[214]) );
  ANDN U130 ( .B(A[213]), .A(S), .Z(O[213]) );
  ANDN U131 ( .B(A[212]), .A(S), .Z(O[212]) );
  ANDN U132 ( .B(A[211]), .A(S), .Z(O[211]) );
  ANDN U133 ( .B(A[210]), .A(S), .Z(O[210]) );
  ANDN U134 ( .B(A[20]), .A(S), .Z(O[20]) );
  ANDN U135 ( .B(A[209]), .A(S), .Z(O[209]) );
  ANDN U136 ( .B(A[208]), .A(S), .Z(O[208]) );
  ANDN U137 ( .B(A[207]), .A(S), .Z(O[207]) );
  ANDN U138 ( .B(A[206]), .A(S), .Z(O[206]) );
  ANDN U139 ( .B(A[205]), .A(S), .Z(O[205]) );
  ANDN U140 ( .B(A[204]), .A(S), .Z(O[204]) );
  ANDN U141 ( .B(A[203]), .A(S), .Z(O[203]) );
  ANDN U142 ( .B(A[202]), .A(S), .Z(O[202]) );
  ANDN U143 ( .B(A[201]), .A(S), .Z(O[201]) );
  ANDN U144 ( .B(A[200]), .A(S), .Z(O[200]) );
  ANDN U145 ( .B(A[1]), .A(S), .Z(O[1]) );
  ANDN U146 ( .B(A[19]), .A(S), .Z(O[19]) );
  ANDN U147 ( .B(A[199]), .A(S), .Z(O[199]) );
  ANDN U148 ( .B(A[198]), .A(S), .Z(O[198]) );
  ANDN U149 ( .B(A[197]), .A(S), .Z(O[197]) );
  ANDN U150 ( .B(A[196]), .A(S), .Z(O[196]) );
  ANDN U151 ( .B(A[195]), .A(S), .Z(O[195]) );
  ANDN U152 ( .B(A[194]), .A(S), .Z(O[194]) );
  ANDN U153 ( .B(A[193]), .A(S), .Z(O[193]) );
  ANDN U154 ( .B(A[192]), .A(S), .Z(O[192]) );
  ANDN U155 ( .B(A[191]), .A(S), .Z(O[191]) );
  ANDN U156 ( .B(A[190]), .A(S), .Z(O[190]) );
  ANDN U157 ( .B(A[18]), .A(S), .Z(O[18]) );
  ANDN U158 ( .B(A[189]), .A(S), .Z(O[189]) );
  ANDN U159 ( .B(A[188]), .A(S), .Z(O[188]) );
  ANDN U160 ( .B(A[187]), .A(S), .Z(O[187]) );
  ANDN U161 ( .B(A[186]), .A(S), .Z(O[186]) );
  ANDN U162 ( .B(A[185]), .A(S), .Z(O[185]) );
  ANDN U163 ( .B(A[184]), .A(S), .Z(O[184]) );
  ANDN U164 ( .B(A[183]), .A(S), .Z(O[183]) );
  ANDN U165 ( .B(A[182]), .A(S), .Z(O[182]) );
  ANDN U166 ( .B(A[181]), .A(S), .Z(O[181]) );
  ANDN U167 ( .B(A[180]), .A(S), .Z(O[180]) );
  ANDN U168 ( .B(A[17]), .A(S), .Z(O[17]) );
  ANDN U169 ( .B(A[179]), .A(S), .Z(O[179]) );
  ANDN U170 ( .B(A[178]), .A(S), .Z(O[178]) );
  ANDN U171 ( .B(A[177]), .A(S), .Z(O[177]) );
  ANDN U172 ( .B(A[176]), .A(S), .Z(O[176]) );
  ANDN U173 ( .B(A[175]), .A(S), .Z(O[175]) );
  ANDN U174 ( .B(A[174]), .A(S), .Z(O[174]) );
  ANDN U175 ( .B(A[173]), .A(S), .Z(O[173]) );
  ANDN U176 ( .B(A[172]), .A(S), .Z(O[172]) );
  ANDN U177 ( .B(A[171]), .A(S), .Z(O[171]) );
  ANDN U178 ( .B(A[170]), .A(S), .Z(O[170]) );
  ANDN U179 ( .B(A[16]), .A(S), .Z(O[16]) );
  ANDN U180 ( .B(A[169]), .A(S), .Z(O[169]) );
  ANDN U181 ( .B(A[168]), .A(S), .Z(O[168]) );
  ANDN U182 ( .B(A[167]), .A(S), .Z(O[167]) );
  ANDN U183 ( .B(A[166]), .A(S), .Z(O[166]) );
  ANDN U184 ( .B(A[165]), .A(S), .Z(O[165]) );
  ANDN U185 ( .B(A[164]), .A(S), .Z(O[164]) );
  ANDN U186 ( .B(A[163]), .A(S), .Z(O[163]) );
  ANDN U187 ( .B(A[162]), .A(S), .Z(O[162]) );
  ANDN U188 ( .B(A[161]), .A(S), .Z(O[161]) );
  ANDN U189 ( .B(A[160]), .A(S), .Z(O[160]) );
  ANDN U190 ( .B(A[15]), .A(S), .Z(O[15]) );
  ANDN U191 ( .B(A[159]), .A(S), .Z(O[159]) );
  ANDN U192 ( .B(A[158]), .A(S), .Z(O[158]) );
  ANDN U193 ( .B(A[157]), .A(S), .Z(O[157]) );
  ANDN U194 ( .B(A[156]), .A(S), .Z(O[156]) );
  ANDN U195 ( .B(A[155]), .A(S), .Z(O[155]) );
  ANDN U196 ( .B(A[154]), .A(S), .Z(O[154]) );
  ANDN U197 ( .B(A[153]), .A(S), .Z(O[153]) );
  ANDN U198 ( .B(A[152]), .A(S), .Z(O[152]) );
  ANDN U199 ( .B(A[151]), .A(S), .Z(O[151]) );
  ANDN U200 ( .B(A[150]), .A(S), .Z(O[150]) );
  ANDN U201 ( .B(A[14]), .A(S), .Z(O[14]) );
  ANDN U202 ( .B(A[149]), .A(S), .Z(O[149]) );
  ANDN U203 ( .B(A[148]), .A(S), .Z(O[148]) );
  ANDN U204 ( .B(A[147]), .A(S), .Z(O[147]) );
  ANDN U205 ( .B(A[146]), .A(S), .Z(O[146]) );
  ANDN U206 ( .B(A[145]), .A(S), .Z(O[145]) );
  ANDN U207 ( .B(A[144]), .A(S), .Z(O[144]) );
  ANDN U208 ( .B(A[143]), .A(S), .Z(O[143]) );
  ANDN U209 ( .B(A[142]), .A(S), .Z(O[142]) );
  ANDN U210 ( .B(A[141]), .A(S), .Z(O[141]) );
  ANDN U211 ( .B(A[140]), .A(S), .Z(O[140]) );
  ANDN U212 ( .B(A[13]), .A(S), .Z(O[13]) );
  ANDN U213 ( .B(A[139]), .A(S), .Z(O[139]) );
  ANDN U214 ( .B(A[138]), .A(S), .Z(O[138]) );
  ANDN U215 ( .B(A[137]), .A(S), .Z(O[137]) );
  ANDN U216 ( .B(A[136]), .A(S), .Z(O[136]) );
  ANDN U217 ( .B(A[135]), .A(S), .Z(O[135]) );
  ANDN U218 ( .B(A[134]), .A(S), .Z(O[134]) );
  ANDN U219 ( .B(A[133]), .A(S), .Z(O[133]) );
  ANDN U220 ( .B(A[132]), .A(S), .Z(O[132]) );
  ANDN U221 ( .B(A[131]), .A(S), .Z(O[131]) );
  ANDN U222 ( .B(A[130]), .A(S), .Z(O[130]) );
  ANDN U223 ( .B(A[12]), .A(S), .Z(O[12]) );
  ANDN U224 ( .B(A[129]), .A(S), .Z(O[129]) );
  ANDN U225 ( .B(A[128]), .A(S), .Z(O[128]) );
  ANDN U226 ( .B(A[127]), .A(S), .Z(O[127]) );
  ANDN U227 ( .B(A[126]), .A(S), .Z(O[126]) );
  ANDN U228 ( .B(A[125]), .A(S), .Z(O[125]) );
  ANDN U229 ( .B(A[124]), .A(S), .Z(O[124]) );
  ANDN U230 ( .B(A[123]), .A(S), .Z(O[123]) );
  ANDN U231 ( .B(A[122]), .A(S), .Z(O[122]) );
  ANDN U232 ( .B(A[121]), .A(S), .Z(O[121]) );
  ANDN U233 ( .B(A[120]), .A(S), .Z(O[120]) );
  ANDN U234 ( .B(A[11]), .A(S), .Z(O[11]) );
  ANDN U235 ( .B(A[119]), .A(S), .Z(O[119]) );
  ANDN U236 ( .B(A[118]), .A(S), .Z(O[118]) );
  ANDN U237 ( .B(A[117]), .A(S), .Z(O[117]) );
  ANDN U238 ( .B(A[116]), .A(S), .Z(O[116]) );
  ANDN U239 ( .B(A[115]), .A(S), .Z(O[115]) );
  ANDN U240 ( .B(A[114]), .A(S), .Z(O[114]) );
  ANDN U241 ( .B(A[113]), .A(S), .Z(O[113]) );
  ANDN U242 ( .B(A[112]), .A(S), .Z(O[112]) );
  ANDN U243 ( .B(A[111]), .A(S), .Z(O[111]) );
  ANDN U244 ( .B(A[110]), .A(S), .Z(O[110]) );
  ANDN U245 ( .B(A[10]), .A(S), .Z(O[10]) );
  ANDN U246 ( .B(A[109]), .A(S), .Z(O[109]) );
  ANDN U247 ( .B(A[108]), .A(S), .Z(O[108]) );
  ANDN U248 ( .B(A[107]), .A(S), .Z(O[107]) );
  ANDN U249 ( .B(A[106]), .A(S), .Z(O[106]) );
  ANDN U250 ( .B(A[105]), .A(S), .Z(O[105]) );
  ANDN U251 ( .B(A[104]), .A(S), .Z(O[104]) );
  ANDN U252 ( .B(A[103]), .A(S), .Z(O[103]) );
  ANDN U253 ( .B(A[102]), .A(S), .Z(O[102]) );
  ANDN U254 ( .B(A[101]), .A(S), .Z(O[101]) );
  ANDN U255 ( .B(A[100]), .A(S), .Z(O[100]) );
  ANDN U256 ( .B(A[0]), .A(S), .Z(O[0]) );
endmodule


module MUX_N258_5 ( A, B, S, O );
  input [257:0] A;
  input [257:0] B;
  output [257:0] O;
  input S;


  ANDN U1 ( .B(A[9]), .A(S), .Z(O[9]) );
  ANDN U2 ( .B(A[99]), .A(S), .Z(O[99]) );
  ANDN U3 ( .B(A[98]), .A(S), .Z(O[98]) );
  ANDN U4 ( .B(A[97]), .A(S), .Z(O[97]) );
  ANDN U5 ( .B(A[96]), .A(S), .Z(O[96]) );
  ANDN U6 ( .B(A[95]), .A(S), .Z(O[95]) );
  ANDN U7 ( .B(A[94]), .A(S), .Z(O[94]) );
  ANDN U8 ( .B(A[93]), .A(S), .Z(O[93]) );
  ANDN U9 ( .B(A[92]), .A(S), .Z(O[92]) );
  ANDN U10 ( .B(A[91]), .A(S), .Z(O[91]) );
  ANDN U11 ( .B(A[90]), .A(S), .Z(O[90]) );
  ANDN U12 ( .B(A[8]), .A(S), .Z(O[8]) );
  ANDN U13 ( .B(A[89]), .A(S), .Z(O[89]) );
  ANDN U14 ( .B(A[88]), .A(S), .Z(O[88]) );
  ANDN U15 ( .B(A[87]), .A(S), .Z(O[87]) );
  ANDN U16 ( .B(A[86]), .A(S), .Z(O[86]) );
  ANDN U17 ( .B(A[85]), .A(S), .Z(O[85]) );
  ANDN U18 ( .B(A[84]), .A(S), .Z(O[84]) );
  ANDN U19 ( .B(A[83]), .A(S), .Z(O[83]) );
  ANDN U20 ( .B(A[82]), .A(S), .Z(O[82]) );
  ANDN U21 ( .B(A[81]), .A(S), .Z(O[81]) );
  ANDN U22 ( .B(A[80]), .A(S), .Z(O[80]) );
  ANDN U23 ( .B(A[7]), .A(S), .Z(O[7]) );
  ANDN U24 ( .B(A[79]), .A(S), .Z(O[79]) );
  ANDN U25 ( .B(A[78]), .A(S), .Z(O[78]) );
  ANDN U26 ( .B(A[77]), .A(S), .Z(O[77]) );
  ANDN U27 ( .B(A[76]), .A(S), .Z(O[76]) );
  ANDN U28 ( .B(A[75]), .A(S), .Z(O[75]) );
  ANDN U29 ( .B(A[74]), .A(S), .Z(O[74]) );
  ANDN U30 ( .B(A[73]), .A(S), .Z(O[73]) );
  ANDN U31 ( .B(A[72]), .A(S), .Z(O[72]) );
  ANDN U32 ( .B(A[71]), .A(S), .Z(O[71]) );
  ANDN U33 ( .B(A[70]), .A(S), .Z(O[70]) );
  ANDN U34 ( .B(A[6]), .A(S), .Z(O[6]) );
  ANDN U35 ( .B(A[69]), .A(S), .Z(O[69]) );
  ANDN U36 ( .B(A[68]), .A(S), .Z(O[68]) );
  ANDN U37 ( .B(A[67]), .A(S), .Z(O[67]) );
  ANDN U38 ( .B(A[66]), .A(S), .Z(O[66]) );
  ANDN U39 ( .B(A[65]), .A(S), .Z(O[65]) );
  ANDN U40 ( .B(A[64]), .A(S), .Z(O[64]) );
  ANDN U41 ( .B(A[63]), .A(S), .Z(O[63]) );
  ANDN U42 ( .B(A[62]), .A(S), .Z(O[62]) );
  ANDN U43 ( .B(A[61]), .A(S), .Z(O[61]) );
  ANDN U44 ( .B(A[60]), .A(S), .Z(O[60]) );
  ANDN U45 ( .B(A[5]), .A(S), .Z(O[5]) );
  ANDN U46 ( .B(A[59]), .A(S), .Z(O[59]) );
  ANDN U47 ( .B(A[58]), .A(S), .Z(O[58]) );
  ANDN U48 ( .B(A[57]), .A(S), .Z(O[57]) );
  ANDN U49 ( .B(A[56]), .A(S), .Z(O[56]) );
  ANDN U50 ( .B(A[55]), .A(S), .Z(O[55]) );
  ANDN U51 ( .B(A[54]), .A(S), .Z(O[54]) );
  ANDN U52 ( .B(A[53]), .A(S), .Z(O[53]) );
  ANDN U53 ( .B(A[52]), .A(S), .Z(O[52]) );
  ANDN U54 ( .B(A[51]), .A(S), .Z(O[51]) );
  ANDN U55 ( .B(A[50]), .A(S), .Z(O[50]) );
  ANDN U56 ( .B(A[4]), .A(S), .Z(O[4]) );
  ANDN U57 ( .B(A[49]), .A(S), .Z(O[49]) );
  ANDN U58 ( .B(A[48]), .A(S), .Z(O[48]) );
  ANDN U59 ( .B(A[47]), .A(S), .Z(O[47]) );
  ANDN U60 ( .B(A[46]), .A(S), .Z(O[46]) );
  ANDN U61 ( .B(A[45]), .A(S), .Z(O[45]) );
  ANDN U62 ( .B(A[44]), .A(S), .Z(O[44]) );
  ANDN U63 ( .B(A[43]), .A(S), .Z(O[43]) );
  ANDN U64 ( .B(A[42]), .A(S), .Z(O[42]) );
  ANDN U65 ( .B(A[41]), .A(S), .Z(O[41]) );
  ANDN U66 ( .B(A[40]), .A(S), .Z(O[40]) );
  ANDN U67 ( .B(A[3]), .A(S), .Z(O[3]) );
  ANDN U68 ( .B(A[39]), .A(S), .Z(O[39]) );
  ANDN U69 ( .B(A[38]), .A(S), .Z(O[38]) );
  ANDN U70 ( .B(A[37]), .A(S), .Z(O[37]) );
  ANDN U71 ( .B(A[36]), .A(S), .Z(O[36]) );
  ANDN U72 ( .B(A[35]), .A(S), .Z(O[35]) );
  ANDN U73 ( .B(A[34]), .A(S), .Z(O[34]) );
  ANDN U74 ( .B(A[33]), .A(S), .Z(O[33]) );
  ANDN U75 ( .B(A[32]), .A(S), .Z(O[32]) );
  ANDN U76 ( .B(A[31]), .A(S), .Z(O[31]) );
  ANDN U77 ( .B(A[30]), .A(S), .Z(O[30]) );
  ANDN U78 ( .B(A[2]), .A(S), .Z(O[2]) );
  ANDN U79 ( .B(A[29]), .A(S), .Z(O[29]) );
  ANDN U80 ( .B(A[28]), .A(S), .Z(O[28]) );
  ANDN U81 ( .B(A[27]), .A(S), .Z(O[27]) );
  ANDN U82 ( .B(A[26]), .A(S), .Z(O[26]) );
  ANDN U83 ( .B(A[25]), .A(S), .Z(O[25]) );
  ANDN U84 ( .B(A[255]), .A(S), .Z(O[255]) );
  ANDN U85 ( .B(A[254]), .A(S), .Z(O[254]) );
  ANDN U86 ( .B(A[253]), .A(S), .Z(O[253]) );
  ANDN U87 ( .B(A[252]), .A(S), .Z(O[252]) );
  ANDN U88 ( .B(A[251]), .A(S), .Z(O[251]) );
  ANDN U89 ( .B(A[250]), .A(S), .Z(O[250]) );
  ANDN U90 ( .B(A[24]), .A(S), .Z(O[24]) );
  ANDN U91 ( .B(A[249]), .A(S), .Z(O[249]) );
  ANDN U92 ( .B(A[248]), .A(S), .Z(O[248]) );
  ANDN U93 ( .B(A[247]), .A(S), .Z(O[247]) );
  ANDN U94 ( .B(A[246]), .A(S), .Z(O[246]) );
  ANDN U95 ( .B(A[245]), .A(S), .Z(O[245]) );
  ANDN U96 ( .B(A[244]), .A(S), .Z(O[244]) );
  ANDN U97 ( .B(A[243]), .A(S), .Z(O[243]) );
  ANDN U98 ( .B(A[242]), .A(S), .Z(O[242]) );
  ANDN U99 ( .B(A[241]), .A(S), .Z(O[241]) );
  ANDN U100 ( .B(A[240]), .A(S), .Z(O[240]) );
  ANDN U101 ( .B(A[23]), .A(S), .Z(O[23]) );
  ANDN U102 ( .B(A[239]), .A(S), .Z(O[239]) );
  ANDN U103 ( .B(A[238]), .A(S), .Z(O[238]) );
  ANDN U104 ( .B(A[237]), .A(S), .Z(O[237]) );
  ANDN U105 ( .B(A[236]), .A(S), .Z(O[236]) );
  ANDN U106 ( .B(A[235]), .A(S), .Z(O[235]) );
  ANDN U107 ( .B(A[234]), .A(S), .Z(O[234]) );
  ANDN U108 ( .B(A[233]), .A(S), .Z(O[233]) );
  ANDN U109 ( .B(A[232]), .A(S), .Z(O[232]) );
  ANDN U110 ( .B(A[231]), .A(S), .Z(O[231]) );
  ANDN U111 ( .B(A[230]), .A(S), .Z(O[230]) );
  ANDN U112 ( .B(A[22]), .A(S), .Z(O[22]) );
  ANDN U113 ( .B(A[229]), .A(S), .Z(O[229]) );
  ANDN U114 ( .B(A[228]), .A(S), .Z(O[228]) );
  ANDN U115 ( .B(A[227]), .A(S), .Z(O[227]) );
  ANDN U116 ( .B(A[226]), .A(S), .Z(O[226]) );
  ANDN U117 ( .B(A[225]), .A(S), .Z(O[225]) );
  ANDN U118 ( .B(A[224]), .A(S), .Z(O[224]) );
  ANDN U119 ( .B(A[223]), .A(S), .Z(O[223]) );
  ANDN U120 ( .B(A[222]), .A(S), .Z(O[222]) );
  ANDN U121 ( .B(A[221]), .A(S), .Z(O[221]) );
  ANDN U122 ( .B(A[220]), .A(S), .Z(O[220]) );
  ANDN U123 ( .B(A[21]), .A(S), .Z(O[21]) );
  ANDN U124 ( .B(A[219]), .A(S), .Z(O[219]) );
  ANDN U125 ( .B(A[218]), .A(S), .Z(O[218]) );
  ANDN U126 ( .B(A[217]), .A(S), .Z(O[217]) );
  ANDN U127 ( .B(A[216]), .A(S), .Z(O[216]) );
  ANDN U128 ( .B(A[215]), .A(S), .Z(O[215]) );
  ANDN U129 ( .B(A[214]), .A(S), .Z(O[214]) );
  ANDN U130 ( .B(A[213]), .A(S), .Z(O[213]) );
  ANDN U131 ( .B(A[212]), .A(S), .Z(O[212]) );
  ANDN U132 ( .B(A[211]), .A(S), .Z(O[211]) );
  ANDN U133 ( .B(A[210]), .A(S), .Z(O[210]) );
  ANDN U134 ( .B(A[20]), .A(S), .Z(O[20]) );
  ANDN U135 ( .B(A[209]), .A(S), .Z(O[209]) );
  ANDN U136 ( .B(A[208]), .A(S), .Z(O[208]) );
  ANDN U137 ( .B(A[207]), .A(S), .Z(O[207]) );
  ANDN U138 ( .B(A[206]), .A(S), .Z(O[206]) );
  ANDN U139 ( .B(A[205]), .A(S), .Z(O[205]) );
  ANDN U140 ( .B(A[204]), .A(S), .Z(O[204]) );
  ANDN U141 ( .B(A[203]), .A(S), .Z(O[203]) );
  ANDN U142 ( .B(A[202]), .A(S), .Z(O[202]) );
  ANDN U143 ( .B(A[201]), .A(S), .Z(O[201]) );
  ANDN U144 ( .B(A[200]), .A(S), .Z(O[200]) );
  ANDN U145 ( .B(A[1]), .A(S), .Z(O[1]) );
  ANDN U146 ( .B(A[19]), .A(S), .Z(O[19]) );
  ANDN U147 ( .B(A[199]), .A(S), .Z(O[199]) );
  ANDN U148 ( .B(A[198]), .A(S), .Z(O[198]) );
  ANDN U149 ( .B(A[197]), .A(S), .Z(O[197]) );
  ANDN U150 ( .B(A[196]), .A(S), .Z(O[196]) );
  ANDN U151 ( .B(A[195]), .A(S), .Z(O[195]) );
  ANDN U152 ( .B(A[194]), .A(S), .Z(O[194]) );
  ANDN U153 ( .B(A[193]), .A(S), .Z(O[193]) );
  ANDN U154 ( .B(A[192]), .A(S), .Z(O[192]) );
  ANDN U155 ( .B(A[191]), .A(S), .Z(O[191]) );
  ANDN U156 ( .B(A[190]), .A(S), .Z(O[190]) );
  ANDN U157 ( .B(A[18]), .A(S), .Z(O[18]) );
  ANDN U158 ( .B(A[189]), .A(S), .Z(O[189]) );
  ANDN U159 ( .B(A[188]), .A(S), .Z(O[188]) );
  ANDN U160 ( .B(A[187]), .A(S), .Z(O[187]) );
  ANDN U161 ( .B(A[186]), .A(S), .Z(O[186]) );
  ANDN U162 ( .B(A[185]), .A(S), .Z(O[185]) );
  ANDN U163 ( .B(A[184]), .A(S), .Z(O[184]) );
  ANDN U164 ( .B(A[183]), .A(S), .Z(O[183]) );
  ANDN U165 ( .B(A[182]), .A(S), .Z(O[182]) );
  ANDN U166 ( .B(A[181]), .A(S), .Z(O[181]) );
  ANDN U167 ( .B(A[180]), .A(S), .Z(O[180]) );
  ANDN U168 ( .B(A[17]), .A(S), .Z(O[17]) );
  ANDN U169 ( .B(A[179]), .A(S), .Z(O[179]) );
  ANDN U170 ( .B(A[178]), .A(S), .Z(O[178]) );
  ANDN U171 ( .B(A[177]), .A(S), .Z(O[177]) );
  ANDN U172 ( .B(A[176]), .A(S), .Z(O[176]) );
  ANDN U173 ( .B(A[175]), .A(S), .Z(O[175]) );
  ANDN U174 ( .B(A[174]), .A(S), .Z(O[174]) );
  ANDN U175 ( .B(A[173]), .A(S), .Z(O[173]) );
  ANDN U176 ( .B(A[172]), .A(S), .Z(O[172]) );
  ANDN U177 ( .B(A[171]), .A(S), .Z(O[171]) );
  ANDN U178 ( .B(A[170]), .A(S), .Z(O[170]) );
  ANDN U179 ( .B(A[16]), .A(S), .Z(O[16]) );
  ANDN U180 ( .B(A[169]), .A(S), .Z(O[169]) );
  ANDN U181 ( .B(A[168]), .A(S), .Z(O[168]) );
  ANDN U182 ( .B(A[167]), .A(S), .Z(O[167]) );
  ANDN U183 ( .B(A[166]), .A(S), .Z(O[166]) );
  ANDN U184 ( .B(A[165]), .A(S), .Z(O[165]) );
  ANDN U185 ( .B(A[164]), .A(S), .Z(O[164]) );
  ANDN U186 ( .B(A[163]), .A(S), .Z(O[163]) );
  ANDN U187 ( .B(A[162]), .A(S), .Z(O[162]) );
  ANDN U188 ( .B(A[161]), .A(S), .Z(O[161]) );
  ANDN U189 ( .B(A[160]), .A(S), .Z(O[160]) );
  ANDN U190 ( .B(A[15]), .A(S), .Z(O[15]) );
  ANDN U191 ( .B(A[159]), .A(S), .Z(O[159]) );
  ANDN U192 ( .B(A[158]), .A(S), .Z(O[158]) );
  ANDN U193 ( .B(A[157]), .A(S), .Z(O[157]) );
  ANDN U194 ( .B(A[156]), .A(S), .Z(O[156]) );
  ANDN U195 ( .B(A[155]), .A(S), .Z(O[155]) );
  ANDN U196 ( .B(A[154]), .A(S), .Z(O[154]) );
  ANDN U197 ( .B(A[153]), .A(S), .Z(O[153]) );
  ANDN U198 ( .B(A[152]), .A(S), .Z(O[152]) );
  ANDN U199 ( .B(A[151]), .A(S), .Z(O[151]) );
  ANDN U200 ( .B(A[150]), .A(S), .Z(O[150]) );
  ANDN U201 ( .B(A[14]), .A(S), .Z(O[14]) );
  ANDN U202 ( .B(A[149]), .A(S), .Z(O[149]) );
  ANDN U203 ( .B(A[148]), .A(S), .Z(O[148]) );
  ANDN U204 ( .B(A[147]), .A(S), .Z(O[147]) );
  ANDN U205 ( .B(A[146]), .A(S), .Z(O[146]) );
  ANDN U206 ( .B(A[145]), .A(S), .Z(O[145]) );
  ANDN U207 ( .B(A[144]), .A(S), .Z(O[144]) );
  ANDN U208 ( .B(A[143]), .A(S), .Z(O[143]) );
  ANDN U209 ( .B(A[142]), .A(S), .Z(O[142]) );
  ANDN U210 ( .B(A[141]), .A(S), .Z(O[141]) );
  ANDN U211 ( .B(A[140]), .A(S), .Z(O[140]) );
  ANDN U212 ( .B(A[13]), .A(S), .Z(O[13]) );
  ANDN U213 ( .B(A[139]), .A(S), .Z(O[139]) );
  ANDN U214 ( .B(A[138]), .A(S), .Z(O[138]) );
  ANDN U215 ( .B(A[137]), .A(S), .Z(O[137]) );
  ANDN U216 ( .B(A[136]), .A(S), .Z(O[136]) );
  ANDN U217 ( .B(A[135]), .A(S), .Z(O[135]) );
  ANDN U218 ( .B(A[134]), .A(S), .Z(O[134]) );
  ANDN U219 ( .B(A[133]), .A(S), .Z(O[133]) );
  ANDN U220 ( .B(A[132]), .A(S), .Z(O[132]) );
  ANDN U221 ( .B(A[131]), .A(S), .Z(O[131]) );
  ANDN U222 ( .B(A[130]), .A(S), .Z(O[130]) );
  ANDN U223 ( .B(A[12]), .A(S), .Z(O[12]) );
  ANDN U224 ( .B(A[129]), .A(S), .Z(O[129]) );
  ANDN U225 ( .B(A[128]), .A(S), .Z(O[128]) );
  ANDN U226 ( .B(A[127]), .A(S), .Z(O[127]) );
  ANDN U227 ( .B(A[126]), .A(S), .Z(O[126]) );
  ANDN U228 ( .B(A[125]), .A(S), .Z(O[125]) );
  ANDN U229 ( .B(A[124]), .A(S), .Z(O[124]) );
  ANDN U230 ( .B(A[123]), .A(S), .Z(O[123]) );
  ANDN U231 ( .B(A[122]), .A(S), .Z(O[122]) );
  ANDN U232 ( .B(A[121]), .A(S), .Z(O[121]) );
  ANDN U233 ( .B(A[120]), .A(S), .Z(O[120]) );
  ANDN U234 ( .B(A[11]), .A(S), .Z(O[11]) );
  ANDN U235 ( .B(A[119]), .A(S), .Z(O[119]) );
  ANDN U236 ( .B(A[118]), .A(S), .Z(O[118]) );
  ANDN U237 ( .B(A[117]), .A(S), .Z(O[117]) );
  ANDN U238 ( .B(A[116]), .A(S), .Z(O[116]) );
  ANDN U239 ( .B(A[115]), .A(S), .Z(O[115]) );
  ANDN U240 ( .B(A[114]), .A(S), .Z(O[114]) );
  ANDN U241 ( .B(A[113]), .A(S), .Z(O[113]) );
  ANDN U242 ( .B(A[112]), .A(S), .Z(O[112]) );
  ANDN U243 ( .B(A[111]), .A(S), .Z(O[111]) );
  ANDN U244 ( .B(A[110]), .A(S), .Z(O[110]) );
  ANDN U245 ( .B(A[10]), .A(S), .Z(O[10]) );
  ANDN U246 ( .B(A[109]), .A(S), .Z(O[109]) );
  ANDN U247 ( .B(A[108]), .A(S), .Z(O[108]) );
  ANDN U248 ( .B(A[107]), .A(S), .Z(O[107]) );
  ANDN U249 ( .B(A[106]), .A(S), .Z(O[106]) );
  ANDN U250 ( .B(A[105]), .A(S), .Z(O[105]) );
  ANDN U251 ( .B(A[104]), .A(S), .Z(O[104]) );
  ANDN U252 ( .B(A[103]), .A(S), .Z(O[103]) );
  ANDN U253 ( .B(A[102]), .A(S), .Z(O[102]) );
  ANDN U254 ( .B(A[101]), .A(S), .Z(O[101]) );
  ANDN U255 ( .B(A[100]), .A(S), .Z(O[100]) );
  ANDN U256 ( .B(A[0]), .A(S), .Z(O[0]) );
endmodule


module MUX_N258_6 ( A, B, S, O );
  input [257:0] A;
  input [257:0] B;
  output [257:0] O;
  input S;


  ANDN U1 ( .B(A[9]), .A(S), .Z(O[9]) );
  ANDN U2 ( .B(A[99]), .A(S), .Z(O[99]) );
  ANDN U3 ( .B(A[98]), .A(S), .Z(O[98]) );
  ANDN U4 ( .B(A[97]), .A(S), .Z(O[97]) );
  ANDN U5 ( .B(A[96]), .A(S), .Z(O[96]) );
  ANDN U6 ( .B(A[95]), .A(S), .Z(O[95]) );
  ANDN U7 ( .B(A[94]), .A(S), .Z(O[94]) );
  ANDN U8 ( .B(A[93]), .A(S), .Z(O[93]) );
  ANDN U9 ( .B(A[92]), .A(S), .Z(O[92]) );
  ANDN U10 ( .B(A[91]), .A(S), .Z(O[91]) );
  ANDN U11 ( .B(A[90]), .A(S), .Z(O[90]) );
  ANDN U12 ( .B(A[8]), .A(S), .Z(O[8]) );
  ANDN U13 ( .B(A[89]), .A(S), .Z(O[89]) );
  ANDN U14 ( .B(A[88]), .A(S), .Z(O[88]) );
  ANDN U15 ( .B(A[87]), .A(S), .Z(O[87]) );
  ANDN U16 ( .B(A[86]), .A(S), .Z(O[86]) );
  ANDN U17 ( .B(A[85]), .A(S), .Z(O[85]) );
  ANDN U18 ( .B(A[84]), .A(S), .Z(O[84]) );
  ANDN U19 ( .B(A[83]), .A(S), .Z(O[83]) );
  ANDN U20 ( .B(A[82]), .A(S), .Z(O[82]) );
  ANDN U21 ( .B(A[81]), .A(S), .Z(O[81]) );
  ANDN U22 ( .B(A[80]), .A(S), .Z(O[80]) );
  ANDN U23 ( .B(A[7]), .A(S), .Z(O[7]) );
  ANDN U24 ( .B(A[79]), .A(S), .Z(O[79]) );
  ANDN U25 ( .B(A[78]), .A(S), .Z(O[78]) );
  ANDN U26 ( .B(A[77]), .A(S), .Z(O[77]) );
  ANDN U27 ( .B(A[76]), .A(S), .Z(O[76]) );
  ANDN U28 ( .B(A[75]), .A(S), .Z(O[75]) );
  ANDN U29 ( .B(A[74]), .A(S), .Z(O[74]) );
  ANDN U30 ( .B(A[73]), .A(S), .Z(O[73]) );
  ANDN U31 ( .B(A[72]), .A(S), .Z(O[72]) );
  ANDN U32 ( .B(A[71]), .A(S), .Z(O[71]) );
  ANDN U33 ( .B(A[70]), .A(S), .Z(O[70]) );
  ANDN U34 ( .B(A[6]), .A(S), .Z(O[6]) );
  ANDN U35 ( .B(A[69]), .A(S), .Z(O[69]) );
  ANDN U36 ( .B(A[68]), .A(S), .Z(O[68]) );
  ANDN U37 ( .B(A[67]), .A(S), .Z(O[67]) );
  ANDN U38 ( .B(A[66]), .A(S), .Z(O[66]) );
  ANDN U39 ( .B(A[65]), .A(S), .Z(O[65]) );
  ANDN U40 ( .B(A[64]), .A(S), .Z(O[64]) );
  ANDN U41 ( .B(A[63]), .A(S), .Z(O[63]) );
  ANDN U42 ( .B(A[62]), .A(S), .Z(O[62]) );
  ANDN U43 ( .B(A[61]), .A(S), .Z(O[61]) );
  ANDN U44 ( .B(A[60]), .A(S), .Z(O[60]) );
  ANDN U45 ( .B(A[5]), .A(S), .Z(O[5]) );
  ANDN U46 ( .B(A[59]), .A(S), .Z(O[59]) );
  ANDN U47 ( .B(A[58]), .A(S), .Z(O[58]) );
  ANDN U48 ( .B(A[57]), .A(S), .Z(O[57]) );
  ANDN U49 ( .B(A[56]), .A(S), .Z(O[56]) );
  ANDN U50 ( .B(A[55]), .A(S), .Z(O[55]) );
  ANDN U51 ( .B(A[54]), .A(S), .Z(O[54]) );
  ANDN U52 ( .B(A[53]), .A(S), .Z(O[53]) );
  ANDN U53 ( .B(A[52]), .A(S), .Z(O[52]) );
  ANDN U54 ( .B(A[51]), .A(S), .Z(O[51]) );
  ANDN U55 ( .B(A[50]), .A(S), .Z(O[50]) );
  ANDN U56 ( .B(A[4]), .A(S), .Z(O[4]) );
  ANDN U57 ( .B(A[49]), .A(S), .Z(O[49]) );
  ANDN U58 ( .B(A[48]), .A(S), .Z(O[48]) );
  ANDN U59 ( .B(A[47]), .A(S), .Z(O[47]) );
  ANDN U60 ( .B(A[46]), .A(S), .Z(O[46]) );
  ANDN U61 ( .B(A[45]), .A(S), .Z(O[45]) );
  ANDN U62 ( .B(A[44]), .A(S), .Z(O[44]) );
  ANDN U63 ( .B(A[43]), .A(S), .Z(O[43]) );
  ANDN U64 ( .B(A[42]), .A(S), .Z(O[42]) );
  ANDN U65 ( .B(A[41]), .A(S), .Z(O[41]) );
  ANDN U66 ( .B(A[40]), .A(S), .Z(O[40]) );
  ANDN U67 ( .B(A[3]), .A(S), .Z(O[3]) );
  ANDN U68 ( .B(A[39]), .A(S), .Z(O[39]) );
  ANDN U69 ( .B(A[38]), .A(S), .Z(O[38]) );
  ANDN U70 ( .B(A[37]), .A(S), .Z(O[37]) );
  ANDN U71 ( .B(A[36]), .A(S), .Z(O[36]) );
  ANDN U72 ( .B(A[35]), .A(S), .Z(O[35]) );
  ANDN U73 ( .B(A[34]), .A(S), .Z(O[34]) );
  ANDN U74 ( .B(A[33]), .A(S), .Z(O[33]) );
  ANDN U75 ( .B(A[32]), .A(S), .Z(O[32]) );
  ANDN U76 ( .B(A[31]), .A(S), .Z(O[31]) );
  ANDN U77 ( .B(A[30]), .A(S), .Z(O[30]) );
  ANDN U78 ( .B(A[2]), .A(S), .Z(O[2]) );
  ANDN U79 ( .B(A[29]), .A(S), .Z(O[29]) );
  ANDN U80 ( .B(A[28]), .A(S), .Z(O[28]) );
  ANDN U81 ( .B(A[27]), .A(S), .Z(O[27]) );
  ANDN U82 ( .B(A[26]), .A(S), .Z(O[26]) );
  ANDN U83 ( .B(A[25]), .A(S), .Z(O[25]) );
  ANDN U84 ( .B(A[255]), .A(S), .Z(O[255]) );
  ANDN U85 ( .B(A[254]), .A(S), .Z(O[254]) );
  ANDN U86 ( .B(A[253]), .A(S), .Z(O[253]) );
  ANDN U87 ( .B(A[252]), .A(S), .Z(O[252]) );
  ANDN U88 ( .B(A[251]), .A(S), .Z(O[251]) );
  ANDN U89 ( .B(A[250]), .A(S), .Z(O[250]) );
  ANDN U90 ( .B(A[24]), .A(S), .Z(O[24]) );
  ANDN U91 ( .B(A[249]), .A(S), .Z(O[249]) );
  ANDN U92 ( .B(A[248]), .A(S), .Z(O[248]) );
  ANDN U93 ( .B(A[247]), .A(S), .Z(O[247]) );
  ANDN U94 ( .B(A[246]), .A(S), .Z(O[246]) );
  ANDN U95 ( .B(A[245]), .A(S), .Z(O[245]) );
  ANDN U96 ( .B(A[244]), .A(S), .Z(O[244]) );
  ANDN U97 ( .B(A[243]), .A(S), .Z(O[243]) );
  ANDN U98 ( .B(A[242]), .A(S), .Z(O[242]) );
  ANDN U99 ( .B(A[241]), .A(S), .Z(O[241]) );
  ANDN U100 ( .B(A[240]), .A(S), .Z(O[240]) );
  ANDN U101 ( .B(A[23]), .A(S), .Z(O[23]) );
  ANDN U102 ( .B(A[239]), .A(S), .Z(O[239]) );
  ANDN U103 ( .B(A[238]), .A(S), .Z(O[238]) );
  ANDN U104 ( .B(A[237]), .A(S), .Z(O[237]) );
  ANDN U105 ( .B(A[236]), .A(S), .Z(O[236]) );
  ANDN U106 ( .B(A[235]), .A(S), .Z(O[235]) );
  ANDN U107 ( .B(A[234]), .A(S), .Z(O[234]) );
  ANDN U108 ( .B(A[233]), .A(S), .Z(O[233]) );
  ANDN U109 ( .B(A[232]), .A(S), .Z(O[232]) );
  ANDN U110 ( .B(A[231]), .A(S), .Z(O[231]) );
  ANDN U111 ( .B(A[230]), .A(S), .Z(O[230]) );
  ANDN U112 ( .B(A[22]), .A(S), .Z(O[22]) );
  ANDN U113 ( .B(A[229]), .A(S), .Z(O[229]) );
  ANDN U114 ( .B(A[228]), .A(S), .Z(O[228]) );
  ANDN U115 ( .B(A[227]), .A(S), .Z(O[227]) );
  ANDN U116 ( .B(A[226]), .A(S), .Z(O[226]) );
  ANDN U117 ( .B(A[225]), .A(S), .Z(O[225]) );
  ANDN U118 ( .B(A[224]), .A(S), .Z(O[224]) );
  ANDN U119 ( .B(A[223]), .A(S), .Z(O[223]) );
  ANDN U120 ( .B(A[222]), .A(S), .Z(O[222]) );
  ANDN U121 ( .B(A[221]), .A(S), .Z(O[221]) );
  ANDN U122 ( .B(A[220]), .A(S), .Z(O[220]) );
  ANDN U123 ( .B(A[21]), .A(S), .Z(O[21]) );
  ANDN U124 ( .B(A[219]), .A(S), .Z(O[219]) );
  ANDN U125 ( .B(A[218]), .A(S), .Z(O[218]) );
  ANDN U126 ( .B(A[217]), .A(S), .Z(O[217]) );
  ANDN U127 ( .B(A[216]), .A(S), .Z(O[216]) );
  ANDN U128 ( .B(A[215]), .A(S), .Z(O[215]) );
  ANDN U129 ( .B(A[214]), .A(S), .Z(O[214]) );
  ANDN U130 ( .B(A[213]), .A(S), .Z(O[213]) );
  ANDN U131 ( .B(A[212]), .A(S), .Z(O[212]) );
  ANDN U132 ( .B(A[211]), .A(S), .Z(O[211]) );
  ANDN U133 ( .B(A[210]), .A(S), .Z(O[210]) );
  ANDN U134 ( .B(A[20]), .A(S), .Z(O[20]) );
  ANDN U135 ( .B(A[209]), .A(S), .Z(O[209]) );
  ANDN U136 ( .B(A[208]), .A(S), .Z(O[208]) );
  ANDN U137 ( .B(A[207]), .A(S), .Z(O[207]) );
  ANDN U138 ( .B(A[206]), .A(S), .Z(O[206]) );
  ANDN U139 ( .B(A[205]), .A(S), .Z(O[205]) );
  ANDN U140 ( .B(A[204]), .A(S), .Z(O[204]) );
  ANDN U141 ( .B(A[203]), .A(S), .Z(O[203]) );
  ANDN U142 ( .B(A[202]), .A(S), .Z(O[202]) );
  ANDN U143 ( .B(A[201]), .A(S), .Z(O[201]) );
  ANDN U144 ( .B(A[200]), .A(S), .Z(O[200]) );
  ANDN U145 ( .B(A[1]), .A(S), .Z(O[1]) );
  ANDN U146 ( .B(A[19]), .A(S), .Z(O[19]) );
  ANDN U147 ( .B(A[199]), .A(S), .Z(O[199]) );
  ANDN U148 ( .B(A[198]), .A(S), .Z(O[198]) );
  ANDN U149 ( .B(A[197]), .A(S), .Z(O[197]) );
  ANDN U150 ( .B(A[196]), .A(S), .Z(O[196]) );
  ANDN U151 ( .B(A[195]), .A(S), .Z(O[195]) );
  ANDN U152 ( .B(A[194]), .A(S), .Z(O[194]) );
  ANDN U153 ( .B(A[193]), .A(S), .Z(O[193]) );
  ANDN U154 ( .B(A[192]), .A(S), .Z(O[192]) );
  ANDN U155 ( .B(A[191]), .A(S), .Z(O[191]) );
  ANDN U156 ( .B(A[190]), .A(S), .Z(O[190]) );
  ANDN U157 ( .B(A[18]), .A(S), .Z(O[18]) );
  ANDN U158 ( .B(A[189]), .A(S), .Z(O[189]) );
  ANDN U159 ( .B(A[188]), .A(S), .Z(O[188]) );
  ANDN U160 ( .B(A[187]), .A(S), .Z(O[187]) );
  ANDN U161 ( .B(A[186]), .A(S), .Z(O[186]) );
  ANDN U162 ( .B(A[185]), .A(S), .Z(O[185]) );
  ANDN U163 ( .B(A[184]), .A(S), .Z(O[184]) );
  ANDN U164 ( .B(A[183]), .A(S), .Z(O[183]) );
  ANDN U165 ( .B(A[182]), .A(S), .Z(O[182]) );
  ANDN U166 ( .B(A[181]), .A(S), .Z(O[181]) );
  ANDN U167 ( .B(A[180]), .A(S), .Z(O[180]) );
  ANDN U168 ( .B(A[17]), .A(S), .Z(O[17]) );
  ANDN U169 ( .B(A[179]), .A(S), .Z(O[179]) );
  ANDN U170 ( .B(A[178]), .A(S), .Z(O[178]) );
  ANDN U171 ( .B(A[177]), .A(S), .Z(O[177]) );
  ANDN U172 ( .B(A[176]), .A(S), .Z(O[176]) );
  ANDN U173 ( .B(A[175]), .A(S), .Z(O[175]) );
  ANDN U174 ( .B(A[174]), .A(S), .Z(O[174]) );
  ANDN U175 ( .B(A[173]), .A(S), .Z(O[173]) );
  ANDN U176 ( .B(A[172]), .A(S), .Z(O[172]) );
  ANDN U177 ( .B(A[171]), .A(S), .Z(O[171]) );
  ANDN U178 ( .B(A[170]), .A(S), .Z(O[170]) );
  ANDN U179 ( .B(A[16]), .A(S), .Z(O[16]) );
  ANDN U180 ( .B(A[169]), .A(S), .Z(O[169]) );
  ANDN U181 ( .B(A[168]), .A(S), .Z(O[168]) );
  ANDN U182 ( .B(A[167]), .A(S), .Z(O[167]) );
  ANDN U183 ( .B(A[166]), .A(S), .Z(O[166]) );
  ANDN U184 ( .B(A[165]), .A(S), .Z(O[165]) );
  ANDN U185 ( .B(A[164]), .A(S), .Z(O[164]) );
  ANDN U186 ( .B(A[163]), .A(S), .Z(O[163]) );
  ANDN U187 ( .B(A[162]), .A(S), .Z(O[162]) );
  ANDN U188 ( .B(A[161]), .A(S), .Z(O[161]) );
  ANDN U189 ( .B(A[160]), .A(S), .Z(O[160]) );
  ANDN U190 ( .B(A[15]), .A(S), .Z(O[15]) );
  ANDN U191 ( .B(A[159]), .A(S), .Z(O[159]) );
  ANDN U192 ( .B(A[158]), .A(S), .Z(O[158]) );
  ANDN U193 ( .B(A[157]), .A(S), .Z(O[157]) );
  ANDN U194 ( .B(A[156]), .A(S), .Z(O[156]) );
  ANDN U195 ( .B(A[155]), .A(S), .Z(O[155]) );
  ANDN U196 ( .B(A[154]), .A(S), .Z(O[154]) );
  ANDN U197 ( .B(A[153]), .A(S), .Z(O[153]) );
  ANDN U198 ( .B(A[152]), .A(S), .Z(O[152]) );
  ANDN U199 ( .B(A[151]), .A(S), .Z(O[151]) );
  ANDN U200 ( .B(A[150]), .A(S), .Z(O[150]) );
  ANDN U201 ( .B(A[14]), .A(S), .Z(O[14]) );
  ANDN U202 ( .B(A[149]), .A(S), .Z(O[149]) );
  ANDN U203 ( .B(A[148]), .A(S), .Z(O[148]) );
  ANDN U204 ( .B(A[147]), .A(S), .Z(O[147]) );
  ANDN U205 ( .B(A[146]), .A(S), .Z(O[146]) );
  ANDN U206 ( .B(A[145]), .A(S), .Z(O[145]) );
  ANDN U207 ( .B(A[144]), .A(S), .Z(O[144]) );
  ANDN U208 ( .B(A[143]), .A(S), .Z(O[143]) );
  ANDN U209 ( .B(A[142]), .A(S), .Z(O[142]) );
  ANDN U210 ( .B(A[141]), .A(S), .Z(O[141]) );
  ANDN U211 ( .B(A[140]), .A(S), .Z(O[140]) );
  ANDN U212 ( .B(A[13]), .A(S), .Z(O[13]) );
  ANDN U213 ( .B(A[139]), .A(S), .Z(O[139]) );
  ANDN U214 ( .B(A[138]), .A(S), .Z(O[138]) );
  ANDN U215 ( .B(A[137]), .A(S), .Z(O[137]) );
  ANDN U216 ( .B(A[136]), .A(S), .Z(O[136]) );
  ANDN U217 ( .B(A[135]), .A(S), .Z(O[135]) );
  ANDN U218 ( .B(A[134]), .A(S), .Z(O[134]) );
  ANDN U219 ( .B(A[133]), .A(S), .Z(O[133]) );
  ANDN U220 ( .B(A[132]), .A(S), .Z(O[132]) );
  ANDN U221 ( .B(A[131]), .A(S), .Z(O[131]) );
  ANDN U222 ( .B(A[130]), .A(S), .Z(O[130]) );
  ANDN U223 ( .B(A[12]), .A(S), .Z(O[12]) );
  ANDN U224 ( .B(A[129]), .A(S), .Z(O[129]) );
  ANDN U225 ( .B(A[128]), .A(S), .Z(O[128]) );
  ANDN U226 ( .B(A[127]), .A(S), .Z(O[127]) );
  ANDN U227 ( .B(A[126]), .A(S), .Z(O[126]) );
  ANDN U228 ( .B(A[125]), .A(S), .Z(O[125]) );
  ANDN U229 ( .B(A[124]), .A(S), .Z(O[124]) );
  ANDN U230 ( .B(A[123]), .A(S), .Z(O[123]) );
  ANDN U231 ( .B(A[122]), .A(S), .Z(O[122]) );
  ANDN U232 ( .B(A[121]), .A(S), .Z(O[121]) );
  ANDN U233 ( .B(A[120]), .A(S), .Z(O[120]) );
  ANDN U234 ( .B(A[11]), .A(S), .Z(O[11]) );
  ANDN U235 ( .B(A[119]), .A(S), .Z(O[119]) );
  ANDN U236 ( .B(A[118]), .A(S), .Z(O[118]) );
  ANDN U237 ( .B(A[117]), .A(S), .Z(O[117]) );
  ANDN U238 ( .B(A[116]), .A(S), .Z(O[116]) );
  ANDN U239 ( .B(A[115]), .A(S), .Z(O[115]) );
  ANDN U240 ( .B(A[114]), .A(S), .Z(O[114]) );
  ANDN U241 ( .B(A[113]), .A(S), .Z(O[113]) );
  ANDN U242 ( .B(A[112]), .A(S), .Z(O[112]) );
  ANDN U243 ( .B(A[111]), .A(S), .Z(O[111]) );
  ANDN U244 ( .B(A[110]), .A(S), .Z(O[110]) );
  ANDN U245 ( .B(A[10]), .A(S), .Z(O[10]) );
  ANDN U246 ( .B(A[109]), .A(S), .Z(O[109]) );
  ANDN U247 ( .B(A[108]), .A(S), .Z(O[108]) );
  ANDN U248 ( .B(A[107]), .A(S), .Z(O[107]) );
  ANDN U249 ( .B(A[106]), .A(S), .Z(O[106]) );
  ANDN U250 ( .B(A[105]), .A(S), .Z(O[105]) );
  ANDN U251 ( .B(A[104]), .A(S), .Z(O[104]) );
  ANDN U252 ( .B(A[103]), .A(S), .Z(O[103]) );
  ANDN U253 ( .B(A[102]), .A(S), .Z(O[102]) );
  ANDN U254 ( .B(A[101]), .A(S), .Z(O[101]) );
  ANDN U255 ( .B(A[100]), .A(S), .Z(O[100]) );
  ANDN U256 ( .B(A[0]), .A(S), .Z(O[0]) );
endmodule


module FA_2322 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(CI), .B(A), .Z(S) );
endmodule


module FA_2323 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  ANDN U1 ( .B(CI), .A(S), .Z(CO) );
  XOR U2 ( .A(A), .B(CI), .Z(S) );
endmodule


module FA_2324 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2325 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2326 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2327 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2328 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2329 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2330 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2331 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2332 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2333 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2334 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2335 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2336 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2337 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2338 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2339 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2340 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2341 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2342 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2343 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2344 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2345 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2346 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2347 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2348 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2349 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2350 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2351 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2352 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2353 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2354 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2355 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2356 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2357 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2358 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2359 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2360 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2361 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2362 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2363 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2364 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2365 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2366 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2367 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2368 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2369 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2370 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2371 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2372 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2373 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2374 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2375 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2376 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2377 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2378 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2379 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2380 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2381 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2382 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2383 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2384 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2385 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2386 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2387 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2388 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2389 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2390 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2391 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2392 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2393 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2394 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2395 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2396 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2397 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2398 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2399 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2400 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2401 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2402 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2403 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2404 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2405 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2406 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2407 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2408 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2409 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2410 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2411 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2412 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2413 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2414 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2415 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2416 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2417 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2418 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2419 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2420 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2421 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2422 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2423 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2424 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2425 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2426 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2427 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2428 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2429 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2430 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2431 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2432 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2433 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2434 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2435 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2436 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2437 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2438 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2439 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2440 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2441 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2442 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2443 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2444 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2445 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2446 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2447 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2448 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2449 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2450 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2451 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2452 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2453 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2454 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2455 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2456 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2457 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2458 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2459 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2460 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2461 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2462 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2463 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2464 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2465 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2466 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2467 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2468 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2469 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2470 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2471 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2472 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2473 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2474 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2475 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2476 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2477 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2478 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2479 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2480 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2481 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2482 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2483 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2484 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2485 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2486 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2487 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2488 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2489 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2490 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2491 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2492 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2493 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2494 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2495 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2496 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2497 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2498 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2499 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2500 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2501 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2502 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2503 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2504 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2505 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2506 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2507 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2508 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2509 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2510 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2511 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2512 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2513 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2514 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2515 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2516 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2517 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2518 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2519 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2520 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2521 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2522 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2523 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2524 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2525 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2526 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2527 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2528 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2529 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2530 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2531 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2532 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2533 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2534 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2535 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2536 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2537 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2538 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2539 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2540 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2541 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2542 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2543 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2544 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2545 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2546 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2547 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2548 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2549 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2550 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2551 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2552 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2553 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2554 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2555 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2556 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2557 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2558 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2559 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2560 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2561 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2562 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2563 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2564 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2565 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2566 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2567 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2568 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2569 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2570 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2571 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2572 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2573 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2574 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2575 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2576 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2577 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2578 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_2579 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N258_1_1 ( A, B, CI, S, CO );
  input [257:0] A;
  input [257:0] B;
  output [257:0] S;
  input CI;
  output CO;

  wire   [257:1] C;

  FA_2579 \FAINST[0].FA_  ( .A(1'b0), .B(B[0]), .CI(1'b0), .S(S[0]) );
  FA_2578 \FAINST[1].FA_  ( .A(A[1]), .B(B[1]), .CI(1'b0), .S(S[1]), .CO(C[2])
         );
  FA_2577 \FAINST[2].FA_  ( .A(A[2]), .B(B[2]), .CI(C[2]), .S(S[2]), .CO(C[3])
         );
  FA_2576 \FAINST[3].FA_  ( .A(A[3]), .B(B[3]), .CI(C[3]), .S(S[3]), .CO(C[4])
         );
  FA_2575 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(C[4]), .S(S[4]), .CO(C[5])
         );
  FA_2574 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_2573 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_2572 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_2571 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_2570 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_2569 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_2568 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_2567 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_2566 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_2565 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_2564 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_2563 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_2562 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_2561 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_2560 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_2559 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_2558 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_2557 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_2556 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_2555 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_2554 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_2553 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_2552 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_2551 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_2550 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_2549 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_2548 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]), .CO(
        C[32]) );
  FA_2547 \FAINST[32].FA_  ( .A(A[32]), .B(B[32]), .CI(C[32]), .S(S[32]), .CO(
        C[33]) );
  FA_2546 \FAINST[33].FA_  ( .A(A[33]), .B(B[33]), .CI(C[33]), .S(S[33]), .CO(
        C[34]) );
  FA_2545 \FAINST[34].FA_  ( .A(A[34]), .B(B[34]), .CI(C[34]), .S(S[34]), .CO(
        C[35]) );
  FA_2544 \FAINST[35].FA_  ( .A(A[35]), .B(B[35]), .CI(C[35]), .S(S[35]), .CO(
        C[36]) );
  FA_2543 \FAINST[36].FA_  ( .A(A[36]), .B(B[36]), .CI(C[36]), .S(S[36]), .CO(
        C[37]) );
  FA_2542 \FAINST[37].FA_  ( .A(A[37]), .B(B[37]), .CI(C[37]), .S(S[37]), .CO(
        C[38]) );
  FA_2541 \FAINST[38].FA_  ( .A(A[38]), .B(B[38]), .CI(C[38]), .S(S[38]), .CO(
        C[39]) );
  FA_2540 \FAINST[39].FA_  ( .A(A[39]), .B(B[39]), .CI(C[39]), .S(S[39]), .CO(
        C[40]) );
  FA_2539 \FAINST[40].FA_  ( .A(A[40]), .B(B[40]), .CI(C[40]), .S(S[40]), .CO(
        C[41]) );
  FA_2538 \FAINST[41].FA_  ( .A(A[41]), .B(B[41]), .CI(C[41]), .S(S[41]), .CO(
        C[42]) );
  FA_2537 \FAINST[42].FA_  ( .A(A[42]), .B(B[42]), .CI(C[42]), .S(S[42]), .CO(
        C[43]) );
  FA_2536 \FAINST[43].FA_  ( .A(A[43]), .B(B[43]), .CI(C[43]), .S(S[43]), .CO(
        C[44]) );
  FA_2535 \FAINST[44].FA_  ( .A(A[44]), .B(B[44]), .CI(C[44]), .S(S[44]), .CO(
        C[45]) );
  FA_2534 \FAINST[45].FA_  ( .A(A[45]), .B(B[45]), .CI(C[45]), .S(S[45]), .CO(
        C[46]) );
  FA_2533 \FAINST[46].FA_  ( .A(A[46]), .B(B[46]), .CI(C[46]), .S(S[46]), .CO(
        C[47]) );
  FA_2532 \FAINST[47].FA_  ( .A(A[47]), .B(B[47]), .CI(C[47]), .S(S[47]), .CO(
        C[48]) );
  FA_2531 \FAINST[48].FA_  ( .A(A[48]), .B(B[48]), .CI(C[48]), .S(S[48]), .CO(
        C[49]) );
  FA_2530 \FAINST[49].FA_  ( .A(A[49]), .B(B[49]), .CI(C[49]), .S(S[49]), .CO(
        C[50]) );
  FA_2529 \FAINST[50].FA_  ( .A(A[50]), .B(B[50]), .CI(C[50]), .S(S[50]), .CO(
        C[51]) );
  FA_2528 \FAINST[51].FA_  ( .A(A[51]), .B(B[51]), .CI(C[51]), .S(S[51]), .CO(
        C[52]) );
  FA_2527 \FAINST[52].FA_  ( .A(A[52]), .B(B[52]), .CI(C[52]), .S(S[52]), .CO(
        C[53]) );
  FA_2526 \FAINST[53].FA_  ( .A(A[53]), .B(B[53]), .CI(C[53]), .S(S[53]), .CO(
        C[54]) );
  FA_2525 \FAINST[54].FA_  ( .A(A[54]), .B(B[54]), .CI(C[54]), .S(S[54]), .CO(
        C[55]) );
  FA_2524 \FAINST[55].FA_  ( .A(A[55]), .B(B[55]), .CI(C[55]), .S(S[55]), .CO(
        C[56]) );
  FA_2523 \FAINST[56].FA_  ( .A(A[56]), .B(B[56]), .CI(C[56]), .S(S[56]), .CO(
        C[57]) );
  FA_2522 \FAINST[57].FA_  ( .A(A[57]), .B(B[57]), .CI(C[57]), .S(S[57]), .CO(
        C[58]) );
  FA_2521 \FAINST[58].FA_  ( .A(A[58]), .B(B[58]), .CI(C[58]), .S(S[58]), .CO(
        C[59]) );
  FA_2520 \FAINST[59].FA_  ( .A(A[59]), .B(B[59]), .CI(C[59]), .S(S[59]), .CO(
        C[60]) );
  FA_2519 \FAINST[60].FA_  ( .A(A[60]), .B(B[60]), .CI(C[60]), .S(S[60]), .CO(
        C[61]) );
  FA_2518 \FAINST[61].FA_  ( .A(A[61]), .B(B[61]), .CI(C[61]), .S(S[61]), .CO(
        C[62]) );
  FA_2517 \FAINST[62].FA_  ( .A(A[62]), .B(B[62]), .CI(C[62]), .S(S[62]), .CO(
        C[63]) );
  FA_2516 \FAINST[63].FA_  ( .A(A[63]), .B(B[63]), .CI(C[63]), .S(S[63]), .CO(
        C[64]) );
  FA_2515 \FAINST[64].FA_  ( .A(A[64]), .B(B[64]), .CI(C[64]), .S(S[64]), .CO(
        C[65]) );
  FA_2514 \FAINST[65].FA_  ( .A(A[65]), .B(B[65]), .CI(C[65]), .S(S[65]), .CO(
        C[66]) );
  FA_2513 \FAINST[66].FA_  ( .A(A[66]), .B(B[66]), .CI(C[66]), .S(S[66]), .CO(
        C[67]) );
  FA_2512 \FAINST[67].FA_  ( .A(A[67]), .B(B[67]), .CI(C[67]), .S(S[67]), .CO(
        C[68]) );
  FA_2511 \FAINST[68].FA_  ( .A(A[68]), .B(B[68]), .CI(C[68]), .S(S[68]), .CO(
        C[69]) );
  FA_2510 \FAINST[69].FA_  ( .A(A[69]), .B(B[69]), .CI(C[69]), .S(S[69]), .CO(
        C[70]) );
  FA_2509 \FAINST[70].FA_  ( .A(A[70]), .B(B[70]), .CI(C[70]), .S(S[70]), .CO(
        C[71]) );
  FA_2508 \FAINST[71].FA_  ( .A(A[71]), .B(B[71]), .CI(C[71]), .S(S[71]), .CO(
        C[72]) );
  FA_2507 \FAINST[72].FA_  ( .A(A[72]), .B(B[72]), .CI(C[72]), .S(S[72]), .CO(
        C[73]) );
  FA_2506 \FAINST[73].FA_  ( .A(A[73]), .B(B[73]), .CI(C[73]), .S(S[73]), .CO(
        C[74]) );
  FA_2505 \FAINST[74].FA_  ( .A(A[74]), .B(B[74]), .CI(C[74]), .S(S[74]), .CO(
        C[75]) );
  FA_2504 \FAINST[75].FA_  ( .A(A[75]), .B(B[75]), .CI(C[75]), .S(S[75]), .CO(
        C[76]) );
  FA_2503 \FAINST[76].FA_  ( .A(A[76]), .B(B[76]), .CI(C[76]), .S(S[76]), .CO(
        C[77]) );
  FA_2502 \FAINST[77].FA_  ( .A(A[77]), .B(B[77]), .CI(C[77]), .S(S[77]), .CO(
        C[78]) );
  FA_2501 \FAINST[78].FA_  ( .A(A[78]), .B(B[78]), .CI(C[78]), .S(S[78]), .CO(
        C[79]) );
  FA_2500 \FAINST[79].FA_  ( .A(A[79]), .B(B[79]), .CI(C[79]), .S(S[79]), .CO(
        C[80]) );
  FA_2499 \FAINST[80].FA_  ( .A(A[80]), .B(B[80]), .CI(C[80]), .S(S[80]), .CO(
        C[81]) );
  FA_2498 \FAINST[81].FA_  ( .A(A[81]), .B(B[81]), .CI(C[81]), .S(S[81]), .CO(
        C[82]) );
  FA_2497 \FAINST[82].FA_  ( .A(A[82]), .B(B[82]), .CI(C[82]), .S(S[82]), .CO(
        C[83]) );
  FA_2496 \FAINST[83].FA_  ( .A(A[83]), .B(B[83]), .CI(C[83]), .S(S[83]), .CO(
        C[84]) );
  FA_2495 \FAINST[84].FA_  ( .A(A[84]), .B(B[84]), .CI(C[84]), .S(S[84]), .CO(
        C[85]) );
  FA_2494 \FAINST[85].FA_  ( .A(A[85]), .B(B[85]), .CI(C[85]), .S(S[85]), .CO(
        C[86]) );
  FA_2493 \FAINST[86].FA_  ( .A(A[86]), .B(B[86]), .CI(C[86]), .S(S[86]), .CO(
        C[87]) );
  FA_2492 \FAINST[87].FA_  ( .A(A[87]), .B(B[87]), .CI(C[87]), .S(S[87]), .CO(
        C[88]) );
  FA_2491 \FAINST[88].FA_  ( .A(A[88]), .B(B[88]), .CI(C[88]), .S(S[88]), .CO(
        C[89]) );
  FA_2490 \FAINST[89].FA_  ( .A(A[89]), .B(B[89]), .CI(C[89]), .S(S[89]), .CO(
        C[90]) );
  FA_2489 \FAINST[90].FA_  ( .A(A[90]), .B(B[90]), .CI(C[90]), .S(S[90]), .CO(
        C[91]) );
  FA_2488 \FAINST[91].FA_  ( .A(A[91]), .B(B[91]), .CI(C[91]), .S(S[91]), .CO(
        C[92]) );
  FA_2487 \FAINST[92].FA_  ( .A(A[92]), .B(B[92]), .CI(C[92]), .S(S[92]), .CO(
        C[93]) );
  FA_2486 \FAINST[93].FA_  ( .A(A[93]), .B(B[93]), .CI(C[93]), .S(S[93]), .CO(
        C[94]) );
  FA_2485 \FAINST[94].FA_  ( .A(A[94]), .B(B[94]), .CI(C[94]), .S(S[94]), .CO(
        C[95]) );
  FA_2484 \FAINST[95].FA_  ( .A(A[95]), .B(B[95]), .CI(C[95]), .S(S[95]), .CO(
        C[96]) );
  FA_2483 \FAINST[96].FA_  ( .A(A[96]), .B(B[96]), .CI(C[96]), .S(S[96]), .CO(
        C[97]) );
  FA_2482 \FAINST[97].FA_  ( .A(A[97]), .B(B[97]), .CI(C[97]), .S(S[97]), .CO(
        C[98]) );
  FA_2481 \FAINST[98].FA_  ( .A(A[98]), .B(B[98]), .CI(C[98]), .S(S[98]), .CO(
        C[99]) );
  FA_2480 \FAINST[99].FA_  ( .A(A[99]), .B(B[99]), .CI(C[99]), .S(S[99]), .CO(
        C[100]) );
  FA_2479 \FAINST[100].FA_  ( .A(A[100]), .B(B[100]), .CI(C[100]), .S(S[100]), 
        .CO(C[101]) );
  FA_2478 \FAINST[101].FA_  ( .A(A[101]), .B(B[101]), .CI(C[101]), .S(S[101]), 
        .CO(C[102]) );
  FA_2477 \FAINST[102].FA_  ( .A(A[102]), .B(B[102]), .CI(C[102]), .S(S[102]), 
        .CO(C[103]) );
  FA_2476 \FAINST[103].FA_  ( .A(A[103]), .B(B[103]), .CI(C[103]), .S(S[103]), 
        .CO(C[104]) );
  FA_2475 \FAINST[104].FA_  ( .A(A[104]), .B(B[104]), .CI(C[104]), .S(S[104]), 
        .CO(C[105]) );
  FA_2474 \FAINST[105].FA_  ( .A(A[105]), .B(B[105]), .CI(C[105]), .S(S[105]), 
        .CO(C[106]) );
  FA_2473 \FAINST[106].FA_  ( .A(A[106]), .B(B[106]), .CI(C[106]), .S(S[106]), 
        .CO(C[107]) );
  FA_2472 \FAINST[107].FA_  ( .A(A[107]), .B(B[107]), .CI(C[107]), .S(S[107]), 
        .CO(C[108]) );
  FA_2471 \FAINST[108].FA_  ( .A(A[108]), .B(B[108]), .CI(C[108]), .S(S[108]), 
        .CO(C[109]) );
  FA_2470 \FAINST[109].FA_  ( .A(A[109]), .B(B[109]), .CI(C[109]), .S(S[109]), 
        .CO(C[110]) );
  FA_2469 \FAINST[110].FA_  ( .A(A[110]), .B(B[110]), .CI(C[110]), .S(S[110]), 
        .CO(C[111]) );
  FA_2468 \FAINST[111].FA_  ( .A(A[111]), .B(B[111]), .CI(C[111]), .S(S[111]), 
        .CO(C[112]) );
  FA_2467 \FAINST[112].FA_  ( .A(A[112]), .B(B[112]), .CI(C[112]), .S(S[112]), 
        .CO(C[113]) );
  FA_2466 \FAINST[113].FA_  ( .A(A[113]), .B(B[113]), .CI(C[113]), .S(S[113]), 
        .CO(C[114]) );
  FA_2465 \FAINST[114].FA_  ( .A(A[114]), .B(B[114]), .CI(C[114]), .S(S[114]), 
        .CO(C[115]) );
  FA_2464 \FAINST[115].FA_  ( .A(A[115]), .B(B[115]), .CI(C[115]), .S(S[115]), 
        .CO(C[116]) );
  FA_2463 \FAINST[116].FA_  ( .A(A[116]), .B(B[116]), .CI(C[116]), .S(S[116]), 
        .CO(C[117]) );
  FA_2462 \FAINST[117].FA_  ( .A(A[117]), .B(B[117]), .CI(C[117]), .S(S[117]), 
        .CO(C[118]) );
  FA_2461 \FAINST[118].FA_  ( .A(A[118]), .B(B[118]), .CI(C[118]), .S(S[118]), 
        .CO(C[119]) );
  FA_2460 \FAINST[119].FA_  ( .A(A[119]), .B(B[119]), .CI(C[119]), .S(S[119]), 
        .CO(C[120]) );
  FA_2459 \FAINST[120].FA_  ( .A(A[120]), .B(B[120]), .CI(C[120]), .S(S[120]), 
        .CO(C[121]) );
  FA_2458 \FAINST[121].FA_  ( .A(A[121]), .B(B[121]), .CI(C[121]), .S(S[121]), 
        .CO(C[122]) );
  FA_2457 \FAINST[122].FA_  ( .A(A[122]), .B(B[122]), .CI(C[122]), .S(S[122]), 
        .CO(C[123]) );
  FA_2456 \FAINST[123].FA_  ( .A(A[123]), .B(B[123]), .CI(C[123]), .S(S[123]), 
        .CO(C[124]) );
  FA_2455 \FAINST[124].FA_  ( .A(A[124]), .B(B[124]), .CI(C[124]), .S(S[124]), 
        .CO(C[125]) );
  FA_2454 \FAINST[125].FA_  ( .A(A[125]), .B(B[125]), .CI(C[125]), .S(S[125]), 
        .CO(C[126]) );
  FA_2453 \FAINST[126].FA_  ( .A(A[126]), .B(B[126]), .CI(C[126]), .S(S[126]), 
        .CO(C[127]) );
  FA_2452 \FAINST[127].FA_  ( .A(A[127]), .B(B[127]), .CI(C[127]), .S(S[127]), 
        .CO(C[128]) );
  FA_2451 \FAINST[128].FA_  ( .A(A[128]), .B(B[128]), .CI(C[128]), .S(S[128]), 
        .CO(C[129]) );
  FA_2450 \FAINST[129].FA_  ( .A(A[129]), .B(B[129]), .CI(C[129]), .S(S[129]), 
        .CO(C[130]) );
  FA_2449 \FAINST[130].FA_  ( .A(A[130]), .B(B[130]), .CI(C[130]), .S(S[130]), 
        .CO(C[131]) );
  FA_2448 \FAINST[131].FA_  ( .A(A[131]), .B(B[131]), .CI(C[131]), .S(S[131]), 
        .CO(C[132]) );
  FA_2447 \FAINST[132].FA_  ( .A(A[132]), .B(B[132]), .CI(C[132]), .S(S[132]), 
        .CO(C[133]) );
  FA_2446 \FAINST[133].FA_  ( .A(A[133]), .B(B[133]), .CI(C[133]), .S(S[133]), 
        .CO(C[134]) );
  FA_2445 \FAINST[134].FA_  ( .A(A[134]), .B(B[134]), .CI(C[134]), .S(S[134]), 
        .CO(C[135]) );
  FA_2444 \FAINST[135].FA_  ( .A(A[135]), .B(B[135]), .CI(C[135]), .S(S[135]), 
        .CO(C[136]) );
  FA_2443 \FAINST[136].FA_  ( .A(A[136]), .B(B[136]), .CI(C[136]), .S(S[136]), 
        .CO(C[137]) );
  FA_2442 \FAINST[137].FA_  ( .A(A[137]), .B(B[137]), .CI(C[137]), .S(S[137]), 
        .CO(C[138]) );
  FA_2441 \FAINST[138].FA_  ( .A(A[138]), .B(B[138]), .CI(C[138]), .S(S[138]), 
        .CO(C[139]) );
  FA_2440 \FAINST[139].FA_  ( .A(A[139]), .B(B[139]), .CI(C[139]), .S(S[139]), 
        .CO(C[140]) );
  FA_2439 \FAINST[140].FA_  ( .A(A[140]), .B(B[140]), .CI(C[140]), .S(S[140]), 
        .CO(C[141]) );
  FA_2438 \FAINST[141].FA_  ( .A(A[141]), .B(B[141]), .CI(C[141]), .S(S[141]), 
        .CO(C[142]) );
  FA_2437 \FAINST[142].FA_  ( .A(A[142]), .B(B[142]), .CI(C[142]), .S(S[142]), 
        .CO(C[143]) );
  FA_2436 \FAINST[143].FA_  ( .A(A[143]), .B(B[143]), .CI(C[143]), .S(S[143]), 
        .CO(C[144]) );
  FA_2435 \FAINST[144].FA_  ( .A(A[144]), .B(B[144]), .CI(C[144]), .S(S[144]), 
        .CO(C[145]) );
  FA_2434 \FAINST[145].FA_  ( .A(A[145]), .B(B[145]), .CI(C[145]), .S(S[145]), 
        .CO(C[146]) );
  FA_2433 \FAINST[146].FA_  ( .A(A[146]), .B(B[146]), .CI(C[146]), .S(S[146]), 
        .CO(C[147]) );
  FA_2432 \FAINST[147].FA_  ( .A(A[147]), .B(B[147]), .CI(C[147]), .S(S[147]), 
        .CO(C[148]) );
  FA_2431 \FAINST[148].FA_  ( .A(A[148]), .B(B[148]), .CI(C[148]), .S(S[148]), 
        .CO(C[149]) );
  FA_2430 \FAINST[149].FA_  ( .A(A[149]), .B(B[149]), .CI(C[149]), .S(S[149]), 
        .CO(C[150]) );
  FA_2429 \FAINST[150].FA_  ( .A(A[150]), .B(B[150]), .CI(C[150]), .S(S[150]), 
        .CO(C[151]) );
  FA_2428 \FAINST[151].FA_  ( .A(A[151]), .B(B[151]), .CI(C[151]), .S(S[151]), 
        .CO(C[152]) );
  FA_2427 \FAINST[152].FA_  ( .A(A[152]), .B(B[152]), .CI(C[152]), .S(S[152]), 
        .CO(C[153]) );
  FA_2426 \FAINST[153].FA_  ( .A(A[153]), .B(B[153]), .CI(C[153]), .S(S[153]), 
        .CO(C[154]) );
  FA_2425 \FAINST[154].FA_  ( .A(A[154]), .B(B[154]), .CI(C[154]), .S(S[154]), 
        .CO(C[155]) );
  FA_2424 \FAINST[155].FA_  ( .A(A[155]), .B(B[155]), .CI(C[155]), .S(S[155]), 
        .CO(C[156]) );
  FA_2423 \FAINST[156].FA_  ( .A(A[156]), .B(B[156]), .CI(C[156]), .S(S[156]), 
        .CO(C[157]) );
  FA_2422 \FAINST[157].FA_  ( .A(A[157]), .B(B[157]), .CI(C[157]), .S(S[157]), 
        .CO(C[158]) );
  FA_2421 \FAINST[158].FA_  ( .A(A[158]), .B(B[158]), .CI(C[158]), .S(S[158]), 
        .CO(C[159]) );
  FA_2420 \FAINST[159].FA_  ( .A(A[159]), .B(B[159]), .CI(C[159]), .S(S[159]), 
        .CO(C[160]) );
  FA_2419 \FAINST[160].FA_  ( .A(A[160]), .B(B[160]), .CI(C[160]), .S(S[160]), 
        .CO(C[161]) );
  FA_2418 \FAINST[161].FA_  ( .A(A[161]), .B(B[161]), .CI(C[161]), .S(S[161]), 
        .CO(C[162]) );
  FA_2417 \FAINST[162].FA_  ( .A(A[162]), .B(B[162]), .CI(C[162]), .S(S[162]), 
        .CO(C[163]) );
  FA_2416 \FAINST[163].FA_  ( .A(A[163]), .B(B[163]), .CI(C[163]), .S(S[163]), 
        .CO(C[164]) );
  FA_2415 \FAINST[164].FA_  ( .A(A[164]), .B(B[164]), .CI(C[164]), .S(S[164]), 
        .CO(C[165]) );
  FA_2414 \FAINST[165].FA_  ( .A(A[165]), .B(B[165]), .CI(C[165]), .S(S[165]), 
        .CO(C[166]) );
  FA_2413 \FAINST[166].FA_  ( .A(A[166]), .B(B[166]), .CI(C[166]), .S(S[166]), 
        .CO(C[167]) );
  FA_2412 \FAINST[167].FA_  ( .A(A[167]), .B(B[167]), .CI(C[167]), .S(S[167]), 
        .CO(C[168]) );
  FA_2411 \FAINST[168].FA_  ( .A(A[168]), .B(B[168]), .CI(C[168]), .S(S[168]), 
        .CO(C[169]) );
  FA_2410 \FAINST[169].FA_  ( .A(A[169]), .B(B[169]), .CI(C[169]), .S(S[169]), 
        .CO(C[170]) );
  FA_2409 \FAINST[170].FA_  ( .A(A[170]), .B(B[170]), .CI(C[170]), .S(S[170]), 
        .CO(C[171]) );
  FA_2408 \FAINST[171].FA_  ( .A(A[171]), .B(B[171]), .CI(C[171]), .S(S[171]), 
        .CO(C[172]) );
  FA_2407 \FAINST[172].FA_  ( .A(A[172]), .B(B[172]), .CI(C[172]), .S(S[172]), 
        .CO(C[173]) );
  FA_2406 \FAINST[173].FA_  ( .A(A[173]), .B(B[173]), .CI(C[173]), .S(S[173]), 
        .CO(C[174]) );
  FA_2405 \FAINST[174].FA_  ( .A(A[174]), .B(B[174]), .CI(C[174]), .S(S[174]), 
        .CO(C[175]) );
  FA_2404 \FAINST[175].FA_  ( .A(A[175]), .B(B[175]), .CI(C[175]), .S(S[175]), 
        .CO(C[176]) );
  FA_2403 \FAINST[176].FA_  ( .A(A[176]), .B(B[176]), .CI(C[176]), .S(S[176]), 
        .CO(C[177]) );
  FA_2402 \FAINST[177].FA_  ( .A(A[177]), .B(B[177]), .CI(C[177]), .S(S[177]), 
        .CO(C[178]) );
  FA_2401 \FAINST[178].FA_  ( .A(A[178]), .B(B[178]), .CI(C[178]), .S(S[178]), 
        .CO(C[179]) );
  FA_2400 \FAINST[179].FA_  ( .A(A[179]), .B(B[179]), .CI(C[179]), .S(S[179]), 
        .CO(C[180]) );
  FA_2399 \FAINST[180].FA_  ( .A(A[180]), .B(B[180]), .CI(C[180]), .S(S[180]), 
        .CO(C[181]) );
  FA_2398 \FAINST[181].FA_  ( .A(A[181]), .B(B[181]), .CI(C[181]), .S(S[181]), 
        .CO(C[182]) );
  FA_2397 \FAINST[182].FA_  ( .A(A[182]), .B(B[182]), .CI(C[182]), .S(S[182]), 
        .CO(C[183]) );
  FA_2396 \FAINST[183].FA_  ( .A(A[183]), .B(B[183]), .CI(C[183]), .S(S[183]), 
        .CO(C[184]) );
  FA_2395 \FAINST[184].FA_  ( .A(A[184]), .B(B[184]), .CI(C[184]), .S(S[184]), 
        .CO(C[185]) );
  FA_2394 \FAINST[185].FA_  ( .A(A[185]), .B(B[185]), .CI(C[185]), .S(S[185]), 
        .CO(C[186]) );
  FA_2393 \FAINST[186].FA_  ( .A(A[186]), .B(B[186]), .CI(C[186]), .S(S[186]), 
        .CO(C[187]) );
  FA_2392 \FAINST[187].FA_  ( .A(A[187]), .B(B[187]), .CI(C[187]), .S(S[187]), 
        .CO(C[188]) );
  FA_2391 \FAINST[188].FA_  ( .A(A[188]), .B(B[188]), .CI(C[188]), .S(S[188]), 
        .CO(C[189]) );
  FA_2390 \FAINST[189].FA_  ( .A(A[189]), .B(B[189]), .CI(C[189]), .S(S[189]), 
        .CO(C[190]) );
  FA_2389 \FAINST[190].FA_  ( .A(A[190]), .B(B[190]), .CI(C[190]), .S(S[190]), 
        .CO(C[191]) );
  FA_2388 \FAINST[191].FA_  ( .A(A[191]), .B(B[191]), .CI(C[191]), .S(S[191]), 
        .CO(C[192]) );
  FA_2387 \FAINST[192].FA_  ( .A(A[192]), .B(B[192]), .CI(C[192]), .S(S[192]), 
        .CO(C[193]) );
  FA_2386 \FAINST[193].FA_  ( .A(A[193]), .B(B[193]), .CI(C[193]), .S(S[193]), 
        .CO(C[194]) );
  FA_2385 \FAINST[194].FA_  ( .A(A[194]), .B(B[194]), .CI(C[194]), .S(S[194]), 
        .CO(C[195]) );
  FA_2384 \FAINST[195].FA_  ( .A(A[195]), .B(B[195]), .CI(C[195]), .S(S[195]), 
        .CO(C[196]) );
  FA_2383 \FAINST[196].FA_  ( .A(A[196]), .B(B[196]), .CI(C[196]), .S(S[196]), 
        .CO(C[197]) );
  FA_2382 \FAINST[197].FA_  ( .A(A[197]), .B(B[197]), .CI(C[197]), .S(S[197]), 
        .CO(C[198]) );
  FA_2381 \FAINST[198].FA_  ( .A(A[198]), .B(B[198]), .CI(C[198]), .S(S[198]), 
        .CO(C[199]) );
  FA_2380 \FAINST[199].FA_  ( .A(A[199]), .B(B[199]), .CI(C[199]), .S(S[199]), 
        .CO(C[200]) );
  FA_2379 \FAINST[200].FA_  ( .A(A[200]), .B(B[200]), .CI(C[200]), .S(S[200]), 
        .CO(C[201]) );
  FA_2378 \FAINST[201].FA_  ( .A(A[201]), .B(B[201]), .CI(C[201]), .S(S[201]), 
        .CO(C[202]) );
  FA_2377 \FAINST[202].FA_  ( .A(A[202]), .B(B[202]), .CI(C[202]), .S(S[202]), 
        .CO(C[203]) );
  FA_2376 \FAINST[203].FA_  ( .A(A[203]), .B(B[203]), .CI(C[203]), .S(S[203]), 
        .CO(C[204]) );
  FA_2375 \FAINST[204].FA_  ( .A(A[204]), .B(B[204]), .CI(C[204]), .S(S[204]), 
        .CO(C[205]) );
  FA_2374 \FAINST[205].FA_  ( .A(A[205]), .B(B[205]), .CI(C[205]), .S(S[205]), 
        .CO(C[206]) );
  FA_2373 \FAINST[206].FA_  ( .A(A[206]), .B(B[206]), .CI(C[206]), .S(S[206]), 
        .CO(C[207]) );
  FA_2372 \FAINST[207].FA_  ( .A(A[207]), .B(B[207]), .CI(C[207]), .S(S[207]), 
        .CO(C[208]) );
  FA_2371 \FAINST[208].FA_  ( .A(A[208]), .B(B[208]), .CI(C[208]), .S(S[208]), 
        .CO(C[209]) );
  FA_2370 \FAINST[209].FA_  ( .A(A[209]), .B(B[209]), .CI(C[209]), .S(S[209]), 
        .CO(C[210]) );
  FA_2369 \FAINST[210].FA_  ( .A(A[210]), .B(B[210]), .CI(C[210]), .S(S[210]), 
        .CO(C[211]) );
  FA_2368 \FAINST[211].FA_  ( .A(A[211]), .B(B[211]), .CI(C[211]), .S(S[211]), 
        .CO(C[212]) );
  FA_2367 \FAINST[212].FA_  ( .A(A[212]), .B(B[212]), .CI(C[212]), .S(S[212]), 
        .CO(C[213]) );
  FA_2366 \FAINST[213].FA_  ( .A(A[213]), .B(B[213]), .CI(C[213]), .S(S[213]), 
        .CO(C[214]) );
  FA_2365 \FAINST[214].FA_  ( .A(A[214]), .B(B[214]), .CI(C[214]), .S(S[214]), 
        .CO(C[215]) );
  FA_2364 \FAINST[215].FA_  ( .A(A[215]), .B(B[215]), .CI(C[215]), .S(S[215]), 
        .CO(C[216]) );
  FA_2363 \FAINST[216].FA_  ( .A(A[216]), .B(B[216]), .CI(C[216]), .S(S[216]), 
        .CO(C[217]) );
  FA_2362 \FAINST[217].FA_  ( .A(A[217]), .B(B[217]), .CI(C[217]), .S(S[217]), 
        .CO(C[218]) );
  FA_2361 \FAINST[218].FA_  ( .A(A[218]), .B(B[218]), .CI(C[218]), .S(S[218]), 
        .CO(C[219]) );
  FA_2360 \FAINST[219].FA_  ( .A(A[219]), .B(B[219]), .CI(C[219]), .S(S[219]), 
        .CO(C[220]) );
  FA_2359 \FAINST[220].FA_  ( .A(A[220]), .B(B[220]), .CI(C[220]), .S(S[220]), 
        .CO(C[221]) );
  FA_2358 \FAINST[221].FA_  ( .A(A[221]), .B(B[221]), .CI(C[221]), .S(S[221]), 
        .CO(C[222]) );
  FA_2357 \FAINST[222].FA_  ( .A(A[222]), .B(B[222]), .CI(C[222]), .S(S[222]), 
        .CO(C[223]) );
  FA_2356 \FAINST[223].FA_  ( .A(A[223]), .B(B[223]), .CI(C[223]), .S(S[223]), 
        .CO(C[224]) );
  FA_2355 \FAINST[224].FA_  ( .A(A[224]), .B(B[224]), .CI(C[224]), .S(S[224]), 
        .CO(C[225]) );
  FA_2354 \FAINST[225].FA_  ( .A(A[225]), .B(B[225]), .CI(C[225]), .S(S[225]), 
        .CO(C[226]) );
  FA_2353 \FAINST[226].FA_  ( .A(A[226]), .B(B[226]), .CI(C[226]), .S(S[226]), 
        .CO(C[227]) );
  FA_2352 \FAINST[227].FA_  ( .A(A[227]), .B(B[227]), .CI(C[227]), .S(S[227]), 
        .CO(C[228]) );
  FA_2351 \FAINST[228].FA_  ( .A(A[228]), .B(B[228]), .CI(C[228]), .S(S[228]), 
        .CO(C[229]) );
  FA_2350 \FAINST[229].FA_  ( .A(A[229]), .B(B[229]), .CI(C[229]), .S(S[229]), 
        .CO(C[230]) );
  FA_2349 \FAINST[230].FA_  ( .A(A[230]), .B(B[230]), .CI(C[230]), .S(S[230]), 
        .CO(C[231]) );
  FA_2348 \FAINST[231].FA_  ( .A(A[231]), .B(B[231]), .CI(C[231]), .S(S[231]), 
        .CO(C[232]) );
  FA_2347 \FAINST[232].FA_  ( .A(A[232]), .B(B[232]), .CI(C[232]), .S(S[232]), 
        .CO(C[233]) );
  FA_2346 \FAINST[233].FA_  ( .A(A[233]), .B(B[233]), .CI(C[233]), .S(S[233]), 
        .CO(C[234]) );
  FA_2345 \FAINST[234].FA_  ( .A(A[234]), .B(B[234]), .CI(C[234]), .S(S[234]), 
        .CO(C[235]) );
  FA_2344 \FAINST[235].FA_  ( .A(A[235]), .B(B[235]), .CI(C[235]), .S(S[235]), 
        .CO(C[236]) );
  FA_2343 \FAINST[236].FA_  ( .A(A[236]), .B(B[236]), .CI(C[236]), .S(S[236]), 
        .CO(C[237]) );
  FA_2342 \FAINST[237].FA_  ( .A(A[237]), .B(B[237]), .CI(C[237]), .S(S[237]), 
        .CO(C[238]) );
  FA_2341 \FAINST[238].FA_  ( .A(A[238]), .B(B[238]), .CI(C[238]), .S(S[238]), 
        .CO(C[239]) );
  FA_2340 \FAINST[239].FA_  ( .A(A[239]), .B(B[239]), .CI(C[239]), .S(S[239]), 
        .CO(C[240]) );
  FA_2339 \FAINST[240].FA_  ( .A(A[240]), .B(B[240]), .CI(C[240]), .S(S[240]), 
        .CO(C[241]) );
  FA_2338 \FAINST[241].FA_  ( .A(A[241]), .B(B[241]), .CI(C[241]), .S(S[241]), 
        .CO(C[242]) );
  FA_2337 \FAINST[242].FA_  ( .A(A[242]), .B(B[242]), .CI(C[242]), .S(S[242]), 
        .CO(C[243]) );
  FA_2336 \FAINST[243].FA_  ( .A(A[243]), .B(B[243]), .CI(C[243]), .S(S[243]), 
        .CO(C[244]) );
  FA_2335 \FAINST[244].FA_  ( .A(A[244]), .B(B[244]), .CI(C[244]), .S(S[244]), 
        .CO(C[245]) );
  FA_2334 \FAINST[245].FA_  ( .A(A[245]), .B(B[245]), .CI(C[245]), .S(S[245]), 
        .CO(C[246]) );
  FA_2333 \FAINST[246].FA_  ( .A(A[246]), .B(B[246]), .CI(C[246]), .S(S[246]), 
        .CO(C[247]) );
  FA_2332 \FAINST[247].FA_  ( .A(A[247]), .B(B[247]), .CI(C[247]), .S(S[247]), 
        .CO(C[248]) );
  FA_2331 \FAINST[248].FA_  ( .A(A[248]), .B(B[248]), .CI(C[248]), .S(S[248]), 
        .CO(C[249]) );
  FA_2330 \FAINST[249].FA_  ( .A(A[249]), .B(B[249]), .CI(C[249]), .S(S[249]), 
        .CO(C[250]) );
  FA_2329 \FAINST[250].FA_  ( .A(A[250]), .B(B[250]), .CI(C[250]), .S(S[250]), 
        .CO(C[251]) );
  FA_2328 \FAINST[251].FA_  ( .A(A[251]), .B(B[251]), .CI(C[251]), .S(S[251]), 
        .CO(C[252]) );
  FA_2327 \FAINST[252].FA_  ( .A(A[252]), .B(B[252]), .CI(C[252]), .S(S[252]), 
        .CO(C[253]) );
  FA_2326 \FAINST[253].FA_  ( .A(A[253]), .B(B[253]), .CI(C[253]), .S(S[253]), 
        .CO(C[254]) );
  FA_2325 \FAINST[254].FA_  ( .A(A[254]), .B(B[254]), .CI(C[254]), .S(S[254]), 
        .CO(C[255]) );
  FA_2324 \FAINST[255].FA_  ( .A(A[255]), .B(B[255]), .CI(C[255]), .S(S[255]), 
        .CO(C[256]) );
  FA_2323 \FAINST[256].FA_  ( .A(A[256]), .B(1'b0), .CI(C[256]), .S(S[256]), 
        .CO(C[257]) );
  FA_2322 \FAINST[257].FA_  ( .A(A[257]), .B(1'b0), .CI(C[257]), .S(S[257]) );
endmodule


module FA_1548 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  AND U1 ( .A(CI), .B(B), .Z(CO) );
endmodule


module FA_1549 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  AND U1 ( .A(CI), .B(B), .Z(CO) );
endmodule


module FA_1550 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1551 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1552 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1553 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1554 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1555 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1556 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1557 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1558 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1559 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1560 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1561 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1562 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1563 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1564 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1565 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1566 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1567 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1568 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1569 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1570 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1571 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1572 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1573 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1574 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1575 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1576 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1577 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1578 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1579 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1580 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1581 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1582 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1583 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1584 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1585 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1586 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1587 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1588 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1589 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1590 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1591 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1592 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1593 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1594 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1595 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1596 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1597 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1598 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1599 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1600 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1601 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1602 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1603 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1604 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1605 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1606 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1607 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1608 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1609 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1610 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1611 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1612 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1613 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1614 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1615 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1616 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1617 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1618 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1619 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1620 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1621 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1622 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1623 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1624 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1625 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1626 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1627 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1628 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1629 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1630 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1631 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1632 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1633 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1634 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1635 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1636 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1637 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1638 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1639 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1640 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1641 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1642 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1643 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1644 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1645 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1646 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1647 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1648 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1649 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1650 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1651 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1652 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1653 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1654 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1655 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1656 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1657 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1658 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1659 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1660 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1661 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1662 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1663 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1664 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1665 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1666 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1667 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1668 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1669 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1670 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1671 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1672 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1673 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1674 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1675 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1676 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1677 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1678 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1679 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1680 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1681 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1682 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1683 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1684 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1685 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1686 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1687 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1688 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1689 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1690 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1691 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1692 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1693 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1694 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1695 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1696 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1697 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1698 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1699 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1700 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1701 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1702 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1703 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1704 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1705 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1706 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1707 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1708 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1709 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1710 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1711 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1712 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1713 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1714 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1715 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1716 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1717 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1718 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1719 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1720 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1721 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1722 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1723 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1724 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1725 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1726 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1727 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1728 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1729 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1730 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1731 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1732 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1733 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1734 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1735 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1736 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1737 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1738 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1739 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1740 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1741 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1742 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1743 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1744 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1745 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1746 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1747 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1748 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1749 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1750 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1751 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1752 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1753 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1754 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1755 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1756 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1757 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1758 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1759 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1760 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1761 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1762 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1763 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1764 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1765 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1766 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1767 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1768 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1769 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1770 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1771 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1772 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1773 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1774 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1775 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1776 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1777 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1778 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1779 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1780 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1781 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1782 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1783 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1784 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1785 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1786 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1787 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1788 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1789 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1790 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1791 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1792 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1793 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1794 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1795 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1796 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1797 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1798 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1799 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1800 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1801 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1802 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1803 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1804 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1805 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  OR U1 ( .A(B), .B(A), .Z(CO) );
endmodule


module COMP_N258_3 ( A, B, O );
  input [257:0] A;
  input [257:0] B;
  output O;
  wire   n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517;
  wire   [257:1] C;

  FA_1805 \FAINST[0].FA_  ( .A(A[0]), .B(n260), .CI(1'b1), .CO(C[1]) );
  FA_1804 \FAINST[1].FA_  ( .A(A[1]), .B(n261), .CI(C[1]), .CO(C[2]) );
  FA_1803 \FAINST[2].FA_  ( .A(A[2]), .B(n262), .CI(C[2]), .CO(C[3]) );
  FA_1802 \FAINST[3].FA_  ( .A(A[3]), .B(n263), .CI(C[3]), .CO(C[4]) );
  FA_1801 \FAINST[4].FA_  ( .A(A[4]), .B(n264), .CI(C[4]), .CO(C[5]) );
  FA_1800 \FAINST[5].FA_  ( .A(A[5]), .B(n265), .CI(C[5]), .CO(C[6]) );
  FA_1799 \FAINST[6].FA_  ( .A(A[6]), .B(n266), .CI(C[6]), .CO(C[7]) );
  FA_1798 \FAINST[7].FA_  ( .A(A[7]), .B(n267), .CI(C[7]), .CO(C[8]) );
  FA_1797 \FAINST[8].FA_  ( .A(A[8]), .B(n268), .CI(C[8]), .CO(C[9]) );
  FA_1796 \FAINST[9].FA_  ( .A(A[9]), .B(n269), .CI(C[9]), .CO(C[10]) );
  FA_1795 \FAINST[10].FA_  ( .A(A[10]), .B(n270), .CI(C[10]), .CO(C[11]) );
  FA_1794 \FAINST[11].FA_  ( .A(A[11]), .B(n271), .CI(C[11]), .CO(C[12]) );
  FA_1793 \FAINST[12].FA_  ( .A(A[12]), .B(n272), .CI(C[12]), .CO(C[13]) );
  FA_1792 \FAINST[13].FA_  ( .A(A[13]), .B(n273), .CI(C[13]), .CO(C[14]) );
  FA_1791 \FAINST[14].FA_  ( .A(A[14]), .B(n274), .CI(C[14]), .CO(C[15]) );
  FA_1790 \FAINST[15].FA_  ( .A(A[15]), .B(n275), .CI(C[15]), .CO(C[16]) );
  FA_1789 \FAINST[16].FA_  ( .A(A[16]), .B(n276), .CI(C[16]), .CO(C[17]) );
  FA_1788 \FAINST[17].FA_  ( .A(A[17]), .B(n277), .CI(C[17]), .CO(C[18]) );
  FA_1787 \FAINST[18].FA_  ( .A(A[18]), .B(n278), .CI(C[18]), .CO(C[19]) );
  FA_1786 \FAINST[19].FA_  ( .A(A[19]), .B(n279), .CI(C[19]), .CO(C[20]) );
  FA_1785 \FAINST[20].FA_  ( .A(A[20]), .B(n280), .CI(C[20]), .CO(C[21]) );
  FA_1784 \FAINST[21].FA_  ( .A(A[21]), .B(n281), .CI(C[21]), .CO(C[22]) );
  FA_1783 \FAINST[22].FA_  ( .A(A[22]), .B(n282), .CI(C[22]), .CO(C[23]) );
  FA_1782 \FAINST[23].FA_  ( .A(A[23]), .B(n283), .CI(C[23]), .CO(C[24]) );
  FA_1781 \FAINST[24].FA_  ( .A(A[24]), .B(n284), .CI(C[24]), .CO(C[25]) );
  FA_1780 \FAINST[25].FA_  ( .A(A[25]), .B(n285), .CI(C[25]), .CO(C[26]) );
  FA_1779 \FAINST[26].FA_  ( .A(A[26]), .B(n286), .CI(C[26]), .CO(C[27]) );
  FA_1778 \FAINST[27].FA_  ( .A(A[27]), .B(n287), .CI(C[27]), .CO(C[28]) );
  FA_1777 \FAINST[28].FA_  ( .A(A[28]), .B(n288), .CI(C[28]), .CO(C[29]) );
  FA_1776 \FAINST[29].FA_  ( .A(A[29]), .B(n289), .CI(C[29]), .CO(C[30]) );
  FA_1775 \FAINST[30].FA_  ( .A(A[30]), .B(n290), .CI(C[30]), .CO(C[31]) );
  FA_1774 \FAINST[31].FA_  ( .A(A[31]), .B(n291), .CI(C[31]), .CO(C[32]) );
  FA_1773 \FAINST[32].FA_  ( .A(A[32]), .B(n292), .CI(C[32]), .CO(C[33]) );
  FA_1772 \FAINST[33].FA_  ( .A(A[33]), .B(n293), .CI(C[33]), .CO(C[34]) );
  FA_1771 \FAINST[34].FA_  ( .A(A[34]), .B(n294), .CI(C[34]), .CO(C[35]) );
  FA_1770 \FAINST[35].FA_  ( .A(A[35]), .B(n295), .CI(C[35]), .CO(C[36]) );
  FA_1769 \FAINST[36].FA_  ( .A(A[36]), .B(n296), .CI(C[36]), .CO(C[37]) );
  FA_1768 \FAINST[37].FA_  ( .A(A[37]), .B(n297), .CI(C[37]), .CO(C[38]) );
  FA_1767 \FAINST[38].FA_  ( .A(A[38]), .B(n298), .CI(C[38]), .CO(C[39]) );
  FA_1766 \FAINST[39].FA_  ( .A(A[39]), .B(n299), .CI(C[39]), .CO(C[40]) );
  FA_1765 \FAINST[40].FA_  ( .A(A[40]), .B(n300), .CI(C[40]), .CO(C[41]) );
  FA_1764 \FAINST[41].FA_  ( .A(A[41]), .B(n301), .CI(C[41]), .CO(C[42]) );
  FA_1763 \FAINST[42].FA_  ( .A(A[42]), .B(n302), .CI(C[42]), .CO(C[43]) );
  FA_1762 \FAINST[43].FA_  ( .A(A[43]), .B(n303), .CI(C[43]), .CO(C[44]) );
  FA_1761 \FAINST[44].FA_  ( .A(A[44]), .B(n304), .CI(C[44]), .CO(C[45]) );
  FA_1760 \FAINST[45].FA_  ( .A(A[45]), .B(n305), .CI(C[45]), .CO(C[46]) );
  FA_1759 \FAINST[46].FA_  ( .A(A[46]), .B(n306), .CI(C[46]), .CO(C[47]) );
  FA_1758 \FAINST[47].FA_  ( .A(A[47]), .B(n307), .CI(C[47]), .CO(C[48]) );
  FA_1757 \FAINST[48].FA_  ( .A(A[48]), .B(n308), .CI(C[48]), .CO(C[49]) );
  FA_1756 \FAINST[49].FA_  ( .A(A[49]), .B(n309), .CI(C[49]), .CO(C[50]) );
  FA_1755 \FAINST[50].FA_  ( .A(A[50]), .B(n310), .CI(C[50]), .CO(C[51]) );
  FA_1754 \FAINST[51].FA_  ( .A(A[51]), .B(n311), .CI(C[51]), .CO(C[52]) );
  FA_1753 \FAINST[52].FA_  ( .A(A[52]), .B(n312), .CI(C[52]), .CO(C[53]) );
  FA_1752 \FAINST[53].FA_  ( .A(A[53]), .B(n313), .CI(C[53]), .CO(C[54]) );
  FA_1751 \FAINST[54].FA_  ( .A(A[54]), .B(n314), .CI(C[54]), .CO(C[55]) );
  FA_1750 \FAINST[55].FA_  ( .A(A[55]), .B(n315), .CI(C[55]), .CO(C[56]) );
  FA_1749 \FAINST[56].FA_  ( .A(A[56]), .B(n316), .CI(C[56]), .CO(C[57]) );
  FA_1748 \FAINST[57].FA_  ( .A(A[57]), .B(n317), .CI(C[57]), .CO(C[58]) );
  FA_1747 \FAINST[58].FA_  ( .A(A[58]), .B(n318), .CI(C[58]), .CO(C[59]) );
  FA_1746 \FAINST[59].FA_  ( .A(A[59]), .B(n319), .CI(C[59]), .CO(C[60]) );
  FA_1745 \FAINST[60].FA_  ( .A(A[60]), .B(n320), .CI(C[60]), .CO(C[61]) );
  FA_1744 \FAINST[61].FA_  ( .A(A[61]), .B(n321), .CI(C[61]), .CO(C[62]) );
  FA_1743 \FAINST[62].FA_  ( .A(A[62]), .B(n322), .CI(C[62]), .CO(C[63]) );
  FA_1742 \FAINST[63].FA_  ( .A(A[63]), .B(n323), .CI(C[63]), .CO(C[64]) );
  FA_1741 \FAINST[64].FA_  ( .A(A[64]), .B(n324), .CI(C[64]), .CO(C[65]) );
  FA_1740 \FAINST[65].FA_  ( .A(A[65]), .B(n325), .CI(C[65]), .CO(C[66]) );
  FA_1739 \FAINST[66].FA_  ( .A(A[66]), .B(n326), .CI(C[66]), .CO(C[67]) );
  FA_1738 \FAINST[67].FA_  ( .A(A[67]), .B(n327), .CI(C[67]), .CO(C[68]) );
  FA_1737 \FAINST[68].FA_  ( .A(A[68]), .B(n328), .CI(C[68]), .CO(C[69]) );
  FA_1736 \FAINST[69].FA_  ( .A(A[69]), .B(n329), .CI(C[69]), .CO(C[70]) );
  FA_1735 \FAINST[70].FA_  ( .A(A[70]), .B(n330), .CI(C[70]), .CO(C[71]) );
  FA_1734 \FAINST[71].FA_  ( .A(A[71]), .B(n331), .CI(C[71]), .CO(C[72]) );
  FA_1733 \FAINST[72].FA_  ( .A(A[72]), .B(n332), .CI(C[72]), .CO(C[73]) );
  FA_1732 \FAINST[73].FA_  ( .A(A[73]), .B(n333), .CI(C[73]), .CO(C[74]) );
  FA_1731 \FAINST[74].FA_  ( .A(A[74]), .B(n334), .CI(C[74]), .CO(C[75]) );
  FA_1730 \FAINST[75].FA_  ( .A(A[75]), .B(n335), .CI(C[75]), .CO(C[76]) );
  FA_1729 \FAINST[76].FA_  ( .A(A[76]), .B(n336), .CI(C[76]), .CO(C[77]) );
  FA_1728 \FAINST[77].FA_  ( .A(A[77]), .B(n337), .CI(C[77]), .CO(C[78]) );
  FA_1727 \FAINST[78].FA_  ( .A(A[78]), .B(n338), .CI(C[78]), .CO(C[79]) );
  FA_1726 \FAINST[79].FA_  ( .A(A[79]), .B(n339), .CI(C[79]), .CO(C[80]) );
  FA_1725 \FAINST[80].FA_  ( .A(A[80]), .B(n340), .CI(C[80]), .CO(C[81]) );
  FA_1724 \FAINST[81].FA_  ( .A(A[81]), .B(n341), .CI(C[81]), .CO(C[82]) );
  FA_1723 \FAINST[82].FA_  ( .A(A[82]), .B(n342), .CI(C[82]), .CO(C[83]) );
  FA_1722 \FAINST[83].FA_  ( .A(A[83]), .B(n343), .CI(C[83]), .CO(C[84]) );
  FA_1721 \FAINST[84].FA_  ( .A(A[84]), .B(n344), .CI(C[84]), .CO(C[85]) );
  FA_1720 \FAINST[85].FA_  ( .A(A[85]), .B(n345), .CI(C[85]), .CO(C[86]) );
  FA_1719 \FAINST[86].FA_  ( .A(A[86]), .B(n346), .CI(C[86]), .CO(C[87]) );
  FA_1718 \FAINST[87].FA_  ( .A(A[87]), .B(n347), .CI(C[87]), .CO(C[88]) );
  FA_1717 \FAINST[88].FA_  ( .A(A[88]), .B(n348), .CI(C[88]), .CO(C[89]) );
  FA_1716 \FAINST[89].FA_  ( .A(A[89]), .B(n349), .CI(C[89]), .CO(C[90]) );
  FA_1715 \FAINST[90].FA_  ( .A(A[90]), .B(n350), .CI(C[90]), .CO(C[91]) );
  FA_1714 \FAINST[91].FA_  ( .A(A[91]), .B(n351), .CI(C[91]), .CO(C[92]) );
  FA_1713 \FAINST[92].FA_  ( .A(A[92]), .B(n352), .CI(C[92]), .CO(C[93]) );
  FA_1712 \FAINST[93].FA_  ( .A(A[93]), .B(n353), .CI(C[93]), .CO(C[94]) );
  FA_1711 \FAINST[94].FA_  ( .A(A[94]), .B(n354), .CI(C[94]), .CO(C[95]) );
  FA_1710 \FAINST[95].FA_  ( .A(A[95]), .B(n355), .CI(C[95]), .CO(C[96]) );
  FA_1709 \FAINST[96].FA_  ( .A(A[96]), .B(n356), .CI(C[96]), .CO(C[97]) );
  FA_1708 \FAINST[97].FA_  ( .A(A[97]), .B(n357), .CI(C[97]), .CO(C[98]) );
  FA_1707 \FAINST[98].FA_  ( .A(A[98]), .B(n358), .CI(C[98]), .CO(C[99]) );
  FA_1706 \FAINST[99].FA_  ( .A(A[99]), .B(n359), .CI(C[99]), .CO(C[100]) );
  FA_1705 \FAINST[100].FA_  ( .A(A[100]), .B(n360), .CI(C[100]), .CO(C[101])
         );
  FA_1704 \FAINST[101].FA_  ( .A(A[101]), .B(n361), .CI(C[101]), .CO(C[102])
         );
  FA_1703 \FAINST[102].FA_  ( .A(A[102]), .B(n362), .CI(C[102]), .CO(C[103])
         );
  FA_1702 \FAINST[103].FA_  ( .A(A[103]), .B(n363), .CI(C[103]), .CO(C[104])
         );
  FA_1701 \FAINST[104].FA_  ( .A(A[104]), .B(n364), .CI(C[104]), .CO(C[105])
         );
  FA_1700 \FAINST[105].FA_  ( .A(A[105]), .B(n365), .CI(C[105]), .CO(C[106])
         );
  FA_1699 \FAINST[106].FA_  ( .A(A[106]), .B(n366), .CI(C[106]), .CO(C[107])
         );
  FA_1698 \FAINST[107].FA_  ( .A(A[107]), .B(n367), .CI(C[107]), .CO(C[108])
         );
  FA_1697 \FAINST[108].FA_  ( .A(A[108]), .B(n368), .CI(C[108]), .CO(C[109])
         );
  FA_1696 \FAINST[109].FA_  ( .A(A[109]), .B(n369), .CI(C[109]), .CO(C[110])
         );
  FA_1695 \FAINST[110].FA_  ( .A(A[110]), .B(n370), .CI(C[110]), .CO(C[111])
         );
  FA_1694 \FAINST[111].FA_  ( .A(A[111]), .B(n371), .CI(C[111]), .CO(C[112])
         );
  FA_1693 \FAINST[112].FA_  ( .A(A[112]), .B(n372), .CI(C[112]), .CO(C[113])
         );
  FA_1692 \FAINST[113].FA_  ( .A(A[113]), .B(n373), .CI(C[113]), .CO(C[114])
         );
  FA_1691 \FAINST[114].FA_  ( .A(A[114]), .B(n374), .CI(C[114]), .CO(C[115])
         );
  FA_1690 \FAINST[115].FA_  ( .A(A[115]), .B(n375), .CI(C[115]), .CO(C[116])
         );
  FA_1689 \FAINST[116].FA_  ( .A(A[116]), .B(n376), .CI(C[116]), .CO(C[117])
         );
  FA_1688 \FAINST[117].FA_  ( .A(A[117]), .B(n377), .CI(C[117]), .CO(C[118])
         );
  FA_1687 \FAINST[118].FA_  ( .A(A[118]), .B(n378), .CI(C[118]), .CO(C[119])
         );
  FA_1686 \FAINST[119].FA_  ( .A(A[119]), .B(n379), .CI(C[119]), .CO(C[120])
         );
  FA_1685 \FAINST[120].FA_  ( .A(A[120]), .B(n380), .CI(C[120]), .CO(C[121])
         );
  FA_1684 \FAINST[121].FA_  ( .A(A[121]), .B(n381), .CI(C[121]), .CO(C[122])
         );
  FA_1683 \FAINST[122].FA_  ( .A(A[122]), .B(n382), .CI(C[122]), .CO(C[123])
         );
  FA_1682 \FAINST[123].FA_  ( .A(A[123]), .B(n383), .CI(C[123]), .CO(C[124])
         );
  FA_1681 \FAINST[124].FA_  ( .A(A[124]), .B(n384), .CI(C[124]), .CO(C[125])
         );
  FA_1680 \FAINST[125].FA_  ( .A(A[125]), .B(n385), .CI(C[125]), .CO(C[126])
         );
  FA_1679 \FAINST[126].FA_  ( .A(A[126]), .B(n386), .CI(C[126]), .CO(C[127])
         );
  FA_1678 \FAINST[127].FA_  ( .A(A[127]), .B(n387), .CI(C[127]), .CO(C[128])
         );
  FA_1677 \FAINST[128].FA_  ( .A(A[128]), .B(n388), .CI(C[128]), .CO(C[129])
         );
  FA_1676 \FAINST[129].FA_  ( .A(A[129]), .B(n389), .CI(C[129]), .CO(C[130])
         );
  FA_1675 \FAINST[130].FA_  ( .A(A[130]), .B(n390), .CI(C[130]), .CO(C[131])
         );
  FA_1674 \FAINST[131].FA_  ( .A(A[131]), .B(n391), .CI(C[131]), .CO(C[132])
         );
  FA_1673 \FAINST[132].FA_  ( .A(A[132]), .B(n392), .CI(C[132]), .CO(C[133])
         );
  FA_1672 \FAINST[133].FA_  ( .A(A[133]), .B(n393), .CI(C[133]), .CO(C[134])
         );
  FA_1671 \FAINST[134].FA_  ( .A(A[134]), .B(n394), .CI(C[134]), .CO(C[135])
         );
  FA_1670 \FAINST[135].FA_  ( .A(A[135]), .B(n395), .CI(C[135]), .CO(C[136])
         );
  FA_1669 \FAINST[136].FA_  ( .A(A[136]), .B(n396), .CI(C[136]), .CO(C[137])
         );
  FA_1668 \FAINST[137].FA_  ( .A(A[137]), .B(n397), .CI(C[137]), .CO(C[138])
         );
  FA_1667 \FAINST[138].FA_  ( .A(A[138]), .B(n398), .CI(C[138]), .CO(C[139])
         );
  FA_1666 \FAINST[139].FA_  ( .A(A[139]), .B(n399), .CI(C[139]), .CO(C[140])
         );
  FA_1665 \FAINST[140].FA_  ( .A(A[140]), .B(n400), .CI(C[140]), .CO(C[141])
         );
  FA_1664 \FAINST[141].FA_  ( .A(A[141]), .B(n401), .CI(C[141]), .CO(C[142])
         );
  FA_1663 \FAINST[142].FA_  ( .A(A[142]), .B(n402), .CI(C[142]), .CO(C[143])
         );
  FA_1662 \FAINST[143].FA_  ( .A(A[143]), .B(n403), .CI(C[143]), .CO(C[144])
         );
  FA_1661 \FAINST[144].FA_  ( .A(A[144]), .B(n404), .CI(C[144]), .CO(C[145])
         );
  FA_1660 \FAINST[145].FA_  ( .A(A[145]), .B(n405), .CI(C[145]), .CO(C[146])
         );
  FA_1659 \FAINST[146].FA_  ( .A(A[146]), .B(n406), .CI(C[146]), .CO(C[147])
         );
  FA_1658 \FAINST[147].FA_  ( .A(A[147]), .B(n407), .CI(C[147]), .CO(C[148])
         );
  FA_1657 \FAINST[148].FA_  ( .A(A[148]), .B(n408), .CI(C[148]), .CO(C[149])
         );
  FA_1656 \FAINST[149].FA_  ( .A(A[149]), .B(n409), .CI(C[149]), .CO(C[150])
         );
  FA_1655 \FAINST[150].FA_  ( .A(A[150]), .B(n410), .CI(C[150]), .CO(C[151])
         );
  FA_1654 \FAINST[151].FA_  ( .A(A[151]), .B(n411), .CI(C[151]), .CO(C[152])
         );
  FA_1653 \FAINST[152].FA_  ( .A(A[152]), .B(n412), .CI(C[152]), .CO(C[153])
         );
  FA_1652 \FAINST[153].FA_  ( .A(A[153]), .B(n413), .CI(C[153]), .CO(C[154])
         );
  FA_1651 \FAINST[154].FA_  ( .A(A[154]), .B(n414), .CI(C[154]), .CO(C[155])
         );
  FA_1650 \FAINST[155].FA_  ( .A(A[155]), .B(n415), .CI(C[155]), .CO(C[156])
         );
  FA_1649 \FAINST[156].FA_  ( .A(A[156]), .B(n416), .CI(C[156]), .CO(C[157])
         );
  FA_1648 \FAINST[157].FA_  ( .A(A[157]), .B(n417), .CI(C[157]), .CO(C[158])
         );
  FA_1647 \FAINST[158].FA_  ( .A(A[158]), .B(n418), .CI(C[158]), .CO(C[159])
         );
  FA_1646 \FAINST[159].FA_  ( .A(A[159]), .B(n419), .CI(C[159]), .CO(C[160])
         );
  FA_1645 \FAINST[160].FA_  ( .A(A[160]), .B(n420), .CI(C[160]), .CO(C[161])
         );
  FA_1644 \FAINST[161].FA_  ( .A(A[161]), .B(n421), .CI(C[161]), .CO(C[162])
         );
  FA_1643 \FAINST[162].FA_  ( .A(A[162]), .B(n422), .CI(C[162]), .CO(C[163])
         );
  FA_1642 \FAINST[163].FA_  ( .A(A[163]), .B(n423), .CI(C[163]), .CO(C[164])
         );
  FA_1641 \FAINST[164].FA_  ( .A(A[164]), .B(n424), .CI(C[164]), .CO(C[165])
         );
  FA_1640 \FAINST[165].FA_  ( .A(A[165]), .B(n425), .CI(C[165]), .CO(C[166])
         );
  FA_1639 \FAINST[166].FA_  ( .A(A[166]), .B(n426), .CI(C[166]), .CO(C[167])
         );
  FA_1638 \FAINST[167].FA_  ( .A(A[167]), .B(n427), .CI(C[167]), .CO(C[168])
         );
  FA_1637 \FAINST[168].FA_  ( .A(A[168]), .B(n428), .CI(C[168]), .CO(C[169])
         );
  FA_1636 \FAINST[169].FA_  ( .A(A[169]), .B(n429), .CI(C[169]), .CO(C[170])
         );
  FA_1635 \FAINST[170].FA_  ( .A(A[170]), .B(n430), .CI(C[170]), .CO(C[171])
         );
  FA_1634 \FAINST[171].FA_  ( .A(A[171]), .B(n431), .CI(C[171]), .CO(C[172])
         );
  FA_1633 \FAINST[172].FA_  ( .A(A[172]), .B(n432), .CI(C[172]), .CO(C[173])
         );
  FA_1632 \FAINST[173].FA_  ( .A(A[173]), .B(n433), .CI(C[173]), .CO(C[174])
         );
  FA_1631 \FAINST[174].FA_  ( .A(A[174]), .B(n434), .CI(C[174]), .CO(C[175])
         );
  FA_1630 \FAINST[175].FA_  ( .A(A[175]), .B(n435), .CI(C[175]), .CO(C[176])
         );
  FA_1629 \FAINST[176].FA_  ( .A(A[176]), .B(n436), .CI(C[176]), .CO(C[177])
         );
  FA_1628 \FAINST[177].FA_  ( .A(A[177]), .B(n437), .CI(C[177]), .CO(C[178])
         );
  FA_1627 \FAINST[178].FA_  ( .A(A[178]), .B(n438), .CI(C[178]), .CO(C[179])
         );
  FA_1626 \FAINST[179].FA_  ( .A(A[179]), .B(n439), .CI(C[179]), .CO(C[180])
         );
  FA_1625 \FAINST[180].FA_  ( .A(A[180]), .B(n440), .CI(C[180]), .CO(C[181])
         );
  FA_1624 \FAINST[181].FA_  ( .A(A[181]), .B(n441), .CI(C[181]), .CO(C[182])
         );
  FA_1623 \FAINST[182].FA_  ( .A(A[182]), .B(n442), .CI(C[182]), .CO(C[183])
         );
  FA_1622 \FAINST[183].FA_  ( .A(A[183]), .B(n443), .CI(C[183]), .CO(C[184])
         );
  FA_1621 \FAINST[184].FA_  ( .A(A[184]), .B(n444), .CI(C[184]), .CO(C[185])
         );
  FA_1620 \FAINST[185].FA_  ( .A(A[185]), .B(n445), .CI(C[185]), .CO(C[186])
         );
  FA_1619 \FAINST[186].FA_  ( .A(A[186]), .B(n446), .CI(C[186]), .CO(C[187])
         );
  FA_1618 \FAINST[187].FA_  ( .A(A[187]), .B(n447), .CI(C[187]), .CO(C[188])
         );
  FA_1617 \FAINST[188].FA_  ( .A(A[188]), .B(n448), .CI(C[188]), .CO(C[189])
         );
  FA_1616 \FAINST[189].FA_  ( .A(A[189]), .B(n449), .CI(C[189]), .CO(C[190])
         );
  FA_1615 \FAINST[190].FA_  ( .A(A[190]), .B(n450), .CI(C[190]), .CO(C[191])
         );
  FA_1614 \FAINST[191].FA_  ( .A(A[191]), .B(n451), .CI(C[191]), .CO(C[192])
         );
  FA_1613 \FAINST[192].FA_  ( .A(A[192]), .B(n452), .CI(C[192]), .CO(C[193])
         );
  FA_1612 \FAINST[193].FA_  ( .A(A[193]), .B(n453), .CI(C[193]), .CO(C[194])
         );
  FA_1611 \FAINST[194].FA_  ( .A(A[194]), .B(n454), .CI(C[194]), .CO(C[195])
         );
  FA_1610 \FAINST[195].FA_  ( .A(A[195]), .B(n455), .CI(C[195]), .CO(C[196])
         );
  FA_1609 \FAINST[196].FA_  ( .A(A[196]), .B(n456), .CI(C[196]), .CO(C[197])
         );
  FA_1608 \FAINST[197].FA_  ( .A(A[197]), .B(n457), .CI(C[197]), .CO(C[198])
         );
  FA_1607 \FAINST[198].FA_  ( .A(A[198]), .B(n458), .CI(C[198]), .CO(C[199])
         );
  FA_1606 \FAINST[199].FA_  ( .A(A[199]), .B(n459), .CI(C[199]), .CO(C[200])
         );
  FA_1605 \FAINST[200].FA_  ( .A(A[200]), .B(n460), .CI(C[200]), .CO(C[201])
         );
  FA_1604 \FAINST[201].FA_  ( .A(A[201]), .B(n461), .CI(C[201]), .CO(C[202])
         );
  FA_1603 \FAINST[202].FA_  ( .A(A[202]), .B(n462), .CI(C[202]), .CO(C[203])
         );
  FA_1602 \FAINST[203].FA_  ( .A(A[203]), .B(n463), .CI(C[203]), .CO(C[204])
         );
  FA_1601 \FAINST[204].FA_  ( .A(A[204]), .B(n464), .CI(C[204]), .CO(C[205])
         );
  FA_1600 \FAINST[205].FA_  ( .A(A[205]), .B(n465), .CI(C[205]), .CO(C[206])
         );
  FA_1599 \FAINST[206].FA_  ( .A(A[206]), .B(n466), .CI(C[206]), .CO(C[207])
         );
  FA_1598 \FAINST[207].FA_  ( .A(A[207]), .B(n467), .CI(C[207]), .CO(C[208])
         );
  FA_1597 \FAINST[208].FA_  ( .A(A[208]), .B(n468), .CI(C[208]), .CO(C[209])
         );
  FA_1596 \FAINST[209].FA_  ( .A(A[209]), .B(n469), .CI(C[209]), .CO(C[210])
         );
  FA_1595 \FAINST[210].FA_  ( .A(A[210]), .B(n470), .CI(C[210]), .CO(C[211])
         );
  FA_1594 \FAINST[211].FA_  ( .A(A[211]), .B(n471), .CI(C[211]), .CO(C[212])
         );
  FA_1593 \FAINST[212].FA_  ( .A(A[212]), .B(n472), .CI(C[212]), .CO(C[213])
         );
  FA_1592 \FAINST[213].FA_  ( .A(A[213]), .B(n473), .CI(C[213]), .CO(C[214])
         );
  FA_1591 \FAINST[214].FA_  ( .A(A[214]), .B(n474), .CI(C[214]), .CO(C[215])
         );
  FA_1590 \FAINST[215].FA_  ( .A(A[215]), .B(n475), .CI(C[215]), .CO(C[216])
         );
  FA_1589 \FAINST[216].FA_  ( .A(A[216]), .B(n476), .CI(C[216]), .CO(C[217])
         );
  FA_1588 \FAINST[217].FA_  ( .A(A[217]), .B(n477), .CI(C[217]), .CO(C[218])
         );
  FA_1587 \FAINST[218].FA_  ( .A(A[218]), .B(n478), .CI(C[218]), .CO(C[219])
         );
  FA_1586 \FAINST[219].FA_  ( .A(A[219]), .B(n479), .CI(C[219]), .CO(C[220])
         );
  FA_1585 \FAINST[220].FA_  ( .A(A[220]), .B(n480), .CI(C[220]), .CO(C[221])
         );
  FA_1584 \FAINST[221].FA_  ( .A(A[221]), .B(n481), .CI(C[221]), .CO(C[222])
         );
  FA_1583 \FAINST[222].FA_  ( .A(A[222]), .B(n482), .CI(C[222]), .CO(C[223])
         );
  FA_1582 \FAINST[223].FA_  ( .A(A[223]), .B(n483), .CI(C[223]), .CO(C[224])
         );
  FA_1581 \FAINST[224].FA_  ( .A(A[224]), .B(n484), .CI(C[224]), .CO(C[225])
         );
  FA_1580 \FAINST[225].FA_  ( .A(A[225]), .B(n485), .CI(C[225]), .CO(C[226])
         );
  FA_1579 \FAINST[226].FA_  ( .A(A[226]), .B(n486), .CI(C[226]), .CO(C[227])
         );
  FA_1578 \FAINST[227].FA_  ( .A(A[227]), .B(n487), .CI(C[227]), .CO(C[228])
         );
  FA_1577 \FAINST[228].FA_  ( .A(A[228]), .B(n488), .CI(C[228]), .CO(C[229])
         );
  FA_1576 \FAINST[229].FA_  ( .A(A[229]), .B(n489), .CI(C[229]), .CO(C[230])
         );
  FA_1575 \FAINST[230].FA_  ( .A(A[230]), .B(n490), .CI(C[230]), .CO(C[231])
         );
  FA_1574 \FAINST[231].FA_  ( .A(A[231]), .B(n491), .CI(C[231]), .CO(C[232])
         );
  FA_1573 \FAINST[232].FA_  ( .A(A[232]), .B(n492), .CI(C[232]), .CO(C[233])
         );
  FA_1572 \FAINST[233].FA_  ( .A(A[233]), .B(n493), .CI(C[233]), .CO(C[234])
         );
  FA_1571 \FAINST[234].FA_  ( .A(A[234]), .B(n494), .CI(C[234]), .CO(C[235])
         );
  FA_1570 \FAINST[235].FA_  ( .A(A[235]), .B(n495), .CI(C[235]), .CO(C[236])
         );
  FA_1569 \FAINST[236].FA_  ( .A(A[236]), .B(n496), .CI(C[236]), .CO(C[237])
         );
  FA_1568 \FAINST[237].FA_  ( .A(A[237]), .B(n497), .CI(C[237]), .CO(C[238])
         );
  FA_1567 \FAINST[238].FA_  ( .A(A[238]), .B(n498), .CI(C[238]), .CO(C[239])
         );
  FA_1566 \FAINST[239].FA_  ( .A(A[239]), .B(n499), .CI(C[239]), .CO(C[240])
         );
  FA_1565 \FAINST[240].FA_  ( .A(A[240]), .B(n500), .CI(C[240]), .CO(C[241])
         );
  FA_1564 \FAINST[241].FA_  ( .A(A[241]), .B(n501), .CI(C[241]), .CO(C[242])
         );
  FA_1563 \FAINST[242].FA_  ( .A(A[242]), .B(n502), .CI(C[242]), .CO(C[243])
         );
  FA_1562 \FAINST[243].FA_  ( .A(A[243]), .B(n503), .CI(C[243]), .CO(C[244])
         );
  FA_1561 \FAINST[244].FA_  ( .A(A[244]), .B(n504), .CI(C[244]), .CO(C[245])
         );
  FA_1560 \FAINST[245].FA_  ( .A(A[245]), .B(n505), .CI(C[245]), .CO(C[246])
         );
  FA_1559 \FAINST[246].FA_  ( .A(A[246]), .B(n506), .CI(C[246]), .CO(C[247])
         );
  FA_1558 \FAINST[247].FA_  ( .A(A[247]), .B(n507), .CI(C[247]), .CO(C[248])
         );
  FA_1557 \FAINST[248].FA_  ( .A(A[248]), .B(n508), .CI(C[248]), .CO(C[249])
         );
  FA_1556 \FAINST[249].FA_  ( .A(A[249]), .B(n509), .CI(C[249]), .CO(C[250])
         );
  FA_1555 \FAINST[250].FA_  ( .A(A[250]), .B(n510), .CI(C[250]), .CO(C[251])
         );
  FA_1554 \FAINST[251].FA_  ( .A(A[251]), .B(n511), .CI(C[251]), .CO(C[252])
         );
  FA_1553 \FAINST[252].FA_  ( .A(A[252]), .B(n512), .CI(C[252]), .CO(C[253])
         );
  FA_1552 \FAINST[253].FA_  ( .A(A[253]), .B(n513), .CI(C[253]), .CO(C[254])
         );
  FA_1551 \FAINST[254].FA_  ( .A(A[254]), .B(n514), .CI(C[254]), .CO(C[255])
         );
  FA_1550 \FAINST[255].FA_  ( .A(A[255]), .B(n515), .CI(C[255]), .CO(C[256])
         );
  FA_1549 \FAINST[256].FA_  ( .A(1'b0), .B(n516), .CI(C[256]), .CO(C[257]) );
  FA_1548 \FAINST[257].FA_  ( .A(1'b0), .B(n517), .CI(C[257]), .CO(O) );
  IV U2 ( .A(B[159]), .Z(n419) );
  IV U3 ( .A(B[160]), .Z(n420) );
  IV U4 ( .A(B[161]), .Z(n421) );
  IV U5 ( .A(B[162]), .Z(n422) );
  IV U6 ( .A(B[163]), .Z(n423) );
  IV U7 ( .A(B[164]), .Z(n424) );
  IV U8 ( .A(B[165]), .Z(n425) );
  IV U9 ( .A(B[166]), .Z(n426) );
  IV U10 ( .A(B[167]), .Z(n427) );
  IV U11 ( .A(B[168]), .Z(n428) );
  IV U12 ( .A(B[249]), .Z(n509) );
  IV U13 ( .A(B[169]), .Z(n429) );
  IV U14 ( .A(B[170]), .Z(n430) );
  IV U15 ( .A(B[171]), .Z(n431) );
  IV U16 ( .A(B[172]), .Z(n432) );
  IV U17 ( .A(B[173]), .Z(n433) );
  IV U18 ( .A(B[174]), .Z(n434) );
  IV U19 ( .A(B[175]), .Z(n435) );
  IV U20 ( .A(B[176]), .Z(n436) );
  IV U21 ( .A(B[177]), .Z(n437) );
  IV U22 ( .A(B[178]), .Z(n438) );
  IV U23 ( .A(B[250]), .Z(n510) );
  IV U24 ( .A(B[179]), .Z(n439) );
  IV U25 ( .A(B[180]), .Z(n440) );
  IV U26 ( .A(B[181]), .Z(n441) );
  IV U27 ( .A(B[182]), .Z(n442) );
  IV U28 ( .A(B[183]), .Z(n443) );
  IV U29 ( .A(B[184]), .Z(n444) );
  IV U30 ( .A(B[185]), .Z(n445) );
  IV U31 ( .A(B[186]), .Z(n446) );
  IV U32 ( .A(B[187]), .Z(n447) );
  IV U33 ( .A(B[188]), .Z(n448) );
  IV U34 ( .A(B[251]), .Z(n511) );
  IV U35 ( .A(B[189]), .Z(n449) );
  IV U36 ( .A(B[190]), .Z(n450) );
  IV U37 ( .A(B[191]), .Z(n451) );
  IV U38 ( .A(B[192]), .Z(n452) );
  IV U39 ( .A(B[193]), .Z(n453) );
  IV U40 ( .A(B[194]), .Z(n454) );
  IV U41 ( .A(B[195]), .Z(n455) );
  IV U42 ( .A(B[196]), .Z(n456) );
  IV U43 ( .A(B[197]), .Z(n457) );
  IV U44 ( .A(B[198]), .Z(n458) );
  IV U45 ( .A(B[252]), .Z(n512) );
  IV U46 ( .A(B[199]), .Z(n459) );
  IV U47 ( .A(B[200]), .Z(n460) );
  IV U48 ( .A(B[201]), .Z(n461) );
  IV U49 ( .A(B[202]), .Z(n462) );
  IV U50 ( .A(B[203]), .Z(n463) );
  IV U51 ( .A(B[204]), .Z(n464) );
  IV U52 ( .A(B[205]), .Z(n465) );
  IV U53 ( .A(B[206]), .Z(n466) );
  IV U54 ( .A(B[207]), .Z(n467) );
  IV U55 ( .A(B[208]), .Z(n468) );
  IV U56 ( .A(B[253]), .Z(n513) );
  IV U57 ( .A(B[209]), .Z(n469) );
  IV U58 ( .A(B[210]), .Z(n470) );
  IV U59 ( .A(B[211]), .Z(n471) );
  IV U60 ( .A(B[212]), .Z(n472) );
  IV U61 ( .A(B[213]), .Z(n473) );
  IV U62 ( .A(B[214]), .Z(n474) );
  IV U63 ( .A(B[215]), .Z(n475) );
  IV U64 ( .A(B[216]), .Z(n476) );
  IV U65 ( .A(B[217]), .Z(n477) );
  IV U66 ( .A(B[218]), .Z(n478) );
  IV U67 ( .A(B[254]), .Z(n514) );
  IV U68 ( .A(B[219]), .Z(n479) );
  IV U69 ( .A(B[220]), .Z(n480) );
  IV U70 ( .A(B[221]), .Z(n481) );
  IV U71 ( .A(B[222]), .Z(n482) );
  IV U72 ( .A(B[223]), .Z(n483) );
  IV U73 ( .A(B[224]), .Z(n484) );
  IV U74 ( .A(B[225]), .Z(n485) );
  IV U75 ( .A(B[226]), .Z(n486) );
  IV U76 ( .A(B[227]), .Z(n487) );
  IV U77 ( .A(B[228]), .Z(n488) );
  IV U78 ( .A(B[255]), .Z(n515) );
  IV U79 ( .A(B[229]), .Z(n489) );
  IV U80 ( .A(B[230]), .Z(n490) );
  IV U81 ( .A(B[231]), .Z(n491) );
  IV U82 ( .A(B[232]), .Z(n492) );
  IV U83 ( .A(B[0]), .Z(n260) );
  IV U84 ( .A(B[1]), .Z(n261) );
  IV U85 ( .A(B[2]), .Z(n262) );
  IV U86 ( .A(B[3]), .Z(n263) );
  IV U87 ( .A(B[4]), .Z(n264) );
  IV U88 ( .A(B[5]), .Z(n265) );
  IV U89 ( .A(B[6]), .Z(n266) );
  IV U90 ( .A(B[7]), .Z(n267) );
  IV U91 ( .A(B[8]), .Z(n268) );
  IV U92 ( .A(B[233]), .Z(n493) );
  IV U93 ( .A(B[9]), .Z(n269) );
  IV U94 ( .A(B[10]), .Z(n270) );
  IV U95 ( .A(B[11]), .Z(n271) );
  IV U96 ( .A(B[12]), .Z(n272) );
  IV U97 ( .A(B[13]), .Z(n273) );
  IV U98 ( .A(B[14]), .Z(n274) );
  IV U99 ( .A(B[15]), .Z(n275) );
  IV U100 ( .A(B[16]), .Z(n276) );
  IV U101 ( .A(B[17]), .Z(n277) );
  IV U102 ( .A(B[18]), .Z(n278) );
  IV U103 ( .A(B[234]), .Z(n494) );
  IV U104 ( .A(B[19]), .Z(n279) );
  IV U105 ( .A(B[20]), .Z(n280) );
  IV U106 ( .A(B[21]), .Z(n281) );
  IV U107 ( .A(B[22]), .Z(n282) );
  IV U108 ( .A(B[23]), .Z(n283) );
  IV U109 ( .A(B[24]), .Z(n284) );
  IV U110 ( .A(B[25]), .Z(n285) );
  IV U111 ( .A(B[26]), .Z(n286) );
  IV U112 ( .A(B[27]), .Z(n287) );
  IV U113 ( .A(B[28]), .Z(n288) );
  IV U114 ( .A(B[235]), .Z(n495) );
  IV U115 ( .A(B[29]), .Z(n289) );
  IV U116 ( .A(B[30]), .Z(n290) );
  IV U117 ( .A(B[31]), .Z(n291) );
  IV U118 ( .A(B[32]), .Z(n292) );
  IV U119 ( .A(B[33]), .Z(n293) );
  IV U120 ( .A(B[34]), .Z(n294) );
  IV U121 ( .A(B[35]), .Z(n295) );
  IV U122 ( .A(B[36]), .Z(n296) );
  IV U123 ( .A(B[37]), .Z(n297) );
  IV U124 ( .A(B[38]), .Z(n298) );
  IV U125 ( .A(B[236]), .Z(n496) );
  IV U126 ( .A(B[39]), .Z(n299) );
  IV U127 ( .A(B[40]), .Z(n300) );
  IV U128 ( .A(B[41]), .Z(n301) );
  IV U129 ( .A(B[42]), .Z(n302) );
  IV U130 ( .A(B[43]), .Z(n303) );
  IV U131 ( .A(B[44]), .Z(n304) );
  IV U132 ( .A(B[45]), .Z(n305) );
  IV U133 ( .A(B[46]), .Z(n306) );
  IV U134 ( .A(B[47]), .Z(n307) );
  IV U135 ( .A(B[48]), .Z(n308) );
  IV U136 ( .A(B[237]), .Z(n497) );
  IV U137 ( .A(B[49]), .Z(n309) );
  IV U138 ( .A(B[50]), .Z(n310) );
  IV U139 ( .A(B[51]), .Z(n311) );
  IV U140 ( .A(B[52]), .Z(n312) );
  IV U141 ( .A(B[53]), .Z(n313) );
  IV U142 ( .A(B[54]), .Z(n314) );
  IV U143 ( .A(B[55]), .Z(n315) );
  IV U144 ( .A(B[56]), .Z(n316) );
  IV U145 ( .A(B[57]), .Z(n317) );
  IV U146 ( .A(B[58]), .Z(n318) );
  IV U147 ( .A(B[238]), .Z(n498) );
  IV U148 ( .A(B[256]), .Z(n516) );
  IV U149 ( .A(B[59]), .Z(n319) );
  IV U150 ( .A(B[60]), .Z(n320) );
  IV U151 ( .A(B[61]), .Z(n321) );
  IV U152 ( .A(B[62]), .Z(n322) );
  IV U153 ( .A(B[63]), .Z(n323) );
  IV U154 ( .A(B[64]), .Z(n324) );
  IV U155 ( .A(B[65]), .Z(n325) );
  IV U156 ( .A(B[66]), .Z(n326) );
  IV U157 ( .A(B[67]), .Z(n327) );
  IV U158 ( .A(B[68]), .Z(n328) );
  IV U159 ( .A(B[239]), .Z(n499) );
  IV U160 ( .A(B[69]), .Z(n329) );
  IV U161 ( .A(B[70]), .Z(n330) );
  IV U162 ( .A(B[71]), .Z(n331) );
  IV U163 ( .A(B[72]), .Z(n332) );
  IV U164 ( .A(B[73]), .Z(n333) );
  IV U165 ( .A(B[74]), .Z(n334) );
  IV U166 ( .A(B[75]), .Z(n335) );
  IV U167 ( .A(B[76]), .Z(n336) );
  IV U168 ( .A(B[77]), .Z(n337) );
  IV U169 ( .A(B[78]), .Z(n338) );
  IV U170 ( .A(B[240]), .Z(n500) );
  IV U171 ( .A(B[79]), .Z(n339) );
  IV U172 ( .A(B[80]), .Z(n340) );
  IV U173 ( .A(B[81]), .Z(n341) );
  IV U174 ( .A(B[82]), .Z(n342) );
  IV U175 ( .A(B[83]), .Z(n343) );
  IV U176 ( .A(B[84]), .Z(n344) );
  IV U177 ( .A(B[85]), .Z(n345) );
  IV U178 ( .A(B[86]), .Z(n346) );
  IV U179 ( .A(B[87]), .Z(n347) );
  IV U180 ( .A(B[88]), .Z(n348) );
  IV U181 ( .A(B[241]), .Z(n501) );
  IV U182 ( .A(B[89]), .Z(n349) );
  IV U183 ( .A(B[90]), .Z(n350) );
  IV U184 ( .A(B[91]), .Z(n351) );
  IV U185 ( .A(B[92]), .Z(n352) );
  IV U186 ( .A(B[93]), .Z(n353) );
  IV U187 ( .A(B[94]), .Z(n354) );
  IV U188 ( .A(B[95]), .Z(n355) );
  IV U189 ( .A(B[96]), .Z(n356) );
  IV U190 ( .A(B[97]), .Z(n357) );
  IV U191 ( .A(B[98]), .Z(n358) );
  IV U192 ( .A(B[242]), .Z(n502) );
  IV U193 ( .A(B[99]), .Z(n359) );
  IV U194 ( .A(B[100]), .Z(n360) );
  IV U195 ( .A(B[101]), .Z(n361) );
  IV U196 ( .A(B[102]), .Z(n362) );
  IV U197 ( .A(B[103]), .Z(n363) );
  IV U198 ( .A(B[104]), .Z(n364) );
  IV U199 ( .A(B[105]), .Z(n365) );
  IV U200 ( .A(B[106]), .Z(n366) );
  IV U201 ( .A(B[107]), .Z(n367) );
  IV U202 ( .A(B[108]), .Z(n368) );
  IV U203 ( .A(B[243]), .Z(n503) );
  IV U204 ( .A(B[109]), .Z(n369) );
  IV U205 ( .A(B[110]), .Z(n370) );
  IV U206 ( .A(B[111]), .Z(n371) );
  IV U207 ( .A(B[112]), .Z(n372) );
  IV U208 ( .A(B[113]), .Z(n373) );
  IV U209 ( .A(B[114]), .Z(n374) );
  IV U210 ( .A(B[115]), .Z(n375) );
  IV U211 ( .A(B[116]), .Z(n376) );
  IV U212 ( .A(B[117]), .Z(n377) );
  IV U213 ( .A(B[118]), .Z(n378) );
  IV U214 ( .A(B[244]), .Z(n504) );
  IV U215 ( .A(B[119]), .Z(n379) );
  IV U216 ( .A(B[120]), .Z(n380) );
  IV U217 ( .A(B[121]), .Z(n381) );
  IV U218 ( .A(B[122]), .Z(n382) );
  IV U219 ( .A(B[123]), .Z(n383) );
  IV U220 ( .A(B[124]), .Z(n384) );
  IV U221 ( .A(B[125]), .Z(n385) );
  IV U222 ( .A(B[126]), .Z(n386) );
  IV U223 ( .A(B[127]), .Z(n387) );
  IV U224 ( .A(B[128]), .Z(n388) );
  IV U225 ( .A(B[245]), .Z(n505) );
  IV U226 ( .A(B[129]), .Z(n389) );
  IV U227 ( .A(B[130]), .Z(n390) );
  IV U228 ( .A(B[131]), .Z(n391) );
  IV U229 ( .A(B[132]), .Z(n392) );
  IV U230 ( .A(B[133]), .Z(n393) );
  IV U231 ( .A(B[134]), .Z(n394) );
  IV U232 ( .A(B[135]), .Z(n395) );
  IV U233 ( .A(B[136]), .Z(n396) );
  IV U234 ( .A(B[137]), .Z(n397) );
  IV U235 ( .A(B[138]), .Z(n398) );
  IV U236 ( .A(B[246]), .Z(n506) );
  IV U237 ( .A(B[139]), .Z(n399) );
  IV U238 ( .A(B[140]), .Z(n400) );
  IV U239 ( .A(B[141]), .Z(n401) );
  IV U240 ( .A(B[142]), .Z(n402) );
  IV U241 ( .A(B[143]), .Z(n403) );
  IV U242 ( .A(B[144]), .Z(n404) );
  IV U243 ( .A(B[145]), .Z(n405) );
  IV U244 ( .A(B[146]), .Z(n406) );
  IV U245 ( .A(B[147]), .Z(n407) );
  IV U246 ( .A(B[148]), .Z(n408) );
  IV U247 ( .A(B[247]), .Z(n507) );
  IV U248 ( .A(B[149]), .Z(n409) );
  IV U249 ( .A(B[150]), .Z(n410) );
  IV U250 ( .A(B[151]), .Z(n411) );
  IV U251 ( .A(B[152]), .Z(n412) );
  IV U252 ( .A(B[153]), .Z(n413) );
  IV U253 ( .A(B[154]), .Z(n414) );
  IV U254 ( .A(B[155]), .Z(n415) );
  IV U255 ( .A(B[156]), .Z(n416) );
  IV U256 ( .A(B[157]), .Z(n417) );
  IV U257 ( .A(B[158]), .Z(n418) );
  IV U258 ( .A(B[248]), .Z(n508) );
  IV U259 ( .A(B[257]), .Z(n517) );
endmodule


module FA_2064 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  OR U1 ( .A(CI), .B(A), .Z(CO) );
endmodule


module FA_2065 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  OR U1 ( .A(CI), .B(A), .Z(CO) );
endmodule


module FA_2066 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2067 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2068 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2069 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2070 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2071 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2072 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2073 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2074 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2075 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2076 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2077 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2078 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2079 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2080 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2081 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2082 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2083 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2084 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2085 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2086 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2087 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2088 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2089 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2090 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2091 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2092 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2093 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2094 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2095 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2096 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2097 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2098 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2099 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2100 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2101 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2102 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2103 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2104 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2105 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2106 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2107 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2108 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2109 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2110 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2111 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2112 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2113 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2114 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2115 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2116 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2117 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2118 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2119 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2120 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2121 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2122 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2123 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2124 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2125 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2126 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2127 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2128 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2129 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2130 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2131 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2132 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2133 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2134 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2135 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2136 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2137 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2138 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2139 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2140 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2141 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2142 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2143 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2144 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2145 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2146 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2147 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2148 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2149 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2150 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2151 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2152 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2153 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2154 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2155 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2156 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2157 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2158 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2159 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2160 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2161 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2162 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2163 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2164 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2165 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2166 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2167 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2168 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2169 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2170 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2171 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2172 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2173 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2174 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2175 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2176 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2177 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2178 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2179 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2180 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2181 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2182 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2183 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2184 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2185 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2186 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2187 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2188 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2189 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2190 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2191 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2192 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2193 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2194 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2195 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2196 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2197 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2198 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2199 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2200 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2201 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2202 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2203 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2204 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2205 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2206 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2207 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2208 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2209 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2210 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2211 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2212 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2213 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2214 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2215 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2216 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2217 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2218 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2219 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2220 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2221 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2222 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2223 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2224 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2225 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2226 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2227 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2228 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2229 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2230 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2231 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2232 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2233 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2234 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2235 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2236 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2237 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2238 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2239 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2240 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2241 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2242 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2243 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2244 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2245 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2246 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2247 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2248 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2249 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2250 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2251 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2252 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2253 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2254 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2255 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2256 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2257 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2258 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2259 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2260 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2261 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2262 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2263 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2264 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2265 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2266 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2267 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2268 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2269 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2270 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2271 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2272 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2273 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2274 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2275 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2276 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2277 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2278 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2279 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2280 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2281 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2282 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2283 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2284 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2285 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2286 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2287 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2288 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2289 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2290 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2291 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2292 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2293 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2294 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2295 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2296 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2297 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2298 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2299 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2300 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2301 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2302 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2303 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2304 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2305 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2306 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2307 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2308 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2309 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2310 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2311 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2312 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2313 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2314 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2315 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2316 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2317 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2318 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2319 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2320 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_2321 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  OR U1 ( .A(B), .B(A), .Z(CO) );
endmodule


module COMP_N258_4 ( A, B, O );
  input [257:0] A;
  input [257:0] B;
  output O;
  wire   n2, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512;
  wire   [257:1] C;

  FA_2321 \FAINST[0].FA_  ( .A(A[0]), .B(n2), .CI(1'b1), .CO(C[1]) );
  FA_2320 \FAINST[1].FA_  ( .A(A[1]), .B(n258), .CI(C[1]), .CO(C[2]) );
  FA_2319 \FAINST[2].FA_  ( .A(A[2]), .B(n259), .CI(C[2]), .CO(C[3]) );
  FA_2318 \FAINST[3].FA_  ( .A(A[3]), .B(n260), .CI(C[3]), .CO(C[4]) );
  FA_2317 \FAINST[4].FA_  ( .A(A[4]), .B(n261), .CI(C[4]), .CO(C[5]) );
  FA_2316 \FAINST[5].FA_  ( .A(A[5]), .B(n262), .CI(C[5]), .CO(C[6]) );
  FA_2315 \FAINST[6].FA_  ( .A(A[6]), .B(n263), .CI(C[6]), .CO(C[7]) );
  FA_2314 \FAINST[7].FA_  ( .A(A[7]), .B(n264), .CI(C[7]), .CO(C[8]) );
  FA_2313 \FAINST[8].FA_  ( .A(A[8]), .B(n265), .CI(C[8]), .CO(C[9]) );
  FA_2312 \FAINST[9].FA_  ( .A(A[9]), .B(n266), .CI(C[9]), .CO(C[10]) );
  FA_2311 \FAINST[10].FA_  ( .A(A[10]), .B(n267), .CI(C[10]), .CO(C[11]) );
  FA_2310 \FAINST[11].FA_  ( .A(A[11]), .B(n268), .CI(C[11]), .CO(C[12]) );
  FA_2309 \FAINST[12].FA_  ( .A(A[12]), .B(n269), .CI(C[12]), .CO(C[13]) );
  FA_2308 \FAINST[13].FA_  ( .A(A[13]), .B(n270), .CI(C[13]), .CO(C[14]) );
  FA_2307 \FAINST[14].FA_  ( .A(A[14]), .B(n271), .CI(C[14]), .CO(C[15]) );
  FA_2306 \FAINST[15].FA_  ( .A(A[15]), .B(n272), .CI(C[15]), .CO(C[16]) );
  FA_2305 \FAINST[16].FA_  ( .A(A[16]), .B(n273), .CI(C[16]), .CO(C[17]) );
  FA_2304 \FAINST[17].FA_  ( .A(A[17]), .B(n274), .CI(C[17]), .CO(C[18]) );
  FA_2303 \FAINST[18].FA_  ( .A(A[18]), .B(n275), .CI(C[18]), .CO(C[19]) );
  FA_2302 \FAINST[19].FA_  ( .A(A[19]), .B(n276), .CI(C[19]), .CO(C[20]) );
  FA_2301 \FAINST[20].FA_  ( .A(A[20]), .B(n277), .CI(C[20]), .CO(C[21]) );
  FA_2300 \FAINST[21].FA_  ( .A(A[21]), .B(n278), .CI(C[21]), .CO(C[22]) );
  FA_2299 \FAINST[22].FA_  ( .A(A[22]), .B(n279), .CI(C[22]), .CO(C[23]) );
  FA_2298 \FAINST[23].FA_  ( .A(A[23]), .B(n280), .CI(C[23]), .CO(C[24]) );
  FA_2297 \FAINST[24].FA_  ( .A(A[24]), .B(n281), .CI(C[24]), .CO(C[25]) );
  FA_2296 \FAINST[25].FA_  ( .A(A[25]), .B(n282), .CI(C[25]), .CO(C[26]) );
  FA_2295 \FAINST[26].FA_  ( .A(A[26]), .B(n283), .CI(C[26]), .CO(C[27]) );
  FA_2294 \FAINST[27].FA_  ( .A(A[27]), .B(n284), .CI(C[27]), .CO(C[28]) );
  FA_2293 \FAINST[28].FA_  ( .A(A[28]), .B(n285), .CI(C[28]), .CO(C[29]) );
  FA_2292 \FAINST[29].FA_  ( .A(A[29]), .B(n286), .CI(C[29]), .CO(C[30]) );
  FA_2291 \FAINST[30].FA_  ( .A(A[30]), .B(n287), .CI(C[30]), .CO(C[31]) );
  FA_2290 \FAINST[31].FA_  ( .A(A[31]), .B(n288), .CI(C[31]), .CO(C[32]) );
  FA_2289 \FAINST[32].FA_  ( .A(A[32]), .B(n289), .CI(C[32]), .CO(C[33]) );
  FA_2288 \FAINST[33].FA_  ( .A(A[33]), .B(n290), .CI(C[33]), .CO(C[34]) );
  FA_2287 \FAINST[34].FA_  ( .A(A[34]), .B(n291), .CI(C[34]), .CO(C[35]) );
  FA_2286 \FAINST[35].FA_  ( .A(A[35]), .B(n292), .CI(C[35]), .CO(C[36]) );
  FA_2285 \FAINST[36].FA_  ( .A(A[36]), .B(n293), .CI(C[36]), .CO(C[37]) );
  FA_2284 \FAINST[37].FA_  ( .A(A[37]), .B(n294), .CI(C[37]), .CO(C[38]) );
  FA_2283 \FAINST[38].FA_  ( .A(A[38]), .B(n295), .CI(C[38]), .CO(C[39]) );
  FA_2282 \FAINST[39].FA_  ( .A(A[39]), .B(n296), .CI(C[39]), .CO(C[40]) );
  FA_2281 \FAINST[40].FA_  ( .A(A[40]), .B(n297), .CI(C[40]), .CO(C[41]) );
  FA_2280 \FAINST[41].FA_  ( .A(A[41]), .B(n298), .CI(C[41]), .CO(C[42]) );
  FA_2279 \FAINST[42].FA_  ( .A(A[42]), .B(n299), .CI(C[42]), .CO(C[43]) );
  FA_2278 \FAINST[43].FA_  ( .A(A[43]), .B(n300), .CI(C[43]), .CO(C[44]) );
  FA_2277 \FAINST[44].FA_  ( .A(A[44]), .B(n301), .CI(C[44]), .CO(C[45]) );
  FA_2276 \FAINST[45].FA_  ( .A(A[45]), .B(n302), .CI(C[45]), .CO(C[46]) );
  FA_2275 \FAINST[46].FA_  ( .A(A[46]), .B(n303), .CI(C[46]), .CO(C[47]) );
  FA_2274 \FAINST[47].FA_  ( .A(A[47]), .B(n304), .CI(C[47]), .CO(C[48]) );
  FA_2273 \FAINST[48].FA_  ( .A(A[48]), .B(n305), .CI(C[48]), .CO(C[49]) );
  FA_2272 \FAINST[49].FA_  ( .A(A[49]), .B(n306), .CI(C[49]), .CO(C[50]) );
  FA_2271 \FAINST[50].FA_  ( .A(A[50]), .B(n307), .CI(C[50]), .CO(C[51]) );
  FA_2270 \FAINST[51].FA_  ( .A(A[51]), .B(n308), .CI(C[51]), .CO(C[52]) );
  FA_2269 \FAINST[52].FA_  ( .A(A[52]), .B(n309), .CI(C[52]), .CO(C[53]) );
  FA_2268 \FAINST[53].FA_  ( .A(A[53]), .B(n310), .CI(C[53]), .CO(C[54]) );
  FA_2267 \FAINST[54].FA_  ( .A(A[54]), .B(n311), .CI(C[54]), .CO(C[55]) );
  FA_2266 \FAINST[55].FA_  ( .A(A[55]), .B(n312), .CI(C[55]), .CO(C[56]) );
  FA_2265 \FAINST[56].FA_  ( .A(A[56]), .B(n313), .CI(C[56]), .CO(C[57]) );
  FA_2264 \FAINST[57].FA_  ( .A(A[57]), .B(n314), .CI(C[57]), .CO(C[58]) );
  FA_2263 \FAINST[58].FA_  ( .A(A[58]), .B(n315), .CI(C[58]), .CO(C[59]) );
  FA_2262 \FAINST[59].FA_  ( .A(A[59]), .B(n316), .CI(C[59]), .CO(C[60]) );
  FA_2261 \FAINST[60].FA_  ( .A(A[60]), .B(n317), .CI(C[60]), .CO(C[61]) );
  FA_2260 \FAINST[61].FA_  ( .A(A[61]), .B(n318), .CI(C[61]), .CO(C[62]) );
  FA_2259 \FAINST[62].FA_  ( .A(A[62]), .B(n319), .CI(C[62]), .CO(C[63]) );
  FA_2258 \FAINST[63].FA_  ( .A(A[63]), .B(n320), .CI(C[63]), .CO(C[64]) );
  FA_2257 \FAINST[64].FA_  ( .A(A[64]), .B(n321), .CI(C[64]), .CO(C[65]) );
  FA_2256 \FAINST[65].FA_  ( .A(A[65]), .B(n322), .CI(C[65]), .CO(C[66]) );
  FA_2255 \FAINST[66].FA_  ( .A(A[66]), .B(n323), .CI(C[66]), .CO(C[67]) );
  FA_2254 \FAINST[67].FA_  ( .A(A[67]), .B(n324), .CI(C[67]), .CO(C[68]) );
  FA_2253 \FAINST[68].FA_  ( .A(A[68]), .B(n325), .CI(C[68]), .CO(C[69]) );
  FA_2252 \FAINST[69].FA_  ( .A(A[69]), .B(n326), .CI(C[69]), .CO(C[70]) );
  FA_2251 \FAINST[70].FA_  ( .A(A[70]), .B(n327), .CI(C[70]), .CO(C[71]) );
  FA_2250 \FAINST[71].FA_  ( .A(A[71]), .B(n328), .CI(C[71]), .CO(C[72]) );
  FA_2249 \FAINST[72].FA_  ( .A(A[72]), .B(n329), .CI(C[72]), .CO(C[73]) );
  FA_2248 \FAINST[73].FA_  ( .A(A[73]), .B(n330), .CI(C[73]), .CO(C[74]) );
  FA_2247 \FAINST[74].FA_  ( .A(A[74]), .B(n331), .CI(C[74]), .CO(C[75]) );
  FA_2246 \FAINST[75].FA_  ( .A(A[75]), .B(n332), .CI(C[75]), .CO(C[76]) );
  FA_2245 \FAINST[76].FA_  ( .A(A[76]), .B(n333), .CI(C[76]), .CO(C[77]) );
  FA_2244 \FAINST[77].FA_  ( .A(A[77]), .B(n334), .CI(C[77]), .CO(C[78]) );
  FA_2243 \FAINST[78].FA_  ( .A(A[78]), .B(n335), .CI(C[78]), .CO(C[79]) );
  FA_2242 \FAINST[79].FA_  ( .A(A[79]), .B(n336), .CI(C[79]), .CO(C[80]) );
  FA_2241 \FAINST[80].FA_  ( .A(A[80]), .B(n337), .CI(C[80]), .CO(C[81]) );
  FA_2240 \FAINST[81].FA_  ( .A(A[81]), .B(n338), .CI(C[81]), .CO(C[82]) );
  FA_2239 \FAINST[82].FA_  ( .A(A[82]), .B(n339), .CI(C[82]), .CO(C[83]) );
  FA_2238 \FAINST[83].FA_  ( .A(A[83]), .B(n340), .CI(C[83]), .CO(C[84]) );
  FA_2237 \FAINST[84].FA_  ( .A(A[84]), .B(n341), .CI(C[84]), .CO(C[85]) );
  FA_2236 \FAINST[85].FA_  ( .A(A[85]), .B(n342), .CI(C[85]), .CO(C[86]) );
  FA_2235 \FAINST[86].FA_  ( .A(A[86]), .B(n343), .CI(C[86]), .CO(C[87]) );
  FA_2234 \FAINST[87].FA_  ( .A(A[87]), .B(n344), .CI(C[87]), .CO(C[88]) );
  FA_2233 \FAINST[88].FA_  ( .A(A[88]), .B(n345), .CI(C[88]), .CO(C[89]) );
  FA_2232 \FAINST[89].FA_  ( .A(A[89]), .B(n346), .CI(C[89]), .CO(C[90]) );
  FA_2231 \FAINST[90].FA_  ( .A(A[90]), .B(n347), .CI(C[90]), .CO(C[91]) );
  FA_2230 \FAINST[91].FA_  ( .A(A[91]), .B(n348), .CI(C[91]), .CO(C[92]) );
  FA_2229 \FAINST[92].FA_  ( .A(A[92]), .B(n349), .CI(C[92]), .CO(C[93]) );
  FA_2228 \FAINST[93].FA_  ( .A(A[93]), .B(n350), .CI(C[93]), .CO(C[94]) );
  FA_2227 \FAINST[94].FA_  ( .A(A[94]), .B(n351), .CI(C[94]), .CO(C[95]) );
  FA_2226 \FAINST[95].FA_  ( .A(A[95]), .B(n352), .CI(C[95]), .CO(C[96]) );
  FA_2225 \FAINST[96].FA_  ( .A(A[96]), .B(n353), .CI(C[96]), .CO(C[97]) );
  FA_2224 \FAINST[97].FA_  ( .A(A[97]), .B(n354), .CI(C[97]), .CO(C[98]) );
  FA_2223 \FAINST[98].FA_  ( .A(A[98]), .B(n355), .CI(C[98]), .CO(C[99]) );
  FA_2222 \FAINST[99].FA_  ( .A(A[99]), .B(n356), .CI(C[99]), .CO(C[100]) );
  FA_2221 \FAINST[100].FA_  ( .A(A[100]), .B(n357), .CI(C[100]), .CO(C[101])
         );
  FA_2220 \FAINST[101].FA_  ( .A(A[101]), .B(n358), .CI(C[101]), .CO(C[102])
         );
  FA_2219 \FAINST[102].FA_  ( .A(A[102]), .B(n359), .CI(C[102]), .CO(C[103])
         );
  FA_2218 \FAINST[103].FA_  ( .A(A[103]), .B(n360), .CI(C[103]), .CO(C[104])
         );
  FA_2217 \FAINST[104].FA_  ( .A(A[104]), .B(n361), .CI(C[104]), .CO(C[105])
         );
  FA_2216 \FAINST[105].FA_  ( .A(A[105]), .B(n362), .CI(C[105]), .CO(C[106])
         );
  FA_2215 \FAINST[106].FA_  ( .A(A[106]), .B(n363), .CI(C[106]), .CO(C[107])
         );
  FA_2214 \FAINST[107].FA_  ( .A(A[107]), .B(n364), .CI(C[107]), .CO(C[108])
         );
  FA_2213 \FAINST[108].FA_  ( .A(A[108]), .B(n365), .CI(C[108]), .CO(C[109])
         );
  FA_2212 \FAINST[109].FA_  ( .A(A[109]), .B(n366), .CI(C[109]), .CO(C[110])
         );
  FA_2211 \FAINST[110].FA_  ( .A(A[110]), .B(n367), .CI(C[110]), .CO(C[111])
         );
  FA_2210 \FAINST[111].FA_  ( .A(A[111]), .B(n368), .CI(C[111]), .CO(C[112])
         );
  FA_2209 \FAINST[112].FA_  ( .A(A[112]), .B(n369), .CI(C[112]), .CO(C[113])
         );
  FA_2208 \FAINST[113].FA_  ( .A(A[113]), .B(n370), .CI(C[113]), .CO(C[114])
         );
  FA_2207 \FAINST[114].FA_  ( .A(A[114]), .B(n371), .CI(C[114]), .CO(C[115])
         );
  FA_2206 \FAINST[115].FA_  ( .A(A[115]), .B(n372), .CI(C[115]), .CO(C[116])
         );
  FA_2205 \FAINST[116].FA_  ( .A(A[116]), .B(n373), .CI(C[116]), .CO(C[117])
         );
  FA_2204 \FAINST[117].FA_  ( .A(A[117]), .B(n374), .CI(C[117]), .CO(C[118])
         );
  FA_2203 \FAINST[118].FA_  ( .A(A[118]), .B(n375), .CI(C[118]), .CO(C[119])
         );
  FA_2202 \FAINST[119].FA_  ( .A(A[119]), .B(n376), .CI(C[119]), .CO(C[120])
         );
  FA_2201 \FAINST[120].FA_  ( .A(A[120]), .B(n377), .CI(C[120]), .CO(C[121])
         );
  FA_2200 \FAINST[121].FA_  ( .A(A[121]), .B(n378), .CI(C[121]), .CO(C[122])
         );
  FA_2199 \FAINST[122].FA_  ( .A(A[122]), .B(n379), .CI(C[122]), .CO(C[123])
         );
  FA_2198 \FAINST[123].FA_  ( .A(A[123]), .B(n380), .CI(C[123]), .CO(C[124])
         );
  FA_2197 \FAINST[124].FA_  ( .A(A[124]), .B(n381), .CI(C[124]), .CO(C[125])
         );
  FA_2196 \FAINST[125].FA_  ( .A(A[125]), .B(n382), .CI(C[125]), .CO(C[126])
         );
  FA_2195 \FAINST[126].FA_  ( .A(A[126]), .B(n383), .CI(C[126]), .CO(C[127])
         );
  FA_2194 \FAINST[127].FA_  ( .A(A[127]), .B(n384), .CI(C[127]), .CO(C[128])
         );
  FA_2193 \FAINST[128].FA_  ( .A(A[128]), .B(n385), .CI(C[128]), .CO(C[129])
         );
  FA_2192 \FAINST[129].FA_  ( .A(A[129]), .B(n386), .CI(C[129]), .CO(C[130])
         );
  FA_2191 \FAINST[130].FA_  ( .A(A[130]), .B(n387), .CI(C[130]), .CO(C[131])
         );
  FA_2190 \FAINST[131].FA_  ( .A(A[131]), .B(n388), .CI(C[131]), .CO(C[132])
         );
  FA_2189 \FAINST[132].FA_  ( .A(A[132]), .B(n389), .CI(C[132]), .CO(C[133])
         );
  FA_2188 \FAINST[133].FA_  ( .A(A[133]), .B(n390), .CI(C[133]), .CO(C[134])
         );
  FA_2187 \FAINST[134].FA_  ( .A(A[134]), .B(n391), .CI(C[134]), .CO(C[135])
         );
  FA_2186 \FAINST[135].FA_  ( .A(A[135]), .B(n392), .CI(C[135]), .CO(C[136])
         );
  FA_2185 \FAINST[136].FA_  ( .A(A[136]), .B(n393), .CI(C[136]), .CO(C[137])
         );
  FA_2184 \FAINST[137].FA_  ( .A(A[137]), .B(n394), .CI(C[137]), .CO(C[138])
         );
  FA_2183 \FAINST[138].FA_  ( .A(A[138]), .B(n395), .CI(C[138]), .CO(C[139])
         );
  FA_2182 \FAINST[139].FA_  ( .A(A[139]), .B(n396), .CI(C[139]), .CO(C[140])
         );
  FA_2181 \FAINST[140].FA_  ( .A(A[140]), .B(n397), .CI(C[140]), .CO(C[141])
         );
  FA_2180 \FAINST[141].FA_  ( .A(A[141]), .B(n398), .CI(C[141]), .CO(C[142])
         );
  FA_2179 \FAINST[142].FA_  ( .A(A[142]), .B(n399), .CI(C[142]), .CO(C[143])
         );
  FA_2178 \FAINST[143].FA_  ( .A(A[143]), .B(n400), .CI(C[143]), .CO(C[144])
         );
  FA_2177 \FAINST[144].FA_  ( .A(A[144]), .B(n401), .CI(C[144]), .CO(C[145])
         );
  FA_2176 \FAINST[145].FA_  ( .A(A[145]), .B(n402), .CI(C[145]), .CO(C[146])
         );
  FA_2175 \FAINST[146].FA_  ( .A(A[146]), .B(n403), .CI(C[146]), .CO(C[147])
         );
  FA_2174 \FAINST[147].FA_  ( .A(A[147]), .B(n404), .CI(C[147]), .CO(C[148])
         );
  FA_2173 \FAINST[148].FA_  ( .A(A[148]), .B(n405), .CI(C[148]), .CO(C[149])
         );
  FA_2172 \FAINST[149].FA_  ( .A(A[149]), .B(n406), .CI(C[149]), .CO(C[150])
         );
  FA_2171 \FAINST[150].FA_  ( .A(A[150]), .B(n407), .CI(C[150]), .CO(C[151])
         );
  FA_2170 \FAINST[151].FA_  ( .A(A[151]), .B(n408), .CI(C[151]), .CO(C[152])
         );
  FA_2169 \FAINST[152].FA_  ( .A(A[152]), .B(n409), .CI(C[152]), .CO(C[153])
         );
  FA_2168 \FAINST[153].FA_  ( .A(A[153]), .B(n410), .CI(C[153]), .CO(C[154])
         );
  FA_2167 \FAINST[154].FA_  ( .A(A[154]), .B(n411), .CI(C[154]), .CO(C[155])
         );
  FA_2166 \FAINST[155].FA_  ( .A(A[155]), .B(n412), .CI(C[155]), .CO(C[156])
         );
  FA_2165 \FAINST[156].FA_  ( .A(A[156]), .B(n413), .CI(C[156]), .CO(C[157])
         );
  FA_2164 \FAINST[157].FA_  ( .A(A[157]), .B(n414), .CI(C[157]), .CO(C[158])
         );
  FA_2163 \FAINST[158].FA_  ( .A(A[158]), .B(n415), .CI(C[158]), .CO(C[159])
         );
  FA_2162 \FAINST[159].FA_  ( .A(A[159]), .B(n416), .CI(C[159]), .CO(C[160])
         );
  FA_2161 \FAINST[160].FA_  ( .A(A[160]), .B(n417), .CI(C[160]), .CO(C[161])
         );
  FA_2160 \FAINST[161].FA_  ( .A(A[161]), .B(n418), .CI(C[161]), .CO(C[162])
         );
  FA_2159 \FAINST[162].FA_  ( .A(A[162]), .B(n419), .CI(C[162]), .CO(C[163])
         );
  FA_2158 \FAINST[163].FA_  ( .A(A[163]), .B(n420), .CI(C[163]), .CO(C[164])
         );
  FA_2157 \FAINST[164].FA_  ( .A(A[164]), .B(n421), .CI(C[164]), .CO(C[165])
         );
  FA_2156 \FAINST[165].FA_  ( .A(A[165]), .B(n422), .CI(C[165]), .CO(C[166])
         );
  FA_2155 \FAINST[166].FA_  ( .A(A[166]), .B(n423), .CI(C[166]), .CO(C[167])
         );
  FA_2154 \FAINST[167].FA_  ( .A(A[167]), .B(n424), .CI(C[167]), .CO(C[168])
         );
  FA_2153 \FAINST[168].FA_  ( .A(A[168]), .B(n425), .CI(C[168]), .CO(C[169])
         );
  FA_2152 \FAINST[169].FA_  ( .A(A[169]), .B(n426), .CI(C[169]), .CO(C[170])
         );
  FA_2151 \FAINST[170].FA_  ( .A(A[170]), .B(n427), .CI(C[170]), .CO(C[171])
         );
  FA_2150 \FAINST[171].FA_  ( .A(A[171]), .B(n428), .CI(C[171]), .CO(C[172])
         );
  FA_2149 \FAINST[172].FA_  ( .A(A[172]), .B(n429), .CI(C[172]), .CO(C[173])
         );
  FA_2148 \FAINST[173].FA_  ( .A(A[173]), .B(n430), .CI(C[173]), .CO(C[174])
         );
  FA_2147 \FAINST[174].FA_  ( .A(A[174]), .B(n431), .CI(C[174]), .CO(C[175])
         );
  FA_2146 \FAINST[175].FA_  ( .A(A[175]), .B(n432), .CI(C[175]), .CO(C[176])
         );
  FA_2145 \FAINST[176].FA_  ( .A(A[176]), .B(n433), .CI(C[176]), .CO(C[177])
         );
  FA_2144 \FAINST[177].FA_  ( .A(A[177]), .B(n434), .CI(C[177]), .CO(C[178])
         );
  FA_2143 \FAINST[178].FA_  ( .A(A[178]), .B(n435), .CI(C[178]), .CO(C[179])
         );
  FA_2142 \FAINST[179].FA_  ( .A(A[179]), .B(n436), .CI(C[179]), .CO(C[180])
         );
  FA_2141 \FAINST[180].FA_  ( .A(A[180]), .B(n437), .CI(C[180]), .CO(C[181])
         );
  FA_2140 \FAINST[181].FA_  ( .A(A[181]), .B(n438), .CI(C[181]), .CO(C[182])
         );
  FA_2139 \FAINST[182].FA_  ( .A(A[182]), .B(n439), .CI(C[182]), .CO(C[183])
         );
  FA_2138 \FAINST[183].FA_  ( .A(A[183]), .B(n440), .CI(C[183]), .CO(C[184])
         );
  FA_2137 \FAINST[184].FA_  ( .A(A[184]), .B(n441), .CI(C[184]), .CO(C[185])
         );
  FA_2136 \FAINST[185].FA_  ( .A(A[185]), .B(n442), .CI(C[185]), .CO(C[186])
         );
  FA_2135 \FAINST[186].FA_  ( .A(A[186]), .B(n443), .CI(C[186]), .CO(C[187])
         );
  FA_2134 \FAINST[187].FA_  ( .A(A[187]), .B(n444), .CI(C[187]), .CO(C[188])
         );
  FA_2133 \FAINST[188].FA_  ( .A(A[188]), .B(n445), .CI(C[188]), .CO(C[189])
         );
  FA_2132 \FAINST[189].FA_  ( .A(A[189]), .B(n446), .CI(C[189]), .CO(C[190])
         );
  FA_2131 \FAINST[190].FA_  ( .A(A[190]), .B(n447), .CI(C[190]), .CO(C[191])
         );
  FA_2130 \FAINST[191].FA_  ( .A(A[191]), .B(n448), .CI(C[191]), .CO(C[192])
         );
  FA_2129 \FAINST[192].FA_  ( .A(A[192]), .B(n449), .CI(C[192]), .CO(C[193])
         );
  FA_2128 \FAINST[193].FA_  ( .A(A[193]), .B(n450), .CI(C[193]), .CO(C[194])
         );
  FA_2127 \FAINST[194].FA_  ( .A(A[194]), .B(n451), .CI(C[194]), .CO(C[195])
         );
  FA_2126 \FAINST[195].FA_  ( .A(A[195]), .B(n452), .CI(C[195]), .CO(C[196])
         );
  FA_2125 \FAINST[196].FA_  ( .A(A[196]), .B(n453), .CI(C[196]), .CO(C[197])
         );
  FA_2124 \FAINST[197].FA_  ( .A(A[197]), .B(n454), .CI(C[197]), .CO(C[198])
         );
  FA_2123 \FAINST[198].FA_  ( .A(A[198]), .B(n455), .CI(C[198]), .CO(C[199])
         );
  FA_2122 \FAINST[199].FA_  ( .A(A[199]), .B(n456), .CI(C[199]), .CO(C[200])
         );
  FA_2121 \FAINST[200].FA_  ( .A(A[200]), .B(n457), .CI(C[200]), .CO(C[201])
         );
  FA_2120 \FAINST[201].FA_  ( .A(A[201]), .B(n458), .CI(C[201]), .CO(C[202])
         );
  FA_2119 \FAINST[202].FA_  ( .A(A[202]), .B(n459), .CI(C[202]), .CO(C[203])
         );
  FA_2118 \FAINST[203].FA_  ( .A(A[203]), .B(n460), .CI(C[203]), .CO(C[204])
         );
  FA_2117 \FAINST[204].FA_  ( .A(A[204]), .B(n461), .CI(C[204]), .CO(C[205])
         );
  FA_2116 \FAINST[205].FA_  ( .A(A[205]), .B(n462), .CI(C[205]), .CO(C[206])
         );
  FA_2115 \FAINST[206].FA_  ( .A(A[206]), .B(n463), .CI(C[206]), .CO(C[207])
         );
  FA_2114 \FAINST[207].FA_  ( .A(A[207]), .B(n464), .CI(C[207]), .CO(C[208])
         );
  FA_2113 \FAINST[208].FA_  ( .A(A[208]), .B(n465), .CI(C[208]), .CO(C[209])
         );
  FA_2112 \FAINST[209].FA_  ( .A(A[209]), .B(n466), .CI(C[209]), .CO(C[210])
         );
  FA_2111 \FAINST[210].FA_  ( .A(A[210]), .B(n467), .CI(C[210]), .CO(C[211])
         );
  FA_2110 \FAINST[211].FA_  ( .A(A[211]), .B(n468), .CI(C[211]), .CO(C[212])
         );
  FA_2109 \FAINST[212].FA_  ( .A(A[212]), .B(n469), .CI(C[212]), .CO(C[213])
         );
  FA_2108 \FAINST[213].FA_  ( .A(A[213]), .B(n470), .CI(C[213]), .CO(C[214])
         );
  FA_2107 \FAINST[214].FA_  ( .A(A[214]), .B(n471), .CI(C[214]), .CO(C[215])
         );
  FA_2106 \FAINST[215].FA_  ( .A(A[215]), .B(n472), .CI(C[215]), .CO(C[216])
         );
  FA_2105 \FAINST[216].FA_  ( .A(A[216]), .B(n473), .CI(C[216]), .CO(C[217])
         );
  FA_2104 \FAINST[217].FA_  ( .A(A[217]), .B(n474), .CI(C[217]), .CO(C[218])
         );
  FA_2103 \FAINST[218].FA_  ( .A(A[218]), .B(n475), .CI(C[218]), .CO(C[219])
         );
  FA_2102 \FAINST[219].FA_  ( .A(A[219]), .B(n476), .CI(C[219]), .CO(C[220])
         );
  FA_2101 \FAINST[220].FA_  ( .A(A[220]), .B(n477), .CI(C[220]), .CO(C[221])
         );
  FA_2100 \FAINST[221].FA_  ( .A(A[221]), .B(n478), .CI(C[221]), .CO(C[222])
         );
  FA_2099 \FAINST[222].FA_  ( .A(A[222]), .B(n479), .CI(C[222]), .CO(C[223])
         );
  FA_2098 \FAINST[223].FA_  ( .A(A[223]), .B(n480), .CI(C[223]), .CO(C[224])
         );
  FA_2097 \FAINST[224].FA_  ( .A(A[224]), .B(n481), .CI(C[224]), .CO(C[225])
         );
  FA_2096 \FAINST[225].FA_  ( .A(A[225]), .B(n482), .CI(C[225]), .CO(C[226])
         );
  FA_2095 \FAINST[226].FA_  ( .A(A[226]), .B(n483), .CI(C[226]), .CO(C[227])
         );
  FA_2094 \FAINST[227].FA_  ( .A(A[227]), .B(n484), .CI(C[227]), .CO(C[228])
         );
  FA_2093 \FAINST[228].FA_  ( .A(A[228]), .B(n485), .CI(C[228]), .CO(C[229])
         );
  FA_2092 \FAINST[229].FA_  ( .A(A[229]), .B(n486), .CI(C[229]), .CO(C[230])
         );
  FA_2091 \FAINST[230].FA_  ( .A(A[230]), .B(n487), .CI(C[230]), .CO(C[231])
         );
  FA_2090 \FAINST[231].FA_  ( .A(A[231]), .B(n488), .CI(C[231]), .CO(C[232])
         );
  FA_2089 \FAINST[232].FA_  ( .A(A[232]), .B(n489), .CI(C[232]), .CO(C[233])
         );
  FA_2088 \FAINST[233].FA_  ( .A(A[233]), .B(n490), .CI(C[233]), .CO(C[234])
         );
  FA_2087 \FAINST[234].FA_  ( .A(A[234]), .B(n491), .CI(C[234]), .CO(C[235])
         );
  FA_2086 \FAINST[235].FA_  ( .A(A[235]), .B(n492), .CI(C[235]), .CO(C[236])
         );
  FA_2085 \FAINST[236].FA_  ( .A(A[236]), .B(n493), .CI(C[236]), .CO(C[237])
         );
  FA_2084 \FAINST[237].FA_  ( .A(A[237]), .B(n494), .CI(C[237]), .CO(C[238])
         );
  FA_2083 \FAINST[238].FA_  ( .A(A[238]), .B(n495), .CI(C[238]), .CO(C[239])
         );
  FA_2082 \FAINST[239].FA_  ( .A(A[239]), .B(n496), .CI(C[239]), .CO(C[240])
         );
  FA_2081 \FAINST[240].FA_  ( .A(A[240]), .B(n497), .CI(C[240]), .CO(C[241])
         );
  FA_2080 \FAINST[241].FA_  ( .A(A[241]), .B(n498), .CI(C[241]), .CO(C[242])
         );
  FA_2079 \FAINST[242].FA_  ( .A(A[242]), .B(n499), .CI(C[242]), .CO(C[243])
         );
  FA_2078 \FAINST[243].FA_  ( .A(A[243]), .B(n500), .CI(C[243]), .CO(C[244])
         );
  FA_2077 \FAINST[244].FA_  ( .A(A[244]), .B(n501), .CI(C[244]), .CO(C[245])
         );
  FA_2076 \FAINST[245].FA_  ( .A(A[245]), .B(n502), .CI(C[245]), .CO(C[246])
         );
  FA_2075 \FAINST[246].FA_  ( .A(A[246]), .B(n503), .CI(C[246]), .CO(C[247])
         );
  FA_2074 \FAINST[247].FA_  ( .A(A[247]), .B(n504), .CI(C[247]), .CO(C[248])
         );
  FA_2073 \FAINST[248].FA_  ( .A(A[248]), .B(n505), .CI(C[248]), .CO(C[249])
         );
  FA_2072 \FAINST[249].FA_  ( .A(A[249]), .B(n506), .CI(C[249]), .CO(C[250])
         );
  FA_2071 \FAINST[250].FA_  ( .A(A[250]), .B(n507), .CI(C[250]), .CO(C[251])
         );
  FA_2070 \FAINST[251].FA_  ( .A(A[251]), .B(n508), .CI(C[251]), .CO(C[252])
         );
  FA_2069 \FAINST[252].FA_  ( .A(A[252]), .B(n509), .CI(C[252]), .CO(C[253])
         );
  FA_2068 \FAINST[253].FA_  ( .A(A[253]), .B(n510), .CI(C[253]), .CO(C[254])
         );
  FA_2067 \FAINST[254].FA_  ( .A(A[254]), .B(n511), .CI(C[254]), .CO(C[255])
         );
  FA_2066 \FAINST[255].FA_  ( .A(A[255]), .B(n512), .CI(C[255]), .CO(C[256])
         );
  FA_2065 \FAINST[256].FA_  ( .A(A[256]), .B(1'b1), .CI(C[256]), .CO(C[257])
         );
  FA_2064 \FAINST[257].FA_  ( .A(A[257]), .B(1'b1), .CI(C[257]), .CO(O) );
  IV U2 ( .A(B[159]), .Z(n416) );
  IV U3 ( .A(B[160]), .Z(n417) );
  IV U4 ( .A(B[161]), .Z(n418) );
  IV U5 ( .A(B[162]), .Z(n419) );
  IV U6 ( .A(B[163]), .Z(n420) );
  IV U7 ( .A(B[164]), .Z(n421) );
  IV U8 ( .A(B[165]), .Z(n422) );
  IV U9 ( .A(B[166]), .Z(n423) );
  IV U10 ( .A(B[167]), .Z(n424) );
  IV U11 ( .A(B[168]), .Z(n425) );
  IV U12 ( .A(B[249]), .Z(n506) );
  IV U13 ( .A(B[169]), .Z(n426) );
  IV U14 ( .A(B[170]), .Z(n427) );
  IV U15 ( .A(B[171]), .Z(n428) );
  IV U16 ( .A(B[172]), .Z(n429) );
  IV U17 ( .A(B[173]), .Z(n430) );
  IV U18 ( .A(B[174]), .Z(n431) );
  IV U19 ( .A(B[175]), .Z(n432) );
  IV U20 ( .A(B[176]), .Z(n433) );
  IV U21 ( .A(B[177]), .Z(n434) );
  IV U22 ( .A(B[178]), .Z(n435) );
  IV U23 ( .A(B[250]), .Z(n507) );
  IV U24 ( .A(B[179]), .Z(n436) );
  IV U25 ( .A(B[180]), .Z(n437) );
  IV U26 ( .A(B[181]), .Z(n438) );
  IV U27 ( .A(B[182]), .Z(n439) );
  IV U28 ( .A(B[183]), .Z(n440) );
  IV U29 ( .A(B[184]), .Z(n441) );
  IV U30 ( .A(B[185]), .Z(n442) );
  IV U31 ( .A(B[186]), .Z(n443) );
  IV U32 ( .A(B[187]), .Z(n444) );
  IV U33 ( .A(B[188]), .Z(n445) );
  IV U34 ( .A(B[251]), .Z(n508) );
  IV U35 ( .A(B[189]), .Z(n446) );
  IV U36 ( .A(B[190]), .Z(n447) );
  IV U37 ( .A(B[191]), .Z(n448) );
  IV U38 ( .A(B[192]), .Z(n449) );
  IV U39 ( .A(B[193]), .Z(n450) );
  IV U40 ( .A(B[194]), .Z(n451) );
  IV U41 ( .A(B[195]), .Z(n452) );
  IV U42 ( .A(B[196]), .Z(n453) );
  IV U43 ( .A(B[197]), .Z(n454) );
  IV U44 ( .A(B[198]), .Z(n455) );
  IV U45 ( .A(B[252]), .Z(n509) );
  IV U46 ( .A(B[199]), .Z(n456) );
  IV U47 ( .A(B[200]), .Z(n457) );
  IV U48 ( .A(B[201]), .Z(n458) );
  IV U49 ( .A(B[202]), .Z(n459) );
  IV U50 ( .A(B[203]), .Z(n460) );
  IV U51 ( .A(B[204]), .Z(n461) );
  IV U52 ( .A(B[205]), .Z(n462) );
  IV U53 ( .A(B[206]), .Z(n463) );
  IV U54 ( .A(B[207]), .Z(n464) );
  IV U55 ( .A(B[208]), .Z(n465) );
  IV U56 ( .A(B[253]), .Z(n510) );
  IV U57 ( .A(B[209]), .Z(n466) );
  IV U58 ( .A(B[210]), .Z(n467) );
  IV U59 ( .A(B[211]), .Z(n468) );
  IV U60 ( .A(B[212]), .Z(n469) );
  IV U61 ( .A(B[213]), .Z(n470) );
  IV U62 ( .A(B[214]), .Z(n471) );
  IV U63 ( .A(B[215]), .Z(n472) );
  IV U64 ( .A(B[216]), .Z(n473) );
  IV U65 ( .A(B[217]), .Z(n474) );
  IV U66 ( .A(B[218]), .Z(n475) );
  IV U67 ( .A(B[254]), .Z(n511) );
  IV U68 ( .A(B[219]), .Z(n476) );
  IV U69 ( .A(B[220]), .Z(n477) );
  IV U70 ( .A(B[221]), .Z(n478) );
  IV U71 ( .A(B[222]), .Z(n479) );
  IV U72 ( .A(B[223]), .Z(n480) );
  IV U73 ( .A(B[224]), .Z(n481) );
  IV U74 ( .A(B[225]), .Z(n482) );
  IV U75 ( .A(B[226]), .Z(n483) );
  IV U76 ( .A(B[227]), .Z(n484) );
  IV U77 ( .A(B[228]), .Z(n485) );
  IV U78 ( .A(B[255]), .Z(n512) );
  IV U79 ( .A(B[229]), .Z(n486) );
  IV U80 ( .A(B[230]), .Z(n487) );
  IV U81 ( .A(B[231]), .Z(n488) );
  IV U82 ( .A(B[232]), .Z(n489) );
  IV U83 ( .A(B[0]), .Z(n2) );
  IV U84 ( .A(B[1]), .Z(n258) );
  IV U85 ( .A(B[2]), .Z(n259) );
  IV U86 ( .A(B[3]), .Z(n260) );
  IV U87 ( .A(B[4]), .Z(n261) );
  IV U88 ( .A(B[5]), .Z(n262) );
  IV U89 ( .A(B[6]), .Z(n263) );
  IV U90 ( .A(B[7]), .Z(n264) );
  IV U91 ( .A(B[8]), .Z(n265) );
  IV U92 ( .A(B[233]), .Z(n490) );
  IV U93 ( .A(B[9]), .Z(n266) );
  IV U94 ( .A(B[10]), .Z(n267) );
  IV U95 ( .A(B[11]), .Z(n268) );
  IV U96 ( .A(B[12]), .Z(n269) );
  IV U97 ( .A(B[13]), .Z(n270) );
  IV U98 ( .A(B[14]), .Z(n271) );
  IV U99 ( .A(B[15]), .Z(n272) );
  IV U100 ( .A(B[16]), .Z(n273) );
  IV U101 ( .A(B[17]), .Z(n274) );
  IV U102 ( .A(B[18]), .Z(n275) );
  IV U103 ( .A(B[234]), .Z(n491) );
  IV U104 ( .A(B[19]), .Z(n276) );
  IV U105 ( .A(B[20]), .Z(n277) );
  IV U106 ( .A(B[21]), .Z(n278) );
  IV U107 ( .A(B[22]), .Z(n279) );
  IV U108 ( .A(B[23]), .Z(n280) );
  IV U109 ( .A(B[24]), .Z(n281) );
  IV U110 ( .A(B[25]), .Z(n282) );
  IV U111 ( .A(B[26]), .Z(n283) );
  IV U112 ( .A(B[27]), .Z(n284) );
  IV U113 ( .A(B[28]), .Z(n285) );
  IV U114 ( .A(B[235]), .Z(n492) );
  IV U115 ( .A(B[29]), .Z(n286) );
  IV U116 ( .A(B[30]), .Z(n287) );
  IV U117 ( .A(B[31]), .Z(n288) );
  IV U118 ( .A(B[32]), .Z(n289) );
  IV U119 ( .A(B[33]), .Z(n290) );
  IV U120 ( .A(B[34]), .Z(n291) );
  IV U121 ( .A(B[35]), .Z(n292) );
  IV U122 ( .A(B[36]), .Z(n293) );
  IV U123 ( .A(B[37]), .Z(n294) );
  IV U124 ( .A(B[38]), .Z(n295) );
  IV U125 ( .A(B[236]), .Z(n493) );
  IV U126 ( .A(B[39]), .Z(n296) );
  IV U127 ( .A(B[40]), .Z(n297) );
  IV U128 ( .A(B[41]), .Z(n298) );
  IV U129 ( .A(B[42]), .Z(n299) );
  IV U130 ( .A(B[43]), .Z(n300) );
  IV U131 ( .A(B[44]), .Z(n301) );
  IV U132 ( .A(B[45]), .Z(n302) );
  IV U133 ( .A(B[46]), .Z(n303) );
  IV U134 ( .A(B[47]), .Z(n304) );
  IV U135 ( .A(B[48]), .Z(n305) );
  IV U136 ( .A(B[237]), .Z(n494) );
  IV U137 ( .A(B[49]), .Z(n306) );
  IV U138 ( .A(B[50]), .Z(n307) );
  IV U139 ( .A(B[51]), .Z(n308) );
  IV U140 ( .A(B[52]), .Z(n309) );
  IV U141 ( .A(B[53]), .Z(n310) );
  IV U142 ( .A(B[54]), .Z(n311) );
  IV U143 ( .A(B[55]), .Z(n312) );
  IV U144 ( .A(B[56]), .Z(n313) );
  IV U145 ( .A(B[57]), .Z(n314) );
  IV U146 ( .A(B[58]), .Z(n315) );
  IV U147 ( .A(B[238]), .Z(n495) );
  IV U148 ( .A(B[59]), .Z(n316) );
  IV U149 ( .A(B[60]), .Z(n317) );
  IV U150 ( .A(B[61]), .Z(n318) );
  IV U151 ( .A(B[62]), .Z(n319) );
  IV U152 ( .A(B[63]), .Z(n320) );
  IV U153 ( .A(B[64]), .Z(n321) );
  IV U154 ( .A(B[65]), .Z(n322) );
  IV U155 ( .A(B[66]), .Z(n323) );
  IV U156 ( .A(B[67]), .Z(n324) );
  IV U157 ( .A(B[68]), .Z(n325) );
  IV U158 ( .A(B[239]), .Z(n496) );
  IV U159 ( .A(B[69]), .Z(n326) );
  IV U160 ( .A(B[70]), .Z(n327) );
  IV U161 ( .A(B[71]), .Z(n328) );
  IV U162 ( .A(B[72]), .Z(n329) );
  IV U163 ( .A(B[73]), .Z(n330) );
  IV U164 ( .A(B[74]), .Z(n331) );
  IV U165 ( .A(B[75]), .Z(n332) );
  IV U166 ( .A(B[76]), .Z(n333) );
  IV U167 ( .A(B[77]), .Z(n334) );
  IV U168 ( .A(B[78]), .Z(n335) );
  IV U169 ( .A(B[240]), .Z(n497) );
  IV U170 ( .A(B[79]), .Z(n336) );
  IV U171 ( .A(B[80]), .Z(n337) );
  IV U172 ( .A(B[81]), .Z(n338) );
  IV U173 ( .A(B[82]), .Z(n339) );
  IV U174 ( .A(B[83]), .Z(n340) );
  IV U175 ( .A(B[84]), .Z(n341) );
  IV U176 ( .A(B[85]), .Z(n342) );
  IV U177 ( .A(B[86]), .Z(n343) );
  IV U178 ( .A(B[87]), .Z(n344) );
  IV U179 ( .A(B[88]), .Z(n345) );
  IV U180 ( .A(B[241]), .Z(n498) );
  IV U181 ( .A(B[89]), .Z(n346) );
  IV U182 ( .A(B[90]), .Z(n347) );
  IV U183 ( .A(B[91]), .Z(n348) );
  IV U184 ( .A(B[92]), .Z(n349) );
  IV U185 ( .A(B[93]), .Z(n350) );
  IV U186 ( .A(B[94]), .Z(n351) );
  IV U187 ( .A(B[95]), .Z(n352) );
  IV U188 ( .A(B[96]), .Z(n353) );
  IV U189 ( .A(B[97]), .Z(n354) );
  IV U190 ( .A(B[98]), .Z(n355) );
  IV U191 ( .A(B[242]), .Z(n499) );
  IV U192 ( .A(B[99]), .Z(n356) );
  IV U193 ( .A(B[100]), .Z(n357) );
  IV U194 ( .A(B[101]), .Z(n358) );
  IV U195 ( .A(B[102]), .Z(n359) );
  IV U196 ( .A(B[103]), .Z(n360) );
  IV U197 ( .A(B[104]), .Z(n361) );
  IV U198 ( .A(B[105]), .Z(n362) );
  IV U199 ( .A(B[106]), .Z(n363) );
  IV U200 ( .A(B[107]), .Z(n364) );
  IV U201 ( .A(B[108]), .Z(n365) );
  IV U202 ( .A(B[243]), .Z(n500) );
  IV U203 ( .A(B[109]), .Z(n366) );
  IV U204 ( .A(B[110]), .Z(n367) );
  IV U205 ( .A(B[111]), .Z(n368) );
  IV U206 ( .A(B[112]), .Z(n369) );
  IV U207 ( .A(B[113]), .Z(n370) );
  IV U208 ( .A(B[114]), .Z(n371) );
  IV U209 ( .A(B[115]), .Z(n372) );
  IV U210 ( .A(B[116]), .Z(n373) );
  IV U211 ( .A(B[117]), .Z(n374) );
  IV U212 ( .A(B[118]), .Z(n375) );
  IV U213 ( .A(B[244]), .Z(n501) );
  IV U214 ( .A(B[119]), .Z(n376) );
  IV U215 ( .A(B[120]), .Z(n377) );
  IV U216 ( .A(B[121]), .Z(n378) );
  IV U217 ( .A(B[122]), .Z(n379) );
  IV U218 ( .A(B[123]), .Z(n380) );
  IV U219 ( .A(B[124]), .Z(n381) );
  IV U220 ( .A(B[125]), .Z(n382) );
  IV U221 ( .A(B[126]), .Z(n383) );
  IV U222 ( .A(B[127]), .Z(n384) );
  IV U223 ( .A(B[128]), .Z(n385) );
  IV U224 ( .A(B[245]), .Z(n502) );
  IV U225 ( .A(B[129]), .Z(n386) );
  IV U226 ( .A(B[130]), .Z(n387) );
  IV U227 ( .A(B[131]), .Z(n388) );
  IV U228 ( .A(B[132]), .Z(n389) );
  IV U229 ( .A(B[133]), .Z(n390) );
  IV U230 ( .A(B[134]), .Z(n391) );
  IV U231 ( .A(B[135]), .Z(n392) );
  IV U232 ( .A(B[136]), .Z(n393) );
  IV U233 ( .A(B[137]), .Z(n394) );
  IV U234 ( .A(B[138]), .Z(n395) );
  IV U235 ( .A(B[246]), .Z(n503) );
  IV U236 ( .A(B[139]), .Z(n396) );
  IV U237 ( .A(B[140]), .Z(n397) );
  IV U238 ( .A(B[141]), .Z(n398) );
  IV U239 ( .A(B[142]), .Z(n399) );
  IV U240 ( .A(B[143]), .Z(n400) );
  IV U241 ( .A(B[144]), .Z(n401) );
  IV U242 ( .A(B[145]), .Z(n402) );
  IV U243 ( .A(B[146]), .Z(n403) );
  IV U244 ( .A(B[147]), .Z(n404) );
  IV U245 ( .A(B[148]), .Z(n405) );
  IV U246 ( .A(B[247]), .Z(n504) );
  IV U247 ( .A(B[149]), .Z(n406) );
  IV U248 ( .A(B[150]), .Z(n407) );
  IV U249 ( .A(B[151]), .Z(n408) );
  IV U250 ( .A(B[152]), .Z(n409) );
  IV U251 ( .A(B[153]), .Z(n410) );
  IV U252 ( .A(B[154]), .Z(n411) );
  IV U253 ( .A(B[155]), .Z(n412) );
  IV U254 ( .A(B[156]), .Z(n413) );
  IV U255 ( .A(B[157]), .Z(n414) );
  IV U256 ( .A(B[158]), .Z(n415) );
  IV U257 ( .A(B[248]), .Z(n505) );
endmodule


module FA_1291 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XNOR U1 ( .A(CI), .B(A), .Z(S) );
endmodule


module FA_1292 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1293 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1294 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1295 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1296 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1297 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1298 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1299 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1300 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1301 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1302 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1303 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1304 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1305 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1306 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1307 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1308 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1309 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1310 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1311 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1312 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1313 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1314 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1315 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1316 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1317 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1318 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1319 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1320 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1321 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1322 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1323 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1324 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1325 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1326 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1327 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1328 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1329 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1330 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1331 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1332 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1333 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1334 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1335 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1336 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1337 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1338 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1339 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1340 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1341 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1342 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1343 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1344 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1345 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1346 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1347 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1348 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1349 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1350 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1351 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1352 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1353 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1354 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1355 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1356 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1357 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1358 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1359 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1360 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1361 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1362 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1363 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1364 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1365 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1366 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1367 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1368 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1369 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1370 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1371 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1372 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1373 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1374 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1375 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1376 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1377 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1378 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1379 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1380 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1381 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1382 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1383 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1384 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1385 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1386 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1387 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1388 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1389 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1390 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1391 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1392 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1393 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1394 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1395 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1396 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1397 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1398 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1399 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1400 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1401 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1402 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1403 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1404 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1405 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1406 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1407 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1408 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1409 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1410 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1411 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1412 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1413 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1414 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1415 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1416 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1417 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1418 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1419 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1420 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1421 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1422 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1423 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1424 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1425 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1426 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1427 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1428 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1429 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1430 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1431 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1432 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1433 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1434 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1435 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1436 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1437 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1438 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1439 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1440 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1441 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1442 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1443 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1444 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1445 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1446 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1447 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1448 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1449 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1450 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1451 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1452 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1453 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1454 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1455 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1456 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1457 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1458 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1459 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1460 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1461 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1462 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1463 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1464 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1465 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1466 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1467 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1468 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1469 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1470 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1471 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1472 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1473 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1474 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1475 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1476 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1477 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1478 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1479 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1480 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1481 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1482 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1483 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1484 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1485 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1486 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1487 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1488 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1489 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1490 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1491 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1492 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1493 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1494 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1495 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1496 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1497 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1498 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1499 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1500 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1501 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1502 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1503 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1504 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1505 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1506 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1507 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1508 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1509 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1510 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1511 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1512 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1513 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1514 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1515 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1516 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1517 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1518 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1519 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1520 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1521 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1522 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1523 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1524 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1525 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1526 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1527 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1528 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1529 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1530 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1531 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1532 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1533 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1534 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1535 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1536 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1537 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1538 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1539 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1540 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1541 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1542 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1543 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1544 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1545 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1546 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1547 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XNOR U1 ( .A(B), .B(A), .Z(S) );
  OR U2 ( .A(B), .B(A), .Z(CO) );
endmodule


module SUB_N258_3 ( A, B, S, CO );
  input [257:0] A;
  input [257:0] B;
  output [257:0] S;
  output CO;
  wire   n2, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512;
  wire   [257:1] C;

  FA_1547 \FAINST[0].FA_  ( .A(A[0]), .B(n2), .CI(1'b1), .S(S[0]), .CO(C[1])
         );
  FA_1546 \FAINST[1].FA_  ( .A(A[1]), .B(n258), .CI(C[1]), .S(S[1]), .CO(C[2])
         );
  FA_1545 \FAINST[2].FA_  ( .A(A[2]), .B(n259), .CI(C[2]), .S(S[2]), .CO(C[3])
         );
  FA_1544 \FAINST[3].FA_  ( .A(A[3]), .B(n260), .CI(C[3]), .S(S[3]), .CO(C[4])
         );
  FA_1543 \FAINST[4].FA_  ( .A(A[4]), .B(n261), .CI(C[4]), .S(S[4]), .CO(C[5])
         );
  FA_1542 \FAINST[5].FA_  ( .A(A[5]), .B(n262), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_1541 \FAINST[6].FA_  ( .A(A[6]), .B(n263), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_1540 \FAINST[7].FA_  ( .A(A[7]), .B(n264), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_1539 \FAINST[8].FA_  ( .A(A[8]), .B(n265), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_1538 \FAINST[9].FA_  ( .A(A[9]), .B(n266), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_1537 \FAINST[10].FA_  ( .A(A[10]), .B(n267), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_1536 \FAINST[11].FA_  ( .A(A[11]), .B(n268), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_1535 \FAINST[12].FA_  ( .A(A[12]), .B(n269), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_1534 \FAINST[13].FA_  ( .A(A[13]), .B(n270), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_1533 \FAINST[14].FA_  ( .A(A[14]), .B(n271), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_1532 \FAINST[15].FA_  ( .A(A[15]), .B(n272), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_1531 \FAINST[16].FA_  ( .A(A[16]), .B(n273), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_1530 \FAINST[17].FA_  ( .A(A[17]), .B(n274), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_1529 \FAINST[18].FA_  ( .A(A[18]), .B(n275), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_1528 \FAINST[19].FA_  ( .A(A[19]), .B(n276), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_1527 \FAINST[20].FA_  ( .A(A[20]), .B(n277), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_1526 \FAINST[21].FA_  ( .A(A[21]), .B(n278), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_1525 \FAINST[22].FA_  ( .A(A[22]), .B(n279), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_1524 \FAINST[23].FA_  ( .A(A[23]), .B(n280), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1523 \FAINST[24].FA_  ( .A(A[24]), .B(n281), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1522 \FAINST[25].FA_  ( .A(A[25]), .B(n282), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1521 \FAINST[26].FA_  ( .A(A[26]), .B(n283), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1520 \FAINST[27].FA_  ( .A(A[27]), .B(n284), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1519 \FAINST[28].FA_  ( .A(A[28]), .B(n285), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1518 \FAINST[29].FA_  ( .A(A[29]), .B(n286), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1517 \FAINST[30].FA_  ( .A(A[30]), .B(n287), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1516 \FAINST[31].FA_  ( .A(A[31]), .B(n288), .CI(C[31]), .S(S[31]), .CO(
        C[32]) );
  FA_1515 \FAINST[32].FA_  ( .A(A[32]), .B(n289), .CI(C[32]), .S(S[32]), .CO(
        C[33]) );
  FA_1514 \FAINST[33].FA_  ( .A(A[33]), .B(n290), .CI(C[33]), .S(S[33]), .CO(
        C[34]) );
  FA_1513 \FAINST[34].FA_  ( .A(A[34]), .B(n291), .CI(C[34]), .S(S[34]), .CO(
        C[35]) );
  FA_1512 \FAINST[35].FA_  ( .A(A[35]), .B(n292), .CI(C[35]), .S(S[35]), .CO(
        C[36]) );
  FA_1511 \FAINST[36].FA_  ( .A(A[36]), .B(n293), .CI(C[36]), .S(S[36]), .CO(
        C[37]) );
  FA_1510 \FAINST[37].FA_  ( .A(A[37]), .B(n294), .CI(C[37]), .S(S[37]), .CO(
        C[38]) );
  FA_1509 \FAINST[38].FA_  ( .A(A[38]), .B(n295), .CI(C[38]), .S(S[38]), .CO(
        C[39]) );
  FA_1508 \FAINST[39].FA_  ( .A(A[39]), .B(n296), .CI(C[39]), .S(S[39]), .CO(
        C[40]) );
  FA_1507 \FAINST[40].FA_  ( .A(A[40]), .B(n297), .CI(C[40]), .S(S[40]), .CO(
        C[41]) );
  FA_1506 \FAINST[41].FA_  ( .A(A[41]), .B(n298), .CI(C[41]), .S(S[41]), .CO(
        C[42]) );
  FA_1505 \FAINST[42].FA_  ( .A(A[42]), .B(n299), .CI(C[42]), .S(S[42]), .CO(
        C[43]) );
  FA_1504 \FAINST[43].FA_  ( .A(A[43]), .B(n300), .CI(C[43]), .S(S[43]), .CO(
        C[44]) );
  FA_1503 \FAINST[44].FA_  ( .A(A[44]), .B(n301), .CI(C[44]), .S(S[44]), .CO(
        C[45]) );
  FA_1502 \FAINST[45].FA_  ( .A(A[45]), .B(n302), .CI(C[45]), .S(S[45]), .CO(
        C[46]) );
  FA_1501 \FAINST[46].FA_  ( .A(A[46]), .B(n303), .CI(C[46]), .S(S[46]), .CO(
        C[47]) );
  FA_1500 \FAINST[47].FA_  ( .A(A[47]), .B(n304), .CI(C[47]), .S(S[47]), .CO(
        C[48]) );
  FA_1499 \FAINST[48].FA_  ( .A(A[48]), .B(n305), .CI(C[48]), .S(S[48]), .CO(
        C[49]) );
  FA_1498 \FAINST[49].FA_  ( .A(A[49]), .B(n306), .CI(C[49]), .S(S[49]), .CO(
        C[50]) );
  FA_1497 \FAINST[50].FA_  ( .A(A[50]), .B(n307), .CI(C[50]), .S(S[50]), .CO(
        C[51]) );
  FA_1496 \FAINST[51].FA_  ( .A(A[51]), .B(n308), .CI(C[51]), .S(S[51]), .CO(
        C[52]) );
  FA_1495 \FAINST[52].FA_  ( .A(A[52]), .B(n309), .CI(C[52]), .S(S[52]), .CO(
        C[53]) );
  FA_1494 \FAINST[53].FA_  ( .A(A[53]), .B(n310), .CI(C[53]), .S(S[53]), .CO(
        C[54]) );
  FA_1493 \FAINST[54].FA_  ( .A(A[54]), .B(n311), .CI(C[54]), .S(S[54]), .CO(
        C[55]) );
  FA_1492 \FAINST[55].FA_  ( .A(A[55]), .B(n312), .CI(C[55]), .S(S[55]), .CO(
        C[56]) );
  FA_1491 \FAINST[56].FA_  ( .A(A[56]), .B(n313), .CI(C[56]), .S(S[56]), .CO(
        C[57]) );
  FA_1490 \FAINST[57].FA_  ( .A(A[57]), .B(n314), .CI(C[57]), .S(S[57]), .CO(
        C[58]) );
  FA_1489 \FAINST[58].FA_  ( .A(A[58]), .B(n315), .CI(C[58]), .S(S[58]), .CO(
        C[59]) );
  FA_1488 \FAINST[59].FA_  ( .A(A[59]), .B(n316), .CI(C[59]), .S(S[59]), .CO(
        C[60]) );
  FA_1487 \FAINST[60].FA_  ( .A(A[60]), .B(n317), .CI(C[60]), .S(S[60]), .CO(
        C[61]) );
  FA_1486 \FAINST[61].FA_  ( .A(A[61]), .B(n318), .CI(C[61]), .S(S[61]), .CO(
        C[62]) );
  FA_1485 \FAINST[62].FA_  ( .A(A[62]), .B(n319), .CI(C[62]), .S(S[62]), .CO(
        C[63]) );
  FA_1484 \FAINST[63].FA_  ( .A(A[63]), .B(n320), .CI(C[63]), .S(S[63]), .CO(
        C[64]) );
  FA_1483 \FAINST[64].FA_  ( .A(A[64]), .B(n321), .CI(C[64]), .S(S[64]), .CO(
        C[65]) );
  FA_1482 \FAINST[65].FA_  ( .A(A[65]), .B(n322), .CI(C[65]), .S(S[65]), .CO(
        C[66]) );
  FA_1481 \FAINST[66].FA_  ( .A(A[66]), .B(n323), .CI(C[66]), .S(S[66]), .CO(
        C[67]) );
  FA_1480 \FAINST[67].FA_  ( .A(A[67]), .B(n324), .CI(C[67]), .S(S[67]), .CO(
        C[68]) );
  FA_1479 \FAINST[68].FA_  ( .A(A[68]), .B(n325), .CI(C[68]), .S(S[68]), .CO(
        C[69]) );
  FA_1478 \FAINST[69].FA_  ( .A(A[69]), .B(n326), .CI(C[69]), .S(S[69]), .CO(
        C[70]) );
  FA_1477 \FAINST[70].FA_  ( .A(A[70]), .B(n327), .CI(C[70]), .S(S[70]), .CO(
        C[71]) );
  FA_1476 \FAINST[71].FA_  ( .A(A[71]), .B(n328), .CI(C[71]), .S(S[71]), .CO(
        C[72]) );
  FA_1475 \FAINST[72].FA_  ( .A(A[72]), .B(n329), .CI(C[72]), .S(S[72]), .CO(
        C[73]) );
  FA_1474 \FAINST[73].FA_  ( .A(A[73]), .B(n330), .CI(C[73]), .S(S[73]), .CO(
        C[74]) );
  FA_1473 \FAINST[74].FA_  ( .A(A[74]), .B(n331), .CI(C[74]), .S(S[74]), .CO(
        C[75]) );
  FA_1472 \FAINST[75].FA_  ( .A(A[75]), .B(n332), .CI(C[75]), .S(S[75]), .CO(
        C[76]) );
  FA_1471 \FAINST[76].FA_  ( .A(A[76]), .B(n333), .CI(C[76]), .S(S[76]), .CO(
        C[77]) );
  FA_1470 \FAINST[77].FA_  ( .A(A[77]), .B(n334), .CI(C[77]), .S(S[77]), .CO(
        C[78]) );
  FA_1469 \FAINST[78].FA_  ( .A(A[78]), .B(n335), .CI(C[78]), .S(S[78]), .CO(
        C[79]) );
  FA_1468 \FAINST[79].FA_  ( .A(A[79]), .B(n336), .CI(C[79]), .S(S[79]), .CO(
        C[80]) );
  FA_1467 \FAINST[80].FA_  ( .A(A[80]), .B(n337), .CI(C[80]), .S(S[80]), .CO(
        C[81]) );
  FA_1466 \FAINST[81].FA_  ( .A(A[81]), .B(n338), .CI(C[81]), .S(S[81]), .CO(
        C[82]) );
  FA_1465 \FAINST[82].FA_  ( .A(A[82]), .B(n339), .CI(C[82]), .S(S[82]), .CO(
        C[83]) );
  FA_1464 \FAINST[83].FA_  ( .A(A[83]), .B(n340), .CI(C[83]), .S(S[83]), .CO(
        C[84]) );
  FA_1463 \FAINST[84].FA_  ( .A(A[84]), .B(n341), .CI(C[84]), .S(S[84]), .CO(
        C[85]) );
  FA_1462 \FAINST[85].FA_  ( .A(A[85]), .B(n342), .CI(C[85]), .S(S[85]), .CO(
        C[86]) );
  FA_1461 \FAINST[86].FA_  ( .A(A[86]), .B(n343), .CI(C[86]), .S(S[86]), .CO(
        C[87]) );
  FA_1460 \FAINST[87].FA_  ( .A(A[87]), .B(n344), .CI(C[87]), .S(S[87]), .CO(
        C[88]) );
  FA_1459 \FAINST[88].FA_  ( .A(A[88]), .B(n345), .CI(C[88]), .S(S[88]), .CO(
        C[89]) );
  FA_1458 \FAINST[89].FA_  ( .A(A[89]), .B(n346), .CI(C[89]), .S(S[89]), .CO(
        C[90]) );
  FA_1457 \FAINST[90].FA_  ( .A(A[90]), .B(n347), .CI(C[90]), .S(S[90]), .CO(
        C[91]) );
  FA_1456 \FAINST[91].FA_  ( .A(A[91]), .B(n348), .CI(C[91]), .S(S[91]), .CO(
        C[92]) );
  FA_1455 \FAINST[92].FA_  ( .A(A[92]), .B(n349), .CI(C[92]), .S(S[92]), .CO(
        C[93]) );
  FA_1454 \FAINST[93].FA_  ( .A(A[93]), .B(n350), .CI(C[93]), .S(S[93]), .CO(
        C[94]) );
  FA_1453 \FAINST[94].FA_  ( .A(A[94]), .B(n351), .CI(C[94]), .S(S[94]), .CO(
        C[95]) );
  FA_1452 \FAINST[95].FA_  ( .A(A[95]), .B(n352), .CI(C[95]), .S(S[95]), .CO(
        C[96]) );
  FA_1451 \FAINST[96].FA_  ( .A(A[96]), .B(n353), .CI(C[96]), .S(S[96]), .CO(
        C[97]) );
  FA_1450 \FAINST[97].FA_  ( .A(A[97]), .B(n354), .CI(C[97]), .S(S[97]), .CO(
        C[98]) );
  FA_1449 \FAINST[98].FA_  ( .A(A[98]), .B(n355), .CI(C[98]), .S(S[98]), .CO(
        C[99]) );
  FA_1448 \FAINST[99].FA_  ( .A(A[99]), .B(n356), .CI(C[99]), .S(S[99]), .CO(
        C[100]) );
  FA_1447 \FAINST[100].FA_  ( .A(A[100]), .B(n357), .CI(C[100]), .S(S[100]), 
        .CO(C[101]) );
  FA_1446 \FAINST[101].FA_  ( .A(A[101]), .B(n358), .CI(C[101]), .S(S[101]), 
        .CO(C[102]) );
  FA_1445 \FAINST[102].FA_  ( .A(A[102]), .B(n359), .CI(C[102]), .S(S[102]), 
        .CO(C[103]) );
  FA_1444 \FAINST[103].FA_  ( .A(A[103]), .B(n360), .CI(C[103]), .S(S[103]), 
        .CO(C[104]) );
  FA_1443 \FAINST[104].FA_  ( .A(A[104]), .B(n361), .CI(C[104]), .S(S[104]), 
        .CO(C[105]) );
  FA_1442 \FAINST[105].FA_  ( .A(A[105]), .B(n362), .CI(C[105]), .S(S[105]), 
        .CO(C[106]) );
  FA_1441 \FAINST[106].FA_  ( .A(A[106]), .B(n363), .CI(C[106]), .S(S[106]), 
        .CO(C[107]) );
  FA_1440 \FAINST[107].FA_  ( .A(A[107]), .B(n364), .CI(C[107]), .S(S[107]), 
        .CO(C[108]) );
  FA_1439 \FAINST[108].FA_  ( .A(A[108]), .B(n365), .CI(C[108]), .S(S[108]), 
        .CO(C[109]) );
  FA_1438 \FAINST[109].FA_  ( .A(A[109]), .B(n366), .CI(C[109]), .S(S[109]), 
        .CO(C[110]) );
  FA_1437 \FAINST[110].FA_  ( .A(A[110]), .B(n367), .CI(C[110]), .S(S[110]), 
        .CO(C[111]) );
  FA_1436 \FAINST[111].FA_  ( .A(A[111]), .B(n368), .CI(C[111]), .S(S[111]), 
        .CO(C[112]) );
  FA_1435 \FAINST[112].FA_  ( .A(A[112]), .B(n369), .CI(C[112]), .S(S[112]), 
        .CO(C[113]) );
  FA_1434 \FAINST[113].FA_  ( .A(A[113]), .B(n370), .CI(C[113]), .S(S[113]), 
        .CO(C[114]) );
  FA_1433 \FAINST[114].FA_  ( .A(A[114]), .B(n371), .CI(C[114]), .S(S[114]), 
        .CO(C[115]) );
  FA_1432 \FAINST[115].FA_  ( .A(A[115]), .B(n372), .CI(C[115]), .S(S[115]), 
        .CO(C[116]) );
  FA_1431 \FAINST[116].FA_  ( .A(A[116]), .B(n373), .CI(C[116]), .S(S[116]), 
        .CO(C[117]) );
  FA_1430 \FAINST[117].FA_  ( .A(A[117]), .B(n374), .CI(C[117]), .S(S[117]), 
        .CO(C[118]) );
  FA_1429 \FAINST[118].FA_  ( .A(A[118]), .B(n375), .CI(C[118]), .S(S[118]), 
        .CO(C[119]) );
  FA_1428 \FAINST[119].FA_  ( .A(A[119]), .B(n376), .CI(C[119]), .S(S[119]), 
        .CO(C[120]) );
  FA_1427 \FAINST[120].FA_  ( .A(A[120]), .B(n377), .CI(C[120]), .S(S[120]), 
        .CO(C[121]) );
  FA_1426 \FAINST[121].FA_  ( .A(A[121]), .B(n378), .CI(C[121]), .S(S[121]), 
        .CO(C[122]) );
  FA_1425 \FAINST[122].FA_  ( .A(A[122]), .B(n379), .CI(C[122]), .S(S[122]), 
        .CO(C[123]) );
  FA_1424 \FAINST[123].FA_  ( .A(A[123]), .B(n380), .CI(C[123]), .S(S[123]), 
        .CO(C[124]) );
  FA_1423 \FAINST[124].FA_  ( .A(A[124]), .B(n381), .CI(C[124]), .S(S[124]), 
        .CO(C[125]) );
  FA_1422 \FAINST[125].FA_  ( .A(A[125]), .B(n382), .CI(C[125]), .S(S[125]), 
        .CO(C[126]) );
  FA_1421 \FAINST[126].FA_  ( .A(A[126]), .B(n383), .CI(C[126]), .S(S[126]), 
        .CO(C[127]) );
  FA_1420 \FAINST[127].FA_  ( .A(A[127]), .B(n384), .CI(C[127]), .S(S[127]), 
        .CO(C[128]) );
  FA_1419 \FAINST[128].FA_  ( .A(A[128]), .B(n385), .CI(C[128]), .S(S[128]), 
        .CO(C[129]) );
  FA_1418 \FAINST[129].FA_  ( .A(A[129]), .B(n386), .CI(C[129]), .S(S[129]), 
        .CO(C[130]) );
  FA_1417 \FAINST[130].FA_  ( .A(A[130]), .B(n387), .CI(C[130]), .S(S[130]), 
        .CO(C[131]) );
  FA_1416 \FAINST[131].FA_  ( .A(A[131]), .B(n388), .CI(C[131]), .S(S[131]), 
        .CO(C[132]) );
  FA_1415 \FAINST[132].FA_  ( .A(A[132]), .B(n389), .CI(C[132]), .S(S[132]), 
        .CO(C[133]) );
  FA_1414 \FAINST[133].FA_  ( .A(A[133]), .B(n390), .CI(C[133]), .S(S[133]), 
        .CO(C[134]) );
  FA_1413 \FAINST[134].FA_  ( .A(A[134]), .B(n391), .CI(C[134]), .S(S[134]), 
        .CO(C[135]) );
  FA_1412 \FAINST[135].FA_  ( .A(A[135]), .B(n392), .CI(C[135]), .S(S[135]), 
        .CO(C[136]) );
  FA_1411 \FAINST[136].FA_  ( .A(A[136]), .B(n393), .CI(C[136]), .S(S[136]), 
        .CO(C[137]) );
  FA_1410 \FAINST[137].FA_  ( .A(A[137]), .B(n394), .CI(C[137]), .S(S[137]), 
        .CO(C[138]) );
  FA_1409 \FAINST[138].FA_  ( .A(A[138]), .B(n395), .CI(C[138]), .S(S[138]), 
        .CO(C[139]) );
  FA_1408 \FAINST[139].FA_  ( .A(A[139]), .B(n396), .CI(C[139]), .S(S[139]), 
        .CO(C[140]) );
  FA_1407 \FAINST[140].FA_  ( .A(A[140]), .B(n397), .CI(C[140]), .S(S[140]), 
        .CO(C[141]) );
  FA_1406 \FAINST[141].FA_  ( .A(A[141]), .B(n398), .CI(C[141]), .S(S[141]), 
        .CO(C[142]) );
  FA_1405 \FAINST[142].FA_  ( .A(A[142]), .B(n399), .CI(C[142]), .S(S[142]), 
        .CO(C[143]) );
  FA_1404 \FAINST[143].FA_  ( .A(A[143]), .B(n400), .CI(C[143]), .S(S[143]), 
        .CO(C[144]) );
  FA_1403 \FAINST[144].FA_  ( .A(A[144]), .B(n401), .CI(C[144]), .S(S[144]), 
        .CO(C[145]) );
  FA_1402 \FAINST[145].FA_  ( .A(A[145]), .B(n402), .CI(C[145]), .S(S[145]), 
        .CO(C[146]) );
  FA_1401 \FAINST[146].FA_  ( .A(A[146]), .B(n403), .CI(C[146]), .S(S[146]), 
        .CO(C[147]) );
  FA_1400 \FAINST[147].FA_  ( .A(A[147]), .B(n404), .CI(C[147]), .S(S[147]), 
        .CO(C[148]) );
  FA_1399 \FAINST[148].FA_  ( .A(A[148]), .B(n405), .CI(C[148]), .S(S[148]), 
        .CO(C[149]) );
  FA_1398 \FAINST[149].FA_  ( .A(A[149]), .B(n406), .CI(C[149]), .S(S[149]), 
        .CO(C[150]) );
  FA_1397 \FAINST[150].FA_  ( .A(A[150]), .B(n407), .CI(C[150]), .S(S[150]), 
        .CO(C[151]) );
  FA_1396 \FAINST[151].FA_  ( .A(A[151]), .B(n408), .CI(C[151]), .S(S[151]), 
        .CO(C[152]) );
  FA_1395 \FAINST[152].FA_  ( .A(A[152]), .B(n409), .CI(C[152]), .S(S[152]), 
        .CO(C[153]) );
  FA_1394 \FAINST[153].FA_  ( .A(A[153]), .B(n410), .CI(C[153]), .S(S[153]), 
        .CO(C[154]) );
  FA_1393 \FAINST[154].FA_  ( .A(A[154]), .B(n411), .CI(C[154]), .S(S[154]), 
        .CO(C[155]) );
  FA_1392 \FAINST[155].FA_  ( .A(A[155]), .B(n412), .CI(C[155]), .S(S[155]), 
        .CO(C[156]) );
  FA_1391 \FAINST[156].FA_  ( .A(A[156]), .B(n413), .CI(C[156]), .S(S[156]), 
        .CO(C[157]) );
  FA_1390 \FAINST[157].FA_  ( .A(A[157]), .B(n414), .CI(C[157]), .S(S[157]), 
        .CO(C[158]) );
  FA_1389 \FAINST[158].FA_  ( .A(A[158]), .B(n415), .CI(C[158]), .S(S[158]), 
        .CO(C[159]) );
  FA_1388 \FAINST[159].FA_  ( .A(A[159]), .B(n416), .CI(C[159]), .S(S[159]), 
        .CO(C[160]) );
  FA_1387 \FAINST[160].FA_  ( .A(A[160]), .B(n417), .CI(C[160]), .S(S[160]), 
        .CO(C[161]) );
  FA_1386 \FAINST[161].FA_  ( .A(A[161]), .B(n418), .CI(C[161]), .S(S[161]), 
        .CO(C[162]) );
  FA_1385 \FAINST[162].FA_  ( .A(A[162]), .B(n419), .CI(C[162]), .S(S[162]), 
        .CO(C[163]) );
  FA_1384 \FAINST[163].FA_  ( .A(A[163]), .B(n420), .CI(C[163]), .S(S[163]), 
        .CO(C[164]) );
  FA_1383 \FAINST[164].FA_  ( .A(A[164]), .B(n421), .CI(C[164]), .S(S[164]), 
        .CO(C[165]) );
  FA_1382 \FAINST[165].FA_  ( .A(A[165]), .B(n422), .CI(C[165]), .S(S[165]), 
        .CO(C[166]) );
  FA_1381 \FAINST[166].FA_  ( .A(A[166]), .B(n423), .CI(C[166]), .S(S[166]), 
        .CO(C[167]) );
  FA_1380 \FAINST[167].FA_  ( .A(A[167]), .B(n424), .CI(C[167]), .S(S[167]), 
        .CO(C[168]) );
  FA_1379 \FAINST[168].FA_  ( .A(A[168]), .B(n425), .CI(C[168]), .S(S[168]), 
        .CO(C[169]) );
  FA_1378 \FAINST[169].FA_  ( .A(A[169]), .B(n426), .CI(C[169]), .S(S[169]), 
        .CO(C[170]) );
  FA_1377 \FAINST[170].FA_  ( .A(A[170]), .B(n427), .CI(C[170]), .S(S[170]), 
        .CO(C[171]) );
  FA_1376 \FAINST[171].FA_  ( .A(A[171]), .B(n428), .CI(C[171]), .S(S[171]), 
        .CO(C[172]) );
  FA_1375 \FAINST[172].FA_  ( .A(A[172]), .B(n429), .CI(C[172]), .S(S[172]), 
        .CO(C[173]) );
  FA_1374 \FAINST[173].FA_  ( .A(A[173]), .B(n430), .CI(C[173]), .S(S[173]), 
        .CO(C[174]) );
  FA_1373 \FAINST[174].FA_  ( .A(A[174]), .B(n431), .CI(C[174]), .S(S[174]), 
        .CO(C[175]) );
  FA_1372 \FAINST[175].FA_  ( .A(A[175]), .B(n432), .CI(C[175]), .S(S[175]), 
        .CO(C[176]) );
  FA_1371 \FAINST[176].FA_  ( .A(A[176]), .B(n433), .CI(C[176]), .S(S[176]), 
        .CO(C[177]) );
  FA_1370 \FAINST[177].FA_  ( .A(A[177]), .B(n434), .CI(C[177]), .S(S[177]), 
        .CO(C[178]) );
  FA_1369 \FAINST[178].FA_  ( .A(A[178]), .B(n435), .CI(C[178]), .S(S[178]), 
        .CO(C[179]) );
  FA_1368 \FAINST[179].FA_  ( .A(A[179]), .B(n436), .CI(C[179]), .S(S[179]), 
        .CO(C[180]) );
  FA_1367 \FAINST[180].FA_  ( .A(A[180]), .B(n437), .CI(C[180]), .S(S[180]), 
        .CO(C[181]) );
  FA_1366 \FAINST[181].FA_  ( .A(A[181]), .B(n438), .CI(C[181]), .S(S[181]), 
        .CO(C[182]) );
  FA_1365 \FAINST[182].FA_  ( .A(A[182]), .B(n439), .CI(C[182]), .S(S[182]), 
        .CO(C[183]) );
  FA_1364 \FAINST[183].FA_  ( .A(A[183]), .B(n440), .CI(C[183]), .S(S[183]), 
        .CO(C[184]) );
  FA_1363 \FAINST[184].FA_  ( .A(A[184]), .B(n441), .CI(C[184]), .S(S[184]), 
        .CO(C[185]) );
  FA_1362 \FAINST[185].FA_  ( .A(A[185]), .B(n442), .CI(C[185]), .S(S[185]), 
        .CO(C[186]) );
  FA_1361 \FAINST[186].FA_  ( .A(A[186]), .B(n443), .CI(C[186]), .S(S[186]), 
        .CO(C[187]) );
  FA_1360 \FAINST[187].FA_  ( .A(A[187]), .B(n444), .CI(C[187]), .S(S[187]), 
        .CO(C[188]) );
  FA_1359 \FAINST[188].FA_  ( .A(A[188]), .B(n445), .CI(C[188]), .S(S[188]), 
        .CO(C[189]) );
  FA_1358 \FAINST[189].FA_  ( .A(A[189]), .B(n446), .CI(C[189]), .S(S[189]), 
        .CO(C[190]) );
  FA_1357 \FAINST[190].FA_  ( .A(A[190]), .B(n447), .CI(C[190]), .S(S[190]), 
        .CO(C[191]) );
  FA_1356 \FAINST[191].FA_  ( .A(A[191]), .B(n448), .CI(C[191]), .S(S[191]), 
        .CO(C[192]) );
  FA_1355 \FAINST[192].FA_  ( .A(A[192]), .B(n449), .CI(C[192]), .S(S[192]), 
        .CO(C[193]) );
  FA_1354 \FAINST[193].FA_  ( .A(A[193]), .B(n450), .CI(C[193]), .S(S[193]), 
        .CO(C[194]) );
  FA_1353 \FAINST[194].FA_  ( .A(A[194]), .B(n451), .CI(C[194]), .S(S[194]), 
        .CO(C[195]) );
  FA_1352 \FAINST[195].FA_  ( .A(A[195]), .B(n452), .CI(C[195]), .S(S[195]), 
        .CO(C[196]) );
  FA_1351 \FAINST[196].FA_  ( .A(A[196]), .B(n453), .CI(C[196]), .S(S[196]), 
        .CO(C[197]) );
  FA_1350 \FAINST[197].FA_  ( .A(A[197]), .B(n454), .CI(C[197]), .S(S[197]), 
        .CO(C[198]) );
  FA_1349 \FAINST[198].FA_  ( .A(A[198]), .B(n455), .CI(C[198]), .S(S[198]), 
        .CO(C[199]) );
  FA_1348 \FAINST[199].FA_  ( .A(A[199]), .B(n456), .CI(C[199]), .S(S[199]), 
        .CO(C[200]) );
  FA_1347 \FAINST[200].FA_  ( .A(A[200]), .B(n457), .CI(C[200]), .S(S[200]), 
        .CO(C[201]) );
  FA_1346 \FAINST[201].FA_  ( .A(A[201]), .B(n458), .CI(C[201]), .S(S[201]), 
        .CO(C[202]) );
  FA_1345 \FAINST[202].FA_  ( .A(A[202]), .B(n459), .CI(C[202]), .S(S[202]), 
        .CO(C[203]) );
  FA_1344 \FAINST[203].FA_  ( .A(A[203]), .B(n460), .CI(C[203]), .S(S[203]), 
        .CO(C[204]) );
  FA_1343 \FAINST[204].FA_  ( .A(A[204]), .B(n461), .CI(C[204]), .S(S[204]), 
        .CO(C[205]) );
  FA_1342 \FAINST[205].FA_  ( .A(A[205]), .B(n462), .CI(C[205]), .S(S[205]), 
        .CO(C[206]) );
  FA_1341 \FAINST[206].FA_  ( .A(A[206]), .B(n463), .CI(C[206]), .S(S[206]), 
        .CO(C[207]) );
  FA_1340 \FAINST[207].FA_  ( .A(A[207]), .B(n464), .CI(C[207]), .S(S[207]), 
        .CO(C[208]) );
  FA_1339 \FAINST[208].FA_  ( .A(A[208]), .B(n465), .CI(C[208]), .S(S[208]), 
        .CO(C[209]) );
  FA_1338 \FAINST[209].FA_  ( .A(A[209]), .B(n466), .CI(C[209]), .S(S[209]), 
        .CO(C[210]) );
  FA_1337 \FAINST[210].FA_  ( .A(A[210]), .B(n467), .CI(C[210]), .S(S[210]), 
        .CO(C[211]) );
  FA_1336 \FAINST[211].FA_  ( .A(A[211]), .B(n468), .CI(C[211]), .S(S[211]), 
        .CO(C[212]) );
  FA_1335 \FAINST[212].FA_  ( .A(A[212]), .B(n469), .CI(C[212]), .S(S[212]), 
        .CO(C[213]) );
  FA_1334 \FAINST[213].FA_  ( .A(A[213]), .B(n470), .CI(C[213]), .S(S[213]), 
        .CO(C[214]) );
  FA_1333 \FAINST[214].FA_  ( .A(A[214]), .B(n471), .CI(C[214]), .S(S[214]), 
        .CO(C[215]) );
  FA_1332 \FAINST[215].FA_  ( .A(A[215]), .B(n472), .CI(C[215]), .S(S[215]), 
        .CO(C[216]) );
  FA_1331 \FAINST[216].FA_  ( .A(A[216]), .B(n473), .CI(C[216]), .S(S[216]), 
        .CO(C[217]) );
  FA_1330 \FAINST[217].FA_  ( .A(A[217]), .B(n474), .CI(C[217]), .S(S[217]), 
        .CO(C[218]) );
  FA_1329 \FAINST[218].FA_  ( .A(A[218]), .B(n475), .CI(C[218]), .S(S[218]), 
        .CO(C[219]) );
  FA_1328 \FAINST[219].FA_  ( .A(A[219]), .B(n476), .CI(C[219]), .S(S[219]), 
        .CO(C[220]) );
  FA_1327 \FAINST[220].FA_  ( .A(A[220]), .B(n477), .CI(C[220]), .S(S[220]), 
        .CO(C[221]) );
  FA_1326 \FAINST[221].FA_  ( .A(A[221]), .B(n478), .CI(C[221]), .S(S[221]), 
        .CO(C[222]) );
  FA_1325 \FAINST[222].FA_  ( .A(A[222]), .B(n479), .CI(C[222]), .S(S[222]), 
        .CO(C[223]) );
  FA_1324 \FAINST[223].FA_  ( .A(A[223]), .B(n480), .CI(C[223]), .S(S[223]), 
        .CO(C[224]) );
  FA_1323 \FAINST[224].FA_  ( .A(A[224]), .B(n481), .CI(C[224]), .S(S[224]), 
        .CO(C[225]) );
  FA_1322 \FAINST[225].FA_  ( .A(A[225]), .B(n482), .CI(C[225]), .S(S[225]), 
        .CO(C[226]) );
  FA_1321 \FAINST[226].FA_  ( .A(A[226]), .B(n483), .CI(C[226]), .S(S[226]), 
        .CO(C[227]) );
  FA_1320 \FAINST[227].FA_  ( .A(A[227]), .B(n484), .CI(C[227]), .S(S[227]), 
        .CO(C[228]) );
  FA_1319 \FAINST[228].FA_  ( .A(A[228]), .B(n485), .CI(C[228]), .S(S[228]), 
        .CO(C[229]) );
  FA_1318 \FAINST[229].FA_  ( .A(A[229]), .B(n486), .CI(C[229]), .S(S[229]), 
        .CO(C[230]) );
  FA_1317 \FAINST[230].FA_  ( .A(A[230]), .B(n487), .CI(C[230]), .S(S[230]), 
        .CO(C[231]) );
  FA_1316 \FAINST[231].FA_  ( .A(A[231]), .B(n488), .CI(C[231]), .S(S[231]), 
        .CO(C[232]) );
  FA_1315 \FAINST[232].FA_  ( .A(A[232]), .B(n489), .CI(C[232]), .S(S[232]), 
        .CO(C[233]) );
  FA_1314 \FAINST[233].FA_  ( .A(A[233]), .B(n490), .CI(C[233]), .S(S[233]), 
        .CO(C[234]) );
  FA_1313 \FAINST[234].FA_  ( .A(A[234]), .B(n491), .CI(C[234]), .S(S[234]), 
        .CO(C[235]) );
  FA_1312 \FAINST[235].FA_  ( .A(A[235]), .B(n492), .CI(C[235]), .S(S[235]), 
        .CO(C[236]) );
  FA_1311 \FAINST[236].FA_  ( .A(A[236]), .B(n493), .CI(C[236]), .S(S[236]), 
        .CO(C[237]) );
  FA_1310 \FAINST[237].FA_  ( .A(A[237]), .B(n494), .CI(C[237]), .S(S[237]), 
        .CO(C[238]) );
  FA_1309 \FAINST[238].FA_  ( .A(A[238]), .B(n495), .CI(C[238]), .S(S[238]), 
        .CO(C[239]) );
  FA_1308 \FAINST[239].FA_  ( .A(A[239]), .B(n496), .CI(C[239]), .S(S[239]), 
        .CO(C[240]) );
  FA_1307 \FAINST[240].FA_  ( .A(A[240]), .B(n497), .CI(C[240]), .S(S[240]), 
        .CO(C[241]) );
  FA_1306 \FAINST[241].FA_  ( .A(A[241]), .B(n498), .CI(C[241]), .S(S[241]), 
        .CO(C[242]) );
  FA_1305 \FAINST[242].FA_  ( .A(A[242]), .B(n499), .CI(C[242]), .S(S[242]), 
        .CO(C[243]) );
  FA_1304 \FAINST[243].FA_  ( .A(A[243]), .B(n500), .CI(C[243]), .S(S[243]), 
        .CO(C[244]) );
  FA_1303 \FAINST[244].FA_  ( .A(A[244]), .B(n501), .CI(C[244]), .S(S[244]), 
        .CO(C[245]) );
  FA_1302 \FAINST[245].FA_  ( .A(A[245]), .B(n502), .CI(C[245]), .S(S[245]), 
        .CO(C[246]) );
  FA_1301 \FAINST[246].FA_  ( .A(A[246]), .B(n503), .CI(C[246]), .S(S[246]), 
        .CO(C[247]) );
  FA_1300 \FAINST[247].FA_  ( .A(A[247]), .B(n504), .CI(C[247]), .S(S[247]), 
        .CO(C[248]) );
  FA_1299 \FAINST[248].FA_  ( .A(A[248]), .B(n505), .CI(C[248]), .S(S[248]), 
        .CO(C[249]) );
  FA_1298 \FAINST[249].FA_  ( .A(A[249]), .B(n506), .CI(C[249]), .S(S[249]), 
        .CO(C[250]) );
  FA_1297 \FAINST[250].FA_  ( .A(A[250]), .B(n507), .CI(C[250]), .S(S[250]), 
        .CO(C[251]) );
  FA_1296 \FAINST[251].FA_  ( .A(A[251]), .B(n508), .CI(C[251]), .S(S[251]), 
        .CO(C[252]) );
  FA_1295 \FAINST[252].FA_  ( .A(A[252]), .B(n509), .CI(C[252]), .S(S[252]), 
        .CO(C[253]) );
  FA_1294 \FAINST[253].FA_  ( .A(A[253]), .B(n510), .CI(C[253]), .S(S[253]), 
        .CO(C[254]) );
  FA_1293 \FAINST[254].FA_  ( .A(A[254]), .B(n511), .CI(C[254]), .S(S[254]), 
        .CO(C[255]) );
  FA_1292 \FAINST[255].FA_  ( .A(A[255]), .B(n512), .CI(C[255]), .S(S[255]), 
        .CO(C[256]) );
  FA_1291 \FAINST[256].FA_  ( .A(A[256]), .B(1'b1), .CI(C[256]), .S(S[256]) );
  IV U2 ( .A(B[159]), .Z(n416) );
  IV U3 ( .A(B[160]), .Z(n417) );
  IV U4 ( .A(B[161]), .Z(n418) );
  IV U5 ( .A(B[162]), .Z(n419) );
  IV U6 ( .A(B[163]), .Z(n420) );
  IV U7 ( .A(B[164]), .Z(n421) );
  IV U8 ( .A(B[165]), .Z(n422) );
  IV U9 ( .A(B[166]), .Z(n423) );
  IV U10 ( .A(B[167]), .Z(n424) );
  IV U11 ( .A(B[168]), .Z(n425) );
  IV U12 ( .A(B[249]), .Z(n506) );
  IV U13 ( .A(B[169]), .Z(n426) );
  IV U14 ( .A(B[170]), .Z(n427) );
  IV U15 ( .A(B[171]), .Z(n428) );
  IV U16 ( .A(B[172]), .Z(n429) );
  IV U17 ( .A(B[173]), .Z(n430) );
  IV U18 ( .A(B[174]), .Z(n431) );
  IV U19 ( .A(B[175]), .Z(n432) );
  IV U20 ( .A(B[176]), .Z(n433) );
  IV U21 ( .A(B[177]), .Z(n434) );
  IV U22 ( .A(B[178]), .Z(n435) );
  IV U23 ( .A(B[250]), .Z(n507) );
  IV U24 ( .A(B[179]), .Z(n436) );
  IV U25 ( .A(B[180]), .Z(n437) );
  IV U26 ( .A(B[181]), .Z(n438) );
  IV U27 ( .A(B[182]), .Z(n439) );
  IV U28 ( .A(B[183]), .Z(n440) );
  IV U29 ( .A(B[184]), .Z(n441) );
  IV U30 ( .A(B[185]), .Z(n442) );
  IV U31 ( .A(B[186]), .Z(n443) );
  IV U32 ( .A(B[187]), .Z(n444) );
  IV U33 ( .A(B[188]), .Z(n445) );
  IV U34 ( .A(B[251]), .Z(n508) );
  IV U35 ( .A(B[189]), .Z(n446) );
  IV U36 ( .A(B[190]), .Z(n447) );
  IV U37 ( .A(B[191]), .Z(n448) );
  IV U38 ( .A(B[192]), .Z(n449) );
  IV U39 ( .A(B[193]), .Z(n450) );
  IV U40 ( .A(B[194]), .Z(n451) );
  IV U41 ( .A(B[195]), .Z(n452) );
  IV U42 ( .A(B[196]), .Z(n453) );
  IV U43 ( .A(B[197]), .Z(n454) );
  IV U44 ( .A(B[198]), .Z(n455) );
  IV U45 ( .A(B[252]), .Z(n509) );
  IV U46 ( .A(B[199]), .Z(n456) );
  IV U47 ( .A(B[200]), .Z(n457) );
  IV U48 ( .A(B[201]), .Z(n458) );
  IV U49 ( .A(B[202]), .Z(n459) );
  IV U50 ( .A(B[203]), .Z(n460) );
  IV U51 ( .A(B[204]), .Z(n461) );
  IV U52 ( .A(B[205]), .Z(n462) );
  IV U53 ( .A(B[206]), .Z(n463) );
  IV U54 ( .A(B[207]), .Z(n464) );
  IV U55 ( .A(B[208]), .Z(n465) );
  IV U56 ( .A(B[253]), .Z(n510) );
  IV U57 ( .A(B[209]), .Z(n466) );
  IV U58 ( .A(B[210]), .Z(n467) );
  IV U59 ( .A(B[211]), .Z(n468) );
  IV U60 ( .A(B[212]), .Z(n469) );
  IV U61 ( .A(B[213]), .Z(n470) );
  IV U62 ( .A(B[214]), .Z(n471) );
  IV U63 ( .A(B[215]), .Z(n472) );
  IV U64 ( .A(B[216]), .Z(n473) );
  IV U65 ( .A(B[217]), .Z(n474) );
  IV U66 ( .A(B[218]), .Z(n475) );
  IV U67 ( .A(B[254]), .Z(n511) );
  IV U68 ( .A(B[219]), .Z(n476) );
  IV U69 ( .A(B[220]), .Z(n477) );
  IV U70 ( .A(B[221]), .Z(n478) );
  IV U71 ( .A(B[222]), .Z(n479) );
  IV U72 ( .A(B[223]), .Z(n480) );
  IV U73 ( .A(B[224]), .Z(n481) );
  IV U74 ( .A(B[225]), .Z(n482) );
  IV U75 ( .A(B[226]), .Z(n483) );
  IV U76 ( .A(B[227]), .Z(n484) );
  IV U77 ( .A(B[228]), .Z(n485) );
  IV U78 ( .A(B[255]), .Z(n512) );
  IV U79 ( .A(B[229]), .Z(n486) );
  IV U80 ( .A(B[230]), .Z(n487) );
  IV U81 ( .A(B[231]), .Z(n488) );
  IV U82 ( .A(B[232]), .Z(n489) );
  IV U83 ( .A(B[0]), .Z(n2) );
  IV U84 ( .A(B[1]), .Z(n258) );
  IV U85 ( .A(B[2]), .Z(n259) );
  IV U86 ( .A(B[3]), .Z(n260) );
  IV U87 ( .A(B[4]), .Z(n261) );
  IV U88 ( .A(B[5]), .Z(n262) );
  IV U89 ( .A(B[6]), .Z(n263) );
  IV U90 ( .A(B[7]), .Z(n264) );
  IV U91 ( .A(B[8]), .Z(n265) );
  IV U92 ( .A(B[233]), .Z(n490) );
  IV U93 ( .A(B[9]), .Z(n266) );
  IV U94 ( .A(B[10]), .Z(n267) );
  IV U95 ( .A(B[11]), .Z(n268) );
  IV U96 ( .A(B[12]), .Z(n269) );
  IV U97 ( .A(B[13]), .Z(n270) );
  IV U98 ( .A(B[14]), .Z(n271) );
  IV U99 ( .A(B[15]), .Z(n272) );
  IV U100 ( .A(B[16]), .Z(n273) );
  IV U101 ( .A(B[17]), .Z(n274) );
  IV U102 ( .A(B[18]), .Z(n275) );
  IV U103 ( .A(B[234]), .Z(n491) );
  IV U104 ( .A(B[19]), .Z(n276) );
  IV U105 ( .A(B[20]), .Z(n277) );
  IV U106 ( .A(B[21]), .Z(n278) );
  IV U107 ( .A(B[22]), .Z(n279) );
  IV U108 ( .A(B[23]), .Z(n280) );
  IV U109 ( .A(B[24]), .Z(n281) );
  IV U110 ( .A(B[25]), .Z(n282) );
  IV U111 ( .A(B[26]), .Z(n283) );
  IV U112 ( .A(B[27]), .Z(n284) );
  IV U113 ( .A(B[28]), .Z(n285) );
  IV U114 ( .A(B[235]), .Z(n492) );
  IV U115 ( .A(B[29]), .Z(n286) );
  IV U116 ( .A(B[30]), .Z(n287) );
  IV U117 ( .A(B[31]), .Z(n288) );
  IV U118 ( .A(B[32]), .Z(n289) );
  IV U119 ( .A(B[33]), .Z(n290) );
  IV U120 ( .A(B[34]), .Z(n291) );
  IV U121 ( .A(B[35]), .Z(n292) );
  IV U122 ( .A(B[36]), .Z(n293) );
  IV U123 ( .A(B[37]), .Z(n294) );
  IV U124 ( .A(B[38]), .Z(n295) );
  IV U125 ( .A(B[236]), .Z(n493) );
  IV U126 ( .A(B[39]), .Z(n296) );
  IV U127 ( .A(B[40]), .Z(n297) );
  IV U128 ( .A(B[41]), .Z(n298) );
  IV U129 ( .A(B[42]), .Z(n299) );
  IV U130 ( .A(B[43]), .Z(n300) );
  IV U131 ( .A(B[44]), .Z(n301) );
  IV U132 ( .A(B[45]), .Z(n302) );
  IV U133 ( .A(B[46]), .Z(n303) );
  IV U134 ( .A(B[47]), .Z(n304) );
  IV U135 ( .A(B[48]), .Z(n305) );
  IV U136 ( .A(B[237]), .Z(n494) );
  IV U137 ( .A(B[49]), .Z(n306) );
  IV U138 ( .A(B[50]), .Z(n307) );
  IV U139 ( .A(B[51]), .Z(n308) );
  IV U140 ( .A(B[52]), .Z(n309) );
  IV U141 ( .A(B[53]), .Z(n310) );
  IV U142 ( .A(B[54]), .Z(n311) );
  IV U143 ( .A(B[55]), .Z(n312) );
  IV U144 ( .A(B[56]), .Z(n313) );
  IV U145 ( .A(B[57]), .Z(n314) );
  IV U146 ( .A(B[58]), .Z(n315) );
  IV U147 ( .A(B[238]), .Z(n495) );
  IV U148 ( .A(B[59]), .Z(n316) );
  IV U149 ( .A(B[60]), .Z(n317) );
  IV U150 ( .A(B[61]), .Z(n318) );
  IV U151 ( .A(B[62]), .Z(n319) );
  IV U152 ( .A(B[63]), .Z(n320) );
  IV U153 ( .A(B[64]), .Z(n321) );
  IV U154 ( .A(B[65]), .Z(n322) );
  IV U155 ( .A(B[66]), .Z(n323) );
  IV U156 ( .A(B[67]), .Z(n324) );
  IV U157 ( .A(B[68]), .Z(n325) );
  IV U158 ( .A(B[239]), .Z(n496) );
  IV U159 ( .A(B[69]), .Z(n326) );
  IV U160 ( .A(B[70]), .Z(n327) );
  IV U161 ( .A(B[71]), .Z(n328) );
  IV U162 ( .A(B[72]), .Z(n329) );
  IV U163 ( .A(B[73]), .Z(n330) );
  IV U164 ( .A(B[74]), .Z(n331) );
  IV U165 ( .A(B[75]), .Z(n332) );
  IV U166 ( .A(B[76]), .Z(n333) );
  IV U167 ( .A(B[77]), .Z(n334) );
  IV U168 ( .A(B[78]), .Z(n335) );
  IV U169 ( .A(B[240]), .Z(n497) );
  IV U170 ( .A(B[79]), .Z(n336) );
  IV U171 ( .A(B[80]), .Z(n337) );
  IV U172 ( .A(B[81]), .Z(n338) );
  IV U173 ( .A(B[82]), .Z(n339) );
  IV U174 ( .A(B[83]), .Z(n340) );
  IV U175 ( .A(B[84]), .Z(n341) );
  IV U176 ( .A(B[85]), .Z(n342) );
  IV U177 ( .A(B[86]), .Z(n343) );
  IV U178 ( .A(B[87]), .Z(n344) );
  IV U179 ( .A(B[88]), .Z(n345) );
  IV U180 ( .A(B[241]), .Z(n498) );
  IV U181 ( .A(B[89]), .Z(n346) );
  IV U182 ( .A(B[90]), .Z(n347) );
  IV U183 ( .A(B[91]), .Z(n348) );
  IV U184 ( .A(B[92]), .Z(n349) );
  IV U185 ( .A(B[93]), .Z(n350) );
  IV U186 ( .A(B[94]), .Z(n351) );
  IV U187 ( .A(B[95]), .Z(n352) );
  IV U188 ( .A(B[96]), .Z(n353) );
  IV U189 ( .A(B[97]), .Z(n354) );
  IV U190 ( .A(B[98]), .Z(n355) );
  IV U191 ( .A(B[242]), .Z(n499) );
  IV U192 ( .A(B[99]), .Z(n356) );
  IV U193 ( .A(B[100]), .Z(n357) );
  IV U194 ( .A(B[101]), .Z(n358) );
  IV U195 ( .A(B[102]), .Z(n359) );
  IV U196 ( .A(B[103]), .Z(n360) );
  IV U197 ( .A(B[104]), .Z(n361) );
  IV U198 ( .A(B[105]), .Z(n362) );
  IV U199 ( .A(B[106]), .Z(n363) );
  IV U200 ( .A(B[107]), .Z(n364) );
  IV U201 ( .A(B[108]), .Z(n365) );
  IV U202 ( .A(B[243]), .Z(n500) );
  IV U203 ( .A(B[109]), .Z(n366) );
  IV U204 ( .A(B[110]), .Z(n367) );
  IV U205 ( .A(B[111]), .Z(n368) );
  IV U206 ( .A(B[112]), .Z(n369) );
  IV U207 ( .A(B[113]), .Z(n370) );
  IV U208 ( .A(B[114]), .Z(n371) );
  IV U209 ( .A(B[115]), .Z(n372) );
  IV U210 ( .A(B[116]), .Z(n373) );
  IV U211 ( .A(B[117]), .Z(n374) );
  IV U212 ( .A(B[118]), .Z(n375) );
  IV U213 ( .A(B[244]), .Z(n501) );
  IV U214 ( .A(B[119]), .Z(n376) );
  IV U215 ( .A(B[120]), .Z(n377) );
  IV U216 ( .A(B[121]), .Z(n378) );
  IV U217 ( .A(B[122]), .Z(n379) );
  IV U218 ( .A(B[123]), .Z(n380) );
  IV U219 ( .A(B[124]), .Z(n381) );
  IV U220 ( .A(B[125]), .Z(n382) );
  IV U221 ( .A(B[126]), .Z(n383) );
  IV U222 ( .A(B[127]), .Z(n384) );
  IV U223 ( .A(B[128]), .Z(n385) );
  IV U224 ( .A(B[245]), .Z(n502) );
  IV U225 ( .A(B[129]), .Z(n386) );
  IV U226 ( .A(B[130]), .Z(n387) );
  IV U227 ( .A(B[131]), .Z(n388) );
  IV U228 ( .A(B[132]), .Z(n389) );
  IV U229 ( .A(B[133]), .Z(n390) );
  IV U230 ( .A(B[134]), .Z(n391) );
  IV U231 ( .A(B[135]), .Z(n392) );
  IV U232 ( .A(B[136]), .Z(n393) );
  IV U233 ( .A(B[137]), .Z(n394) );
  IV U234 ( .A(B[138]), .Z(n395) );
  IV U235 ( .A(B[246]), .Z(n503) );
  IV U236 ( .A(B[139]), .Z(n396) );
  IV U237 ( .A(B[140]), .Z(n397) );
  IV U238 ( .A(B[141]), .Z(n398) );
  IV U239 ( .A(B[142]), .Z(n399) );
  IV U240 ( .A(B[143]), .Z(n400) );
  IV U241 ( .A(B[144]), .Z(n401) );
  IV U242 ( .A(B[145]), .Z(n402) );
  IV U243 ( .A(B[146]), .Z(n403) );
  IV U244 ( .A(B[147]), .Z(n404) );
  IV U245 ( .A(B[148]), .Z(n405) );
  IV U246 ( .A(B[247]), .Z(n504) );
  IV U247 ( .A(B[149]), .Z(n406) );
  IV U248 ( .A(B[150]), .Z(n407) );
  IV U249 ( .A(B[151]), .Z(n408) );
  IV U250 ( .A(B[152]), .Z(n409) );
  IV U251 ( .A(B[153]), .Z(n410) );
  IV U252 ( .A(B[154]), .Z(n411) );
  IV U253 ( .A(B[155]), .Z(n412) );
  IV U254 ( .A(B[156]), .Z(n413) );
  IV U255 ( .A(B[157]), .Z(n414) );
  IV U256 ( .A(B[158]), .Z(n415) );
  IV U257 ( .A(B[248]), .Z(n505) );
endmodule


module FA_1806 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XNOR U1 ( .A(CI), .B(A), .Z(S) );
endmodule


module FA_1807 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  NANDN U1 ( .A(CI), .B(S), .Z(CO) );
  XNOR U2 ( .A(A), .B(CI), .Z(S) );
endmodule


module FA_1808 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1809 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1810 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1811 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1812 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1813 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1814 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1815 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1816 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1817 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1818 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1819 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1820 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1821 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1822 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1823 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1824 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1825 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1826 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1827 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1828 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1829 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1830 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1831 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1832 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1833 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1834 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1835 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1836 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1837 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1838 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1839 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1840 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1841 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1842 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1843 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1844 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1845 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1846 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1847 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1848 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1849 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1850 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1851 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1852 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1853 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1854 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1855 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1856 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1857 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1858 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1859 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1860 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1861 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1862 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1863 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1864 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1865 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1866 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1867 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1868 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1869 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1870 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1871 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1872 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1873 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1874 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1875 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1876 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1877 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1878 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1879 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1880 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1881 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1882 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1883 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1884 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1885 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1886 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1887 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1888 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1889 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1890 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1891 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1892 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1893 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1894 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1895 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1896 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1897 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1898 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1899 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1900 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1901 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1902 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1903 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1904 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1905 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1906 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1907 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1908 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1909 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1910 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1911 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1912 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1913 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1914 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1915 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1916 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1917 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1918 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1919 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1920 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1921 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1922 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1923 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1924 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1925 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1926 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1927 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1928 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1929 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1930 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1931 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1932 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1933 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1934 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1935 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1936 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1937 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1938 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1939 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1940 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1941 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1942 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1943 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1944 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1945 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1946 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1947 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1948 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1949 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1950 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1951 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1952 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1953 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1954 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1955 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1956 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1957 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1958 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1959 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1960 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1961 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1962 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1963 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1964 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1965 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1966 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1967 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1968 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1969 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1970 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1971 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1972 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1973 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1974 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1975 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1976 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1977 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1978 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1979 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1980 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1981 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1982 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1983 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1984 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1985 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1986 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1987 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1988 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1989 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1990 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1991 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1992 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1993 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1994 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1995 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1996 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1997 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1998 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1999 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2000 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2001 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2002 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2003 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2004 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2005 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2006 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2007 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2008 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2009 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2010 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2011 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2012 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2013 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2014 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2015 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2016 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2017 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2018 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2019 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2020 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2021 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2022 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2023 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2024 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2025 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2026 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2027 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2028 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2029 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2030 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2031 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2032 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2033 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2034 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2035 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2036 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2037 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2038 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2039 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2040 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2041 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2042 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2043 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2044 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2045 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2046 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2047 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2048 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2049 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2050 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2051 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2052 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2053 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2054 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2055 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2056 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2057 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2058 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2059 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2060 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2061 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2062 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_2063 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XNOR U1 ( .A(B), .B(A), .Z(S) );
  OR U2 ( .A(B), .B(A), .Z(CO) );
endmodule


module SUB_N258_4 ( A, B, S, CO );
  input [257:0] A;
  input [257:0] B;
  output [257:0] S;
  output CO;
  wire   n2, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512;
  wire   [257:1] C;

  FA_2063 \FAINST[0].FA_  ( .A(A[0]), .B(n2), .CI(1'b1), .S(S[0]), .CO(C[1])
         );
  FA_2062 \FAINST[1].FA_  ( .A(A[1]), .B(n258), .CI(C[1]), .S(S[1]), .CO(C[2])
         );
  FA_2061 \FAINST[2].FA_  ( .A(A[2]), .B(n259), .CI(C[2]), .S(S[2]), .CO(C[3])
         );
  FA_2060 \FAINST[3].FA_  ( .A(A[3]), .B(n260), .CI(C[3]), .S(S[3]), .CO(C[4])
         );
  FA_2059 \FAINST[4].FA_  ( .A(A[4]), .B(n261), .CI(C[4]), .S(S[4]), .CO(C[5])
         );
  FA_2058 \FAINST[5].FA_  ( .A(A[5]), .B(n262), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_2057 \FAINST[6].FA_  ( .A(A[6]), .B(n263), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_2056 \FAINST[7].FA_  ( .A(A[7]), .B(n264), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_2055 \FAINST[8].FA_  ( .A(A[8]), .B(n265), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_2054 \FAINST[9].FA_  ( .A(A[9]), .B(n266), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_2053 \FAINST[10].FA_  ( .A(A[10]), .B(n267), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_2052 \FAINST[11].FA_  ( .A(A[11]), .B(n268), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_2051 \FAINST[12].FA_  ( .A(A[12]), .B(n269), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_2050 \FAINST[13].FA_  ( .A(A[13]), .B(n270), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_2049 \FAINST[14].FA_  ( .A(A[14]), .B(n271), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_2048 \FAINST[15].FA_  ( .A(A[15]), .B(n272), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_2047 \FAINST[16].FA_  ( .A(A[16]), .B(n273), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_2046 \FAINST[17].FA_  ( .A(A[17]), .B(n274), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_2045 \FAINST[18].FA_  ( .A(A[18]), .B(n275), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_2044 \FAINST[19].FA_  ( .A(A[19]), .B(n276), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_2043 \FAINST[20].FA_  ( .A(A[20]), .B(n277), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_2042 \FAINST[21].FA_  ( .A(A[21]), .B(n278), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_2041 \FAINST[22].FA_  ( .A(A[22]), .B(n279), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_2040 \FAINST[23].FA_  ( .A(A[23]), .B(n280), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_2039 \FAINST[24].FA_  ( .A(A[24]), .B(n281), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_2038 \FAINST[25].FA_  ( .A(A[25]), .B(n282), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_2037 \FAINST[26].FA_  ( .A(A[26]), .B(n283), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_2036 \FAINST[27].FA_  ( .A(A[27]), .B(n284), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_2035 \FAINST[28].FA_  ( .A(A[28]), .B(n285), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_2034 \FAINST[29].FA_  ( .A(A[29]), .B(n286), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_2033 \FAINST[30].FA_  ( .A(A[30]), .B(n287), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_2032 \FAINST[31].FA_  ( .A(A[31]), .B(n288), .CI(C[31]), .S(S[31]), .CO(
        C[32]) );
  FA_2031 \FAINST[32].FA_  ( .A(A[32]), .B(n289), .CI(C[32]), .S(S[32]), .CO(
        C[33]) );
  FA_2030 \FAINST[33].FA_  ( .A(A[33]), .B(n290), .CI(C[33]), .S(S[33]), .CO(
        C[34]) );
  FA_2029 \FAINST[34].FA_  ( .A(A[34]), .B(n291), .CI(C[34]), .S(S[34]), .CO(
        C[35]) );
  FA_2028 \FAINST[35].FA_  ( .A(A[35]), .B(n292), .CI(C[35]), .S(S[35]), .CO(
        C[36]) );
  FA_2027 \FAINST[36].FA_  ( .A(A[36]), .B(n293), .CI(C[36]), .S(S[36]), .CO(
        C[37]) );
  FA_2026 \FAINST[37].FA_  ( .A(A[37]), .B(n294), .CI(C[37]), .S(S[37]), .CO(
        C[38]) );
  FA_2025 \FAINST[38].FA_  ( .A(A[38]), .B(n295), .CI(C[38]), .S(S[38]), .CO(
        C[39]) );
  FA_2024 \FAINST[39].FA_  ( .A(A[39]), .B(n296), .CI(C[39]), .S(S[39]), .CO(
        C[40]) );
  FA_2023 \FAINST[40].FA_  ( .A(A[40]), .B(n297), .CI(C[40]), .S(S[40]), .CO(
        C[41]) );
  FA_2022 \FAINST[41].FA_  ( .A(A[41]), .B(n298), .CI(C[41]), .S(S[41]), .CO(
        C[42]) );
  FA_2021 \FAINST[42].FA_  ( .A(A[42]), .B(n299), .CI(C[42]), .S(S[42]), .CO(
        C[43]) );
  FA_2020 \FAINST[43].FA_  ( .A(A[43]), .B(n300), .CI(C[43]), .S(S[43]), .CO(
        C[44]) );
  FA_2019 \FAINST[44].FA_  ( .A(A[44]), .B(n301), .CI(C[44]), .S(S[44]), .CO(
        C[45]) );
  FA_2018 \FAINST[45].FA_  ( .A(A[45]), .B(n302), .CI(C[45]), .S(S[45]), .CO(
        C[46]) );
  FA_2017 \FAINST[46].FA_  ( .A(A[46]), .B(n303), .CI(C[46]), .S(S[46]), .CO(
        C[47]) );
  FA_2016 \FAINST[47].FA_  ( .A(A[47]), .B(n304), .CI(C[47]), .S(S[47]), .CO(
        C[48]) );
  FA_2015 \FAINST[48].FA_  ( .A(A[48]), .B(n305), .CI(C[48]), .S(S[48]), .CO(
        C[49]) );
  FA_2014 \FAINST[49].FA_  ( .A(A[49]), .B(n306), .CI(C[49]), .S(S[49]), .CO(
        C[50]) );
  FA_2013 \FAINST[50].FA_  ( .A(A[50]), .B(n307), .CI(C[50]), .S(S[50]), .CO(
        C[51]) );
  FA_2012 \FAINST[51].FA_  ( .A(A[51]), .B(n308), .CI(C[51]), .S(S[51]), .CO(
        C[52]) );
  FA_2011 \FAINST[52].FA_  ( .A(A[52]), .B(n309), .CI(C[52]), .S(S[52]), .CO(
        C[53]) );
  FA_2010 \FAINST[53].FA_  ( .A(A[53]), .B(n310), .CI(C[53]), .S(S[53]), .CO(
        C[54]) );
  FA_2009 \FAINST[54].FA_  ( .A(A[54]), .B(n311), .CI(C[54]), .S(S[54]), .CO(
        C[55]) );
  FA_2008 \FAINST[55].FA_  ( .A(A[55]), .B(n312), .CI(C[55]), .S(S[55]), .CO(
        C[56]) );
  FA_2007 \FAINST[56].FA_  ( .A(A[56]), .B(n313), .CI(C[56]), .S(S[56]), .CO(
        C[57]) );
  FA_2006 \FAINST[57].FA_  ( .A(A[57]), .B(n314), .CI(C[57]), .S(S[57]), .CO(
        C[58]) );
  FA_2005 \FAINST[58].FA_  ( .A(A[58]), .B(n315), .CI(C[58]), .S(S[58]), .CO(
        C[59]) );
  FA_2004 \FAINST[59].FA_  ( .A(A[59]), .B(n316), .CI(C[59]), .S(S[59]), .CO(
        C[60]) );
  FA_2003 \FAINST[60].FA_  ( .A(A[60]), .B(n317), .CI(C[60]), .S(S[60]), .CO(
        C[61]) );
  FA_2002 \FAINST[61].FA_  ( .A(A[61]), .B(n318), .CI(C[61]), .S(S[61]), .CO(
        C[62]) );
  FA_2001 \FAINST[62].FA_  ( .A(A[62]), .B(n319), .CI(C[62]), .S(S[62]), .CO(
        C[63]) );
  FA_2000 \FAINST[63].FA_  ( .A(A[63]), .B(n320), .CI(C[63]), .S(S[63]), .CO(
        C[64]) );
  FA_1999 \FAINST[64].FA_  ( .A(A[64]), .B(n321), .CI(C[64]), .S(S[64]), .CO(
        C[65]) );
  FA_1998 \FAINST[65].FA_  ( .A(A[65]), .B(n322), .CI(C[65]), .S(S[65]), .CO(
        C[66]) );
  FA_1997 \FAINST[66].FA_  ( .A(A[66]), .B(n323), .CI(C[66]), .S(S[66]), .CO(
        C[67]) );
  FA_1996 \FAINST[67].FA_  ( .A(A[67]), .B(n324), .CI(C[67]), .S(S[67]), .CO(
        C[68]) );
  FA_1995 \FAINST[68].FA_  ( .A(A[68]), .B(n325), .CI(C[68]), .S(S[68]), .CO(
        C[69]) );
  FA_1994 \FAINST[69].FA_  ( .A(A[69]), .B(n326), .CI(C[69]), .S(S[69]), .CO(
        C[70]) );
  FA_1993 \FAINST[70].FA_  ( .A(A[70]), .B(n327), .CI(C[70]), .S(S[70]), .CO(
        C[71]) );
  FA_1992 \FAINST[71].FA_  ( .A(A[71]), .B(n328), .CI(C[71]), .S(S[71]), .CO(
        C[72]) );
  FA_1991 \FAINST[72].FA_  ( .A(A[72]), .B(n329), .CI(C[72]), .S(S[72]), .CO(
        C[73]) );
  FA_1990 \FAINST[73].FA_  ( .A(A[73]), .B(n330), .CI(C[73]), .S(S[73]), .CO(
        C[74]) );
  FA_1989 \FAINST[74].FA_  ( .A(A[74]), .B(n331), .CI(C[74]), .S(S[74]), .CO(
        C[75]) );
  FA_1988 \FAINST[75].FA_  ( .A(A[75]), .B(n332), .CI(C[75]), .S(S[75]), .CO(
        C[76]) );
  FA_1987 \FAINST[76].FA_  ( .A(A[76]), .B(n333), .CI(C[76]), .S(S[76]), .CO(
        C[77]) );
  FA_1986 \FAINST[77].FA_  ( .A(A[77]), .B(n334), .CI(C[77]), .S(S[77]), .CO(
        C[78]) );
  FA_1985 \FAINST[78].FA_  ( .A(A[78]), .B(n335), .CI(C[78]), .S(S[78]), .CO(
        C[79]) );
  FA_1984 \FAINST[79].FA_  ( .A(A[79]), .B(n336), .CI(C[79]), .S(S[79]), .CO(
        C[80]) );
  FA_1983 \FAINST[80].FA_  ( .A(A[80]), .B(n337), .CI(C[80]), .S(S[80]), .CO(
        C[81]) );
  FA_1982 \FAINST[81].FA_  ( .A(A[81]), .B(n338), .CI(C[81]), .S(S[81]), .CO(
        C[82]) );
  FA_1981 \FAINST[82].FA_  ( .A(A[82]), .B(n339), .CI(C[82]), .S(S[82]), .CO(
        C[83]) );
  FA_1980 \FAINST[83].FA_  ( .A(A[83]), .B(n340), .CI(C[83]), .S(S[83]), .CO(
        C[84]) );
  FA_1979 \FAINST[84].FA_  ( .A(A[84]), .B(n341), .CI(C[84]), .S(S[84]), .CO(
        C[85]) );
  FA_1978 \FAINST[85].FA_  ( .A(A[85]), .B(n342), .CI(C[85]), .S(S[85]), .CO(
        C[86]) );
  FA_1977 \FAINST[86].FA_  ( .A(A[86]), .B(n343), .CI(C[86]), .S(S[86]), .CO(
        C[87]) );
  FA_1976 \FAINST[87].FA_  ( .A(A[87]), .B(n344), .CI(C[87]), .S(S[87]), .CO(
        C[88]) );
  FA_1975 \FAINST[88].FA_  ( .A(A[88]), .B(n345), .CI(C[88]), .S(S[88]), .CO(
        C[89]) );
  FA_1974 \FAINST[89].FA_  ( .A(A[89]), .B(n346), .CI(C[89]), .S(S[89]), .CO(
        C[90]) );
  FA_1973 \FAINST[90].FA_  ( .A(A[90]), .B(n347), .CI(C[90]), .S(S[90]), .CO(
        C[91]) );
  FA_1972 \FAINST[91].FA_  ( .A(A[91]), .B(n348), .CI(C[91]), .S(S[91]), .CO(
        C[92]) );
  FA_1971 \FAINST[92].FA_  ( .A(A[92]), .B(n349), .CI(C[92]), .S(S[92]), .CO(
        C[93]) );
  FA_1970 \FAINST[93].FA_  ( .A(A[93]), .B(n350), .CI(C[93]), .S(S[93]), .CO(
        C[94]) );
  FA_1969 \FAINST[94].FA_  ( .A(A[94]), .B(n351), .CI(C[94]), .S(S[94]), .CO(
        C[95]) );
  FA_1968 \FAINST[95].FA_  ( .A(A[95]), .B(n352), .CI(C[95]), .S(S[95]), .CO(
        C[96]) );
  FA_1967 \FAINST[96].FA_  ( .A(A[96]), .B(n353), .CI(C[96]), .S(S[96]), .CO(
        C[97]) );
  FA_1966 \FAINST[97].FA_  ( .A(A[97]), .B(n354), .CI(C[97]), .S(S[97]), .CO(
        C[98]) );
  FA_1965 \FAINST[98].FA_  ( .A(A[98]), .B(n355), .CI(C[98]), .S(S[98]), .CO(
        C[99]) );
  FA_1964 \FAINST[99].FA_  ( .A(A[99]), .B(n356), .CI(C[99]), .S(S[99]), .CO(
        C[100]) );
  FA_1963 \FAINST[100].FA_  ( .A(A[100]), .B(n357), .CI(C[100]), .S(S[100]), 
        .CO(C[101]) );
  FA_1962 \FAINST[101].FA_  ( .A(A[101]), .B(n358), .CI(C[101]), .S(S[101]), 
        .CO(C[102]) );
  FA_1961 \FAINST[102].FA_  ( .A(A[102]), .B(n359), .CI(C[102]), .S(S[102]), 
        .CO(C[103]) );
  FA_1960 \FAINST[103].FA_  ( .A(A[103]), .B(n360), .CI(C[103]), .S(S[103]), 
        .CO(C[104]) );
  FA_1959 \FAINST[104].FA_  ( .A(A[104]), .B(n361), .CI(C[104]), .S(S[104]), 
        .CO(C[105]) );
  FA_1958 \FAINST[105].FA_  ( .A(A[105]), .B(n362), .CI(C[105]), .S(S[105]), 
        .CO(C[106]) );
  FA_1957 \FAINST[106].FA_  ( .A(A[106]), .B(n363), .CI(C[106]), .S(S[106]), 
        .CO(C[107]) );
  FA_1956 \FAINST[107].FA_  ( .A(A[107]), .B(n364), .CI(C[107]), .S(S[107]), 
        .CO(C[108]) );
  FA_1955 \FAINST[108].FA_  ( .A(A[108]), .B(n365), .CI(C[108]), .S(S[108]), 
        .CO(C[109]) );
  FA_1954 \FAINST[109].FA_  ( .A(A[109]), .B(n366), .CI(C[109]), .S(S[109]), 
        .CO(C[110]) );
  FA_1953 \FAINST[110].FA_  ( .A(A[110]), .B(n367), .CI(C[110]), .S(S[110]), 
        .CO(C[111]) );
  FA_1952 \FAINST[111].FA_  ( .A(A[111]), .B(n368), .CI(C[111]), .S(S[111]), 
        .CO(C[112]) );
  FA_1951 \FAINST[112].FA_  ( .A(A[112]), .B(n369), .CI(C[112]), .S(S[112]), 
        .CO(C[113]) );
  FA_1950 \FAINST[113].FA_  ( .A(A[113]), .B(n370), .CI(C[113]), .S(S[113]), 
        .CO(C[114]) );
  FA_1949 \FAINST[114].FA_  ( .A(A[114]), .B(n371), .CI(C[114]), .S(S[114]), 
        .CO(C[115]) );
  FA_1948 \FAINST[115].FA_  ( .A(A[115]), .B(n372), .CI(C[115]), .S(S[115]), 
        .CO(C[116]) );
  FA_1947 \FAINST[116].FA_  ( .A(A[116]), .B(n373), .CI(C[116]), .S(S[116]), 
        .CO(C[117]) );
  FA_1946 \FAINST[117].FA_  ( .A(A[117]), .B(n374), .CI(C[117]), .S(S[117]), 
        .CO(C[118]) );
  FA_1945 \FAINST[118].FA_  ( .A(A[118]), .B(n375), .CI(C[118]), .S(S[118]), 
        .CO(C[119]) );
  FA_1944 \FAINST[119].FA_  ( .A(A[119]), .B(n376), .CI(C[119]), .S(S[119]), 
        .CO(C[120]) );
  FA_1943 \FAINST[120].FA_  ( .A(A[120]), .B(n377), .CI(C[120]), .S(S[120]), 
        .CO(C[121]) );
  FA_1942 \FAINST[121].FA_  ( .A(A[121]), .B(n378), .CI(C[121]), .S(S[121]), 
        .CO(C[122]) );
  FA_1941 \FAINST[122].FA_  ( .A(A[122]), .B(n379), .CI(C[122]), .S(S[122]), 
        .CO(C[123]) );
  FA_1940 \FAINST[123].FA_  ( .A(A[123]), .B(n380), .CI(C[123]), .S(S[123]), 
        .CO(C[124]) );
  FA_1939 \FAINST[124].FA_  ( .A(A[124]), .B(n381), .CI(C[124]), .S(S[124]), 
        .CO(C[125]) );
  FA_1938 \FAINST[125].FA_  ( .A(A[125]), .B(n382), .CI(C[125]), .S(S[125]), 
        .CO(C[126]) );
  FA_1937 \FAINST[126].FA_  ( .A(A[126]), .B(n383), .CI(C[126]), .S(S[126]), 
        .CO(C[127]) );
  FA_1936 \FAINST[127].FA_  ( .A(A[127]), .B(n384), .CI(C[127]), .S(S[127]), 
        .CO(C[128]) );
  FA_1935 \FAINST[128].FA_  ( .A(A[128]), .B(n385), .CI(C[128]), .S(S[128]), 
        .CO(C[129]) );
  FA_1934 \FAINST[129].FA_  ( .A(A[129]), .B(n386), .CI(C[129]), .S(S[129]), 
        .CO(C[130]) );
  FA_1933 \FAINST[130].FA_  ( .A(A[130]), .B(n387), .CI(C[130]), .S(S[130]), 
        .CO(C[131]) );
  FA_1932 \FAINST[131].FA_  ( .A(A[131]), .B(n388), .CI(C[131]), .S(S[131]), 
        .CO(C[132]) );
  FA_1931 \FAINST[132].FA_  ( .A(A[132]), .B(n389), .CI(C[132]), .S(S[132]), 
        .CO(C[133]) );
  FA_1930 \FAINST[133].FA_  ( .A(A[133]), .B(n390), .CI(C[133]), .S(S[133]), 
        .CO(C[134]) );
  FA_1929 \FAINST[134].FA_  ( .A(A[134]), .B(n391), .CI(C[134]), .S(S[134]), 
        .CO(C[135]) );
  FA_1928 \FAINST[135].FA_  ( .A(A[135]), .B(n392), .CI(C[135]), .S(S[135]), 
        .CO(C[136]) );
  FA_1927 \FAINST[136].FA_  ( .A(A[136]), .B(n393), .CI(C[136]), .S(S[136]), 
        .CO(C[137]) );
  FA_1926 \FAINST[137].FA_  ( .A(A[137]), .B(n394), .CI(C[137]), .S(S[137]), 
        .CO(C[138]) );
  FA_1925 \FAINST[138].FA_  ( .A(A[138]), .B(n395), .CI(C[138]), .S(S[138]), 
        .CO(C[139]) );
  FA_1924 \FAINST[139].FA_  ( .A(A[139]), .B(n396), .CI(C[139]), .S(S[139]), 
        .CO(C[140]) );
  FA_1923 \FAINST[140].FA_  ( .A(A[140]), .B(n397), .CI(C[140]), .S(S[140]), 
        .CO(C[141]) );
  FA_1922 \FAINST[141].FA_  ( .A(A[141]), .B(n398), .CI(C[141]), .S(S[141]), 
        .CO(C[142]) );
  FA_1921 \FAINST[142].FA_  ( .A(A[142]), .B(n399), .CI(C[142]), .S(S[142]), 
        .CO(C[143]) );
  FA_1920 \FAINST[143].FA_  ( .A(A[143]), .B(n400), .CI(C[143]), .S(S[143]), 
        .CO(C[144]) );
  FA_1919 \FAINST[144].FA_  ( .A(A[144]), .B(n401), .CI(C[144]), .S(S[144]), 
        .CO(C[145]) );
  FA_1918 \FAINST[145].FA_  ( .A(A[145]), .B(n402), .CI(C[145]), .S(S[145]), 
        .CO(C[146]) );
  FA_1917 \FAINST[146].FA_  ( .A(A[146]), .B(n403), .CI(C[146]), .S(S[146]), 
        .CO(C[147]) );
  FA_1916 \FAINST[147].FA_  ( .A(A[147]), .B(n404), .CI(C[147]), .S(S[147]), 
        .CO(C[148]) );
  FA_1915 \FAINST[148].FA_  ( .A(A[148]), .B(n405), .CI(C[148]), .S(S[148]), 
        .CO(C[149]) );
  FA_1914 \FAINST[149].FA_  ( .A(A[149]), .B(n406), .CI(C[149]), .S(S[149]), 
        .CO(C[150]) );
  FA_1913 \FAINST[150].FA_  ( .A(A[150]), .B(n407), .CI(C[150]), .S(S[150]), 
        .CO(C[151]) );
  FA_1912 \FAINST[151].FA_  ( .A(A[151]), .B(n408), .CI(C[151]), .S(S[151]), 
        .CO(C[152]) );
  FA_1911 \FAINST[152].FA_  ( .A(A[152]), .B(n409), .CI(C[152]), .S(S[152]), 
        .CO(C[153]) );
  FA_1910 \FAINST[153].FA_  ( .A(A[153]), .B(n410), .CI(C[153]), .S(S[153]), 
        .CO(C[154]) );
  FA_1909 \FAINST[154].FA_  ( .A(A[154]), .B(n411), .CI(C[154]), .S(S[154]), 
        .CO(C[155]) );
  FA_1908 \FAINST[155].FA_  ( .A(A[155]), .B(n412), .CI(C[155]), .S(S[155]), 
        .CO(C[156]) );
  FA_1907 \FAINST[156].FA_  ( .A(A[156]), .B(n413), .CI(C[156]), .S(S[156]), 
        .CO(C[157]) );
  FA_1906 \FAINST[157].FA_  ( .A(A[157]), .B(n414), .CI(C[157]), .S(S[157]), 
        .CO(C[158]) );
  FA_1905 \FAINST[158].FA_  ( .A(A[158]), .B(n415), .CI(C[158]), .S(S[158]), 
        .CO(C[159]) );
  FA_1904 \FAINST[159].FA_  ( .A(A[159]), .B(n416), .CI(C[159]), .S(S[159]), 
        .CO(C[160]) );
  FA_1903 \FAINST[160].FA_  ( .A(A[160]), .B(n417), .CI(C[160]), .S(S[160]), 
        .CO(C[161]) );
  FA_1902 \FAINST[161].FA_  ( .A(A[161]), .B(n418), .CI(C[161]), .S(S[161]), 
        .CO(C[162]) );
  FA_1901 \FAINST[162].FA_  ( .A(A[162]), .B(n419), .CI(C[162]), .S(S[162]), 
        .CO(C[163]) );
  FA_1900 \FAINST[163].FA_  ( .A(A[163]), .B(n420), .CI(C[163]), .S(S[163]), 
        .CO(C[164]) );
  FA_1899 \FAINST[164].FA_  ( .A(A[164]), .B(n421), .CI(C[164]), .S(S[164]), 
        .CO(C[165]) );
  FA_1898 \FAINST[165].FA_  ( .A(A[165]), .B(n422), .CI(C[165]), .S(S[165]), 
        .CO(C[166]) );
  FA_1897 \FAINST[166].FA_  ( .A(A[166]), .B(n423), .CI(C[166]), .S(S[166]), 
        .CO(C[167]) );
  FA_1896 \FAINST[167].FA_  ( .A(A[167]), .B(n424), .CI(C[167]), .S(S[167]), 
        .CO(C[168]) );
  FA_1895 \FAINST[168].FA_  ( .A(A[168]), .B(n425), .CI(C[168]), .S(S[168]), 
        .CO(C[169]) );
  FA_1894 \FAINST[169].FA_  ( .A(A[169]), .B(n426), .CI(C[169]), .S(S[169]), 
        .CO(C[170]) );
  FA_1893 \FAINST[170].FA_  ( .A(A[170]), .B(n427), .CI(C[170]), .S(S[170]), 
        .CO(C[171]) );
  FA_1892 \FAINST[171].FA_  ( .A(A[171]), .B(n428), .CI(C[171]), .S(S[171]), 
        .CO(C[172]) );
  FA_1891 \FAINST[172].FA_  ( .A(A[172]), .B(n429), .CI(C[172]), .S(S[172]), 
        .CO(C[173]) );
  FA_1890 \FAINST[173].FA_  ( .A(A[173]), .B(n430), .CI(C[173]), .S(S[173]), 
        .CO(C[174]) );
  FA_1889 \FAINST[174].FA_  ( .A(A[174]), .B(n431), .CI(C[174]), .S(S[174]), 
        .CO(C[175]) );
  FA_1888 \FAINST[175].FA_  ( .A(A[175]), .B(n432), .CI(C[175]), .S(S[175]), 
        .CO(C[176]) );
  FA_1887 \FAINST[176].FA_  ( .A(A[176]), .B(n433), .CI(C[176]), .S(S[176]), 
        .CO(C[177]) );
  FA_1886 \FAINST[177].FA_  ( .A(A[177]), .B(n434), .CI(C[177]), .S(S[177]), 
        .CO(C[178]) );
  FA_1885 \FAINST[178].FA_  ( .A(A[178]), .B(n435), .CI(C[178]), .S(S[178]), 
        .CO(C[179]) );
  FA_1884 \FAINST[179].FA_  ( .A(A[179]), .B(n436), .CI(C[179]), .S(S[179]), 
        .CO(C[180]) );
  FA_1883 \FAINST[180].FA_  ( .A(A[180]), .B(n437), .CI(C[180]), .S(S[180]), 
        .CO(C[181]) );
  FA_1882 \FAINST[181].FA_  ( .A(A[181]), .B(n438), .CI(C[181]), .S(S[181]), 
        .CO(C[182]) );
  FA_1881 \FAINST[182].FA_  ( .A(A[182]), .B(n439), .CI(C[182]), .S(S[182]), 
        .CO(C[183]) );
  FA_1880 \FAINST[183].FA_  ( .A(A[183]), .B(n440), .CI(C[183]), .S(S[183]), 
        .CO(C[184]) );
  FA_1879 \FAINST[184].FA_  ( .A(A[184]), .B(n441), .CI(C[184]), .S(S[184]), 
        .CO(C[185]) );
  FA_1878 \FAINST[185].FA_  ( .A(A[185]), .B(n442), .CI(C[185]), .S(S[185]), 
        .CO(C[186]) );
  FA_1877 \FAINST[186].FA_  ( .A(A[186]), .B(n443), .CI(C[186]), .S(S[186]), 
        .CO(C[187]) );
  FA_1876 \FAINST[187].FA_  ( .A(A[187]), .B(n444), .CI(C[187]), .S(S[187]), 
        .CO(C[188]) );
  FA_1875 \FAINST[188].FA_  ( .A(A[188]), .B(n445), .CI(C[188]), .S(S[188]), 
        .CO(C[189]) );
  FA_1874 \FAINST[189].FA_  ( .A(A[189]), .B(n446), .CI(C[189]), .S(S[189]), 
        .CO(C[190]) );
  FA_1873 \FAINST[190].FA_  ( .A(A[190]), .B(n447), .CI(C[190]), .S(S[190]), 
        .CO(C[191]) );
  FA_1872 \FAINST[191].FA_  ( .A(A[191]), .B(n448), .CI(C[191]), .S(S[191]), 
        .CO(C[192]) );
  FA_1871 \FAINST[192].FA_  ( .A(A[192]), .B(n449), .CI(C[192]), .S(S[192]), 
        .CO(C[193]) );
  FA_1870 \FAINST[193].FA_  ( .A(A[193]), .B(n450), .CI(C[193]), .S(S[193]), 
        .CO(C[194]) );
  FA_1869 \FAINST[194].FA_  ( .A(A[194]), .B(n451), .CI(C[194]), .S(S[194]), 
        .CO(C[195]) );
  FA_1868 \FAINST[195].FA_  ( .A(A[195]), .B(n452), .CI(C[195]), .S(S[195]), 
        .CO(C[196]) );
  FA_1867 \FAINST[196].FA_  ( .A(A[196]), .B(n453), .CI(C[196]), .S(S[196]), 
        .CO(C[197]) );
  FA_1866 \FAINST[197].FA_  ( .A(A[197]), .B(n454), .CI(C[197]), .S(S[197]), 
        .CO(C[198]) );
  FA_1865 \FAINST[198].FA_  ( .A(A[198]), .B(n455), .CI(C[198]), .S(S[198]), 
        .CO(C[199]) );
  FA_1864 \FAINST[199].FA_  ( .A(A[199]), .B(n456), .CI(C[199]), .S(S[199]), 
        .CO(C[200]) );
  FA_1863 \FAINST[200].FA_  ( .A(A[200]), .B(n457), .CI(C[200]), .S(S[200]), 
        .CO(C[201]) );
  FA_1862 \FAINST[201].FA_  ( .A(A[201]), .B(n458), .CI(C[201]), .S(S[201]), 
        .CO(C[202]) );
  FA_1861 \FAINST[202].FA_  ( .A(A[202]), .B(n459), .CI(C[202]), .S(S[202]), 
        .CO(C[203]) );
  FA_1860 \FAINST[203].FA_  ( .A(A[203]), .B(n460), .CI(C[203]), .S(S[203]), 
        .CO(C[204]) );
  FA_1859 \FAINST[204].FA_  ( .A(A[204]), .B(n461), .CI(C[204]), .S(S[204]), 
        .CO(C[205]) );
  FA_1858 \FAINST[205].FA_  ( .A(A[205]), .B(n462), .CI(C[205]), .S(S[205]), 
        .CO(C[206]) );
  FA_1857 \FAINST[206].FA_  ( .A(A[206]), .B(n463), .CI(C[206]), .S(S[206]), 
        .CO(C[207]) );
  FA_1856 \FAINST[207].FA_  ( .A(A[207]), .B(n464), .CI(C[207]), .S(S[207]), 
        .CO(C[208]) );
  FA_1855 \FAINST[208].FA_  ( .A(A[208]), .B(n465), .CI(C[208]), .S(S[208]), 
        .CO(C[209]) );
  FA_1854 \FAINST[209].FA_  ( .A(A[209]), .B(n466), .CI(C[209]), .S(S[209]), 
        .CO(C[210]) );
  FA_1853 \FAINST[210].FA_  ( .A(A[210]), .B(n467), .CI(C[210]), .S(S[210]), 
        .CO(C[211]) );
  FA_1852 \FAINST[211].FA_  ( .A(A[211]), .B(n468), .CI(C[211]), .S(S[211]), 
        .CO(C[212]) );
  FA_1851 \FAINST[212].FA_  ( .A(A[212]), .B(n469), .CI(C[212]), .S(S[212]), 
        .CO(C[213]) );
  FA_1850 \FAINST[213].FA_  ( .A(A[213]), .B(n470), .CI(C[213]), .S(S[213]), 
        .CO(C[214]) );
  FA_1849 \FAINST[214].FA_  ( .A(A[214]), .B(n471), .CI(C[214]), .S(S[214]), 
        .CO(C[215]) );
  FA_1848 \FAINST[215].FA_  ( .A(A[215]), .B(n472), .CI(C[215]), .S(S[215]), 
        .CO(C[216]) );
  FA_1847 \FAINST[216].FA_  ( .A(A[216]), .B(n473), .CI(C[216]), .S(S[216]), 
        .CO(C[217]) );
  FA_1846 \FAINST[217].FA_  ( .A(A[217]), .B(n474), .CI(C[217]), .S(S[217]), 
        .CO(C[218]) );
  FA_1845 \FAINST[218].FA_  ( .A(A[218]), .B(n475), .CI(C[218]), .S(S[218]), 
        .CO(C[219]) );
  FA_1844 \FAINST[219].FA_  ( .A(A[219]), .B(n476), .CI(C[219]), .S(S[219]), 
        .CO(C[220]) );
  FA_1843 \FAINST[220].FA_  ( .A(A[220]), .B(n477), .CI(C[220]), .S(S[220]), 
        .CO(C[221]) );
  FA_1842 \FAINST[221].FA_  ( .A(A[221]), .B(n478), .CI(C[221]), .S(S[221]), 
        .CO(C[222]) );
  FA_1841 \FAINST[222].FA_  ( .A(A[222]), .B(n479), .CI(C[222]), .S(S[222]), 
        .CO(C[223]) );
  FA_1840 \FAINST[223].FA_  ( .A(A[223]), .B(n480), .CI(C[223]), .S(S[223]), 
        .CO(C[224]) );
  FA_1839 \FAINST[224].FA_  ( .A(A[224]), .B(n481), .CI(C[224]), .S(S[224]), 
        .CO(C[225]) );
  FA_1838 \FAINST[225].FA_  ( .A(A[225]), .B(n482), .CI(C[225]), .S(S[225]), 
        .CO(C[226]) );
  FA_1837 \FAINST[226].FA_  ( .A(A[226]), .B(n483), .CI(C[226]), .S(S[226]), 
        .CO(C[227]) );
  FA_1836 \FAINST[227].FA_  ( .A(A[227]), .B(n484), .CI(C[227]), .S(S[227]), 
        .CO(C[228]) );
  FA_1835 \FAINST[228].FA_  ( .A(A[228]), .B(n485), .CI(C[228]), .S(S[228]), 
        .CO(C[229]) );
  FA_1834 \FAINST[229].FA_  ( .A(A[229]), .B(n486), .CI(C[229]), .S(S[229]), 
        .CO(C[230]) );
  FA_1833 \FAINST[230].FA_  ( .A(A[230]), .B(n487), .CI(C[230]), .S(S[230]), 
        .CO(C[231]) );
  FA_1832 \FAINST[231].FA_  ( .A(A[231]), .B(n488), .CI(C[231]), .S(S[231]), 
        .CO(C[232]) );
  FA_1831 \FAINST[232].FA_  ( .A(A[232]), .B(n489), .CI(C[232]), .S(S[232]), 
        .CO(C[233]) );
  FA_1830 \FAINST[233].FA_  ( .A(A[233]), .B(n490), .CI(C[233]), .S(S[233]), 
        .CO(C[234]) );
  FA_1829 \FAINST[234].FA_  ( .A(A[234]), .B(n491), .CI(C[234]), .S(S[234]), 
        .CO(C[235]) );
  FA_1828 \FAINST[235].FA_  ( .A(A[235]), .B(n492), .CI(C[235]), .S(S[235]), 
        .CO(C[236]) );
  FA_1827 \FAINST[236].FA_  ( .A(A[236]), .B(n493), .CI(C[236]), .S(S[236]), 
        .CO(C[237]) );
  FA_1826 \FAINST[237].FA_  ( .A(A[237]), .B(n494), .CI(C[237]), .S(S[237]), 
        .CO(C[238]) );
  FA_1825 \FAINST[238].FA_  ( .A(A[238]), .B(n495), .CI(C[238]), .S(S[238]), 
        .CO(C[239]) );
  FA_1824 \FAINST[239].FA_  ( .A(A[239]), .B(n496), .CI(C[239]), .S(S[239]), 
        .CO(C[240]) );
  FA_1823 \FAINST[240].FA_  ( .A(A[240]), .B(n497), .CI(C[240]), .S(S[240]), 
        .CO(C[241]) );
  FA_1822 \FAINST[241].FA_  ( .A(A[241]), .B(n498), .CI(C[241]), .S(S[241]), 
        .CO(C[242]) );
  FA_1821 \FAINST[242].FA_  ( .A(A[242]), .B(n499), .CI(C[242]), .S(S[242]), 
        .CO(C[243]) );
  FA_1820 \FAINST[243].FA_  ( .A(A[243]), .B(n500), .CI(C[243]), .S(S[243]), 
        .CO(C[244]) );
  FA_1819 \FAINST[244].FA_  ( .A(A[244]), .B(n501), .CI(C[244]), .S(S[244]), 
        .CO(C[245]) );
  FA_1818 \FAINST[245].FA_  ( .A(A[245]), .B(n502), .CI(C[245]), .S(S[245]), 
        .CO(C[246]) );
  FA_1817 \FAINST[246].FA_  ( .A(A[246]), .B(n503), .CI(C[246]), .S(S[246]), 
        .CO(C[247]) );
  FA_1816 \FAINST[247].FA_  ( .A(A[247]), .B(n504), .CI(C[247]), .S(S[247]), 
        .CO(C[248]) );
  FA_1815 \FAINST[248].FA_  ( .A(A[248]), .B(n505), .CI(C[248]), .S(S[248]), 
        .CO(C[249]) );
  FA_1814 \FAINST[249].FA_  ( .A(A[249]), .B(n506), .CI(C[249]), .S(S[249]), 
        .CO(C[250]) );
  FA_1813 \FAINST[250].FA_  ( .A(A[250]), .B(n507), .CI(C[250]), .S(S[250]), 
        .CO(C[251]) );
  FA_1812 \FAINST[251].FA_  ( .A(A[251]), .B(n508), .CI(C[251]), .S(S[251]), 
        .CO(C[252]) );
  FA_1811 \FAINST[252].FA_  ( .A(A[252]), .B(n509), .CI(C[252]), .S(S[252]), 
        .CO(C[253]) );
  FA_1810 \FAINST[253].FA_  ( .A(A[253]), .B(n510), .CI(C[253]), .S(S[253]), 
        .CO(C[254]) );
  FA_1809 \FAINST[254].FA_  ( .A(A[254]), .B(n511), .CI(C[254]), .S(S[254]), 
        .CO(C[255]) );
  FA_1808 \FAINST[255].FA_  ( .A(A[255]), .B(n512), .CI(C[255]), .S(S[255]), 
        .CO(C[256]) );
  FA_1807 \FAINST[256].FA_  ( .A(A[256]), .B(1'b1), .CI(C[256]), .S(S[256]), 
        .CO(C[257]) );
  FA_1806 \FAINST[257].FA_  ( .A(A[257]), .B(1'b1), .CI(C[257]), .S(S[257]) );
  IV U2 ( .A(B[159]), .Z(n416) );
  IV U3 ( .A(B[160]), .Z(n417) );
  IV U4 ( .A(B[161]), .Z(n418) );
  IV U5 ( .A(B[162]), .Z(n419) );
  IV U6 ( .A(B[163]), .Z(n420) );
  IV U7 ( .A(B[164]), .Z(n421) );
  IV U8 ( .A(B[165]), .Z(n422) );
  IV U9 ( .A(B[166]), .Z(n423) );
  IV U10 ( .A(B[167]), .Z(n424) );
  IV U11 ( .A(B[168]), .Z(n425) );
  IV U12 ( .A(B[249]), .Z(n506) );
  IV U13 ( .A(B[169]), .Z(n426) );
  IV U14 ( .A(B[170]), .Z(n427) );
  IV U15 ( .A(B[171]), .Z(n428) );
  IV U16 ( .A(B[172]), .Z(n429) );
  IV U17 ( .A(B[173]), .Z(n430) );
  IV U18 ( .A(B[174]), .Z(n431) );
  IV U19 ( .A(B[175]), .Z(n432) );
  IV U20 ( .A(B[176]), .Z(n433) );
  IV U21 ( .A(B[177]), .Z(n434) );
  IV U22 ( .A(B[178]), .Z(n435) );
  IV U23 ( .A(B[250]), .Z(n507) );
  IV U24 ( .A(B[179]), .Z(n436) );
  IV U25 ( .A(B[180]), .Z(n437) );
  IV U26 ( .A(B[181]), .Z(n438) );
  IV U27 ( .A(B[182]), .Z(n439) );
  IV U28 ( .A(B[183]), .Z(n440) );
  IV U29 ( .A(B[184]), .Z(n441) );
  IV U30 ( .A(B[185]), .Z(n442) );
  IV U31 ( .A(B[186]), .Z(n443) );
  IV U32 ( .A(B[187]), .Z(n444) );
  IV U33 ( .A(B[188]), .Z(n445) );
  IV U34 ( .A(B[251]), .Z(n508) );
  IV U35 ( .A(B[189]), .Z(n446) );
  IV U36 ( .A(B[190]), .Z(n447) );
  IV U37 ( .A(B[191]), .Z(n448) );
  IV U38 ( .A(B[192]), .Z(n449) );
  IV U39 ( .A(B[193]), .Z(n450) );
  IV U40 ( .A(B[194]), .Z(n451) );
  IV U41 ( .A(B[195]), .Z(n452) );
  IV U42 ( .A(B[196]), .Z(n453) );
  IV U43 ( .A(B[197]), .Z(n454) );
  IV U44 ( .A(B[198]), .Z(n455) );
  IV U45 ( .A(B[252]), .Z(n509) );
  IV U46 ( .A(B[199]), .Z(n456) );
  IV U47 ( .A(B[200]), .Z(n457) );
  IV U48 ( .A(B[201]), .Z(n458) );
  IV U49 ( .A(B[202]), .Z(n459) );
  IV U50 ( .A(B[203]), .Z(n460) );
  IV U51 ( .A(B[204]), .Z(n461) );
  IV U52 ( .A(B[205]), .Z(n462) );
  IV U53 ( .A(B[206]), .Z(n463) );
  IV U54 ( .A(B[207]), .Z(n464) );
  IV U55 ( .A(B[208]), .Z(n465) );
  IV U56 ( .A(B[253]), .Z(n510) );
  IV U57 ( .A(B[209]), .Z(n466) );
  IV U58 ( .A(B[210]), .Z(n467) );
  IV U59 ( .A(B[211]), .Z(n468) );
  IV U60 ( .A(B[212]), .Z(n469) );
  IV U61 ( .A(B[213]), .Z(n470) );
  IV U62 ( .A(B[214]), .Z(n471) );
  IV U63 ( .A(B[215]), .Z(n472) );
  IV U64 ( .A(B[216]), .Z(n473) );
  IV U65 ( .A(B[217]), .Z(n474) );
  IV U66 ( .A(B[218]), .Z(n475) );
  IV U67 ( .A(B[254]), .Z(n511) );
  IV U68 ( .A(B[219]), .Z(n476) );
  IV U69 ( .A(B[220]), .Z(n477) );
  IV U70 ( .A(B[221]), .Z(n478) );
  IV U71 ( .A(B[222]), .Z(n479) );
  IV U72 ( .A(B[223]), .Z(n480) );
  IV U73 ( .A(B[224]), .Z(n481) );
  IV U74 ( .A(B[225]), .Z(n482) );
  IV U75 ( .A(B[226]), .Z(n483) );
  IV U76 ( .A(B[227]), .Z(n484) );
  IV U77 ( .A(B[228]), .Z(n485) );
  IV U78 ( .A(B[255]), .Z(n512) );
  IV U79 ( .A(B[229]), .Z(n486) );
  IV U80 ( .A(B[230]), .Z(n487) );
  IV U81 ( .A(B[231]), .Z(n488) );
  IV U82 ( .A(B[232]), .Z(n489) );
  IV U83 ( .A(B[0]), .Z(n2) );
  IV U84 ( .A(B[1]), .Z(n258) );
  IV U85 ( .A(B[2]), .Z(n259) );
  IV U86 ( .A(B[3]), .Z(n260) );
  IV U87 ( .A(B[4]), .Z(n261) );
  IV U88 ( .A(B[5]), .Z(n262) );
  IV U89 ( .A(B[6]), .Z(n263) );
  IV U90 ( .A(B[7]), .Z(n264) );
  IV U91 ( .A(B[8]), .Z(n265) );
  IV U92 ( .A(B[233]), .Z(n490) );
  IV U93 ( .A(B[9]), .Z(n266) );
  IV U94 ( .A(B[10]), .Z(n267) );
  IV U95 ( .A(B[11]), .Z(n268) );
  IV U96 ( .A(B[12]), .Z(n269) );
  IV U97 ( .A(B[13]), .Z(n270) );
  IV U98 ( .A(B[14]), .Z(n271) );
  IV U99 ( .A(B[15]), .Z(n272) );
  IV U100 ( .A(B[16]), .Z(n273) );
  IV U101 ( .A(B[17]), .Z(n274) );
  IV U102 ( .A(B[18]), .Z(n275) );
  IV U103 ( .A(B[234]), .Z(n491) );
  IV U104 ( .A(B[19]), .Z(n276) );
  IV U105 ( .A(B[20]), .Z(n277) );
  IV U106 ( .A(B[21]), .Z(n278) );
  IV U107 ( .A(B[22]), .Z(n279) );
  IV U108 ( .A(B[23]), .Z(n280) );
  IV U109 ( .A(B[24]), .Z(n281) );
  IV U110 ( .A(B[25]), .Z(n282) );
  IV U111 ( .A(B[26]), .Z(n283) );
  IV U112 ( .A(B[27]), .Z(n284) );
  IV U113 ( .A(B[28]), .Z(n285) );
  IV U114 ( .A(B[235]), .Z(n492) );
  IV U115 ( .A(B[29]), .Z(n286) );
  IV U116 ( .A(B[30]), .Z(n287) );
  IV U117 ( .A(B[31]), .Z(n288) );
  IV U118 ( .A(B[32]), .Z(n289) );
  IV U119 ( .A(B[33]), .Z(n290) );
  IV U120 ( .A(B[34]), .Z(n291) );
  IV U121 ( .A(B[35]), .Z(n292) );
  IV U122 ( .A(B[36]), .Z(n293) );
  IV U123 ( .A(B[37]), .Z(n294) );
  IV U124 ( .A(B[38]), .Z(n295) );
  IV U125 ( .A(B[236]), .Z(n493) );
  IV U126 ( .A(B[39]), .Z(n296) );
  IV U127 ( .A(B[40]), .Z(n297) );
  IV U128 ( .A(B[41]), .Z(n298) );
  IV U129 ( .A(B[42]), .Z(n299) );
  IV U130 ( .A(B[43]), .Z(n300) );
  IV U131 ( .A(B[44]), .Z(n301) );
  IV U132 ( .A(B[45]), .Z(n302) );
  IV U133 ( .A(B[46]), .Z(n303) );
  IV U134 ( .A(B[47]), .Z(n304) );
  IV U135 ( .A(B[48]), .Z(n305) );
  IV U136 ( .A(B[237]), .Z(n494) );
  IV U137 ( .A(B[49]), .Z(n306) );
  IV U138 ( .A(B[50]), .Z(n307) );
  IV U139 ( .A(B[51]), .Z(n308) );
  IV U140 ( .A(B[52]), .Z(n309) );
  IV U141 ( .A(B[53]), .Z(n310) );
  IV U142 ( .A(B[54]), .Z(n311) );
  IV U143 ( .A(B[55]), .Z(n312) );
  IV U144 ( .A(B[56]), .Z(n313) );
  IV U145 ( .A(B[57]), .Z(n314) );
  IV U146 ( .A(B[58]), .Z(n315) );
  IV U147 ( .A(B[238]), .Z(n495) );
  IV U148 ( .A(B[59]), .Z(n316) );
  IV U149 ( .A(B[60]), .Z(n317) );
  IV U150 ( .A(B[61]), .Z(n318) );
  IV U151 ( .A(B[62]), .Z(n319) );
  IV U152 ( .A(B[63]), .Z(n320) );
  IV U153 ( .A(B[64]), .Z(n321) );
  IV U154 ( .A(B[65]), .Z(n322) );
  IV U155 ( .A(B[66]), .Z(n323) );
  IV U156 ( .A(B[67]), .Z(n324) );
  IV U157 ( .A(B[68]), .Z(n325) );
  IV U158 ( .A(B[239]), .Z(n496) );
  IV U159 ( .A(B[69]), .Z(n326) );
  IV U160 ( .A(B[70]), .Z(n327) );
  IV U161 ( .A(B[71]), .Z(n328) );
  IV U162 ( .A(B[72]), .Z(n329) );
  IV U163 ( .A(B[73]), .Z(n330) );
  IV U164 ( .A(B[74]), .Z(n331) );
  IV U165 ( .A(B[75]), .Z(n332) );
  IV U166 ( .A(B[76]), .Z(n333) );
  IV U167 ( .A(B[77]), .Z(n334) );
  IV U168 ( .A(B[78]), .Z(n335) );
  IV U169 ( .A(B[240]), .Z(n497) );
  IV U170 ( .A(B[79]), .Z(n336) );
  IV U171 ( .A(B[80]), .Z(n337) );
  IV U172 ( .A(B[81]), .Z(n338) );
  IV U173 ( .A(B[82]), .Z(n339) );
  IV U174 ( .A(B[83]), .Z(n340) );
  IV U175 ( .A(B[84]), .Z(n341) );
  IV U176 ( .A(B[85]), .Z(n342) );
  IV U177 ( .A(B[86]), .Z(n343) );
  IV U178 ( .A(B[87]), .Z(n344) );
  IV U179 ( .A(B[88]), .Z(n345) );
  IV U180 ( .A(B[241]), .Z(n498) );
  IV U181 ( .A(B[89]), .Z(n346) );
  IV U182 ( .A(B[90]), .Z(n347) );
  IV U183 ( .A(B[91]), .Z(n348) );
  IV U184 ( .A(B[92]), .Z(n349) );
  IV U185 ( .A(B[93]), .Z(n350) );
  IV U186 ( .A(B[94]), .Z(n351) );
  IV U187 ( .A(B[95]), .Z(n352) );
  IV U188 ( .A(B[96]), .Z(n353) );
  IV U189 ( .A(B[97]), .Z(n354) );
  IV U190 ( .A(B[98]), .Z(n355) );
  IV U191 ( .A(B[242]), .Z(n499) );
  IV U192 ( .A(B[99]), .Z(n356) );
  IV U193 ( .A(B[100]), .Z(n357) );
  IV U194 ( .A(B[101]), .Z(n358) );
  IV U195 ( .A(B[102]), .Z(n359) );
  IV U196 ( .A(B[103]), .Z(n360) );
  IV U197 ( .A(B[104]), .Z(n361) );
  IV U198 ( .A(B[105]), .Z(n362) );
  IV U199 ( .A(B[106]), .Z(n363) );
  IV U200 ( .A(B[107]), .Z(n364) );
  IV U201 ( .A(B[108]), .Z(n365) );
  IV U202 ( .A(B[243]), .Z(n500) );
  IV U203 ( .A(B[109]), .Z(n366) );
  IV U204 ( .A(B[110]), .Z(n367) );
  IV U205 ( .A(B[111]), .Z(n368) );
  IV U206 ( .A(B[112]), .Z(n369) );
  IV U207 ( .A(B[113]), .Z(n370) );
  IV U208 ( .A(B[114]), .Z(n371) );
  IV U209 ( .A(B[115]), .Z(n372) );
  IV U210 ( .A(B[116]), .Z(n373) );
  IV U211 ( .A(B[117]), .Z(n374) );
  IV U212 ( .A(B[118]), .Z(n375) );
  IV U213 ( .A(B[244]), .Z(n501) );
  IV U214 ( .A(B[119]), .Z(n376) );
  IV U215 ( .A(B[120]), .Z(n377) );
  IV U216 ( .A(B[121]), .Z(n378) );
  IV U217 ( .A(B[122]), .Z(n379) );
  IV U218 ( .A(B[123]), .Z(n380) );
  IV U219 ( .A(B[124]), .Z(n381) );
  IV U220 ( .A(B[125]), .Z(n382) );
  IV U221 ( .A(B[126]), .Z(n383) );
  IV U222 ( .A(B[127]), .Z(n384) );
  IV U223 ( .A(B[128]), .Z(n385) );
  IV U224 ( .A(B[245]), .Z(n502) );
  IV U225 ( .A(B[129]), .Z(n386) );
  IV U226 ( .A(B[130]), .Z(n387) );
  IV U227 ( .A(B[131]), .Z(n388) );
  IV U228 ( .A(B[132]), .Z(n389) );
  IV U229 ( .A(B[133]), .Z(n390) );
  IV U230 ( .A(B[134]), .Z(n391) );
  IV U231 ( .A(B[135]), .Z(n392) );
  IV U232 ( .A(B[136]), .Z(n393) );
  IV U233 ( .A(B[137]), .Z(n394) );
  IV U234 ( .A(B[138]), .Z(n395) );
  IV U235 ( .A(B[246]), .Z(n503) );
  IV U236 ( .A(B[139]), .Z(n396) );
  IV U237 ( .A(B[140]), .Z(n397) );
  IV U238 ( .A(B[141]), .Z(n398) );
  IV U239 ( .A(B[142]), .Z(n399) );
  IV U240 ( .A(B[143]), .Z(n400) );
  IV U241 ( .A(B[144]), .Z(n401) );
  IV U242 ( .A(B[145]), .Z(n402) );
  IV U243 ( .A(B[146]), .Z(n403) );
  IV U244 ( .A(B[147]), .Z(n404) );
  IV U245 ( .A(B[148]), .Z(n405) );
  IV U246 ( .A(B[247]), .Z(n504) );
  IV U247 ( .A(B[149]), .Z(n406) );
  IV U248 ( .A(B[150]), .Z(n407) );
  IV U249 ( .A(B[151]), .Z(n408) );
  IV U250 ( .A(B[152]), .Z(n409) );
  IV U251 ( .A(B[153]), .Z(n410) );
  IV U252 ( .A(B[154]), .Z(n411) );
  IV U253 ( .A(B[155]), .Z(n412) );
  IV U254 ( .A(B[156]), .Z(n413) );
  IV U255 ( .A(B[157]), .Z(n414) );
  IV U256 ( .A(B[158]), .Z(n415) );
  IV U257 ( .A(B[248]), .Z(n505) );
endmodule


module modmult_step_N256_1_1 ( xregN_1, y, n, zin, zout );
  input [255:0] y;
  input [255:0] n;
  input [257:0] zin;
  output [257:0] zout;
  input xregN_1;
  wire   c1, c2, n4;
  wire   [257:0] w1;
  wire   [257:0] w2;
  wire   [257:0] w3;
  wire   [257:0] z2;
  wire   [257:0] z3;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6;

  MUX_N258_6 MUX_1 ( .A({1'b0, 1'b0, y}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .S(xregN_1), .O({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, w1[255:0]}) );
  MUX_N258_5 MUX_2 ( .A({1'b0, 1'b0, n}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .S(c1), .O({SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        w2[255:0]}) );
  MUX_N258_4 MUX_3 ( .A({1'b0, 1'b0, n}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .S(n4), .O({SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        w3[255:0]}) );
  ADD_N258_1_1 ADD_1 ( .A({zin[256:0], 1'b0}), .B({1'b0, 1'b0, w1[255:0]}), 
        .CI(1'b0), .S(z2) );
  COMP_N258_4 COMP_1 ( .A(z2), .B({1'b0, 1'b0, n}), .O(c1) );
  SUB_N258_4 SUB_1 ( .A(z2), .B({1'b0, 1'b0, w2[255:0]}), .S(z3) );
  COMP_N258_3 COMP_2 ( .A({1'b0, 1'b0, n}), .B(z3), .O(c2) );
  SUB_N258_3 SUB_2 ( .A({1'b0, z3[256:0]}), .B({1'b0, 1'b0, w3[255:0]}), .S({
        SYNOPSYS_UNCONNECTED__6, zout[256:0]}) );
  IV U2 ( .A(c2), .Z(n4) );
endmodule


module modmult_N256_CC128 ( clk, rst, start, x, y, n, o );
  input [255:0] x;
  input [255:0] y;
  input [255:0] n;
  output [255:0] o;
  input clk, rst, start;
  wire   \zout[1][256] , \zin[1][256] , \zin[1][255] , \zin[1][254] ,
         \zin[1][253] , \zin[1][252] , \zin[1][251] , \zin[1][250] ,
         \zin[1][249] , \zin[1][248] , \zin[1][247] , \zin[1][246] ,
         \zin[1][245] , \zin[1][244] , \zin[1][243] , \zin[1][242] ,
         \zin[1][241] , \zin[1][240] , \zin[1][239] , \zin[1][238] ,
         \zin[1][237] , \zin[1][236] , \zin[1][235] , \zin[1][234] ,
         \zin[1][233] , \zin[1][232] , \zin[1][231] , \zin[1][230] ,
         \zin[1][229] , \zin[1][228] , \zin[1][227] , \zin[1][226] ,
         \zin[1][225] , \zin[1][224] , \zin[1][223] , \zin[1][222] ,
         \zin[1][221] , \zin[1][220] , \zin[1][219] , \zin[1][218] ,
         \zin[1][217] , \zin[1][216] , \zin[1][215] , \zin[1][214] ,
         \zin[1][213] , \zin[1][212] , \zin[1][211] , \zin[1][210] ,
         \zin[1][209] , \zin[1][208] , \zin[1][207] , \zin[1][206] ,
         \zin[1][205] , \zin[1][204] , \zin[1][203] , \zin[1][202] ,
         \zin[1][201] , \zin[1][200] , \zin[1][199] , \zin[1][198] ,
         \zin[1][197] , \zin[1][196] , \zin[1][195] , \zin[1][194] ,
         \zin[1][193] , \zin[1][192] , \zin[1][191] , \zin[1][190] ,
         \zin[1][189] , \zin[1][188] , \zin[1][187] , \zin[1][186] ,
         \zin[1][185] , \zin[1][184] , \zin[1][183] , \zin[1][182] ,
         \zin[1][181] , \zin[1][180] , \zin[1][179] , \zin[1][178] ,
         \zin[1][177] , \zin[1][176] , \zin[1][175] , \zin[1][174] ,
         \zin[1][173] , \zin[1][172] , \zin[1][171] , \zin[1][170] ,
         \zin[1][169] , \zin[1][168] , \zin[1][167] , \zin[1][166] ,
         \zin[1][165] , \zin[1][164] , \zin[1][163] , \zin[1][162] ,
         \zin[1][161] , \zin[1][160] , \zin[1][159] , \zin[1][158] ,
         \zin[1][157] , \zin[1][156] , \zin[1][155] , \zin[1][154] ,
         \zin[1][153] , \zin[1][152] , \zin[1][151] , \zin[1][150] ,
         \zin[1][149] , \zin[1][148] , \zin[1][147] , \zin[1][146] ,
         \zin[1][145] , \zin[1][144] , \zin[1][143] , \zin[1][142] ,
         \zin[1][141] , \zin[1][140] , \zin[1][139] , \zin[1][138] ,
         \zin[1][137] , \zin[1][136] , \zin[1][135] , \zin[1][134] ,
         \zin[1][133] , \zin[1][132] , \zin[1][131] , \zin[1][130] ,
         \zin[1][129] , \zin[1][128] , \zin[1][127] , \zin[1][126] ,
         \zin[1][125] , \zin[1][124] , \zin[1][123] , \zin[1][122] ,
         \zin[1][121] , \zin[1][120] , \zin[1][119] , \zin[1][118] ,
         \zin[1][117] , \zin[1][116] , \zin[1][115] , \zin[1][114] ,
         \zin[1][113] , \zin[1][112] , \zin[1][111] , \zin[1][110] ,
         \zin[1][109] , \zin[1][108] , \zin[1][107] , \zin[1][106] ,
         \zin[1][105] , \zin[1][104] , \zin[1][103] , \zin[1][102] ,
         \zin[1][101] , \zin[1][100] , \zin[1][99] , \zin[1][98] ,
         \zin[1][97] , \zin[1][96] , \zin[1][95] , \zin[1][94] , \zin[1][93] ,
         \zin[1][92] , \zin[1][91] , \zin[1][90] , \zin[1][89] , \zin[1][88] ,
         \zin[1][87] , \zin[1][86] , \zin[1][85] , \zin[1][84] , \zin[1][83] ,
         \zin[1][82] , \zin[1][81] , \zin[1][80] , \zin[1][79] , \zin[1][78] ,
         \zin[1][77] , \zin[1][76] , \zin[1][75] , \zin[1][74] , \zin[1][73] ,
         \zin[1][72] , \zin[1][71] , \zin[1][70] , \zin[1][69] , \zin[1][68] ,
         \zin[1][67] , \zin[1][66] , \zin[1][65] , \zin[1][64] , \zin[1][63] ,
         \zin[1][62] , \zin[1][61] , \zin[1][60] , \zin[1][59] , \zin[1][58] ,
         \zin[1][57] , \zin[1][56] , \zin[1][55] , \zin[1][54] , \zin[1][53] ,
         \zin[1][52] , \zin[1][51] , \zin[1][50] , \zin[1][49] , \zin[1][48] ,
         \zin[1][47] , \zin[1][46] , \zin[1][45] , \zin[1][44] , \zin[1][43] ,
         \zin[1][42] , \zin[1][41] , \zin[1][40] , \zin[1][39] , \zin[1][38] ,
         \zin[1][37] , \zin[1][36] , \zin[1][35] , \zin[1][34] , \zin[1][33] ,
         \zin[1][32] , \zin[1][31] , \zin[1][30] , \zin[1][29] , \zin[1][28] ,
         \zin[1][27] , \zin[1][26] , \zin[1][25] , \zin[1][24] , \zin[1][23] ,
         \zin[1][22] , \zin[1][21] , \zin[1][20] , \zin[1][19] , \zin[1][18] ,
         \zin[1][17] , \zin[1][16] , \zin[1][15] , \zin[1][14] , \zin[1][13] ,
         \zin[1][12] , \zin[1][11] , \zin[1][10] , \zin[1][9] , \zin[1][8] ,
         \zin[1][7] , \zin[1][6] , \zin[1][5] , \zin[1][4] , \zin[1][3] ,
         \zin[1][2] , \zin[1][1] , \zin[1][0] , \zin[0][256] , \zin[0][255] ,
         \zin[0][254] , \zin[0][253] , \zin[0][252] , \zin[0][251] ,
         \zin[0][250] , \zin[0][249] , \zin[0][248] , \zin[0][247] ,
         \zin[0][246] , \zin[0][245] , \zin[0][244] , \zin[0][243] ,
         \zin[0][242] , \zin[0][241] , \zin[0][240] , \zin[0][239] ,
         \zin[0][238] , \zin[0][237] , \zin[0][236] , \zin[0][235] ,
         \zin[0][234] , \zin[0][233] , \zin[0][232] , \zin[0][231] ,
         \zin[0][230] , \zin[0][229] , \zin[0][228] , \zin[0][227] ,
         \zin[0][226] , \zin[0][225] , \zin[0][224] , \zin[0][223] ,
         \zin[0][222] , \zin[0][221] , \zin[0][220] , \zin[0][219] ,
         \zin[0][218] , \zin[0][217] , \zin[0][216] , \zin[0][215] ,
         \zin[0][214] , \zin[0][213] , \zin[0][212] , \zin[0][211] ,
         \zin[0][210] , \zin[0][209] , \zin[0][208] , \zin[0][207] ,
         \zin[0][206] , \zin[0][205] , \zin[0][204] , \zin[0][203] ,
         \zin[0][202] , \zin[0][201] , \zin[0][200] , \zin[0][199] ,
         \zin[0][198] , \zin[0][197] , \zin[0][196] , \zin[0][195] ,
         \zin[0][194] , \zin[0][193] , \zin[0][192] , \zin[0][191] ,
         \zin[0][190] , \zin[0][189] , \zin[0][188] , \zin[0][187] ,
         \zin[0][186] , \zin[0][185] , \zin[0][184] , \zin[0][183] ,
         \zin[0][182] , \zin[0][181] , \zin[0][180] , \zin[0][179] ,
         \zin[0][178] , \zin[0][177] , \zin[0][176] , \zin[0][175] ,
         \zin[0][174] , \zin[0][173] , \zin[0][172] , \zin[0][171] ,
         \zin[0][170] , \zin[0][169] , \zin[0][168] , \zin[0][167] ,
         \zin[0][166] , \zin[0][165] , \zin[0][164] , \zin[0][163] ,
         \zin[0][162] , \zin[0][161] , \zin[0][160] , \zin[0][159] ,
         \zin[0][158] , \zin[0][157] , \zin[0][156] , \zin[0][155] ,
         \zin[0][154] , \zin[0][153] , \zin[0][152] , \zin[0][151] ,
         \zin[0][150] , \zin[0][149] , \zin[0][148] , \zin[0][147] ,
         \zin[0][146] , \zin[0][145] , \zin[0][144] , \zin[0][143] ,
         \zin[0][142] , \zin[0][141] , \zin[0][140] , \zin[0][139] ,
         \zin[0][138] , \zin[0][137] , \zin[0][136] , \zin[0][135] ,
         \zin[0][134] , \zin[0][133] , \zin[0][132] , \zin[0][131] ,
         \zin[0][130] , \zin[0][129] , \zin[0][128] , \zin[0][127] ,
         \zin[0][126] , \zin[0][125] , \zin[0][124] , \zin[0][123] ,
         \zin[0][122] , \zin[0][121] , \zin[0][120] , \zin[0][119] ,
         \zin[0][118] , \zin[0][117] , \zin[0][116] , \zin[0][115] ,
         \zin[0][114] , \zin[0][113] , \zin[0][112] , \zin[0][111] ,
         \zin[0][110] , \zin[0][109] , \zin[0][108] , \zin[0][107] ,
         \zin[0][106] , \zin[0][105] , \zin[0][104] , \zin[0][103] ,
         \zin[0][102] , \zin[0][101] , \zin[0][100] , \zin[0][99] ,
         \zin[0][98] , \zin[0][97] , \zin[0][96] , \zin[0][95] , \zin[0][94] ,
         \zin[0][93] , \zin[0][92] , \zin[0][91] , \zin[0][90] , \zin[0][89] ,
         \zin[0][88] , \zin[0][87] , \zin[0][86] , \zin[0][85] , \zin[0][84] ,
         \zin[0][83] , \zin[0][82] , \zin[0][81] , \zin[0][80] , \zin[0][79] ,
         \zin[0][78] , \zin[0][77] , \zin[0][76] , \zin[0][75] , \zin[0][74] ,
         \zin[0][73] , \zin[0][72] , \zin[0][71] , \zin[0][70] , \zin[0][69] ,
         \zin[0][68] , \zin[0][67] , \zin[0][66] , \zin[0][65] , \zin[0][64] ,
         \zin[0][63] , \zin[0][62] , \zin[0][61] , \zin[0][60] , \zin[0][59] ,
         \zin[0][58] , \zin[0][57] , \zin[0][56] , \zin[0][55] , \zin[0][54] ,
         \zin[0][53] , \zin[0][52] , \zin[0][51] , \zin[0][50] , \zin[0][49] ,
         \zin[0][48] , \zin[0][47] , \zin[0][46] , \zin[0][45] , \zin[0][44] ,
         \zin[0][43] , \zin[0][42] , \zin[0][41] , \zin[0][40] , \zin[0][39] ,
         \zin[0][38] , \zin[0][37] , \zin[0][36] , \zin[0][35] , \zin[0][34] ,
         \zin[0][33] , \zin[0][32] , \zin[0][31] , \zin[0][30] , \zin[0][29] ,
         \zin[0][28] , \zin[0][27] , \zin[0][26] , \zin[0][25] , \zin[0][24] ,
         \zin[0][23] , \zin[0][22] , \zin[0][21] , \zin[0][20] , \zin[0][19] ,
         \zin[0][18] , \zin[0][17] , \zin[0][16] , \zin[0][15] , \zin[0][14] ,
         \zin[0][13] , \zin[0][12] , \zin[0][11] , \zin[0][10] , \zin[0][9] ,
         \zin[0][8] , \zin[0][7] , \zin[0][6] , \zin[0][5] , \zin[0][4] ,
         \zin[0][3] , \zin[0][2] , \zin[0][1] , \zin[0][0] ;
  wire   [255:0] xin;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;

  modmult_step_N256_1_0 \MODMULT_STEP[0].modmult_step_  ( .xregN_1(xin[255]), 
        .y(y), .n(n), .zin({1'b0, \zin[0][256] , \zin[0][255] , \zin[0][254] , 
        \zin[0][253] , \zin[0][252] , \zin[0][251] , \zin[0][250] , 
        \zin[0][249] , \zin[0][248] , \zin[0][247] , \zin[0][246] , 
        \zin[0][245] , \zin[0][244] , \zin[0][243] , \zin[0][242] , 
        \zin[0][241] , \zin[0][240] , \zin[0][239] , \zin[0][238] , 
        \zin[0][237] , \zin[0][236] , \zin[0][235] , \zin[0][234] , 
        \zin[0][233] , \zin[0][232] , \zin[0][231] , \zin[0][230] , 
        \zin[0][229] , \zin[0][228] , \zin[0][227] , \zin[0][226] , 
        \zin[0][225] , \zin[0][224] , \zin[0][223] , \zin[0][222] , 
        \zin[0][221] , \zin[0][220] , \zin[0][219] , \zin[0][218] , 
        \zin[0][217] , \zin[0][216] , \zin[0][215] , \zin[0][214] , 
        \zin[0][213] , \zin[0][212] , \zin[0][211] , \zin[0][210] , 
        \zin[0][209] , \zin[0][208] , \zin[0][207] , \zin[0][206] , 
        \zin[0][205] , \zin[0][204] , \zin[0][203] , \zin[0][202] , 
        \zin[0][201] , \zin[0][200] , \zin[0][199] , \zin[0][198] , 
        \zin[0][197] , \zin[0][196] , \zin[0][195] , \zin[0][194] , 
        \zin[0][193] , \zin[0][192] , \zin[0][191] , \zin[0][190] , 
        \zin[0][189] , \zin[0][188] , \zin[0][187] , \zin[0][186] , 
        \zin[0][185] , \zin[0][184] , \zin[0][183] , \zin[0][182] , 
        \zin[0][181] , \zin[0][180] , \zin[0][179] , \zin[0][178] , 
        \zin[0][177] , \zin[0][176] , \zin[0][175] , \zin[0][174] , 
        \zin[0][173] , \zin[0][172] , \zin[0][171] , \zin[0][170] , 
        \zin[0][169] , \zin[0][168] , \zin[0][167] , \zin[0][166] , 
        \zin[0][165] , \zin[0][164] , \zin[0][163] , \zin[0][162] , 
        \zin[0][161] , \zin[0][160] , \zin[0][159] , \zin[0][158] , 
        \zin[0][157] , \zin[0][156] , \zin[0][155] , \zin[0][154] , 
        \zin[0][153] , \zin[0][152] , \zin[0][151] , \zin[0][150] , 
        \zin[0][149] , \zin[0][148] , \zin[0][147] , \zin[0][146] , 
        \zin[0][145] , \zin[0][144] , \zin[0][143] , \zin[0][142] , 
        \zin[0][141] , \zin[0][140] , \zin[0][139] , \zin[0][138] , 
        \zin[0][137] , \zin[0][136] , \zin[0][135] , \zin[0][134] , 
        \zin[0][133] , \zin[0][132] , \zin[0][131] , \zin[0][130] , 
        \zin[0][129] , \zin[0][128] , \zin[0][127] , \zin[0][126] , 
        \zin[0][125] , \zin[0][124] , \zin[0][123] , \zin[0][122] , 
        \zin[0][121] , \zin[0][120] , \zin[0][119] , \zin[0][118] , 
        \zin[0][117] , \zin[0][116] , \zin[0][115] , \zin[0][114] , 
        \zin[0][113] , \zin[0][112] , \zin[0][111] , \zin[0][110] , 
        \zin[0][109] , \zin[0][108] , \zin[0][107] , \zin[0][106] , 
        \zin[0][105] , \zin[0][104] , \zin[0][103] , \zin[0][102] , 
        \zin[0][101] , \zin[0][100] , \zin[0][99] , \zin[0][98] , \zin[0][97] , 
        \zin[0][96] , \zin[0][95] , \zin[0][94] , \zin[0][93] , \zin[0][92] , 
        \zin[0][91] , \zin[0][90] , \zin[0][89] , \zin[0][88] , \zin[0][87] , 
        \zin[0][86] , \zin[0][85] , \zin[0][84] , \zin[0][83] , \zin[0][82] , 
        \zin[0][81] , \zin[0][80] , \zin[0][79] , \zin[0][78] , \zin[0][77] , 
        \zin[0][76] , \zin[0][75] , \zin[0][74] , \zin[0][73] , \zin[0][72] , 
        \zin[0][71] , \zin[0][70] , \zin[0][69] , \zin[0][68] , \zin[0][67] , 
        \zin[0][66] , \zin[0][65] , \zin[0][64] , \zin[0][63] , \zin[0][62] , 
        \zin[0][61] , \zin[0][60] , \zin[0][59] , \zin[0][58] , \zin[0][57] , 
        \zin[0][56] , \zin[0][55] , \zin[0][54] , \zin[0][53] , \zin[0][52] , 
        \zin[0][51] , \zin[0][50] , \zin[0][49] , \zin[0][48] , \zin[0][47] , 
        \zin[0][46] , \zin[0][45] , \zin[0][44] , \zin[0][43] , \zin[0][42] , 
        \zin[0][41] , \zin[0][40] , \zin[0][39] , \zin[0][38] , \zin[0][37] , 
        \zin[0][36] , \zin[0][35] , \zin[0][34] , \zin[0][33] , \zin[0][32] , 
        \zin[0][31] , \zin[0][30] , \zin[0][29] , \zin[0][28] , \zin[0][27] , 
        \zin[0][26] , \zin[0][25] , \zin[0][24] , \zin[0][23] , \zin[0][22] , 
        \zin[0][21] , \zin[0][20] , \zin[0][19] , \zin[0][18] , \zin[0][17] , 
        \zin[0][16] , \zin[0][15] , \zin[0][14] , \zin[0][13] , \zin[0][12] , 
        \zin[0][11] , \zin[0][10] , \zin[0][9] , \zin[0][8] , \zin[0][7] , 
        \zin[0][6] , \zin[0][5] , \zin[0][4] , \zin[0][3] , \zin[0][2] , 
        \zin[0][1] , \zin[0][0] }), .zout({SYNOPSYS_UNCONNECTED__0, 
        \zin[1][256] , \zin[1][255] , \zin[1][254] , \zin[1][253] , 
        \zin[1][252] , \zin[1][251] , \zin[1][250] , \zin[1][249] , 
        \zin[1][248] , \zin[1][247] , \zin[1][246] , \zin[1][245] , 
        \zin[1][244] , \zin[1][243] , \zin[1][242] , \zin[1][241] , 
        \zin[1][240] , \zin[1][239] , \zin[1][238] , \zin[1][237] , 
        \zin[1][236] , \zin[1][235] , \zin[1][234] , \zin[1][233] , 
        \zin[1][232] , \zin[1][231] , \zin[1][230] , \zin[1][229] , 
        \zin[1][228] , \zin[1][227] , \zin[1][226] , \zin[1][225] , 
        \zin[1][224] , \zin[1][223] , \zin[1][222] , \zin[1][221] , 
        \zin[1][220] , \zin[1][219] , \zin[1][218] , \zin[1][217] , 
        \zin[1][216] , \zin[1][215] , \zin[1][214] , \zin[1][213] , 
        \zin[1][212] , \zin[1][211] , \zin[1][210] , \zin[1][209] , 
        \zin[1][208] , \zin[1][207] , \zin[1][206] , \zin[1][205] , 
        \zin[1][204] , \zin[1][203] , \zin[1][202] , \zin[1][201] , 
        \zin[1][200] , \zin[1][199] , \zin[1][198] , \zin[1][197] , 
        \zin[1][196] , \zin[1][195] , \zin[1][194] , \zin[1][193] , 
        \zin[1][192] , \zin[1][191] , \zin[1][190] , \zin[1][189] , 
        \zin[1][188] , \zin[1][187] , \zin[1][186] , \zin[1][185] , 
        \zin[1][184] , \zin[1][183] , \zin[1][182] , \zin[1][181] , 
        \zin[1][180] , \zin[1][179] , \zin[1][178] , \zin[1][177] , 
        \zin[1][176] , \zin[1][175] , \zin[1][174] , \zin[1][173] , 
        \zin[1][172] , \zin[1][171] , \zin[1][170] , \zin[1][169] , 
        \zin[1][168] , \zin[1][167] , \zin[1][166] , \zin[1][165] , 
        \zin[1][164] , \zin[1][163] , \zin[1][162] , \zin[1][161] , 
        \zin[1][160] , \zin[1][159] , \zin[1][158] , \zin[1][157] , 
        \zin[1][156] , \zin[1][155] , \zin[1][154] , \zin[1][153] , 
        \zin[1][152] , \zin[1][151] , \zin[1][150] , \zin[1][149] , 
        \zin[1][148] , \zin[1][147] , \zin[1][146] , \zin[1][145] , 
        \zin[1][144] , \zin[1][143] , \zin[1][142] , \zin[1][141] , 
        \zin[1][140] , \zin[1][139] , \zin[1][138] , \zin[1][137] , 
        \zin[1][136] , \zin[1][135] , \zin[1][134] , \zin[1][133] , 
        \zin[1][132] , \zin[1][131] , \zin[1][130] , \zin[1][129] , 
        \zin[1][128] , \zin[1][127] , \zin[1][126] , \zin[1][125] , 
        \zin[1][124] , \zin[1][123] , \zin[1][122] , \zin[1][121] , 
        \zin[1][120] , \zin[1][119] , \zin[1][118] , \zin[1][117] , 
        \zin[1][116] , \zin[1][115] , \zin[1][114] , \zin[1][113] , 
        \zin[1][112] , \zin[1][111] , \zin[1][110] , \zin[1][109] , 
        \zin[1][108] , \zin[1][107] , \zin[1][106] , \zin[1][105] , 
        \zin[1][104] , \zin[1][103] , \zin[1][102] , \zin[1][101] , 
        \zin[1][100] , \zin[1][99] , \zin[1][98] , \zin[1][97] , \zin[1][96] , 
        \zin[1][95] , \zin[1][94] , \zin[1][93] , \zin[1][92] , \zin[1][91] , 
        \zin[1][90] , \zin[1][89] , \zin[1][88] , \zin[1][87] , \zin[1][86] , 
        \zin[1][85] , \zin[1][84] , \zin[1][83] , \zin[1][82] , \zin[1][81] , 
        \zin[1][80] , \zin[1][79] , \zin[1][78] , \zin[1][77] , \zin[1][76] , 
        \zin[1][75] , \zin[1][74] , \zin[1][73] , \zin[1][72] , \zin[1][71] , 
        \zin[1][70] , \zin[1][69] , \zin[1][68] , \zin[1][67] , \zin[1][66] , 
        \zin[1][65] , \zin[1][64] , \zin[1][63] , \zin[1][62] , \zin[1][61] , 
        \zin[1][60] , \zin[1][59] , \zin[1][58] , \zin[1][57] , \zin[1][56] , 
        \zin[1][55] , \zin[1][54] , \zin[1][53] , \zin[1][52] , \zin[1][51] , 
        \zin[1][50] , \zin[1][49] , \zin[1][48] , \zin[1][47] , \zin[1][46] , 
        \zin[1][45] , \zin[1][44] , \zin[1][43] , \zin[1][42] , \zin[1][41] , 
        \zin[1][40] , \zin[1][39] , \zin[1][38] , \zin[1][37] , \zin[1][36] , 
        \zin[1][35] , \zin[1][34] , \zin[1][33] , \zin[1][32] , \zin[1][31] , 
        \zin[1][30] , \zin[1][29] , \zin[1][28] , \zin[1][27] , \zin[1][26] , 
        \zin[1][25] , \zin[1][24] , \zin[1][23] , \zin[1][22] , \zin[1][21] , 
        \zin[1][20] , \zin[1][19] , \zin[1][18] , \zin[1][17] , \zin[1][16] , 
        \zin[1][15] , \zin[1][14] , \zin[1][13] , \zin[1][12] , \zin[1][11] , 
        \zin[1][10] , \zin[1][9] , \zin[1][8] , \zin[1][7] , \zin[1][6] , 
        \zin[1][5] , \zin[1][4] , \zin[1][3] , \zin[1][2] , \zin[1][1] , 
        \zin[1][0] }) );
  modmult_step_N256_1_1 \MODMULT_STEP[1].modmult_step_  ( .xregN_1(xin[254]), 
        .y(y), .n(n), .zin({1'b0, \zin[1][256] , \zin[1][255] , \zin[1][254] , 
        \zin[1][253] , \zin[1][252] , \zin[1][251] , \zin[1][250] , 
        \zin[1][249] , \zin[1][248] , \zin[1][247] , \zin[1][246] , 
        \zin[1][245] , \zin[1][244] , \zin[1][243] , \zin[1][242] , 
        \zin[1][241] , \zin[1][240] , \zin[1][239] , \zin[1][238] , 
        \zin[1][237] , \zin[1][236] , \zin[1][235] , \zin[1][234] , 
        \zin[1][233] , \zin[1][232] , \zin[1][231] , \zin[1][230] , 
        \zin[1][229] , \zin[1][228] , \zin[1][227] , \zin[1][226] , 
        \zin[1][225] , \zin[1][224] , \zin[1][223] , \zin[1][222] , 
        \zin[1][221] , \zin[1][220] , \zin[1][219] , \zin[1][218] , 
        \zin[1][217] , \zin[1][216] , \zin[1][215] , \zin[1][214] , 
        \zin[1][213] , \zin[1][212] , \zin[1][211] , \zin[1][210] , 
        \zin[1][209] , \zin[1][208] , \zin[1][207] , \zin[1][206] , 
        \zin[1][205] , \zin[1][204] , \zin[1][203] , \zin[1][202] , 
        \zin[1][201] , \zin[1][200] , \zin[1][199] , \zin[1][198] , 
        \zin[1][197] , \zin[1][196] , \zin[1][195] , \zin[1][194] , 
        \zin[1][193] , \zin[1][192] , \zin[1][191] , \zin[1][190] , 
        \zin[1][189] , \zin[1][188] , \zin[1][187] , \zin[1][186] , 
        \zin[1][185] , \zin[1][184] , \zin[1][183] , \zin[1][182] , 
        \zin[1][181] , \zin[1][180] , \zin[1][179] , \zin[1][178] , 
        \zin[1][177] , \zin[1][176] , \zin[1][175] , \zin[1][174] , 
        \zin[1][173] , \zin[1][172] , \zin[1][171] , \zin[1][170] , 
        \zin[1][169] , \zin[1][168] , \zin[1][167] , \zin[1][166] , 
        \zin[1][165] , \zin[1][164] , \zin[1][163] , \zin[1][162] , 
        \zin[1][161] , \zin[1][160] , \zin[1][159] , \zin[1][158] , 
        \zin[1][157] , \zin[1][156] , \zin[1][155] , \zin[1][154] , 
        \zin[1][153] , \zin[1][152] , \zin[1][151] , \zin[1][150] , 
        \zin[1][149] , \zin[1][148] , \zin[1][147] , \zin[1][146] , 
        \zin[1][145] , \zin[1][144] , \zin[1][143] , \zin[1][142] , 
        \zin[1][141] , \zin[1][140] , \zin[1][139] , \zin[1][138] , 
        \zin[1][137] , \zin[1][136] , \zin[1][135] , \zin[1][134] , 
        \zin[1][133] , \zin[1][132] , \zin[1][131] , \zin[1][130] , 
        \zin[1][129] , \zin[1][128] , \zin[1][127] , \zin[1][126] , 
        \zin[1][125] , \zin[1][124] , \zin[1][123] , \zin[1][122] , 
        \zin[1][121] , \zin[1][120] , \zin[1][119] , \zin[1][118] , 
        \zin[1][117] , \zin[1][116] , \zin[1][115] , \zin[1][114] , 
        \zin[1][113] , \zin[1][112] , \zin[1][111] , \zin[1][110] , 
        \zin[1][109] , \zin[1][108] , \zin[1][107] , \zin[1][106] , 
        \zin[1][105] , \zin[1][104] , \zin[1][103] , \zin[1][102] , 
        \zin[1][101] , \zin[1][100] , \zin[1][99] , \zin[1][98] , \zin[1][97] , 
        \zin[1][96] , \zin[1][95] , \zin[1][94] , \zin[1][93] , \zin[1][92] , 
        \zin[1][91] , \zin[1][90] , \zin[1][89] , \zin[1][88] , \zin[1][87] , 
        \zin[1][86] , \zin[1][85] , \zin[1][84] , \zin[1][83] , \zin[1][82] , 
        \zin[1][81] , \zin[1][80] , \zin[1][79] , \zin[1][78] , \zin[1][77] , 
        \zin[1][76] , \zin[1][75] , \zin[1][74] , \zin[1][73] , \zin[1][72] , 
        \zin[1][71] , \zin[1][70] , \zin[1][69] , \zin[1][68] , \zin[1][67] , 
        \zin[1][66] , \zin[1][65] , \zin[1][64] , \zin[1][63] , \zin[1][62] , 
        \zin[1][61] , \zin[1][60] , \zin[1][59] , \zin[1][58] , \zin[1][57] , 
        \zin[1][56] , \zin[1][55] , \zin[1][54] , \zin[1][53] , \zin[1][52] , 
        \zin[1][51] , \zin[1][50] , \zin[1][49] , \zin[1][48] , \zin[1][47] , 
        \zin[1][46] , \zin[1][45] , \zin[1][44] , \zin[1][43] , \zin[1][42] , 
        \zin[1][41] , \zin[1][40] , \zin[1][39] , \zin[1][38] , \zin[1][37] , 
        \zin[1][36] , \zin[1][35] , \zin[1][34] , \zin[1][33] , \zin[1][32] , 
        \zin[1][31] , \zin[1][30] , \zin[1][29] , \zin[1][28] , \zin[1][27] , 
        \zin[1][26] , \zin[1][25] , \zin[1][24] , \zin[1][23] , \zin[1][22] , 
        \zin[1][21] , \zin[1][20] , \zin[1][19] , \zin[1][18] , \zin[1][17] , 
        \zin[1][16] , \zin[1][15] , \zin[1][14] , \zin[1][13] , \zin[1][12] , 
        \zin[1][11] , \zin[1][10] , \zin[1][9] , \zin[1][8] , \zin[1][7] , 
        \zin[1][6] , \zin[1][5] , \zin[1][4] , \zin[1][3] , \zin[1][2] , 
        \zin[1][1] , \zin[1][0] }), .zout({SYNOPSYS_UNCONNECTED__1, 
        \zout[1][256] , o}) );
  DFF \xreg_reg[1]  ( .D(1'b0), .CLK(clk), .RST(start), .I(x[1]), .Q(xin[1])
         );
  DFF \xreg_reg[3]  ( .D(xin[1]), .CLK(clk), .RST(start), .I(x[3]), .Q(xin[3])
         );
  DFF \xreg_reg[5]  ( .D(xin[3]), .CLK(clk), .RST(start), .I(x[5]), .Q(xin[5])
         );
  DFF \xreg_reg[7]  ( .D(xin[5]), .CLK(clk), .RST(start), .I(x[7]), .Q(xin[7])
         );
  DFF \xreg_reg[9]  ( .D(xin[7]), .CLK(clk), .RST(start), .I(x[9]), .Q(xin[9])
         );
  DFF \xreg_reg[11]  ( .D(xin[9]), .CLK(clk), .RST(start), .I(x[11]), .Q(
        xin[11]) );
  DFF \xreg_reg[13]  ( .D(xin[11]), .CLK(clk), .RST(start), .I(x[13]), .Q(
        xin[13]) );
  DFF \xreg_reg[15]  ( .D(xin[13]), .CLK(clk), .RST(start), .I(x[15]), .Q(
        xin[15]) );
  DFF \xreg_reg[17]  ( .D(xin[15]), .CLK(clk), .RST(start), .I(x[17]), .Q(
        xin[17]) );
  DFF \xreg_reg[19]  ( .D(xin[17]), .CLK(clk), .RST(start), .I(x[19]), .Q(
        xin[19]) );
  DFF \xreg_reg[21]  ( .D(xin[19]), .CLK(clk), .RST(start), .I(x[21]), .Q(
        xin[21]) );
  DFF \xreg_reg[23]  ( .D(xin[21]), .CLK(clk), .RST(start), .I(x[23]), .Q(
        xin[23]) );
  DFF \xreg_reg[25]  ( .D(xin[23]), .CLK(clk), .RST(start), .I(x[25]), .Q(
        xin[25]) );
  DFF \xreg_reg[27]  ( .D(xin[25]), .CLK(clk), .RST(start), .I(x[27]), .Q(
        xin[27]) );
  DFF \xreg_reg[29]  ( .D(xin[27]), .CLK(clk), .RST(start), .I(x[29]), .Q(
        xin[29]) );
  DFF \xreg_reg[31]  ( .D(xin[29]), .CLK(clk), .RST(start), .I(x[31]), .Q(
        xin[31]) );
  DFF \xreg_reg[33]  ( .D(xin[31]), .CLK(clk), .RST(start), .I(x[33]), .Q(
        xin[33]) );
  DFF \xreg_reg[35]  ( .D(xin[33]), .CLK(clk), .RST(start), .I(x[35]), .Q(
        xin[35]) );
  DFF \xreg_reg[37]  ( .D(xin[35]), .CLK(clk), .RST(start), .I(x[37]), .Q(
        xin[37]) );
  DFF \xreg_reg[39]  ( .D(xin[37]), .CLK(clk), .RST(start), .I(x[39]), .Q(
        xin[39]) );
  DFF \xreg_reg[41]  ( .D(xin[39]), .CLK(clk), .RST(start), .I(x[41]), .Q(
        xin[41]) );
  DFF \xreg_reg[43]  ( .D(xin[41]), .CLK(clk), .RST(start), .I(x[43]), .Q(
        xin[43]) );
  DFF \xreg_reg[45]  ( .D(xin[43]), .CLK(clk), .RST(start), .I(x[45]), .Q(
        xin[45]) );
  DFF \xreg_reg[47]  ( .D(xin[45]), .CLK(clk), .RST(start), .I(x[47]), .Q(
        xin[47]) );
  DFF \xreg_reg[49]  ( .D(xin[47]), .CLK(clk), .RST(start), .I(x[49]), .Q(
        xin[49]) );
  DFF \xreg_reg[51]  ( .D(xin[49]), .CLK(clk), .RST(start), .I(x[51]), .Q(
        xin[51]) );
  DFF \xreg_reg[53]  ( .D(xin[51]), .CLK(clk), .RST(start), .I(x[53]), .Q(
        xin[53]) );
  DFF \xreg_reg[55]  ( .D(xin[53]), .CLK(clk), .RST(start), .I(x[55]), .Q(
        xin[55]) );
  DFF \xreg_reg[57]  ( .D(xin[55]), .CLK(clk), .RST(start), .I(x[57]), .Q(
        xin[57]) );
  DFF \xreg_reg[59]  ( .D(xin[57]), .CLK(clk), .RST(start), .I(x[59]), .Q(
        xin[59]) );
  DFF \xreg_reg[61]  ( .D(xin[59]), .CLK(clk), .RST(start), .I(x[61]), .Q(
        xin[61]) );
  DFF \xreg_reg[63]  ( .D(xin[61]), .CLK(clk), .RST(start), .I(x[63]), .Q(
        xin[63]) );
  DFF \xreg_reg[65]  ( .D(xin[63]), .CLK(clk), .RST(start), .I(x[65]), .Q(
        xin[65]) );
  DFF \xreg_reg[67]  ( .D(xin[65]), .CLK(clk), .RST(start), .I(x[67]), .Q(
        xin[67]) );
  DFF \xreg_reg[69]  ( .D(xin[67]), .CLK(clk), .RST(start), .I(x[69]), .Q(
        xin[69]) );
  DFF \xreg_reg[71]  ( .D(xin[69]), .CLK(clk), .RST(start), .I(x[71]), .Q(
        xin[71]) );
  DFF \xreg_reg[73]  ( .D(xin[71]), .CLK(clk), .RST(start), .I(x[73]), .Q(
        xin[73]) );
  DFF \xreg_reg[75]  ( .D(xin[73]), .CLK(clk), .RST(start), .I(x[75]), .Q(
        xin[75]) );
  DFF \xreg_reg[77]  ( .D(xin[75]), .CLK(clk), .RST(start), .I(x[77]), .Q(
        xin[77]) );
  DFF \xreg_reg[79]  ( .D(xin[77]), .CLK(clk), .RST(start), .I(x[79]), .Q(
        xin[79]) );
  DFF \xreg_reg[81]  ( .D(xin[79]), .CLK(clk), .RST(start), .I(x[81]), .Q(
        xin[81]) );
  DFF \xreg_reg[83]  ( .D(xin[81]), .CLK(clk), .RST(start), .I(x[83]), .Q(
        xin[83]) );
  DFF \xreg_reg[85]  ( .D(xin[83]), .CLK(clk), .RST(start), .I(x[85]), .Q(
        xin[85]) );
  DFF \xreg_reg[87]  ( .D(xin[85]), .CLK(clk), .RST(start), .I(x[87]), .Q(
        xin[87]) );
  DFF \xreg_reg[89]  ( .D(xin[87]), .CLK(clk), .RST(start), .I(x[89]), .Q(
        xin[89]) );
  DFF \xreg_reg[91]  ( .D(xin[89]), .CLK(clk), .RST(start), .I(x[91]), .Q(
        xin[91]) );
  DFF \xreg_reg[93]  ( .D(xin[91]), .CLK(clk), .RST(start), .I(x[93]), .Q(
        xin[93]) );
  DFF \xreg_reg[95]  ( .D(xin[93]), .CLK(clk), .RST(start), .I(x[95]), .Q(
        xin[95]) );
  DFF \xreg_reg[97]  ( .D(xin[95]), .CLK(clk), .RST(start), .I(x[97]), .Q(
        xin[97]) );
  DFF \xreg_reg[99]  ( .D(xin[97]), .CLK(clk), .RST(start), .I(x[99]), .Q(
        xin[99]) );
  DFF \xreg_reg[101]  ( .D(xin[99]), .CLK(clk), .RST(start), .I(x[101]), .Q(
        xin[101]) );
  DFF \xreg_reg[103]  ( .D(xin[101]), .CLK(clk), .RST(start), .I(x[103]), .Q(
        xin[103]) );
  DFF \xreg_reg[105]  ( .D(xin[103]), .CLK(clk), .RST(start), .I(x[105]), .Q(
        xin[105]) );
  DFF \xreg_reg[107]  ( .D(xin[105]), .CLK(clk), .RST(start), .I(x[107]), .Q(
        xin[107]) );
  DFF \xreg_reg[109]  ( .D(xin[107]), .CLK(clk), .RST(start), .I(x[109]), .Q(
        xin[109]) );
  DFF \xreg_reg[111]  ( .D(xin[109]), .CLK(clk), .RST(start), .I(x[111]), .Q(
        xin[111]) );
  DFF \xreg_reg[113]  ( .D(xin[111]), .CLK(clk), .RST(start), .I(x[113]), .Q(
        xin[113]) );
  DFF \xreg_reg[115]  ( .D(xin[113]), .CLK(clk), .RST(start), .I(x[115]), .Q(
        xin[115]) );
  DFF \xreg_reg[117]  ( .D(xin[115]), .CLK(clk), .RST(start), .I(x[117]), .Q(
        xin[117]) );
  DFF \xreg_reg[119]  ( .D(xin[117]), .CLK(clk), .RST(start), .I(x[119]), .Q(
        xin[119]) );
  DFF \xreg_reg[121]  ( .D(xin[119]), .CLK(clk), .RST(start), .I(x[121]), .Q(
        xin[121]) );
  DFF \xreg_reg[123]  ( .D(xin[121]), .CLK(clk), .RST(start), .I(x[123]), .Q(
        xin[123]) );
  DFF \xreg_reg[125]  ( .D(xin[123]), .CLK(clk), .RST(start), .I(x[125]), .Q(
        xin[125]) );
  DFF \xreg_reg[127]  ( .D(xin[125]), .CLK(clk), .RST(start), .I(x[127]), .Q(
        xin[127]) );
  DFF \xreg_reg[129]  ( .D(xin[127]), .CLK(clk), .RST(start), .I(x[129]), .Q(
        xin[129]) );
  DFF \xreg_reg[131]  ( .D(xin[129]), .CLK(clk), .RST(start), .I(x[131]), .Q(
        xin[131]) );
  DFF \xreg_reg[133]  ( .D(xin[131]), .CLK(clk), .RST(start), .I(x[133]), .Q(
        xin[133]) );
  DFF \xreg_reg[135]  ( .D(xin[133]), .CLK(clk), .RST(start), .I(x[135]), .Q(
        xin[135]) );
  DFF \xreg_reg[137]  ( .D(xin[135]), .CLK(clk), .RST(start), .I(x[137]), .Q(
        xin[137]) );
  DFF \xreg_reg[139]  ( .D(xin[137]), .CLK(clk), .RST(start), .I(x[139]), .Q(
        xin[139]) );
  DFF \xreg_reg[141]  ( .D(xin[139]), .CLK(clk), .RST(start), .I(x[141]), .Q(
        xin[141]) );
  DFF \xreg_reg[143]  ( .D(xin[141]), .CLK(clk), .RST(start), .I(x[143]), .Q(
        xin[143]) );
  DFF \xreg_reg[145]  ( .D(xin[143]), .CLK(clk), .RST(start), .I(x[145]), .Q(
        xin[145]) );
  DFF \xreg_reg[147]  ( .D(xin[145]), .CLK(clk), .RST(start), .I(x[147]), .Q(
        xin[147]) );
  DFF \xreg_reg[149]  ( .D(xin[147]), .CLK(clk), .RST(start), .I(x[149]), .Q(
        xin[149]) );
  DFF \xreg_reg[151]  ( .D(xin[149]), .CLK(clk), .RST(start), .I(x[151]), .Q(
        xin[151]) );
  DFF \xreg_reg[153]  ( .D(xin[151]), .CLK(clk), .RST(start), .I(x[153]), .Q(
        xin[153]) );
  DFF \xreg_reg[155]  ( .D(xin[153]), .CLK(clk), .RST(start), .I(x[155]), .Q(
        xin[155]) );
  DFF \xreg_reg[157]  ( .D(xin[155]), .CLK(clk), .RST(start), .I(x[157]), .Q(
        xin[157]) );
  DFF \xreg_reg[159]  ( .D(xin[157]), .CLK(clk), .RST(start), .I(x[159]), .Q(
        xin[159]) );
  DFF \xreg_reg[161]  ( .D(xin[159]), .CLK(clk), .RST(start), .I(x[161]), .Q(
        xin[161]) );
  DFF \xreg_reg[163]  ( .D(xin[161]), .CLK(clk), .RST(start), .I(x[163]), .Q(
        xin[163]) );
  DFF \xreg_reg[165]  ( .D(xin[163]), .CLK(clk), .RST(start), .I(x[165]), .Q(
        xin[165]) );
  DFF \xreg_reg[167]  ( .D(xin[165]), .CLK(clk), .RST(start), .I(x[167]), .Q(
        xin[167]) );
  DFF \xreg_reg[169]  ( .D(xin[167]), .CLK(clk), .RST(start), .I(x[169]), .Q(
        xin[169]) );
  DFF \xreg_reg[171]  ( .D(xin[169]), .CLK(clk), .RST(start), .I(x[171]), .Q(
        xin[171]) );
  DFF \xreg_reg[173]  ( .D(xin[171]), .CLK(clk), .RST(start), .I(x[173]), .Q(
        xin[173]) );
  DFF \xreg_reg[175]  ( .D(xin[173]), .CLK(clk), .RST(start), .I(x[175]), .Q(
        xin[175]) );
  DFF \xreg_reg[177]  ( .D(xin[175]), .CLK(clk), .RST(start), .I(x[177]), .Q(
        xin[177]) );
  DFF \xreg_reg[179]  ( .D(xin[177]), .CLK(clk), .RST(start), .I(x[179]), .Q(
        xin[179]) );
  DFF \xreg_reg[181]  ( .D(xin[179]), .CLK(clk), .RST(start), .I(x[181]), .Q(
        xin[181]) );
  DFF \xreg_reg[183]  ( .D(xin[181]), .CLK(clk), .RST(start), .I(x[183]), .Q(
        xin[183]) );
  DFF \xreg_reg[185]  ( .D(xin[183]), .CLK(clk), .RST(start), .I(x[185]), .Q(
        xin[185]) );
  DFF \xreg_reg[187]  ( .D(xin[185]), .CLK(clk), .RST(start), .I(x[187]), .Q(
        xin[187]) );
  DFF \xreg_reg[189]  ( .D(xin[187]), .CLK(clk), .RST(start), .I(x[189]), .Q(
        xin[189]) );
  DFF \xreg_reg[191]  ( .D(xin[189]), .CLK(clk), .RST(start), .I(x[191]), .Q(
        xin[191]) );
  DFF \xreg_reg[193]  ( .D(xin[191]), .CLK(clk), .RST(start), .I(x[193]), .Q(
        xin[193]) );
  DFF \xreg_reg[195]  ( .D(xin[193]), .CLK(clk), .RST(start), .I(x[195]), .Q(
        xin[195]) );
  DFF \xreg_reg[197]  ( .D(xin[195]), .CLK(clk), .RST(start), .I(x[197]), .Q(
        xin[197]) );
  DFF \xreg_reg[199]  ( .D(xin[197]), .CLK(clk), .RST(start), .I(x[199]), .Q(
        xin[199]) );
  DFF \xreg_reg[201]  ( .D(xin[199]), .CLK(clk), .RST(start), .I(x[201]), .Q(
        xin[201]) );
  DFF \xreg_reg[203]  ( .D(xin[201]), .CLK(clk), .RST(start), .I(x[203]), .Q(
        xin[203]) );
  DFF \xreg_reg[205]  ( .D(xin[203]), .CLK(clk), .RST(start), .I(x[205]), .Q(
        xin[205]) );
  DFF \xreg_reg[207]  ( .D(xin[205]), .CLK(clk), .RST(start), .I(x[207]), .Q(
        xin[207]) );
  DFF \xreg_reg[209]  ( .D(xin[207]), .CLK(clk), .RST(start), .I(x[209]), .Q(
        xin[209]) );
  DFF \xreg_reg[211]  ( .D(xin[209]), .CLK(clk), .RST(start), .I(x[211]), .Q(
        xin[211]) );
  DFF \xreg_reg[213]  ( .D(xin[211]), .CLK(clk), .RST(start), .I(x[213]), .Q(
        xin[213]) );
  DFF \xreg_reg[215]  ( .D(xin[213]), .CLK(clk), .RST(start), .I(x[215]), .Q(
        xin[215]) );
  DFF \xreg_reg[217]  ( .D(xin[215]), .CLK(clk), .RST(start), .I(x[217]), .Q(
        xin[217]) );
  DFF \xreg_reg[219]  ( .D(xin[217]), .CLK(clk), .RST(start), .I(x[219]), .Q(
        xin[219]) );
  DFF \xreg_reg[221]  ( .D(xin[219]), .CLK(clk), .RST(start), .I(x[221]), .Q(
        xin[221]) );
  DFF \xreg_reg[223]  ( .D(xin[221]), .CLK(clk), .RST(start), .I(x[223]), .Q(
        xin[223]) );
  DFF \xreg_reg[225]  ( .D(xin[223]), .CLK(clk), .RST(start), .I(x[225]), .Q(
        xin[225]) );
  DFF \xreg_reg[227]  ( .D(xin[225]), .CLK(clk), .RST(start), .I(x[227]), .Q(
        xin[227]) );
  DFF \xreg_reg[229]  ( .D(xin[227]), .CLK(clk), .RST(start), .I(x[229]), .Q(
        xin[229]) );
  DFF \xreg_reg[231]  ( .D(xin[229]), .CLK(clk), .RST(start), .I(x[231]), .Q(
        xin[231]) );
  DFF \xreg_reg[233]  ( .D(xin[231]), .CLK(clk), .RST(start), .I(x[233]), .Q(
        xin[233]) );
  DFF \xreg_reg[235]  ( .D(xin[233]), .CLK(clk), .RST(start), .I(x[235]), .Q(
        xin[235]) );
  DFF \xreg_reg[237]  ( .D(xin[235]), .CLK(clk), .RST(start), .I(x[237]), .Q(
        xin[237]) );
  DFF \xreg_reg[239]  ( .D(xin[237]), .CLK(clk), .RST(start), .I(x[239]), .Q(
        xin[239]) );
  DFF \xreg_reg[241]  ( .D(xin[239]), .CLK(clk), .RST(start), .I(x[241]), .Q(
        xin[241]) );
  DFF \xreg_reg[243]  ( .D(xin[241]), .CLK(clk), .RST(start), .I(x[243]), .Q(
        xin[243]) );
  DFF \xreg_reg[245]  ( .D(xin[243]), .CLK(clk), .RST(start), .I(x[245]), .Q(
        xin[245]) );
  DFF \xreg_reg[247]  ( .D(xin[245]), .CLK(clk), .RST(start), .I(x[247]), .Q(
        xin[247]) );
  DFF \xreg_reg[249]  ( .D(xin[247]), .CLK(clk), .RST(start), .I(x[249]), .Q(
        xin[249]) );
  DFF \xreg_reg[251]  ( .D(xin[249]), .CLK(clk), .RST(start), .I(x[251]), .Q(
        xin[251]) );
  DFF \xreg_reg[253]  ( .D(xin[251]), .CLK(clk), .RST(start), .I(x[253]), .Q(
        xin[253]) );
  DFF \xreg_reg[255]  ( .D(xin[253]), .CLK(clk), .RST(start), .I(x[255]), .Q(
        xin[255]) );
  DFF \xreg_reg[0]  ( .D(1'b0), .CLK(clk), .RST(start), .I(x[0]), .Q(xin[0])
         );
  DFF \xreg_reg[2]  ( .D(xin[0]), .CLK(clk), .RST(start), .I(x[2]), .Q(xin[2])
         );
  DFF \xreg_reg[4]  ( .D(xin[2]), .CLK(clk), .RST(start), .I(x[4]), .Q(xin[4])
         );
  DFF \xreg_reg[6]  ( .D(xin[4]), .CLK(clk), .RST(start), .I(x[6]), .Q(xin[6])
         );
  DFF \xreg_reg[8]  ( .D(xin[6]), .CLK(clk), .RST(start), .I(x[8]), .Q(xin[8])
         );
  DFF \xreg_reg[10]  ( .D(xin[8]), .CLK(clk), .RST(start), .I(x[10]), .Q(
        xin[10]) );
  DFF \xreg_reg[12]  ( .D(xin[10]), .CLK(clk), .RST(start), .I(x[12]), .Q(
        xin[12]) );
  DFF \xreg_reg[14]  ( .D(xin[12]), .CLK(clk), .RST(start), .I(x[14]), .Q(
        xin[14]) );
  DFF \xreg_reg[16]  ( .D(xin[14]), .CLK(clk), .RST(start), .I(x[16]), .Q(
        xin[16]) );
  DFF \xreg_reg[18]  ( .D(xin[16]), .CLK(clk), .RST(start), .I(x[18]), .Q(
        xin[18]) );
  DFF \xreg_reg[20]  ( .D(xin[18]), .CLK(clk), .RST(start), .I(x[20]), .Q(
        xin[20]) );
  DFF \xreg_reg[22]  ( .D(xin[20]), .CLK(clk), .RST(start), .I(x[22]), .Q(
        xin[22]) );
  DFF \xreg_reg[24]  ( .D(xin[22]), .CLK(clk), .RST(start), .I(x[24]), .Q(
        xin[24]) );
  DFF \xreg_reg[26]  ( .D(xin[24]), .CLK(clk), .RST(start), .I(x[26]), .Q(
        xin[26]) );
  DFF \xreg_reg[28]  ( .D(xin[26]), .CLK(clk), .RST(start), .I(x[28]), .Q(
        xin[28]) );
  DFF \xreg_reg[30]  ( .D(xin[28]), .CLK(clk), .RST(start), .I(x[30]), .Q(
        xin[30]) );
  DFF \xreg_reg[32]  ( .D(xin[30]), .CLK(clk), .RST(start), .I(x[32]), .Q(
        xin[32]) );
  DFF \xreg_reg[34]  ( .D(xin[32]), .CLK(clk), .RST(start), .I(x[34]), .Q(
        xin[34]) );
  DFF \xreg_reg[36]  ( .D(xin[34]), .CLK(clk), .RST(start), .I(x[36]), .Q(
        xin[36]) );
  DFF \xreg_reg[38]  ( .D(xin[36]), .CLK(clk), .RST(start), .I(x[38]), .Q(
        xin[38]) );
  DFF \xreg_reg[40]  ( .D(xin[38]), .CLK(clk), .RST(start), .I(x[40]), .Q(
        xin[40]) );
  DFF \xreg_reg[42]  ( .D(xin[40]), .CLK(clk), .RST(start), .I(x[42]), .Q(
        xin[42]) );
  DFF \xreg_reg[44]  ( .D(xin[42]), .CLK(clk), .RST(start), .I(x[44]), .Q(
        xin[44]) );
  DFF \xreg_reg[46]  ( .D(xin[44]), .CLK(clk), .RST(start), .I(x[46]), .Q(
        xin[46]) );
  DFF \xreg_reg[48]  ( .D(xin[46]), .CLK(clk), .RST(start), .I(x[48]), .Q(
        xin[48]) );
  DFF \xreg_reg[50]  ( .D(xin[48]), .CLK(clk), .RST(start), .I(x[50]), .Q(
        xin[50]) );
  DFF \xreg_reg[52]  ( .D(xin[50]), .CLK(clk), .RST(start), .I(x[52]), .Q(
        xin[52]) );
  DFF \xreg_reg[54]  ( .D(xin[52]), .CLK(clk), .RST(start), .I(x[54]), .Q(
        xin[54]) );
  DFF \xreg_reg[56]  ( .D(xin[54]), .CLK(clk), .RST(start), .I(x[56]), .Q(
        xin[56]) );
  DFF \xreg_reg[58]  ( .D(xin[56]), .CLK(clk), .RST(start), .I(x[58]), .Q(
        xin[58]) );
  DFF \xreg_reg[60]  ( .D(xin[58]), .CLK(clk), .RST(start), .I(x[60]), .Q(
        xin[60]) );
  DFF \xreg_reg[62]  ( .D(xin[60]), .CLK(clk), .RST(start), .I(x[62]), .Q(
        xin[62]) );
  DFF \xreg_reg[64]  ( .D(xin[62]), .CLK(clk), .RST(start), .I(x[64]), .Q(
        xin[64]) );
  DFF \xreg_reg[66]  ( .D(xin[64]), .CLK(clk), .RST(start), .I(x[66]), .Q(
        xin[66]) );
  DFF \xreg_reg[68]  ( .D(xin[66]), .CLK(clk), .RST(start), .I(x[68]), .Q(
        xin[68]) );
  DFF \xreg_reg[70]  ( .D(xin[68]), .CLK(clk), .RST(start), .I(x[70]), .Q(
        xin[70]) );
  DFF \xreg_reg[72]  ( .D(xin[70]), .CLK(clk), .RST(start), .I(x[72]), .Q(
        xin[72]) );
  DFF \xreg_reg[74]  ( .D(xin[72]), .CLK(clk), .RST(start), .I(x[74]), .Q(
        xin[74]) );
  DFF \xreg_reg[76]  ( .D(xin[74]), .CLK(clk), .RST(start), .I(x[76]), .Q(
        xin[76]) );
  DFF \xreg_reg[78]  ( .D(xin[76]), .CLK(clk), .RST(start), .I(x[78]), .Q(
        xin[78]) );
  DFF \xreg_reg[80]  ( .D(xin[78]), .CLK(clk), .RST(start), .I(x[80]), .Q(
        xin[80]) );
  DFF \xreg_reg[82]  ( .D(xin[80]), .CLK(clk), .RST(start), .I(x[82]), .Q(
        xin[82]) );
  DFF \xreg_reg[84]  ( .D(xin[82]), .CLK(clk), .RST(start), .I(x[84]), .Q(
        xin[84]) );
  DFF \xreg_reg[86]  ( .D(xin[84]), .CLK(clk), .RST(start), .I(x[86]), .Q(
        xin[86]) );
  DFF \xreg_reg[88]  ( .D(xin[86]), .CLK(clk), .RST(start), .I(x[88]), .Q(
        xin[88]) );
  DFF \xreg_reg[90]  ( .D(xin[88]), .CLK(clk), .RST(start), .I(x[90]), .Q(
        xin[90]) );
  DFF \xreg_reg[92]  ( .D(xin[90]), .CLK(clk), .RST(start), .I(x[92]), .Q(
        xin[92]) );
  DFF \xreg_reg[94]  ( .D(xin[92]), .CLK(clk), .RST(start), .I(x[94]), .Q(
        xin[94]) );
  DFF \xreg_reg[96]  ( .D(xin[94]), .CLK(clk), .RST(start), .I(x[96]), .Q(
        xin[96]) );
  DFF \xreg_reg[98]  ( .D(xin[96]), .CLK(clk), .RST(start), .I(x[98]), .Q(
        xin[98]) );
  DFF \xreg_reg[100]  ( .D(xin[98]), .CLK(clk), .RST(start), .I(x[100]), .Q(
        xin[100]) );
  DFF \xreg_reg[102]  ( .D(xin[100]), .CLK(clk), .RST(start), .I(x[102]), .Q(
        xin[102]) );
  DFF \xreg_reg[104]  ( .D(xin[102]), .CLK(clk), .RST(start), .I(x[104]), .Q(
        xin[104]) );
  DFF \xreg_reg[106]  ( .D(xin[104]), .CLK(clk), .RST(start), .I(x[106]), .Q(
        xin[106]) );
  DFF \xreg_reg[108]  ( .D(xin[106]), .CLK(clk), .RST(start), .I(x[108]), .Q(
        xin[108]) );
  DFF \xreg_reg[110]  ( .D(xin[108]), .CLK(clk), .RST(start), .I(x[110]), .Q(
        xin[110]) );
  DFF \xreg_reg[112]  ( .D(xin[110]), .CLK(clk), .RST(start), .I(x[112]), .Q(
        xin[112]) );
  DFF \xreg_reg[114]  ( .D(xin[112]), .CLK(clk), .RST(start), .I(x[114]), .Q(
        xin[114]) );
  DFF \xreg_reg[116]  ( .D(xin[114]), .CLK(clk), .RST(start), .I(x[116]), .Q(
        xin[116]) );
  DFF \xreg_reg[118]  ( .D(xin[116]), .CLK(clk), .RST(start), .I(x[118]), .Q(
        xin[118]) );
  DFF \xreg_reg[120]  ( .D(xin[118]), .CLK(clk), .RST(start), .I(x[120]), .Q(
        xin[120]) );
  DFF \xreg_reg[122]  ( .D(xin[120]), .CLK(clk), .RST(start), .I(x[122]), .Q(
        xin[122]) );
  DFF \xreg_reg[124]  ( .D(xin[122]), .CLK(clk), .RST(start), .I(x[124]), .Q(
        xin[124]) );
  DFF \xreg_reg[126]  ( .D(xin[124]), .CLK(clk), .RST(start), .I(x[126]), .Q(
        xin[126]) );
  DFF \xreg_reg[128]  ( .D(xin[126]), .CLK(clk), .RST(start), .I(x[128]), .Q(
        xin[128]) );
  DFF \xreg_reg[130]  ( .D(xin[128]), .CLK(clk), .RST(start), .I(x[130]), .Q(
        xin[130]) );
  DFF \xreg_reg[132]  ( .D(xin[130]), .CLK(clk), .RST(start), .I(x[132]), .Q(
        xin[132]) );
  DFF \xreg_reg[134]  ( .D(xin[132]), .CLK(clk), .RST(start), .I(x[134]), .Q(
        xin[134]) );
  DFF \xreg_reg[136]  ( .D(xin[134]), .CLK(clk), .RST(start), .I(x[136]), .Q(
        xin[136]) );
  DFF \xreg_reg[138]  ( .D(xin[136]), .CLK(clk), .RST(start), .I(x[138]), .Q(
        xin[138]) );
  DFF \xreg_reg[140]  ( .D(xin[138]), .CLK(clk), .RST(start), .I(x[140]), .Q(
        xin[140]) );
  DFF \xreg_reg[142]  ( .D(xin[140]), .CLK(clk), .RST(start), .I(x[142]), .Q(
        xin[142]) );
  DFF \xreg_reg[144]  ( .D(xin[142]), .CLK(clk), .RST(start), .I(x[144]), .Q(
        xin[144]) );
  DFF \xreg_reg[146]  ( .D(xin[144]), .CLK(clk), .RST(start), .I(x[146]), .Q(
        xin[146]) );
  DFF \xreg_reg[148]  ( .D(xin[146]), .CLK(clk), .RST(start), .I(x[148]), .Q(
        xin[148]) );
  DFF \xreg_reg[150]  ( .D(xin[148]), .CLK(clk), .RST(start), .I(x[150]), .Q(
        xin[150]) );
  DFF \xreg_reg[152]  ( .D(xin[150]), .CLK(clk), .RST(start), .I(x[152]), .Q(
        xin[152]) );
  DFF \xreg_reg[154]  ( .D(xin[152]), .CLK(clk), .RST(start), .I(x[154]), .Q(
        xin[154]) );
  DFF \xreg_reg[156]  ( .D(xin[154]), .CLK(clk), .RST(start), .I(x[156]), .Q(
        xin[156]) );
  DFF \xreg_reg[158]  ( .D(xin[156]), .CLK(clk), .RST(start), .I(x[158]), .Q(
        xin[158]) );
  DFF \xreg_reg[160]  ( .D(xin[158]), .CLK(clk), .RST(start), .I(x[160]), .Q(
        xin[160]) );
  DFF \xreg_reg[162]  ( .D(xin[160]), .CLK(clk), .RST(start), .I(x[162]), .Q(
        xin[162]) );
  DFF \xreg_reg[164]  ( .D(xin[162]), .CLK(clk), .RST(start), .I(x[164]), .Q(
        xin[164]) );
  DFF \xreg_reg[166]  ( .D(xin[164]), .CLK(clk), .RST(start), .I(x[166]), .Q(
        xin[166]) );
  DFF \xreg_reg[168]  ( .D(xin[166]), .CLK(clk), .RST(start), .I(x[168]), .Q(
        xin[168]) );
  DFF \xreg_reg[170]  ( .D(xin[168]), .CLK(clk), .RST(start), .I(x[170]), .Q(
        xin[170]) );
  DFF \xreg_reg[172]  ( .D(xin[170]), .CLK(clk), .RST(start), .I(x[172]), .Q(
        xin[172]) );
  DFF \xreg_reg[174]  ( .D(xin[172]), .CLK(clk), .RST(start), .I(x[174]), .Q(
        xin[174]) );
  DFF \xreg_reg[176]  ( .D(xin[174]), .CLK(clk), .RST(start), .I(x[176]), .Q(
        xin[176]) );
  DFF \xreg_reg[178]  ( .D(xin[176]), .CLK(clk), .RST(start), .I(x[178]), .Q(
        xin[178]) );
  DFF \xreg_reg[180]  ( .D(xin[178]), .CLK(clk), .RST(start), .I(x[180]), .Q(
        xin[180]) );
  DFF \xreg_reg[182]  ( .D(xin[180]), .CLK(clk), .RST(start), .I(x[182]), .Q(
        xin[182]) );
  DFF \xreg_reg[184]  ( .D(xin[182]), .CLK(clk), .RST(start), .I(x[184]), .Q(
        xin[184]) );
  DFF \xreg_reg[186]  ( .D(xin[184]), .CLK(clk), .RST(start), .I(x[186]), .Q(
        xin[186]) );
  DFF \xreg_reg[188]  ( .D(xin[186]), .CLK(clk), .RST(start), .I(x[188]), .Q(
        xin[188]) );
  DFF \xreg_reg[190]  ( .D(xin[188]), .CLK(clk), .RST(start), .I(x[190]), .Q(
        xin[190]) );
  DFF \xreg_reg[192]  ( .D(xin[190]), .CLK(clk), .RST(start), .I(x[192]), .Q(
        xin[192]) );
  DFF \xreg_reg[194]  ( .D(xin[192]), .CLK(clk), .RST(start), .I(x[194]), .Q(
        xin[194]) );
  DFF \xreg_reg[196]  ( .D(xin[194]), .CLK(clk), .RST(start), .I(x[196]), .Q(
        xin[196]) );
  DFF \xreg_reg[198]  ( .D(xin[196]), .CLK(clk), .RST(start), .I(x[198]), .Q(
        xin[198]) );
  DFF \xreg_reg[200]  ( .D(xin[198]), .CLK(clk), .RST(start), .I(x[200]), .Q(
        xin[200]) );
  DFF \xreg_reg[202]  ( .D(xin[200]), .CLK(clk), .RST(start), .I(x[202]), .Q(
        xin[202]) );
  DFF \xreg_reg[204]  ( .D(xin[202]), .CLK(clk), .RST(start), .I(x[204]), .Q(
        xin[204]) );
  DFF \xreg_reg[206]  ( .D(xin[204]), .CLK(clk), .RST(start), .I(x[206]), .Q(
        xin[206]) );
  DFF \xreg_reg[208]  ( .D(xin[206]), .CLK(clk), .RST(start), .I(x[208]), .Q(
        xin[208]) );
  DFF \xreg_reg[210]  ( .D(xin[208]), .CLK(clk), .RST(start), .I(x[210]), .Q(
        xin[210]) );
  DFF \xreg_reg[212]  ( .D(xin[210]), .CLK(clk), .RST(start), .I(x[212]), .Q(
        xin[212]) );
  DFF \xreg_reg[214]  ( .D(xin[212]), .CLK(clk), .RST(start), .I(x[214]), .Q(
        xin[214]) );
  DFF \xreg_reg[216]  ( .D(xin[214]), .CLK(clk), .RST(start), .I(x[216]), .Q(
        xin[216]) );
  DFF \xreg_reg[218]  ( .D(xin[216]), .CLK(clk), .RST(start), .I(x[218]), .Q(
        xin[218]) );
  DFF \xreg_reg[220]  ( .D(xin[218]), .CLK(clk), .RST(start), .I(x[220]), .Q(
        xin[220]) );
  DFF \xreg_reg[222]  ( .D(xin[220]), .CLK(clk), .RST(start), .I(x[222]), .Q(
        xin[222]) );
  DFF \xreg_reg[224]  ( .D(xin[222]), .CLK(clk), .RST(start), .I(x[224]), .Q(
        xin[224]) );
  DFF \xreg_reg[226]  ( .D(xin[224]), .CLK(clk), .RST(start), .I(x[226]), .Q(
        xin[226]) );
  DFF \xreg_reg[228]  ( .D(xin[226]), .CLK(clk), .RST(start), .I(x[228]), .Q(
        xin[228]) );
  DFF \xreg_reg[230]  ( .D(xin[228]), .CLK(clk), .RST(start), .I(x[230]), .Q(
        xin[230]) );
  DFF \xreg_reg[232]  ( .D(xin[230]), .CLK(clk), .RST(start), .I(x[232]), .Q(
        xin[232]) );
  DFF \xreg_reg[234]  ( .D(xin[232]), .CLK(clk), .RST(start), .I(x[234]), .Q(
        xin[234]) );
  DFF \xreg_reg[236]  ( .D(xin[234]), .CLK(clk), .RST(start), .I(x[236]), .Q(
        xin[236]) );
  DFF \xreg_reg[238]  ( .D(xin[236]), .CLK(clk), .RST(start), .I(x[238]), .Q(
        xin[238]) );
  DFF \xreg_reg[240]  ( .D(xin[238]), .CLK(clk), .RST(start), .I(x[240]), .Q(
        xin[240]) );
  DFF \xreg_reg[242]  ( .D(xin[240]), .CLK(clk), .RST(start), .I(x[242]), .Q(
        xin[242]) );
  DFF \xreg_reg[244]  ( .D(xin[242]), .CLK(clk), .RST(start), .I(x[244]), .Q(
        xin[244]) );
  DFF \xreg_reg[246]  ( .D(xin[244]), .CLK(clk), .RST(start), .I(x[246]), .Q(
        xin[246]) );
  DFF \xreg_reg[248]  ( .D(xin[246]), .CLK(clk), .RST(start), .I(x[248]), .Q(
        xin[248]) );
  DFF \xreg_reg[250]  ( .D(xin[248]), .CLK(clk), .RST(start), .I(x[250]), .Q(
        xin[250]) );
  DFF \xreg_reg[252]  ( .D(xin[250]), .CLK(clk), .RST(start), .I(x[252]), .Q(
        xin[252]) );
  DFF \xreg_reg[254]  ( .D(xin[252]), .CLK(clk), .RST(start), .I(x[254]), .Q(
        xin[254]) );
  DFF \zreg_reg[0]  ( .D(o[0]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][0] ) );
  DFF \zreg_reg[1]  ( .D(o[1]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][1] ) );
  DFF \zreg_reg[2]  ( .D(o[2]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][2] ) );
  DFF \zreg_reg[3]  ( .D(o[3]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][3] ) );
  DFF \zreg_reg[4]  ( .D(o[4]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][4] ) );
  DFF \zreg_reg[5]  ( .D(o[5]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][5] ) );
  DFF \zreg_reg[6]  ( .D(o[6]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][6] ) );
  DFF \zreg_reg[7]  ( .D(o[7]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][7] ) );
  DFF \zreg_reg[8]  ( .D(o[8]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][8] ) );
  DFF \zreg_reg[9]  ( .D(o[9]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][9] ) );
  DFF \zreg_reg[10]  ( .D(o[10]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][10] ) );
  DFF \zreg_reg[11]  ( .D(o[11]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][11] ) );
  DFF \zreg_reg[12]  ( .D(o[12]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][12] ) );
  DFF \zreg_reg[13]  ( .D(o[13]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][13] ) );
  DFF \zreg_reg[14]  ( .D(o[14]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][14] ) );
  DFF \zreg_reg[15]  ( .D(o[15]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][15] ) );
  DFF \zreg_reg[16]  ( .D(o[16]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][16] ) );
  DFF \zreg_reg[17]  ( .D(o[17]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][17] ) );
  DFF \zreg_reg[18]  ( .D(o[18]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][18] ) );
  DFF \zreg_reg[19]  ( .D(o[19]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][19] ) );
  DFF \zreg_reg[20]  ( .D(o[20]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][20] ) );
  DFF \zreg_reg[21]  ( .D(o[21]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][21] ) );
  DFF \zreg_reg[22]  ( .D(o[22]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][22] ) );
  DFF \zreg_reg[23]  ( .D(o[23]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][23] ) );
  DFF \zreg_reg[24]  ( .D(o[24]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][24] ) );
  DFF \zreg_reg[25]  ( .D(o[25]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][25] ) );
  DFF \zreg_reg[26]  ( .D(o[26]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][26] ) );
  DFF \zreg_reg[27]  ( .D(o[27]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][27] ) );
  DFF \zreg_reg[28]  ( .D(o[28]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][28] ) );
  DFF \zreg_reg[29]  ( .D(o[29]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][29] ) );
  DFF \zreg_reg[30]  ( .D(o[30]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][30] ) );
  DFF \zreg_reg[31]  ( .D(o[31]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][31] ) );
  DFF \zreg_reg[32]  ( .D(o[32]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][32] ) );
  DFF \zreg_reg[33]  ( .D(o[33]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][33] ) );
  DFF \zreg_reg[34]  ( .D(o[34]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][34] ) );
  DFF \zreg_reg[35]  ( .D(o[35]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][35] ) );
  DFF \zreg_reg[36]  ( .D(o[36]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][36] ) );
  DFF \zreg_reg[37]  ( .D(o[37]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][37] ) );
  DFF \zreg_reg[38]  ( .D(o[38]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][38] ) );
  DFF \zreg_reg[39]  ( .D(o[39]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][39] ) );
  DFF \zreg_reg[40]  ( .D(o[40]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][40] ) );
  DFF \zreg_reg[41]  ( .D(o[41]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][41] ) );
  DFF \zreg_reg[42]  ( .D(o[42]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][42] ) );
  DFF \zreg_reg[43]  ( .D(o[43]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][43] ) );
  DFF \zreg_reg[44]  ( .D(o[44]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][44] ) );
  DFF \zreg_reg[45]  ( .D(o[45]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][45] ) );
  DFF \zreg_reg[46]  ( .D(o[46]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][46] ) );
  DFF \zreg_reg[47]  ( .D(o[47]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][47] ) );
  DFF \zreg_reg[48]  ( .D(o[48]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][48] ) );
  DFF \zreg_reg[49]  ( .D(o[49]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][49] ) );
  DFF \zreg_reg[50]  ( .D(o[50]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][50] ) );
  DFF \zreg_reg[51]  ( .D(o[51]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][51] ) );
  DFF \zreg_reg[52]  ( .D(o[52]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][52] ) );
  DFF \zreg_reg[53]  ( .D(o[53]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][53] ) );
  DFF \zreg_reg[54]  ( .D(o[54]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][54] ) );
  DFF \zreg_reg[55]  ( .D(o[55]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][55] ) );
  DFF \zreg_reg[56]  ( .D(o[56]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][56] ) );
  DFF \zreg_reg[57]  ( .D(o[57]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][57] ) );
  DFF \zreg_reg[58]  ( .D(o[58]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][58] ) );
  DFF \zreg_reg[59]  ( .D(o[59]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][59] ) );
  DFF \zreg_reg[60]  ( .D(o[60]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][60] ) );
  DFF \zreg_reg[61]  ( .D(o[61]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][61] ) );
  DFF \zreg_reg[62]  ( .D(o[62]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][62] ) );
  DFF \zreg_reg[63]  ( .D(o[63]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][63] ) );
  DFF \zreg_reg[64]  ( .D(o[64]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][64] ) );
  DFF \zreg_reg[65]  ( .D(o[65]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][65] ) );
  DFF \zreg_reg[66]  ( .D(o[66]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][66] ) );
  DFF \zreg_reg[67]  ( .D(o[67]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][67] ) );
  DFF \zreg_reg[68]  ( .D(o[68]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][68] ) );
  DFF \zreg_reg[69]  ( .D(o[69]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][69] ) );
  DFF \zreg_reg[70]  ( .D(o[70]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][70] ) );
  DFF \zreg_reg[71]  ( .D(o[71]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][71] ) );
  DFF \zreg_reg[72]  ( .D(o[72]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][72] ) );
  DFF \zreg_reg[73]  ( .D(o[73]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][73] ) );
  DFF \zreg_reg[74]  ( .D(o[74]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][74] ) );
  DFF \zreg_reg[75]  ( .D(o[75]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][75] ) );
  DFF \zreg_reg[76]  ( .D(o[76]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][76] ) );
  DFF \zreg_reg[77]  ( .D(o[77]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][77] ) );
  DFF \zreg_reg[78]  ( .D(o[78]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][78] ) );
  DFF \zreg_reg[79]  ( .D(o[79]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][79] ) );
  DFF \zreg_reg[80]  ( .D(o[80]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][80] ) );
  DFF \zreg_reg[81]  ( .D(o[81]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][81] ) );
  DFF \zreg_reg[82]  ( .D(o[82]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][82] ) );
  DFF \zreg_reg[83]  ( .D(o[83]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][83] ) );
  DFF \zreg_reg[84]  ( .D(o[84]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][84] ) );
  DFF \zreg_reg[85]  ( .D(o[85]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][85] ) );
  DFF \zreg_reg[86]  ( .D(o[86]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][86] ) );
  DFF \zreg_reg[87]  ( .D(o[87]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][87] ) );
  DFF \zreg_reg[88]  ( .D(o[88]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][88] ) );
  DFF \zreg_reg[89]  ( .D(o[89]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][89] ) );
  DFF \zreg_reg[90]  ( .D(o[90]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][90] ) );
  DFF \zreg_reg[91]  ( .D(o[91]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][91] ) );
  DFF \zreg_reg[92]  ( .D(o[92]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][92] ) );
  DFF \zreg_reg[93]  ( .D(o[93]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][93] ) );
  DFF \zreg_reg[94]  ( .D(o[94]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][94] ) );
  DFF \zreg_reg[95]  ( .D(o[95]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][95] ) );
  DFF \zreg_reg[96]  ( .D(o[96]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][96] ) );
  DFF \zreg_reg[97]  ( .D(o[97]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][97] ) );
  DFF \zreg_reg[98]  ( .D(o[98]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][98] ) );
  DFF \zreg_reg[99]  ( .D(o[99]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][99] ) );
  DFF \zreg_reg[100]  ( .D(o[100]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][100] ) );
  DFF \zreg_reg[101]  ( .D(o[101]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][101] ) );
  DFF \zreg_reg[102]  ( .D(o[102]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][102] ) );
  DFF \zreg_reg[103]  ( .D(o[103]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][103] ) );
  DFF \zreg_reg[104]  ( .D(o[104]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][104] ) );
  DFF \zreg_reg[105]  ( .D(o[105]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][105] ) );
  DFF \zreg_reg[106]  ( .D(o[106]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][106] ) );
  DFF \zreg_reg[107]  ( .D(o[107]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][107] ) );
  DFF \zreg_reg[108]  ( .D(o[108]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][108] ) );
  DFF \zreg_reg[109]  ( .D(o[109]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][109] ) );
  DFF \zreg_reg[110]  ( .D(o[110]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][110] ) );
  DFF \zreg_reg[111]  ( .D(o[111]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][111] ) );
  DFF \zreg_reg[112]  ( .D(o[112]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][112] ) );
  DFF \zreg_reg[113]  ( .D(o[113]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][113] ) );
  DFF \zreg_reg[114]  ( .D(o[114]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][114] ) );
  DFF \zreg_reg[115]  ( .D(o[115]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][115] ) );
  DFF \zreg_reg[116]  ( .D(o[116]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][116] ) );
  DFF \zreg_reg[117]  ( .D(o[117]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][117] ) );
  DFF \zreg_reg[118]  ( .D(o[118]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][118] ) );
  DFF \zreg_reg[119]  ( .D(o[119]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][119] ) );
  DFF \zreg_reg[120]  ( .D(o[120]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][120] ) );
  DFF \zreg_reg[121]  ( .D(o[121]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][121] ) );
  DFF \zreg_reg[122]  ( .D(o[122]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][122] ) );
  DFF \zreg_reg[123]  ( .D(o[123]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][123] ) );
  DFF \zreg_reg[124]  ( .D(o[124]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][124] ) );
  DFF \zreg_reg[125]  ( .D(o[125]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][125] ) );
  DFF \zreg_reg[126]  ( .D(o[126]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][126] ) );
  DFF \zreg_reg[127]  ( .D(o[127]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][127] ) );
  DFF \zreg_reg[128]  ( .D(o[128]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][128] ) );
  DFF \zreg_reg[129]  ( .D(o[129]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][129] ) );
  DFF \zreg_reg[130]  ( .D(o[130]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][130] ) );
  DFF \zreg_reg[131]  ( .D(o[131]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][131] ) );
  DFF \zreg_reg[132]  ( .D(o[132]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][132] ) );
  DFF \zreg_reg[133]  ( .D(o[133]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][133] ) );
  DFF \zreg_reg[134]  ( .D(o[134]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][134] ) );
  DFF \zreg_reg[135]  ( .D(o[135]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][135] ) );
  DFF \zreg_reg[136]  ( .D(o[136]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][136] ) );
  DFF \zreg_reg[137]  ( .D(o[137]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][137] ) );
  DFF \zreg_reg[138]  ( .D(o[138]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][138] ) );
  DFF \zreg_reg[139]  ( .D(o[139]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][139] ) );
  DFF \zreg_reg[140]  ( .D(o[140]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][140] ) );
  DFF \zreg_reg[141]  ( .D(o[141]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][141] ) );
  DFF \zreg_reg[142]  ( .D(o[142]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][142] ) );
  DFF \zreg_reg[143]  ( .D(o[143]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][143] ) );
  DFF \zreg_reg[144]  ( .D(o[144]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][144] ) );
  DFF \zreg_reg[145]  ( .D(o[145]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][145] ) );
  DFF \zreg_reg[146]  ( .D(o[146]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][146] ) );
  DFF \zreg_reg[147]  ( .D(o[147]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][147] ) );
  DFF \zreg_reg[148]  ( .D(o[148]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][148] ) );
  DFF \zreg_reg[149]  ( .D(o[149]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][149] ) );
  DFF \zreg_reg[150]  ( .D(o[150]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][150] ) );
  DFF \zreg_reg[151]  ( .D(o[151]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][151] ) );
  DFF \zreg_reg[152]  ( .D(o[152]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][152] ) );
  DFF \zreg_reg[153]  ( .D(o[153]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][153] ) );
  DFF \zreg_reg[154]  ( .D(o[154]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][154] ) );
  DFF \zreg_reg[155]  ( .D(o[155]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][155] ) );
  DFF \zreg_reg[156]  ( .D(o[156]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][156] ) );
  DFF \zreg_reg[157]  ( .D(o[157]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][157] ) );
  DFF \zreg_reg[158]  ( .D(o[158]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][158] ) );
  DFF \zreg_reg[159]  ( .D(o[159]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][159] ) );
  DFF \zreg_reg[160]  ( .D(o[160]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][160] ) );
  DFF \zreg_reg[161]  ( .D(o[161]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][161] ) );
  DFF \zreg_reg[162]  ( .D(o[162]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][162] ) );
  DFF \zreg_reg[163]  ( .D(o[163]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][163] ) );
  DFF \zreg_reg[164]  ( .D(o[164]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][164] ) );
  DFF \zreg_reg[165]  ( .D(o[165]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][165] ) );
  DFF \zreg_reg[166]  ( .D(o[166]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][166] ) );
  DFF \zreg_reg[167]  ( .D(o[167]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][167] ) );
  DFF \zreg_reg[168]  ( .D(o[168]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][168] ) );
  DFF \zreg_reg[169]  ( .D(o[169]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][169] ) );
  DFF \zreg_reg[170]  ( .D(o[170]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][170] ) );
  DFF \zreg_reg[171]  ( .D(o[171]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][171] ) );
  DFF \zreg_reg[172]  ( .D(o[172]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][172] ) );
  DFF \zreg_reg[173]  ( .D(o[173]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][173] ) );
  DFF \zreg_reg[174]  ( .D(o[174]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][174] ) );
  DFF \zreg_reg[175]  ( .D(o[175]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][175] ) );
  DFF \zreg_reg[176]  ( .D(o[176]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][176] ) );
  DFF \zreg_reg[177]  ( .D(o[177]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][177] ) );
  DFF \zreg_reg[178]  ( .D(o[178]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][178] ) );
  DFF \zreg_reg[179]  ( .D(o[179]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][179] ) );
  DFF \zreg_reg[180]  ( .D(o[180]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][180] ) );
  DFF \zreg_reg[181]  ( .D(o[181]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][181] ) );
  DFF \zreg_reg[182]  ( .D(o[182]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][182] ) );
  DFF \zreg_reg[183]  ( .D(o[183]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][183] ) );
  DFF \zreg_reg[184]  ( .D(o[184]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][184] ) );
  DFF \zreg_reg[185]  ( .D(o[185]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][185] ) );
  DFF \zreg_reg[186]  ( .D(o[186]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][186] ) );
  DFF \zreg_reg[187]  ( .D(o[187]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][187] ) );
  DFF \zreg_reg[188]  ( .D(o[188]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][188] ) );
  DFF \zreg_reg[189]  ( .D(o[189]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][189] ) );
  DFF \zreg_reg[190]  ( .D(o[190]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][190] ) );
  DFF \zreg_reg[191]  ( .D(o[191]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][191] ) );
  DFF \zreg_reg[192]  ( .D(o[192]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][192] ) );
  DFF \zreg_reg[193]  ( .D(o[193]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][193] ) );
  DFF \zreg_reg[194]  ( .D(o[194]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][194] ) );
  DFF \zreg_reg[195]  ( .D(o[195]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][195] ) );
  DFF \zreg_reg[196]  ( .D(o[196]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][196] ) );
  DFF \zreg_reg[197]  ( .D(o[197]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][197] ) );
  DFF \zreg_reg[198]  ( .D(o[198]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][198] ) );
  DFF \zreg_reg[199]  ( .D(o[199]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][199] ) );
  DFF \zreg_reg[200]  ( .D(o[200]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][200] ) );
  DFF \zreg_reg[201]  ( .D(o[201]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][201] ) );
  DFF \zreg_reg[202]  ( .D(o[202]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][202] ) );
  DFF \zreg_reg[203]  ( .D(o[203]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][203] ) );
  DFF \zreg_reg[204]  ( .D(o[204]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][204] ) );
  DFF \zreg_reg[205]  ( .D(o[205]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][205] ) );
  DFF \zreg_reg[206]  ( .D(o[206]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][206] ) );
  DFF \zreg_reg[207]  ( .D(o[207]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][207] ) );
  DFF \zreg_reg[208]  ( .D(o[208]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][208] ) );
  DFF \zreg_reg[209]  ( .D(o[209]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][209] ) );
  DFF \zreg_reg[210]  ( .D(o[210]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][210] ) );
  DFF \zreg_reg[211]  ( .D(o[211]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][211] ) );
  DFF \zreg_reg[212]  ( .D(o[212]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][212] ) );
  DFF \zreg_reg[213]  ( .D(o[213]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][213] ) );
  DFF \zreg_reg[214]  ( .D(o[214]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][214] ) );
  DFF \zreg_reg[215]  ( .D(o[215]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][215] ) );
  DFF \zreg_reg[216]  ( .D(o[216]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][216] ) );
  DFF \zreg_reg[217]  ( .D(o[217]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][217] ) );
  DFF \zreg_reg[218]  ( .D(o[218]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][218] ) );
  DFF \zreg_reg[219]  ( .D(o[219]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][219] ) );
  DFF \zreg_reg[220]  ( .D(o[220]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][220] ) );
  DFF \zreg_reg[221]  ( .D(o[221]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][221] ) );
  DFF \zreg_reg[222]  ( .D(o[222]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][222] ) );
  DFF \zreg_reg[223]  ( .D(o[223]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][223] ) );
  DFF \zreg_reg[224]  ( .D(o[224]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][224] ) );
  DFF \zreg_reg[225]  ( .D(o[225]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][225] ) );
  DFF \zreg_reg[226]  ( .D(o[226]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][226] ) );
  DFF \zreg_reg[227]  ( .D(o[227]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][227] ) );
  DFF \zreg_reg[228]  ( .D(o[228]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][228] ) );
  DFF \zreg_reg[229]  ( .D(o[229]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][229] ) );
  DFF \zreg_reg[230]  ( .D(o[230]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][230] ) );
  DFF \zreg_reg[231]  ( .D(o[231]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][231] ) );
  DFF \zreg_reg[232]  ( .D(o[232]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][232] ) );
  DFF \zreg_reg[233]  ( .D(o[233]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][233] ) );
  DFF \zreg_reg[234]  ( .D(o[234]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][234] ) );
  DFF \zreg_reg[235]  ( .D(o[235]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][235] ) );
  DFF \zreg_reg[236]  ( .D(o[236]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][236] ) );
  DFF \zreg_reg[237]  ( .D(o[237]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][237] ) );
  DFF \zreg_reg[238]  ( .D(o[238]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][238] ) );
  DFF \zreg_reg[239]  ( .D(o[239]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][239] ) );
  DFF \zreg_reg[240]  ( .D(o[240]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][240] ) );
  DFF \zreg_reg[241]  ( .D(o[241]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][241] ) );
  DFF \zreg_reg[242]  ( .D(o[242]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][242] ) );
  DFF \zreg_reg[243]  ( .D(o[243]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][243] ) );
  DFF \zreg_reg[244]  ( .D(o[244]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][244] ) );
  DFF \zreg_reg[245]  ( .D(o[245]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][245] ) );
  DFF \zreg_reg[246]  ( .D(o[246]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][246] ) );
  DFF \zreg_reg[247]  ( .D(o[247]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][247] ) );
  DFF \zreg_reg[248]  ( .D(o[248]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][248] ) );
  DFF \zreg_reg[249]  ( .D(o[249]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][249] ) );
  DFF \zreg_reg[250]  ( .D(o[250]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][250] ) );
  DFF \zreg_reg[251]  ( .D(o[251]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][251] ) );
  DFF \zreg_reg[252]  ( .D(o[252]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][252] ) );
  DFF \zreg_reg[253]  ( .D(o[253]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][253] ) );
  DFF \zreg_reg[254]  ( .D(o[254]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][254] ) );
  DFF \zreg_reg[255]  ( .D(o[255]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][255] ) );
  DFF \zreg_reg[256]  ( .D(\zout[1][256] ), .CLK(clk), .RST(start), .I(1'b0), 
        .Q(\zin[0][256] ) );
endmodule


module MUX_N256_4 ( A, B, S, O );
  input [255:0] A;
  input [255:0] B;
  output [255:0] O;
  input S;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512;

  XOR U1 ( .A(A[9]), .B(n1), .Z(O[9]) );
  AND U2 ( .A(S), .B(n2), .Z(n1) );
  XOR U3 ( .A(B[9]), .B(A[9]), .Z(n2) );
  XOR U4 ( .A(A[99]), .B(n3), .Z(O[99]) );
  AND U5 ( .A(S), .B(n4), .Z(n3) );
  XOR U6 ( .A(B[99]), .B(A[99]), .Z(n4) );
  XOR U7 ( .A(A[98]), .B(n5), .Z(O[98]) );
  AND U8 ( .A(S), .B(n6), .Z(n5) );
  XOR U9 ( .A(B[98]), .B(A[98]), .Z(n6) );
  XOR U10 ( .A(A[97]), .B(n7), .Z(O[97]) );
  AND U11 ( .A(S), .B(n8), .Z(n7) );
  XOR U12 ( .A(B[97]), .B(A[97]), .Z(n8) );
  XOR U13 ( .A(A[96]), .B(n9), .Z(O[96]) );
  AND U14 ( .A(S), .B(n10), .Z(n9) );
  XOR U15 ( .A(B[96]), .B(A[96]), .Z(n10) );
  XOR U16 ( .A(A[95]), .B(n11), .Z(O[95]) );
  AND U17 ( .A(S), .B(n12), .Z(n11) );
  XOR U18 ( .A(B[95]), .B(A[95]), .Z(n12) );
  XOR U19 ( .A(A[94]), .B(n13), .Z(O[94]) );
  AND U20 ( .A(S), .B(n14), .Z(n13) );
  XOR U21 ( .A(B[94]), .B(A[94]), .Z(n14) );
  XOR U22 ( .A(A[93]), .B(n15), .Z(O[93]) );
  AND U23 ( .A(S), .B(n16), .Z(n15) );
  XOR U24 ( .A(B[93]), .B(A[93]), .Z(n16) );
  XOR U25 ( .A(A[92]), .B(n17), .Z(O[92]) );
  AND U26 ( .A(S), .B(n18), .Z(n17) );
  XOR U27 ( .A(B[92]), .B(A[92]), .Z(n18) );
  XOR U28 ( .A(A[91]), .B(n19), .Z(O[91]) );
  AND U29 ( .A(S), .B(n20), .Z(n19) );
  XOR U30 ( .A(B[91]), .B(A[91]), .Z(n20) );
  XOR U31 ( .A(A[90]), .B(n21), .Z(O[90]) );
  AND U32 ( .A(S), .B(n22), .Z(n21) );
  XOR U33 ( .A(B[90]), .B(A[90]), .Z(n22) );
  XOR U34 ( .A(A[8]), .B(n23), .Z(O[8]) );
  AND U35 ( .A(S), .B(n24), .Z(n23) );
  XOR U36 ( .A(B[8]), .B(A[8]), .Z(n24) );
  XOR U37 ( .A(A[89]), .B(n25), .Z(O[89]) );
  AND U38 ( .A(S), .B(n26), .Z(n25) );
  XOR U39 ( .A(B[89]), .B(A[89]), .Z(n26) );
  XOR U40 ( .A(A[88]), .B(n27), .Z(O[88]) );
  AND U41 ( .A(S), .B(n28), .Z(n27) );
  XOR U42 ( .A(B[88]), .B(A[88]), .Z(n28) );
  XOR U43 ( .A(A[87]), .B(n29), .Z(O[87]) );
  AND U44 ( .A(S), .B(n30), .Z(n29) );
  XOR U45 ( .A(B[87]), .B(A[87]), .Z(n30) );
  XOR U46 ( .A(A[86]), .B(n31), .Z(O[86]) );
  AND U47 ( .A(S), .B(n32), .Z(n31) );
  XOR U48 ( .A(B[86]), .B(A[86]), .Z(n32) );
  XOR U49 ( .A(A[85]), .B(n33), .Z(O[85]) );
  AND U50 ( .A(S), .B(n34), .Z(n33) );
  XOR U51 ( .A(B[85]), .B(A[85]), .Z(n34) );
  XOR U52 ( .A(A[84]), .B(n35), .Z(O[84]) );
  AND U53 ( .A(S), .B(n36), .Z(n35) );
  XOR U54 ( .A(B[84]), .B(A[84]), .Z(n36) );
  XOR U55 ( .A(A[83]), .B(n37), .Z(O[83]) );
  AND U56 ( .A(S), .B(n38), .Z(n37) );
  XOR U57 ( .A(B[83]), .B(A[83]), .Z(n38) );
  XOR U58 ( .A(A[82]), .B(n39), .Z(O[82]) );
  AND U59 ( .A(S), .B(n40), .Z(n39) );
  XOR U60 ( .A(B[82]), .B(A[82]), .Z(n40) );
  XOR U61 ( .A(A[81]), .B(n41), .Z(O[81]) );
  AND U62 ( .A(S), .B(n42), .Z(n41) );
  XOR U63 ( .A(B[81]), .B(A[81]), .Z(n42) );
  XOR U64 ( .A(A[80]), .B(n43), .Z(O[80]) );
  AND U65 ( .A(S), .B(n44), .Z(n43) );
  XOR U66 ( .A(B[80]), .B(A[80]), .Z(n44) );
  XOR U67 ( .A(A[7]), .B(n45), .Z(O[7]) );
  AND U68 ( .A(S), .B(n46), .Z(n45) );
  XOR U69 ( .A(B[7]), .B(A[7]), .Z(n46) );
  XOR U70 ( .A(A[79]), .B(n47), .Z(O[79]) );
  AND U71 ( .A(S), .B(n48), .Z(n47) );
  XOR U72 ( .A(B[79]), .B(A[79]), .Z(n48) );
  XOR U73 ( .A(A[78]), .B(n49), .Z(O[78]) );
  AND U74 ( .A(S), .B(n50), .Z(n49) );
  XOR U75 ( .A(B[78]), .B(A[78]), .Z(n50) );
  XOR U76 ( .A(A[77]), .B(n51), .Z(O[77]) );
  AND U77 ( .A(S), .B(n52), .Z(n51) );
  XOR U78 ( .A(B[77]), .B(A[77]), .Z(n52) );
  XOR U79 ( .A(A[76]), .B(n53), .Z(O[76]) );
  AND U80 ( .A(S), .B(n54), .Z(n53) );
  XOR U81 ( .A(B[76]), .B(A[76]), .Z(n54) );
  XOR U82 ( .A(A[75]), .B(n55), .Z(O[75]) );
  AND U83 ( .A(S), .B(n56), .Z(n55) );
  XOR U84 ( .A(B[75]), .B(A[75]), .Z(n56) );
  XOR U85 ( .A(A[74]), .B(n57), .Z(O[74]) );
  AND U86 ( .A(S), .B(n58), .Z(n57) );
  XOR U87 ( .A(B[74]), .B(A[74]), .Z(n58) );
  XOR U88 ( .A(A[73]), .B(n59), .Z(O[73]) );
  AND U89 ( .A(S), .B(n60), .Z(n59) );
  XOR U90 ( .A(B[73]), .B(A[73]), .Z(n60) );
  XOR U91 ( .A(A[72]), .B(n61), .Z(O[72]) );
  AND U92 ( .A(S), .B(n62), .Z(n61) );
  XOR U93 ( .A(B[72]), .B(A[72]), .Z(n62) );
  XOR U94 ( .A(A[71]), .B(n63), .Z(O[71]) );
  AND U95 ( .A(S), .B(n64), .Z(n63) );
  XOR U96 ( .A(B[71]), .B(A[71]), .Z(n64) );
  XOR U97 ( .A(A[70]), .B(n65), .Z(O[70]) );
  AND U98 ( .A(S), .B(n66), .Z(n65) );
  XOR U99 ( .A(B[70]), .B(A[70]), .Z(n66) );
  XOR U100 ( .A(A[6]), .B(n67), .Z(O[6]) );
  AND U101 ( .A(S), .B(n68), .Z(n67) );
  XOR U102 ( .A(B[6]), .B(A[6]), .Z(n68) );
  XOR U103 ( .A(A[69]), .B(n69), .Z(O[69]) );
  AND U104 ( .A(S), .B(n70), .Z(n69) );
  XOR U105 ( .A(B[69]), .B(A[69]), .Z(n70) );
  XOR U106 ( .A(A[68]), .B(n71), .Z(O[68]) );
  AND U107 ( .A(S), .B(n72), .Z(n71) );
  XOR U108 ( .A(B[68]), .B(A[68]), .Z(n72) );
  XOR U109 ( .A(A[67]), .B(n73), .Z(O[67]) );
  AND U110 ( .A(S), .B(n74), .Z(n73) );
  XOR U111 ( .A(B[67]), .B(A[67]), .Z(n74) );
  XOR U112 ( .A(A[66]), .B(n75), .Z(O[66]) );
  AND U113 ( .A(S), .B(n76), .Z(n75) );
  XOR U114 ( .A(B[66]), .B(A[66]), .Z(n76) );
  XOR U115 ( .A(A[65]), .B(n77), .Z(O[65]) );
  AND U116 ( .A(S), .B(n78), .Z(n77) );
  XOR U117 ( .A(B[65]), .B(A[65]), .Z(n78) );
  XOR U118 ( .A(A[64]), .B(n79), .Z(O[64]) );
  AND U119 ( .A(S), .B(n80), .Z(n79) );
  XOR U120 ( .A(B[64]), .B(A[64]), .Z(n80) );
  XOR U121 ( .A(A[63]), .B(n81), .Z(O[63]) );
  AND U122 ( .A(S), .B(n82), .Z(n81) );
  XOR U123 ( .A(B[63]), .B(A[63]), .Z(n82) );
  XOR U124 ( .A(A[62]), .B(n83), .Z(O[62]) );
  AND U125 ( .A(S), .B(n84), .Z(n83) );
  XOR U126 ( .A(B[62]), .B(A[62]), .Z(n84) );
  XOR U127 ( .A(A[61]), .B(n85), .Z(O[61]) );
  AND U128 ( .A(S), .B(n86), .Z(n85) );
  XOR U129 ( .A(B[61]), .B(A[61]), .Z(n86) );
  XOR U130 ( .A(A[60]), .B(n87), .Z(O[60]) );
  AND U131 ( .A(S), .B(n88), .Z(n87) );
  XOR U132 ( .A(B[60]), .B(A[60]), .Z(n88) );
  XOR U133 ( .A(A[5]), .B(n89), .Z(O[5]) );
  AND U134 ( .A(S), .B(n90), .Z(n89) );
  XOR U135 ( .A(B[5]), .B(A[5]), .Z(n90) );
  XOR U136 ( .A(A[59]), .B(n91), .Z(O[59]) );
  AND U137 ( .A(S), .B(n92), .Z(n91) );
  XOR U138 ( .A(B[59]), .B(A[59]), .Z(n92) );
  XOR U139 ( .A(A[58]), .B(n93), .Z(O[58]) );
  AND U140 ( .A(S), .B(n94), .Z(n93) );
  XOR U141 ( .A(B[58]), .B(A[58]), .Z(n94) );
  XOR U142 ( .A(A[57]), .B(n95), .Z(O[57]) );
  AND U143 ( .A(S), .B(n96), .Z(n95) );
  XOR U144 ( .A(B[57]), .B(A[57]), .Z(n96) );
  XOR U145 ( .A(A[56]), .B(n97), .Z(O[56]) );
  AND U146 ( .A(S), .B(n98), .Z(n97) );
  XOR U147 ( .A(B[56]), .B(A[56]), .Z(n98) );
  XOR U148 ( .A(A[55]), .B(n99), .Z(O[55]) );
  AND U149 ( .A(S), .B(n100), .Z(n99) );
  XOR U150 ( .A(B[55]), .B(A[55]), .Z(n100) );
  XOR U151 ( .A(A[54]), .B(n101), .Z(O[54]) );
  AND U152 ( .A(S), .B(n102), .Z(n101) );
  XOR U153 ( .A(B[54]), .B(A[54]), .Z(n102) );
  XOR U154 ( .A(A[53]), .B(n103), .Z(O[53]) );
  AND U155 ( .A(S), .B(n104), .Z(n103) );
  XOR U156 ( .A(B[53]), .B(A[53]), .Z(n104) );
  XOR U157 ( .A(A[52]), .B(n105), .Z(O[52]) );
  AND U158 ( .A(S), .B(n106), .Z(n105) );
  XOR U159 ( .A(B[52]), .B(A[52]), .Z(n106) );
  XOR U160 ( .A(A[51]), .B(n107), .Z(O[51]) );
  AND U161 ( .A(S), .B(n108), .Z(n107) );
  XOR U162 ( .A(B[51]), .B(A[51]), .Z(n108) );
  XOR U163 ( .A(A[50]), .B(n109), .Z(O[50]) );
  AND U164 ( .A(S), .B(n110), .Z(n109) );
  XOR U165 ( .A(B[50]), .B(A[50]), .Z(n110) );
  XOR U166 ( .A(A[4]), .B(n111), .Z(O[4]) );
  AND U167 ( .A(S), .B(n112), .Z(n111) );
  XOR U168 ( .A(B[4]), .B(A[4]), .Z(n112) );
  XOR U169 ( .A(A[49]), .B(n113), .Z(O[49]) );
  AND U170 ( .A(S), .B(n114), .Z(n113) );
  XOR U171 ( .A(B[49]), .B(A[49]), .Z(n114) );
  XOR U172 ( .A(A[48]), .B(n115), .Z(O[48]) );
  AND U173 ( .A(S), .B(n116), .Z(n115) );
  XOR U174 ( .A(B[48]), .B(A[48]), .Z(n116) );
  XOR U175 ( .A(A[47]), .B(n117), .Z(O[47]) );
  AND U176 ( .A(S), .B(n118), .Z(n117) );
  XOR U177 ( .A(B[47]), .B(A[47]), .Z(n118) );
  XOR U178 ( .A(A[46]), .B(n119), .Z(O[46]) );
  AND U179 ( .A(S), .B(n120), .Z(n119) );
  XOR U180 ( .A(B[46]), .B(A[46]), .Z(n120) );
  XOR U181 ( .A(A[45]), .B(n121), .Z(O[45]) );
  AND U182 ( .A(S), .B(n122), .Z(n121) );
  XOR U183 ( .A(B[45]), .B(A[45]), .Z(n122) );
  XOR U184 ( .A(A[44]), .B(n123), .Z(O[44]) );
  AND U185 ( .A(S), .B(n124), .Z(n123) );
  XOR U186 ( .A(B[44]), .B(A[44]), .Z(n124) );
  XOR U187 ( .A(A[43]), .B(n125), .Z(O[43]) );
  AND U188 ( .A(S), .B(n126), .Z(n125) );
  XOR U189 ( .A(B[43]), .B(A[43]), .Z(n126) );
  XOR U190 ( .A(A[42]), .B(n127), .Z(O[42]) );
  AND U191 ( .A(S), .B(n128), .Z(n127) );
  XOR U192 ( .A(B[42]), .B(A[42]), .Z(n128) );
  XOR U193 ( .A(A[41]), .B(n129), .Z(O[41]) );
  AND U194 ( .A(S), .B(n130), .Z(n129) );
  XOR U195 ( .A(B[41]), .B(A[41]), .Z(n130) );
  XOR U196 ( .A(A[40]), .B(n131), .Z(O[40]) );
  AND U197 ( .A(S), .B(n132), .Z(n131) );
  XOR U198 ( .A(B[40]), .B(A[40]), .Z(n132) );
  XOR U199 ( .A(A[3]), .B(n133), .Z(O[3]) );
  AND U200 ( .A(S), .B(n134), .Z(n133) );
  XOR U201 ( .A(B[3]), .B(A[3]), .Z(n134) );
  XOR U202 ( .A(A[39]), .B(n135), .Z(O[39]) );
  AND U203 ( .A(S), .B(n136), .Z(n135) );
  XOR U204 ( .A(B[39]), .B(A[39]), .Z(n136) );
  XOR U205 ( .A(A[38]), .B(n137), .Z(O[38]) );
  AND U206 ( .A(S), .B(n138), .Z(n137) );
  XOR U207 ( .A(B[38]), .B(A[38]), .Z(n138) );
  XOR U208 ( .A(A[37]), .B(n139), .Z(O[37]) );
  AND U209 ( .A(S), .B(n140), .Z(n139) );
  XOR U210 ( .A(B[37]), .B(A[37]), .Z(n140) );
  XOR U211 ( .A(A[36]), .B(n141), .Z(O[36]) );
  AND U212 ( .A(S), .B(n142), .Z(n141) );
  XOR U213 ( .A(B[36]), .B(A[36]), .Z(n142) );
  XOR U214 ( .A(A[35]), .B(n143), .Z(O[35]) );
  AND U215 ( .A(S), .B(n144), .Z(n143) );
  XOR U216 ( .A(B[35]), .B(A[35]), .Z(n144) );
  XOR U217 ( .A(A[34]), .B(n145), .Z(O[34]) );
  AND U218 ( .A(S), .B(n146), .Z(n145) );
  XOR U219 ( .A(B[34]), .B(A[34]), .Z(n146) );
  XOR U220 ( .A(A[33]), .B(n147), .Z(O[33]) );
  AND U221 ( .A(S), .B(n148), .Z(n147) );
  XOR U222 ( .A(B[33]), .B(A[33]), .Z(n148) );
  XOR U223 ( .A(A[32]), .B(n149), .Z(O[32]) );
  AND U224 ( .A(S), .B(n150), .Z(n149) );
  XOR U225 ( .A(B[32]), .B(A[32]), .Z(n150) );
  XOR U226 ( .A(A[31]), .B(n151), .Z(O[31]) );
  AND U227 ( .A(S), .B(n152), .Z(n151) );
  XOR U228 ( .A(B[31]), .B(A[31]), .Z(n152) );
  XOR U229 ( .A(A[30]), .B(n153), .Z(O[30]) );
  AND U230 ( .A(S), .B(n154), .Z(n153) );
  XOR U231 ( .A(B[30]), .B(A[30]), .Z(n154) );
  XOR U232 ( .A(A[2]), .B(n155), .Z(O[2]) );
  AND U233 ( .A(S), .B(n156), .Z(n155) );
  XOR U234 ( .A(B[2]), .B(A[2]), .Z(n156) );
  XOR U235 ( .A(A[29]), .B(n157), .Z(O[29]) );
  AND U236 ( .A(S), .B(n158), .Z(n157) );
  XOR U237 ( .A(B[29]), .B(A[29]), .Z(n158) );
  XOR U238 ( .A(A[28]), .B(n159), .Z(O[28]) );
  AND U239 ( .A(S), .B(n160), .Z(n159) );
  XOR U240 ( .A(B[28]), .B(A[28]), .Z(n160) );
  XOR U241 ( .A(A[27]), .B(n161), .Z(O[27]) );
  AND U242 ( .A(S), .B(n162), .Z(n161) );
  XOR U243 ( .A(B[27]), .B(A[27]), .Z(n162) );
  XOR U244 ( .A(A[26]), .B(n163), .Z(O[26]) );
  AND U245 ( .A(S), .B(n164), .Z(n163) );
  XOR U246 ( .A(B[26]), .B(A[26]), .Z(n164) );
  XOR U247 ( .A(A[25]), .B(n165), .Z(O[25]) );
  AND U248 ( .A(S), .B(n166), .Z(n165) );
  XOR U249 ( .A(B[25]), .B(A[25]), .Z(n166) );
  XOR U250 ( .A(A[255]), .B(n167), .Z(O[255]) );
  AND U251 ( .A(S), .B(n168), .Z(n167) );
  XOR U252 ( .A(B[255]), .B(A[255]), .Z(n168) );
  XOR U253 ( .A(A[254]), .B(n169), .Z(O[254]) );
  AND U254 ( .A(S), .B(n170), .Z(n169) );
  XOR U255 ( .A(B[254]), .B(A[254]), .Z(n170) );
  XOR U256 ( .A(A[253]), .B(n171), .Z(O[253]) );
  AND U257 ( .A(S), .B(n172), .Z(n171) );
  XOR U258 ( .A(B[253]), .B(A[253]), .Z(n172) );
  XOR U259 ( .A(A[252]), .B(n173), .Z(O[252]) );
  AND U260 ( .A(S), .B(n174), .Z(n173) );
  XOR U261 ( .A(B[252]), .B(A[252]), .Z(n174) );
  XOR U262 ( .A(A[251]), .B(n175), .Z(O[251]) );
  AND U263 ( .A(S), .B(n176), .Z(n175) );
  XOR U264 ( .A(B[251]), .B(A[251]), .Z(n176) );
  XOR U265 ( .A(A[250]), .B(n177), .Z(O[250]) );
  AND U266 ( .A(S), .B(n178), .Z(n177) );
  XOR U267 ( .A(B[250]), .B(A[250]), .Z(n178) );
  XOR U268 ( .A(A[24]), .B(n179), .Z(O[24]) );
  AND U269 ( .A(S), .B(n180), .Z(n179) );
  XOR U270 ( .A(B[24]), .B(A[24]), .Z(n180) );
  XOR U271 ( .A(A[249]), .B(n181), .Z(O[249]) );
  AND U272 ( .A(S), .B(n182), .Z(n181) );
  XOR U273 ( .A(B[249]), .B(A[249]), .Z(n182) );
  XOR U274 ( .A(A[248]), .B(n183), .Z(O[248]) );
  AND U275 ( .A(S), .B(n184), .Z(n183) );
  XOR U276 ( .A(B[248]), .B(A[248]), .Z(n184) );
  XOR U277 ( .A(A[247]), .B(n185), .Z(O[247]) );
  AND U278 ( .A(S), .B(n186), .Z(n185) );
  XOR U279 ( .A(B[247]), .B(A[247]), .Z(n186) );
  XOR U280 ( .A(A[246]), .B(n187), .Z(O[246]) );
  AND U281 ( .A(S), .B(n188), .Z(n187) );
  XOR U282 ( .A(B[246]), .B(A[246]), .Z(n188) );
  XOR U283 ( .A(A[245]), .B(n189), .Z(O[245]) );
  AND U284 ( .A(S), .B(n190), .Z(n189) );
  XOR U285 ( .A(B[245]), .B(A[245]), .Z(n190) );
  XOR U286 ( .A(A[244]), .B(n191), .Z(O[244]) );
  AND U287 ( .A(S), .B(n192), .Z(n191) );
  XOR U288 ( .A(B[244]), .B(A[244]), .Z(n192) );
  XOR U289 ( .A(A[243]), .B(n193), .Z(O[243]) );
  AND U290 ( .A(S), .B(n194), .Z(n193) );
  XOR U291 ( .A(B[243]), .B(A[243]), .Z(n194) );
  XOR U292 ( .A(A[242]), .B(n195), .Z(O[242]) );
  AND U293 ( .A(S), .B(n196), .Z(n195) );
  XOR U294 ( .A(B[242]), .B(A[242]), .Z(n196) );
  XOR U295 ( .A(A[241]), .B(n197), .Z(O[241]) );
  AND U296 ( .A(S), .B(n198), .Z(n197) );
  XOR U297 ( .A(B[241]), .B(A[241]), .Z(n198) );
  XOR U298 ( .A(A[240]), .B(n199), .Z(O[240]) );
  AND U299 ( .A(S), .B(n200), .Z(n199) );
  XOR U300 ( .A(B[240]), .B(A[240]), .Z(n200) );
  XOR U301 ( .A(A[23]), .B(n201), .Z(O[23]) );
  AND U302 ( .A(S), .B(n202), .Z(n201) );
  XOR U303 ( .A(B[23]), .B(A[23]), .Z(n202) );
  XOR U304 ( .A(A[239]), .B(n203), .Z(O[239]) );
  AND U305 ( .A(S), .B(n204), .Z(n203) );
  XOR U306 ( .A(B[239]), .B(A[239]), .Z(n204) );
  XOR U307 ( .A(A[238]), .B(n205), .Z(O[238]) );
  AND U308 ( .A(S), .B(n206), .Z(n205) );
  XOR U309 ( .A(B[238]), .B(A[238]), .Z(n206) );
  XOR U310 ( .A(A[237]), .B(n207), .Z(O[237]) );
  AND U311 ( .A(S), .B(n208), .Z(n207) );
  XOR U312 ( .A(B[237]), .B(A[237]), .Z(n208) );
  XOR U313 ( .A(A[236]), .B(n209), .Z(O[236]) );
  AND U314 ( .A(S), .B(n210), .Z(n209) );
  XOR U315 ( .A(B[236]), .B(A[236]), .Z(n210) );
  XOR U316 ( .A(A[235]), .B(n211), .Z(O[235]) );
  AND U317 ( .A(S), .B(n212), .Z(n211) );
  XOR U318 ( .A(B[235]), .B(A[235]), .Z(n212) );
  XOR U319 ( .A(A[234]), .B(n213), .Z(O[234]) );
  AND U320 ( .A(S), .B(n214), .Z(n213) );
  XOR U321 ( .A(B[234]), .B(A[234]), .Z(n214) );
  XOR U322 ( .A(A[233]), .B(n215), .Z(O[233]) );
  AND U323 ( .A(S), .B(n216), .Z(n215) );
  XOR U324 ( .A(B[233]), .B(A[233]), .Z(n216) );
  XOR U325 ( .A(A[232]), .B(n217), .Z(O[232]) );
  AND U326 ( .A(S), .B(n218), .Z(n217) );
  XOR U327 ( .A(B[232]), .B(A[232]), .Z(n218) );
  XOR U328 ( .A(A[231]), .B(n219), .Z(O[231]) );
  AND U329 ( .A(S), .B(n220), .Z(n219) );
  XOR U330 ( .A(B[231]), .B(A[231]), .Z(n220) );
  XOR U331 ( .A(A[230]), .B(n221), .Z(O[230]) );
  AND U332 ( .A(S), .B(n222), .Z(n221) );
  XOR U333 ( .A(B[230]), .B(A[230]), .Z(n222) );
  XOR U334 ( .A(A[22]), .B(n223), .Z(O[22]) );
  AND U335 ( .A(S), .B(n224), .Z(n223) );
  XOR U336 ( .A(B[22]), .B(A[22]), .Z(n224) );
  XOR U337 ( .A(A[229]), .B(n225), .Z(O[229]) );
  AND U338 ( .A(S), .B(n226), .Z(n225) );
  XOR U339 ( .A(B[229]), .B(A[229]), .Z(n226) );
  XOR U340 ( .A(A[228]), .B(n227), .Z(O[228]) );
  AND U341 ( .A(S), .B(n228), .Z(n227) );
  XOR U342 ( .A(B[228]), .B(A[228]), .Z(n228) );
  XOR U343 ( .A(A[227]), .B(n229), .Z(O[227]) );
  AND U344 ( .A(S), .B(n230), .Z(n229) );
  XOR U345 ( .A(B[227]), .B(A[227]), .Z(n230) );
  XOR U346 ( .A(A[226]), .B(n231), .Z(O[226]) );
  AND U347 ( .A(S), .B(n232), .Z(n231) );
  XOR U348 ( .A(B[226]), .B(A[226]), .Z(n232) );
  XOR U349 ( .A(A[225]), .B(n233), .Z(O[225]) );
  AND U350 ( .A(S), .B(n234), .Z(n233) );
  XOR U351 ( .A(B[225]), .B(A[225]), .Z(n234) );
  XOR U352 ( .A(A[224]), .B(n235), .Z(O[224]) );
  AND U353 ( .A(S), .B(n236), .Z(n235) );
  XOR U354 ( .A(B[224]), .B(A[224]), .Z(n236) );
  XOR U355 ( .A(A[223]), .B(n237), .Z(O[223]) );
  AND U356 ( .A(S), .B(n238), .Z(n237) );
  XOR U357 ( .A(B[223]), .B(A[223]), .Z(n238) );
  XOR U358 ( .A(A[222]), .B(n239), .Z(O[222]) );
  AND U359 ( .A(S), .B(n240), .Z(n239) );
  XOR U360 ( .A(B[222]), .B(A[222]), .Z(n240) );
  XOR U361 ( .A(A[221]), .B(n241), .Z(O[221]) );
  AND U362 ( .A(S), .B(n242), .Z(n241) );
  XOR U363 ( .A(B[221]), .B(A[221]), .Z(n242) );
  XOR U364 ( .A(A[220]), .B(n243), .Z(O[220]) );
  AND U365 ( .A(S), .B(n244), .Z(n243) );
  XOR U366 ( .A(B[220]), .B(A[220]), .Z(n244) );
  XOR U367 ( .A(A[21]), .B(n245), .Z(O[21]) );
  AND U368 ( .A(S), .B(n246), .Z(n245) );
  XOR U369 ( .A(B[21]), .B(A[21]), .Z(n246) );
  XOR U370 ( .A(A[219]), .B(n247), .Z(O[219]) );
  AND U371 ( .A(S), .B(n248), .Z(n247) );
  XOR U372 ( .A(B[219]), .B(A[219]), .Z(n248) );
  XOR U373 ( .A(A[218]), .B(n249), .Z(O[218]) );
  AND U374 ( .A(S), .B(n250), .Z(n249) );
  XOR U375 ( .A(B[218]), .B(A[218]), .Z(n250) );
  XOR U376 ( .A(A[217]), .B(n251), .Z(O[217]) );
  AND U377 ( .A(S), .B(n252), .Z(n251) );
  XOR U378 ( .A(B[217]), .B(A[217]), .Z(n252) );
  XOR U379 ( .A(A[216]), .B(n253), .Z(O[216]) );
  AND U380 ( .A(S), .B(n254), .Z(n253) );
  XOR U381 ( .A(B[216]), .B(A[216]), .Z(n254) );
  XOR U382 ( .A(A[215]), .B(n255), .Z(O[215]) );
  AND U383 ( .A(S), .B(n256), .Z(n255) );
  XOR U384 ( .A(B[215]), .B(A[215]), .Z(n256) );
  XOR U385 ( .A(A[214]), .B(n257), .Z(O[214]) );
  AND U386 ( .A(S), .B(n258), .Z(n257) );
  XOR U387 ( .A(B[214]), .B(A[214]), .Z(n258) );
  XOR U388 ( .A(A[213]), .B(n259), .Z(O[213]) );
  AND U389 ( .A(S), .B(n260), .Z(n259) );
  XOR U390 ( .A(B[213]), .B(A[213]), .Z(n260) );
  XOR U391 ( .A(A[212]), .B(n261), .Z(O[212]) );
  AND U392 ( .A(S), .B(n262), .Z(n261) );
  XOR U393 ( .A(B[212]), .B(A[212]), .Z(n262) );
  XOR U394 ( .A(A[211]), .B(n263), .Z(O[211]) );
  AND U395 ( .A(S), .B(n264), .Z(n263) );
  XOR U396 ( .A(B[211]), .B(A[211]), .Z(n264) );
  XOR U397 ( .A(A[210]), .B(n265), .Z(O[210]) );
  AND U398 ( .A(S), .B(n266), .Z(n265) );
  XOR U399 ( .A(B[210]), .B(A[210]), .Z(n266) );
  XOR U400 ( .A(A[20]), .B(n267), .Z(O[20]) );
  AND U401 ( .A(S), .B(n268), .Z(n267) );
  XOR U402 ( .A(B[20]), .B(A[20]), .Z(n268) );
  XOR U403 ( .A(A[209]), .B(n269), .Z(O[209]) );
  AND U404 ( .A(S), .B(n270), .Z(n269) );
  XOR U405 ( .A(B[209]), .B(A[209]), .Z(n270) );
  XOR U406 ( .A(A[208]), .B(n271), .Z(O[208]) );
  AND U407 ( .A(S), .B(n272), .Z(n271) );
  XOR U408 ( .A(B[208]), .B(A[208]), .Z(n272) );
  XOR U409 ( .A(A[207]), .B(n273), .Z(O[207]) );
  AND U410 ( .A(S), .B(n274), .Z(n273) );
  XOR U411 ( .A(B[207]), .B(A[207]), .Z(n274) );
  XOR U412 ( .A(A[206]), .B(n275), .Z(O[206]) );
  AND U413 ( .A(S), .B(n276), .Z(n275) );
  XOR U414 ( .A(B[206]), .B(A[206]), .Z(n276) );
  XOR U415 ( .A(A[205]), .B(n277), .Z(O[205]) );
  AND U416 ( .A(S), .B(n278), .Z(n277) );
  XOR U417 ( .A(B[205]), .B(A[205]), .Z(n278) );
  XOR U418 ( .A(A[204]), .B(n279), .Z(O[204]) );
  AND U419 ( .A(S), .B(n280), .Z(n279) );
  XOR U420 ( .A(B[204]), .B(A[204]), .Z(n280) );
  XOR U421 ( .A(A[203]), .B(n281), .Z(O[203]) );
  AND U422 ( .A(S), .B(n282), .Z(n281) );
  XOR U423 ( .A(B[203]), .B(A[203]), .Z(n282) );
  XOR U424 ( .A(A[202]), .B(n283), .Z(O[202]) );
  AND U425 ( .A(S), .B(n284), .Z(n283) );
  XOR U426 ( .A(B[202]), .B(A[202]), .Z(n284) );
  XOR U427 ( .A(A[201]), .B(n285), .Z(O[201]) );
  AND U428 ( .A(S), .B(n286), .Z(n285) );
  XOR U429 ( .A(B[201]), .B(A[201]), .Z(n286) );
  XOR U430 ( .A(A[200]), .B(n287), .Z(O[200]) );
  AND U431 ( .A(S), .B(n288), .Z(n287) );
  XOR U432 ( .A(B[200]), .B(A[200]), .Z(n288) );
  XOR U433 ( .A(A[1]), .B(n289), .Z(O[1]) );
  AND U434 ( .A(S), .B(n290), .Z(n289) );
  XOR U435 ( .A(B[1]), .B(A[1]), .Z(n290) );
  XOR U436 ( .A(A[19]), .B(n291), .Z(O[19]) );
  AND U437 ( .A(S), .B(n292), .Z(n291) );
  XOR U438 ( .A(B[19]), .B(A[19]), .Z(n292) );
  XOR U439 ( .A(A[199]), .B(n293), .Z(O[199]) );
  AND U440 ( .A(S), .B(n294), .Z(n293) );
  XOR U441 ( .A(B[199]), .B(A[199]), .Z(n294) );
  XOR U442 ( .A(A[198]), .B(n295), .Z(O[198]) );
  AND U443 ( .A(S), .B(n296), .Z(n295) );
  XOR U444 ( .A(B[198]), .B(A[198]), .Z(n296) );
  XOR U445 ( .A(A[197]), .B(n297), .Z(O[197]) );
  AND U446 ( .A(S), .B(n298), .Z(n297) );
  XOR U447 ( .A(B[197]), .B(A[197]), .Z(n298) );
  XOR U448 ( .A(A[196]), .B(n299), .Z(O[196]) );
  AND U449 ( .A(S), .B(n300), .Z(n299) );
  XOR U450 ( .A(B[196]), .B(A[196]), .Z(n300) );
  XOR U451 ( .A(A[195]), .B(n301), .Z(O[195]) );
  AND U452 ( .A(S), .B(n302), .Z(n301) );
  XOR U453 ( .A(B[195]), .B(A[195]), .Z(n302) );
  XOR U454 ( .A(A[194]), .B(n303), .Z(O[194]) );
  AND U455 ( .A(S), .B(n304), .Z(n303) );
  XOR U456 ( .A(B[194]), .B(A[194]), .Z(n304) );
  XOR U457 ( .A(A[193]), .B(n305), .Z(O[193]) );
  AND U458 ( .A(S), .B(n306), .Z(n305) );
  XOR U459 ( .A(B[193]), .B(A[193]), .Z(n306) );
  XOR U460 ( .A(A[192]), .B(n307), .Z(O[192]) );
  AND U461 ( .A(S), .B(n308), .Z(n307) );
  XOR U462 ( .A(B[192]), .B(A[192]), .Z(n308) );
  XOR U463 ( .A(A[191]), .B(n309), .Z(O[191]) );
  AND U464 ( .A(S), .B(n310), .Z(n309) );
  XOR U465 ( .A(B[191]), .B(A[191]), .Z(n310) );
  XOR U466 ( .A(A[190]), .B(n311), .Z(O[190]) );
  AND U467 ( .A(S), .B(n312), .Z(n311) );
  XOR U468 ( .A(B[190]), .B(A[190]), .Z(n312) );
  XOR U469 ( .A(A[18]), .B(n313), .Z(O[18]) );
  AND U470 ( .A(S), .B(n314), .Z(n313) );
  XOR U471 ( .A(B[18]), .B(A[18]), .Z(n314) );
  XOR U472 ( .A(A[189]), .B(n315), .Z(O[189]) );
  AND U473 ( .A(S), .B(n316), .Z(n315) );
  XOR U474 ( .A(B[189]), .B(A[189]), .Z(n316) );
  XOR U475 ( .A(A[188]), .B(n317), .Z(O[188]) );
  AND U476 ( .A(S), .B(n318), .Z(n317) );
  XOR U477 ( .A(B[188]), .B(A[188]), .Z(n318) );
  XOR U478 ( .A(A[187]), .B(n319), .Z(O[187]) );
  AND U479 ( .A(S), .B(n320), .Z(n319) );
  XOR U480 ( .A(B[187]), .B(A[187]), .Z(n320) );
  XOR U481 ( .A(A[186]), .B(n321), .Z(O[186]) );
  AND U482 ( .A(S), .B(n322), .Z(n321) );
  XOR U483 ( .A(B[186]), .B(A[186]), .Z(n322) );
  XOR U484 ( .A(A[185]), .B(n323), .Z(O[185]) );
  AND U485 ( .A(S), .B(n324), .Z(n323) );
  XOR U486 ( .A(B[185]), .B(A[185]), .Z(n324) );
  XOR U487 ( .A(A[184]), .B(n325), .Z(O[184]) );
  AND U488 ( .A(S), .B(n326), .Z(n325) );
  XOR U489 ( .A(B[184]), .B(A[184]), .Z(n326) );
  XOR U490 ( .A(A[183]), .B(n327), .Z(O[183]) );
  AND U491 ( .A(S), .B(n328), .Z(n327) );
  XOR U492 ( .A(B[183]), .B(A[183]), .Z(n328) );
  XOR U493 ( .A(A[182]), .B(n329), .Z(O[182]) );
  AND U494 ( .A(S), .B(n330), .Z(n329) );
  XOR U495 ( .A(B[182]), .B(A[182]), .Z(n330) );
  XOR U496 ( .A(A[181]), .B(n331), .Z(O[181]) );
  AND U497 ( .A(S), .B(n332), .Z(n331) );
  XOR U498 ( .A(B[181]), .B(A[181]), .Z(n332) );
  XOR U499 ( .A(A[180]), .B(n333), .Z(O[180]) );
  AND U500 ( .A(S), .B(n334), .Z(n333) );
  XOR U501 ( .A(B[180]), .B(A[180]), .Z(n334) );
  XOR U502 ( .A(A[17]), .B(n335), .Z(O[17]) );
  AND U503 ( .A(S), .B(n336), .Z(n335) );
  XOR U504 ( .A(B[17]), .B(A[17]), .Z(n336) );
  XOR U505 ( .A(A[179]), .B(n337), .Z(O[179]) );
  AND U506 ( .A(S), .B(n338), .Z(n337) );
  XOR U507 ( .A(B[179]), .B(A[179]), .Z(n338) );
  XOR U508 ( .A(A[178]), .B(n339), .Z(O[178]) );
  AND U509 ( .A(S), .B(n340), .Z(n339) );
  XOR U510 ( .A(B[178]), .B(A[178]), .Z(n340) );
  XOR U511 ( .A(A[177]), .B(n341), .Z(O[177]) );
  AND U512 ( .A(S), .B(n342), .Z(n341) );
  XOR U513 ( .A(B[177]), .B(A[177]), .Z(n342) );
  XOR U514 ( .A(A[176]), .B(n343), .Z(O[176]) );
  AND U515 ( .A(S), .B(n344), .Z(n343) );
  XOR U516 ( .A(B[176]), .B(A[176]), .Z(n344) );
  XOR U517 ( .A(A[175]), .B(n345), .Z(O[175]) );
  AND U518 ( .A(S), .B(n346), .Z(n345) );
  XOR U519 ( .A(B[175]), .B(A[175]), .Z(n346) );
  XOR U520 ( .A(A[174]), .B(n347), .Z(O[174]) );
  AND U521 ( .A(S), .B(n348), .Z(n347) );
  XOR U522 ( .A(B[174]), .B(A[174]), .Z(n348) );
  XOR U523 ( .A(A[173]), .B(n349), .Z(O[173]) );
  AND U524 ( .A(S), .B(n350), .Z(n349) );
  XOR U525 ( .A(B[173]), .B(A[173]), .Z(n350) );
  XOR U526 ( .A(A[172]), .B(n351), .Z(O[172]) );
  AND U527 ( .A(S), .B(n352), .Z(n351) );
  XOR U528 ( .A(B[172]), .B(A[172]), .Z(n352) );
  XOR U529 ( .A(A[171]), .B(n353), .Z(O[171]) );
  AND U530 ( .A(S), .B(n354), .Z(n353) );
  XOR U531 ( .A(B[171]), .B(A[171]), .Z(n354) );
  XOR U532 ( .A(A[170]), .B(n355), .Z(O[170]) );
  AND U533 ( .A(S), .B(n356), .Z(n355) );
  XOR U534 ( .A(B[170]), .B(A[170]), .Z(n356) );
  XOR U535 ( .A(A[16]), .B(n357), .Z(O[16]) );
  AND U536 ( .A(S), .B(n358), .Z(n357) );
  XOR U537 ( .A(B[16]), .B(A[16]), .Z(n358) );
  XOR U538 ( .A(A[169]), .B(n359), .Z(O[169]) );
  AND U539 ( .A(S), .B(n360), .Z(n359) );
  XOR U540 ( .A(B[169]), .B(A[169]), .Z(n360) );
  XOR U541 ( .A(A[168]), .B(n361), .Z(O[168]) );
  AND U542 ( .A(S), .B(n362), .Z(n361) );
  XOR U543 ( .A(B[168]), .B(A[168]), .Z(n362) );
  XOR U544 ( .A(A[167]), .B(n363), .Z(O[167]) );
  AND U545 ( .A(S), .B(n364), .Z(n363) );
  XOR U546 ( .A(B[167]), .B(A[167]), .Z(n364) );
  XOR U547 ( .A(A[166]), .B(n365), .Z(O[166]) );
  AND U548 ( .A(S), .B(n366), .Z(n365) );
  XOR U549 ( .A(B[166]), .B(A[166]), .Z(n366) );
  XOR U550 ( .A(A[165]), .B(n367), .Z(O[165]) );
  AND U551 ( .A(S), .B(n368), .Z(n367) );
  XOR U552 ( .A(B[165]), .B(A[165]), .Z(n368) );
  XOR U553 ( .A(A[164]), .B(n369), .Z(O[164]) );
  AND U554 ( .A(S), .B(n370), .Z(n369) );
  XOR U555 ( .A(B[164]), .B(A[164]), .Z(n370) );
  XOR U556 ( .A(A[163]), .B(n371), .Z(O[163]) );
  AND U557 ( .A(S), .B(n372), .Z(n371) );
  XOR U558 ( .A(B[163]), .B(A[163]), .Z(n372) );
  XOR U559 ( .A(A[162]), .B(n373), .Z(O[162]) );
  AND U560 ( .A(S), .B(n374), .Z(n373) );
  XOR U561 ( .A(B[162]), .B(A[162]), .Z(n374) );
  XOR U562 ( .A(A[161]), .B(n375), .Z(O[161]) );
  AND U563 ( .A(S), .B(n376), .Z(n375) );
  XOR U564 ( .A(B[161]), .B(A[161]), .Z(n376) );
  XOR U565 ( .A(A[160]), .B(n377), .Z(O[160]) );
  AND U566 ( .A(S), .B(n378), .Z(n377) );
  XOR U567 ( .A(B[160]), .B(A[160]), .Z(n378) );
  XOR U568 ( .A(A[15]), .B(n379), .Z(O[15]) );
  AND U569 ( .A(S), .B(n380), .Z(n379) );
  XOR U570 ( .A(B[15]), .B(A[15]), .Z(n380) );
  XOR U571 ( .A(A[159]), .B(n381), .Z(O[159]) );
  AND U572 ( .A(S), .B(n382), .Z(n381) );
  XOR U573 ( .A(B[159]), .B(A[159]), .Z(n382) );
  XOR U574 ( .A(A[158]), .B(n383), .Z(O[158]) );
  AND U575 ( .A(S), .B(n384), .Z(n383) );
  XOR U576 ( .A(B[158]), .B(A[158]), .Z(n384) );
  XOR U577 ( .A(A[157]), .B(n385), .Z(O[157]) );
  AND U578 ( .A(S), .B(n386), .Z(n385) );
  XOR U579 ( .A(B[157]), .B(A[157]), .Z(n386) );
  XOR U580 ( .A(A[156]), .B(n387), .Z(O[156]) );
  AND U581 ( .A(S), .B(n388), .Z(n387) );
  XOR U582 ( .A(B[156]), .B(A[156]), .Z(n388) );
  XOR U583 ( .A(A[155]), .B(n389), .Z(O[155]) );
  AND U584 ( .A(S), .B(n390), .Z(n389) );
  XOR U585 ( .A(B[155]), .B(A[155]), .Z(n390) );
  XOR U586 ( .A(A[154]), .B(n391), .Z(O[154]) );
  AND U587 ( .A(S), .B(n392), .Z(n391) );
  XOR U588 ( .A(B[154]), .B(A[154]), .Z(n392) );
  XOR U589 ( .A(A[153]), .B(n393), .Z(O[153]) );
  AND U590 ( .A(S), .B(n394), .Z(n393) );
  XOR U591 ( .A(B[153]), .B(A[153]), .Z(n394) );
  XOR U592 ( .A(A[152]), .B(n395), .Z(O[152]) );
  AND U593 ( .A(S), .B(n396), .Z(n395) );
  XOR U594 ( .A(B[152]), .B(A[152]), .Z(n396) );
  XOR U595 ( .A(A[151]), .B(n397), .Z(O[151]) );
  AND U596 ( .A(S), .B(n398), .Z(n397) );
  XOR U597 ( .A(B[151]), .B(A[151]), .Z(n398) );
  XOR U598 ( .A(A[150]), .B(n399), .Z(O[150]) );
  AND U599 ( .A(S), .B(n400), .Z(n399) );
  XOR U600 ( .A(B[150]), .B(A[150]), .Z(n400) );
  XOR U601 ( .A(A[14]), .B(n401), .Z(O[14]) );
  AND U602 ( .A(S), .B(n402), .Z(n401) );
  XOR U603 ( .A(B[14]), .B(A[14]), .Z(n402) );
  XOR U604 ( .A(A[149]), .B(n403), .Z(O[149]) );
  AND U605 ( .A(S), .B(n404), .Z(n403) );
  XOR U606 ( .A(B[149]), .B(A[149]), .Z(n404) );
  XOR U607 ( .A(A[148]), .B(n405), .Z(O[148]) );
  AND U608 ( .A(S), .B(n406), .Z(n405) );
  XOR U609 ( .A(B[148]), .B(A[148]), .Z(n406) );
  XOR U610 ( .A(A[147]), .B(n407), .Z(O[147]) );
  AND U611 ( .A(S), .B(n408), .Z(n407) );
  XOR U612 ( .A(B[147]), .B(A[147]), .Z(n408) );
  XOR U613 ( .A(A[146]), .B(n409), .Z(O[146]) );
  AND U614 ( .A(S), .B(n410), .Z(n409) );
  XOR U615 ( .A(B[146]), .B(A[146]), .Z(n410) );
  XOR U616 ( .A(A[145]), .B(n411), .Z(O[145]) );
  AND U617 ( .A(S), .B(n412), .Z(n411) );
  XOR U618 ( .A(B[145]), .B(A[145]), .Z(n412) );
  XOR U619 ( .A(A[144]), .B(n413), .Z(O[144]) );
  AND U620 ( .A(S), .B(n414), .Z(n413) );
  XOR U621 ( .A(B[144]), .B(A[144]), .Z(n414) );
  XOR U622 ( .A(A[143]), .B(n415), .Z(O[143]) );
  AND U623 ( .A(S), .B(n416), .Z(n415) );
  XOR U624 ( .A(B[143]), .B(A[143]), .Z(n416) );
  XOR U625 ( .A(A[142]), .B(n417), .Z(O[142]) );
  AND U626 ( .A(S), .B(n418), .Z(n417) );
  XOR U627 ( .A(B[142]), .B(A[142]), .Z(n418) );
  XOR U628 ( .A(A[141]), .B(n419), .Z(O[141]) );
  AND U629 ( .A(S), .B(n420), .Z(n419) );
  XOR U630 ( .A(B[141]), .B(A[141]), .Z(n420) );
  XOR U631 ( .A(A[140]), .B(n421), .Z(O[140]) );
  AND U632 ( .A(S), .B(n422), .Z(n421) );
  XOR U633 ( .A(B[140]), .B(A[140]), .Z(n422) );
  XOR U634 ( .A(A[13]), .B(n423), .Z(O[13]) );
  AND U635 ( .A(S), .B(n424), .Z(n423) );
  XOR U636 ( .A(B[13]), .B(A[13]), .Z(n424) );
  XOR U637 ( .A(A[139]), .B(n425), .Z(O[139]) );
  AND U638 ( .A(S), .B(n426), .Z(n425) );
  XOR U639 ( .A(B[139]), .B(A[139]), .Z(n426) );
  XOR U640 ( .A(A[138]), .B(n427), .Z(O[138]) );
  AND U641 ( .A(S), .B(n428), .Z(n427) );
  XOR U642 ( .A(B[138]), .B(A[138]), .Z(n428) );
  XOR U643 ( .A(A[137]), .B(n429), .Z(O[137]) );
  AND U644 ( .A(S), .B(n430), .Z(n429) );
  XOR U645 ( .A(B[137]), .B(A[137]), .Z(n430) );
  XOR U646 ( .A(A[136]), .B(n431), .Z(O[136]) );
  AND U647 ( .A(S), .B(n432), .Z(n431) );
  XOR U648 ( .A(B[136]), .B(A[136]), .Z(n432) );
  XOR U649 ( .A(A[135]), .B(n433), .Z(O[135]) );
  AND U650 ( .A(S), .B(n434), .Z(n433) );
  XOR U651 ( .A(B[135]), .B(A[135]), .Z(n434) );
  XOR U652 ( .A(A[134]), .B(n435), .Z(O[134]) );
  AND U653 ( .A(S), .B(n436), .Z(n435) );
  XOR U654 ( .A(B[134]), .B(A[134]), .Z(n436) );
  XOR U655 ( .A(A[133]), .B(n437), .Z(O[133]) );
  AND U656 ( .A(S), .B(n438), .Z(n437) );
  XOR U657 ( .A(B[133]), .B(A[133]), .Z(n438) );
  XOR U658 ( .A(A[132]), .B(n439), .Z(O[132]) );
  AND U659 ( .A(S), .B(n440), .Z(n439) );
  XOR U660 ( .A(B[132]), .B(A[132]), .Z(n440) );
  XOR U661 ( .A(A[131]), .B(n441), .Z(O[131]) );
  AND U662 ( .A(S), .B(n442), .Z(n441) );
  XOR U663 ( .A(B[131]), .B(A[131]), .Z(n442) );
  XOR U664 ( .A(A[130]), .B(n443), .Z(O[130]) );
  AND U665 ( .A(S), .B(n444), .Z(n443) );
  XOR U666 ( .A(B[130]), .B(A[130]), .Z(n444) );
  XOR U667 ( .A(A[12]), .B(n445), .Z(O[12]) );
  AND U668 ( .A(S), .B(n446), .Z(n445) );
  XOR U669 ( .A(B[12]), .B(A[12]), .Z(n446) );
  XOR U670 ( .A(A[129]), .B(n447), .Z(O[129]) );
  AND U671 ( .A(S), .B(n448), .Z(n447) );
  XOR U672 ( .A(B[129]), .B(A[129]), .Z(n448) );
  XOR U673 ( .A(A[128]), .B(n449), .Z(O[128]) );
  AND U674 ( .A(S), .B(n450), .Z(n449) );
  XOR U675 ( .A(B[128]), .B(A[128]), .Z(n450) );
  XOR U676 ( .A(A[127]), .B(n451), .Z(O[127]) );
  AND U677 ( .A(S), .B(n452), .Z(n451) );
  XOR U678 ( .A(B[127]), .B(A[127]), .Z(n452) );
  XOR U679 ( .A(A[126]), .B(n453), .Z(O[126]) );
  AND U680 ( .A(S), .B(n454), .Z(n453) );
  XOR U681 ( .A(B[126]), .B(A[126]), .Z(n454) );
  XOR U682 ( .A(A[125]), .B(n455), .Z(O[125]) );
  AND U683 ( .A(S), .B(n456), .Z(n455) );
  XOR U684 ( .A(B[125]), .B(A[125]), .Z(n456) );
  XOR U685 ( .A(A[124]), .B(n457), .Z(O[124]) );
  AND U686 ( .A(S), .B(n458), .Z(n457) );
  XOR U687 ( .A(B[124]), .B(A[124]), .Z(n458) );
  XOR U688 ( .A(A[123]), .B(n459), .Z(O[123]) );
  AND U689 ( .A(S), .B(n460), .Z(n459) );
  XOR U690 ( .A(B[123]), .B(A[123]), .Z(n460) );
  XOR U691 ( .A(A[122]), .B(n461), .Z(O[122]) );
  AND U692 ( .A(S), .B(n462), .Z(n461) );
  XOR U693 ( .A(B[122]), .B(A[122]), .Z(n462) );
  XOR U694 ( .A(A[121]), .B(n463), .Z(O[121]) );
  AND U695 ( .A(S), .B(n464), .Z(n463) );
  XOR U696 ( .A(B[121]), .B(A[121]), .Z(n464) );
  XOR U697 ( .A(A[120]), .B(n465), .Z(O[120]) );
  AND U698 ( .A(S), .B(n466), .Z(n465) );
  XOR U699 ( .A(B[120]), .B(A[120]), .Z(n466) );
  XOR U700 ( .A(A[11]), .B(n467), .Z(O[11]) );
  AND U701 ( .A(S), .B(n468), .Z(n467) );
  XOR U702 ( .A(B[11]), .B(A[11]), .Z(n468) );
  XOR U703 ( .A(A[119]), .B(n469), .Z(O[119]) );
  AND U704 ( .A(S), .B(n470), .Z(n469) );
  XOR U705 ( .A(B[119]), .B(A[119]), .Z(n470) );
  XOR U706 ( .A(A[118]), .B(n471), .Z(O[118]) );
  AND U707 ( .A(S), .B(n472), .Z(n471) );
  XOR U708 ( .A(B[118]), .B(A[118]), .Z(n472) );
  XOR U709 ( .A(A[117]), .B(n473), .Z(O[117]) );
  AND U710 ( .A(S), .B(n474), .Z(n473) );
  XOR U711 ( .A(B[117]), .B(A[117]), .Z(n474) );
  XOR U712 ( .A(A[116]), .B(n475), .Z(O[116]) );
  AND U713 ( .A(S), .B(n476), .Z(n475) );
  XOR U714 ( .A(B[116]), .B(A[116]), .Z(n476) );
  XOR U715 ( .A(A[115]), .B(n477), .Z(O[115]) );
  AND U716 ( .A(S), .B(n478), .Z(n477) );
  XOR U717 ( .A(B[115]), .B(A[115]), .Z(n478) );
  XOR U718 ( .A(A[114]), .B(n479), .Z(O[114]) );
  AND U719 ( .A(S), .B(n480), .Z(n479) );
  XOR U720 ( .A(B[114]), .B(A[114]), .Z(n480) );
  XOR U721 ( .A(A[113]), .B(n481), .Z(O[113]) );
  AND U722 ( .A(S), .B(n482), .Z(n481) );
  XOR U723 ( .A(B[113]), .B(A[113]), .Z(n482) );
  XOR U724 ( .A(A[112]), .B(n483), .Z(O[112]) );
  AND U725 ( .A(S), .B(n484), .Z(n483) );
  XOR U726 ( .A(B[112]), .B(A[112]), .Z(n484) );
  XOR U727 ( .A(A[111]), .B(n485), .Z(O[111]) );
  AND U728 ( .A(S), .B(n486), .Z(n485) );
  XOR U729 ( .A(B[111]), .B(A[111]), .Z(n486) );
  XOR U730 ( .A(A[110]), .B(n487), .Z(O[110]) );
  AND U731 ( .A(S), .B(n488), .Z(n487) );
  XOR U732 ( .A(B[110]), .B(A[110]), .Z(n488) );
  XOR U733 ( .A(A[10]), .B(n489), .Z(O[10]) );
  AND U734 ( .A(S), .B(n490), .Z(n489) );
  XOR U735 ( .A(B[10]), .B(A[10]), .Z(n490) );
  XOR U736 ( .A(A[109]), .B(n491), .Z(O[109]) );
  AND U737 ( .A(S), .B(n492), .Z(n491) );
  XOR U738 ( .A(B[109]), .B(A[109]), .Z(n492) );
  XOR U739 ( .A(A[108]), .B(n493), .Z(O[108]) );
  AND U740 ( .A(S), .B(n494), .Z(n493) );
  XOR U741 ( .A(B[108]), .B(A[108]), .Z(n494) );
  XOR U742 ( .A(A[107]), .B(n495), .Z(O[107]) );
  AND U743 ( .A(S), .B(n496), .Z(n495) );
  XOR U744 ( .A(B[107]), .B(A[107]), .Z(n496) );
  XOR U745 ( .A(A[106]), .B(n497), .Z(O[106]) );
  AND U746 ( .A(S), .B(n498), .Z(n497) );
  XOR U747 ( .A(B[106]), .B(A[106]), .Z(n498) );
  XOR U748 ( .A(A[105]), .B(n499), .Z(O[105]) );
  AND U749 ( .A(S), .B(n500), .Z(n499) );
  XOR U750 ( .A(B[105]), .B(A[105]), .Z(n500) );
  XOR U751 ( .A(A[104]), .B(n501), .Z(O[104]) );
  AND U752 ( .A(S), .B(n502), .Z(n501) );
  XOR U753 ( .A(B[104]), .B(A[104]), .Z(n502) );
  XOR U754 ( .A(A[103]), .B(n503), .Z(O[103]) );
  AND U755 ( .A(S), .B(n504), .Z(n503) );
  XOR U756 ( .A(B[103]), .B(A[103]), .Z(n504) );
  XOR U757 ( .A(A[102]), .B(n505), .Z(O[102]) );
  AND U758 ( .A(S), .B(n506), .Z(n505) );
  XOR U759 ( .A(B[102]), .B(A[102]), .Z(n506) );
  XOR U760 ( .A(A[101]), .B(n507), .Z(O[101]) );
  AND U761 ( .A(S), .B(n508), .Z(n507) );
  XOR U762 ( .A(B[101]), .B(A[101]), .Z(n508) );
  XOR U763 ( .A(A[100]), .B(n509), .Z(O[100]) );
  AND U764 ( .A(S), .B(n510), .Z(n509) );
  XOR U765 ( .A(B[100]), .B(A[100]), .Z(n510) );
  XOR U766 ( .A(A[0]), .B(n511), .Z(O[0]) );
  AND U767 ( .A(S), .B(n512), .Z(n511) );
  XOR U768 ( .A(B[0]), .B(A[0]), .Z(n512) );
endmodule


module MUX_N256_5 ( A, B, S, O );
  input [255:0] A;
  input [255:0] B;
  output [255:0] O;
  input S;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510;

  XOR U1 ( .A(B[8]), .B(n1), .Z(O[9]) );
  AND U2 ( .A(S), .B(n2), .Z(n1) );
  XOR U3 ( .A(B[9]), .B(B[8]), .Z(n2) );
  XOR U4 ( .A(B[98]), .B(n3), .Z(O[99]) );
  AND U5 ( .A(S), .B(n4), .Z(n3) );
  XOR U6 ( .A(B[99]), .B(B[98]), .Z(n4) );
  XOR U7 ( .A(B[97]), .B(n5), .Z(O[98]) );
  AND U8 ( .A(S), .B(n6), .Z(n5) );
  XOR U9 ( .A(B[98]), .B(B[97]), .Z(n6) );
  XOR U10 ( .A(B[96]), .B(n7), .Z(O[97]) );
  AND U11 ( .A(S), .B(n8), .Z(n7) );
  XOR U12 ( .A(B[97]), .B(B[96]), .Z(n8) );
  XOR U13 ( .A(B[95]), .B(n9), .Z(O[96]) );
  AND U14 ( .A(S), .B(n10), .Z(n9) );
  XOR U15 ( .A(B[96]), .B(B[95]), .Z(n10) );
  XOR U16 ( .A(B[94]), .B(n11), .Z(O[95]) );
  AND U17 ( .A(S), .B(n12), .Z(n11) );
  XOR U18 ( .A(B[95]), .B(B[94]), .Z(n12) );
  XOR U19 ( .A(B[93]), .B(n13), .Z(O[94]) );
  AND U20 ( .A(S), .B(n14), .Z(n13) );
  XOR U21 ( .A(B[94]), .B(B[93]), .Z(n14) );
  XOR U22 ( .A(B[92]), .B(n15), .Z(O[93]) );
  AND U23 ( .A(S), .B(n16), .Z(n15) );
  XOR U24 ( .A(B[93]), .B(B[92]), .Z(n16) );
  XOR U25 ( .A(B[91]), .B(n17), .Z(O[92]) );
  AND U26 ( .A(S), .B(n18), .Z(n17) );
  XOR U27 ( .A(B[92]), .B(B[91]), .Z(n18) );
  XOR U28 ( .A(B[90]), .B(n19), .Z(O[91]) );
  AND U29 ( .A(S), .B(n20), .Z(n19) );
  XOR U30 ( .A(B[91]), .B(B[90]), .Z(n20) );
  XOR U31 ( .A(B[89]), .B(n21), .Z(O[90]) );
  AND U32 ( .A(S), .B(n22), .Z(n21) );
  XOR U33 ( .A(B[90]), .B(B[89]), .Z(n22) );
  XOR U34 ( .A(B[7]), .B(n23), .Z(O[8]) );
  AND U35 ( .A(S), .B(n24), .Z(n23) );
  XOR U36 ( .A(B[8]), .B(B[7]), .Z(n24) );
  XOR U37 ( .A(B[88]), .B(n25), .Z(O[89]) );
  AND U38 ( .A(S), .B(n26), .Z(n25) );
  XOR U39 ( .A(B[89]), .B(B[88]), .Z(n26) );
  XOR U40 ( .A(B[87]), .B(n27), .Z(O[88]) );
  AND U41 ( .A(S), .B(n28), .Z(n27) );
  XOR U42 ( .A(B[88]), .B(B[87]), .Z(n28) );
  XOR U43 ( .A(B[86]), .B(n29), .Z(O[87]) );
  AND U44 ( .A(S), .B(n30), .Z(n29) );
  XOR U45 ( .A(B[87]), .B(B[86]), .Z(n30) );
  XOR U46 ( .A(B[85]), .B(n31), .Z(O[86]) );
  AND U47 ( .A(S), .B(n32), .Z(n31) );
  XOR U48 ( .A(B[86]), .B(B[85]), .Z(n32) );
  XOR U49 ( .A(B[84]), .B(n33), .Z(O[85]) );
  AND U50 ( .A(S), .B(n34), .Z(n33) );
  XOR U51 ( .A(B[85]), .B(B[84]), .Z(n34) );
  XOR U52 ( .A(B[83]), .B(n35), .Z(O[84]) );
  AND U53 ( .A(S), .B(n36), .Z(n35) );
  XOR U54 ( .A(B[84]), .B(B[83]), .Z(n36) );
  XOR U55 ( .A(B[82]), .B(n37), .Z(O[83]) );
  AND U56 ( .A(S), .B(n38), .Z(n37) );
  XOR U57 ( .A(B[83]), .B(B[82]), .Z(n38) );
  XOR U58 ( .A(B[81]), .B(n39), .Z(O[82]) );
  AND U59 ( .A(S), .B(n40), .Z(n39) );
  XOR U60 ( .A(B[82]), .B(B[81]), .Z(n40) );
  XOR U61 ( .A(B[80]), .B(n41), .Z(O[81]) );
  AND U62 ( .A(S), .B(n42), .Z(n41) );
  XOR U63 ( .A(B[81]), .B(B[80]), .Z(n42) );
  XOR U64 ( .A(B[79]), .B(n43), .Z(O[80]) );
  AND U65 ( .A(S), .B(n44), .Z(n43) );
  XOR U66 ( .A(B[80]), .B(B[79]), .Z(n44) );
  XOR U67 ( .A(B[6]), .B(n45), .Z(O[7]) );
  AND U68 ( .A(S), .B(n46), .Z(n45) );
  XOR U69 ( .A(B[7]), .B(B[6]), .Z(n46) );
  XOR U70 ( .A(B[78]), .B(n47), .Z(O[79]) );
  AND U71 ( .A(S), .B(n48), .Z(n47) );
  XOR U72 ( .A(B[79]), .B(B[78]), .Z(n48) );
  XOR U73 ( .A(B[77]), .B(n49), .Z(O[78]) );
  AND U74 ( .A(S), .B(n50), .Z(n49) );
  XOR U75 ( .A(B[78]), .B(B[77]), .Z(n50) );
  XOR U76 ( .A(B[76]), .B(n51), .Z(O[77]) );
  AND U77 ( .A(S), .B(n52), .Z(n51) );
  XOR U78 ( .A(B[77]), .B(B[76]), .Z(n52) );
  XOR U79 ( .A(B[75]), .B(n53), .Z(O[76]) );
  AND U80 ( .A(S), .B(n54), .Z(n53) );
  XOR U81 ( .A(B[76]), .B(B[75]), .Z(n54) );
  XOR U82 ( .A(B[74]), .B(n55), .Z(O[75]) );
  AND U83 ( .A(S), .B(n56), .Z(n55) );
  XOR U84 ( .A(B[75]), .B(B[74]), .Z(n56) );
  XOR U85 ( .A(B[73]), .B(n57), .Z(O[74]) );
  AND U86 ( .A(S), .B(n58), .Z(n57) );
  XOR U87 ( .A(B[74]), .B(B[73]), .Z(n58) );
  XOR U88 ( .A(B[72]), .B(n59), .Z(O[73]) );
  AND U89 ( .A(S), .B(n60), .Z(n59) );
  XOR U90 ( .A(B[73]), .B(B[72]), .Z(n60) );
  XOR U91 ( .A(B[71]), .B(n61), .Z(O[72]) );
  AND U92 ( .A(S), .B(n62), .Z(n61) );
  XOR U93 ( .A(B[72]), .B(B[71]), .Z(n62) );
  XOR U94 ( .A(B[70]), .B(n63), .Z(O[71]) );
  AND U95 ( .A(S), .B(n64), .Z(n63) );
  XOR U96 ( .A(B[71]), .B(B[70]), .Z(n64) );
  XOR U97 ( .A(B[69]), .B(n65), .Z(O[70]) );
  AND U98 ( .A(S), .B(n66), .Z(n65) );
  XOR U99 ( .A(B[70]), .B(B[69]), .Z(n66) );
  XOR U100 ( .A(B[5]), .B(n67), .Z(O[6]) );
  AND U101 ( .A(S), .B(n68), .Z(n67) );
  XOR U102 ( .A(B[6]), .B(B[5]), .Z(n68) );
  XOR U103 ( .A(B[68]), .B(n69), .Z(O[69]) );
  AND U104 ( .A(S), .B(n70), .Z(n69) );
  XOR U105 ( .A(B[69]), .B(B[68]), .Z(n70) );
  XOR U106 ( .A(B[67]), .B(n71), .Z(O[68]) );
  AND U107 ( .A(S), .B(n72), .Z(n71) );
  XOR U108 ( .A(B[68]), .B(B[67]), .Z(n72) );
  XOR U109 ( .A(B[66]), .B(n73), .Z(O[67]) );
  AND U110 ( .A(S), .B(n74), .Z(n73) );
  XOR U111 ( .A(B[67]), .B(B[66]), .Z(n74) );
  XOR U112 ( .A(B[65]), .B(n75), .Z(O[66]) );
  AND U113 ( .A(S), .B(n76), .Z(n75) );
  XOR U114 ( .A(B[66]), .B(B[65]), .Z(n76) );
  XOR U115 ( .A(B[64]), .B(n77), .Z(O[65]) );
  AND U116 ( .A(S), .B(n78), .Z(n77) );
  XOR U117 ( .A(B[65]), .B(B[64]), .Z(n78) );
  XOR U118 ( .A(B[63]), .B(n79), .Z(O[64]) );
  AND U119 ( .A(S), .B(n80), .Z(n79) );
  XOR U120 ( .A(B[64]), .B(B[63]), .Z(n80) );
  XOR U121 ( .A(B[62]), .B(n81), .Z(O[63]) );
  AND U122 ( .A(S), .B(n82), .Z(n81) );
  XOR U123 ( .A(B[63]), .B(B[62]), .Z(n82) );
  XOR U124 ( .A(B[61]), .B(n83), .Z(O[62]) );
  AND U125 ( .A(S), .B(n84), .Z(n83) );
  XOR U126 ( .A(B[62]), .B(B[61]), .Z(n84) );
  XOR U127 ( .A(B[60]), .B(n85), .Z(O[61]) );
  AND U128 ( .A(S), .B(n86), .Z(n85) );
  XOR U129 ( .A(B[61]), .B(B[60]), .Z(n86) );
  XOR U130 ( .A(B[59]), .B(n87), .Z(O[60]) );
  AND U131 ( .A(S), .B(n88), .Z(n87) );
  XOR U132 ( .A(B[60]), .B(B[59]), .Z(n88) );
  XOR U133 ( .A(B[4]), .B(n89), .Z(O[5]) );
  AND U134 ( .A(S), .B(n90), .Z(n89) );
  XOR U135 ( .A(B[5]), .B(B[4]), .Z(n90) );
  XOR U136 ( .A(B[58]), .B(n91), .Z(O[59]) );
  AND U137 ( .A(S), .B(n92), .Z(n91) );
  XOR U138 ( .A(B[59]), .B(B[58]), .Z(n92) );
  XOR U139 ( .A(B[57]), .B(n93), .Z(O[58]) );
  AND U140 ( .A(S), .B(n94), .Z(n93) );
  XOR U141 ( .A(B[58]), .B(B[57]), .Z(n94) );
  XOR U142 ( .A(B[56]), .B(n95), .Z(O[57]) );
  AND U143 ( .A(S), .B(n96), .Z(n95) );
  XOR U144 ( .A(B[57]), .B(B[56]), .Z(n96) );
  XOR U145 ( .A(B[55]), .B(n97), .Z(O[56]) );
  AND U146 ( .A(S), .B(n98), .Z(n97) );
  XOR U147 ( .A(B[56]), .B(B[55]), .Z(n98) );
  XOR U148 ( .A(B[54]), .B(n99), .Z(O[55]) );
  AND U149 ( .A(S), .B(n100), .Z(n99) );
  XOR U150 ( .A(B[55]), .B(B[54]), .Z(n100) );
  XOR U151 ( .A(B[53]), .B(n101), .Z(O[54]) );
  AND U152 ( .A(S), .B(n102), .Z(n101) );
  XOR U153 ( .A(B[54]), .B(B[53]), .Z(n102) );
  XOR U154 ( .A(B[52]), .B(n103), .Z(O[53]) );
  AND U155 ( .A(S), .B(n104), .Z(n103) );
  XOR U156 ( .A(B[53]), .B(B[52]), .Z(n104) );
  XOR U157 ( .A(B[51]), .B(n105), .Z(O[52]) );
  AND U158 ( .A(S), .B(n106), .Z(n105) );
  XOR U159 ( .A(B[52]), .B(B[51]), .Z(n106) );
  XOR U160 ( .A(B[50]), .B(n107), .Z(O[51]) );
  AND U161 ( .A(S), .B(n108), .Z(n107) );
  XOR U162 ( .A(B[51]), .B(B[50]), .Z(n108) );
  XOR U163 ( .A(B[49]), .B(n109), .Z(O[50]) );
  AND U164 ( .A(S), .B(n110), .Z(n109) );
  XOR U165 ( .A(B[50]), .B(B[49]), .Z(n110) );
  XOR U166 ( .A(B[3]), .B(n111), .Z(O[4]) );
  AND U167 ( .A(S), .B(n112), .Z(n111) );
  XOR U168 ( .A(B[4]), .B(B[3]), .Z(n112) );
  XOR U169 ( .A(B[48]), .B(n113), .Z(O[49]) );
  AND U170 ( .A(S), .B(n114), .Z(n113) );
  XOR U171 ( .A(B[49]), .B(B[48]), .Z(n114) );
  XOR U172 ( .A(B[47]), .B(n115), .Z(O[48]) );
  AND U173 ( .A(S), .B(n116), .Z(n115) );
  XOR U174 ( .A(B[48]), .B(B[47]), .Z(n116) );
  XOR U175 ( .A(B[46]), .B(n117), .Z(O[47]) );
  AND U176 ( .A(S), .B(n118), .Z(n117) );
  XOR U177 ( .A(B[47]), .B(B[46]), .Z(n118) );
  XOR U178 ( .A(B[45]), .B(n119), .Z(O[46]) );
  AND U179 ( .A(S), .B(n120), .Z(n119) );
  XOR U180 ( .A(B[46]), .B(B[45]), .Z(n120) );
  XOR U181 ( .A(B[44]), .B(n121), .Z(O[45]) );
  AND U182 ( .A(S), .B(n122), .Z(n121) );
  XOR U183 ( .A(B[45]), .B(B[44]), .Z(n122) );
  XOR U184 ( .A(B[43]), .B(n123), .Z(O[44]) );
  AND U185 ( .A(S), .B(n124), .Z(n123) );
  XOR U186 ( .A(B[44]), .B(B[43]), .Z(n124) );
  XOR U187 ( .A(B[42]), .B(n125), .Z(O[43]) );
  AND U188 ( .A(S), .B(n126), .Z(n125) );
  XOR U189 ( .A(B[43]), .B(B[42]), .Z(n126) );
  XOR U190 ( .A(B[41]), .B(n127), .Z(O[42]) );
  AND U191 ( .A(S), .B(n128), .Z(n127) );
  XOR U192 ( .A(B[42]), .B(B[41]), .Z(n128) );
  XOR U193 ( .A(B[40]), .B(n129), .Z(O[41]) );
  AND U194 ( .A(S), .B(n130), .Z(n129) );
  XOR U195 ( .A(B[41]), .B(B[40]), .Z(n130) );
  XOR U196 ( .A(B[39]), .B(n131), .Z(O[40]) );
  AND U197 ( .A(S), .B(n132), .Z(n131) );
  XOR U198 ( .A(B[40]), .B(B[39]), .Z(n132) );
  XOR U199 ( .A(B[2]), .B(n133), .Z(O[3]) );
  AND U200 ( .A(S), .B(n134), .Z(n133) );
  XOR U201 ( .A(B[3]), .B(B[2]), .Z(n134) );
  XOR U202 ( .A(B[38]), .B(n135), .Z(O[39]) );
  AND U203 ( .A(S), .B(n136), .Z(n135) );
  XOR U204 ( .A(B[39]), .B(B[38]), .Z(n136) );
  XOR U205 ( .A(B[37]), .B(n137), .Z(O[38]) );
  AND U206 ( .A(S), .B(n138), .Z(n137) );
  XOR U207 ( .A(B[38]), .B(B[37]), .Z(n138) );
  XOR U208 ( .A(B[36]), .B(n139), .Z(O[37]) );
  AND U209 ( .A(S), .B(n140), .Z(n139) );
  XOR U210 ( .A(B[37]), .B(B[36]), .Z(n140) );
  XOR U211 ( .A(B[35]), .B(n141), .Z(O[36]) );
  AND U212 ( .A(S), .B(n142), .Z(n141) );
  XOR U213 ( .A(B[36]), .B(B[35]), .Z(n142) );
  XOR U214 ( .A(B[34]), .B(n143), .Z(O[35]) );
  AND U215 ( .A(S), .B(n144), .Z(n143) );
  XOR U216 ( .A(B[35]), .B(B[34]), .Z(n144) );
  XOR U217 ( .A(B[33]), .B(n145), .Z(O[34]) );
  AND U218 ( .A(S), .B(n146), .Z(n145) );
  XOR U219 ( .A(B[34]), .B(B[33]), .Z(n146) );
  XOR U220 ( .A(B[32]), .B(n147), .Z(O[33]) );
  AND U221 ( .A(S), .B(n148), .Z(n147) );
  XOR U222 ( .A(B[33]), .B(B[32]), .Z(n148) );
  XOR U223 ( .A(B[31]), .B(n149), .Z(O[32]) );
  AND U224 ( .A(S), .B(n150), .Z(n149) );
  XOR U225 ( .A(B[32]), .B(B[31]), .Z(n150) );
  XOR U226 ( .A(B[30]), .B(n151), .Z(O[31]) );
  AND U227 ( .A(S), .B(n152), .Z(n151) );
  XOR U228 ( .A(B[31]), .B(B[30]), .Z(n152) );
  XOR U229 ( .A(B[29]), .B(n153), .Z(O[30]) );
  AND U230 ( .A(S), .B(n154), .Z(n153) );
  XOR U231 ( .A(B[30]), .B(B[29]), .Z(n154) );
  XOR U232 ( .A(B[1]), .B(n155), .Z(O[2]) );
  AND U233 ( .A(S), .B(n156), .Z(n155) );
  XOR U234 ( .A(B[2]), .B(B[1]), .Z(n156) );
  XOR U235 ( .A(B[28]), .B(n157), .Z(O[29]) );
  AND U236 ( .A(S), .B(n158), .Z(n157) );
  XOR U237 ( .A(B[29]), .B(B[28]), .Z(n158) );
  XOR U238 ( .A(B[27]), .B(n159), .Z(O[28]) );
  AND U239 ( .A(S), .B(n160), .Z(n159) );
  XOR U240 ( .A(B[28]), .B(B[27]), .Z(n160) );
  XOR U241 ( .A(B[26]), .B(n161), .Z(O[27]) );
  AND U242 ( .A(S), .B(n162), .Z(n161) );
  XOR U243 ( .A(B[27]), .B(B[26]), .Z(n162) );
  XOR U244 ( .A(B[25]), .B(n163), .Z(O[26]) );
  AND U245 ( .A(S), .B(n164), .Z(n163) );
  XOR U246 ( .A(B[26]), .B(B[25]), .Z(n164) );
  XOR U247 ( .A(B[24]), .B(n165), .Z(O[25]) );
  AND U248 ( .A(S), .B(n166), .Z(n165) );
  XOR U249 ( .A(B[25]), .B(B[24]), .Z(n166) );
  XOR U250 ( .A(B[254]), .B(n167), .Z(O[255]) );
  AND U251 ( .A(S), .B(n168), .Z(n167) );
  XOR U252 ( .A(B[255]), .B(B[254]), .Z(n168) );
  XOR U253 ( .A(B[253]), .B(n169), .Z(O[254]) );
  AND U254 ( .A(S), .B(n170), .Z(n169) );
  XOR U255 ( .A(B[254]), .B(B[253]), .Z(n170) );
  XOR U256 ( .A(B[252]), .B(n171), .Z(O[253]) );
  AND U257 ( .A(S), .B(n172), .Z(n171) );
  XOR U258 ( .A(B[253]), .B(B[252]), .Z(n172) );
  XOR U259 ( .A(B[251]), .B(n173), .Z(O[252]) );
  AND U260 ( .A(S), .B(n174), .Z(n173) );
  XOR U261 ( .A(B[252]), .B(B[251]), .Z(n174) );
  XOR U262 ( .A(B[250]), .B(n175), .Z(O[251]) );
  AND U263 ( .A(S), .B(n176), .Z(n175) );
  XOR U264 ( .A(B[251]), .B(B[250]), .Z(n176) );
  XOR U265 ( .A(B[249]), .B(n177), .Z(O[250]) );
  AND U266 ( .A(S), .B(n178), .Z(n177) );
  XOR U267 ( .A(B[250]), .B(B[249]), .Z(n178) );
  XOR U268 ( .A(B[23]), .B(n179), .Z(O[24]) );
  AND U269 ( .A(S), .B(n180), .Z(n179) );
  XOR U270 ( .A(B[24]), .B(B[23]), .Z(n180) );
  XOR U271 ( .A(B[248]), .B(n181), .Z(O[249]) );
  AND U272 ( .A(S), .B(n182), .Z(n181) );
  XOR U273 ( .A(B[249]), .B(B[248]), .Z(n182) );
  XOR U274 ( .A(B[247]), .B(n183), .Z(O[248]) );
  AND U275 ( .A(S), .B(n184), .Z(n183) );
  XOR U276 ( .A(B[248]), .B(B[247]), .Z(n184) );
  XOR U277 ( .A(B[246]), .B(n185), .Z(O[247]) );
  AND U278 ( .A(S), .B(n186), .Z(n185) );
  XOR U279 ( .A(B[247]), .B(B[246]), .Z(n186) );
  XOR U280 ( .A(B[245]), .B(n187), .Z(O[246]) );
  AND U281 ( .A(S), .B(n188), .Z(n187) );
  XOR U282 ( .A(B[246]), .B(B[245]), .Z(n188) );
  XOR U283 ( .A(B[244]), .B(n189), .Z(O[245]) );
  AND U284 ( .A(S), .B(n190), .Z(n189) );
  XOR U285 ( .A(B[245]), .B(B[244]), .Z(n190) );
  XOR U286 ( .A(B[243]), .B(n191), .Z(O[244]) );
  AND U287 ( .A(S), .B(n192), .Z(n191) );
  XOR U288 ( .A(B[244]), .B(B[243]), .Z(n192) );
  XOR U289 ( .A(B[242]), .B(n193), .Z(O[243]) );
  AND U290 ( .A(S), .B(n194), .Z(n193) );
  XOR U291 ( .A(B[243]), .B(B[242]), .Z(n194) );
  XOR U292 ( .A(B[241]), .B(n195), .Z(O[242]) );
  AND U293 ( .A(S), .B(n196), .Z(n195) );
  XOR U294 ( .A(B[242]), .B(B[241]), .Z(n196) );
  XOR U295 ( .A(B[240]), .B(n197), .Z(O[241]) );
  AND U296 ( .A(S), .B(n198), .Z(n197) );
  XOR U297 ( .A(B[241]), .B(B[240]), .Z(n198) );
  XOR U298 ( .A(B[239]), .B(n199), .Z(O[240]) );
  AND U299 ( .A(S), .B(n200), .Z(n199) );
  XOR U300 ( .A(B[240]), .B(B[239]), .Z(n200) );
  XOR U301 ( .A(B[22]), .B(n201), .Z(O[23]) );
  AND U302 ( .A(S), .B(n202), .Z(n201) );
  XOR U303 ( .A(B[23]), .B(B[22]), .Z(n202) );
  XOR U304 ( .A(B[238]), .B(n203), .Z(O[239]) );
  AND U305 ( .A(S), .B(n204), .Z(n203) );
  XOR U306 ( .A(B[239]), .B(B[238]), .Z(n204) );
  XOR U307 ( .A(B[237]), .B(n205), .Z(O[238]) );
  AND U308 ( .A(S), .B(n206), .Z(n205) );
  XOR U309 ( .A(B[238]), .B(B[237]), .Z(n206) );
  XOR U310 ( .A(B[236]), .B(n207), .Z(O[237]) );
  AND U311 ( .A(S), .B(n208), .Z(n207) );
  XOR U312 ( .A(B[237]), .B(B[236]), .Z(n208) );
  XOR U313 ( .A(B[235]), .B(n209), .Z(O[236]) );
  AND U314 ( .A(S), .B(n210), .Z(n209) );
  XOR U315 ( .A(B[236]), .B(B[235]), .Z(n210) );
  XOR U316 ( .A(B[234]), .B(n211), .Z(O[235]) );
  AND U317 ( .A(S), .B(n212), .Z(n211) );
  XOR U318 ( .A(B[235]), .B(B[234]), .Z(n212) );
  XOR U319 ( .A(B[233]), .B(n213), .Z(O[234]) );
  AND U320 ( .A(S), .B(n214), .Z(n213) );
  XOR U321 ( .A(B[234]), .B(B[233]), .Z(n214) );
  XOR U322 ( .A(B[232]), .B(n215), .Z(O[233]) );
  AND U323 ( .A(S), .B(n216), .Z(n215) );
  XOR U324 ( .A(B[233]), .B(B[232]), .Z(n216) );
  XOR U325 ( .A(B[231]), .B(n217), .Z(O[232]) );
  AND U326 ( .A(S), .B(n218), .Z(n217) );
  XOR U327 ( .A(B[232]), .B(B[231]), .Z(n218) );
  XOR U328 ( .A(B[230]), .B(n219), .Z(O[231]) );
  AND U329 ( .A(S), .B(n220), .Z(n219) );
  XOR U330 ( .A(B[231]), .B(B[230]), .Z(n220) );
  XOR U331 ( .A(B[229]), .B(n221), .Z(O[230]) );
  AND U332 ( .A(S), .B(n222), .Z(n221) );
  XOR U333 ( .A(B[230]), .B(B[229]), .Z(n222) );
  XOR U334 ( .A(B[21]), .B(n223), .Z(O[22]) );
  AND U335 ( .A(S), .B(n224), .Z(n223) );
  XOR U336 ( .A(B[22]), .B(B[21]), .Z(n224) );
  XOR U337 ( .A(B[228]), .B(n225), .Z(O[229]) );
  AND U338 ( .A(S), .B(n226), .Z(n225) );
  XOR U339 ( .A(B[229]), .B(B[228]), .Z(n226) );
  XOR U340 ( .A(B[227]), .B(n227), .Z(O[228]) );
  AND U341 ( .A(S), .B(n228), .Z(n227) );
  XOR U342 ( .A(B[228]), .B(B[227]), .Z(n228) );
  XOR U343 ( .A(B[226]), .B(n229), .Z(O[227]) );
  AND U344 ( .A(S), .B(n230), .Z(n229) );
  XOR U345 ( .A(B[227]), .B(B[226]), .Z(n230) );
  XOR U346 ( .A(B[225]), .B(n231), .Z(O[226]) );
  AND U347 ( .A(S), .B(n232), .Z(n231) );
  XOR U348 ( .A(B[226]), .B(B[225]), .Z(n232) );
  XOR U349 ( .A(B[224]), .B(n233), .Z(O[225]) );
  AND U350 ( .A(S), .B(n234), .Z(n233) );
  XOR U351 ( .A(B[225]), .B(B[224]), .Z(n234) );
  XOR U352 ( .A(B[223]), .B(n235), .Z(O[224]) );
  AND U353 ( .A(S), .B(n236), .Z(n235) );
  XOR U354 ( .A(B[224]), .B(B[223]), .Z(n236) );
  XOR U355 ( .A(B[222]), .B(n237), .Z(O[223]) );
  AND U356 ( .A(S), .B(n238), .Z(n237) );
  XOR U357 ( .A(B[223]), .B(B[222]), .Z(n238) );
  XOR U358 ( .A(B[221]), .B(n239), .Z(O[222]) );
  AND U359 ( .A(S), .B(n240), .Z(n239) );
  XOR U360 ( .A(B[222]), .B(B[221]), .Z(n240) );
  XOR U361 ( .A(B[220]), .B(n241), .Z(O[221]) );
  AND U362 ( .A(S), .B(n242), .Z(n241) );
  XOR U363 ( .A(B[221]), .B(B[220]), .Z(n242) );
  XOR U364 ( .A(B[219]), .B(n243), .Z(O[220]) );
  AND U365 ( .A(S), .B(n244), .Z(n243) );
  XOR U366 ( .A(B[220]), .B(B[219]), .Z(n244) );
  XOR U367 ( .A(B[20]), .B(n245), .Z(O[21]) );
  AND U368 ( .A(S), .B(n246), .Z(n245) );
  XOR U369 ( .A(B[21]), .B(B[20]), .Z(n246) );
  XOR U370 ( .A(B[218]), .B(n247), .Z(O[219]) );
  AND U371 ( .A(S), .B(n248), .Z(n247) );
  XOR U372 ( .A(B[219]), .B(B[218]), .Z(n248) );
  XOR U373 ( .A(B[217]), .B(n249), .Z(O[218]) );
  AND U374 ( .A(S), .B(n250), .Z(n249) );
  XOR U375 ( .A(B[218]), .B(B[217]), .Z(n250) );
  XOR U376 ( .A(B[216]), .B(n251), .Z(O[217]) );
  AND U377 ( .A(S), .B(n252), .Z(n251) );
  XOR U378 ( .A(B[217]), .B(B[216]), .Z(n252) );
  XOR U379 ( .A(B[215]), .B(n253), .Z(O[216]) );
  AND U380 ( .A(S), .B(n254), .Z(n253) );
  XOR U381 ( .A(B[216]), .B(B[215]), .Z(n254) );
  XOR U382 ( .A(B[214]), .B(n255), .Z(O[215]) );
  AND U383 ( .A(S), .B(n256), .Z(n255) );
  XOR U384 ( .A(B[215]), .B(B[214]), .Z(n256) );
  XOR U385 ( .A(B[213]), .B(n257), .Z(O[214]) );
  AND U386 ( .A(S), .B(n258), .Z(n257) );
  XOR U387 ( .A(B[214]), .B(B[213]), .Z(n258) );
  XOR U388 ( .A(B[212]), .B(n259), .Z(O[213]) );
  AND U389 ( .A(S), .B(n260), .Z(n259) );
  XOR U390 ( .A(B[213]), .B(B[212]), .Z(n260) );
  XOR U391 ( .A(B[211]), .B(n261), .Z(O[212]) );
  AND U392 ( .A(S), .B(n262), .Z(n261) );
  XOR U393 ( .A(B[212]), .B(B[211]), .Z(n262) );
  XOR U394 ( .A(B[210]), .B(n263), .Z(O[211]) );
  AND U395 ( .A(S), .B(n264), .Z(n263) );
  XOR U396 ( .A(B[211]), .B(B[210]), .Z(n264) );
  XOR U397 ( .A(B[209]), .B(n265), .Z(O[210]) );
  AND U398 ( .A(S), .B(n266), .Z(n265) );
  XOR U399 ( .A(B[210]), .B(B[209]), .Z(n266) );
  XOR U400 ( .A(B[19]), .B(n267), .Z(O[20]) );
  AND U401 ( .A(S), .B(n268), .Z(n267) );
  XOR U402 ( .A(B[20]), .B(B[19]), .Z(n268) );
  XOR U403 ( .A(B[208]), .B(n269), .Z(O[209]) );
  AND U404 ( .A(S), .B(n270), .Z(n269) );
  XOR U405 ( .A(B[209]), .B(B[208]), .Z(n270) );
  XOR U406 ( .A(B[207]), .B(n271), .Z(O[208]) );
  AND U407 ( .A(S), .B(n272), .Z(n271) );
  XOR U408 ( .A(B[208]), .B(B[207]), .Z(n272) );
  XOR U409 ( .A(B[206]), .B(n273), .Z(O[207]) );
  AND U410 ( .A(S), .B(n274), .Z(n273) );
  XOR U411 ( .A(B[207]), .B(B[206]), .Z(n274) );
  XOR U412 ( .A(B[205]), .B(n275), .Z(O[206]) );
  AND U413 ( .A(S), .B(n276), .Z(n275) );
  XOR U414 ( .A(B[206]), .B(B[205]), .Z(n276) );
  XOR U415 ( .A(B[204]), .B(n277), .Z(O[205]) );
  AND U416 ( .A(S), .B(n278), .Z(n277) );
  XOR U417 ( .A(B[205]), .B(B[204]), .Z(n278) );
  XOR U418 ( .A(B[203]), .B(n279), .Z(O[204]) );
  AND U419 ( .A(S), .B(n280), .Z(n279) );
  XOR U420 ( .A(B[204]), .B(B[203]), .Z(n280) );
  XOR U421 ( .A(B[202]), .B(n281), .Z(O[203]) );
  AND U422 ( .A(S), .B(n282), .Z(n281) );
  XOR U423 ( .A(B[203]), .B(B[202]), .Z(n282) );
  XOR U424 ( .A(B[201]), .B(n283), .Z(O[202]) );
  AND U425 ( .A(S), .B(n284), .Z(n283) );
  XOR U426 ( .A(B[202]), .B(B[201]), .Z(n284) );
  XOR U427 ( .A(B[200]), .B(n285), .Z(O[201]) );
  AND U428 ( .A(S), .B(n286), .Z(n285) );
  XOR U429 ( .A(B[201]), .B(B[200]), .Z(n286) );
  XOR U430 ( .A(B[199]), .B(n287), .Z(O[200]) );
  AND U431 ( .A(S), .B(n288), .Z(n287) );
  XOR U432 ( .A(B[200]), .B(B[199]), .Z(n288) );
  XOR U433 ( .A(B[0]), .B(n289), .Z(O[1]) );
  AND U434 ( .A(S), .B(n290), .Z(n289) );
  XOR U435 ( .A(B[1]), .B(B[0]), .Z(n290) );
  XOR U436 ( .A(B[18]), .B(n291), .Z(O[19]) );
  AND U437 ( .A(S), .B(n292), .Z(n291) );
  XOR U438 ( .A(B[19]), .B(B[18]), .Z(n292) );
  XOR U439 ( .A(B[198]), .B(n293), .Z(O[199]) );
  AND U440 ( .A(S), .B(n294), .Z(n293) );
  XOR U441 ( .A(B[199]), .B(B[198]), .Z(n294) );
  XOR U442 ( .A(B[197]), .B(n295), .Z(O[198]) );
  AND U443 ( .A(S), .B(n296), .Z(n295) );
  XOR U444 ( .A(B[198]), .B(B[197]), .Z(n296) );
  XOR U445 ( .A(B[196]), .B(n297), .Z(O[197]) );
  AND U446 ( .A(S), .B(n298), .Z(n297) );
  XOR U447 ( .A(B[197]), .B(B[196]), .Z(n298) );
  XOR U448 ( .A(B[195]), .B(n299), .Z(O[196]) );
  AND U449 ( .A(S), .B(n300), .Z(n299) );
  XOR U450 ( .A(B[196]), .B(B[195]), .Z(n300) );
  XOR U451 ( .A(B[194]), .B(n301), .Z(O[195]) );
  AND U452 ( .A(S), .B(n302), .Z(n301) );
  XOR U453 ( .A(B[195]), .B(B[194]), .Z(n302) );
  XOR U454 ( .A(B[193]), .B(n303), .Z(O[194]) );
  AND U455 ( .A(S), .B(n304), .Z(n303) );
  XOR U456 ( .A(B[194]), .B(B[193]), .Z(n304) );
  XOR U457 ( .A(B[192]), .B(n305), .Z(O[193]) );
  AND U458 ( .A(S), .B(n306), .Z(n305) );
  XOR U459 ( .A(B[193]), .B(B[192]), .Z(n306) );
  XOR U460 ( .A(B[191]), .B(n307), .Z(O[192]) );
  AND U461 ( .A(S), .B(n308), .Z(n307) );
  XOR U462 ( .A(B[192]), .B(B[191]), .Z(n308) );
  XOR U463 ( .A(B[190]), .B(n309), .Z(O[191]) );
  AND U464 ( .A(S), .B(n310), .Z(n309) );
  XOR U465 ( .A(B[191]), .B(B[190]), .Z(n310) );
  XOR U466 ( .A(B[189]), .B(n311), .Z(O[190]) );
  AND U467 ( .A(S), .B(n312), .Z(n311) );
  XOR U468 ( .A(B[190]), .B(B[189]), .Z(n312) );
  XOR U469 ( .A(B[17]), .B(n313), .Z(O[18]) );
  AND U470 ( .A(S), .B(n314), .Z(n313) );
  XOR U471 ( .A(B[18]), .B(B[17]), .Z(n314) );
  XOR U472 ( .A(B[188]), .B(n315), .Z(O[189]) );
  AND U473 ( .A(S), .B(n316), .Z(n315) );
  XOR U474 ( .A(B[189]), .B(B[188]), .Z(n316) );
  XOR U475 ( .A(B[187]), .B(n317), .Z(O[188]) );
  AND U476 ( .A(S), .B(n318), .Z(n317) );
  XOR U477 ( .A(B[188]), .B(B[187]), .Z(n318) );
  XOR U478 ( .A(B[186]), .B(n319), .Z(O[187]) );
  AND U479 ( .A(S), .B(n320), .Z(n319) );
  XOR U480 ( .A(B[187]), .B(B[186]), .Z(n320) );
  XOR U481 ( .A(B[185]), .B(n321), .Z(O[186]) );
  AND U482 ( .A(S), .B(n322), .Z(n321) );
  XOR U483 ( .A(B[186]), .B(B[185]), .Z(n322) );
  XOR U484 ( .A(B[184]), .B(n323), .Z(O[185]) );
  AND U485 ( .A(S), .B(n324), .Z(n323) );
  XOR U486 ( .A(B[185]), .B(B[184]), .Z(n324) );
  XOR U487 ( .A(B[183]), .B(n325), .Z(O[184]) );
  AND U488 ( .A(S), .B(n326), .Z(n325) );
  XOR U489 ( .A(B[184]), .B(B[183]), .Z(n326) );
  XOR U490 ( .A(B[182]), .B(n327), .Z(O[183]) );
  AND U491 ( .A(S), .B(n328), .Z(n327) );
  XOR U492 ( .A(B[183]), .B(B[182]), .Z(n328) );
  XOR U493 ( .A(B[181]), .B(n329), .Z(O[182]) );
  AND U494 ( .A(S), .B(n330), .Z(n329) );
  XOR U495 ( .A(B[182]), .B(B[181]), .Z(n330) );
  XOR U496 ( .A(B[180]), .B(n331), .Z(O[181]) );
  AND U497 ( .A(S), .B(n332), .Z(n331) );
  XOR U498 ( .A(B[181]), .B(B[180]), .Z(n332) );
  XOR U499 ( .A(B[179]), .B(n333), .Z(O[180]) );
  AND U500 ( .A(S), .B(n334), .Z(n333) );
  XOR U501 ( .A(B[180]), .B(B[179]), .Z(n334) );
  XOR U502 ( .A(B[16]), .B(n335), .Z(O[17]) );
  AND U503 ( .A(S), .B(n336), .Z(n335) );
  XOR U504 ( .A(B[17]), .B(B[16]), .Z(n336) );
  XOR U505 ( .A(B[178]), .B(n337), .Z(O[179]) );
  AND U506 ( .A(S), .B(n338), .Z(n337) );
  XOR U507 ( .A(B[179]), .B(B[178]), .Z(n338) );
  XOR U508 ( .A(B[177]), .B(n339), .Z(O[178]) );
  AND U509 ( .A(S), .B(n340), .Z(n339) );
  XOR U510 ( .A(B[178]), .B(B[177]), .Z(n340) );
  XOR U511 ( .A(B[176]), .B(n341), .Z(O[177]) );
  AND U512 ( .A(S), .B(n342), .Z(n341) );
  XOR U513 ( .A(B[177]), .B(B[176]), .Z(n342) );
  XOR U514 ( .A(B[175]), .B(n343), .Z(O[176]) );
  AND U515 ( .A(S), .B(n344), .Z(n343) );
  XOR U516 ( .A(B[176]), .B(B[175]), .Z(n344) );
  XOR U517 ( .A(B[174]), .B(n345), .Z(O[175]) );
  AND U518 ( .A(S), .B(n346), .Z(n345) );
  XOR U519 ( .A(B[175]), .B(B[174]), .Z(n346) );
  XOR U520 ( .A(B[173]), .B(n347), .Z(O[174]) );
  AND U521 ( .A(S), .B(n348), .Z(n347) );
  XOR U522 ( .A(B[174]), .B(B[173]), .Z(n348) );
  XOR U523 ( .A(B[172]), .B(n349), .Z(O[173]) );
  AND U524 ( .A(S), .B(n350), .Z(n349) );
  XOR U525 ( .A(B[173]), .B(B[172]), .Z(n350) );
  XOR U526 ( .A(B[171]), .B(n351), .Z(O[172]) );
  AND U527 ( .A(S), .B(n352), .Z(n351) );
  XOR U528 ( .A(B[172]), .B(B[171]), .Z(n352) );
  XOR U529 ( .A(B[170]), .B(n353), .Z(O[171]) );
  AND U530 ( .A(S), .B(n354), .Z(n353) );
  XOR U531 ( .A(B[171]), .B(B[170]), .Z(n354) );
  XOR U532 ( .A(B[169]), .B(n355), .Z(O[170]) );
  AND U533 ( .A(S), .B(n356), .Z(n355) );
  XOR U534 ( .A(B[170]), .B(B[169]), .Z(n356) );
  XOR U535 ( .A(B[15]), .B(n357), .Z(O[16]) );
  AND U536 ( .A(S), .B(n358), .Z(n357) );
  XOR U537 ( .A(B[16]), .B(B[15]), .Z(n358) );
  XOR U538 ( .A(B[168]), .B(n359), .Z(O[169]) );
  AND U539 ( .A(S), .B(n360), .Z(n359) );
  XOR U540 ( .A(B[169]), .B(B[168]), .Z(n360) );
  XOR U541 ( .A(B[167]), .B(n361), .Z(O[168]) );
  AND U542 ( .A(S), .B(n362), .Z(n361) );
  XOR U543 ( .A(B[168]), .B(B[167]), .Z(n362) );
  XOR U544 ( .A(B[166]), .B(n363), .Z(O[167]) );
  AND U545 ( .A(S), .B(n364), .Z(n363) );
  XOR U546 ( .A(B[167]), .B(B[166]), .Z(n364) );
  XOR U547 ( .A(B[165]), .B(n365), .Z(O[166]) );
  AND U548 ( .A(S), .B(n366), .Z(n365) );
  XOR U549 ( .A(B[166]), .B(B[165]), .Z(n366) );
  XOR U550 ( .A(B[164]), .B(n367), .Z(O[165]) );
  AND U551 ( .A(S), .B(n368), .Z(n367) );
  XOR U552 ( .A(B[165]), .B(B[164]), .Z(n368) );
  XOR U553 ( .A(B[163]), .B(n369), .Z(O[164]) );
  AND U554 ( .A(S), .B(n370), .Z(n369) );
  XOR U555 ( .A(B[164]), .B(B[163]), .Z(n370) );
  XOR U556 ( .A(B[162]), .B(n371), .Z(O[163]) );
  AND U557 ( .A(S), .B(n372), .Z(n371) );
  XOR U558 ( .A(B[163]), .B(B[162]), .Z(n372) );
  XOR U559 ( .A(B[161]), .B(n373), .Z(O[162]) );
  AND U560 ( .A(S), .B(n374), .Z(n373) );
  XOR U561 ( .A(B[162]), .B(B[161]), .Z(n374) );
  XOR U562 ( .A(B[160]), .B(n375), .Z(O[161]) );
  AND U563 ( .A(S), .B(n376), .Z(n375) );
  XOR U564 ( .A(B[161]), .B(B[160]), .Z(n376) );
  XOR U565 ( .A(B[159]), .B(n377), .Z(O[160]) );
  AND U566 ( .A(S), .B(n378), .Z(n377) );
  XOR U567 ( .A(B[160]), .B(B[159]), .Z(n378) );
  XOR U568 ( .A(B[14]), .B(n379), .Z(O[15]) );
  AND U569 ( .A(S), .B(n380), .Z(n379) );
  XOR U570 ( .A(B[15]), .B(B[14]), .Z(n380) );
  XOR U571 ( .A(B[158]), .B(n381), .Z(O[159]) );
  AND U572 ( .A(S), .B(n382), .Z(n381) );
  XOR U573 ( .A(B[159]), .B(B[158]), .Z(n382) );
  XOR U574 ( .A(B[157]), .B(n383), .Z(O[158]) );
  AND U575 ( .A(S), .B(n384), .Z(n383) );
  XOR U576 ( .A(B[158]), .B(B[157]), .Z(n384) );
  XOR U577 ( .A(B[156]), .B(n385), .Z(O[157]) );
  AND U578 ( .A(S), .B(n386), .Z(n385) );
  XOR U579 ( .A(B[157]), .B(B[156]), .Z(n386) );
  XOR U580 ( .A(B[155]), .B(n387), .Z(O[156]) );
  AND U581 ( .A(S), .B(n388), .Z(n387) );
  XOR U582 ( .A(B[156]), .B(B[155]), .Z(n388) );
  XOR U583 ( .A(B[154]), .B(n389), .Z(O[155]) );
  AND U584 ( .A(S), .B(n390), .Z(n389) );
  XOR U585 ( .A(B[155]), .B(B[154]), .Z(n390) );
  XOR U586 ( .A(B[153]), .B(n391), .Z(O[154]) );
  AND U587 ( .A(S), .B(n392), .Z(n391) );
  XOR U588 ( .A(B[154]), .B(B[153]), .Z(n392) );
  XOR U589 ( .A(B[152]), .B(n393), .Z(O[153]) );
  AND U590 ( .A(S), .B(n394), .Z(n393) );
  XOR U591 ( .A(B[153]), .B(B[152]), .Z(n394) );
  XOR U592 ( .A(B[151]), .B(n395), .Z(O[152]) );
  AND U593 ( .A(S), .B(n396), .Z(n395) );
  XOR U594 ( .A(B[152]), .B(B[151]), .Z(n396) );
  XOR U595 ( .A(B[150]), .B(n397), .Z(O[151]) );
  AND U596 ( .A(S), .B(n398), .Z(n397) );
  XOR U597 ( .A(B[151]), .B(B[150]), .Z(n398) );
  XOR U598 ( .A(B[149]), .B(n399), .Z(O[150]) );
  AND U599 ( .A(S), .B(n400), .Z(n399) );
  XOR U600 ( .A(B[150]), .B(B[149]), .Z(n400) );
  XOR U601 ( .A(B[13]), .B(n401), .Z(O[14]) );
  AND U602 ( .A(S), .B(n402), .Z(n401) );
  XOR U603 ( .A(B[14]), .B(B[13]), .Z(n402) );
  XOR U604 ( .A(B[148]), .B(n403), .Z(O[149]) );
  AND U605 ( .A(S), .B(n404), .Z(n403) );
  XOR U606 ( .A(B[149]), .B(B[148]), .Z(n404) );
  XOR U607 ( .A(B[147]), .B(n405), .Z(O[148]) );
  AND U608 ( .A(S), .B(n406), .Z(n405) );
  XOR U609 ( .A(B[148]), .B(B[147]), .Z(n406) );
  XOR U610 ( .A(B[146]), .B(n407), .Z(O[147]) );
  AND U611 ( .A(S), .B(n408), .Z(n407) );
  XOR U612 ( .A(B[147]), .B(B[146]), .Z(n408) );
  XOR U613 ( .A(B[145]), .B(n409), .Z(O[146]) );
  AND U614 ( .A(S), .B(n410), .Z(n409) );
  XOR U615 ( .A(B[146]), .B(B[145]), .Z(n410) );
  XOR U616 ( .A(B[144]), .B(n411), .Z(O[145]) );
  AND U617 ( .A(S), .B(n412), .Z(n411) );
  XOR U618 ( .A(B[145]), .B(B[144]), .Z(n412) );
  XOR U619 ( .A(B[143]), .B(n413), .Z(O[144]) );
  AND U620 ( .A(S), .B(n414), .Z(n413) );
  XOR U621 ( .A(B[144]), .B(B[143]), .Z(n414) );
  XOR U622 ( .A(B[142]), .B(n415), .Z(O[143]) );
  AND U623 ( .A(S), .B(n416), .Z(n415) );
  XOR U624 ( .A(B[143]), .B(B[142]), .Z(n416) );
  XOR U625 ( .A(B[141]), .B(n417), .Z(O[142]) );
  AND U626 ( .A(S), .B(n418), .Z(n417) );
  XOR U627 ( .A(B[142]), .B(B[141]), .Z(n418) );
  XOR U628 ( .A(B[140]), .B(n419), .Z(O[141]) );
  AND U629 ( .A(S), .B(n420), .Z(n419) );
  XOR U630 ( .A(B[141]), .B(B[140]), .Z(n420) );
  XOR U631 ( .A(B[139]), .B(n421), .Z(O[140]) );
  AND U632 ( .A(S), .B(n422), .Z(n421) );
  XOR U633 ( .A(B[140]), .B(B[139]), .Z(n422) );
  XOR U634 ( .A(B[12]), .B(n423), .Z(O[13]) );
  AND U635 ( .A(S), .B(n424), .Z(n423) );
  XOR U636 ( .A(B[13]), .B(B[12]), .Z(n424) );
  XOR U637 ( .A(B[138]), .B(n425), .Z(O[139]) );
  AND U638 ( .A(S), .B(n426), .Z(n425) );
  XOR U639 ( .A(B[139]), .B(B[138]), .Z(n426) );
  XOR U640 ( .A(B[137]), .B(n427), .Z(O[138]) );
  AND U641 ( .A(S), .B(n428), .Z(n427) );
  XOR U642 ( .A(B[138]), .B(B[137]), .Z(n428) );
  XOR U643 ( .A(B[136]), .B(n429), .Z(O[137]) );
  AND U644 ( .A(S), .B(n430), .Z(n429) );
  XOR U645 ( .A(B[137]), .B(B[136]), .Z(n430) );
  XOR U646 ( .A(B[135]), .B(n431), .Z(O[136]) );
  AND U647 ( .A(S), .B(n432), .Z(n431) );
  XOR U648 ( .A(B[136]), .B(B[135]), .Z(n432) );
  XOR U649 ( .A(B[134]), .B(n433), .Z(O[135]) );
  AND U650 ( .A(S), .B(n434), .Z(n433) );
  XOR U651 ( .A(B[135]), .B(B[134]), .Z(n434) );
  XOR U652 ( .A(B[133]), .B(n435), .Z(O[134]) );
  AND U653 ( .A(S), .B(n436), .Z(n435) );
  XOR U654 ( .A(B[134]), .B(B[133]), .Z(n436) );
  XOR U655 ( .A(B[132]), .B(n437), .Z(O[133]) );
  AND U656 ( .A(S), .B(n438), .Z(n437) );
  XOR U657 ( .A(B[133]), .B(B[132]), .Z(n438) );
  XOR U658 ( .A(B[131]), .B(n439), .Z(O[132]) );
  AND U659 ( .A(S), .B(n440), .Z(n439) );
  XOR U660 ( .A(B[132]), .B(B[131]), .Z(n440) );
  XOR U661 ( .A(B[130]), .B(n441), .Z(O[131]) );
  AND U662 ( .A(S), .B(n442), .Z(n441) );
  XOR U663 ( .A(B[131]), .B(B[130]), .Z(n442) );
  XOR U664 ( .A(B[129]), .B(n443), .Z(O[130]) );
  AND U665 ( .A(S), .B(n444), .Z(n443) );
  XOR U666 ( .A(B[130]), .B(B[129]), .Z(n444) );
  XOR U667 ( .A(B[11]), .B(n445), .Z(O[12]) );
  AND U668 ( .A(S), .B(n446), .Z(n445) );
  XOR U669 ( .A(B[12]), .B(B[11]), .Z(n446) );
  XOR U670 ( .A(B[128]), .B(n447), .Z(O[129]) );
  AND U671 ( .A(S), .B(n448), .Z(n447) );
  XOR U672 ( .A(B[129]), .B(B[128]), .Z(n448) );
  XOR U673 ( .A(B[127]), .B(n449), .Z(O[128]) );
  AND U674 ( .A(S), .B(n450), .Z(n449) );
  XOR U675 ( .A(B[128]), .B(B[127]), .Z(n450) );
  XOR U676 ( .A(B[126]), .B(n451), .Z(O[127]) );
  AND U677 ( .A(S), .B(n452), .Z(n451) );
  XOR U678 ( .A(B[127]), .B(B[126]), .Z(n452) );
  XOR U679 ( .A(B[125]), .B(n453), .Z(O[126]) );
  AND U680 ( .A(S), .B(n454), .Z(n453) );
  XOR U681 ( .A(B[126]), .B(B[125]), .Z(n454) );
  XOR U682 ( .A(B[124]), .B(n455), .Z(O[125]) );
  AND U683 ( .A(S), .B(n456), .Z(n455) );
  XOR U684 ( .A(B[125]), .B(B[124]), .Z(n456) );
  XOR U685 ( .A(B[123]), .B(n457), .Z(O[124]) );
  AND U686 ( .A(S), .B(n458), .Z(n457) );
  XOR U687 ( .A(B[124]), .B(B[123]), .Z(n458) );
  XOR U688 ( .A(B[122]), .B(n459), .Z(O[123]) );
  AND U689 ( .A(S), .B(n460), .Z(n459) );
  XOR U690 ( .A(B[123]), .B(B[122]), .Z(n460) );
  XOR U691 ( .A(B[121]), .B(n461), .Z(O[122]) );
  AND U692 ( .A(S), .B(n462), .Z(n461) );
  XOR U693 ( .A(B[122]), .B(B[121]), .Z(n462) );
  XOR U694 ( .A(B[120]), .B(n463), .Z(O[121]) );
  AND U695 ( .A(S), .B(n464), .Z(n463) );
  XOR U696 ( .A(B[121]), .B(B[120]), .Z(n464) );
  XOR U697 ( .A(B[119]), .B(n465), .Z(O[120]) );
  AND U698 ( .A(S), .B(n466), .Z(n465) );
  XOR U699 ( .A(B[120]), .B(B[119]), .Z(n466) );
  XOR U700 ( .A(B[10]), .B(n467), .Z(O[11]) );
  AND U701 ( .A(S), .B(n468), .Z(n467) );
  XOR U702 ( .A(B[11]), .B(B[10]), .Z(n468) );
  XOR U703 ( .A(B[118]), .B(n469), .Z(O[119]) );
  AND U704 ( .A(S), .B(n470), .Z(n469) );
  XOR U705 ( .A(B[119]), .B(B[118]), .Z(n470) );
  XOR U706 ( .A(B[117]), .B(n471), .Z(O[118]) );
  AND U707 ( .A(S), .B(n472), .Z(n471) );
  XOR U708 ( .A(B[118]), .B(B[117]), .Z(n472) );
  XOR U709 ( .A(B[116]), .B(n473), .Z(O[117]) );
  AND U710 ( .A(S), .B(n474), .Z(n473) );
  XOR U711 ( .A(B[117]), .B(B[116]), .Z(n474) );
  XOR U712 ( .A(B[115]), .B(n475), .Z(O[116]) );
  AND U713 ( .A(S), .B(n476), .Z(n475) );
  XOR U714 ( .A(B[116]), .B(B[115]), .Z(n476) );
  XOR U715 ( .A(B[114]), .B(n477), .Z(O[115]) );
  AND U716 ( .A(S), .B(n478), .Z(n477) );
  XOR U717 ( .A(B[115]), .B(B[114]), .Z(n478) );
  XOR U718 ( .A(B[113]), .B(n479), .Z(O[114]) );
  AND U719 ( .A(S), .B(n480), .Z(n479) );
  XOR U720 ( .A(B[114]), .B(B[113]), .Z(n480) );
  XOR U721 ( .A(B[112]), .B(n481), .Z(O[113]) );
  AND U722 ( .A(S), .B(n482), .Z(n481) );
  XOR U723 ( .A(B[113]), .B(B[112]), .Z(n482) );
  XOR U724 ( .A(B[111]), .B(n483), .Z(O[112]) );
  AND U725 ( .A(S), .B(n484), .Z(n483) );
  XOR U726 ( .A(B[112]), .B(B[111]), .Z(n484) );
  XOR U727 ( .A(B[110]), .B(n485), .Z(O[111]) );
  AND U728 ( .A(S), .B(n486), .Z(n485) );
  XOR U729 ( .A(B[111]), .B(B[110]), .Z(n486) );
  XOR U730 ( .A(B[109]), .B(n487), .Z(O[110]) );
  AND U731 ( .A(S), .B(n488), .Z(n487) );
  XOR U732 ( .A(B[110]), .B(B[109]), .Z(n488) );
  XOR U733 ( .A(B[9]), .B(n489), .Z(O[10]) );
  AND U734 ( .A(S), .B(n490), .Z(n489) );
  XOR U735 ( .A(B[9]), .B(B[10]), .Z(n490) );
  XOR U736 ( .A(B[108]), .B(n491), .Z(O[109]) );
  AND U737 ( .A(S), .B(n492), .Z(n491) );
  XOR U738 ( .A(B[109]), .B(B[108]), .Z(n492) );
  XOR U739 ( .A(B[107]), .B(n493), .Z(O[108]) );
  AND U740 ( .A(S), .B(n494), .Z(n493) );
  XOR U741 ( .A(B[108]), .B(B[107]), .Z(n494) );
  XOR U742 ( .A(B[106]), .B(n495), .Z(O[107]) );
  AND U743 ( .A(S), .B(n496), .Z(n495) );
  XOR U744 ( .A(B[107]), .B(B[106]), .Z(n496) );
  XOR U745 ( .A(B[105]), .B(n497), .Z(O[106]) );
  AND U746 ( .A(S), .B(n498), .Z(n497) );
  XOR U747 ( .A(B[106]), .B(B[105]), .Z(n498) );
  XOR U748 ( .A(B[104]), .B(n499), .Z(O[105]) );
  AND U749 ( .A(S), .B(n500), .Z(n499) );
  XOR U750 ( .A(B[105]), .B(B[104]), .Z(n500) );
  XOR U751 ( .A(B[103]), .B(n501), .Z(O[104]) );
  AND U752 ( .A(S), .B(n502), .Z(n501) );
  XOR U753 ( .A(B[104]), .B(B[103]), .Z(n502) );
  XOR U754 ( .A(B[102]), .B(n503), .Z(O[103]) );
  AND U755 ( .A(S), .B(n504), .Z(n503) );
  XOR U756 ( .A(B[103]), .B(B[102]), .Z(n504) );
  XOR U757 ( .A(B[101]), .B(n505), .Z(O[102]) );
  AND U758 ( .A(S), .B(n506), .Z(n505) );
  XOR U759 ( .A(B[102]), .B(B[101]), .Z(n506) );
  XOR U760 ( .A(B[100]), .B(n507), .Z(O[101]) );
  AND U761 ( .A(S), .B(n508), .Z(n507) );
  XOR U762 ( .A(B[101]), .B(B[100]), .Z(n508) );
  XOR U763 ( .A(B[99]), .B(n509), .Z(O[100]) );
  AND U764 ( .A(S), .B(n510), .Z(n509) );
  XOR U765 ( .A(B[99]), .B(B[100]), .Z(n510) );
  AND U766 ( .A(B[0]), .B(S), .Z(O[0]) );
endmodule


module modexp_2N_NN_N256_CC65536 ( clk, rst, m, e, n, c );
  input [255:0] m;
  input [255:0] e;
  input [255:0] n;
  output [255:0] c;
  input clk, rst;
  wire   _0_net_, first_one, mul_pow, n6, n8, n137, n138, n139, n140;
  wire   [127:0] start_in;
  wire   [255:0] ein;
  wire   [255:0] creg_next;
  wire   [255:0] o;
  wire   [255:0] ereg_next;
  wire   [255:0] y;

  MUX_N256_3 MUX_4 ( .A(o), .B(c), .S(_0_net_), .O(creg_next) );
  MUX_N256_5 MUX_6 ( .A({ein[254:0], 1'b0}), .B(ein), .S(mul_pow), .O(
        ereg_next) );
  MUX_N256_4 MUX_9 ( .A(m), .B(c), .S(mul_pow), .O(y) );
  modmult_N256_CC128 modmult_1 ( .clk(clk), .rst(1'b0), .start(start_in[0]), 
        .x(c), .y(y), .n(n), .o(o) );
  DFF \start_reg_reg[0]  ( .D(start_in[127]), .CLK(clk), .RST(rst), .I(1'b1), 
        .Q(start_in[0]) );
  DFF \start_reg_reg[1]  ( .D(start_in[0]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[1]) );
  DFF \start_reg_reg[2]  ( .D(start_in[1]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[2]) );
  DFF \start_reg_reg[3]  ( .D(start_in[2]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[3]) );
  DFF \start_reg_reg[4]  ( .D(start_in[3]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[4]) );
  DFF \start_reg_reg[5]  ( .D(start_in[4]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[5]) );
  DFF \start_reg_reg[6]  ( .D(start_in[5]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[6]) );
  DFF \start_reg_reg[7]  ( .D(start_in[6]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[7]) );
  DFF \start_reg_reg[8]  ( .D(start_in[7]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[8]) );
  DFF \start_reg_reg[9]  ( .D(start_in[8]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[9]) );
  DFF \start_reg_reg[10]  ( .D(start_in[9]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[10]) );
  DFF \start_reg_reg[11]  ( .D(start_in[10]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[11]) );
  DFF \start_reg_reg[12]  ( .D(start_in[11]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[12]) );
  DFF \start_reg_reg[13]  ( .D(start_in[12]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[13]) );
  DFF \start_reg_reg[14]  ( .D(start_in[13]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[14]) );
  DFF \start_reg_reg[15]  ( .D(start_in[14]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[15]) );
  DFF \start_reg_reg[16]  ( .D(start_in[15]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[16]) );
  DFF \start_reg_reg[17]  ( .D(start_in[16]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[17]) );
  DFF \start_reg_reg[18]  ( .D(start_in[17]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[18]) );
  DFF \start_reg_reg[19]  ( .D(start_in[18]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[19]) );
  DFF \start_reg_reg[20]  ( .D(start_in[19]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[20]) );
  DFF \start_reg_reg[21]  ( .D(start_in[20]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[21]) );
  DFF \start_reg_reg[22]  ( .D(start_in[21]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[22]) );
  DFF \start_reg_reg[23]  ( .D(start_in[22]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[23]) );
  DFF \start_reg_reg[24]  ( .D(start_in[23]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[24]) );
  DFF \start_reg_reg[25]  ( .D(start_in[24]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[25]) );
  DFF \start_reg_reg[26]  ( .D(start_in[25]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[26]) );
  DFF \start_reg_reg[27]  ( .D(start_in[26]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[27]) );
  DFF \start_reg_reg[28]  ( .D(start_in[27]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[28]) );
  DFF \start_reg_reg[29]  ( .D(start_in[28]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[29]) );
  DFF \start_reg_reg[30]  ( .D(start_in[29]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[30]) );
  DFF \start_reg_reg[31]  ( .D(start_in[30]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[31]) );
  DFF \start_reg_reg[32]  ( .D(start_in[31]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[32]) );
  DFF \start_reg_reg[33]  ( .D(start_in[32]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[33]) );
  DFF \start_reg_reg[34]  ( .D(start_in[33]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[34]) );
  DFF \start_reg_reg[35]  ( .D(start_in[34]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[35]) );
  DFF \start_reg_reg[36]  ( .D(start_in[35]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[36]) );
  DFF \start_reg_reg[37]  ( .D(start_in[36]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[37]) );
  DFF \start_reg_reg[38]  ( .D(start_in[37]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[38]) );
  DFF \start_reg_reg[39]  ( .D(start_in[38]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[39]) );
  DFF \start_reg_reg[40]  ( .D(start_in[39]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[40]) );
  DFF \start_reg_reg[41]  ( .D(start_in[40]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[41]) );
  DFF \start_reg_reg[42]  ( .D(start_in[41]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[42]) );
  DFF \start_reg_reg[43]  ( .D(start_in[42]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[43]) );
  DFF \start_reg_reg[44]  ( .D(start_in[43]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[44]) );
  DFF \start_reg_reg[45]  ( .D(start_in[44]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[45]) );
  DFF \start_reg_reg[46]  ( .D(start_in[45]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[46]) );
  DFF \start_reg_reg[47]  ( .D(start_in[46]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[47]) );
  DFF \start_reg_reg[48]  ( .D(start_in[47]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[48]) );
  DFF \start_reg_reg[49]  ( .D(start_in[48]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[49]) );
  DFF \start_reg_reg[50]  ( .D(start_in[49]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[50]) );
  DFF \start_reg_reg[51]  ( .D(start_in[50]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[51]) );
  DFF \start_reg_reg[52]  ( .D(start_in[51]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[52]) );
  DFF \start_reg_reg[53]  ( .D(start_in[52]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[53]) );
  DFF \start_reg_reg[54]  ( .D(start_in[53]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[54]) );
  DFF \start_reg_reg[55]  ( .D(start_in[54]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[55]) );
  DFF \start_reg_reg[56]  ( .D(start_in[55]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[56]) );
  DFF \start_reg_reg[57]  ( .D(start_in[56]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[57]) );
  DFF \start_reg_reg[58]  ( .D(start_in[57]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[58]) );
  DFF \start_reg_reg[59]  ( .D(start_in[58]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[59]) );
  DFF \start_reg_reg[60]  ( .D(start_in[59]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[60]) );
  DFF \start_reg_reg[61]  ( .D(start_in[60]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[61]) );
  DFF \start_reg_reg[62]  ( .D(start_in[61]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[62]) );
  DFF \start_reg_reg[63]  ( .D(start_in[62]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[63]) );
  DFF \start_reg_reg[64]  ( .D(start_in[63]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[64]) );
  DFF \start_reg_reg[65]  ( .D(start_in[64]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[65]) );
  DFF \start_reg_reg[66]  ( .D(start_in[65]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[66]) );
  DFF \start_reg_reg[67]  ( .D(start_in[66]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[67]) );
  DFF \start_reg_reg[68]  ( .D(start_in[67]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[68]) );
  DFF \start_reg_reg[69]  ( .D(start_in[68]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[69]) );
  DFF \start_reg_reg[70]  ( .D(start_in[69]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[70]) );
  DFF \start_reg_reg[71]  ( .D(start_in[70]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[71]) );
  DFF \start_reg_reg[72]  ( .D(start_in[71]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[72]) );
  DFF \start_reg_reg[73]  ( .D(start_in[72]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[73]) );
  DFF \start_reg_reg[74]  ( .D(start_in[73]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[74]) );
  DFF \start_reg_reg[75]  ( .D(start_in[74]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[75]) );
  DFF \start_reg_reg[76]  ( .D(start_in[75]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[76]) );
  DFF \start_reg_reg[77]  ( .D(start_in[76]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[77]) );
  DFF \start_reg_reg[78]  ( .D(start_in[77]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[78]) );
  DFF \start_reg_reg[79]  ( .D(start_in[78]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[79]) );
  DFF \start_reg_reg[80]  ( .D(start_in[79]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[80]) );
  DFF \start_reg_reg[81]  ( .D(start_in[80]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[81]) );
  DFF \start_reg_reg[82]  ( .D(start_in[81]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[82]) );
  DFF \start_reg_reg[83]  ( .D(start_in[82]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[83]) );
  DFF \start_reg_reg[84]  ( .D(start_in[83]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[84]) );
  DFF \start_reg_reg[85]  ( .D(start_in[84]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[85]) );
  DFF \start_reg_reg[86]  ( .D(start_in[85]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[86]) );
  DFF \start_reg_reg[87]  ( .D(start_in[86]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[87]) );
  DFF \start_reg_reg[88]  ( .D(start_in[87]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[88]) );
  DFF \start_reg_reg[89]  ( .D(start_in[88]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[89]) );
  DFF \start_reg_reg[90]  ( .D(start_in[89]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[90]) );
  DFF \start_reg_reg[91]  ( .D(start_in[90]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[91]) );
  DFF \start_reg_reg[92]  ( .D(start_in[91]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[92]) );
  DFF \start_reg_reg[93]  ( .D(start_in[92]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[93]) );
  DFF \start_reg_reg[94]  ( .D(start_in[93]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[94]) );
  DFF \start_reg_reg[95]  ( .D(start_in[94]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[95]) );
  DFF \start_reg_reg[96]  ( .D(start_in[95]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[96]) );
  DFF \start_reg_reg[97]  ( .D(start_in[96]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[97]) );
  DFF \start_reg_reg[98]  ( .D(start_in[97]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[98]) );
  DFF \start_reg_reg[99]  ( .D(start_in[98]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[99]) );
  DFF \start_reg_reg[100]  ( .D(start_in[99]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[100]) );
  DFF \start_reg_reg[101]  ( .D(start_in[100]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[101]) );
  DFF \start_reg_reg[102]  ( .D(start_in[101]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[102]) );
  DFF \start_reg_reg[103]  ( .D(start_in[102]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[103]) );
  DFF \start_reg_reg[104]  ( .D(start_in[103]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[104]) );
  DFF \start_reg_reg[105]  ( .D(start_in[104]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[105]) );
  DFF \start_reg_reg[106]  ( .D(start_in[105]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[106]) );
  DFF \start_reg_reg[107]  ( .D(start_in[106]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[107]) );
  DFF \start_reg_reg[108]  ( .D(start_in[107]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[108]) );
  DFF \start_reg_reg[109]  ( .D(start_in[108]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[109]) );
  DFF \start_reg_reg[110]  ( .D(start_in[109]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[110]) );
  DFF \start_reg_reg[111]  ( .D(start_in[110]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[111]) );
  DFF \start_reg_reg[112]  ( .D(start_in[111]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[112]) );
  DFF \start_reg_reg[113]  ( .D(start_in[112]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[113]) );
  DFF \start_reg_reg[114]  ( .D(start_in[113]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[114]) );
  DFF \start_reg_reg[115]  ( .D(start_in[114]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[115]) );
  DFF \start_reg_reg[116]  ( .D(start_in[115]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[116]) );
  DFF \start_reg_reg[117]  ( .D(start_in[116]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[117]) );
  DFF \start_reg_reg[118]  ( .D(start_in[117]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[118]) );
  DFF \start_reg_reg[119]  ( .D(start_in[118]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[119]) );
  DFF \start_reg_reg[120]  ( .D(start_in[119]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[120]) );
  DFF \start_reg_reg[121]  ( .D(start_in[120]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[121]) );
  DFF \start_reg_reg[122]  ( .D(start_in[121]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[122]) );
  DFF \start_reg_reg[123]  ( .D(start_in[122]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[123]) );
  DFF \start_reg_reg[124]  ( .D(start_in[123]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[124]) );
  DFF \start_reg_reg[125]  ( .D(start_in[124]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[125]) );
  DFF \start_reg_reg[126]  ( .D(start_in[125]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[126]) );
  DFF \start_reg_reg[127]  ( .D(start_in[126]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[127]) );
  DFF mul_pow_reg ( .D(n8), .CLK(clk), .RST(rst), .I(1'b0), .Q(mul_pow) );
  DFF \ereg_reg[0]  ( .D(ereg_next[0]), .CLK(clk), .RST(rst), .I(e[0]), .Q(
        ein[0]) );
  DFF \ereg_reg[1]  ( .D(ereg_next[1]), .CLK(clk), .RST(rst), .I(e[1]), .Q(
        ein[1]) );
  DFF \ereg_reg[2]  ( .D(ereg_next[2]), .CLK(clk), .RST(rst), .I(e[2]), .Q(
        ein[2]) );
  DFF \ereg_reg[3]  ( .D(ereg_next[3]), .CLK(clk), .RST(rst), .I(e[3]), .Q(
        ein[3]) );
  DFF \ereg_reg[4]  ( .D(ereg_next[4]), .CLK(clk), .RST(rst), .I(e[4]), .Q(
        ein[4]) );
  DFF \ereg_reg[5]  ( .D(ereg_next[5]), .CLK(clk), .RST(rst), .I(e[5]), .Q(
        ein[5]) );
  DFF \ereg_reg[6]  ( .D(ereg_next[6]), .CLK(clk), .RST(rst), .I(e[6]), .Q(
        ein[6]) );
  DFF \ereg_reg[7]  ( .D(ereg_next[7]), .CLK(clk), .RST(rst), .I(e[7]), .Q(
        ein[7]) );
  DFF \ereg_reg[8]  ( .D(ereg_next[8]), .CLK(clk), .RST(rst), .I(e[8]), .Q(
        ein[8]) );
  DFF \ereg_reg[9]  ( .D(ereg_next[9]), .CLK(clk), .RST(rst), .I(e[9]), .Q(
        ein[9]) );
  DFF \ereg_reg[10]  ( .D(ereg_next[10]), .CLK(clk), .RST(rst), .I(e[10]), .Q(
        ein[10]) );
  DFF \ereg_reg[11]  ( .D(ereg_next[11]), .CLK(clk), .RST(rst), .I(e[11]), .Q(
        ein[11]) );
  DFF \ereg_reg[12]  ( .D(ereg_next[12]), .CLK(clk), .RST(rst), .I(e[12]), .Q(
        ein[12]) );
  DFF \ereg_reg[13]  ( .D(ereg_next[13]), .CLK(clk), .RST(rst), .I(e[13]), .Q(
        ein[13]) );
  DFF \ereg_reg[14]  ( .D(ereg_next[14]), .CLK(clk), .RST(rst), .I(e[14]), .Q(
        ein[14]) );
  DFF \ereg_reg[15]  ( .D(ereg_next[15]), .CLK(clk), .RST(rst), .I(e[15]), .Q(
        ein[15]) );
  DFF \ereg_reg[16]  ( .D(ereg_next[16]), .CLK(clk), .RST(rst), .I(e[16]), .Q(
        ein[16]) );
  DFF \ereg_reg[17]  ( .D(ereg_next[17]), .CLK(clk), .RST(rst), .I(e[17]), .Q(
        ein[17]) );
  DFF \ereg_reg[18]  ( .D(ereg_next[18]), .CLK(clk), .RST(rst), .I(e[18]), .Q(
        ein[18]) );
  DFF \ereg_reg[19]  ( .D(ereg_next[19]), .CLK(clk), .RST(rst), .I(e[19]), .Q(
        ein[19]) );
  DFF \ereg_reg[20]  ( .D(ereg_next[20]), .CLK(clk), .RST(rst), .I(e[20]), .Q(
        ein[20]) );
  DFF \ereg_reg[21]  ( .D(ereg_next[21]), .CLK(clk), .RST(rst), .I(e[21]), .Q(
        ein[21]) );
  DFF \ereg_reg[22]  ( .D(ereg_next[22]), .CLK(clk), .RST(rst), .I(e[22]), .Q(
        ein[22]) );
  DFF \ereg_reg[23]  ( .D(ereg_next[23]), .CLK(clk), .RST(rst), .I(e[23]), .Q(
        ein[23]) );
  DFF \ereg_reg[24]  ( .D(ereg_next[24]), .CLK(clk), .RST(rst), .I(e[24]), .Q(
        ein[24]) );
  DFF \ereg_reg[25]  ( .D(ereg_next[25]), .CLK(clk), .RST(rst), .I(e[25]), .Q(
        ein[25]) );
  DFF \ereg_reg[26]  ( .D(ereg_next[26]), .CLK(clk), .RST(rst), .I(e[26]), .Q(
        ein[26]) );
  DFF \ereg_reg[27]  ( .D(ereg_next[27]), .CLK(clk), .RST(rst), .I(e[27]), .Q(
        ein[27]) );
  DFF \ereg_reg[28]  ( .D(ereg_next[28]), .CLK(clk), .RST(rst), .I(e[28]), .Q(
        ein[28]) );
  DFF \ereg_reg[29]  ( .D(ereg_next[29]), .CLK(clk), .RST(rst), .I(e[29]), .Q(
        ein[29]) );
  DFF \ereg_reg[30]  ( .D(ereg_next[30]), .CLK(clk), .RST(rst), .I(e[30]), .Q(
        ein[30]) );
  DFF \ereg_reg[31]  ( .D(ereg_next[31]), .CLK(clk), .RST(rst), .I(e[31]), .Q(
        ein[31]) );
  DFF \ereg_reg[32]  ( .D(ereg_next[32]), .CLK(clk), .RST(rst), .I(e[32]), .Q(
        ein[32]) );
  DFF \ereg_reg[33]  ( .D(ereg_next[33]), .CLK(clk), .RST(rst), .I(e[33]), .Q(
        ein[33]) );
  DFF \ereg_reg[34]  ( .D(ereg_next[34]), .CLK(clk), .RST(rst), .I(e[34]), .Q(
        ein[34]) );
  DFF \ereg_reg[35]  ( .D(ereg_next[35]), .CLK(clk), .RST(rst), .I(e[35]), .Q(
        ein[35]) );
  DFF \ereg_reg[36]  ( .D(ereg_next[36]), .CLK(clk), .RST(rst), .I(e[36]), .Q(
        ein[36]) );
  DFF \ereg_reg[37]  ( .D(ereg_next[37]), .CLK(clk), .RST(rst), .I(e[37]), .Q(
        ein[37]) );
  DFF \ereg_reg[38]  ( .D(ereg_next[38]), .CLK(clk), .RST(rst), .I(e[38]), .Q(
        ein[38]) );
  DFF \ereg_reg[39]  ( .D(ereg_next[39]), .CLK(clk), .RST(rst), .I(e[39]), .Q(
        ein[39]) );
  DFF \ereg_reg[40]  ( .D(ereg_next[40]), .CLK(clk), .RST(rst), .I(e[40]), .Q(
        ein[40]) );
  DFF \ereg_reg[41]  ( .D(ereg_next[41]), .CLK(clk), .RST(rst), .I(e[41]), .Q(
        ein[41]) );
  DFF \ereg_reg[42]  ( .D(ereg_next[42]), .CLK(clk), .RST(rst), .I(e[42]), .Q(
        ein[42]) );
  DFF \ereg_reg[43]  ( .D(ereg_next[43]), .CLK(clk), .RST(rst), .I(e[43]), .Q(
        ein[43]) );
  DFF \ereg_reg[44]  ( .D(ereg_next[44]), .CLK(clk), .RST(rst), .I(e[44]), .Q(
        ein[44]) );
  DFF \ereg_reg[45]  ( .D(ereg_next[45]), .CLK(clk), .RST(rst), .I(e[45]), .Q(
        ein[45]) );
  DFF \ereg_reg[46]  ( .D(ereg_next[46]), .CLK(clk), .RST(rst), .I(e[46]), .Q(
        ein[46]) );
  DFF \ereg_reg[47]  ( .D(ereg_next[47]), .CLK(clk), .RST(rst), .I(e[47]), .Q(
        ein[47]) );
  DFF \ereg_reg[48]  ( .D(ereg_next[48]), .CLK(clk), .RST(rst), .I(e[48]), .Q(
        ein[48]) );
  DFF \ereg_reg[49]  ( .D(ereg_next[49]), .CLK(clk), .RST(rst), .I(e[49]), .Q(
        ein[49]) );
  DFF \ereg_reg[50]  ( .D(ereg_next[50]), .CLK(clk), .RST(rst), .I(e[50]), .Q(
        ein[50]) );
  DFF \ereg_reg[51]  ( .D(ereg_next[51]), .CLK(clk), .RST(rst), .I(e[51]), .Q(
        ein[51]) );
  DFF \ereg_reg[52]  ( .D(ereg_next[52]), .CLK(clk), .RST(rst), .I(e[52]), .Q(
        ein[52]) );
  DFF \ereg_reg[53]  ( .D(ereg_next[53]), .CLK(clk), .RST(rst), .I(e[53]), .Q(
        ein[53]) );
  DFF \ereg_reg[54]  ( .D(ereg_next[54]), .CLK(clk), .RST(rst), .I(e[54]), .Q(
        ein[54]) );
  DFF \ereg_reg[55]  ( .D(ereg_next[55]), .CLK(clk), .RST(rst), .I(e[55]), .Q(
        ein[55]) );
  DFF \ereg_reg[56]  ( .D(ereg_next[56]), .CLK(clk), .RST(rst), .I(e[56]), .Q(
        ein[56]) );
  DFF \ereg_reg[57]  ( .D(ereg_next[57]), .CLK(clk), .RST(rst), .I(e[57]), .Q(
        ein[57]) );
  DFF \ereg_reg[58]  ( .D(ereg_next[58]), .CLK(clk), .RST(rst), .I(e[58]), .Q(
        ein[58]) );
  DFF \ereg_reg[59]  ( .D(ereg_next[59]), .CLK(clk), .RST(rst), .I(e[59]), .Q(
        ein[59]) );
  DFF \ereg_reg[60]  ( .D(ereg_next[60]), .CLK(clk), .RST(rst), .I(e[60]), .Q(
        ein[60]) );
  DFF \ereg_reg[61]  ( .D(ereg_next[61]), .CLK(clk), .RST(rst), .I(e[61]), .Q(
        ein[61]) );
  DFF \ereg_reg[62]  ( .D(ereg_next[62]), .CLK(clk), .RST(rst), .I(e[62]), .Q(
        ein[62]) );
  DFF \ereg_reg[63]  ( .D(ereg_next[63]), .CLK(clk), .RST(rst), .I(e[63]), .Q(
        ein[63]) );
  DFF \ereg_reg[64]  ( .D(ereg_next[64]), .CLK(clk), .RST(rst), .I(e[64]), .Q(
        ein[64]) );
  DFF \ereg_reg[65]  ( .D(ereg_next[65]), .CLK(clk), .RST(rst), .I(e[65]), .Q(
        ein[65]) );
  DFF \ereg_reg[66]  ( .D(ereg_next[66]), .CLK(clk), .RST(rst), .I(e[66]), .Q(
        ein[66]) );
  DFF \ereg_reg[67]  ( .D(ereg_next[67]), .CLK(clk), .RST(rst), .I(e[67]), .Q(
        ein[67]) );
  DFF \ereg_reg[68]  ( .D(ereg_next[68]), .CLK(clk), .RST(rst), .I(e[68]), .Q(
        ein[68]) );
  DFF \ereg_reg[69]  ( .D(ereg_next[69]), .CLK(clk), .RST(rst), .I(e[69]), .Q(
        ein[69]) );
  DFF \ereg_reg[70]  ( .D(ereg_next[70]), .CLK(clk), .RST(rst), .I(e[70]), .Q(
        ein[70]) );
  DFF \ereg_reg[71]  ( .D(ereg_next[71]), .CLK(clk), .RST(rst), .I(e[71]), .Q(
        ein[71]) );
  DFF \ereg_reg[72]  ( .D(ereg_next[72]), .CLK(clk), .RST(rst), .I(e[72]), .Q(
        ein[72]) );
  DFF \ereg_reg[73]  ( .D(ereg_next[73]), .CLK(clk), .RST(rst), .I(e[73]), .Q(
        ein[73]) );
  DFF \ereg_reg[74]  ( .D(ereg_next[74]), .CLK(clk), .RST(rst), .I(e[74]), .Q(
        ein[74]) );
  DFF \ereg_reg[75]  ( .D(ereg_next[75]), .CLK(clk), .RST(rst), .I(e[75]), .Q(
        ein[75]) );
  DFF \ereg_reg[76]  ( .D(ereg_next[76]), .CLK(clk), .RST(rst), .I(e[76]), .Q(
        ein[76]) );
  DFF \ereg_reg[77]  ( .D(ereg_next[77]), .CLK(clk), .RST(rst), .I(e[77]), .Q(
        ein[77]) );
  DFF \ereg_reg[78]  ( .D(ereg_next[78]), .CLK(clk), .RST(rst), .I(e[78]), .Q(
        ein[78]) );
  DFF \ereg_reg[79]  ( .D(ereg_next[79]), .CLK(clk), .RST(rst), .I(e[79]), .Q(
        ein[79]) );
  DFF \ereg_reg[80]  ( .D(ereg_next[80]), .CLK(clk), .RST(rst), .I(e[80]), .Q(
        ein[80]) );
  DFF \ereg_reg[81]  ( .D(ereg_next[81]), .CLK(clk), .RST(rst), .I(e[81]), .Q(
        ein[81]) );
  DFF \ereg_reg[82]  ( .D(ereg_next[82]), .CLK(clk), .RST(rst), .I(e[82]), .Q(
        ein[82]) );
  DFF \ereg_reg[83]  ( .D(ereg_next[83]), .CLK(clk), .RST(rst), .I(e[83]), .Q(
        ein[83]) );
  DFF \ereg_reg[84]  ( .D(ereg_next[84]), .CLK(clk), .RST(rst), .I(e[84]), .Q(
        ein[84]) );
  DFF \ereg_reg[85]  ( .D(ereg_next[85]), .CLK(clk), .RST(rst), .I(e[85]), .Q(
        ein[85]) );
  DFF \ereg_reg[86]  ( .D(ereg_next[86]), .CLK(clk), .RST(rst), .I(e[86]), .Q(
        ein[86]) );
  DFF \ereg_reg[87]  ( .D(ereg_next[87]), .CLK(clk), .RST(rst), .I(e[87]), .Q(
        ein[87]) );
  DFF \ereg_reg[88]  ( .D(ereg_next[88]), .CLK(clk), .RST(rst), .I(e[88]), .Q(
        ein[88]) );
  DFF \ereg_reg[89]  ( .D(ereg_next[89]), .CLK(clk), .RST(rst), .I(e[89]), .Q(
        ein[89]) );
  DFF \ereg_reg[90]  ( .D(ereg_next[90]), .CLK(clk), .RST(rst), .I(e[90]), .Q(
        ein[90]) );
  DFF \ereg_reg[91]  ( .D(ereg_next[91]), .CLK(clk), .RST(rst), .I(e[91]), .Q(
        ein[91]) );
  DFF \ereg_reg[92]  ( .D(ereg_next[92]), .CLK(clk), .RST(rst), .I(e[92]), .Q(
        ein[92]) );
  DFF \ereg_reg[93]  ( .D(ereg_next[93]), .CLK(clk), .RST(rst), .I(e[93]), .Q(
        ein[93]) );
  DFF \ereg_reg[94]  ( .D(ereg_next[94]), .CLK(clk), .RST(rst), .I(e[94]), .Q(
        ein[94]) );
  DFF \ereg_reg[95]  ( .D(ereg_next[95]), .CLK(clk), .RST(rst), .I(e[95]), .Q(
        ein[95]) );
  DFF \ereg_reg[96]  ( .D(ereg_next[96]), .CLK(clk), .RST(rst), .I(e[96]), .Q(
        ein[96]) );
  DFF \ereg_reg[97]  ( .D(ereg_next[97]), .CLK(clk), .RST(rst), .I(e[97]), .Q(
        ein[97]) );
  DFF \ereg_reg[98]  ( .D(ereg_next[98]), .CLK(clk), .RST(rst), .I(e[98]), .Q(
        ein[98]) );
  DFF \ereg_reg[99]  ( .D(ereg_next[99]), .CLK(clk), .RST(rst), .I(e[99]), .Q(
        ein[99]) );
  DFF \ereg_reg[100]  ( .D(ereg_next[100]), .CLK(clk), .RST(rst), .I(e[100]), 
        .Q(ein[100]) );
  DFF \ereg_reg[101]  ( .D(ereg_next[101]), .CLK(clk), .RST(rst), .I(e[101]), 
        .Q(ein[101]) );
  DFF \ereg_reg[102]  ( .D(ereg_next[102]), .CLK(clk), .RST(rst), .I(e[102]), 
        .Q(ein[102]) );
  DFF \ereg_reg[103]  ( .D(ereg_next[103]), .CLK(clk), .RST(rst), .I(e[103]), 
        .Q(ein[103]) );
  DFF \ereg_reg[104]  ( .D(ereg_next[104]), .CLK(clk), .RST(rst), .I(e[104]), 
        .Q(ein[104]) );
  DFF \ereg_reg[105]  ( .D(ereg_next[105]), .CLK(clk), .RST(rst), .I(e[105]), 
        .Q(ein[105]) );
  DFF \ereg_reg[106]  ( .D(ereg_next[106]), .CLK(clk), .RST(rst), .I(e[106]), 
        .Q(ein[106]) );
  DFF \ereg_reg[107]  ( .D(ereg_next[107]), .CLK(clk), .RST(rst), .I(e[107]), 
        .Q(ein[107]) );
  DFF \ereg_reg[108]  ( .D(ereg_next[108]), .CLK(clk), .RST(rst), .I(e[108]), 
        .Q(ein[108]) );
  DFF \ereg_reg[109]  ( .D(ereg_next[109]), .CLK(clk), .RST(rst), .I(e[109]), 
        .Q(ein[109]) );
  DFF \ereg_reg[110]  ( .D(ereg_next[110]), .CLK(clk), .RST(rst), .I(e[110]), 
        .Q(ein[110]) );
  DFF \ereg_reg[111]  ( .D(ereg_next[111]), .CLK(clk), .RST(rst), .I(e[111]), 
        .Q(ein[111]) );
  DFF \ereg_reg[112]  ( .D(ereg_next[112]), .CLK(clk), .RST(rst), .I(e[112]), 
        .Q(ein[112]) );
  DFF \ereg_reg[113]  ( .D(ereg_next[113]), .CLK(clk), .RST(rst), .I(e[113]), 
        .Q(ein[113]) );
  DFF \ereg_reg[114]  ( .D(ereg_next[114]), .CLK(clk), .RST(rst), .I(e[114]), 
        .Q(ein[114]) );
  DFF \ereg_reg[115]  ( .D(ereg_next[115]), .CLK(clk), .RST(rst), .I(e[115]), 
        .Q(ein[115]) );
  DFF \ereg_reg[116]  ( .D(ereg_next[116]), .CLK(clk), .RST(rst), .I(e[116]), 
        .Q(ein[116]) );
  DFF \ereg_reg[117]  ( .D(ereg_next[117]), .CLK(clk), .RST(rst), .I(e[117]), 
        .Q(ein[117]) );
  DFF \ereg_reg[118]  ( .D(ereg_next[118]), .CLK(clk), .RST(rst), .I(e[118]), 
        .Q(ein[118]) );
  DFF \ereg_reg[119]  ( .D(ereg_next[119]), .CLK(clk), .RST(rst), .I(e[119]), 
        .Q(ein[119]) );
  DFF \ereg_reg[120]  ( .D(ereg_next[120]), .CLK(clk), .RST(rst), .I(e[120]), 
        .Q(ein[120]) );
  DFF \ereg_reg[121]  ( .D(ereg_next[121]), .CLK(clk), .RST(rst), .I(e[121]), 
        .Q(ein[121]) );
  DFF \ereg_reg[122]  ( .D(ereg_next[122]), .CLK(clk), .RST(rst), .I(e[122]), 
        .Q(ein[122]) );
  DFF \ereg_reg[123]  ( .D(ereg_next[123]), .CLK(clk), .RST(rst), .I(e[123]), 
        .Q(ein[123]) );
  DFF \ereg_reg[124]  ( .D(ereg_next[124]), .CLK(clk), .RST(rst), .I(e[124]), 
        .Q(ein[124]) );
  DFF \ereg_reg[125]  ( .D(ereg_next[125]), .CLK(clk), .RST(rst), .I(e[125]), 
        .Q(ein[125]) );
  DFF \ereg_reg[126]  ( .D(ereg_next[126]), .CLK(clk), .RST(rst), .I(e[126]), 
        .Q(ein[126]) );
  DFF \ereg_reg[127]  ( .D(ereg_next[127]), .CLK(clk), .RST(rst), .I(e[127]), 
        .Q(ein[127]) );
  DFF \ereg_reg[128]  ( .D(ereg_next[128]), .CLK(clk), .RST(rst), .I(e[128]), 
        .Q(ein[128]) );
  DFF \ereg_reg[129]  ( .D(ereg_next[129]), .CLK(clk), .RST(rst), .I(e[129]), 
        .Q(ein[129]) );
  DFF \ereg_reg[130]  ( .D(ereg_next[130]), .CLK(clk), .RST(rst), .I(e[130]), 
        .Q(ein[130]) );
  DFF \ereg_reg[131]  ( .D(ereg_next[131]), .CLK(clk), .RST(rst), .I(e[131]), 
        .Q(ein[131]) );
  DFF \ereg_reg[132]  ( .D(ereg_next[132]), .CLK(clk), .RST(rst), .I(e[132]), 
        .Q(ein[132]) );
  DFF \ereg_reg[133]  ( .D(ereg_next[133]), .CLK(clk), .RST(rst), .I(e[133]), 
        .Q(ein[133]) );
  DFF \ereg_reg[134]  ( .D(ereg_next[134]), .CLK(clk), .RST(rst), .I(e[134]), 
        .Q(ein[134]) );
  DFF \ereg_reg[135]  ( .D(ereg_next[135]), .CLK(clk), .RST(rst), .I(e[135]), 
        .Q(ein[135]) );
  DFF \ereg_reg[136]  ( .D(ereg_next[136]), .CLK(clk), .RST(rst), .I(e[136]), 
        .Q(ein[136]) );
  DFF \ereg_reg[137]  ( .D(ereg_next[137]), .CLK(clk), .RST(rst), .I(e[137]), 
        .Q(ein[137]) );
  DFF \ereg_reg[138]  ( .D(ereg_next[138]), .CLK(clk), .RST(rst), .I(e[138]), 
        .Q(ein[138]) );
  DFF \ereg_reg[139]  ( .D(ereg_next[139]), .CLK(clk), .RST(rst), .I(e[139]), 
        .Q(ein[139]) );
  DFF \ereg_reg[140]  ( .D(ereg_next[140]), .CLK(clk), .RST(rst), .I(e[140]), 
        .Q(ein[140]) );
  DFF \ereg_reg[141]  ( .D(ereg_next[141]), .CLK(clk), .RST(rst), .I(e[141]), 
        .Q(ein[141]) );
  DFF \ereg_reg[142]  ( .D(ereg_next[142]), .CLK(clk), .RST(rst), .I(e[142]), 
        .Q(ein[142]) );
  DFF \ereg_reg[143]  ( .D(ereg_next[143]), .CLK(clk), .RST(rst), .I(e[143]), 
        .Q(ein[143]) );
  DFF \ereg_reg[144]  ( .D(ereg_next[144]), .CLK(clk), .RST(rst), .I(e[144]), 
        .Q(ein[144]) );
  DFF \ereg_reg[145]  ( .D(ereg_next[145]), .CLK(clk), .RST(rst), .I(e[145]), 
        .Q(ein[145]) );
  DFF \ereg_reg[146]  ( .D(ereg_next[146]), .CLK(clk), .RST(rst), .I(e[146]), 
        .Q(ein[146]) );
  DFF \ereg_reg[147]  ( .D(ereg_next[147]), .CLK(clk), .RST(rst), .I(e[147]), 
        .Q(ein[147]) );
  DFF \ereg_reg[148]  ( .D(ereg_next[148]), .CLK(clk), .RST(rst), .I(e[148]), 
        .Q(ein[148]) );
  DFF \ereg_reg[149]  ( .D(ereg_next[149]), .CLK(clk), .RST(rst), .I(e[149]), 
        .Q(ein[149]) );
  DFF \ereg_reg[150]  ( .D(ereg_next[150]), .CLK(clk), .RST(rst), .I(e[150]), 
        .Q(ein[150]) );
  DFF \ereg_reg[151]  ( .D(ereg_next[151]), .CLK(clk), .RST(rst), .I(e[151]), 
        .Q(ein[151]) );
  DFF \ereg_reg[152]  ( .D(ereg_next[152]), .CLK(clk), .RST(rst), .I(e[152]), 
        .Q(ein[152]) );
  DFF \ereg_reg[153]  ( .D(ereg_next[153]), .CLK(clk), .RST(rst), .I(e[153]), 
        .Q(ein[153]) );
  DFF \ereg_reg[154]  ( .D(ereg_next[154]), .CLK(clk), .RST(rst), .I(e[154]), 
        .Q(ein[154]) );
  DFF \ereg_reg[155]  ( .D(ereg_next[155]), .CLK(clk), .RST(rst), .I(e[155]), 
        .Q(ein[155]) );
  DFF \ereg_reg[156]  ( .D(ereg_next[156]), .CLK(clk), .RST(rst), .I(e[156]), 
        .Q(ein[156]) );
  DFF \ereg_reg[157]  ( .D(ereg_next[157]), .CLK(clk), .RST(rst), .I(e[157]), 
        .Q(ein[157]) );
  DFF \ereg_reg[158]  ( .D(ereg_next[158]), .CLK(clk), .RST(rst), .I(e[158]), 
        .Q(ein[158]) );
  DFF \ereg_reg[159]  ( .D(ereg_next[159]), .CLK(clk), .RST(rst), .I(e[159]), 
        .Q(ein[159]) );
  DFF \ereg_reg[160]  ( .D(ereg_next[160]), .CLK(clk), .RST(rst), .I(e[160]), 
        .Q(ein[160]) );
  DFF \ereg_reg[161]  ( .D(ereg_next[161]), .CLK(clk), .RST(rst), .I(e[161]), 
        .Q(ein[161]) );
  DFF \ereg_reg[162]  ( .D(ereg_next[162]), .CLK(clk), .RST(rst), .I(e[162]), 
        .Q(ein[162]) );
  DFF \ereg_reg[163]  ( .D(ereg_next[163]), .CLK(clk), .RST(rst), .I(e[163]), 
        .Q(ein[163]) );
  DFF \ereg_reg[164]  ( .D(ereg_next[164]), .CLK(clk), .RST(rst), .I(e[164]), 
        .Q(ein[164]) );
  DFF \ereg_reg[165]  ( .D(ereg_next[165]), .CLK(clk), .RST(rst), .I(e[165]), 
        .Q(ein[165]) );
  DFF \ereg_reg[166]  ( .D(ereg_next[166]), .CLK(clk), .RST(rst), .I(e[166]), 
        .Q(ein[166]) );
  DFF \ereg_reg[167]  ( .D(ereg_next[167]), .CLK(clk), .RST(rst), .I(e[167]), 
        .Q(ein[167]) );
  DFF \ereg_reg[168]  ( .D(ereg_next[168]), .CLK(clk), .RST(rst), .I(e[168]), 
        .Q(ein[168]) );
  DFF \ereg_reg[169]  ( .D(ereg_next[169]), .CLK(clk), .RST(rst), .I(e[169]), 
        .Q(ein[169]) );
  DFF \ereg_reg[170]  ( .D(ereg_next[170]), .CLK(clk), .RST(rst), .I(e[170]), 
        .Q(ein[170]) );
  DFF \ereg_reg[171]  ( .D(ereg_next[171]), .CLK(clk), .RST(rst), .I(e[171]), 
        .Q(ein[171]) );
  DFF \ereg_reg[172]  ( .D(ereg_next[172]), .CLK(clk), .RST(rst), .I(e[172]), 
        .Q(ein[172]) );
  DFF \ereg_reg[173]  ( .D(ereg_next[173]), .CLK(clk), .RST(rst), .I(e[173]), 
        .Q(ein[173]) );
  DFF \ereg_reg[174]  ( .D(ereg_next[174]), .CLK(clk), .RST(rst), .I(e[174]), 
        .Q(ein[174]) );
  DFF \ereg_reg[175]  ( .D(ereg_next[175]), .CLK(clk), .RST(rst), .I(e[175]), 
        .Q(ein[175]) );
  DFF \ereg_reg[176]  ( .D(ereg_next[176]), .CLK(clk), .RST(rst), .I(e[176]), 
        .Q(ein[176]) );
  DFF \ereg_reg[177]  ( .D(ereg_next[177]), .CLK(clk), .RST(rst), .I(e[177]), 
        .Q(ein[177]) );
  DFF \ereg_reg[178]  ( .D(ereg_next[178]), .CLK(clk), .RST(rst), .I(e[178]), 
        .Q(ein[178]) );
  DFF \ereg_reg[179]  ( .D(ereg_next[179]), .CLK(clk), .RST(rst), .I(e[179]), 
        .Q(ein[179]) );
  DFF \ereg_reg[180]  ( .D(ereg_next[180]), .CLK(clk), .RST(rst), .I(e[180]), 
        .Q(ein[180]) );
  DFF \ereg_reg[181]  ( .D(ereg_next[181]), .CLK(clk), .RST(rst), .I(e[181]), 
        .Q(ein[181]) );
  DFF \ereg_reg[182]  ( .D(ereg_next[182]), .CLK(clk), .RST(rst), .I(e[182]), 
        .Q(ein[182]) );
  DFF \ereg_reg[183]  ( .D(ereg_next[183]), .CLK(clk), .RST(rst), .I(e[183]), 
        .Q(ein[183]) );
  DFF \ereg_reg[184]  ( .D(ereg_next[184]), .CLK(clk), .RST(rst), .I(e[184]), 
        .Q(ein[184]) );
  DFF \ereg_reg[185]  ( .D(ereg_next[185]), .CLK(clk), .RST(rst), .I(e[185]), 
        .Q(ein[185]) );
  DFF \ereg_reg[186]  ( .D(ereg_next[186]), .CLK(clk), .RST(rst), .I(e[186]), 
        .Q(ein[186]) );
  DFF \ereg_reg[187]  ( .D(ereg_next[187]), .CLK(clk), .RST(rst), .I(e[187]), 
        .Q(ein[187]) );
  DFF \ereg_reg[188]  ( .D(ereg_next[188]), .CLK(clk), .RST(rst), .I(e[188]), 
        .Q(ein[188]) );
  DFF \ereg_reg[189]  ( .D(ereg_next[189]), .CLK(clk), .RST(rst), .I(e[189]), 
        .Q(ein[189]) );
  DFF \ereg_reg[190]  ( .D(ereg_next[190]), .CLK(clk), .RST(rst), .I(e[190]), 
        .Q(ein[190]) );
  DFF \ereg_reg[191]  ( .D(ereg_next[191]), .CLK(clk), .RST(rst), .I(e[191]), 
        .Q(ein[191]) );
  DFF \ereg_reg[192]  ( .D(ereg_next[192]), .CLK(clk), .RST(rst), .I(e[192]), 
        .Q(ein[192]) );
  DFF \ereg_reg[193]  ( .D(ereg_next[193]), .CLK(clk), .RST(rst), .I(e[193]), 
        .Q(ein[193]) );
  DFF \ereg_reg[194]  ( .D(ereg_next[194]), .CLK(clk), .RST(rst), .I(e[194]), 
        .Q(ein[194]) );
  DFF \ereg_reg[195]  ( .D(ereg_next[195]), .CLK(clk), .RST(rst), .I(e[195]), 
        .Q(ein[195]) );
  DFF \ereg_reg[196]  ( .D(ereg_next[196]), .CLK(clk), .RST(rst), .I(e[196]), 
        .Q(ein[196]) );
  DFF \ereg_reg[197]  ( .D(ereg_next[197]), .CLK(clk), .RST(rst), .I(e[197]), 
        .Q(ein[197]) );
  DFF \ereg_reg[198]  ( .D(ereg_next[198]), .CLK(clk), .RST(rst), .I(e[198]), 
        .Q(ein[198]) );
  DFF \ereg_reg[199]  ( .D(ereg_next[199]), .CLK(clk), .RST(rst), .I(e[199]), 
        .Q(ein[199]) );
  DFF \ereg_reg[200]  ( .D(ereg_next[200]), .CLK(clk), .RST(rst), .I(e[200]), 
        .Q(ein[200]) );
  DFF \ereg_reg[201]  ( .D(ereg_next[201]), .CLK(clk), .RST(rst), .I(e[201]), 
        .Q(ein[201]) );
  DFF \ereg_reg[202]  ( .D(ereg_next[202]), .CLK(clk), .RST(rst), .I(e[202]), 
        .Q(ein[202]) );
  DFF \ereg_reg[203]  ( .D(ereg_next[203]), .CLK(clk), .RST(rst), .I(e[203]), 
        .Q(ein[203]) );
  DFF \ereg_reg[204]  ( .D(ereg_next[204]), .CLK(clk), .RST(rst), .I(e[204]), 
        .Q(ein[204]) );
  DFF \ereg_reg[205]  ( .D(ereg_next[205]), .CLK(clk), .RST(rst), .I(e[205]), 
        .Q(ein[205]) );
  DFF \ereg_reg[206]  ( .D(ereg_next[206]), .CLK(clk), .RST(rst), .I(e[206]), 
        .Q(ein[206]) );
  DFF \ereg_reg[207]  ( .D(ereg_next[207]), .CLK(clk), .RST(rst), .I(e[207]), 
        .Q(ein[207]) );
  DFF \ereg_reg[208]  ( .D(ereg_next[208]), .CLK(clk), .RST(rst), .I(e[208]), 
        .Q(ein[208]) );
  DFF \ereg_reg[209]  ( .D(ereg_next[209]), .CLK(clk), .RST(rst), .I(e[209]), 
        .Q(ein[209]) );
  DFF \ereg_reg[210]  ( .D(ereg_next[210]), .CLK(clk), .RST(rst), .I(e[210]), 
        .Q(ein[210]) );
  DFF \ereg_reg[211]  ( .D(ereg_next[211]), .CLK(clk), .RST(rst), .I(e[211]), 
        .Q(ein[211]) );
  DFF \ereg_reg[212]  ( .D(ereg_next[212]), .CLK(clk), .RST(rst), .I(e[212]), 
        .Q(ein[212]) );
  DFF \ereg_reg[213]  ( .D(ereg_next[213]), .CLK(clk), .RST(rst), .I(e[213]), 
        .Q(ein[213]) );
  DFF \ereg_reg[214]  ( .D(ereg_next[214]), .CLK(clk), .RST(rst), .I(e[214]), 
        .Q(ein[214]) );
  DFF \ereg_reg[215]  ( .D(ereg_next[215]), .CLK(clk), .RST(rst), .I(e[215]), 
        .Q(ein[215]) );
  DFF \ereg_reg[216]  ( .D(ereg_next[216]), .CLK(clk), .RST(rst), .I(e[216]), 
        .Q(ein[216]) );
  DFF \ereg_reg[217]  ( .D(ereg_next[217]), .CLK(clk), .RST(rst), .I(e[217]), 
        .Q(ein[217]) );
  DFF \ereg_reg[218]  ( .D(ereg_next[218]), .CLK(clk), .RST(rst), .I(e[218]), 
        .Q(ein[218]) );
  DFF \ereg_reg[219]  ( .D(ereg_next[219]), .CLK(clk), .RST(rst), .I(e[219]), 
        .Q(ein[219]) );
  DFF \ereg_reg[220]  ( .D(ereg_next[220]), .CLK(clk), .RST(rst), .I(e[220]), 
        .Q(ein[220]) );
  DFF \ereg_reg[221]  ( .D(ereg_next[221]), .CLK(clk), .RST(rst), .I(e[221]), 
        .Q(ein[221]) );
  DFF \ereg_reg[222]  ( .D(ereg_next[222]), .CLK(clk), .RST(rst), .I(e[222]), 
        .Q(ein[222]) );
  DFF \ereg_reg[223]  ( .D(ereg_next[223]), .CLK(clk), .RST(rst), .I(e[223]), 
        .Q(ein[223]) );
  DFF \ereg_reg[224]  ( .D(ereg_next[224]), .CLK(clk), .RST(rst), .I(e[224]), 
        .Q(ein[224]) );
  DFF \ereg_reg[225]  ( .D(ereg_next[225]), .CLK(clk), .RST(rst), .I(e[225]), 
        .Q(ein[225]) );
  DFF \ereg_reg[226]  ( .D(ereg_next[226]), .CLK(clk), .RST(rst), .I(e[226]), 
        .Q(ein[226]) );
  DFF \ereg_reg[227]  ( .D(ereg_next[227]), .CLK(clk), .RST(rst), .I(e[227]), 
        .Q(ein[227]) );
  DFF \ereg_reg[228]  ( .D(ereg_next[228]), .CLK(clk), .RST(rst), .I(e[228]), 
        .Q(ein[228]) );
  DFF \ereg_reg[229]  ( .D(ereg_next[229]), .CLK(clk), .RST(rst), .I(e[229]), 
        .Q(ein[229]) );
  DFF \ereg_reg[230]  ( .D(ereg_next[230]), .CLK(clk), .RST(rst), .I(e[230]), 
        .Q(ein[230]) );
  DFF \ereg_reg[231]  ( .D(ereg_next[231]), .CLK(clk), .RST(rst), .I(e[231]), 
        .Q(ein[231]) );
  DFF \ereg_reg[232]  ( .D(ereg_next[232]), .CLK(clk), .RST(rst), .I(e[232]), 
        .Q(ein[232]) );
  DFF \ereg_reg[233]  ( .D(ereg_next[233]), .CLK(clk), .RST(rst), .I(e[233]), 
        .Q(ein[233]) );
  DFF \ereg_reg[234]  ( .D(ereg_next[234]), .CLK(clk), .RST(rst), .I(e[234]), 
        .Q(ein[234]) );
  DFF \ereg_reg[235]  ( .D(ereg_next[235]), .CLK(clk), .RST(rst), .I(e[235]), 
        .Q(ein[235]) );
  DFF \ereg_reg[236]  ( .D(ereg_next[236]), .CLK(clk), .RST(rst), .I(e[236]), 
        .Q(ein[236]) );
  DFF \ereg_reg[237]  ( .D(ereg_next[237]), .CLK(clk), .RST(rst), .I(e[237]), 
        .Q(ein[237]) );
  DFF \ereg_reg[238]  ( .D(ereg_next[238]), .CLK(clk), .RST(rst), .I(e[238]), 
        .Q(ein[238]) );
  DFF \ereg_reg[239]  ( .D(ereg_next[239]), .CLK(clk), .RST(rst), .I(e[239]), 
        .Q(ein[239]) );
  DFF \ereg_reg[240]  ( .D(ereg_next[240]), .CLK(clk), .RST(rst), .I(e[240]), 
        .Q(ein[240]) );
  DFF \ereg_reg[241]  ( .D(ereg_next[241]), .CLK(clk), .RST(rst), .I(e[241]), 
        .Q(ein[241]) );
  DFF \ereg_reg[242]  ( .D(ereg_next[242]), .CLK(clk), .RST(rst), .I(e[242]), 
        .Q(ein[242]) );
  DFF \ereg_reg[243]  ( .D(ereg_next[243]), .CLK(clk), .RST(rst), .I(e[243]), 
        .Q(ein[243]) );
  DFF \ereg_reg[244]  ( .D(ereg_next[244]), .CLK(clk), .RST(rst), .I(e[244]), 
        .Q(ein[244]) );
  DFF \ereg_reg[245]  ( .D(ereg_next[245]), .CLK(clk), .RST(rst), .I(e[245]), 
        .Q(ein[245]) );
  DFF \ereg_reg[246]  ( .D(ereg_next[246]), .CLK(clk), .RST(rst), .I(e[246]), 
        .Q(ein[246]) );
  DFF \ereg_reg[247]  ( .D(ereg_next[247]), .CLK(clk), .RST(rst), .I(e[247]), 
        .Q(ein[247]) );
  DFF \ereg_reg[248]  ( .D(ereg_next[248]), .CLK(clk), .RST(rst), .I(e[248]), 
        .Q(ein[248]) );
  DFF \ereg_reg[249]  ( .D(ereg_next[249]), .CLK(clk), .RST(rst), .I(e[249]), 
        .Q(ein[249]) );
  DFF \ereg_reg[250]  ( .D(ereg_next[250]), .CLK(clk), .RST(rst), .I(e[250]), 
        .Q(ein[250]) );
  DFF \ereg_reg[251]  ( .D(ereg_next[251]), .CLK(clk), .RST(rst), .I(e[251]), 
        .Q(ein[251]) );
  DFF \ereg_reg[252]  ( .D(ereg_next[252]), .CLK(clk), .RST(rst), .I(e[252]), 
        .Q(ein[252]) );
  DFF \ereg_reg[253]  ( .D(ereg_next[253]), .CLK(clk), .RST(rst), .I(e[253]), 
        .Q(ein[253]) );
  DFF \ereg_reg[254]  ( .D(ereg_next[254]), .CLK(clk), .RST(rst), .I(e[254]), 
        .Q(ein[254]) );
  DFF \ereg_reg[255]  ( .D(ereg_next[255]), .CLK(clk), .RST(rst), .I(e[255]), 
        .Q(ein[255]) );
  DFF first_one_reg ( .D(n6), .CLK(clk), .RST(rst), .I(1'b0), .Q(first_one) );
  DFF \creg_reg[0]  ( .D(creg_next[0]), .CLK(clk), .RST(rst), .I(m[0]), .Q(
        c[0]) );
  DFF \creg_reg[1]  ( .D(creg_next[1]), .CLK(clk), .RST(rst), .I(m[1]), .Q(
        c[1]) );
  DFF \creg_reg[2]  ( .D(creg_next[2]), .CLK(clk), .RST(rst), .I(m[2]), .Q(
        c[2]) );
  DFF \creg_reg[3]  ( .D(creg_next[3]), .CLK(clk), .RST(rst), .I(m[3]), .Q(
        c[3]) );
  DFF \creg_reg[4]  ( .D(creg_next[4]), .CLK(clk), .RST(rst), .I(m[4]), .Q(
        c[4]) );
  DFF \creg_reg[5]  ( .D(creg_next[5]), .CLK(clk), .RST(rst), .I(m[5]), .Q(
        c[5]) );
  DFF \creg_reg[6]  ( .D(creg_next[6]), .CLK(clk), .RST(rst), .I(m[6]), .Q(
        c[6]) );
  DFF \creg_reg[7]  ( .D(creg_next[7]), .CLK(clk), .RST(rst), .I(m[7]), .Q(
        c[7]) );
  DFF \creg_reg[8]  ( .D(creg_next[8]), .CLK(clk), .RST(rst), .I(m[8]), .Q(
        c[8]) );
  DFF \creg_reg[9]  ( .D(creg_next[9]), .CLK(clk), .RST(rst), .I(m[9]), .Q(
        c[9]) );
  DFF \creg_reg[10]  ( .D(creg_next[10]), .CLK(clk), .RST(rst), .I(m[10]), .Q(
        c[10]) );
  DFF \creg_reg[11]  ( .D(creg_next[11]), .CLK(clk), .RST(rst), .I(m[11]), .Q(
        c[11]) );
  DFF \creg_reg[12]  ( .D(creg_next[12]), .CLK(clk), .RST(rst), .I(m[12]), .Q(
        c[12]) );
  DFF \creg_reg[13]  ( .D(creg_next[13]), .CLK(clk), .RST(rst), .I(m[13]), .Q(
        c[13]) );
  DFF \creg_reg[14]  ( .D(creg_next[14]), .CLK(clk), .RST(rst), .I(m[14]), .Q(
        c[14]) );
  DFF \creg_reg[15]  ( .D(creg_next[15]), .CLK(clk), .RST(rst), .I(m[15]), .Q(
        c[15]) );
  DFF \creg_reg[16]  ( .D(creg_next[16]), .CLK(clk), .RST(rst), .I(m[16]), .Q(
        c[16]) );
  DFF \creg_reg[17]  ( .D(creg_next[17]), .CLK(clk), .RST(rst), .I(m[17]), .Q(
        c[17]) );
  DFF \creg_reg[18]  ( .D(creg_next[18]), .CLK(clk), .RST(rst), .I(m[18]), .Q(
        c[18]) );
  DFF \creg_reg[19]  ( .D(creg_next[19]), .CLK(clk), .RST(rst), .I(m[19]), .Q(
        c[19]) );
  DFF \creg_reg[20]  ( .D(creg_next[20]), .CLK(clk), .RST(rst), .I(m[20]), .Q(
        c[20]) );
  DFF \creg_reg[21]  ( .D(creg_next[21]), .CLK(clk), .RST(rst), .I(m[21]), .Q(
        c[21]) );
  DFF \creg_reg[22]  ( .D(creg_next[22]), .CLK(clk), .RST(rst), .I(m[22]), .Q(
        c[22]) );
  DFF \creg_reg[23]  ( .D(creg_next[23]), .CLK(clk), .RST(rst), .I(m[23]), .Q(
        c[23]) );
  DFF \creg_reg[24]  ( .D(creg_next[24]), .CLK(clk), .RST(rst), .I(m[24]), .Q(
        c[24]) );
  DFF \creg_reg[25]  ( .D(creg_next[25]), .CLK(clk), .RST(rst), .I(m[25]), .Q(
        c[25]) );
  DFF \creg_reg[26]  ( .D(creg_next[26]), .CLK(clk), .RST(rst), .I(m[26]), .Q(
        c[26]) );
  DFF \creg_reg[27]  ( .D(creg_next[27]), .CLK(clk), .RST(rst), .I(m[27]), .Q(
        c[27]) );
  DFF \creg_reg[28]  ( .D(creg_next[28]), .CLK(clk), .RST(rst), .I(m[28]), .Q(
        c[28]) );
  DFF \creg_reg[29]  ( .D(creg_next[29]), .CLK(clk), .RST(rst), .I(m[29]), .Q(
        c[29]) );
  DFF \creg_reg[30]  ( .D(creg_next[30]), .CLK(clk), .RST(rst), .I(m[30]), .Q(
        c[30]) );
  DFF \creg_reg[31]  ( .D(creg_next[31]), .CLK(clk), .RST(rst), .I(m[31]), .Q(
        c[31]) );
  DFF \creg_reg[32]  ( .D(creg_next[32]), .CLK(clk), .RST(rst), .I(m[32]), .Q(
        c[32]) );
  DFF \creg_reg[33]  ( .D(creg_next[33]), .CLK(clk), .RST(rst), .I(m[33]), .Q(
        c[33]) );
  DFF \creg_reg[34]  ( .D(creg_next[34]), .CLK(clk), .RST(rst), .I(m[34]), .Q(
        c[34]) );
  DFF \creg_reg[35]  ( .D(creg_next[35]), .CLK(clk), .RST(rst), .I(m[35]), .Q(
        c[35]) );
  DFF \creg_reg[36]  ( .D(creg_next[36]), .CLK(clk), .RST(rst), .I(m[36]), .Q(
        c[36]) );
  DFF \creg_reg[37]  ( .D(creg_next[37]), .CLK(clk), .RST(rst), .I(m[37]), .Q(
        c[37]) );
  DFF \creg_reg[38]  ( .D(creg_next[38]), .CLK(clk), .RST(rst), .I(m[38]), .Q(
        c[38]) );
  DFF \creg_reg[39]  ( .D(creg_next[39]), .CLK(clk), .RST(rst), .I(m[39]), .Q(
        c[39]) );
  DFF \creg_reg[40]  ( .D(creg_next[40]), .CLK(clk), .RST(rst), .I(m[40]), .Q(
        c[40]) );
  DFF \creg_reg[41]  ( .D(creg_next[41]), .CLK(clk), .RST(rst), .I(m[41]), .Q(
        c[41]) );
  DFF \creg_reg[42]  ( .D(creg_next[42]), .CLK(clk), .RST(rst), .I(m[42]), .Q(
        c[42]) );
  DFF \creg_reg[43]  ( .D(creg_next[43]), .CLK(clk), .RST(rst), .I(m[43]), .Q(
        c[43]) );
  DFF \creg_reg[44]  ( .D(creg_next[44]), .CLK(clk), .RST(rst), .I(m[44]), .Q(
        c[44]) );
  DFF \creg_reg[45]  ( .D(creg_next[45]), .CLK(clk), .RST(rst), .I(m[45]), .Q(
        c[45]) );
  DFF \creg_reg[46]  ( .D(creg_next[46]), .CLK(clk), .RST(rst), .I(m[46]), .Q(
        c[46]) );
  DFF \creg_reg[47]  ( .D(creg_next[47]), .CLK(clk), .RST(rst), .I(m[47]), .Q(
        c[47]) );
  DFF \creg_reg[48]  ( .D(creg_next[48]), .CLK(clk), .RST(rst), .I(m[48]), .Q(
        c[48]) );
  DFF \creg_reg[49]  ( .D(creg_next[49]), .CLK(clk), .RST(rst), .I(m[49]), .Q(
        c[49]) );
  DFF \creg_reg[50]  ( .D(creg_next[50]), .CLK(clk), .RST(rst), .I(m[50]), .Q(
        c[50]) );
  DFF \creg_reg[51]  ( .D(creg_next[51]), .CLK(clk), .RST(rst), .I(m[51]), .Q(
        c[51]) );
  DFF \creg_reg[52]  ( .D(creg_next[52]), .CLK(clk), .RST(rst), .I(m[52]), .Q(
        c[52]) );
  DFF \creg_reg[53]  ( .D(creg_next[53]), .CLK(clk), .RST(rst), .I(m[53]), .Q(
        c[53]) );
  DFF \creg_reg[54]  ( .D(creg_next[54]), .CLK(clk), .RST(rst), .I(m[54]), .Q(
        c[54]) );
  DFF \creg_reg[55]  ( .D(creg_next[55]), .CLK(clk), .RST(rst), .I(m[55]), .Q(
        c[55]) );
  DFF \creg_reg[56]  ( .D(creg_next[56]), .CLK(clk), .RST(rst), .I(m[56]), .Q(
        c[56]) );
  DFF \creg_reg[57]  ( .D(creg_next[57]), .CLK(clk), .RST(rst), .I(m[57]), .Q(
        c[57]) );
  DFF \creg_reg[58]  ( .D(creg_next[58]), .CLK(clk), .RST(rst), .I(m[58]), .Q(
        c[58]) );
  DFF \creg_reg[59]  ( .D(creg_next[59]), .CLK(clk), .RST(rst), .I(m[59]), .Q(
        c[59]) );
  DFF \creg_reg[60]  ( .D(creg_next[60]), .CLK(clk), .RST(rst), .I(m[60]), .Q(
        c[60]) );
  DFF \creg_reg[61]  ( .D(creg_next[61]), .CLK(clk), .RST(rst), .I(m[61]), .Q(
        c[61]) );
  DFF \creg_reg[62]  ( .D(creg_next[62]), .CLK(clk), .RST(rst), .I(m[62]), .Q(
        c[62]) );
  DFF \creg_reg[63]  ( .D(creg_next[63]), .CLK(clk), .RST(rst), .I(m[63]), .Q(
        c[63]) );
  DFF \creg_reg[64]  ( .D(creg_next[64]), .CLK(clk), .RST(rst), .I(m[64]), .Q(
        c[64]) );
  DFF \creg_reg[65]  ( .D(creg_next[65]), .CLK(clk), .RST(rst), .I(m[65]), .Q(
        c[65]) );
  DFF \creg_reg[66]  ( .D(creg_next[66]), .CLK(clk), .RST(rst), .I(m[66]), .Q(
        c[66]) );
  DFF \creg_reg[67]  ( .D(creg_next[67]), .CLK(clk), .RST(rst), .I(m[67]), .Q(
        c[67]) );
  DFF \creg_reg[68]  ( .D(creg_next[68]), .CLK(clk), .RST(rst), .I(m[68]), .Q(
        c[68]) );
  DFF \creg_reg[69]  ( .D(creg_next[69]), .CLK(clk), .RST(rst), .I(m[69]), .Q(
        c[69]) );
  DFF \creg_reg[70]  ( .D(creg_next[70]), .CLK(clk), .RST(rst), .I(m[70]), .Q(
        c[70]) );
  DFF \creg_reg[71]  ( .D(creg_next[71]), .CLK(clk), .RST(rst), .I(m[71]), .Q(
        c[71]) );
  DFF \creg_reg[72]  ( .D(creg_next[72]), .CLK(clk), .RST(rst), .I(m[72]), .Q(
        c[72]) );
  DFF \creg_reg[73]  ( .D(creg_next[73]), .CLK(clk), .RST(rst), .I(m[73]), .Q(
        c[73]) );
  DFF \creg_reg[74]  ( .D(creg_next[74]), .CLK(clk), .RST(rst), .I(m[74]), .Q(
        c[74]) );
  DFF \creg_reg[75]  ( .D(creg_next[75]), .CLK(clk), .RST(rst), .I(m[75]), .Q(
        c[75]) );
  DFF \creg_reg[76]  ( .D(creg_next[76]), .CLK(clk), .RST(rst), .I(m[76]), .Q(
        c[76]) );
  DFF \creg_reg[77]  ( .D(creg_next[77]), .CLK(clk), .RST(rst), .I(m[77]), .Q(
        c[77]) );
  DFF \creg_reg[78]  ( .D(creg_next[78]), .CLK(clk), .RST(rst), .I(m[78]), .Q(
        c[78]) );
  DFF \creg_reg[79]  ( .D(creg_next[79]), .CLK(clk), .RST(rst), .I(m[79]), .Q(
        c[79]) );
  DFF \creg_reg[80]  ( .D(creg_next[80]), .CLK(clk), .RST(rst), .I(m[80]), .Q(
        c[80]) );
  DFF \creg_reg[81]  ( .D(creg_next[81]), .CLK(clk), .RST(rst), .I(m[81]), .Q(
        c[81]) );
  DFF \creg_reg[82]  ( .D(creg_next[82]), .CLK(clk), .RST(rst), .I(m[82]), .Q(
        c[82]) );
  DFF \creg_reg[83]  ( .D(creg_next[83]), .CLK(clk), .RST(rst), .I(m[83]), .Q(
        c[83]) );
  DFF \creg_reg[84]  ( .D(creg_next[84]), .CLK(clk), .RST(rst), .I(m[84]), .Q(
        c[84]) );
  DFF \creg_reg[85]  ( .D(creg_next[85]), .CLK(clk), .RST(rst), .I(m[85]), .Q(
        c[85]) );
  DFF \creg_reg[86]  ( .D(creg_next[86]), .CLK(clk), .RST(rst), .I(m[86]), .Q(
        c[86]) );
  DFF \creg_reg[87]  ( .D(creg_next[87]), .CLK(clk), .RST(rst), .I(m[87]), .Q(
        c[87]) );
  DFF \creg_reg[88]  ( .D(creg_next[88]), .CLK(clk), .RST(rst), .I(m[88]), .Q(
        c[88]) );
  DFF \creg_reg[89]  ( .D(creg_next[89]), .CLK(clk), .RST(rst), .I(m[89]), .Q(
        c[89]) );
  DFF \creg_reg[90]  ( .D(creg_next[90]), .CLK(clk), .RST(rst), .I(m[90]), .Q(
        c[90]) );
  DFF \creg_reg[91]  ( .D(creg_next[91]), .CLK(clk), .RST(rst), .I(m[91]), .Q(
        c[91]) );
  DFF \creg_reg[92]  ( .D(creg_next[92]), .CLK(clk), .RST(rst), .I(m[92]), .Q(
        c[92]) );
  DFF \creg_reg[93]  ( .D(creg_next[93]), .CLK(clk), .RST(rst), .I(m[93]), .Q(
        c[93]) );
  DFF \creg_reg[94]  ( .D(creg_next[94]), .CLK(clk), .RST(rst), .I(m[94]), .Q(
        c[94]) );
  DFF \creg_reg[95]  ( .D(creg_next[95]), .CLK(clk), .RST(rst), .I(m[95]), .Q(
        c[95]) );
  DFF \creg_reg[96]  ( .D(creg_next[96]), .CLK(clk), .RST(rst), .I(m[96]), .Q(
        c[96]) );
  DFF \creg_reg[97]  ( .D(creg_next[97]), .CLK(clk), .RST(rst), .I(m[97]), .Q(
        c[97]) );
  DFF \creg_reg[98]  ( .D(creg_next[98]), .CLK(clk), .RST(rst), .I(m[98]), .Q(
        c[98]) );
  DFF \creg_reg[99]  ( .D(creg_next[99]), .CLK(clk), .RST(rst), .I(m[99]), .Q(
        c[99]) );
  DFF \creg_reg[100]  ( .D(creg_next[100]), .CLK(clk), .RST(rst), .I(m[100]), 
        .Q(c[100]) );
  DFF \creg_reg[101]  ( .D(creg_next[101]), .CLK(clk), .RST(rst), .I(m[101]), 
        .Q(c[101]) );
  DFF \creg_reg[102]  ( .D(creg_next[102]), .CLK(clk), .RST(rst), .I(m[102]), 
        .Q(c[102]) );
  DFF \creg_reg[103]  ( .D(creg_next[103]), .CLK(clk), .RST(rst), .I(m[103]), 
        .Q(c[103]) );
  DFF \creg_reg[104]  ( .D(creg_next[104]), .CLK(clk), .RST(rst), .I(m[104]), 
        .Q(c[104]) );
  DFF \creg_reg[105]  ( .D(creg_next[105]), .CLK(clk), .RST(rst), .I(m[105]), 
        .Q(c[105]) );
  DFF \creg_reg[106]  ( .D(creg_next[106]), .CLK(clk), .RST(rst), .I(m[106]), 
        .Q(c[106]) );
  DFF \creg_reg[107]  ( .D(creg_next[107]), .CLK(clk), .RST(rst), .I(m[107]), 
        .Q(c[107]) );
  DFF \creg_reg[108]  ( .D(creg_next[108]), .CLK(clk), .RST(rst), .I(m[108]), 
        .Q(c[108]) );
  DFF \creg_reg[109]  ( .D(creg_next[109]), .CLK(clk), .RST(rst), .I(m[109]), 
        .Q(c[109]) );
  DFF \creg_reg[110]  ( .D(creg_next[110]), .CLK(clk), .RST(rst), .I(m[110]), 
        .Q(c[110]) );
  DFF \creg_reg[111]  ( .D(creg_next[111]), .CLK(clk), .RST(rst), .I(m[111]), 
        .Q(c[111]) );
  DFF \creg_reg[112]  ( .D(creg_next[112]), .CLK(clk), .RST(rst), .I(m[112]), 
        .Q(c[112]) );
  DFF \creg_reg[113]  ( .D(creg_next[113]), .CLK(clk), .RST(rst), .I(m[113]), 
        .Q(c[113]) );
  DFF \creg_reg[114]  ( .D(creg_next[114]), .CLK(clk), .RST(rst), .I(m[114]), 
        .Q(c[114]) );
  DFF \creg_reg[115]  ( .D(creg_next[115]), .CLK(clk), .RST(rst), .I(m[115]), 
        .Q(c[115]) );
  DFF \creg_reg[116]  ( .D(creg_next[116]), .CLK(clk), .RST(rst), .I(m[116]), 
        .Q(c[116]) );
  DFF \creg_reg[117]  ( .D(creg_next[117]), .CLK(clk), .RST(rst), .I(m[117]), 
        .Q(c[117]) );
  DFF \creg_reg[118]  ( .D(creg_next[118]), .CLK(clk), .RST(rst), .I(m[118]), 
        .Q(c[118]) );
  DFF \creg_reg[119]  ( .D(creg_next[119]), .CLK(clk), .RST(rst), .I(m[119]), 
        .Q(c[119]) );
  DFF \creg_reg[120]  ( .D(creg_next[120]), .CLK(clk), .RST(rst), .I(m[120]), 
        .Q(c[120]) );
  DFF \creg_reg[121]  ( .D(creg_next[121]), .CLK(clk), .RST(rst), .I(m[121]), 
        .Q(c[121]) );
  DFF \creg_reg[122]  ( .D(creg_next[122]), .CLK(clk), .RST(rst), .I(m[122]), 
        .Q(c[122]) );
  DFF \creg_reg[123]  ( .D(creg_next[123]), .CLK(clk), .RST(rst), .I(m[123]), 
        .Q(c[123]) );
  DFF \creg_reg[124]  ( .D(creg_next[124]), .CLK(clk), .RST(rst), .I(m[124]), 
        .Q(c[124]) );
  DFF \creg_reg[125]  ( .D(creg_next[125]), .CLK(clk), .RST(rst), .I(m[125]), 
        .Q(c[125]) );
  DFF \creg_reg[126]  ( .D(creg_next[126]), .CLK(clk), .RST(rst), .I(m[126]), 
        .Q(c[126]) );
  DFF \creg_reg[127]  ( .D(creg_next[127]), .CLK(clk), .RST(rst), .I(m[127]), 
        .Q(c[127]) );
  DFF \creg_reg[128]  ( .D(creg_next[128]), .CLK(clk), .RST(rst), .I(m[128]), 
        .Q(c[128]) );
  DFF \creg_reg[129]  ( .D(creg_next[129]), .CLK(clk), .RST(rst), .I(m[129]), 
        .Q(c[129]) );
  DFF \creg_reg[130]  ( .D(creg_next[130]), .CLK(clk), .RST(rst), .I(m[130]), 
        .Q(c[130]) );
  DFF \creg_reg[131]  ( .D(creg_next[131]), .CLK(clk), .RST(rst), .I(m[131]), 
        .Q(c[131]) );
  DFF \creg_reg[132]  ( .D(creg_next[132]), .CLK(clk), .RST(rst), .I(m[132]), 
        .Q(c[132]) );
  DFF \creg_reg[133]  ( .D(creg_next[133]), .CLK(clk), .RST(rst), .I(m[133]), 
        .Q(c[133]) );
  DFF \creg_reg[134]  ( .D(creg_next[134]), .CLK(clk), .RST(rst), .I(m[134]), 
        .Q(c[134]) );
  DFF \creg_reg[135]  ( .D(creg_next[135]), .CLK(clk), .RST(rst), .I(m[135]), 
        .Q(c[135]) );
  DFF \creg_reg[136]  ( .D(creg_next[136]), .CLK(clk), .RST(rst), .I(m[136]), 
        .Q(c[136]) );
  DFF \creg_reg[137]  ( .D(creg_next[137]), .CLK(clk), .RST(rst), .I(m[137]), 
        .Q(c[137]) );
  DFF \creg_reg[138]  ( .D(creg_next[138]), .CLK(clk), .RST(rst), .I(m[138]), 
        .Q(c[138]) );
  DFF \creg_reg[139]  ( .D(creg_next[139]), .CLK(clk), .RST(rst), .I(m[139]), 
        .Q(c[139]) );
  DFF \creg_reg[140]  ( .D(creg_next[140]), .CLK(clk), .RST(rst), .I(m[140]), 
        .Q(c[140]) );
  DFF \creg_reg[141]  ( .D(creg_next[141]), .CLK(clk), .RST(rst), .I(m[141]), 
        .Q(c[141]) );
  DFF \creg_reg[142]  ( .D(creg_next[142]), .CLK(clk), .RST(rst), .I(m[142]), 
        .Q(c[142]) );
  DFF \creg_reg[143]  ( .D(creg_next[143]), .CLK(clk), .RST(rst), .I(m[143]), 
        .Q(c[143]) );
  DFF \creg_reg[144]  ( .D(creg_next[144]), .CLK(clk), .RST(rst), .I(m[144]), 
        .Q(c[144]) );
  DFF \creg_reg[145]  ( .D(creg_next[145]), .CLK(clk), .RST(rst), .I(m[145]), 
        .Q(c[145]) );
  DFF \creg_reg[146]  ( .D(creg_next[146]), .CLK(clk), .RST(rst), .I(m[146]), 
        .Q(c[146]) );
  DFF \creg_reg[147]  ( .D(creg_next[147]), .CLK(clk), .RST(rst), .I(m[147]), 
        .Q(c[147]) );
  DFF \creg_reg[148]  ( .D(creg_next[148]), .CLK(clk), .RST(rst), .I(m[148]), 
        .Q(c[148]) );
  DFF \creg_reg[149]  ( .D(creg_next[149]), .CLK(clk), .RST(rst), .I(m[149]), 
        .Q(c[149]) );
  DFF \creg_reg[150]  ( .D(creg_next[150]), .CLK(clk), .RST(rst), .I(m[150]), 
        .Q(c[150]) );
  DFF \creg_reg[151]  ( .D(creg_next[151]), .CLK(clk), .RST(rst), .I(m[151]), 
        .Q(c[151]) );
  DFF \creg_reg[152]  ( .D(creg_next[152]), .CLK(clk), .RST(rst), .I(m[152]), 
        .Q(c[152]) );
  DFF \creg_reg[153]  ( .D(creg_next[153]), .CLK(clk), .RST(rst), .I(m[153]), 
        .Q(c[153]) );
  DFF \creg_reg[154]  ( .D(creg_next[154]), .CLK(clk), .RST(rst), .I(m[154]), 
        .Q(c[154]) );
  DFF \creg_reg[155]  ( .D(creg_next[155]), .CLK(clk), .RST(rst), .I(m[155]), 
        .Q(c[155]) );
  DFF \creg_reg[156]  ( .D(creg_next[156]), .CLK(clk), .RST(rst), .I(m[156]), 
        .Q(c[156]) );
  DFF \creg_reg[157]  ( .D(creg_next[157]), .CLK(clk), .RST(rst), .I(m[157]), 
        .Q(c[157]) );
  DFF \creg_reg[158]  ( .D(creg_next[158]), .CLK(clk), .RST(rst), .I(m[158]), 
        .Q(c[158]) );
  DFF \creg_reg[159]  ( .D(creg_next[159]), .CLK(clk), .RST(rst), .I(m[159]), 
        .Q(c[159]) );
  DFF \creg_reg[160]  ( .D(creg_next[160]), .CLK(clk), .RST(rst), .I(m[160]), 
        .Q(c[160]) );
  DFF \creg_reg[161]  ( .D(creg_next[161]), .CLK(clk), .RST(rst), .I(m[161]), 
        .Q(c[161]) );
  DFF \creg_reg[162]  ( .D(creg_next[162]), .CLK(clk), .RST(rst), .I(m[162]), 
        .Q(c[162]) );
  DFF \creg_reg[163]  ( .D(creg_next[163]), .CLK(clk), .RST(rst), .I(m[163]), 
        .Q(c[163]) );
  DFF \creg_reg[164]  ( .D(creg_next[164]), .CLK(clk), .RST(rst), .I(m[164]), 
        .Q(c[164]) );
  DFF \creg_reg[165]  ( .D(creg_next[165]), .CLK(clk), .RST(rst), .I(m[165]), 
        .Q(c[165]) );
  DFF \creg_reg[166]  ( .D(creg_next[166]), .CLK(clk), .RST(rst), .I(m[166]), 
        .Q(c[166]) );
  DFF \creg_reg[167]  ( .D(creg_next[167]), .CLK(clk), .RST(rst), .I(m[167]), 
        .Q(c[167]) );
  DFF \creg_reg[168]  ( .D(creg_next[168]), .CLK(clk), .RST(rst), .I(m[168]), 
        .Q(c[168]) );
  DFF \creg_reg[169]  ( .D(creg_next[169]), .CLK(clk), .RST(rst), .I(m[169]), 
        .Q(c[169]) );
  DFF \creg_reg[170]  ( .D(creg_next[170]), .CLK(clk), .RST(rst), .I(m[170]), 
        .Q(c[170]) );
  DFF \creg_reg[171]  ( .D(creg_next[171]), .CLK(clk), .RST(rst), .I(m[171]), 
        .Q(c[171]) );
  DFF \creg_reg[172]  ( .D(creg_next[172]), .CLK(clk), .RST(rst), .I(m[172]), 
        .Q(c[172]) );
  DFF \creg_reg[173]  ( .D(creg_next[173]), .CLK(clk), .RST(rst), .I(m[173]), 
        .Q(c[173]) );
  DFF \creg_reg[174]  ( .D(creg_next[174]), .CLK(clk), .RST(rst), .I(m[174]), 
        .Q(c[174]) );
  DFF \creg_reg[175]  ( .D(creg_next[175]), .CLK(clk), .RST(rst), .I(m[175]), 
        .Q(c[175]) );
  DFF \creg_reg[176]  ( .D(creg_next[176]), .CLK(clk), .RST(rst), .I(m[176]), 
        .Q(c[176]) );
  DFF \creg_reg[177]  ( .D(creg_next[177]), .CLK(clk), .RST(rst), .I(m[177]), 
        .Q(c[177]) );
  DFF \creg_reg[178]  ( .D(creg_next[178]), .CLK(clk), .RST(rst), .I(m[178]), 
        .Q(c[178]) );
  DFF \creg_reg[179]  ( .D(creg_next[179]), .CLK(clk), .RST(rst), .I(m[179]), 
        .Q(c[179]) );
  DFF \creg_reg[180]  ( .D(creg_next[180]), .CLK(clk), .RST(rst), .I(m[180]), 
        .Q(c[180]) );
  DFF \creg_reg[181]  ( .D(creg_next[181]), .CLK(clk), .RST(rst), .I(m[181]), 
        .Q(c[181]) );
  DFF \creg_reg[182]  ( .D(creg_next[182]), .CLK(clk), .RST(rst), .I(m[182]), 
        .Q(c[182]) );
  DFF \creg_reg[183]  ( .D(creg_next[183]), .CLK(clk), .RST(rst), .I(m[183]), 
        .Q(c[183]) );
  DFF \creg_reg[184]  ( .D(creg_next[184]), .CLK(clk), .RST(rst), .I(m[184]), 
        .Q(c[184]) );
  DFF \creg_reg[185]  ( .D(creg_next[185]), .CLK(clk), .RST(rst), .I(m[185]), 
        .Q(c[185]) );
  DFF \creg_reg[186]  ( .D(creg_next[186]), .CLK(clk), .RST(rst), .I(m[186]), 
        .Q(c[186]) );
  DFF \creg_reg[187]  ( .D(creg_next[187]), .CLK(clk), .RST(rst), .I(m[187]), 
        .Q(c[187]) );
  DFF \creg_reg[188]  ( .D(creg_next[188]), .CLK(clk), .RST(rst), .I(m[188]), 
        .Q(c[188]) );
  DFF \creg_reg[189]  ( .D(creg_next[189]), .CLK(clk), .RST(rst), .I(m[189]), 
        .Q(c[189]) );
  DFF \creg_reg[190]  ( .D(creg_next[190]), .CLK(clk), .RST(rst), .I(m[190]), 
        .Q(c[190]) );
  DFF \creg_reg[191]  ( .D(creg_next[191]), .CLK(clk), .RST(rst), .I(m[191]), 
        .Q(c[191]) );
  DFF \creg_reg[192]  ( .D(creg_next[192]), .CLK(clk), .RST(rst), .I(m[192]), 
        .Q(c[192]) );
  DFF \creg_reg[193]  ( .D(creg_next[193]), .CLK(clk), .RST(rst), .I(m[193]), 
        .Q(c[193]) );
  DFF \creg_reg[194]  ( .D(creg_next[194]), .CLK(clk), .RST(rst), .I(m[194]), 
        .Q(c[194]) );
  DFF \creg_reg[195]  ( .D(creg_next[195]), .CLK(clk), .RST(rst), .I(m[195]), 
        .Q(c[195]) );
  DFF \creg_reg[196]  ( .D(creg_next[196]), .CLK(clk), .RST(rst), .I(m[196]), 
        .Q(c[196]) );
  DFF \creg_reg[197]  ( .D(creg_next[197]), .CLK(clk), .RST(rst), .I(m[197]), 
        .Q(c[197]) );
  DFF \creg_reg[198]  ( .D(creg_next[198]), .CLK(clk), .RST(rst), .I(m[198]), 
        .Q(c[198]) );
  DFF \creg_reg[199]  ( .D(creg_next[199]), .CLK(clk), .RST(rst), .I(m[199]), 
        .Q(c[199]) );
  DFF \creg_reg[200]  ( .D(creg_next[200]), .CLK(clk), .RST(rst), .I(m[200]), 
        .Q(c[200]) );
  DFF \creg_reg[201]  ( .D(creg_next[201]), .CLK(clk), .RST(rst), .I(m[201]), 
        .Q(c[201]) );
  DFF \creg_reg[202]  ( .D(creg_next[202]), .CLK(clk), .RST(rst), .I(m[202]), 
        .Q(c[202]) );
  DFF \creg_reg[203]  ( .D(creg_next[203]), .CLK(clk), .RST(rst), .I(m[203]), 
        .Q(c[203]) );
  DFF \creg_reg[204]  ( .D(creg_next[204]), .CLK(clk), .RST(rst), .I(m[204]), 
        .Q(c[204]) );
  DFF \creg_reg[205]  ( .D(creg_next[205]), .CLK(clk), .RST(rst), .I(m[205]), 
        .Q(c[205]) );
  DFF \creg_reg[206]  ( .D(creg_next[206]), .CLK(clk), .RST(rst), .I(m[206]), 
        .Q(c[206]) );
  DFF \creg_reg[207]  ( .D(creg_next[207]), .CLK(clk), .RST(rst), .I(m[207]), 
        .Q(c[207]) );
  DFF \creg_reg[208]  ( .D(creg_next[208]), .CLK(clk), .RST(rst), .I(m[208]), 
        .Q(c[208]) );
  DFF \creg_reg[209]  ( .D(creg_next[209]), .CLK(clk), .RST(rst), .I(m[209]), 
        .Q(c[209]) );
  DFF \creg_reg[210]  ( .D(creg_next[210]), .CLK(clk), .RST(rst), .I(m[210]), 
        .Q(c[210]) );
  DFF \creg_reg[211]  ( .D(creg_next[211]), .CLK(clk), .RST(rst), .I(m[211]), 
        .Q(c[211]) );
  DFF \creg_reg[212]  ( .D(creg_next[212]), .CLK(clk), .RST(rst), .I(m[212]), 
        .Q(c[212]) );
  DFF \creg_reg[213]  ( .D(creg_next[213]), .CLK(clk), .RST(rst), .I(m[213]), 
        .Q(c[213]) );
  DFF \creg_reg[214]  ( .D(creg_next[214]), .CLK(clk), .RST(rst), .I(m[214]), 
        .Q(c[214]) );
  DFF \creg_reg[215]  ( .D(creg_next[215]), .CLK(clk), .RST(rst), .I(m[215]), 
        .Q(c[215]) );
  DFF \creg_reg[216]  ( .D(creg_next[216]), .CLK(clk), .RST(rst), .I(m[216]), 
        .Q(c[216]) );
  DFF \creg_reg[217]  ( .D(creg_next[217]), .CLK(clk), .RST(rst), .I(m[217]), 
        .Q(c[217]) );
  DFF \creg_reg[218]  ( .D(creg_next[218]), .CLK(clk), .RST(rst), .I(m[218]), 
        .Q(c[218]) );
  DFF \creg_reg[219]  ( .D(creg_next[219]), .CLK(clk), .RST(rst), .I(m[219]), 
        .Q(c[219]) );
  DFF \creg_reg[220]  ( .D(creg_next[220]), .CLK(clk), .RST(rst), .I(m[220]), 
        .Q(c[220]) );
  DFF \creg_reg[221]  ( .D(creg_next[221]), .CLK(clk), .RST(rst), .I(m[221]), 
        .Q(c[221]) );
  DFF \creg_reg[222]  ( .D(creg_next[222]), .CLK(clk), .RST(rst), .I(m[222]), 
        .Q(c[222]) );
  DFF \creg_reg[223]  ( .D(creg_next[223]), .CLK(clk), .RST(rst), .I(m[223]), 
        .Q(c[223]) );
  DFF \creg_reg[224]  ( .D(creg_next[224]), .CLK(clk), .RST(rst), .I(m[224]), 
        .Q(c[224]) );
  DFF \creg_reg[225]  ( .D(creg_next[225]), .CLK(clk), .RST(rst), .I(m[225]), 
        .Q(c[225]) );
  DFF \creg_reg[226]  ( .D(creg_next[226]), .CLK(clk), .RST(rst), .I(m[226]), 
        .Q(c[226]) );
  DFF \creg_reg[227]  ( .D(creg_next[227]), .CLK(clk), .RST(rst), .I(m[227]), 
        .Q(c[227]) );
  DFF \creg_reg[228]  ( .D(creg_next[228]), .CLK(clk), .RST(rst), .I(m[228]), 
        .Q(c[228]) );
  DFF \creg_reg[229]  ( .D(creg_next[229]), .CLK(clk), .RST(rst), .I(m[229]), 
        .Q(c[229]) );
  DFF \creg_reg[230]  ( .D(creg_next[230]), .CLK(clk), .RST(rst), .I(m[230]), 
        .Q(c[230]) );
  DFF \creg_reg[231]  ( .D(creg_next[231]), .CLK(clk), .RST(rst), .I(m[231]), 
        .Q(c[231]) );
  DFF \creg_reg[232]  ( .D(creg_next[232]), .CLK(clk), .RST(rst), .I(m[232]), 
        .Q(c[232]) );
  DFF \creg_reg[233]  ( .D(creg_next[233]), .CLK(clk), .RST(rst), .I(m[233]), 
        .Q(c[233]) );
  DFF \creg_reg[234]  ( .D(creg_next[234]), .CLK(clk), .RST(rst), .I(m[234]), 
        .Q(c[234]) );
  DFF \creg_reg[235]  ( .D(creg_next[235]), .CLK(clk), .RST(rst), .I(m[235]), 
        .Q(c[235]) );
  DFF \creg_reg[236]  ( .D(creg_next[236]), .CLK(clk), .RST(rst), .I(m[236]), 
        .Q(c[236]) );
  DFF \creg_reg[237]  ( .D(creg_next[237]), .CLK(clk), .RST(rst), .I(m[237]), 
        .Q(c[237]) );
  DFF \creg_reg[238]  ( .D(creg_next[238]), .CLK(clk), .RST(rst), .I(m[238]), 
        .Q(c[238]) );
  DFF \creg_reg[239]  ( .D(creg_next[239]), .CLK(clk), .RST(rst), .I(m[239]), 
        .Q(c[239]) );
  DFF \creg_reg[240]  ( .D(creg_next[240]), .CLK(clk), .RST(rst), .I(m[240]), 
        .Q(c[240]) );
  DFF \creg_reg[241]  ( .D(creg_next[241]), .CLK(clk), .RST(rst), .I(m[241]), 
        .Q(c[241]) );
  DFF \creg_reg[242]  ( .D(creg_next[242]), .CLK(clk), .RST(rst), .I(m[242]), 
        .Q(c[242]) );
  DFF \creg_reg[243]  ( .D(creg_next[243]), .CLK(clk), .RST(rst), .I(m[243]), 
        .Q(c[243]) );
  DFF \creg_reg[244]  ( .D(creg_next[244]), .CLK(clk), .RST(rst), .I(m[244]), 
        .Q(c[244]) );
  DFF \creg_reg[245]  ( .D(creg_next[245]), .CLK(clk), .RST(rst), .I(m[245]), 
        .Q(c[245]) );
  DFF \creg_reg[246]  ( .D(creg_next[246]), .CLK(clk), .RST(rst), .I(m[246]), 
        .Q(c[246]) );
  DFF \creg_reg[247]  ( .D(creg_next[247]), .CLK(clk), .RST(rst), .I(m[247]), 
        .Q(c[247]) );
  DFF \creg_reg[248]  ( .D(creg_next[248]), .CLK(clk), .RST(rst), .I(m[248]), 
        .Q(c[248]) );
  DFF \creg_reg[249]  ( .D(creg_next[249]), .CLK(clk), .RST(rst), .I(m[249]), 
        .Q(c[249]) );
  DFF \creg_reg[250]  ( .D(creg_next[250]), .CLK(clk), .RST(rst), .I(m[250]), 
        .Q(c[250]) );
  DFF \creg_reg[251]  ( .D(creg_next[251]), .CLK(clk), .RST(rst), .I(m[251]), 
        .Q(c[251]) );
  DFF \creg_reg[252]  ( .D(creg_next[252]), .CLK(clk), .RST(rst), .I(m[252]), 
        .Q(c[252]) );
  DFF \creg_reg[253]  ( .D(creg_next[253]), .CLK(clk), .RST(rst), .I(m[253]), 
        .Q(c[253]) );
  DFF \creg_reg[254]  ( .D(creg_next[254]), .CLK(clk), .RST(rst), .I(m[254]), 
        .Q(c[254]) );
  DFF \creg_reg[255]  ( .D(creg_next[255]), .CLK(clk), .RST(rst), .I(m[255]), 
        .Q(c[255]) );
  XOR U140 ( .A(start_in[127]), .B(mul_pow), .Z(n8) );
  NANDN U141 ( .A(first_one), .B(n137), .Z(n6) );
  NAND U142 ( .A(n138), .B(ein[255]), .Z(n137) );
  AND U143 ( .A(mul_pow), .B(start_in[127]), .Z(n138) );
  NAND U144 ( .A(n139), .B(n140), .Z(_0_net_) );
  NANDN U145 ( .A(mul_pow), .B(first_one), .Z(n140) );
  NAND U146 ( .A(first_one), .B(ein[255]), .Z(n139) );
endmodule

