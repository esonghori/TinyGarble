
module round_2 ( in, round_const, out );
  input [1599:0] in;
  input [63:0] round_const;
  output [1599:0] out;
  wire   round_const_63, round_const_31, round_const_15, round_const_7,
         round_const_3, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
         n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
         n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
         n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
         n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
         n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
         n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
         n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
         n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
         n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
         n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
         n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
         n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807;
  assign round_const_63 = round_const[63];
  assign round_const_31 = round_const[31];
  assign round_const_15 = round_const[15];
  assign round_const_7 = round_const[7];
  assign round_const_3 = round_const[3];

  XOR U1 ( .A(in[1469]), .B(in[509]), .Z(n2) );
  XNOR U2 ( .A(in[829]), .B(in[189]), .Z(n1) );
  XNOR U3 ( .A(n2), .B(n1), .Z(n3) );
  XOR U4 ( .A(in[1149]), .B(n3), .Z(n872) );
  XOR U5 ( .A(in[1598]), .B(in[638]), .Z(n5) );
  XNOR U6 ( .A(in[958]), .B(in[318]), .Z(n4) );
  XNOR U7 ( .A(n5), .B(n4), .Z(n6) );
  XOR U8 ( .A(in[1278]), .B(n6), .Z(n1473) );
  XNOR U9 ( .A(n872), .B(n1473), .Z(n3815) );
  XNOR U10 ( .A(in[254]), .B(n3815), .Z(n3577) );
  XOR U11 ( .A(in[1345]), .B(in[65]), .Z(n8) );
  XNOR U12 ( .A(in[1025]), .B(in[385]), .Z(n7) );
  XNOR U13 ( .A(n8), .B(n7), .Z(n9) );
  XOR U14 ( .A(in[705]), .B(n9), .Z(n1481) );
  XOR U15 ( .A(in[1474]), .B(in[514]), .Z(n11) );
  XNOR U16 ( .A(in[834]), .B(in[194]), .Z(n10) );
  XNOR U17 ( .A(n11), .B(n10), .Z(n12) );
  XNOR U18 ( .A(in[1154]), .B(n12), .Z(n1188) );
  XNOR U19 ( .A(n1481), .B(n1188), .Z(n3570) );
  XNOR U20 ( .A(in[1410]), .B(n3570), .Z(n3576) );
  XOR U21 ( .A(in[328]), .B(in[8]), .Z(n14) );
  XNOR U22 ( .A(in[968]), .B(in[648]), .Z(n13) );
  XNOR U23 ( .A(n14), .B(n13), .Z(n15) );
  XOR U24 ( .A(in[1288]), .B(n15), .Z(n1209) );
  XOR U25 ( .A(in[137]), .B(in[457]), .Z(n17) );
  XNOR U26 ( .A(in[777]), .B(in[1417]), .Z(n16) );
  XNOR U27 ( .A(n17), .B(n16), .Z(n18) );
  XOR U28 ( .A(in[1097]), .B(n18), .Z(n1141) );
  XNOR U29 ( .A(n1209), .B(n1141), .Z(n4086) );
  XNOR U30 ( .A(in[1033]), .B(n4086), .Z(n2609) );
  NAND U31 ( .A(n3576), .B(n2609), .Z(n19) );
  XNOR U32 ( .A(n3577), .B(n19), .Z(out[0]) );
  XOR U33 ( .A(in[1515]), .B(in[555]), .Z(n21) );
  XNOR U34 ( .A(in[875]), .B(in[235]), .Z(n20) );
  XNOR U35 ( .A(n21), .B(n20), .Z(n22) );
  XOR U36 ( .A(in[1195]), .B(n22), .Z(n1329) );
  XOR U37 ( .A(in[1386]), .B(in[106]), .Z(n24) );
  XNOR U38 ( .A(in[1066]), .B(in[746]), .Z(n23) );
  XNOR U39 ( .A(n24), .B(n23), .Z(n25) );
  XOR U40 ( .A(in[426]), .B(n25), .Z(n475) );
  XNOR U41 ( .A(n1329), .B(n475), .Z(n3750) );
  XNOR U42 ( .A(in[171]), .B(n3750), .Z(n1301) );
  XOR U43 ( .A(in[140]), .B(in[460]), .Z(n27) );
  XNOR U44 ( .A(in[1100]), .B(in[1420]), .Z(n26) );
  XNOR U45 ( .A(n27), .B(n26), .Z(n28) );
  XOR U46 ( .A(in[780]), .B(n28), .Z(n1159) );
  XOR U47 ( .A(in[971]), .B(in[1291]), .Z(n30) );
  XNOR U48 ( .A(in[11]), .B(in[331]), .Z(n29) );
  XNOR U49 ( .A(n30), .B(n29), .Z(n31) );
  XNOR U50 ( .A(in[651]), .B(n31), .Z(n1220) );
  XNOR U51 ( .A(n1159), .B(n1220), .Z(n4095) );
  XNOR U52 ( .A(in[1356]), .B(n4095), .Z(n1696) );
  XOR U53 ( .A(in[1364]), .B(in[724]), .Z(n33) );
  XNOR U54 ( .A(in[84]), .B(in[404]), .Z(n32) );
  XNOR U55 ( .A(n33), .B(n32), .Z(n34) );
  XOR U56 ( .A(in[1044]), .B(n34), .Z(n777) );
  XOR U57 ( .A(in[1555]), .B(in[595]), .Z(n36) );
  XNOR U58 ( .A(in[915]), .B(in[275]), .Z(n35) );
  XNOR U59 ( .A(n36), .B(n35), .Z(n37) );
  XOR U60 ( .A(in[1235]), .B(n37), .Z(n489) );
  XNOR U61 ( .A(n777), .B(n489), .Z(n3882) );
  XNOR U62 ( .A(in[980]), .B(n3882), .Z(n1693) );
  NAND U63 ( .A(n1696), .B(n1693), .Z(n38) );
  XNOR U64 ( .A(n1301), .B(n38), .Z(out[1000]) );
  XOR U65 ( .A(in[1516]), .B(in[556]), .Z(n40) );
  XNOR U66 ( .A(in[876]), .B(in[236]), .Z(n39) );
  XNOR U67 ( .A(n40), .B(n39), .Z(n41) );
  XOR U68 ( .A(in[1196]), .B(n41), .Z(n1333) );
  XOR U69 ( .A(in[1387]), .B(in[107]), .Z(n43) );
  XNOR U70 ( .A(in[1067]), .B(in[747]), .Z(n42) );
  XNOR U71 ( .A(n43), .B(n42), .Z(n44) );
  XOR U72 ( .A(in[427]), .B(n44), .Z(n486) );
  XNOR U73 ( .A(n1333), .B(n486), .Z(n3758) );
  XNOR U74 ( .A(in[172]), .B(n3758), .Z(n1305) );
  XOR U75 ( .A(in[972]), .B(in[12]), .Z(n46) );
  XNOR U76 ( .A(in[1292]), .B(in[332]), .Z(n45) );
  XNOR U77 ( .A(n46), .B(n45), .Z(n47) );
  XOR U78 ( .A(in[652]), .B(n47), .Z(n1223) );
  XOR U79 ( .A(in[141]), .B(in[461]), .Z(n49) );
  XNOR U80 ( .A(in[1101]), .B(in[1421]), .Z(n48) );
  XNOR U81 ( .A(n49), .B(n48), .Z(n50) );
  XNOR U82 ( .A(in[781]), .B(n50), .Z(n1164) );
  XNOR U83 ( .A(n1223), .B(n1164), .Z(n4098) );
  XNOR U84 ( .A(in[1357]), .B(n4098), .Z(n1700) );
  XOR U85 ( .A(in[1365]), .B(in[725]), .Z(n52) );
  XNOR U86 ( .A(in[85]), .B(in[405]), .Z(n51) );
  XNOR U87 ( .A(n52), .B(n51), .Z(n53) );
  XOR U88 ( .A(in[1045]), .B(n53), .Z(n790) );
  XOR U89 ( .A(in[1556]), .B(in[596]), .Z(n55) );
  XNOR U90 ( .A(in[916]), .B(in[276]), .Z(n54) );
  XNOR U91 ( .A(n55), .B(n54), .Z(n56) );
  XOR U92 ( .A(in[1236]), .B(n56), .Z(n504) );
  XNOR U93 ( .A(n790), .B(n504), .Z(n3884) );
  XNOR U94 ( .A(in[981]), .B(n3884), .Z(n1697) );
  NAND U95 ( .A(n1700), .B(n1697), .Z(n57) );
  XNOR U96 ( .A(n1305), .B(n57), .Z(out[1001]) );
  XOR U97 ( .A(in[1388]), .B(in[108]), .Z(n59) );
  XNOR U98 ( .A(in[1068]), .B(in[748]), .Z(n58) );
  XNOR U99 ( .A(n59), .B(n58), .Z(n60) );
  XOR U100 ( .A(in[428]), .B(n60), .Z(n1395) );
  XOR U101 ( .A(in[1517]), .B(in[557]), .Z(n62) );
  XNOR U102 ( .A(in[877]), .B(in[237]), .Z(n61) );
  XNOR U103 ( .A(n62), .B(n61), .Z(n63) );
  XOR U104 ( .A(in[1197]), .B(n63), .Z(n1337) );
  XNOR U105 ( .A(n1395), .B(n1337), .Z(n3762) );
  XNOR U106 ( .A(in[173]), .B(n3762), .Z(n1310) );
  XOR U107 ( .A(in[973]), .B(in[13]), .Z(n65) );
  XNOR U108 ( .A(in[1293]), .B(in[333]), .Z(n64) );
  XNOR U109 ( .A(n65), .B(n64), .Z(n66) );
  XOR U110 ( .A(in[653]), .B(n66), .Z(n1226) );
  XOR U111 ( .A(in[142]), .B(in[1422]), .Z(n68) );
  XNOR U112 ( .A(in[1102]), .B(in[782]), .Z(n67) );
  XNOR U113 ( .A(n68), .B(n67), .Z(n69) );
  XNOR U114 ( .A(in[462]), .B(n69), .Z(n1169) );
  XNOR U115 ( .A(n1226), .B(n1169), .Z(n4101) );
  XNOR U116 ( .A(in[1358]), .B(n4101), .Z(n1704) );
  XOR U117 ( .A(in[1366]), .B(in[726]), .Z(n71) );
  XNOR U118 ( .A(in[86]), .B(in[406]), .Z(n70) );
  XNOR U119 ( .A(n71), .B(n70), .Z(n72) );
  XOR U120 ( .A(in[1046]), .B(n72), .Z(n803) );
  XOR U121 ( .A(in[1557]), .B(in[597]), .Z(n74) );
  XNOR U122 ( .A(in[917]), .B(in[277]), .Z(n73) );
  XNOR U123 ( .A(n74), .B(n73), .Z(n75) );
  XOR U124 ( .A(in[1237]), .B(n75), .Z(n519) );
  XNOR U125 ( .A(n803), .B(n519), .Z(n3886) );
  XNOR U126 ( .A(in[982]), .B(n3886), .Z(n1701) );
  NAND U127 ( .A(n1704), .B(n1701), .Z(n76) );
  XNOR U128 ( .A(n1310), .B(n76), .Z(out[1002]) );
  XOR U129 ( .A(in[1389]), .B(in[109]), .Z(n78) );
  XNOR U130 ( .A(in[1069]), .B(in[749]), .Z(n77) );
  XNOR U131 ( .A(n78), .B(n77), .Z(n79) );
  XOR U132 ( .A(in[429]), .B(n79), .Z(n1399) );
  XOR U133 ( .A(in[1518]), .B(in[558]), .Z(n81) );
  XNOR U134 ( .A(in[878]), .B(in[238]), .Z(n80) );
  XNOR U135 ( .A(n81), .B(n80), .Z(n82) );
  XOR U136 ( .A(in[1198]), .B(n82), .Z(n1341) );
  XNOR U137 ( .A(n1399), .B(n1341), .Z(n3766) );
  XNOR U138 ( .A(in[174]), .B(n3766), .Z(n1314) );
  XOR U139 ( .A(in[143]), .B(in[1423]), .Z(n84) );
  XNOR U140 ( .A(in[1103]), .B(in[783]), .Z(n83) );
  XNOR U141 ( .A(n84), .B(n83), .Z(n85) );
  XOR U142 ( .A(in[463]), .B(n85), .Z(n1174) );
  XOR U143 ( .A(in[974]), .B(in[14]), .Z(n87) );
  XNOR U144 ( .A(in[1294]), .B(in[334]), .Z(n86) );
  XNOR U145 ( .A(n87), .B(n86), .Z(n88) );
  XNOR U146 ( .A(in[654]), .B(n88), .Z(n1229) );
  XNOR U147 ( .A(n1174), .B(n1229), .Z(n4104) );
  XNOR U148 ( .A(in[1359]), .B(n4104), .Z(n1708) );
  XOR U149 ( .A(in[1367]), .B(in[727]), .Z(n90) );
  XNOR U150 ( .A(in[87]), .B(in[407]), .Z(n89) );
  XNOR U151 ( .A(n90), .B(n89), .Z(n91) );
  XOR U152 ( .A(in[1047]), .B(n91), .Z(n816) );
  XOR U153 ( .A(in[1558]), .B(in[598]), .Z(n93) );
  XNOR U154 ( .A(in[918]), .B(in[278]), .Z(n92) );
  XNOR U155 ( .A(n93), .B(n92), .Z(n94) );
  XOR U156 ( .A(in[1238]), .B(n94), .Z(n534) );
  XNOR U157 ( .A(n816), .B(n534), .Z(n3888) );
  XNOR U158 ( .A(in[983]), .B(n3888), .Z(n1705) );
  NAND U159 ( .A(n1708), .B(n1705), .Z(n95) );
  XNOR U160 ( .A(n1314), .B(n95), .Z(out[1003]) );
  XOR U161 ( .A(in[1390]), .B(in[110]), .Z(n97) );
  XNOR U162 ( .A(in[1070]), .B(in[750]), .Z(n96) );
  XNOR U163 ( .A(n97), .B(n96), .Z(n98) );
  XOR U164 ( .A(in[430]), .B(n98), .Z(n1403) );
  XOR U165 ( .A(in[1519]), .B(in[559]), .Z(n100) );
  XNOR U166 ( .A(in[879]), .B(in[239]), .Z(n99) );
  XNOR U167 ( .A(n100), .B(n99), .Z(n101) );
  XOR U168 ( .A(in[1199]), .B(n101), .Z(n1345) );
  XNOR U169 ( .A(n1403), .B(n1345), .Z(n3770) );
  XNOR U170 ( .A(in[175]), .B(n3770), .Z(n1318) );
  XOR U171 ( .A(in[144]), .B(in[1424]), .Z(n103) );
  XNOR U172 ( .A(in[1104]), .B(in[784]), .Z(n102) );
  XNOR U173 ( .A(n103), .B(n102), .Z(n104) );
  XOR U174 ( .A(in[464]), .B(n104), .Z(n1179) );
  XOR U175 ( .A(in[975]), .B(in[15]), .Z(n106) );
  XNOR U176 ( .A(in[1295]), .B(in[335]), .Z(n105) );
  XNOR U177 ( .A(n106), .B(n105), .Z(n107) );
  XNOR U178 ( .A(in[655]), .B(n107), .Z(n1232) );
  XNOR U179 ( .A(n1179), .B(n1232), .Z(n4107) );
  XNOR U180 ( .A(in[1360]), .B(n4107), .Z(n1713) );
  XOR U181 ( .A(in[1368]), .B(in[728]), .Z(n109) );
  XNOR U182 ( .A(in[88]), .B(in[408]), .Z(n108) );
  XNOR U183 ( .A(n109), .B(n108), .Z(n110) );
  XOR U184 ( .A(in[1048]), .B(n110), .Z(n829) );
  XOR U185 ( .A(in[1559]), .B(in[599]), .Z(n112) );
  XNOR U186 ( .A(in[919]), .B(in[279]), .Z(n111) );
  XNOR U187 ( .A(n112), .B(n111), .Z(n113) );
  XOR U188 ( .A(in[1239]), .B(n113), .Z(n549) );
  XNOR U189 ( .A(n829), .B(n549), .Z(n3890) );
  XNOR U190 ( .A(in[984]), .B(n3890), .Z(n1710) );
  NAND U191 ( .A(n1713), .B(n1710), .Z(n114) );
  XNOR U192 ( .A(n1318), .B(n114), .Z(out[1004]) );
  XOR U193 ( .A(in[1391]), .B(in[111]), .Z(n116) );
  XNOR U194 ( .A(in[1071]), .B(in[751]), .Z(n115) );
  XNOR U195 ( .A(n116), .B(n115), .Z(n117) );
  XOR U196 ( .A(in[431]), .B(n117), .Z(n1407) );
  XOR U197 ( .A(in[1520]), .B(in[560]), .Z(n119) );
  XNOR U198 ( .A(in[880]), .B(in[240]), .Z(n118) );
  XNOR U199 ( .A(n119), .B(n118), .Z(n120) );
  XOR U200 ( .A(in[1200]), .B(n120), .Z(n1350) );
  XNOR U201 ( .A(n1407), .B(n1350), .Z(n3774) );
  XNOR U202 ( .A(in[176]), .B(n3774), .Z(n1322) );
  XOR U203 ( .A(in[976]), .B(in[16]), .Z(n122) );
  XNOR U204 ( .A(in[1296]), .B(in[336]), .Z(n121) );
  XNOR U205 ( .A(n122), .B(n121), .Z(n123) );
  XOR U206 ( .A(in[656]), .B(n123), .Z(n1235) );
  XOR U207 ( .A(in[145]), .B(in[1425]), .Z(n125) );
  XNOR U208 ( .A(in[1105]), .B(in[785]), .Z(n124) );
  XNOR U209 ( .A(n125), .B(n124), .Z(n126) );
  XNOR U210 ( .A(in[465]), .B(n126), .Z(n1184) );
  XNOR U211 ( .A(n1235), .B(n1184), .Z(n4114) );
  XNOR U212 ( .A(in[1361]), .B(n4114), .Z(n1717) );
  XOR U213 ( .A(in[1369]), .B(in[729]), .Z(n128) );
  XNOR U214 ( .A(in[89]), .B(in[409]), .Z(n127) );
  XNOR U215 ( .A(n128), .B(n127), .Z(n129) );
  XOR U216 ( .A(in[1049]), .B(n129), .Z(n842) );
  XOR U217 ( .A(in[1560]), .B(in[600]), .Z(n131) );
  XNOR U218 ( .A(in[920]), .B(in[280]), .Z(n130) );
  XNOR U219 ( .A(n131), .B(n130), .Z(n132) );
  XOR U220 ( .A(in[1240]), .B(n132), .Z(n564) );
  XNOR U221 ( .A(n842), .B(n564), .Z(n3892) );
  XNOR U222 ( .A(in[985]), .B(n3892), .Z(n1714) );
  NAND U223 ( .A(n1717), .B(n1714), .Z(n133) );
  XNOR U224 ( .A(n1322), .B(n133), .Z(out[1005]) );
  XOR U225 ( .A(in[1392]), .B(in[112]), .Z(n135) );
  XNOR U226 ( .A(in[1072]), .B(in[752]), .Z(n134) );
  XNOR U227 ( .A(n135), .B(n134), .Z(n136) );
  XOR U228 ( .A(in[432]), .B(n136), .Z(n1411) );
  XOR U229 ( .A(in[1521]), .B(in[561]), .Z(n138) );
  XNOR U230 ( .A(in[881]), .B(in[241]), .Z(n137) );
  XNOR U231 ( .A(n138), .B(n137), .Z(n139) );
  XOR U232 ( .A(in[1201]), .B(n139), .Z(n1354) );
  XNOR U233 ( .A(n1411), .B(n1354), .Z(n3778) );
  XNOR U234 ( .A(in[177]), .B(n3778), .Z(n1326) );
  XOR U235 ( .A(in[1426]), .B(in[466]), .Z(n141) );
  XNOR U236 ( .A(in[786]), .B(in[146]), .Z(n140) );
  XNOR U237 ( .A(n141), .B(n140), .Z(n142) );
  XOR U238 ( .A(in[1106]), .B(n142), .Z(n488) );
  XOR U239 ( .A(in[17]), .B(in[657]), .Z(n144) );
  XNOR U240 ( .A(in[977]), .B(in[337]), .Z(n143) );
  XNOR U241 ( .A(n144), .B(n143), .Z(n145) );
  XNOR U242 ( .A(in[1297]), .B(n145), .Z(n1238) );
  XNOR U243 ( .A(n488), .B(n1238), .Z(n4117) );
  XNOR U244 ( .A(n4117), .B(in[1362]), .Z(n1721) );
  XOR U245 ( .A(in[1370]), .B(in[730]), .Z(n147) );
  XNOR U246 ( .A(in[90]), .B(in[410]), .Z(n146) );
  XNOR U247 ( .A(n147), .B(n146), .Z(n148) );
  XOR U248 ( .A(in[1050]), .B(n148), .Z(n857) );
  XOR U249 ( .A(in[1561]), .B(in[601]), .Z(n150) );
  XNOR U250 ( .A(in[921]), .B(in[281]), .Z(n149) );
  XNOR U251 ( .A(n150), .B(n149), .Z(n151) );
  XOR U252 ( .A(in[1241]), .B(n151), .Z(n590) );
  XNOR U253 ( .A(n857), .B(n590), .Z(n3894) );
  XNOR U254 ( .A(in[986]), .B(n3894), .Z(n1718) );
  NAND U255 ( .A(n1721), .B(n1718), .Z(n152) );
  XNOR U256 ( .A(n1326), .B(n152), .Z(out[1006]) );
  XOR U257 ( .A(in[1393]), .B(in[113]), .Z(n154) );
  XNOR U258 ( .A(in[1073]), .B(in[753]), .Z(n153) );
  XNOR U259 ( .A(n154), .B(n153), .Z(n155) );
  XOR U260 ( .A(in[433]), .B(n155), .Z(n1415) );
  XOR U261 ( .A(in[1522]), .B(in[562]), .Z(n157) );
  XNOR U262 ( .A(in[882]), .B(in[242]), .Z(n156) );
  XNOR U263 ( .A(n157), .B(n156), .Z(n158) );
  XOR U264 ( .A(in[1202]), .B(n158), .Z(n1358) );
  XNOR U265 ( .A(n1415), .B(n1358), .Z(n3782) );
  XNOR U266 ( .A(in[178]), .B(n3782), .Z(n1330) );
  XOR U267 ( .A(in[978]), .B(in[18]), .Z(n160) );
  XNOR U268 ( .A(in[1298]), .B(in[338]), .Z(n159) );
  XNOR U269 ( .A(n160), .B(n159), .Z(n161) );
  XOR U270 ( .A(in[658]), .B(n161), .Z(n1241) );
  XOR U271 ( .A(in[147]), .B(in[1427]), .Z(n163) );
  XNOR U272 ( .A(in[1107]), .B(in[787]), .Z(n162) );
  XNOR U273 ( .A(n163), .B(n162), .Z(n164) );
  XNOR U274 ( .A(in[467]), .B(n164), .Z(n503) );
  XNOR U275 ( .A(n1241), .B(n503), .Z(n4120) );
  XNOR U276 ( .A(in[1363]), .B(n4120), .Z(n1725) );
  XOR U277 ( .A(in[1371]), .B(in[731]), .Z(n166) );
  XNOR U278 ( .A(in[91]), .B(in[411]), .Z(n165) );
  XNOR U279 ( .A(n166), .B(n165), .Z(n167) );
  XOR U280 ( .A(in[1051]), .B(n167), .Z(n870) );
  XOR U281 ( .A(in[1562]), .B(in[602]), .Z(n169) );
  XNOR U282 ( .A(in[922]), .B(in[282]), .Z(n168) );
  XNOR U283 ( .A(n169), .B(n168), .Z(n170) );
  XOR U284 ( .A(in[1242]), .B(n170), .Z(n605) );
  XNOR U285 ( .A(n870), .B(n605), .Z(n3896) );
  XNOR U286 ( .A(in[987]), .B(n3896), .Z(n1722) );
  NAND U287 ( .A(n1725), .B(n1722), .Z(n171) );
  XNOR U288 ( .A(n1330), .B(n171), .Z(out[1007]) );
  XOR U289 ( .A(in[1394]), .B(in[114]), .Z(n173) );
  XNOR U290 ( .A(in[1074]), .B(in[754]), .Z(n172) );
  XNOR U291 ( .A(n173), .B(n172), .Z(n174) );
  XOR U292 ( .A(in[434]), .B(n174), .Z(n1419) );
  XOR U293 ( .A(in[1523]), .B(in[563]), .Z(n176) );
  XNOR U294 ( .A(in[883]), .B(in[243]), .Z(n175) );
  XNOR U295 ( .A(n176), .B(n175), .Z(n177) );
  XOR U296 ( .A(in[1203]), .B(n177), .Z(n1362) );
  XNOR U297 ( .A(n1419), .B(n1362), .Z(n3786) );
  XNOR U298 ( .A(in[179]), .B(n3786), .Z(n1334) );
  XOR U299 ( .A(in[148]), .B(in[1428]), .Z(n179) );
  XNOR U300 ( .A(in[1108]), .B(in[788]), .Z(n178) );
  XNOR U301 ( .A(n179), .B(n178), .Z(n180) );
  XOR U302 ( .A(in[468]), .B(n180), .Z(n518) );
  XOR U303 ( .A(in[979]), .B(in[19]), .Z(n182) );
  XNOR U304 ( .A(in[1299]), .B(in[339]), .Z(n181) );
  XNOR U305 ( .A(n182), .B(n181), .Z(n183) );
  XNOR U306 ( .A(in[659]), .B(n183), .Z(n1245) );
  XNOR U307 ( .A(n518), .B(n1245), .Z(n4123) );
  XNOR U308 ( .A(in[1364]), .B(n4123), .Z(n1729) );
  XOR U309 ( .A(in[1372]), .B(in[732]), .Z(n185) );
  XNOR U310 ( .A(in[92]), .B(in[412]), .Z(n184) );
  XNOR U311 ( .A(n185), .B(n184), .Z(n186) );
  XOR U312 ( .A(in[1052]), .B(n186), .Z(n890) );
  XOR U313 ( .A(in[1563]), .B(in[603]), .Z(n188) );
  XNOR U314 ( .A(in[923]), .B(in[283]), .Z(n187) );
  XNOR U315 ( .A(n188), .B(n187), .Z(n189) );
  XOR U316 ( .A(in[1243]), .B(n189), .Z(n620) );
  XNOR U317 ( .A(n890), .B(n620), .Z(n3900) );
  XNOR U318 ( .A(in[988]), .B(n3900), .Z(n1726) );
  NAND U319 ( .A(n1729), .B(n1726), .Z(n190) );
  XNOR U320 ( .A(n1334), .B(n190), .Z(out[1008]) );
  XOR U321 ( .A(in[1395]), .B(in[115]), .Z(n192) );
  XNOR U322 ( .A(in[1075]), .B(in[755]), .Z(n191) );
  XNOR U323 ( .A(n192), .B(n191), .Z(n193) );
  XOR U324 ( .A(in[435]), .B(n193), .Z(n1423) );
  XOR U325 ( .A(in[1524]), .B(in[564]), .Z(n195) );
  XNOR U326 ( .A(in[884]), .B(in[244]), .Z(n194) );
  XNOR U327 ( .A(n195), .B(n194), .Z(n196) );
  XOR U328 ( .A(in[1204]), .B(n196), .Z(n1366) );
  XNOR U329 ( .A(n1423), .B(n1366), .Z(n3790) );
  XNOR U330 ( .A(in[180]), .B(n3790), .Z(n1338) );
  XOR U331 ( .A(in[340]), .B(in[660]), .Z(n198) );
  XNOR U332 ( .A(in[20]), .B(in[1300]), .Z(n197) );
  XNOR U333 ( .A(n198), .B(n197), .Z(n199) );
  XOR U334 ( .A(in[980]), .B(n199), .Z(n1248) );
  XOR U335 ( .A(in[149]), .B(in[1429]), .Z(n201) );
  XNOR U336 ( .A(in[1109]), .B(in[789]), .Z(n200) );
  XNOR U337 ( .A(n201), .B(n200), .Z(n202) );
  XNOR U338 ( .A(in[469]), .B(n202), .Z(n533) );
  XNOR U339 ( .A(n1248), .B(n533), .Z(n4126) );
  XNOR U340 ( .A(in[1365]), .B(n4126), .Z(n1733) );
  XOR U341 ( .A(in[1373]), .B(in[733]), .Z(n204) );
  XNOR U342 ( .A(in[93]), .B(in[413]), .Z(n203) );
  XNOR U343 ( .A(n204), .B(n203), .Z(n205) );
  XOR U344 ( .A(in[1053]), .B(n205), .Z(n903) );
  XOR U345 ( .A(in[1564]), .B(in[604]), .Z(n207) );
  XNOR U346 ( .A(in[924]), .B(in[284]), .Z(n206) );
  XNOR U347 ( .A(n207), .B(n206), .Z(n208) );
  XOR U348 ( .A(in[1244]), .B(n208), .Z(n635) );
  XNOR U349 ( .A(n903), .B(n635), .Z(n3902) );
  XNOR U350 ( .A(in[989]), .B(n3902), .Z(n1730) );
  NAND U351 ( .A(n1733), .B(n1730), .Z(n209) );
  XNOR U352 ( .A(n1338), .B(n209), .Z(out[1009]) );
  XOR U353 ( .A(in[1339]), .B(in[59]), .Z(n211) );
  XNOR U354 ( .A(in[699]), .B(in[379]), .Z(n210) );
  XNOR U355 ( .A(n211), .B(n210), .Z(n212) );
  XOR U356 ( .A(in[1019]), .B(n212), .Z(n861) );
  XOR U357 ( .A(in[1530]), .B(in[570]), .Z(n214) );
  XNOR U358 ( .A(in[1210]), .B(in[250]), .Z(n213) );
  XNOR U359 ( .A(n214), .B(n213), .Z(n215) );
  XOR U360 ( .A(in[890]), .B(n215), .Z(n327) );
  XNOR U361 ( .A(n861), .B(n327), .Z(n3592) );
  XNOR U362 ( .A(in[635]), .B(n3592), .Z(n2550) );
  XOR U363 ( .A(in[161]), .B(in[1441]), .Z(n217) );
  XNOR U364 ( .A(in[801]), .B(in[1121]), .Z(n216) );
  XNOR U365 ( .A(n217), .B(n216), .Z(n218) );
  XOR U366 ( .A(in[481]), .B(n218), .Z(n454) );
  XOR U367 ( .A(in[1570]), .B(in[610]), .Z(n220) );
  XNOR U368 ( .A(in[930]), .B(in[290]), .Z(n219) );
  XNOR U369 ( .A(n220), .B(n219), .Z(n221) );
  XNOR U370 ( .A(in[1250]), .B(n221), .Z(n337) );
  XNOR U371 ( .A(n454), .B(n337), .Z(n3689) );
  XNOR U372 ( .A(in[226]), .B(n3689), .Z(n2831) );
  XOR U373 ( .A(in[1510]), .B(in[550]), .Z(n223) );
  XNOR U374 ( .A(in[870]), .B(in[230]), .Z(n222) );
  XNOR U375 ( .A(n223), .B(n222), .Z(n224) );
  XOR U376 ( .A(in[1190]), .B(n224), .Z(n1309) );
  XOR U377 ( .A(in[1061]), .B(in[421]), .Z(n226) );
  XNOR U378 ( .A(in[741]), .B(in[1381]), .Z(n225) );
  XNOR U379 ( .A(n226), .B(n225), .Z(n227) );
  XOR U380 ( .A(in[101]), .B(n227), .Z(n373) );
  XNOR U381 ( .A(n1309), .B(n373), .Z(n3730) );
  XNOR U382 ( .A(in[1446]), .B(n3730), .Z(n2828) );
  NAND U383 ( .A(n2831), .B(n2828), .Z(n228) );
  XNOR U384 ( .A(n2550), .B(n228), .Z(out[100]) );
  XOR U385 ( .A(in[1396]), .B(in[116]), .Z(n230) );
  XNOR U386 ( .A(in[1076]), .B(in[756]), .Z(n229) );
  XNOR U387 ( .A(n230), .B(n229), .Z(n231) );
  XOR U388 ( .A(in[436]), .B(n231), .Z(n1428) );
  XOR U389 ( .A(in[1525]), .B(in[565]), .Z(n233) );
  XNOR U390 ( .A(in[885]), .B(in[245]), .Z(n232) );
  XNOR U391 ( .A(n233), .B(n232), .Z(n234) );
  XOR U392 ( .A(in[1205]), .B(n234), .Z(n1370) );
  XNOR U393 ( .A(n1428), .B(n1370), .Z(n3794) );
  XNOR U394 ( .A(in[181]), .B(n3794), .Z(n1342) );
  XOR U395 ( .A(in[341]), .B(in[661]), .Z(n236) );
  XNOR U396 ( .A(in[21]), .B(in[1301]), .Z(n235) );
  XNOR U397 ( .A(n236), .B(n235), .Z(n237) );
  XOR U398 ( .A(in[981]), .B(n237), .Z(n1251) );
  XOR U399 ( .A(in[150]), .B(in[1430]), .Z(n239) );
  XNOR U400 ( .A(in[1110]), .B(in[790]), .Z(n238) );
  XNOR U401 ( .A(n239), .B(n238), .Z(n240) );
  XNOR U402 ( .A(in[470]), .B(n240), .Z(n548) );
  XNOR U403 ( .A(n1251), .B(n548), .Z(n4129) );
  XNOR U404 ( .A(in[1366]), .B(n4129), .Z(n1737) );
  XOR U405 ( .A(in[1374]), .B(in[734]), .Z(n242) );
  XNOR U406 ( .A(in[94]), .B(in[414]), .Z(n241) );
  XNOR U407 ( .A(n242), .B(n241), .Z(n243) );
  XOR U408 ( .A(in[1054]), .B(n243), .Z(n916) );
  XOR U409 ( .A(in[1565]), .B(in[605]), .Z(n245) );
  XNOR U410 ( .A(in[925]), .B(in[285]), .Z(n244) );
  XNOR U411 ( .A(n245), .B(n244), .Z(n246) );
  XOR U412 ( .A(in[1245]), .B(n246), .Z(n650) );
  XNOR U413 ( .A(n916), .B(n650), .Z(n3904) );
  XNOR U414 ( .A(in[990]), .B(n3904), .Z(n1734) );
  NAND U415 ( .A(n1737), .B(n1734), .Z(n247) );
  XNOR U416 ( .A(n1342), .B(n247), .Z(out[1010]) );
  XOR U417 ( .A(in[1526]), .B(in[566]), .Z(n249) );
  XNOR U418 ( .A(in[886]), .B(in[246]), .Z(n248) );
  XNOR U419 ( .A(n249), .B(n248), .Z(n250) );
  XOR U420 ( .A(in[1206]), .B(n250), .Z(n1374) );
  XOR U421 ( .A(in[1397]), .B(in[117]), .Z(n252) );
  XNOR U422 ( .A(in[1077]), .B(in[757]), .Z(n251) );
  XNOR U423 ( .A(n252), .B(n251), .Z(n253) );
  XOR U424 ( .A(in[437]), .B(n253), .Z(n1432) );
  XNOR U425 ( .A(n1374), .B(n1432), .Z(n3804) );
  XNOR U426 ( .A(in[182]), .B(n3804), .Z(n1346) );
  XOR U427 ( .A(in[151]), .B(in[1431]), .Z(n255) );
  XNOR U428 ( .A(in[1111]), .B(in[791]), .Z(n254) );
  XNOR U429 ( .A(n255), .B(n254), .Z(n256) );
  XOR U430 ( .A(in[471]), .B(n256), .Z(n563) );
  XOR U431 ( .A(in[342]), .B(in[662]), .Z(n258) );
  XNOR U432 ( .A(in[22]), .B(in[1302]), .Z(n257) );
  XNOR U433 ( .A(n258), .B(n257), .Z(n259) );
  XNOR U434 ( .A(in[982]), .B(n259), .Z(n1254) );
  XNOR U435 ( .A(n563), .B(n1254), .Z(n4132) );
  XNOR U436 ( .A(in[1367]), .B(n4132), .Z(n1741) );
  XOR U437 ( .A(in[1375]), .B(in[735]), .Z(n261) );
  XNOR U438 ( .A(in[95]), .B(in[415]), .Z(n260) );
  XNOR U439 ( .A(n261), .B(n260), .Z(n262) );
  XOR U440 ( .A(in[1055]), .B(n262), .Z(n929) );
  XOR U441 ( .A(in[1566]), .B(in[606]), .Z(n264) );
  XNOR U442 ( .A(in[926]), .B(in[286]), .Z(n263) );
  XNOR U443 ( .A(n264), .B(n263), .Z(n265) );
  XOR U444 ( .A(in[1246]), .B(n265), .Z(n665) );
  XNOR U445 ( .A(n929), .B(n665), .Z(n3906) );
  XNOR U446 ( .A(in[991]), .B(n3906), .Z(n1738) );
  NAND U447 ( .A(n1741), .B(n1738), .Z(n266) );
  XNOR U448 ( .A(n1346), .B(n266), .Z(out[1011]) );
  XOR U449 ( .A(in[1527]), .B(in[567]), .Z(n268) );
  XNOR U450 ( .A(in[887]), .B(in[247]), .Z(n267) );
  XNOR U451 ( .A(n268), .B(n267), .Z(n269) );
  XOR U452 ( .A(in[1207]), .B(n269), .Z(n1378) );
  XOR U453 ( .A(in[1398]), .B(in[118]), .Z(n271) );
  XNOR U454 ( .A(in[1078]), .B(in[758]), .Z(n270) );
  XNOR U455 ( .A(n271), .B(n270), .Z(n272) );
  XOR U456 ( .A(in[438]), .B(n272), .Z(n1436) );
  XNOR U457 ( .A(n1378), .B(n1436), .Z(n3808) );
  XNOR U458 ( .A(in[183]), .B(n3808), .Z(n1351) );
  XOR U459 ( .A(in[343]), .B(in[663]), .Z(n274) );
  XNOR U460 ( .A(in[23]), .B(in[1303]), .Z(n273) );
  XNOR U461 ( .A(n274), .B(n273), .Z(n275) );
  XOR U462 ( .A(in[983]), .B(n275), .Z(n1257) );
  XOR U463 ( .A(in[152]), .B(in[1432]), .Z(n277) );
  XNOR U464 ( .A(in[1112]), .B(in[792]), .Z(n276) );
  XNOR U465 ( .A(n277), .B(n276), .Z(n278) );
  XNOR U466 ( .A(in[472]), .B(n278), .Z(n589) );
  XNOR U467 ( .A(n1257), .B(n589), .Z(n4135) );
  XNOR U468 ( .A(in[1368]), .B(n4135), .Z(n1745) );
  XOR U469 ( .A(in[1376]), .B(in[736]), .Z(n280) );
  XNOR U470 ( .A(in[96]), .B(in[416]), .Z(n279) );
  XNOR U471 ( .A(n280), .B(n279), .Z(n281) );
  XOR U472 ( .A(in[1056]), .B(n281), .Z(n944) );
  XOR U473 ( .A(in[1567]), .B(in[607]), .Z(n283) );
  XNOR U474 ( .A(in[927]), .B(in[287]), .Z(n282) );
  XNOR U475 ( .A(n283), .B(n282), .Z(n284) );
  XOR U476 ( .A(in[1247]), .B(n284), .Z(n680) );
  XNOR U477 ( .A(n944), .B(n680), .Z(n3908) );
  XNOR U478 ( .A(in[992]), .B(n3908), .Z(n1742) );
  NAND U479 ( .A(n1745), .B(n1742), .Z(n285) );
  XNOR U480 ( .A(n1351), .B(n285), .Z(out[1012]) );
  XOR U481 ( .A(in[1528]), .B(in[568]), .Z(n287) );
  XNOR U482 ( .A(in[888]), .B(in[248]), .Z(n286) );
  XNOR U483 ( .A(n287), .B(n286), .Z(n288) );
  XOR U484 ( .A(in[1208]), .B(n288), .Z(n1382) );
  XOR U485 ( .A(in[1399]), .B(in[119]), .Z(n290) );
  XNOR U486 ( .A(in[1079]), .B(in[759]), .Z(n289) );
  XNOR U487 ( .A(n290), .B(n289), .Z(n291) );
  XOR U488 ( .A(in[439]), .B(n291), .Z(n1440) );
  XNOR U489 ( .A(n1382), .B(n1440), .Z(n3812) );
  XNOR U490 ( .A(in[184]), .B(n3812), .Z(n1355) );
  XOR U491 ( .A(in[153]), .B(in[1433]), .Z(n293) );
  XNOR U492 ( .A(in[1113]), .B(in[793]), .Z(n292) );
  XNOR U493 ( .A(n293), .B(n292), .Z(n294) );
  XOR U494 ( .A(in[473]), .B(n294), .Z(n604) );
  XOR U495 ( .A(in[344]), .B(in[664]), .Z(n296) );
  XNOR U496 ( .A(in[24]), .B(in[1304]), .Z(n295) );
  XNOR U497 ( .A(n296), .B(n295), .Z(n297) );
  XNOR U498 ( .A(in[984]), .B(n297), .Z(n1260) );
  XNOR U499 ( .A(n604), .B(n1260), .Z(n4138) );
  XNOR U500 ( .A(in[1369]), .B(n4138), .Z(n1749) );
  XOR U501 ( .A(in[1377]), .B(in[737]), .Z(n299) );
  XNOR U502 ( .A(in[97]), .B(in[417]), .Z(n298) );
  XNOR U503 ( .A(n299), .B(n298), .Z(n300) );
  XOR U504 ( .A(in[1057]), .B(n300), .Z(n959) );
  XOR U505 ( .A(in[1568]), .B(in[608]), .Z(n302) );
  XNOR U506 ( .A(in[928]), .B(in[288]), .Z(n301) );
  XNOR U507 ( .A(n302), .B(n301), .Z(n303) );
  XOR U508 ( .A(in[1248]), .B(n303), .Z(n695) );
  XNOR U509 ( .A(n959), .B(n695), .Z(n3910) );
  XNOR U510 ( .A(in[993]), .B(n3910), .Z(n1746) );
  NAND U511 ( .A(n1749), .B(n1746), .Z(n304) );
  XNOR U512 ( .A(n1355), .B(n304), .Z(out[1013]) );
  XOR U513 ( .A(in[1529]), .B(in[569]), .Z(n306) );
  XNOR U514 ( .A(in[889]), .B(in[249]), .Z(n305) );
  XNOR U515 ( .A(n306), .B(n305), .Z(n307) );
  XOR U516 ( .A(in[1209]), .B(n307), .Z(n1386) );
  XOR U517 ( .A(in[1400]), .B(in[120]), .Z(n309) );
  XNOR U518 ( .A(in[1080]), .B(in[760]), .Z(n308) );
  XNOR U519 ( .A(n309), .B(n308), .Z(n310) );
  XOR U520 ( .A(in[440]), .B(n310), .Z(n1444) );
  XNOR U521 ( .A(n1386), .B(n1444), .Z(n3816) );
  XNOR U522 ( .A(in[185]), .B(n3816), .Z(n1359) );
  XOR U523 ( .A(in[345]), .B(in[665]), .Z(n312) );
  XNOR U524 ( .A(in[25]), .B(in[1305]), .Z(n311) );
  XNOR U525 ( .A(n312), .B(n311), .Z(n313) );
  XOR U526 ( .A(in[985]), .B(n313), .Z(n1263) );
  XOR U527 ( .A(in[154]), .B(in[1434]), .Z(n315) );
  XNOR U528 ( .A(in[1114]), .B(in[794]), .Z(n314) );
  XNOR U529 ( .A(n315), .B(n314), .Z(n316) );
  XNOR U530 ( .A(in[474]), .B(n316), .Z(n619) );
  XNOR U531 ( .A(n1263), .B(n619), .Z(n4141) );
  XNOR U532 ( .A(in[1370]), .B(n4141), .Z(n1754) );
  XOR U533 ( .A(in[1569]), .B(in[609]), .Z(n318) );
  XNOR U534 ( .A(in[929]), .B(in[289]), .Z(n317) );
  XNOR U535 ( .A(n318), .B(n317), .Z(n319) );
  XOR U536 ( .A(in[1249]), .B(n319), .Z(n710) );
  XOR U537 ( .A(in[1378]), .B(in[738]), .Z(n321) );
  XNOR U538 ( .A(in[98]), .B(in[418]), .Z(n320) );
  XNOR U539 ( .A(n321), .B(n320), .Z(n322) );
  XOR U540 ( .A(in[1058]), .B(n322), .Z(n974) );
  XNOR U541 ( .A(n710), .B(n974), .Z(n3912) );
  XNOR U542 ( .A(in[994]), .B(n3912), .Z(n1751) );
  NAND U543 ( .A(n1754), .B(n1751), .Z(n323) );
  XNOR U544 ( .A(n1359), .B(n323), .Z(out[1014]) );
  XOR U545 ( .A(in[1401]), .B(in[121]), .Z(n325) );
  XNOR U546 ( .A(in[1081]), .B(in[761]), .Z(n324) );
  XNOR U547 ( .A(n325), .B(n324), .Z(n326) );
  XOR U548 ( .A(in[441]), .B(n326), .Z(n1448) );
  XNOR U549 ( .A(n327), .B(n1448), .Z(n3538) );
  XNOR U550 ( .A(in[186]), .B(n3538), .Z(n1363) );
  XOR U551 ( .A(in[155]), .B(in[1435]), .Z(n329) );
  XNOR U552 ( .A(in[1115]), .B(in[795]), .Z(n328) );
  XNOR U553 ( .A(n329), .B(n328), .Z(n330) );
  XOR U554 ( .A(in[475]), .B(n330), .Z(n634) );
  XOR U555 ( .A(in[346]), .B(in[666]), .Z(n332) );
  XNOR U556 ( .A(in[26]), .B(in[1306]), .Z(n331) );
  XNOR U557 ( .A(n332), .B(n331), .Z(n333) );
  XNOR U558 ( .A(in[986]), .B(n333), .Z(n1266) );
  XNOR U559 ( .A(n634), .B(n1266), .Z(n4148) );
  XNOR U560 ( .A(in[1371]), .B(n4148), .Z(n1758) );
  XOR U561 ( .A(in[1379]), .B(in[739]), .Z(n335) );
  XNOR U562 ( .A(in[99]), .B(in[419]), .Z(n334) );
  XNOR U563 ( .A(n335), .B(n334), .Z(n336) );
  XNOR U564 ( .A(in[1059]), .B(n336), .Z(n989) );
  XNOR U565 ( .A(n337), .B(n989), .Z(n3914) );
  XNOR U566 ( .A(in[995]), .B(n3914), .Z(n1755) );
  NAND U567 ( .A(n1758), .B(n1755), .Z(n338) );
  XNOR U568 ( .A(n1363), .B(n338), .Z(out[1015]) );
  XOR U569 ( .A(in[1402]), .B(in[122]), .Z(n340) );
  XNOR U570 ( .A(in[1082]), .B(in[762]), .Z(n339) );
  XNOR U571 ( .A(n340), .B(n339), .Z(n341) );
  XOR U572 ( .A(in[442]), .B(n341), .Z(n1452) );
  XOR U573 ( .A(in[1531]), .B(in[571]), .Z(n343) );
  XNOR U574 ( .A(in[1211]), .B(in[251]), .Z(n342) );
  XNOR U575 ( .A(n343), .B(n342), .Z(n344) );
  XOR U576 ( .A(in[891]), .B(n344), .Z(n416) );
  XNOR U577 ( .A(n1452), .B(n416), .Z(n3542) );
  XNOR U578 ( .A(in[187]), .B(n3542), .Z(n1367) );
  XOR U579 ( .A(in[156]), .B(in[1436]), .Z(n346) );
  XNOR U580 ( .A(in[1116]), .B(in[796]), .Z(n345) );
  XNOR U581 ( .A(n346), .B(n345), .Z(n347) );
  XOR U582 ( .A(in[476]), .B(n347), .Z(n649) );
  XOR U583 ( .A(in[347]), .B(in[667]), .Z(n349) );
  XNOR U584 ( .A(in[27]), .B(in[1307]), .Z(n348) );
  XNOR U585 ( .A(n349), .B(n348), .Z(n350) );
  XNOR U586 ( .A(in[987]), .B(n350), .Z(n1269) );
  XNOR U587 ( .A(n649), .B(n1269), .Z(n4151) );
  XNOR U588 ( .A(in[1372]), .B(n4151), .Z(n1762) );
  XOR U589 ( .A(in[1060]), .B(in[420]), .Z(n352) );
  XNOR U590 ( .A(in[740]), .B(in[1380]), .Z(n351) );
  XNOR U591 ( .A(n352), .B(n351), .Z(n353) );
  XOR U592 ( .A(in[100]), .B(n353), .Z(n1004) );
  XOR U593 ( .A(in[1571]), .B(in[611]), .Z(n355) );
  XNOR U594 ( .A(in[931]), .B(in[291]), .Z(n354) );
  XNOR U595 ( .A(n355), .B(n354), .Z(n356) );
  XOR U596 ( .A(in[1251]), .B(n356), .Z(n420) );
  XNOR U597 ( .A(n1004), .B(n420), .Z(n3916) );
  XNOR U598 ( .A(in[996]), .B(n3916), .Z(n1759) );
  NAND U599 ( .A(n1762), .B(n1759), .Z(n357) );
  XNOR U600 ( .A(n1367), .B(n357), .Z(out[1016]) );
  XOR U601 ( .A(in[1403]), .B(in[123]), .Z(n359) );
  XNOR U602 ( .A(in[1083]), .B(in[763]), .Z(n358) );
  XNOR U603 ( .A(n359), .B(n358), .Z(n360) );
  XOR U604 ( .A(in[443]), .B(n360), .Z(n1456) );
  XOR U605 ( .A(in[1532]), .B(in[572]), .Z(n362) );
  XNOR U606 ( .A(in[1212]), .B(in[252]), .Z(n361) );
  XNOR U607 ( .A(n362), .B(n361), .Z(n363) );
  XOR U608 ( .A(in[892]), .B(n363), .Z(n581) );
  XNOR U609 ( .A(n1456), .B(n581), .Z(n3546) );
  XNOR U610 ( .A(in[188]), .B(n3546), .Z(n1371) );
  XOR U611 ( .A(in[157]), .B(in[1437]), .Z(n365) );
  XNOR U612 ( .A(in[1117]), .B(in[797]), .Z(n364) );
  XNOR U613 ( .A(n365), .B(n364), .Z(n366) );
  XOR U614 ( .A(in[477]), .B(n366), .Z(n664) );
  XOR U615 ( .A(in[348]), .B(in[668]), .Z(n368) );
  XNOR U616 ( .A(in[28]), .B(in[1308]), .Z(n367) );
  XNOR U617 ( .A(n368), .B(n367), .Z(n369) );
  XNOR U618 ( .A(in[988]), .B(n369), .Z(n1272) );
  XNOR U619 ( .A(n664), .B(n1272), .Z(n4154) );
  XNOR U620 ( .A(in[1373]), .B(n4154), .Z(n1766) );
  XOR U621 ( .A(in[1572]), .B(in[612]), .Z(n371) );
  XNOR U622 ( .A(in[932]), .B(in[292]), .Z(n370) );
  XNOR U623 ( .A(n371), .B(n370), .Z(n372) );
  XOR U624 ( .A(in[1252]), .B(n372), .Z(n583) );
  XNOR U625 ( .A(n373), .B(n583), .Z(n3918) );
  XNOR U626 ( .A(in[997]), .B(n3918), .Z(n1763) );
  NAND U627 ( .A(n1766), .B(n1763), .Z(n374) );
  XNOR U628 ( .A(n1371), .B(n374), .Z(out[1017]) );
  XOR U629 ( .A(in[1404]), .B(in[124]), .Z(n376) );
  XNOR U630 ( .A(in[1084]), .B(in[764]), .Z(n375) );
  XNOR U631 ( .A(n376), .B(n375), .Z(n377) );
  XOR U632 ( .A(in[444]), .B(n377), .Z(n1460) );
  XOR U633 ( .A(in[1533]), .B(in[573]), .Z(n379) );
  XNOR U634 ( .A(in[1213]), .B(in[253]), .Z(n378) );
  XNOR U635 ( .A(n379), .B(n378), .Z(n380) );
  XOR U636 ( .A(in[893]), .B(n380), .Z(n740) );
  XNOR U637 ( .A(n1460), .B(n740), .Z(n3550) );
  XNOR U638 ( .A(in[189]), .B(n3550), .Z(n1375) );
  XOR U639 ( .A(in[158]), .B(in[1438]), .Z(n382) );
  XNOR U640 ( .A(in[1118]), .B(in[798]), .Z(n381) );
  XNOR U641 ( .A(n382), .B(n381), .Z(n383) );
  XOR U642 ( .A(in[478]), .B(n383), .Z(n679) );
  XOR U643 ( .A(in[349]), .B(in[669]), .Z(n385) );
  XNOR U644 ( .A(in[29]), .B(in[1309]), .Z(n384) );
  XNOR U645 ( .A(n385), .B(n384), .Z(n386) );
  XNOR U646 ( .A(in[989]), .B(n386), .Z(n1276) );
  XNOR U647 ( .A(n679), .B(n1276), .Z(n4157) );
  XNOR U648 ( .A(in[1374]), .B(n4157), .Z(n1770) );
  XOR U649 ( .A(in[1062]), .B(in[422]), .Z(n388) );
  XNOR U650 ( .A(in[742]), .B(in[1382]), .Z(n387) );
  XNOR U651 ( .A(n388), .B(n387), .Z(n389) );
  XOR U652 ( .A(in[102]), .B(n389), .Z(n424) );
  XOR U653 ( .A(in[1573]), .B(in[613]), .Z(n391) );
  XNOR U654 ( .A(in[933]), .B(in[293]), .Z(n390) );
  XNOR U655 ( .A(n391), .B(n390), .Z(n392) );
  XOR U656 ( .A(in[1253]), .B(n392), .Z(n742) );
  XNOR U657 ( .A(n424), .B(n742), .Z(n3924) );
  XNOR U658 ( .A(in[998]), .B(n3924), .Z(n1767) );
  NAND U659 ( .A(n1770), .B(n1767), .Z(n393) );
  XNOR U660 ( .A(n1375), .B(n393), .Z(out[1018]) );
  XOR U661 ( .A(in[1405]), .B(in[125]), .Z(n395) );
  XNOR U662 ( .A(in[1085]), .B(in[765]), .Z(n394) );
  XNOR U663 ( .A(n395), .B(n394), .Z(n396) );
  XOR U664 ( .A(in[445]), .B(n396), .Z(n1464) );
  XOR U665 ( .A(in[1534]), .B(in[894]), .Z(n398) );
  XNOR U666 ( .A(in[574]), .B(in[1214]), .Z(n397) );
  XNOR U667 ( .A(n398), .B(n397), .Z(n399) );
  XOR U668 ( .A(in[254]), .B(n399), .Z(n877) );
  XNOR U669 ( .A(n1464), .B(n877), .Z(n3554) );
  XNOR U670 ( .A(in[190]), .B(n3554), .Z(n1379) );
  XOR U671 ( .A(in[1439]), .B(in[479]), .Z(n401) );
  XNOR U672 ( .A(in[799]), .B(in[159]), .Z(n400) );
  XNOR U673 ( .A(n401), .B(n400), .Z(n402) );
  XOR U674 ( .A(in[1119]), .B(n402), .Z(n694) );
  XOR U675 ( .A(in[350]), .B(in[670]), .Z(n404) );
  XNOR U676 ( .A(in[30]), .B(in[1310]), .Z(n403) );
  XNOR U677 ( .A(n404), .B(n403), .Z(n405) );
  XNOR U678 ( .A(in[990]), .B(n405), .Z(n1279) );
  XNOR U679 ( .A(n694), .B(n1279), .Z(n4160) );
  XNOR U680 ( .A(in[1375]), .B(n4160), .Z(n1774) );
  XOR U681 ( .A(in[1063]), .B(in[423]), .Z(n407) );
  XNOR U682 ( .A(in[743]), .B(in[1383]), .Z(n406) );
  XNOR U683 ( .A(n407), .B(n406), .Z(n408) );
  XOR U684 ( .A(in[103]), .B(n408), .Z(n587) );
  XOR U685 ( .A(in[1574]), .B(in[614]), .Z(n410) );
  XNOR U686 ( .A(in[934]), .B(in[294]), .Z(n409) );
  XNOR U687 ( .A(n410), .B(n409), .Z(n411) );
  XOR U688 ( .A(in[1254]), .B(n411), .Z(n786) );
  XNOR U689 ( .A(n587), .B(n786), .Z(n3926) );
  XNOR U690 ( .A(in[999]), .B(n3926), .Z(n1771) );
  NAND U691 ( .A(n1774), .B(n1771), .Z(n412) );
  XNOR U692 ( .A(n1379), .B(n412), .Z(out[1019]) );
  XOR U693 ( .A(in[1340]), .B(in[60]), .Z(n414) );
  XNOR U694 ( .A(in[700]), .B(in[380]), .Z(n413) );
  XNOR U695 ( .A(n414), .B(n413), .Z(n415) );
  XOR U696 ( .A(in[1020]), .B(n415), .Z(n871) );
  XNOR U697 ( .A(n416), .B(n871), .Z(n3596) );
  XNOR U698 ( .A(in[636]), .B(n3596), .Z(n2552) );
  XOR U699 ( .A(in[162]), .B(in[1442]), .Z(n418) );
  XNOR U700 ( .A(in[802]), .B(in[1122]), .Z(n417) );
  XNOR U701 ( .A(n418), .B(n417), .Z(n419) );
  XNOR U702 ( .A(in[482]), .B(n419), .Z(n471) );
  XNOR U703 ( .A(n420), .B(n471), .Z(n3693) );
  XNOR U704 ( .A(in[227]), .B(n3693), .Z(n2845) );
  XOR U705 ( .A(in[1511]), .B(in[551]), .Z(n422) );
  XNOR U706 ( .A(in[871]), .B(in[231]), .Z(n421) );
  XNOR U707 ( .A(n422), .B(n421), .Z(n423) );
  XOR U708 ( .A(in[1191]), .B(n423), .Z(n1313) );
  XNOR U709 ( .A(n424), .B(n1313), .Z(n3734) );
  XNOR U710 ( .A(in[1447]), .B(n3734), .Z(n2842) );
  NAND U711 ( .A(n2845), .B(n2842), .Z(n425) );
  XNOR U712 ( .A(n2552), .B(n425), .Z(out[101]) );
  XOR U713 ( .A(in[1406]), .B(in[126]), .Z(n427) );
  XNOR U714 ( .A(in[1086]), .B(in[766]), .Z(n426) );
  XNOR U715 ( .A(n427), .B(n426), .Z(n428) );
  XOR U716 ( .A(in[446]), .B(n428), .Z(n1469) );
  XOR U717 ( .A(in[1535]), .B(in[575]), .Z(n430) );
  XNOR U718 ( .A(in[895]), .B(in[255]), .Z(n429) );
  XNOR U719 ( .A(n430), .B(n429), .Z(n431) );
  XOR U720 ( .A(in[1215]), .B(n431), .Z(n1024) );
  XNOR U721 ( .A(n1469), .B(n1024), .Z(n3558) );
  XNOR U722 ( .A(in[191]), .B(n3558), .Z(n1383) );
  XOR U723 ( .A(in[1440]), .B(in[480]), .Z(n433) );
  XNOR U724 ( .A(in[800]), .B(in[160]), .Z(n432) );
  XNOR U725 ( .A(n433), .B(n432), .Z(n434) );
  XOR U726 ( .A(in[1120]), .B(n434), .Z(n709) );
  XOR U727 ( .A(in[351]), .B(in[671]), .Z(n436) );
  XNOR U728 ( .A(in[31]), .B(in[1311]), .Z(n435) );
  XNOR U729 ( .A(n436), .B(n435), .Z(n437) );
  XNOR U730 ( .A(in[991]), .B(n437), .Z(n1282) );
  XNOR U731 ( .A(n709), .B(n1282), .Z(n4163) );
  XNOR U732 ( .A(in[1376]), .B(n4163), .Z(n1778) );
  XOR U733 ( .A(in[1064]), .B(in[424]), .Z(n439) );
  XNOR U734 ( .A(in[744]), .B(in[1384]), .Z(n438) );
  XNOR U735 ( .A(n439), .B(n438), .Z(n440) );
  XOR U736 ( .A(in[104]), .B(n440), .Z(n746) );
  XOR U737 ( .A(in[1575]), .B(in[615]), .Z(n442) );
  XNOR U738 ( .A(in[935]), .B(in[295]), .Z(n441) );
  XNOR U739 ( .A(n442), .B(n441), .Z(n443) );
  XOR U740 ( .A(in[1255]), .B(n443), .Z(n799) );
  XNOR U741 ( .A(n746), .B(n799), .Z(n3928) );
  XNOR U742 ( .A(in[1000]), .B(n3928), .Z(n1775) );
  NAND U743 ( .A(n1778), .B(n1775), .Z(n444) );
  XNOR U744 ( .A(n1383), .B(n444), .Z(out[1020]) );
  XOR U745 ( .A(in[1407]), .B(in[127]), .Z(n446) );
  XNOR U746 ( .A(in[1087]), .B(in[767]), .Z(n445) );
  XNOR U747 ( .A(n446), .B(n445), .Z(n447) );
  XOR U748 ( .A(in[447]), .B(n447), .Z(n1472) );
  XOR U749 ( .A(in[1472]), .B(in[512]), .Z(n449) );
  XNOR U750 ( .A(in[832]), .B(in[192]), .Z(n448) );
  XNOR U751 ( .A(n449), .B(n448), .Z(n450) );
  XOR U752 ( .A(in[1152]), .B(n450), .Z(n1091) );
  XNOR U753 ( .A(n1472), .B(n1091), .Z(n3562) );
  XNOR U754 ( .A(in[128]), .B(n3562), .Z(n1387) );
  XOR U755 ( .A(in[352]), .B(in[672]), .Z(n452) );
  XNOR U756 ( .A(in[32]), .B(in[1312]), .Z(n451) );
  XNOR U757 ( .A(n452), .B(n451), .Z(n453) );
  XNOR U758 ( .A(in[992]), .B(n453), .Z(n1285) );
  XNOR U759 ( .A(n454), .B(n1285), .Z(n4166) );
  XNOR U760 ( .A(in[1377]), .B(n4166), .Z(n1782) );
  XOR U761 ( .A(in[1065]), .B(in[425]), .Z(n456) );
  XNOR U762 ( .A(in[745]), .B(in[1385]), .Z(n455) );
  XNOR U763 ( .A(n456), .B(n455), .Z(n457) );
  XOR U764 ( .A(in[105]), .B(n457), .Z(n881) );
  XOR U765 ( .A(in[1576]), .B(in[616]), .Z(n459) );
  XNOR U766 ( .A(in[936]), .B(in[296]), .Z(n458) );
  XNOR U767 ( .A(n459), .B(n458), .Z(n460) );
  XOR U768 ( .A(in[1256]), .B(n460), .Z(n812) );
  XNOR U769 ( .A(n881), .B(n812), .Z(n3930) );
  XNOR U770 ( .A(in[1001]), .B(n3930), .Z(n1779) );
  NAND U771 ( .A(n1782), .B(n1779), .Z(n461) );
  XNOR U772 ( .A(n1387), .B(n461), .Z(out[1021]) );
  XOR U773 ( .A(in[1344]), .B(in[64]), .Z(n463) );
  XNOR U774 ( .A(in[1024]), .B(in[384]), .Z(n462) );
  XNOR U775 ( .A(n463), .B(n462), .Z(n464) );
  XOR U776 ( .A(in[704]), .B(n464), .Z(n1477) );
  XOR U777 ( .A(in[1473]), .B(in[513]), .Z(n466) );
  XNOR U778 ( .A(in[833]), .B(in[193]), .Z(n465) );
  XNOR U779 ( .A(n466), .B(n465), .Z(n467) );
  XOR U780 ( .A(in[1153]), .B(n467), .Z(n1144) );
  XNOR U781 ( .A(n1477), .B(n1144), .Z(n3566) );
  XNOR U782 ( .A(in[129]), .B(n3566), .Z(n1390) );
  XOR U783 ( .A(in[353]), .B(in[673]), .Z(n469) );
  XNOR U784 ( .A(in[33]), .B(in[1313]), .Z(n468) );
  XNOR U785 ( .A(n469), .B(n468), .Z(n470) );
  XOR U786 ( .A(in[993]), .B(n470), .Z(n1288) );
  XNOR U787 ( .A(n1288), .B(n471), .Z(n4169) );
  XNOR U788 ( .A(in[1378]), .B(n4169), .Z(n1786) );
  XOR U789 ( .A(in[1577]), .B(in[617]), .Z(n473) );
  XNOR U790 ( .A(in[937]), .B(in[297]), .Z(n472) );
  XNOR U791 ( .A(n473), .B(n472), .Z(n474) );
  XOR U792 ( .A(in[1257]), .B(n474), .Z(n825) );
  XNOR U793 ( .A(n475), .B(n825), .Z(n3932) );
  XNOR U794 ( .A(in[1002]), .B(n3932), .Z(n1783) );
  NAND U795 ( .A(n1786), .B(n1783), .Z(n476) );
  XNOR U796 ( .A(n1390), .B(n476), .Z(out[1022]) );
  XOR U797 ( .A(n3570), .B(in[130]), .Z(n1392) );
  XOR U798 ( .A(in[163]), .B(in[1443]), .Z(n478) );
  XNOR U799 ( .A(in[803]), .B(in[1123]), .Z(n477) );
  XNOR U800 ( .A(n478), .B(n477), .Z(n479) );
  XOR U801 ( .A(in[483]), .B(n479), .Z(n582) );
  XOR U802 ( .A(in[354]), .B(in[674]), .Z(n481) );
  XNOR U803 ( .A(in[34]), .B(in[1314]), .Z(n480) );
  XNOR U804 ( .A(n481), .B(n480), .Z(n482) );
  XNOR U805 ( .A(in[994]), .B(n482), .Z(n1291) );
  XNOR U806 ( .A(n582), .B(n1291), .Z(n4172) );
  XNOR U807 ( .A(in[1379]), .B(n4172), .Z(n1790) );
  XOR U808 ( .A(in[1578]), .B(in[618]), .Z(n484) );
  XNOR U809 ( .A(in[938]), .B(in[298]), .Z(n483) );
  XNOR U810 ( .A(n484), .B(n483), .Z(n485) );
  XOR U811 ( .A(in[1258]), .B(n485), .Z(n838) );
  XNOR U812 ( .A(n486), .B(n838), .Z(n3934) );
  XNOR U813 ( .A(in[1003]), .B(n3934), .Z(n1787) );
  NAND U814 ( .A(n1790), .B(n1787), .Z(n487) );
  XNOR U815 ( .A(n1392), .B(n487), .Z(out[1023]) );
  XNOR U816 ( .A(n489), .B(n488), .Z(n3625) );
  XNOR U817 ( .A(in[531]), .B(n3625), .Z(n1396) );
  XOR U818 ( .A(in[1346]), .B(in[66]), .Z(n491) );
  XNOR U819 ( .A(in[1026]), .B(in[386]), .Z(n490) );
  XNOR U820 ( .A(n491), .B(n490), .Z(n492) );
  XOR U821 ( .A(in[706]), .B(n492), .Z(n1485) );
  XOR U822 ( .A(in[1475]), .B(in[515]), .Z(n494) );
  XNOR U823 ( .A(in[835]), .B(in[195]), .Z(n493) );
  XNOR U824 ( .A(n494), .B(n493), .Z(n495) );
  XNOR U825 ( .A(in[1155]), .B(n495), .Z(n1196) );
  XNOR U826 ( .A(n1485), .B(n1196), .Z(n3574) );
  XNOR U827 ( .A(in[131]), .B(n3574), .Z(n4631) );
  XOR U828 ( .A(in[35]), .B(in[675]), .Z(n497) );
  XNOR U829 ( .A(in[355]), .B(in[1315]), .Z(n496) );
  XNOR U830 ( .A(n497), .B(n496), .Z(n498) );
  XOR U831 ( .A(in[995]), .B(n498), .Z(n1294) );
  XOR U832 ( .A(in[164]), .B(in[1444]), .Z(n500) );
  XNOR U833 ( .A(in[804]), .B(in[1124]), .Z(n499) );
  XNOR U834 ( .A(n500), .B(n499), .Z(n501) );
  XOR U835 ( .A(in[484]), .B(n501), .Z(n741) );
  XNOR U836 ( .A(n1294), .B(n741), .Z(n4175) );
  XNOR U837 ( .A(in[1380]), .B(n4175), .Z(n4628) );
  NAND U838 ( .A(n4631), .B(n4628), .Z(n502) );
  XNOR U839 ( .A(n1396), .B(n502), .Z(out[1024]) );
  XOR U840 ( .A(n504), .B(n503), .Z(n3629) );
  XNOR U841 ( .A(in[532]), .B(n3629), .Z(n1400) );
  XOR U842 ( .A(in[1347]), .B(in[67]), .Z(n506) );
  XNOR U843 ( .A(in[1027]), .B(in[387]), .Z(n505) );
  XNOR U844 ( .A(n506), .B(n505), .Z(n507) );
  XOR U845 ( .A(in[707]), .B(n507), .Z(n1489) );
  XOR U846 ( .A(in[1476]), .B(in[516]), .Z(n509) );
  XNOR U847 ( .A(in[836]), .B(in[196]), .Z(n508) );
  XNOR U848 ( .A(n509), .B(n508), .Z(n510) );
  XNOR U849 ( .A(in[1156]), .B(n510), .Z(n1199) );
  XNOR U850 ( .A(n1489), .B(n1199), .Z(n3582) );
  XNOR U851 ( .A(in[132]), .B(n3582), .Z(n4635) );
  XOR U852 ( .A(in[1445]), .B(in[165]), .Z(n512) );
  XNOR U853 ( .A(in[805]), .B(in[1125]), .Z(n511) );
  XNOR U854 ( .A(n512), .B(n511), .Z(n513) );
  XOR U855 ( .A(in[485]), .B(n513), .Z(n785) );
  XOR U856 ( .A(in[36]), .B(in[676]), .Z(n515) );
  XNOR U857 ( .A(in[356]), .B(in[1316]), .Z(n514) );
  XNOR U858 ( .A(n515), .B(n514), .Z(n516) );
  XOR U859 ( .A(in[996]), .B(n516), .Z(n1297) );
  XNOR U860 ( .A(n785), .B(n1297), .Z(n4182) );
  XNOR U861 ( .A(in[1381]), .B(n4182), .Z(n4632) );
  NAND U862 ( .A(n4635), .B(n4632), .Z(n517) );
  XNOR U863 ( .A(n1400), .B(n517), .Z(out[1025]) );
  XNOR U864 ( .A(n519), .B(n518), .Z(n3633) );
  XNOR U865 ( .A(in[533]), .B(n3633), .Z(n1404) );
  XOR U866 ( .A(in[1348]), .B(in[68]), .Z(n521) );
  XNOR U867 ( .A(in[1028]), .B(in[388]), .Z(n520) );
  XNOR U868 ( .A(n521), .B(n520), .Z(n522) );
  XOR U869 ( .A(in[708]), .B(n522), .Z(n1493) );
  XOR U870 ( .A(in[1477]), .B(in[517]), .Z(n524) );
  XNOR U871 ( .A(in[837]), .B(in[197]), .Z(n523) );
  XNOR U872 ( .A(n524), .B(n523), .Z(n525) );
  XNOR U873 ( .A(in[1157]), .B(n525), .Z(n1202) );
  XNOR U874 ( .A(n1493), .B(n1202), .Z(n3586) );
  XNOR U875 ( .A(in[133]), .B(n3586), .Z(n4639) );
  XOR U876 ( .A(in[37]), .B(in[677]), .Z(n527) );
  XNOR U877 ( .A(in[357]), .B(in[1317]), .Z(n526) );
  XNOR U878 ( .A(n527), .B(n526), .Z(n528) );
  XOR U879 ( .A(in[997]), .B(n528), .Z(n1300) );
  XOR U880 ( .A(in[166]), .B(in[806]), .Z(n530) );
  XNOR U881 ( .A(in[1126]), .B(in[486]), .Z(n529) );
  XNOR U882 ( .A(n530), .B(n529), .Z(n531) );
  XOR U883 ( .A(in[1446]), .B(n531), .Z(n798) );
  XNOR U884 ( .A(n1300), .B(n798), .Z(n4185) );
  XNOR U885 ( .A(in[1382]), .B(n4185), .Z(n4636) );
  NAND U886 ( .A(n4639), .B(n4636), .Z(n532) );
  XNOR U887 ( .A(n1404), .B(n532), .Z(out[1026]) );
  XOR U888 ( .A(n534), .B(n533), .Z(n3637) );
  XNOR U889 ( .A(in[534]), .B(n3637), .Z(n1408) );
  XOR U890 ( .A(in[1349]), .B(in[69]), .Z(n536) );
  XNOR U891 ( .A(in[1029]), .B(in[389]), .Z(n535) );
  XNOR U892 ( .A(n536), .B(n535), .Z(n537) );
  XOR U893 ( .A(in[709]), .B(n537), .Z(n1497) );
  XOR U894 ( .A(in[1478]), .B(in[518]), .Z(n539) );
  XNOR U895 ( .A(in[838]), .B(in[198]), .Z(n538) );
  XNOR U896 ( .A(n539), .B(n538), .Z(n540) );
  XNOR U897 ( .A(in[1158]), .B(n540), .Z(n1205) );
  XNOR U898 ( .A(n1497), .B(n1205), .Z(n3590) );
  XNOR U899 ( .A(in[134]), .B(n3590), .Z(n4643) );
  XOR U900 ( .A(in[38]), .B(in[678]), .Z(n542) );
  XNOR U901 ( .A(in[358]), .B(in[1318]), .Z(n541) );
  XNOR U902 ( .A(n542), .B(n541), .Z(n543) );
  XOR U903 ( .A(in[998]), .B(n543), .Z(n1304) );
  XOR U904 ( .A(in[167]), .B(in[807]), .Z(n545) );
  XNOR U905 ( .A(in[1127]), .B(in[487]), .Z(n544) );
  XNOR U906 ( .A(n545), .B(n544), .Z(n546) );
  XOR U907 ( .A(in[1447]), .B(n546), .Z(n811) );
  XNOR U908 ( .A(n1304), .B(n811), .Z(n3964) );
  XNOR U909 ( .A(in[1383]), .B(n3964), .Z(n4640) );
  NAND U910 ( .A(n4643), .B(n4640), .Z(n547) );
  XNOR U911 ( .A(n1408), .B(n547), .Z(out[1027]) );
  XOR U912 ( .A(n549), .B(n548), .Z(n3641) );
  XNOR U913 ( .A(in[535]), .B(n3641), .Z(n1412) );
  XOR U914 ( .A(in[1350]), .B(in[70]), .Z(n551) );
  XNOR U915 ( .A(in[1030]), .B(in[390]), .Z(n550) );
  XNOR U916 ( .A(n551), .B(n550), .Z(n552) );
  XOR U917 ( .A(in[710]), .B(n552), .Z(n1501) );
  XOR U918 ( .A(in[199]), .B(in[1479]), .Z(n554) );
  XNOR U919 ( .A(in[1159]), .B(in[839]), .Z(n553) );
  XNOR U920 ( .A(n554), .B(n553), .Z(n555) );
  XNOR U921 ( .A(in[519]), .B(n555), .Z(n1208) );
  XNOR U922 ( .A(n1501), .B(n1208), .Z(n3594) );
  XNOR U923 ( .A(in[135]), .B(n3594), .Z(n4647) );
  XOR U924 ( .A(in[39]), .B(in[679]), .Z(n557) );
  XNOR U925 ( .A(in[359]), .B(in[1319]), .Z(n556) );
  XNOR U926 ( .A(n557), .B(n556), .Z(n558) );
  XOR U927 ( .A(in[999]), .B(n558), .Z(n1308) );
  XOR U928 ( .A(in[168]), .B(in[1448]), .Z(n560) );
  XNOR U929 ( .A(in[1128]), .B(in[808]), .Z(n559) );
  XNOR U930 ( .A(n560), .B(n559), .Z(n561) );
  XOR U931 ( .A(in[488]), .B(n561), .Z(n824) );
  XNOR U932 ( .A(n1308), .B(n824), .Z(n3967) );
  XNOR U933 ( .A(in[1384]), .B(n3967), .Z(n4644) );
  NAND U934 ( .A(n4647), .B(n4644), .Z(n562) );
  XNOR U935 ( .A(n1412), .B(n562), .Z(out[1028]) );
  XNOR U936 ( .A(n564), .B(n563), .Z(n3645) );
  XNOR U937 ( .A(in[536]), .B(n3645), .Z(n1416) );
  XOR U938 ( .A(in[1351]), .B(in[711]), .Z(n566) );
  XNOR U939 ( .A(in[1031]), .B(in[391]), .Z(n565) );
  XNOR U940 ( .A(n566), .B(n565), .Z(n567) );
  XOR U941 ( .A(in[71]), .B(n567), .Z(n1505) );
  XOR U942 ( .A(in[1480]), .B(in[520]), .Z(n569) );
  XNOR U943 ( .A(in[840]), .B(in[200]), .Z(n568) );
  XNOR U944 ( .A(n569), .B(n568), .Z(n570) );
  XNOR U945 ( .A(in[1160]), .B(n570), .Z(n1213) );
  XNOR U946 ( .A(n1505), .B(n1213), .Z(n3598) );
  XNOR U947 ( .A(in[136]), .B(n3598), .Z(n4651) );
  XOR U948 ( .A(in[169]), .B(in[1449]), .Z(n572) );
  XNOR U949 ( .A(in[1129]), .B(in[809]), .Z(n571) );
  XNOR U950 ( .A(n572), .B(n571), .Z(n573) );
  XOR U951 ( .A(in[489]), .B(n573), .Z(n837) );
  XOR U952 ( .A(in[680]), .B(in[1320]), .Z(n575) );
  XNOR U953 ( .A(in[40]), .B(in[360]), .Z(n574) );
  XNOR U954 ( .A(n575), .B(n574), .Z(n576) );
  XOR U955 ( .A(in[1000]), .B(n576), .Z(n1312) );
  XNOR U956 ( .A(n837), .B(n1312), .Z(n3974) );
  XNOR U957 ( .A(in[1385]), .B(n3974), .Z(n4648) );
  NAND U958 ( .A(n4651), .B(n4648), .Z(n577) );
  XNOR U959 ( .A(n1416), .B(n577), .Z(out[1029]) );
  XOR U960 ( .A(in[1341]), .B(in[61]), .Z(n579) );
  XNOR U961 ( .A(in[701]), .B(in[381]), .Z(n578) );
  XNOR U962 ( .A(n579), .B(n578), .Z(n580) );
  XOR U963 ( .A(in[1021]), .B(n580), .Z(n894) );
  XNOR U964 ( .A(n581), .B(n894), .Z(n3600) );
  XNOR U965 ( .A(in[637]), .B(n3600), .Z(n2555) );
  XOR U966 ( .A(n583), .B(n582), .Z(n3697) );
  XNOR U967 ( .A(in[228]), .B(n3697), .Z(n2859) );
  XOR U968 ( .A(in[1512]), .B(in[552]), .Z(n585) );
  XNOR U969 ( .A(in[872]), .B(in[232]), .Z(n584) );
  XNOR U970 ( .A(n585), .B(n584), .Z(n586) );
  XOR U971 ( .A(in[1192]), .B(n586), .Z(n1317) );
  XNOR U972 ( .A(n587), .B(n1317), .Z(n3738) );
  XNOR U973 ( .A(in[1448]), .B(n3738), .Z(n2856) );
  NAND U974 ( .A(n2859), .B(n2856), .Z(n588) );
  XNOR U975 ( .A(n2555), .B(n588), .Z(out[102]) );
  XOR U976 ( .A(n590), .B(n589), .Z(n3649) );
  XNOR U977 ( .A(in[537]), .B(n3649), .Z(n1420) );
  XOR U978 ( .A(in[1352]), .B(in[712]), .Z(n592) );
  XNOR U979 ( .A(in[1032]), .B(in[392]), .Z(n591) );
  XNOR U980 ( .A(n592), .B(n591), .Z(n593) );
  XOR U981 ( .A(in[72]), .B(n593), .Z(n1510) );
  XOR U982 ( .A(in[1481]), .B(in[521]), .Z(n595) );
  XNOR U983 ( .A(in[841]), .B(in[201]), .Z(n594) );
  XNOR U984 ( .A(n595), .B(n594), .Z(n596) );
  XNOR U985 ( .A(in[1161]), .B(n596), .Z(n1216) );
  XNOR U986 ( .A(n1510), .B(n1216), .Z(n3602) );
  XNOR U987 ( .A(in[137]), .B(n3602), .Z(n4655) );
  XOR U988 ( .A(in[170]), .B(in[1450]), .Z(n598) );
  XNOR U989 ( .A(in[1130]), .B(in[810]), .Z(n597) );
  XNOR U990 ( .A(n598), .B(n597), .Z(n599) );
  XOR U991 ( .A(in[490]), .B(n599), .Z(n853) );
  XOR U992 ( .A(in[681]), .B(in[1321]), .Z(n601) );
  XNOR U993 ( .A(in[41]), .B(in[361]), .Z(n600) );
  XNOR U994 ( .A(n601), .B(n600), .Z(n602) );
  XOR U995 ( .A(in[1001]), .B(n602), .Z(n1316) );
  XNOR U996 ( .A(n853), .B(n1316), .Z(n3977) );
  XNOR U997 ( .A(in[1386]), .B(n3977), .Z(n4652) );
  NAND U998 ( .A(n4655), .B(n4652), .Z(n603) );
  XNOR U999 ( .A(n1420), .B(n603), .Z(out[1030]) );
  XNOR U1000 ( .A(n605), .B(n604), .Z(n3653) );
  XNOR U1001 ( .A(in[538]), .B(n3653), .Z(n1424) );
  XOR U1002 ( .A(in[1353]), .B(in[393]), .Z(n607) );
  XNOR U1003 ( .A(in[713]), .B(in[73]), .Z(n606) );
  XNOR U1004 ( .A(n607), .B(n606), .Z(n608) );
  XOR U1005 ( .A(in[1033]), .B(n608), .Z(n1514) );
  XOR U1006 ( .A(in[1482]), .B(in[522]), .Z(n610) );
  XNOR U1007 ( .A(in[842]), .B(in[202]), .Z(n609) );
  XNOR U1008 ( .A(n610), .B(n609), .Z(n611) );
  XNOR U1009 ( .A(in[1162]), .B(n611), .Z(n1219) );
  XNOR U1010 ( .A(n1514), .B(n1219), .Z(n3606) );
  XNOR U1011 ( .A(in[138]), .B(n3606), .Z(n4659) );
  XOR U1012 ( .A(in[811]), .B(in[491]), .Z(n613) );
  XNOR U1013 ( .A(in[1451]), .B(in[1131]), .Z(n612) );
  XNOR U1014 ( .A(n613), .B(n612), .Z(n614) );
  XOR U1015 ( .A(in[171]), .B(n614), .Z(n866) );
  XOR U1016 ( .A(in[682]), .B(in[1322]), .Z(n616) );
  XNOR U1017 ( .A(in[42]), .B(in[362]), .Z(n615) );
  XNOR U1018 ( .A(n616), .B(n615), .Z(n617) );
  XOR U1019 ( .A(in[1002]), .B(n617), .Z(n1321) );
  XNOR U1020 ( .A(n866), .B(n1321), .Z(n3980) );
  XNOR U1021 ( .A(in[1387]), .B(n3980), .Z(n4656) );
  NAND U1022 ( .A(n4659), .B(n4656), .Z(n618) );
  XNOR U1023 ( .A(n1424), .B(n618), .Z(out[1031]) );
  XOR U1024 ( .A(n620), .B(n619), .Z(n3657) );
  XNOR U1025 ( .A(in[539]), .B(n3657), .Z(n1429) );
  XOR U1026 ( .A(in[1483]), .B(in[523]), .Z(n622) );
  XNOR U1027 ( .A(in[843]), .B(in[203]), .Z(n621) );
  XNOR U1028 ( .A(n622), .B(n621), .Z(n623) );
  XOR U1029 ( .A(in[1163]), .B(n623), .Z(n1222) );
  XOR U1030 ( .A(in[1354]), .B(in[714]), .Z(n625) );
  XNOR U1031 ( .A(in[74]), .B(in[394]), .Z(n624) );
  XNOR U1032 ( .A(n625), .B(n624), .Z(n626) );
  XNOR U1033 ( .A(in[1034]), .B(n626), .Z(n1518) );
  XNOR U1034 ( .A(n1222), .B(n1518), .Z(n3610) );
  XNOR U1035 ( .A(n3610), .B(in[139]), .Z(n4663) );
  XOR U1036 ( .A(in[683]), .B(in[1323]), .Z(n628) );
  XNOR U1037 ( .A(in[43]), .B(in[363]), .Z(n627) );
  XNOR U1038 ( .A(n628), .B(n627), .Z(n629) );
  XOR U1039 ( .A(in[1003]), .B(n629), .Z(n1325) );
  XOR U1040 ( .A(in[812]), .B(in[492]), .Z(n631) );
  XNOR U1041 ( .A(in[1452]), .B(in[1132]), .Z(n630) );
  XNOR U1042 ( .A(n631), .B(n630), .Z(n632) );
  XOR U1043 ( .A(in[172]), .B(n632), .Z(n886) );
  XNOR U1044 ( .A(n1325), .B(n886), .Z(n3983) );
  XNOR U1045 ( .A(in[1388]), .B(n3983), .Z(n4660) );
  NAND U1046 ( .A(n4663), .B(n4660), .Z(n633) );
  XNOR U1047 ( .A(n1429), .B(n633), .Z(out[1032]) );
  XNOR U1048 ( .A(n635), .B(n634), .Z(n3661) );
  XNOR U1049 ( .A(in[540]), .B(n3661), .Z(n1433) );
  XOR U1050 ( .A(in[1355]), .B(in[715]), .Z(n637) );
  XNOR U1051 ( .A(in[1035]), .B(in[395]), .Z(n636) );
  XNOR U1052 ( .A(n637), .B(n636), .Z(n638) );
  XOR U1053 ( .A(in[75]), .B(n638), .Z(n1522) );
  XOR U1054 ( .A(in[1484]), .B(in[524]), .Z(n640) );
  XNOR U1055 ( .A(in[844]), .B(in[204]), .Z(n639) );
  XNOR U1056 ( .A(n640), .B(n639), .Z(n641) );
  XNOR U1057 ( .A(in[1164]), .B(n641), .Z(n1225) );
  XNOR U1058 ( .A(n1522), .B(n1225), .Z(n3614) );
  XNOR U1059 ( .A(in[140]), .B(n3614), .Z(n4667) );
  XOR U1060 ( .A(in[813]), .B(in[493]), .Z(n643) );
  XNOR U1061 ( .A(in[1453]), .B(in[1133]), .Z(n642) );
  XNOR U1062 ( .A(n643), .B(n642), .Z(n644) );
  XOR U1063 ( .A(in[173]), .B(n644), .Z(n899) );
  XOR U1064 ( .A(in[1324]), .B(in[44]), .Z(n646) );
  XNOR U1065 ( .A(in[684]), .B(in[364]), .Z(n645) );
  XNOR U1066 ( .A(n646), .B(n645), .Z(n647) );
  XOR U1067 ( .A(in[1004]), .B(n647), .Z(n1328) );
  XNOR U1068 ( .A(n899), .B(n1328), .Z(n3986) );
  XNOR U1069 ( .A(in[1389]), .B(n3986), .Z(n4664) );
  NAND U1070 ( .A(n4667), .B(n4664), .Z(n648) );
  XNOR U1071 ( .A(n1433), .B(n648), .Z(out[1033]) );
  XNOR U1072 ( .A(n650), .B(n649), .Z(n3669) );
  XNOR U1073 ( .A(in[541]), .B(n3669), .Z(n1437) );
  XOR U1074 ( .A(in[76]), .B(in[1036]), .Z(n652) );
  XNOR U1075 ( .A(in[716]), .B(in[396]), .Z(n651) );
  XNOR U1076 ( .A(n652), .B(n651), .Z(n653) );
  XOR U1077 ( .A(in[1356]), .B(n653), .Z(n1526) );
  XOR U1078 ( .A(in[1485]), .B(in[525]), .Z(n655) );
  XNOR U1079 ( .A(in[845]), .B(in[205]), .Z(n654) );
  XNOR U1080 ( .A(n655), .B(n654), .Z(n656) );
  XNOR U1081 ( .A(in[1165]), .B(n656), .Z(n1228) );
  XNOR U1082 ( .A(n1526), .B(n1228), .Z(n3618) );
  XNOR U1083 ( .A(in[141]), .B(n3618), .Z(n4675) );
  XOR U1084 ( .A(in[814]), .B(in[494]), .Z(n658) );
  XNOR U1085 ( .A(in[1454]), .B(in[1134]), .Z(n657) );
  XNOR U1086 ( .A(n658), .B(n657), .Z(n659) );
  XOR U1087 ( .A(in[174]), .B(n659), .Z(n912) );
  XOR U1088 ( .A(in[1325]), .B(in[45]), .Z(n661) );
  XNOR U1089 ( .A(in[685]), .B(in[365]), .Z(n660) );
  XNOR U1090 ( .A(n661), .B(n660), .Z(n662) );
  XOR U1091 ( .A(in[1005]), .B(n662), .Z(n1332) );
  XNOR U1092 ( .A(n912), .B(n1332), .Z(n3989) );
  XNOR U1093 ( .A(in[1390]), .B(n3989), .Z(n4672) );
  NAND U1094 ( .A(n4675), .B(n4672), .Z(n663) );
  XNOR U1095 ( .A(n1437), .B(n663), .Z(out[1034]) );
  XNOR U1096 ( .A(n665), .B(n664), .Z(n3673) );
  XNOR U1097 ( .A(in[542]), .B(n3673), .Z(n1441) );
  XOR U1098 ( .A(in[77]), .B(in[1037]), .Z(n667) );
  XNOR U1099 ( .A(in[717]), .B(in[397]), .Z(n666) );
  XNOR U1100 ( .A(n667), .B(n666), .Z(n668) );
  XOR U1101 ( .A(in[1357]), .B(n668), .Z(n1530) );
  XOR U1102 ( .A(in[1486]), .B(in[526]), .Z(n670) );
  XNOR U1103 ( .A(in[846]), .B(in[206]), .Z(n669) );
  XNOR U1104 ( .A(n670), .B(n669), .Z(n671) );
  XNOR U1105 ( .A(in[1166]), .B(n671), .Z(n1231) );
  XNOR U1106 ( .A(n1530), .B(n1231), .Z(n3626) );
  XNOR U1107 ( .A(in[142]), .B(n3626), .Z(n4679) );
  XOR U1108 ( .A(in[815]), .B(in[495]), .Z(n673) );
  XNOR U1109 ( .A(in[1455]), .B(in[1135]), .Z(n672) );
  XNOR U1110 ( .A(n673), .B(n672), .Z(n674) );
  XOR U1111 ( .A(in[175]), .B(n674), .Z(n925) );
  XOR U1112 ( .A(in[1326]), .B(in[46]), .Z(n676) );
  XNOR U1113 ( .A(in[686]), .B(in[366]), .Z(n675) );
  XNOR U1114 ( .A(n676), .B(n675), .Z(n677) );
  XOR U1115 ( .A(in[1006]), .B(n677), .Z(n1336) );
  XNOR U1116 ( .A(n925), .B(n1336), .Z(n3992) );
  XNOR U1117 ( .A(in[1391]), .B(n3992), .Z(n4676) );
  NAND U1118 ( .A(n4679), .B(n4676), .Z(n678) );
  XNOR U1119 ( .A(n1441), .B(n678), .Z(out[1035]) );
  XNOR U1120 ( .A(n680), .B(n679), .Z(n3677) );
  XNOR U1121 ( .A(in[543]), .B(n3677), .Z(n1445) );
  XOR U1122 ( .A(in[78]), .B(in[1038]), .Z(n682) );
  XNOR U1123 ( .A(in[718]), .B(in[398]), .Z(n681) );
  XNOR U1124 ( .A(n682), .B(n681), .Z(n683) );
  XOR U1125 ( .A(in[1358]), .B(n683), .Z(n1534) );
  XOR U1126 ( .A(in[1487]), .B(in[527]), .Z(n685) );
  XNOR U1127 ( .A(in[847]), .B(in[207]), .Z(n684) );
  XNOR U1128 ( .A(n685), .B(n684), .Z(n686) );
  XNOR U1129 ( .A(in[1167]), .B(n686), .Z(n1234) );
  XNOR U1130 ( .A(n1534), .B(n1234), .Z(n3630) );
  XNOR U1131 ( .A(in[143]), .B(n3630), .Z(n4683) );
  XOR U1132 ( .A(in[1327]), .B(in[47]), .Z(n688) );
  XNOR U1133 ( .A(in[687]), .B(in[367]), .Z(n687) );
  XNOR U1134 ( .A(n688), .B(n687), .Z(n689) );
  XOR U1135 ( .A(in[1007]), .B(n689), .Z(n1340) );
  XOR U1136 ( .A(in[816]), .B(in[496]), .Z(n691) );
  XNOR U1137 ( .A(in[1456]), .B(in[1136]), .Z(n690) );
  XNOR U1138 ( .A(n691), .B(n690), .Z(n692) );
  XOR U1139 ( .A(in[176]), .B(n692), .Z(n940) );
  XNOR U1140 ( .A(n1340), .B(n940), .Z(n3995) );
  XNOR U1141 ( .A(in[1392]), .B(n3995), .Z(n4680) );
  NAND U1142 ( .A(n4683), .B(n4680), .Z(n693) );
  XNOR U1143 ( .A(n1445), .B(n693), .Z(out[1036]) );
  XNOR U1144 ( .A(n695), .B(n694), .Z(n3681) );
  XNOR U1145 ( .A(in[544]), .B(n3681), .Z(n1449) );
  XOR U1146 ( .A(in[79]), .B(in[1039]), .Z(n697) );
  XNOR U1147 ( .A(in[719]), .B(in[399]), .Z(n696) );
  XNOR U1148 ( .A(n697), .B(n696), .Z(n698) );
  XOR U1149 ( .A(in[1359]), .B(n698), .Z(n1538) );
  XOR U1150 ( .A(in[1488]), .B(in[528]), .Z(n700) );
  XNOR U1151 ( .A(in[848]), .B(in[208]), .Z(n699) );
  XNOR U1152 ( .A(n700), .B(n699), .Z(n701) );
  XNOR U1153 ( .A(in[1168]), .B(n701), .Z(n1237) );
  XNOR U1154 ( .A(n1538), .B(n1237), .Z(n3634) );
  XNOR U1155 ( .A(in[144]), .B(n3634), .Z(n4687) );
  XOR U1156 ( .A(in[817]), .B(in[497]), .Z(n703) );
  XNOR U1157 ( .A(in[1457]), .B(in[1137]), .Z(n702) );
  XNOR U1158 ( .A(n703), .B(n702), .Z(n704) );
  XOR U1159 ( .A(in[177]), .B(n704), .Z(n955) );
  XOR U1160 ( .A(in[1328]), .B(in[48]), .Z(n706) );
  XNOR U1161 ( .A(in[688]), .B(in[368]), .Z(n705) );
  XNOR U1162 ( .A(n706), .B(n705), .Z(n707) );
  XOR U1163 ( .A(in[1008]), .B(n707), .Z(n1344) );
  XNOR U1164 ( .A(n955), .B(n1344), .Z(n3998) );
  XNOR U1165 ( .A(in[1393]), .B(n3998), .Z(n4684) );
  NAND U1166 ( .A(n4687), .B(n4684), .Z(n708) );
  XNOR U1167 ( .A(n1449), .B(n708), .Z(out[1037]) );
  XNOR U1168 ( .A(n710), .B(n709), .Z(n3685) );
  XNOR U1169 ( .A(in[545]), .B(n3685), .Z(n1453) );
  XOR U1170 ( .A(in[80]), .B(in[1040]), .Z(n712) );
  XNOR U1171 ( .A(in[720]), .B(in[400]), .Z(n711) );
  XNOR U1172 ( .A(n712), .B(n711), .Z(n713) );
  XOR U1173 ( .A(in[1360]), .B(n713), .Z(n1542) );
  XOR U1174 ( .A(in[1489]), .B(in[529]), .Z(n715) );
  XNOR U1175 ( .A(in[849]), .B(in[209]), .Z(n714) );
  XNOR U1176 ( .A(n715), .B(n714), .Z(n716) );
  XNOR U1177 ( .A(in[1169]), .B(n716), .Z(n1240) );
  XNOR U1178 ( .A(n1542), .B(n1240), .Z(n3638) );
  XNOR U1179 ( .A(in[145]), .B(n3638), .Z(n4691) );
  XOR U1180 ( .A(in[1329]), .B(in[49]), .Z(n718) );
  XNOR U1181 ( .A(in[689]), .B(in[369]), .Z(n717) );
  XNOR U1182 ( .A(n718), .B(n717), .Z(n719) );
  XOR U1183 ( .A(in[1009]), .B(n719), .Z(n1349) );
  XOR U1184 ( .A(in[818]), .B(in[498]), .Z(n721) );
  XNOR U1185 ( .A(in[1458]), .B(in[1138]), .Z(n720) );
  XNOR U1186 ( .A(n721), .B(n720), .Z(n722) );
  XOR U1187 ( .A(in[178]), .B(n722), .Z(n970) );
  XNOR U1188 ( .A(n1349), .B(n970), .Z(n4001) );
  XNOR U1189 ( .A(in[1394]), .B(n4001), .Z(n4688) );
  NAND U1190 ( .A(n4691), .B(n4688), .Z(n723) );
  XNOR U1191 ( .A(n1453), .B(n723), .Z(out[1038]) );
  XOR U1192 ( .A(n3689), .B(in[546]), .Z(n1457) );
  XOR U1193 ( .A(in[81]), .B(in[1041]), .Z(n725) );
  XNOR U1194 ( .A(in[721]), .B(in[401]), .Z(n724) );
  XNOR U1195 ( .A(n725), .B(n724), .Z(n726) );
  XOR U1196 ( .A(in[1361]), .B(n726), .Z(n1546) );
  XOR U1197 ( .A(in[1490]), .B(in[530]), .Z(n728) );
  XNOR U1198 ( .A(in[850]), .B(in[210]), .Z(n727) );
  XNOR U1199 ( .A(n728), .B(n727), .Z(n729) );
  XNOR U1200 ( .A(in[1170]), .B(n729), .Z(n1244) );
  XNOR U1201 ( .A(n1546), .B(n1244), .Z(n3642) );
  XNOR U1202 ( .A(in[146]), .B(n3642), .Z(n4695) );
  XOR U1203 ( .A(in[819]), .B(in[499]), .Z(n731) );
  XNOR U1204 ( .A(in[1459]), .B(in[1139]), .Z(n730) );
  XNOR U1205 ( .A(n731), .B(n730), .Z(n732) );
  XOR U1206 ( .A(in[179]), .B(n732), .Z(n985) );
  XOR U1207 ( .A(in[1330]), .B(in[50]), .Z(n734) );
  XNOR U1208 ( .A(in[690]), .B(in[370]), .Z(n733) );
  XNOR U1209 ( .A(n734), .B(n733), .Z(n735) );
  XOR U1210 ( .A(in[1010]), .B(n735), .Z(n1353) );
  XNOR U1211 ( .A(n985), .B(n1353), .Z(n4008) );
  XNOR U1212 ( .A(in[1395]), .B(n4008), .Z(n4692) );
  NAND U1213 ( .A(n4695), .B(n4692), .Z(n736) );
  XNOR U1214 ( .A(n1457), .B(n736), .Z(out[1039]) );
  XOR U1215 ( .A(in[1342]), .B(in[62]), .Z(n738) );
  XNOR U1216 ( .A(in[702]), .B(in[382]), .Z(n737) );
  XNOR U1217 ( .A(n738), .B(n737), .Z(n739) );
  XOR U1218 ( .A(in[1022]), .B(n739), .Z(n907) );
  XNOR U1219 ( .A(n740), .B(n907), .Z(n3604) );
  XNOR U1220 ( .A(in[638]), .B(n3604), .Z(n2557) );
  XOR U1221 ( .A(n742), .B(n741), .Z(n3701) );
  XNOR U1222 ( .A(in[229]), .B(n3701), .Z(n2873) );
  XOR U1223 ( .A(in[1513]), .B(in[553]), .Z(n744) );
  XNOR U1224 ( .A(in[873]), .B(in[233]), .Z(n743) );
  XNOR U1225 ( .A(n744), .B(n743), .Z(n745) );
  XOR U1226 ( .A(in[1193]), .B(n745), .Z(n1320) );
  XNOR U1227 ( .A(n746), .B(n1320), .Z(n3742) );
  XNOR U1228 ( .A(in[1449]), .B(n3742), .Z(n2870) );
  NAND U1229 ( .A(n2873), .B(n2870), .Z(n747) );
  XNOR U1230 ( .A(n2557), .B(n747), .Z(out[103]) );
  XOR U1231 ( .A(n3693), .B(in[547]), .Z(n1461) );
  XOR U1232 ( .A(in[1042]), .B(in[402]), .Z(n749) );
  XNOR U1233 ( .A(in[722]), .B(in[82]), .Z(n748) );
  XNOR U1234 ( .A(n749), .B(n748), .Z(n750) );
  XOR U1235 ( .A(in[1362]), .B(n750), .Z(n1551) );
  XOR U1236 ( .A(in[851]), .B(in[1171]), .Z(n752) );
  XNOR U1237 ( .A(in[1491]), .B(in[211]), .Z(n751) );
  XNOR U1238 ( .A(n752), .B(n751), .Z(n753) );
  XNOR U1239 ( .A(in[531]), .B(n753), .Z(n1247) );
  XNOR U1240 ( .A(n1551), .B(n1247), .Z(n3646) );
  XNOR U1241 ( .A(in[147]), .B(n3646), .Z(n4699) );
  XOR U1242 ( .A(in[820]), .B(in[500]), .Z(n755) );
  XNOR U1243 ( .A(in[1460]), .B(in[1140]), .Z(n754) );
  XNOR U1244 ( .A(n755), .B(n754), .Z(n756) );
  XOR U1245 ( .A(in[180]), .B(n756), .Z(n1000) );
  XOR U1246 ( .A(in[1331]), .B(in[51]), .Z(n758) );
  XNOR U1247 ( .A(in[691]), .B(in[371]), .Z(n757) );
  XNOR U1248 ( .A(n758), .B(n757), .Z(n759) );
  XOR U1249 ( .A(in[1011]), .B(n759), .Z(n1357) );
  XNOR U1250 ( .A(n1000), .B(n1357), .Z(n4011) );
  XNOR U1251 ( .A(in[1396]), .B(n4011), .Z(n4696) );
  NAND U1252 ( .A(n4699), .B(n4696), .Z(n760) );
  XNOR U1253 ( .A(n1461), .B(n760), .Z(out[1040]) );
  XOR U1254 ( .A(n3697), .B(in[548]), .Z(n1465) );
  XOR U1255 ( .A(in[83]), .B(in[1043]), .Z(n762) );
  XNOR U1256 ( .A(in[723]), .B(in[403]), .Z(n761) );
  XNOR U1257 ( .A(n762), .B(n761), .Z(n763) );
  XOR U1258 ( .A(in[1363]), .B(n763), .Z(n1555) );
  XOR U1259 ( .A(in[852]), .B(in[1172]), .Z(n765) );
  XNOR U1260 ( .A(in[1492]), .B(in[212]), .Z(n764) );
  XNOR U1261 ( .A(n765), .B(n764), .Z(n766) );
  XNOR U1262 ( .A(in[532]), .B(n766), .Z(n1250) );
  XNOR U1263 ( .A(n1555), .B(n1250), .Z(n3650) );
  XNOR U1264 ( .A(in[148]), .B(n3650), .Z(n4703) );
  XOR U1265 ( .A(in[1332]), .B(in[52]), .Z(n768) );
  XNOR U1266 ( .A(in[692]), .B(in[372]), .Z(n767) );
  XNOR U1267 ( .A(n768), .B(n767), .Z(n769) );
  XOR U1268 ( .A(in[1012]), .B(n769), .Z(n1361) );
  XOR U1269 ( .A(in[821]), .B(in[501]), .Z(n771) );
  XNOR U1270 ( .A(in[1461]), .B(in[1141]), .Z(n770) );
  XNOR U1271 ( .A(n771), .B(n770), .Z(n772) );
  XOR U1272 ( .A(in[181]), .B(n772), .Z(n1015) );
  XNOR U1273 ( .A(n1361), .B(n1015), .Z(n4014) );
  XNOR U1274 ( .A(in[1397]), .B(n4014), .Z(n4700) );
  NAND U1275 ( .A(n4703), .B(n4700), .Z(n773) );
  XNOR U1276 ( .A(n1465), .B(n773), .Z(out[1041]) );
  XOR U1277 ( .A(n3701), .B(in[549]), .Z(n1470) );
  XOR U1278 ( .A(in[853]), .B(in[1173]), .Z(n775) );
  XNOR U1279 ( .A(in[1493]), .B(in[213]), .Z(n774) );
  XNOR U1280 ( .A(n775), .B(n774), .Z(n776) );
  XNOR U1281 ( .A(in[533]), .B(n776), .Z(n1253) );
  XNOR U1282 ( .A(n777), .B(n1253), .Z(n3654) );
  XNOR U1283 ( .A(in[149]), .B(n3654), .Z(n4707) );
  XOR U1284 ( .A(in[822]), .B(in[502]), .Z(n779) );
  XNOR U1285 ( .A(in[1462]), .B(in[1142]), .Z(n778) );
  XNOR U1286 ( .A(n779), .B(n778), .Z(n780) );
  XOR U1287 ( .A(in[182]), .B(n780), .Z(n1029) );
  XOR U1288 ( .A(in[1333]), .B(in[53]), .Z(n782) );
  XNOR U1289 ( .A(in[693]), .B(in[373]), .Z(n781) );
  XNOR U1290 ( .A(n782), .B(n781), .Z(n783) );
  XOR U1291 ( .A(in[1013]), .B(n783), .Z(n1365) );
  XNOR U1292 ( .A(n1029), .B(n1365), .Z(n4017) );
  XNOR U1293 ( .A(in[1398]), .B(n4017), .Z(n4704) );
  NAND U1294 ( .A(n4707), .B(n4704), .Z(n784) );
  XNOR U1295 ( .A(n1470), .B(n784), .Z(out[1042]) );
  XNOR U1296 ( .A(n786), .B(n785), .Z(n3705) );
  XNOR U1297 ( .A(in[550]), .B(n3705), .Z(n1474) );
  XOR U1298 ( .A(in[854]), .B(in[1174]), .Z(n788) );
  XNOR U1299 ( .A(in[1494]), .B(in[214]), .Z(n787) );
  XNOR U1300 ( .A(n788), .B(n787), .Z(n789) );
  XNOR U1301 ( .A(in[534]), .B(n789), .Z(n1256) );
  XNOR U1302 ( .A(n790), .B(n1256), .Z(n3658) );
  XNOR U1303 ( .A(in[150]), .B(n3658), .Z(n4711) );
  XOR U1304 ( .A(in[823]), .B(in[503]), .Z(n792) );
  XNOR U1305 ( .A(in[1463]), .B(in[1143]), .Z(n791) );
  XNOR U1306 ( .A(n792), .B(n791), .Z(n793) );
  XOR U1307 ( .A(in[183]), .B(n793), .Z(n1040) );
  XOR U1308 ( .A(in[1334]), .B(in[54]), .Z(n795) );
  XNOR U1309 ( .A(in[694]), .B(in[374]), .Z(n794) );
  XNOR U1310 ( .A(n795), .B(n794), .Z(n796) );
  XOR U1311 ( .A(in[1014]), .B(n796), .Z(n1369) );
  XNOR U1312 ( .A(n1040), .B(n1369), .Z(n4020) );
  XNOR U1313 ( .A(in[1399]), .B(n4020), .Z(n4708) );
  NAND U1314 ( .A(n4711), .B(n4708), .Z(n797) );
  XNOR U1315 ( .A(n1474), .B(n797), .Z(out[1043]) );
  XNOR U1316 ( .A(n799), .B(n798), .Z(n3713) );
  XNOR U1317 ( .A(in[551]), .B(n3713), .Z(n1478) );
  XOR U1318 ( .A(in[855]), .B(in[1175]), .Z(n801) );
  XNOR U1319 ( .A(in[1495]), .B(in[215]), .Z(n800) );
  XNOR U1320 ( .A(n801), .B(n800), .Z(n802) );
  XNOR U1321 ( .A(in[535]), .B(n802), .Z(n1259) );
  XNOR U1322 ( .A(n803), .B(n1259), .Z(n3662) );
  XNOR U1323 ( .A(in[151]), .B(n3662), .Z(n4719) );
  XOR U1324 ( .A(in[824]), .B(in[504]), .Z(n805) );
  XNOR U1325 ( .A(in[1464]), .B(in[1144]), .Z(n804) );
  XNOR U1326 ( .A(n805), .B(n804), .Z(n806) );
  XOR U1327 ( .A(in[184]), .B(n806), .Z(n1045) );
  XOR U1328 ( .A(in[1335]), .B(in[55]), .Z(n808) );
  XNOR U1329 ( .A(in[695]), .B(in[375]), .Z(n807) );
  XNOR U1330 ( .A(n808), .B(n807), .Z(n809) );
  XOR U1331 ( .A(in[1015]), .B(n809), .Z(n1373) );
  XNOR U1332 ( .A(n1045), .B(n1373), .Z(n4023) );
  XNOR U1333 ( .A(in[1400]), .B(n4023), .Z(n4716) );
  NAND U1334 ( .A(n4719), .B(n4716), .Z(n810) );
  XNOR U1335 ( .A(n1478), .B(n810), .Z(out[1044]) );
  XNOR U1336 ( .A(n812), .B(n811), .Z(n3717) );
  XNOR U1337 ( .A(in[552]), .B(n3717), .Z(n1482) );
  XOR U1338 ( .A(in[856]), .B(in[1176]), .Z(n814) );
  XNOR U1339 ( .A(in[1496]), .B(in[216]), .Z(n813) );
  XNOR U1340 ( .A(n814), .B(n813), .Z(n815) );
  XNOR U1341 ( .A(in[536]), .B(n815), .Z(n1262) );
  XNOR U1342 ( .A(n816), .B(n1262), .Z(n3670) );
  XNOR U1343 ( .A(in[152]), .B(n3670), .Z(n4723) );
  XOR U1344 ( .A(in[1336]), .B(in[56]), .Z(n818) );
  XNOR U1345 ( .A(in[696]), .B(in[376]), .Z(n817) );
  XNOR U1346 ( .A(n818), .B(n817), .Z(n819) );
  XOR U1347 ( .A(in[1016]), .B(n819), .Z(n1377) );
  XOR U1348 ( .A(in[825]), .B(in[505]), .Z(n821) );
  XNOR U1349 ( .A(in[1465]), .B(in[1145]), .Z(n820) );
  XNOR U1350 ( .A(n821), .B(n820), .Z(n822) );
  XOR U1351 ( .A(in[185]), .B(n822), .Z(n1056) );
  XNOR U1352 ( .A(n1377), .B(n1056), .Z(n4026) );
  XNOR U1353 ( .A(in[1401]), .B(n4026), .Z(n4720) );
  NAND U1354 ( .A(n4723), .B(n4720), .Z(n823) );
  XNOR U1355 ( .A(n1482), .B(n823), .Z(out[1045]) );
  XNOR U1356 ( .A(n825), .B(n824), .Z(n3721) );
  XNOR U1357 ( .A(in[553]), .B(n3721), .Z(n1486) );
  XOR U1358 ( .A(in[857]), .B(in[1177]), .Z(n827) );
  XNOR U1359 ( .A(in[1497]), .B(in[217]), .Z(n826) );
  XNOR U1360 ( .A(n827), .B(n826), .Z(n828) );
  XNOR U1361 ( .A(in[537]), .B(n828), .Z(n1265) );
  XNOR U1362 ( .A(n829), .B(n1265), .Z(n3674) );
  XNOR U1363 ( .A(in[153]), .B(n3674), .Z(n4727) );
  XOR U1364 ( .A(in[1337]), .B(in[57]), .Z(n831) );
  XNOR U1365 ( .A(in[697]), .B(in[377]), .Z(n830) );
  XNOR U1366 ( .A(n831), .B(n830), .Z(n832) );
  XOR U1367 ( .A(in[1017]), .B(n832), .Z(n1381) );
  XOR U1368 ( .A(in[826]), .B(in[506]), .Z(n834) );
  XNOR U1369 ( .A(in[1466]), .B(in[1146]), .Z(n833) );
  XNOR U1370 ( .A(n834), .B(n833), .Z(n835) );
  XOR U1371 ( .A(in[186]), .B(n835), .Z(n1067) );
  XNOR U1372 ( .A(n1381), .B(n1067), .Z(n4029) );
  XNOR U1373 ( .A(in[1402]), .B(n4029), .Z(n4724) );
  NAND U1374 ( .A(n4727), .B(n4724), .Z(n836) );
  XNOR U1375 ( .A(n1486), .B(n836), .Z(out[1046]) );
  XNOR U1376 ( .A(n838), .B(n837), .Z(n3725) );
  XNOR U1377 ( .A(in[554]), .B(n3725), .Z(n1490) );
  XOR U1378 ( .A(in[858]), .B(in[1178]), .Z(n840) );
  XNOR U1379 ( .A(in[1498]), .B(in[218]), .Z(n839) );
  XNOR U1380 ( .A(n840), .B(n839), .Z(n841) );
  XNOR U1381 ( .A(in[538]), .B(n841), .Z(n1268) );
  XNOR U1382 ( .A(n842), .B(n1268), .Z(n3678) );
  XNOR U1383 ( .A(in[154]), .B(n3678), .Z(n4731) );
  XOR U1384 ( .A(in[1338]), .B(in[58]), .Z(n844) );
  XNOR U1385 ( .A(in[698]), .B(in[378]), .Z(n843) );
  XNOR U1386 ( .A(n844), .B(n843), .Z(n845) );
  XOR U1387 ( .A(in[1018]), .B(n845), .Z(n1385) );
  XOR U1388 ( .A(in[827]), .B(in[507]), .Z(n847) );
  XNOR U1389 ( .A(in[1467]), .B(in[1147]), .Z(n846) );
  XNOR U1390 ( .A(n847), .B(n846), .Z(n848) );
  XOR U1391 ( .A(in[187]), .B(n848), .Z(n1072) );
  XNOR U1392 ( .A(n1385), .B(n1072), .Z(n4032) );
  XNOR U1393 ( .A(in[1403]), .B(n4032), .Z(n4728) );
  NAND U1394 ( .A(n4731), .B(n4728), .Z(n849) );
  XNOR U1395 ( .A(n1490), .B(n849), .Z(out[1047]) );
  XOR U1396 ( .A(in[1579]), .B(in[619]), .Z(n851) );
  XNOR U1397 ( .A(in[939]), .B(in[299]), .Z(n850) );
  XNOR U1398 ( .A(n851), .B(n850), .Z(n852) );
  XOR U1399 ( .A(in[1259]), .B(n852), .Z(n1394) );
  XNOR U1400 ( .A(n853), .B(n1394), .Z(n3729) );
  XNOR U1401 ( .A(in[555]), .B(n3729), .Z(n1494) );
  XOR U1402 ( .A(in[859]), .B(in[1179]), .Z(n855) );
  XNOR U1403 ( .A(in[1499]), .B(in[219]), .Z(n854) );
  XNOR U1404 ( .A(n855), .B(n854), .Z(n856) );
  XNOR U1405 ( .A(in[539]), .B(n856), .Z(n1271) );
  XNOR U1406 ( .A(n857), .B(n1271), .Z(n3682) );
  XNOR U1407 ( .A(in[155]), .B(n3682), .Z(n4735) );
  XOR U1408 ( .A(in[828]), .B(in[508]), .Z(n859) );
  XNOR U1409 ( .A(in[1468]), .B(in[1148]), .Z(n858) );
  XNOR U1410 ( .A(n859), .B(n858), .Z(n860) );
  XOR U1411 ( .A(in[188]), .B(n860), .Z(n1077) );
  XNOR U1412 ( .A(n861), .B(n1077), .Z(n4035) );
  XNOR U1413 ( .A(in[1404]), .B(n4035), .Z(n4732) );
  NAND U1414 ( .A(n4735), .B(n4732), .Z(n862) );
  XNOR U1415 ( .A(n1494), .B(n862), .Z(out[1048]) );
  XOR U1416 ( .A(in[1580]), .B(in[620]), .Z(n864) );
  XNOR U1417 ( .A(in[940]), .B(in[300]), .Z(n863) );
  XNOR U1418 ( .A(n864), .B(n863), .Z(n865) );
  XOR U1419 ( .A(in[1260]), .B(n865), .Z(n1398) );
  XNOR U1420 ( .A(n866), .B(n1398), .Z(n3733) );
  XNOR U1421 ( .A(in[556]), .B(n3733), .Z(n1498) );
  XOR U1422 ( .A(in[860]), .B(in[1180]), .Z(n868) );
  XNOR U1423 ( .A(in[1500]), .B(in[220]), .Z(n867) );
  XNOR U1424 ( .A(n868), .B(n867), .Z(n869) );
  XNOR U1425 ( .A(in[540]), .B(n869), .Z(n1275) );
  XNOR U1426 ( .A(n870), .B(n1275), .Z(n3686) );
  XNOR U1427 ( .A(in[156]), .B(n3686), .Z(n4739) );
  XNOR U1428 ( .A(n872), .B(n871), .Z(n4042) );
  XNOR U1429 ( .A(in[1405]), .B(n4042), .Z(n4736) );
  NAND U1430 ( .A(n4739), .B(n4736), .Z(n873) );
  XNOR U1431 ( .A(n1498), .B(n873), .Z(out[1049]) );
  XOR U1432 ( .A(in[1343]), .B(in[63]), .Z(n875) );
  XNOR U1433 ( .A(in[703]), .B(in[383]), .Z(n874) );
  XNOR U1434 ( .A(n875), .B(n874), .Z(n876) );
  XOR U1435 ( .A(in[1023]), .B(n876), .Z(n920) );
  XNOR U1436 ( .A(n877), .B(n920), .Z(n3608) );
  XNOR U1437 ( .A(in[639]), .B(n3608), .Z(n2559) );
  XOR U1438 ( .A(in[230]), .B(n3705), .Z(n2889) );
  XOR U1439 ( .A(in[874]), .B(in[1194]), .Z(n879) );
  XNOR U1440 ( .A(in[1514]), .B(in[234]), .Z(n878) );
  XNOR U1441 ( .A(n879), .B(n878), .Z(n880) );
  XOR U1442 ( .A(in[554]), .B(n880), .Z(n1324) );
  XNOR U1443 ( .A(n881), .B(n1324), .Z(n3746) );
  XNOR U1444 ( .A(in[1450]), .B(n3746), .Z(n2886) );
  NAND U1445 ( .A(n2889), .B(n2886), .Z(n882) );
  XNOR U1446 ( .A(n2559), .B(n882), .Z(out[104]) );
  XOR U1447 ( .A(in[1581]), .B(in[621]), .Z(n884) );
  XNOR U1448 ( .A(in[941]), .B(in[301]), .Z(n883) );
  XNOR U1449 ( .A(n884), .B(n883), .Z(n885) );
  XOR U1450 ( .A(in[1261]), .B(n885), .Z(n1402) );
  XNOR U1451 ( .A(n886), .B(n1402), .Z(n3737) );
  XNOR U1452 ( .A(in[557]), .B(n3737), .Z(n1502) );
  XOR U1453 ( .A(in[861]), .B(in[1181]), .Z(n888) );
  XNOR U1454 ( .A(in[1501]), .B(in[221]), .Z(n887) );
  XNOR U1455 ( .A(n888), .B(n887), .Z(n889) );
  XNOR U1456 ( .A(in[541]), .B(n889), .Z(n1278) );
  XNOR U1457 ( .A(n890), .B(n1278), .Z(n3690) );
  XNOR U1458 ( .A(in[157]), .B(n3690), .Z(n4743) );
  XOR U1459 ( .A(in[830]), .B(in[510]), .Z(n892) );
  XNOR U1460 ( .A(in[1470]), .B(in[1150]), .Z(n891) );
  XNOR U1461 ( .A(n892), .B(n891), .Z(n893) );
  XOR U1462 ( .A(in[190]), .B(n893), .Z(n1083) );
  XNOR U1463 ( .A(n894), .B(n1083), .Z(n4045) );
  XNOR U1464 ( .A(in[1406]), .B(n4045), .Z(n4740) );
  NAND U1465 ( .A(n4743), .B(n4740), .Z(n895) );
  XNOR U1466 ( .A(n1502), .B(n895), .Z(out[1050]) );
  XOR U1467 ( .A(in[1582]), .B(in[622]), .Z(n897) );
  XNOR U1468 ( .A(in[942]), .B(in[302]), .Z(n896) );
  XNOR U1469 ( .A(n897), .B(n896), .Z(n898) );
  XOR U1470 ( .A(in[1262]), .B(n898), .Z(n1406) );
  XNOR U1471 ( .A(n899), .B(n1406), .Z(n3741) );
  XNOR U1472 ( .A(in[558]), .B(n3741), .Z(n1506) );
  XOR U1473 ( .A(in[862]), .B(in[1182]), .Z(n901) );
  XNOR U1474 ( .A(in[1502]), .B(in[222]), .Z(n900) );
  XNOR U1475 ( .A(n901), .B(n900), .Z(n902) );
  XNOR U1476 ( .A(in[542]), .B(n902), .Z(n1281) );
  XNOR U1477 ( .A(n903), .B(n1281), .Z(n3694) );
  XNOR U1478 ( .A(in[158]), .B(n3694), .Z(n4747) );
  XOR U1479 ( .A(in[831]), .B(in[511]), .Z(n905) );
  XNOR U1480 ( .A(in[1471]), .B(in[1151]), .Z(n904) );
  XNOR U1481 ( .A(n905), .B(n904), .Z(n906) );
  XOR U1482 ( .A(in[191]), .B(n906), .Z(n1088) );
  XNOR U1483 ( .A(n907), .B(n1088), .Z(n4048) );
  XNOR U1484 ( .A(in[1407]), .B(n4048), .Z(n4744) );
  NAND U1485 ( .A(n4747), .B(n4744), .Z(n908) );
  XNOR U1486 ( .A(n1506), .B(n908), .Z(out[1051]) );
  XOR U1487 ( .A(in[1583]), .B(in[623]), .Z(n910) );
  XNOR U1488 ( .A(in[943]), .B(in[303]), .Z(n909) );
  XNOR U1489 ( .A(n910), .B(n909), .Z(n911) );
  XOR U1490 ( .A(in[1263]), .B(n911), .Z(n1410) );
  XNOR U1491 ( .A(n912), .B(n1410), .Z(n3745) );
  XNOR U1492 ( .A(in[559]), .B(n3745), .Z(n1511) );
  XOR U1493 ( .A(in[863]), .B(in[1183]), .Z(n914) );
  XNOR U1494 ( .A(in[1503]), .B(in[223]), .Z(n913) );
  XNOR U1495 ( .A(n914), .B(n913), .Z(n915) );
  XNOR U1496 ( .A(in[543]), .B(n915), .Z(n1284) );
  XNOR U1497 ( .A(n916), .B(n1284), .Z(n3698) );
  XNOR U1498 ( .A(in[159]), .B(n3698), .Z(n4751) );
  XOR U1499 ( .A(in[768]), .B(in[1088]), .Z(n918) );
  XNOR U1500 ( .A(in[448]), .B(in[1408]), .Z(n917) );
  XNOR U1501 ( .A(n918), .B(n917), .Z(n919) );
  XOR U1502 ( .A(in[128]), .B(n919), .Z(n1096) );
  XNOR U1503 ( .A(n920), .B(n1096), .Z(n4051) );
  XNOR U1504 ( .A(in[1344]), .B(n4051), .Z(n4748) );
  NAND U1505 ( .A(n4751), .B(n4748), .Z(n921) );
  XNOR U1506 ( .A(n1511), .B(n921), .Z(out[1052]) );
  XOR U1507 ( .A(in[1584]), .B(in[624]), .Z(n923) );
  XNOR U1508 ( .A(in[944]), .B(in[304]), .Z(n922) );
  XNOR U1509 ( .A(n923), .B(n922), .Z(n924) );
  XOR U1510 ( .A(in[1264]), .B(n924), .Z(n1414) );
  XNOR U1511 ( .A(n925), .B(n1414), .Z(n3749) );
  XNOR U1512 ( .A(in[560]), .B(n3749), .Z(n1515) );
  XOR U1513 ( .A(in[224]), .B(in[864]), .Z(n927) );
  XNOR U1514 ( .A(in[1184]), .B(in[1504]), .Z(n926) );
  XNOR U1515 ( .A(n927), .B(n926), .Z(n928) );
  XNOR U1516 ( .A(in[544]), .B(n928), .Z(n1287) );
  XNOR U1517 ( .A(n929), .B(n1287), .Z(n3702) );
  XNOR U1518 ( .A(in[160]), .B(n3702), .Z(n4755) );
  XOR U1519 ( .A(in[1280]), .B(in[640]), .Z(n931) );
  XNOR U1520 ( .A(in[960]), .B(in[320]), .Z(n930) );
  XNOR U1521 ( .A(n931), .B(n930), .Z(n932) );
  XOR U1522 ( .A(in[0]), .B(n932), .Z(n1023) );
  XOR U1523 ( .A(in[769]), .B(in[1089]), .Z(n934) );
  XNOR U1524 ( .A(in[449]), .B(in[1409]), .Z(n933) );
  XNOR U1525 ( .A(n934), .B(n933), .Z(n935) );
  XOR U1526 ( .A(in[129]), .B(n935), .Z(n1101) );
  XNOR U1527 ( .A(n1023), .B(n1101), .Z(n4054) );
  XNOR U1528 ( .A(in[1345]), .B(n4054), .Z(n4752) );
  NAND U1529 ( .A(n4755), .B(n4752), .Z(n936) );
  XNOR U1530 ( .A(n1515), .B(n936), .Z(out[1053]) );
  XOR U1531 ( .A(in[1585]), .B(in[625]), .Z(n938) );
  XNOR U1532 ( .A(in[945]), .B(in[305]), .Z(n937) );
  XNOR U1533 ( .A(n938), .B(n937), .Z(n939) );
  XOR U1534 ( .A(in[1265]), .B(n939), .Z(n1418) );
  XNOR U1535 ( .A(n940), .B(n1418), .Z(n3757) );
  XNOR U1536 ( .A(in[561]), .B(n3757), .Z(n1519) );
  XOR U1537 ( .A(in[225]), .B(in[865]), .Z(n942) );
  XNOR U1538 ( .A(in[1185]), .B(in[1505]), .Z(n941) );
  XNOR U1539 ( .A(n942), .B(n941), .Z(n943) );
  XNOR U1540 ( .A(in[545]), .B(n943), .Z(n1290) );
  XNOR U1541 ( .A(n944), .B(n1290), .Z(n3706) );
  XNOR U1542 ( .A(in[161]), .B(n3706), .Z(n4763) );
  XOR U1543 ( .A(in[1]), .B(in[641]), .Z(n946) );
  XNOR U1544 ( .A(in[961]), .B(in[321]), .Z(n945) );
  XNOR U1545 ( .A(n946), .B(n945), .Z(n947) );
  XOR U1546 ( .A(in[1281]), .B(n947), .Z(n1090) );
  XOR U1547 ( .A(in[1090]), .B(in[450]), .Z(n949) );
  XNOR U1548 ( .A(in[130]), .B(in[770]), .Z(n948) );
  XNOR U1549 ( .A(n949), .B(n948), .Z(n950) );
  XOR U1550 ( .A(in[1410]), .B(n950), .Z(n1106) );
  XNOR U1551 ( .A(n1090), .B(n1106), .Z(n4057) );
  XNOR U1552 ( .A(in[1346]), .B(n4057), .Z(n4760) );
  NAND U1553 ( .A(n4763), .B(n4760), .Z(n951) );
  XNOR U1554 ( .A(n1519), .B(n951), .Z(out[1054]) );
  XOR U1555 ( .A(in[1586]), .B(in[626]), .Z(n953) );
  XNOR U1556 ( .A(in[946]), .B(in[306]), .Z(n952) );
  XNOR U1557 ( .A(n953), .B(n952), .Z(n954) );
  XOR U1558 ( .A(in[1266]), .B(n954), .Z(n1422) );
  XNOR U1559 ( .A(n955), .B(n1422), .Z(n3761) );
  XNOR U1560 ( .A(in[562]), .B(n3761), .Z(n1523) );
  XOR U1561 ( .A(in[1186]), .B(in[1506]), .Z(n957) );
  XNOR U1562 ( .A(in[546]), .B(in[866]), .Z(n956) );
  XNOR U1563 ( .A(n957), .B(n956), .Z(n958) );
  XNOR U1564 ( .A(in[226]), .B(n958), .Z(n1293) );
  XNOR U1565 ( .A(n959), .B(n1293), .Z(n3714) );
  XNOR U1566 ( .A(in[162]), .B(n3714), .Z(n4767) );
  XOR U1567 ( .A(in[771]), .B(in[1091]), .Z(n961) );
  XNOR U1568 ( .A(in[451]), .B(in[1411]), .Z(n960) );
  XNOR U1569 ( .A(n961), .B(n960), .Z(n962) );
  XOR U1570 ( .A(in[131]), .B(n962), .Z(n1111) );
  XOR U1571 ( .A(in[2]), .B(in[642]), .Z(n964) );
  XNOR U1572 ( .A(in[962]), .B(in[322]), .Z(n963) );
  XNOR U1573 ( .A(n964), .B(n963), .Z(n965) );
  XOR U1574 ( .A(in[1282]), .B(n965), .Z(n1143) );
  XNOR U1575 ( .A(n1111), .B(n1143), .Z(n4060) );
  XNOR U1576 ( .A(in[1347]), .B(n4060), .Z(n4764) );
  NAND U1577 ( .A(n4767), .B(n4764), .Z(n966) );
  XNOR U1578 ( .A(n1523), .B(n966), .Z(out[1055]) );
  XOR U1579 ( .A(in[1587]), .B(in[627]), .Z(n968) );
  XNOR U1580 ( .A(in[947]), .B(in[307]), .Z(n967) );
  XNOR U1581 ( .A(n968), .B(n967), .Z(n969) );
  XOR U1582 ( .A(in[1267]), .B(n969), .Z(n1427) );
  XNOR U1583 ( .A(n970), .B(n1427), .Z(n3765) );
  XNOR U1584 ( .A(in[563]), .B(n3765), .Z(n1527) );
  XOR U1585 ( .A(in[1187]), .B(in[1507]), .Z(n972) );
  XNOR U1586 ( .A(in[547]), .B(in[867]), .Z(n971) );
  XNOR U1587 ( .A(n972), .B(n971), .Z(n973) );
  XNOR U1588 ( .A(in[227]), .B(n973), .Z(n1296) );
  XNOR U1589 ( .A(n974), .B(n1296), .Z(n3718) );
  XNOR U1590 ( .A(in[163]), .B(n3718), .Z(n4771) );
  XOR U1591 ( .A(in[323]), .B(in[643]), .Z(n976) );
  XNOR U1592 ( .A(in[963]), .B(in[3]), .Z(n975) );
  XNOR U1593 ( .A(n976), .B(n975), .Z(n977) );
  XOR U1594 ( .A(in[1283]), .B(n977), .Z(n1189) );
  XOR U1595 ( .A(in[772]), .B(in[1092]), .Z(n979) );
  XNOR U1596 ( .A(in[452]), .B(in[1412]), .Z(n978) );
  XNOR U1597 ( .A(n979), .B(n978), .Z(n980) );
  XOR U1598 ( .A(in[132]), .B(n980), .Z(n1116) );
  XNOR U1599 ( .A(n1189), .B(n1116), .Z(n4063) );
  XNOR U1600 ( .A(in[1348]), .B(n4063), .Z(n4768) );
  NAND U1601 ( .A(n4771), .B(n4768), .Z(n981) );
  XNOR U1602 ( .A(n1527), .B(n981), .Z(out[1056]) );
  XOR U1603 ( .A(in[1588]), .B(in[628]), .Z(n983) );
  XNOR U1604 ( .A(in[948]), .B(in[308]), .Z(n982) );
  XNOR U1605 ( .A(n983), .B(n982), .Z(n984) );
  XOR U1606 ( .A(in[1268]), .B(n984), .Z(n1431) );
  XNOR U1607 ( .A(n985), .B(n1431), .Z(n3769) );
  XNOR U1608 ( .A(in[564]), .B(n3769), .Z(n1531) );
  XOR U1609 ( .A(in[1188]), .B(in[1508]), .Z(n987) );
  XNOR U1610 ( .A(in[548]), .B(in[868]), .Z(n986) );
  XNOR U1611 ( .A(n987), .B(n986), .Z(n988) );
  XOR U1612 ( .A(in[228]), .B(n988), .Z(n1299) );
  XNOR U1613 ( .A(n1299), .B(n989), .Z(n3722) );
  XNOR U1614 ( .A(in[164]), .B(n3722), .Z(n4775) );
  XOR U1615 ( .A(in[324]), .B(in[644]), .Z(n991) );
  XNOR U1616 ( .A(in[964]), .B(in[4]), .Z(n990) );
  XNOR U1617 ( .A(n991), .B(n990), .Z(n992) );
  XOR U1618 ( .A(in[1284]), .B(n992), .Z(n1197) );
  XOR U1619 ( .A(in[773]), .B(in[1093]), .Z(n994) );
  XNOR U1620 ( .A(in[453]), .B(in[1413]), .Z(n993) );
  XNOR U1621 ( .A(n994), .B(n993), .Z(n995) );
  XOR U1622 ( .A(in[133]), .B(n995), .Z(n1121) );
  XNOR U1623 ( .A(n1197), .B(n1121), .Z(n4066) );
  XNOR U1624 ( .A(in[1349]), .B(n4066), .Z(n4772) );
  NAND U1625 ( .A(n4775), .B(n4772), .Z(n996) );
  XNOR U1626 ( .A(n1531), .B(n996), .Z(out[1057]) );
  XOR U1627 ( .A(in[1589]), .B(in[629]), .Z(n998) );
  XNOR U1628 ( .A(in[949]), .B(in[309]), .Z(n997) );
  XNOR U1629 ( .A(n998), .B(n997), .Z(n999) );
  XOR U1630 ( .A(in[1269]), .B(n999), .Z(n1435) );
  XNOR U1631 ( .A(n1000), .B(n1435), .Z(n3773) );
  XNOR U1632 ( .A(in[565]), .B(n3773), .Z(n1535) );
  XOR U1633 ( .A(in[1189]), .B(in[1509]), .Z(n1002) );
  XNOR U1634 ( .A(in[549]), .B(in[869]), .Z(n1001) );
  XNOR U1635 ( .A(n1002), .B(n1001), .Z(n1003) );
  XNOR U1636 ( .A(in[229]), .B(n1003), .Z(n1303) );
  XNOR U1637 ( .A(n1004), .B(n1303), .Z(n3726) );
  XNOR U1638 ( .A(in[165]), .B(n3726), .Z(n4779) );
  XOR U1639 ( .A(in[774]), .B(in[1094]), .Z(n1006) );
  XNOR U1640 ( .A(in[454]), .B(in[1414]), .Z(n1005) );
  XNOR U1641 ( .A(n1006), .B(n1005), .Z(n1007) );
  XOR U1642 ( .A(in[134]), .B(n1007), .Z(n1126) );
  XOR U1643 ( .A(in[325]), .B(in[645]), .Z(n1009) );
  XNOR U1644 ( .A(in[965]), .B(in[5]), .Z(n1008) );
  XNOR U1645 ( .A(n1009), .B(n1008), .Z(n1010) );
  XOR U1646 ( .A(in[1285]), .B(n1010), .Z(n1200) );
  XNOR U1647 ( .A(n1126), .B(n1200), .Z(n4069) );
  XNOR U1648 ( .A(in[1350]), .B(n4069), .Z(n4776) );
  NAND U1649 ( .A(n4779), .B(n4776), .Z(n1011) );
  XNOR U1650 ( .A(n1535), .B(n1011), .Z(out[1058]) );
  XOR U1651 ( .A(in[1590]), .B(in[630]), .Z(n1013) );
  XNOR U1652 ( .A(in[950]), .B(in[310]), .Z(n1012) );
  XNOR U1653 ( .A(n1013), .B(n1012), .Z(n1014) );
  XOR U1654 ( .A(in[1270]), .B(n1014), .Z(n1439) );
  XNOR U1655 ( .A(n1015), .B(n1439), .Z(n3777) );
  XNOR U1656 ( .A(in[566]), .B(n3777), .Z(n1539) );
  XOR U1657 ( .A(in[166]), .B(n3730), .Z(n4783) );
  XOR U1658 ( .A(in[326]), .B(in[6]), .Z(n1017) );
  XNOR U1659 ( .A(in[966]), .B(in[646]), .Z(n1016) );
  XNOR U1660 ( .A(n1017), .B(n1016), .Z(n1018) );
  XOR U1661 ( .A(in[1286]), .B(n1018), .Z(n1203) );
  XOR U1662 ( .A(in[775]), .B(in[1095]), .Z(n1020) );
  XNOR U1663 ( .A(in[455]), .B(in[1415]), .Z(n1019) );
  XNOR U1664 ( .A(n1020), .B(n1019), .Z(n1021) );
  XOR U1665 ( .A(in[135]), .B(n1021), .Z(n1131) );
  XNOR U1666 ( .A(n1203), .B(n1131), .Z(n4080) );
  XNOR U1667 ( .A(in[1351]), .B(n4080), .Z(n4780) );
  NAND U1668 ( .A(n4783), .B(n4780), .Z(n1022) );
  XNOR U1669 ( .A(n1539), .B(n1022), .Z(out[1059]) );
  XNOR U1670 ( .A(n1024), .B(n1023), .Z(n3612) );
  XNOR U1671 ( .A(in[576]), .B(n3612), .Z(n2561) );
  XOR U1672 ( .A(in[231]), .B(n3713), .Z(n2903) );
  XNOR U1673 ( .A(in[1451]), .B(n3750), .Z(n2900) );
  NAND U1674 ( .A(n2903), .B(n2900), .Z(n1025) );
  XNOR U1675 ( .A(n2561), .B(n1025), .Z(out[105]) );
  XOR U1676 ( .A(in[1591]), .B(in[631]), .Z(n1027) );
  XNOR U1677 ( .A(in[951]), .B(in[311]), .Z(n1026) );
  XNOR U1678 ( .A(n1027), .B(n1026), .Z(n1028) );
  XOR U1679 ( .A(in[1271]), .B(n1028), .Z(n1443) );
  XNOR U1680 ( .A(n1029), .B(n1443), .Z(n3781) );
  XNOR U1681 ( .A(in[567]), .B(n3781), .Z(n1543) );
  XOR U1682 ( .A(in[167]), .B(n3734), .Z(n4787) );
  XOR U1683 ( .A(in[776]), .B(in[1096]), .Z(n1031) );
  XNOR U1684 ( .A(in[456]), .B(in[1416]), .Z(n1030) );
  XNOR U1685 ( .A(n1031), .B(n1030), .Z(n1032) );
  XOR U1686 ( .A(in[136]), .B(n1032), .Z(n1136) );
  XOR U1687 ( .A(in[327]), .B(in[7]), .Z(n1034) );
  XNOR U1688 ( .A(in[967]), .B(in[647]), .Z(n1033) );
  XNOR U1689 ( .A(n1034), .B(n1033), .Z(n1035) );
  XOR U1690 ( .A(in[1287]), .B(n1035), .Z(n1206) );
  XNOR U1691 ( .A(n1136), .B(n1206), .Z(n4083) );
  XNOR U1692 ( .A(in[1352]), .B(n4083), .Z(n4784) );
  NAND U1693 ( .A(n4787), .B(n4784), .Z(n1036) );
  XNOR U1694 ( .A(n1543), .B(n1036), .Z(out[1060]) );
  XOR U1695 ( .A(in[632]), .B(in[1592]), .Z(n1038) );
  XNOR U1696 ( .A(in[1272]), .B(in[312]), .Z(n1037) );
  XNOR U1697 ( .A(n1038), .B(n1037), .Z(n1039) );
  XOR U1698 ( .A(in[952]), .B(n1039), .Z(n1447) );
  XNOR U1699 ( .A(n1040), .B(n1447), .Z(n3785) );
  XNOR U1700 ( .A(in[568]), .B(n3785), .Z(n1547) );
  XOR U1701 ( .A(in[168]), .B(n3738), .Z(n4791) );
  XNOR U1702 ( .A(in[1353]), .B(n4086), .Z(n4788) );
  NAND U1703 ( .A(n4791), .B(n4788), .Z(n1041) );
  XNOR U1704 ( .A(n1547), .B(n1041), .Z(out[1061]) );
  XOR U1705 ( .A(in[633]), .B(in[1593]), .Z(n1043) );
  XNOR U1706 ( .A(in[1273]), .B(in[313]), .Z(n1042) );
  XNOR U1707 ( .A(n1043), .B(n1042), .Z(n1044) );
  XOR U1708 ( .A(in[953]), .B(n1044), .Z(n1451) );
  XNOR U1709 ( .A(n1045), .B(n1451), .Z(n3789) );
  XNOR U1710 ( .A(in[569]), .B(n3789), .Z(n1552) );
  XOR U1711 ( .A(in[169]), .B(n3742), .Z(n4795) );
  XOR U1712 ( .A(in[329]), .B(in[969]), .Z(n1047) );
  XNOR U1713 ( .A(in[9]), .B(in[649]), .Z(n1046) );
  XNOR U1714 ( .A(n1047), .B(n1046), .Z(n1048) );
  XOR U1715 ( .A(in[1289]), .B(n1048), .Z(n1214) );
  XOR U1716 ( .A(in[778]), .B(in[1098]), .Z(n1050) );
  XNOR U1717 ( .A(in[458]), .B(in[1418]), .Z(n1049) );
  XNOR U1718 ( .A(n1050), .B(n1049), .Z(n1051) );
  XOR U1719 ( .A(in[138]), .B(n1051), .Z(n1149) );
  XNOR U1720 ( .A(n1214), .B(n1149), .Z(n4089) );
  XNOR U1721 ( .A(in[1354]), .B(n4089), .Z(n4792) );
  NAND U1722 ( .A(n4795), .B(n4792), .Z(n1052) );
  XNOR U1723 ( .A(n1552), .B(n1052), .Z(out[1062]) );
  XOR U1724 ( .A(in[634]), .B(in[1594]), .Z(n1054) );
  XNOR U1725 ( .A(in[1274]), .B(in[314]), .Z(n1053) );
  XNOR U1726 ( .A(n1054), .B(n1053), .Z(n1055) );
  XOR U1727 ( .A(in[954]), .B(n1055), .Z(n1455) );
  XNOR U1728 ( .A(n1056), .B(n1455), .Z(n3793) );
  XNOR U1729 ( .A(in[570]), .B(n3793), .Z(n1556) );
  XOR U1730 ( .A(in[170]), .B(n3746), .Z(n4799) );
  XOR U1731 ( .A(in[1419]), .B(in[779]), .Z(n1058) );
  XNOR U1732 ( .A(in[1099]), .B(in[459]), .Z(n1057) );
  XNOR U1733 ( .A(n1058), .B(n1057), .Z(n1059) );
  XOR U1734 ( .A(in[139]), .B(n1059), .Z(n1154) );
  XOR U1735 ( .A(in[1290]), .B(in[650]), .Z(n1061) );
  XNOR U1736 ( .A(in[970]), .B(in[330]), .Z(n1060) );
  XNOR U1737 ( .A(n1061), .B(n1060), .Z(n1062) );
  XOR U1738 ( .A(in[10]), .B(n1062), .Z(n1217) );
  XNOR U1739 ( .A(n1154), .B(n1217), .Z(n4092) );
  XNOR U1740 ( .A(in[1355]), .B(n4092), .Z(n4796) );
  NAND U1741 ( .A(n4799), .B(n4796), .Z(n1063) );
  XNOR U1742 ( .A(n1556), .B(n1063), .Z(out[1063]) );
  XOR U1743 ( .A(in[955]), .B(in[1275]), .Z(n1065) );
  XNOR U1744 ( .A(in[1595]), .B(in[315]), .Z(n1064) );
  XNOR U1745 ( .A(n1065), .B(n1064), .Z(n1066) );
  XNOR U1746 ( .A(in[635]), .B(n1066), .Z(n1459) );
  XNOR U1747 ( .A(n1067), .B(n1459), .Z(n3803) );
  XNOR U1748 ( .A(in[571]), .B(n3803), .Z(n1558) );
  NOR U1749 ( .A(n1301), .B(n1696), .Z(n1068) );
  XNOR U1750 ( .A(n1558), .B(n1068), .Z(out[1064]) );
  XOR U1751 ( .A(in[956]), .B(in[1276]), .Z(n1070) );
  XNOR U1752 ( .A(in[1596]), .B(in[316]), .Z(n1069) );
  XNOR U1753 ( .A(n1070), .B(n1069), .Z(n1071) );
  XNOR U1754 ( .A(in[636]), .B(n1071), .Z(n1463) );
  XNOR U1755 ( .A(n1072), .B(n1463), .Z(n3807) );
  XNOR U1756 ( .A(in[572]), .B(n3807), .Z(n1560) );
  NOR U1757 ( .A(n1305), .B(n1700), .Z(n1073) );
  XNOR U1758 ( .A(n1560), .B(n1073), .Z(out[1065]) );
  XOR U1759 ( .A(in[957]), .B(in[1277]), .Z(n1075) );
  XNOR U1760 ( .A(in[1597]), .B(in[317]), .Z(n1074) );
  XNOR U1761 ( .A(n1075), .B(n1074), .Z(n1076) );
  XNOR U1762 ( .A(in[637]), .B(n1076), .Z(n1468) );
  XNOR U1763 ( .A(n1077), .B(n1468), .Z(n3811) );
  XNOR U1764 ( .A(in[573]), .B(n3811), .Z(n1562) );
  NOR U1765 ( .A(n1310), .B(n1704), .Z(n1078) );
  XNOR U1766 ( .A(n1562), .B(n1078), .Z(out[1066]) );
  XOR U1767 ( .A(in[574]), .B(n3815), .Z(n1564) );
  NOR U1768 ( .A(n1314), .B(n1708), .Z(n1079) );
  XNOR U1769 ( .A(n1564), .B(n1079), .Z(out[1067]) );
  XOR U1770 ( .A(in[959]), .B(in[1279]), .Z(n1081) );
  XNOR U1771 ( .A(in[1599]), .B(in[319]), .Z(n1080) );
  XNOR U1772 ( .A(n1081), .B(n1080), .Z(n1082) );
  XNOR U1773 ( .A(in[639]), .B(n1082), .Z(n1476) );
  XNOR U1774 ( .A(n1083), .B(n1476), .Z(n3537) );
  XNOR U1775 ( .A(in[575]), .B(n3537), .Z(n1566) );
  NOR U1776 ( .A(n1318), .B(n1713), .Z(n1084) );
  XNOR U1777 ( .A(n1566), .B(n1084), .Z(out[1068]) );
  XOR U1778 ( .A(in[896]), .B(in[1216]), .Z(n1086) );
  XNOR U1779 ( .A(in[1536]), .B(in[256]), .Z(n1085) );
  XNOR U1780 ( .A(n1086), .B(n1085), .Z(n1087) );
  XNOR U1781 ( .A(in[576]), .B(n1087), .Z(n1480) );
  XNOR U1782 ( .A(n1088), .B(n1480), .Z(n3541) );
  XNOR U1783 ( .A(in[512]), .B(n3541), .Z(n1568) );
  NOR U1784 ( .A(n1322), .B(n1717), .Z(n1089) );
  XNOR U1785 ( .A(n1568), .B(n1089), .Z(out[1069]) );
  XNOR U1786 ( .A(n1091), .B(n1090), .Z(n3616) );
  XNOR U1787 ( .A(in[577]), .B(n3616), .Z(n2563) );
  XOR U1788 ( .A(in[232]), .B(n3717), .Z(n2917) );
  XNOR U1789 ( .A(in[1452]), .B(n3758), .Z(n2914) );
  NAND U1790 ( .A(n2917), .B(n2914), .Z(n1092) );
  XNOR U1791 ( .A(n2563), .B(n1092), .Z(out[106]) );
  XOR U1792 ( .A(in[897]), .B(in[1217]), .Z(n1094) );
  XNOR U1793 ( .A(in[1537]), .B(in[257]), .Z(n1093) );
  XNOR U1794 ( .A(n1094), .B(n1093), .Z(n1095) );
  XNOR U1795 ( .A(in[577]), .B(n1095), .Z(n1484) );
  XNOR U1796 ( .A(n1096), .B(n1484), .Z(n3545) );
  XNOR U1797 ( .A(in[513]), .B(n3545), .Z(n1570) );
  NOR U1798 ( .A(n1326), .B(n1721), .Z(n1097) );
  XNOR U1799 ( .A(n1570), .B(n1097), .Z(out[1070]) );
  XOR U1800 ( .A(in[1538]), .B(in[578]), .Z(n1099) );
  XNOR U1801 ( .A(in[898]), .B(in[258]), .Z(n1098) );
  XNOR U1802 ( .A(n1099), .B(n1098), .Z(n1100) );
  XNOR U1803 ( .A(in[1218]), .B(n1100), .Z(n1488) );
  XNOR U1804 ( .A(n1101), .B(n1488), .Z(n3549) );
  XNOR U1805 ( .A(in[514]), .B(n3549), .Z(n1572) );
  NOR U1806 ( .A(n1330), .B(n1725), .Z(n1102) );
  XNOR U1807 ( .A(n1572), .B(n1102), .Z(out[1071]) );
  XOR U1808 ( .A(in[1539]), .B(in[579]), .Z(n1104) );
  XNOR U1809 ( .A(in[899]), .B(in[259]), .Z(n1103) );
  XNOR U1810 ( .A(n1104), .B(n1103), .Z(n1105) );
  XNOR U1811 ( .A(in[1219]), .B(n1105), .Z(n1492) );
  XNOR U1812 ( .A(n1106), .B(n1492), .Z(n3553) );
  XNOR U1813 ( .A(in[515]), .B(n3553), .Z(n1576) );
  NOR U1814 ( .A(n1334), .B(n1729), .Z(n1107) );
  XNOR U1815 ( .A(n1576), .B(n1107), .Z(out[1072]) );
  XOR U1816 ( .A(in[1540]), .B(in[580]), .Z(n1109) );
  XNOR U1817 ( .A(in[900]), .B(in[260]), .Z(n1108) );
  XNOR U1818 ( .A(n1109), .B(n1108), .Z(n1110) );
  XNOR U1819 ( .A(in[1220]), .B(n1110), .Z(n1496) );
  XNOR U1820 ( .A(n1111), .B(n1496), .Z(n3557) );
  XNOR U1821 ( .A(in[516]), .B(n3557), .Z(n1578) );
  NOR U1822 ( .A(n1338), .B(n1733), .Z(n1112) );
  XNOR U1823 ( .A(n1578), .B(n1112), .Z(out[1073]) );
  XOR U1824 ( .A(in[1541]), .B(in[581]), .Z(n1114) );
  XNOR U1825 ( .A(in[901]), .B(in[261]), .Z(n1113) );
  XNOR U1826 ( .A(n1114), .B(n1113), .Z(n1115) );
  XNOR U1827 ( .A(in[1221]), .B(n1115), .Z(n1500) );
  XNOR U1828 ( .A(n1116), .B(n1500), .Z(n3561) );
  XNOR U1829 ( .A(in[517]), .B(n3561), .Z(n1580) );
  NOR U1830 ( .A(n1342), .B(n1737), .Z(n1117) );
  XNOR U1831 ( .A(n1580), .B(n1117), .Z(out[1074]) );
  XOR U1832 ( .A(in[1542]), .B(in[582]), .Z(n1119) );
  XNOR U1833 ( .A(in[902]), .B(in[262]), .Z(n1118) );
  XNOR U1834 ( .A(n1119), .B(n1118), .Z(n1120) );
  XNOR U1835 ( .A(in[1222]), .B(n1120), .Z(n1504) );
  XNOR U1836 ( .A(n1121), .B(n1504), .Z(n3565) );
  XNOR U1837 ( .A(in[518]), .B(n3565), .Z(n1582) );
  NOR U1838 ( .A(n1346), .B(n1741), .Z(n1122) );
  XNOR U1839 ( .A(n1582), .B(n1122), .Z(out[1075]) );
  XOR U1840 ( .A(in[1543]), .B(in[583]), .Z(n1124) );
  XNOR U1841 ( .A(in[903]), .B(in[263]), .Z(n1123) );
  XNOR U1842 ( .A(n1124), .B(n1123), .Z(n1125) );
  XNOR U1843 ( .A(in[1223]), .B(n1125), .Z(n1509) );
  XNOR U1844 ( .A(n1126), .B(n1509), .Z(n3569) );
  XNOR U1845 ( .A(in[519]), .B(n3569), .Z(n1584) );
  NOR U1846 ( .A(n1351), .B(n1745), .Z(n1127) );
  XNOR U1847 ( .A(n1584), .B(n1127), .Z(out[1076]) );
  XOR U1848 ( .A(in[1544]), .B(in[584]), .Z(n1129) );
  XNOR U1849 ( .A(in[904]), .B(in[264]), .Z(n1128) );
  XNOR U1850 ( .A(n1129), .B(n1128), .Z(n1130) );
  XNOR U1851 ( .A(in[1224]), .B(n1130), .Z(n1513) );
  XNOR U1852 ( .A(n1131), .B(n1513), .Z(n3573) );
  XNOR U1853 ( .A(in[520]), .B(n3573), .Z(n1586) );
  NOR U1854 ( .A(n1355), .B(n1749), .Z(n1132) );
  XNOR U1855 ( .A(n1586), .B(n1132), .Z(out[1077]) );
  XOR U1856 ( .A(in[1545]), .B(in[585]), .Z(n1134) );
  XNOR U1857 ( .A(in[905]), .B(in[265]), .Z(n1133) );
  XNOR U1858 ( .A(n1134), .B(n1133), .Z(n1135) );
  XNOR U1859 ( .A(in[1225]), .B(n1135), .Z(n1517) );
  XNOR U1860 ( .A(n1136), .B(n1517), .Z(n3581) );
  XNOR U1861 ( .A(in[521]), .B(n3581), .Z(n1588) );
  NOR U1862 ( .A(n1359), .B(n1754), .Z(n1137) );
  XNOR U1863 ( .A(n1588), .B(n1137), .Z(out[1078]) );
  XOR U1864 ( .A(in[1546]), .B(in[586]), .Z(n1139) );
  XNOR U1865 ( .A(in[906]), .B(in[266]), .Z(n1138) );
  XNOR U1866 ( .A(n1139), .B(n1138), .Z(n1140) );
  XNOR U1867 ( .A(in[1226]), .B(n1140), .Z(n1521) );
  XNOR U1868 ( .A(n1141), .B(n1521), .Z(n3585) );
  XNOR U1869 ( .A(in[522]), .B(n3585), .Z(n1590) );
  NOR U1870 ( .A(n1363), .B(n1758), .Z(n1142) );
  XNOR U1871 ( .A(n1590), .B(n1142), .Z(out[1079]) );
  XNOR U1872 ( .A(n1144), .B(n1143), .Z(n3624) );
  XNOR U1873 ( .A(in[578]), .B(n3624), .Z(n2565) );
  XOR U1874 ( .A(in[233]), .B(n3721), .Z(n2931) );
  XNOR U1875 ( .A(in[1453]), .B(n3762), .Z(n2928) );
  NAND U1876 ( .A(n2931), .B(n2928), .Z(n1145) );
  XNOR U1877 ( .A(n2565), .B(n1145), .Z(out[107]) );
  XOR U1878 ( .A(in[1547]), .B(in[587]), .Z(n1147) );
  XNOR U1879 ( .A(in[907]), .B(in[267]), .Z(n1146) );
  XNOR U1880 ( .A(n1147), .B(n1146), .Z(n1148) );
  XNOR U1881 ( .A(in[1227]), .B(n1148), .Z(n1525) );
  XNOR U1882 ( .A(n1149), .B(n1525), .Z(n3589) );
  XNOR U1883 ( .A(in[523]), .B(n3589), .Z(n1592) );
  NOR U1884 ( .A(n1367), .B(n1762), .Z(n1150) );
  XNOR U1885 ( .A(n1592), .B(n1150), .Z(out[1080]) );
  XOR U1886 ( .A(in[1548]), .B(in[588]), .Z(n1152) );
  XNOR U1887 ( .A(in[908]), .B(in[268]), .Z(n1151) );
  XNOR U1888 ( .A(n1152), .B(n1151), .Z(n1153) );
  XNOR U1889 ( .A(in[1228]), .B(n1153), .Z(n1529) );
  XNOR U1890 ( .A(n1154), .B(n1529), .Z(n3593) );
  XNOR U1891 ( .A(in[524]), .B(n3593), .Z(n1594) );
  NOR U1892 ( .A(n1371), .B(n1766), .Z(n1155) );
  XNOR U1893 ( .A(n1594), .B(n1155), .Z(out[1081]) );
  XOR U1894 ( .A(in[1549]), .B(in[589]), .Z(n1157) );
  XNOR U1895 ( .A(in[909]), .B(in[269]), .Z(n1156) );
  XNOR U1896 ( .A(n1157), .B(n1156), .Z(n1158) );
  XNOR U1897 ( .A(in[1229]), .B(n1158), .Z(n1533) );
  XNOR U1898 ( .A(n1159), .B(n1533), .Z(n3597) );
  XNOR U1899 ( .A(in[525]), .B(n3597), .Z(n1597) );
  NOR U1900 ( .A(n1375), .B(n1770), .Z(n1160) );
  XNOR U1901 ( .A(n1597), .B(n1160), .Z(out[1082]) );
  XOR U1902 ( .A(in[1550]), .B(in[590]), .Z(n1162) );
  XNOR U1903 ( .A(in[910]), .B(in[270]), .Z(n1161) );
  XNOR U1904 ( .A(n1162), .B(n1161), .Z(n1163) );
  XOR U1905 ( .A(in[1230]), .B(n1163), .Z(n1537) );
  XNOR U1906 ( .A(n1537), .B(n1164), .Z(n3601) );
  XNOR U1907 ( .A(in[526]), .B(n3601), .Z(n1599) );
  NOR U1908 ( .A(n1379), .B(n1774), .Z(n1165) );
  XNOR U1909 ( .A(n1599), .B(n1165), .Z(out[1083]) );
  XOR U1910 ( .A(in[1551]), .B(in[591]), .Z(n1167) );
  XNOR U1911 ( .A(in[911]), .B(in[271]), .Z(n1166) );
  XNOR U1912 ( .A(n1167), .B(n1166), .Z(n1168) );
  XOR U1913 ( .A(in[1231]), .B(n1168), .Z(n1541) );
  XNOR U1914 ( .A(n1541), .B(n1169), .Z(n3605) );
  XNOR U1915 ( .A(in[527]), .B(n3605), .Z(n1601) );
  NOR U1916 ( .A(n1383), .B(n1778), .Z(n1170) );
  XNOR U1917 ( .A(n1601), .B(n1170), .Z(out[1084]) );
  XOR U1918 ( .A(in[1552]), .B(in[592]), .Z(n1172) );
  XNOR U1919 ( .A(in[912]), .B(in[272]), .Z(n1171) );
  XNOR U1920 ( .A(n1172), .B(n1171), .Z(n1173) );
  XNOR U1921 ( .A(in[1232]), .B(n1173), .Z(n1545) );
  XNOR U1922 ( .A(n1174), .B(n1545), .Z(n3609) );
  XNOR U1923 ( .A(in[528]), .B(n3609), .Z(n1603) );
  NOR U1924 ( .A(n1387), .B(n1782), .Z(n1175) );
  XNOR U1925 ( .A(n1603), .B(n1175), .Z(out[1085]) );
  XOR U1926 ( .A(in[1553]), .B(in[593]), .Z(n1177) );
  XNOR U1927 ( .A(in[913]), .B(in[273]), .Z(n1176) );
  XNOR U1928 ( .A(n1177), .B(n1176), .Z(n1178) );
  XNOR U1929 ( .A(in[1233]), .B(n1178), .Z(n1550) );
  XNOR U1930 ( .A(n1179), .B(n1550), .Z(n3613) );
  XNOR U1931 ( .A(in[529]), .B(n3613), .Z(n1605) );
  NOR U1932 ( .A(n1390), .B(n1786), .Z(n1180) );
  XNOR U1933 ( .A(n1605), .B(n1180), .Z(out[1086]) );
  XOR U1934 ( .A(in[1554]), .B(in[594]), .Z(n1182) );
  XNOR U1935 ( .A(in[914]), .B(in[274]), .Z(n1181) );
  XNOR U1936 ( .A(n1182), .B(n1181), .Z(n1183) );
  XOR U1937 ( .A(in[1234]), .B(n1183), .Z(n1554) );
  XNOR U1938 ( .A(n1554), .B(n1184), .Z(n3617) );
  XNOR U1939 ( .A(in[530]), .B(n3617), .Z(n1607) );
  NOR U1940 ( .A(n1392), .B(n1790), .Z(n1185) );
  XNOR U1941 ( .A(n1607), .B(n1185), .Z(out[1087]) );
  XOR U1942 ( .A(in[957]), .B(n3600), .Z(n1609) );
  NOR U1943 ( .A(n1396), .B(n4631), .Z(n1186) );
  XNOR U1944 ( .A(n1609), .B(n1186), .Z(out[1088]) );
  XOR U1945 ( .A(in[958]), .B(n3604), .Z(n1611) );
  NOR U1946 ( .A(n1400), .B(n4635), .Z(n1187) );
  XNOR U1947 ( .A(n1611), .B(n1187), .Z(out[1089]) );
  XOR U1948 ( .A(n1189), .B(n1188), .Z(n3628) );
  XNOR U1949 ( .A(in[579]), .B(n3628), .Z(n2567) );
  XOR U1950 ( .A(in[234]), .B(n3725), .Z(n2947) );
  XNOR U1951 ( .A(in[1454]), .B(n3766), .Z(n2944) );
  NAND U1952 ( .A(n2947), .B(n2944), .Z(n1190) );
  XNOR U1953 ( .A(n2567), .B(n1190), .Z(out[108]) );
  XOR U1954 ( .A(in[959]), .B(n3608), .Z(n1613) );
  NOR U1955 ( .A(n1404), .B(n4639), .Z(n1191) );
  XNOR U1956 ( .A(n1613), .B(n1191), .Z(out[1090]) );
  XOR U1957 ( .A(in[896]), .B(n3612), .Z(n1615) );
  NOR U1958 ( .A(n1408), .B(n4643), .Z(n1192) );
  XNOR U1959 ( .A(n1615), .B(n1192), .Z(out[1091]) );
  XOR U1960 ( .A(in[897]), .B(n3616), .Z(n1618) );
  NOR U1961 ( .A(n1412), .B(n4647), .Z(n1193) );
  XNOR U1962 ( .A(n1618), .B(n1193), .Z(out[1092]) );
  XOR U1963 ( .A(in[898]), .B(n3624), .Z(n1620) );
  NOR U1964 ( .A(n1416), .B(n4651), .Z(n1194) );
  XNOR U1965 ( .A(n1620), .B(n1194), .Z(out[1093]) );
  XOR U1966 ( .A(in[899]), .B(n3628), .Z(n1622) );
  NOR U1967 ( .A(n1420), .B(n4655), .Z(n1195) );
  XNOR U1968 ( .A(n1622), .B(n1195), .Z(out[1094]) );
  XNOR U1969 ( .A(n1197), .B(n1196), .Z(n3632) );
  XNOR U1970 ( .A(in[900]), .B(n3632), .Z(n1624) );
  NOR U1971 ( .A(n1424), .B(n4659), .Z(n1198) );
  XNOR U1972 ( .A(n1624), .B(n1198), .Z(out[1095]) );
  XNOR U1973 ( .A(n1200), .B(n1199), .Z(n3636) );
  XNOR U1974 ( .A(in[901]), .B(n3636), .Z(n1626) );
  NOR U1975 ( .A(n1429), .B(n4663), .Z(n1201) );
  XNOR U1976 ( .A(n1626), .B(n1201), .Z(out[1096]) );
  XNOR U1977 ( .A(n1203), .B(n1202), .Z(n3640) );
  XNOR U1978 ( .A(in[902]), .B(n3640), .Z(n1628) );
  NOR U1979 ( .A(n1433), .B(n4667), .Z(n1204) );
  XNOR U1980 ( .A(n1628), .B(n1204), .Z(out[1097]) );
  XNOR U1981 ( .A(n1206), .B(n1205), .Z(n3644) );
  XNOR U1982 ( .A(in[903]), .B(n3644), .Z(n1630) );
  NOR U1983 ( .A(n1437), .B(n4675), .Z(n1207) );
  XNOR U1984 ( .A(n1630), .B(n1207), .Z(out[1098]) );
  XNOR U1985 ( .A(n1209), .B(n1208), .Z(n3648) );
  XNOR U1986 ( .A(in[904]), .B(n3648), .Z(n1632) );
  NOR U1987 ( .A(n1441), .B(n4679), .Z(n1210) );
  XNOR U1988 ( .A(n1632), .B(n1210), .Z(out[1099]) );
  XOR U1989 ( .A(in[580]), .B(n3632), .Z(n2569) );
  XOR U1990 ( .A(in[235]), .B(n3729), .Z(n2971) );
  XNOR U1991 ( .A(in[1455]), .B(n3770), .Z(n2968) );
  NAND U1992 ( .A(n2971), .B(n2968), .Z(n1211) );
  XNOR U1993 ( .A(n2569), .B(n1211), .Z(out[109]) );
  XOR U1994 ( .A(in[200]), .B(n3573), .Z(n3921) );
  XNOR U1995 ( .A(in[1420]), .B(n3614), .Z(n3920) );
  XOR U1996 ( .A(n4120), .B(in[1043]), .Z(n2632) );
  NAND U1997 ( .A(n3920), .B(n2632), .Z(n1212) );
  XNOR U1998 ( .A(n3921), .B(n1212), .Z(out[10]) );
  XNOR U1999 ( .A(n1214), .B(n1213), .Z(n3652) );
  XNOR U2000 ( .A(in[905]), .B(n3652), .Z(n1634) );
  NOR U2001 ( .A(n1445), .B(n4683), .Z(n1215) );
  XNOR U2002 ( .A(n1634), .B(n1215), .Z(out[1100]) );
  XNOR U2003 ( .A(n1217), .B(n1216), .Z(n3656) );
  XNOR U2004 ( .A(in[906]), .B(n3656), .Z(n1636) );
  NOR U2005 ( .A(n1449), .B(n4687), .Z(n1218) );
  XNOR U2006 ( .A(n1636), .B(n1218), .Z(out[1101]) );
  XOR U2007 ( .A(n1220), .B(n1219), .Z(n3660) );
  XNOR U2008 ( .A(in[907]), .B(n3660), .Z(n1639) );
  NOR U2009 ( .A(n1453), .B(n4691), .Z(n1221) );
  XNOR U2010 ( .A(n1639), .B(n1221), .Z(out[1102]) );
  XOR U2011 ( .A(n1223), .B(n1222), .Z(n3668) );
  XNOR U2012 ( .A(in[908]), .B(n3668), .Z(n1641) );
  NOR U2013 ( .A(n1457), .B(n4695), .Z(n1224) );
  XNOR U2014 ( .A(n1641), .B(n1224), .Z(out[1103]) );
  XNOR U2015 ( .A(n1226), .B(n1225), .Z(n3672) );
  XNOR U2016 ( .A(in[909]), .B(n3672), .Z(n1643) );
  NOR U2017 ( .A(n1461), .B(n4699), .Z(n1227) );
  XNOR U2018 ( .A(n1643), .B(n1227), .Z(out[1104]) );
  XOR U2019 ( .A(n1229), .B(n1228), .Z(n3676) );
  XNOR U2020 ( .A(in[910]), .B(n3676), .Z(n1645) );
  NOR U2021 ( .A(n1465), .B(n4703), .Z(n1230) );
  XNOR U2022 ( .A(n1645), .B(n1230), .Z(out[1105]) );
  XOR U2023 ( .A(n1232), .B(n1231), .Z(n3680) );
  XNOR U2024 ( .A(in[911]), .B(n3680), .Z(n1647) );
  NOR U2025 ( .A(n1470), .B(n4707), .Z(n1233) );
  XNOR U2026 ( .A(n1647), .B(n1233), .Z(out[1106]) );
  XNOR U2027 ( .A(n1235), .B(n1234), .Z(n3684) );
  XNOR U2028 ( .A(in[912]), .B(n3684), .Z(n1649) );
  NOR U2029 ( .A(n1474), .B(n4711), .Z(n1236) );
  XNOR U2030 ( .A(n1649), .B(n1236), .Z(out[1107]) );
  XOR U2031 ( .A(n1238), .B(n1237), .Z(n3688) );
  XNOR U2032 ( .A(in[913]), .B(n3688), .Z(n1651) );
  NOR U2033 ( .A(n1478), .B(n4719), .Z(n1239) );
  XNOR U2034 ( .A(n1651), .B(n1239), .Z(out[1108]) );
  XNOR U2035 ( .A(n1241), .B(n1240), .Z(n3692) );
  XNOR U2036 ( .A(in[914]), .B(n3692), .Z(n1653) );
  NOR U2037 ( .A(n1482), .B(n4723), .Z(n1242) );
  XNOR U2038 ( .A(n1653), .B(n1242), .Z(out[1109]) );
  XOR U2039 ( .A(in[581]), .B(n3636), .Z(n2571) );
  XOR U2040 ( .A(in[236]), .B(n3733), .Z(n2995) );
  XNOR U2041 ( .A(in[1456]), .B(n3774), .Z(n2992) );
  NAND U2042 ( .A(n2995), .B(n2992), .Z(n1243) );
  XNOR U2043 ( .A(n2571), .B(n1243), .Z(out[110]) );
  XOR U2044 ( .A(n1245), .B(n1244), .Z(n3696) );
  XNOR U2045 ( .A(in[915]), .B(n3696), .Z(n1655) );
  NOR U2046 ( .A(n1486), .B(n4727), .Z(n1246) );
  XNOR U2047 ( .A(n1655), .B(n1246), .Z(out[1110]) );
  XNOR U2048 ( .A(n1248), .B(n1247), .Z(n3700) );
  XNOR U2049 ( .A(in[916]), .B(n3700), .Z(n1657) );
  NOR U2050 ( .A(n1490), .B(n4731), .Z(n1249) );
  XNOR U2051 ( .A(n1657), .B(n1249), .Z(out[1111]) );
  XNOR U2052 ( .A(n1251), .B(n1250), .Z(n3704) );
  XNOR U2053 ( .A(in[917]), .B(n3704), .Z(n1660) );
  NOR U2054 ( .A(n1494), .B(n4735), .Z(n1252) );
  XNOR U2055 ( .A(n1660), .B(n1252), .Z(out[1112]) );
  XOR U2056 ( .A(n1254), .B(n1253), .Z(n3712) );
  XNOR U2057 ( .A(in[918]), .B(n3712), .Z(n1662) );
  NOR U2058 ( .A(n1498), .B(n4739), .Z(n1255) );
  XNOR U2059 ( .A(n1662), .B(n1255), .Z(out[1113]) );
  XNOR U2060 ( .A(n1257), .B(n1256), .Z(n3716) );
  XNOR U2061 ( .A(in[919]), .B(n3716), .Z(n1664) );
  NOR U2062 ( .A(n1502), .B(n4743), .Z(n1258) );
  XNOR U2063 ( .A(n1664), .B(n1258), .Z(out[1114]) );
  XOR U2064 ( .A(n1260), .B(n1259), .Z(n3720) );
  XNOR U2065 ( .A(in[920]), .B(n3720), .Z(n1666) );
  NOR U2066 ( .A(n1506), .B(n4747), .Z(n1261) );
  XNOR U2067 ( .A(n1666), .B(n1261), .Z(out[1115]) );
  XNOR U2068 ( .A(n1263), .B(n1262), .Z(n3724) );
  XNOR U2069 ( .A(in[921]), .B(n3724), .Z(n1668) );
  NOR U2070 ( .A(n1511), .B(n4751), .Z(n1264) );
  XNOR U2071 ( .A(n1668), .B(n1264), .Z(out[1116]) );
  XOR U2072 ( .A(n1266), .B(n1265), .Z(n3728) );
  XNOR U2073 ( .A(in[922]), .B(n3728), .Z(n1670) );
  NOR U2074 ( .A(n1515), .B(n4755), .Z(n1267) );
  XNOR U2075 ( .A(n1670), .B(n1267), .Z(out[1117]) );
  XOR U2076 ( .A(n1269), .B(n1268), .Z(n3732) );
  XNOR U2077 ( .A(in[923]), .B(n3732), .Z(n1672) );
  NOR U2078 ( .A(n1519), .B(n4763), .Z(n1270) );
  XNOR U2079 ( .A(n1672), .B(n1270), .Z(out[1118]) );
  XOR U2080 ( .A(n1272), .B(n1271), .Z(n3736) );
  XNOR U2081 ( .A(in[924]), .B(n3736), .Z(n1674) );
  NOR U2082 ( .A(n1523), .B(n4767), .Z(n1273) );
  XNOR U2083 ( .A(n1674), .B(n1273), .Z(out[1119]) );
  XOR U2084 ( .A(in[582]), .B(n3640), .Z(n2573) );
  XOR U2085 ( .A(in[237]), .B(n3737), .Z(n3019) );
  XNOR U2086 ( .A(in[1457]), .B(n3778), .Z(n3016) );
  NAND U2087 ( .A(n3019), .B(n3016), .Z(n1274) );
  XNOR U2088 ( .A(n2573), .B(n1274), .Z(out[111]) );
  XOR U2089 ( .A(n1276), .B(n1275), .Z(n3740) );
  XNOR U2090 ( .A(in[925]), .B(n3740), .Z(n1676) );
  NOR U2091 ( .A(n1527), .B(n4771), .Z(n1277) );
  XNOR U2092 ( .A(n1676), .B(n1277), .Z(out[1120]) );
  XOR U2093 ( .A(n1279), .B(n1278), .Z(n3744) );
  XNOR U2094 ( .A(in[926]), .B(n3744), .Z(n1678) );
  NOR U2095 ( .A(n1531), .B(n4775), .Z(n1280) );
  XNOR U2096 ( .A(n1678), .B(n1280), .Z(out[1121]) );
  XOR U2097 ( .A(n1282), .B(n1281), .Z(n3748) );
  XNOR U2098 ( .A(in[927]), .B(n3748), .Z(n1681) );
  NOR U2099 ( .A(n1535), .B(n4779), .Z(n1283) );
  XNOR U2100 ( .A(n1681), .B(n1283), .Z(out[1122]) );
  XOR U2101 ( .A(n1285), .B(n1284), .Z(n3756) );
  XNOR U2102 ( .A(in[928]), .B(n3756), .Z(n1683) );
  NOR U2103 ( .A(n1539), .B(n4783), .Z(n1286) );
  XNOR U2104 ( .A(n1683), .B(n1286), .Z(out[1123]) );
  XNOR U2105 ( .A(n1288), .B(n1287), .Z(n3760) );
  XNOR U2106 ( .A(in[929]), .B(n3760), .Z(n1685) );
  NOR U2107 ( .A(n1543), .B(n4787), .Z(n1289) );
  XNOR U2108 ( .A(n1685), .B(n1289), .Z(out[1124]) );
  XOR U2109 ( .A(n1291), .B(n1290), .Z(n3764) );
  XNOR U2110 ( .A(in[930]), .B(n3764), .Z(n1687) );
  NOR U2111 ( .A(n1547), .B(n4791), .Z(n1292) );
  XNOR U2112 ( .A(n1687), .B(n1292), .Z(out[1125]) );
  XNOR U2113 ( .A(n1294), .B(n1293), .Z(n3768) );
  XNOR U2114 ( .A(in[931]), .B(n3768), .Z(n1689) );
  NOR U2115 ( .A(n1552), .B(n4795), .Z(n1295) );
  XNOR U2116 ( .A(n1689), .B(n1295), .Z(out[1126]) );
  XNOR U2117 ( .A(n1297), .B(n1296), .Z(n3772) );
  XNOR U2118 ( .A(in[932]), .B(n3772), .Z(n1691) );
  NOR U2119 ( .A(n1556), .B(n4799), .Z(n1298) );
  XNOR U2120 ( .A(n1691), .B(n1298), .Z(out[1127]) );
  XNOR U2121 ( .A(n1300), .B(n1299), .Z(n3776) );
  XNOR U2122 ( .A(in[933]), .B(n3776), .Z(n1694) );
  NAND U2123 ( .A(n1558), .B(n1301), .Z(n1302) );
  XNOR U2124 ( .A(n1694), .B(n1302), .Z(out[1128]) );
  XOR U2125 ( .A(n1304), .B(n1303), .Z(n3780) );
  XNOR U2126 ( .A(in[934]), .B(n3780), .Z(n1698) );
  NAND U2127 ( .A(n1560), .B(n1305), .Z(n1306) );
  XNOR U2128 ( .A(n1698), .B(n1306), .Z(out[1129]) );
  XOR U2129 ( .A(in[583]), .B(n3644), .Z(n2576) );
  XOR U2130 ( .A(in[238]), .B(n3741), .Z(n3043) );
  XNOR U2131 ( .A(in[1458]), .B(n3782), .Z(n3040) );
  NAND U2132 ( .A(n3043), .B(n3040), .Z(n1307) );
  XNOR U2133 ( .A(n2576), .B(n1307), .Z(out[112]) );
  XNOR U2134 ( .A(n1309), .B(n1308), .Z(n3784) );
  XNOR U2135 ( .A(in[935]), .B(n3784), .Z(n1702) );
  NAND U2136 ( .A(n1562), .B(n1310), .Z(n1311) );
  XNOR U2137 ( .A(n1702), .B(n1311), .Z(out[1130]) );
  XNOR U2138 ( .A(n1313), .B(n1312), .Z(n3788) );
  XNOR U2139 ( .A(in[936]), .B(n3788), .Z(n1706) );
  NAND U2140 ( .A(n1564), .B(n1314), .Z(n1315) );
  XNOR U2141 ( .A(n1706), .B(n1315), .Z(out[1131]) );
  XNOR U2142 ( .A(n1317), .B(n1316), .Z(n3792) );
  XNOR U2143 ( .A(in[937]), .B(n3792), .Z(n1711) );
  NAND U2144 ( .A(n1566), .B(n1318), .Z(n1319) );
  XNOR U2145 ( .A(n1711), .B(n1319), .Z(out[1132]) );
  XNOR U2146 ( .A(n1321), .B(n1320), .Z(n3802) );
  XNOR U2147 ( .A(in[938]), .B(n3802), .Z(n1715) );
  NAND U2148 ( .A(n1568), .B(n1322), .Z(n1323) );
  XNOR U2149 ( .A(n1715), .B(n1323), .Z(out[1133]) );
  XNOR U2150 ( .A(n1325), .B(n1324), .Z(n3806) );
  XNOR U2151 ( .A(in[939]), .B(n3806), .Z(n1719) );
  NAND U2152 ( .A(n1570), .B(n1326), .Z(n1327) );
  XNOR U2153 ( .A(n1719), .B(n1327), .Z(out[1134]) );
  XNOR U2154 ( .A(n1329), .B(n1328), .Z(n3810) );
  XNOR U2155 ( .A(in[940]), .B(n3810), .Z(n1723) );
  NAND U2156 ( .A(n1572), .B(n1330), .Z(n1331) );
  XNOR U2157 ( .A(n1723), .B(n1331), .Z(out[1135]) );
  XNOR U2158 ( .A(n1333), .B(n1332), .Z(n3814) );
  XNOR U2159 ( .A(in[941]), .B(n3814), .Z(n1727) );
  NAND U2160 ( .A(n1576), .B(n1334), .Z(n1335) );
  XNOR U2161 ( .A(n1727), .B(n1335), .Z(out[1136]) );
  XNOR U2162 ( .A(n1337), .B(n1336), .Z(n3536) );
  XNOR U2163 ( .A(in[942]), .B(n3536), .Z(n1731) );
  NAND U2164 ( .A(n1578), .B(n1338), .Z(n1339) );
  XNOR U2165 ( .A(n1731), .B(n1339), .Z(out[1137]) );
  XNOR U2166 ( .A(n1341), .B(n1340), .Z(n3540) );
  XNOR U2167 ( .A(in[943]), .B(n3540), .Z(n1735) );
  NAND U2168 ( .A(n1580), .B(n1342), .Z(n1343) );
  XNOR U2169 ( .A(n1735), .B(n1343), .Z(out[1138]) );
  XNOR U2170 ( .A(n1345), .B(n1344), .Z(n3544) );
  XNOR U2171 ( .A(in[944]), .B(n3544), .Z(n1739) );
  NAND U2172 ( .A(n1582), .B(n1346), .Z(n1347) );
  XNOR U2173 ( .A(n1739), .B(n1347), .Z(out[1139]) );
  XOR U2174 ( .A(in[584]), .B(n3648), .Z(n2578) );
  XOR U2175 ( .A(in[239]), .B(n3745), .Z(n3067) );
  XNOR U2176 ( .A(in[1459]), .B(n3786), .Z(n3064) );
  NAND U2177 ( .A(n3067), .B(n3064), .Z(n1348) );
  XNOR U2178 ( .A(n2578), .B(n1348), .Z(out[113]) );
  XNOR U2179 ( .A(n1350), .B(n1349), .Z(n3548) );
  XNOR U2180 ( .A(in[945]), .B(n3548), .Z(n1743) );
  NAND U2181 ( .A(n1584), .B(n1351), .Z(n1352) );
  XNOR U2182 ( .A(n1743), .B(n1352), .Z(out[1140]) );
  XNOR U2183 ( .A(n1354), .B(n1353), .Z(n3552) );
  XNOR U2184 ( .A(in[946]), .B(n3552), .Z(n1747) );
  NAND U2185 ( .A(n1586), .B(n1355), .Z(n1356) );
  XNOR U2186 ( .A(n1747), .B(n1356), .Z(out[1141]) );
  XNOR U2187 ( .A(n1358), .B(n1357), .Z(n3556) );
  XNOR U2188 ( .A(in[947]), .B(n3556), .Z(n1752) );
  NAND U2189 ( .A(n1588), .B(n1359), .Z(n1360) );
  XNOR U2190 ( .A(n1752), .B(n1360), .Z(out[1142]) );
  XNOR U2191 ( .A(n1362), .B(n1361), .Z(n3560) );
  XNOR U2192 ( .A(in[948]), .B(n3560), .Z(n1756) );
  NAND U2193 ( .A(n1590), .B(n1363), .Z(n1364) );
  XNOR U2194 ( .A(n1756), .B(n1364), .Z(out[1143]) );
  XNOR U2195 ( .A(n1366), .B(n1365), .Z(n3564) );
  XNOR U2196 ( .A(in[949]), .B(n3564), .Z(n1760) );
  NAND U2197 ( .A(n1592), .B(n1367), .Z(n1368) );
  XNOR U2198 ( .A(n1760), .B(n1368), .Z(out[1144]) );
  XNOR U2199 ( .A(n1370), .B(n1369), .Z(n3568) );
  XNOR U2200 ( .A(in[950]), .B(n3568), .Z(n1764) );
  NAND U2201 ( .A(n1594), .B(n1371), .Z(n1372) );
  XNOR U2202 ( .A(n1764), .B(n1372), .Z(out[1145]) );
  XNOR U2203 ( .A(n1374), .B(n1373), .Z(n3572) );
  XNOR U2204 ( .A(in[951]), .B(n3572), .Z(n1768) );
  NAND U2205 ( .A(n1597), .B(n1375), .Z(n1376) );
  XNOR U2206 ( .A(n1768), .B(n1376), .Z(out[1146]) );
  XNOR U2207 ( .A(n1378), .B(n1377), .Z(n3580) );
  XNOR U2208 ( .A(in[952]), .B(n3580), .Z(n1772) );
  NAND U2209 ( .A(n1599), .B(n1379), .Z(n1380) );
  XNOR U2210 ( .A(n1772), .B(n1380), .Z(out[1147]) );
  XNOR U2211 ( .A(n1382), .B(n1381), .Z(n3584) );
  XNOR U2212 ( .A(in[953]), .B(n3584), .Z(n1776) );
  NAND U2213 ( .A(n1601), .B(n1383), .Z(n1384) );
  XNOR U2214 ( .A(n1776), .B(n1384), .Z(out[1148]) );
  XNOR U2215 ( .A(n1386), .B(n1385), .Z(n3588) );
  XNOR U2216 ( .A(in[954]), .B(n3588), .Z(n1780) );
  NAND U2217 ( .A(n1603), .B(n1387), .Z(n1388) );
  XNOR U2218 ( .A(n1780), .B(n1388), .Z(out[1149]) );
  XOR U2219 ( .A(in[585]), .B(n3652), .Z(n2580) );
  XOR U2220 ( .A(in[240]), .B(n3749), .Z(n3093) );
  XNOR U2221 ( .A(in[1460]), .B(n3790), .Z(n3090) );
  NAND U2222 ( .A(n3093), .B(n3090), .Z(n1389) );
  XNOR U2223 ( .A(n2580), .B(n1389), .Z(out[114]) );
  XNOR U2224 ( .A(in[955]), .B(n3592), .Z(n1784) );
  NAND U2225 ( .A(n1605), .B(n1390), .Z(n1391) );
  XNOR U2226 ( .A(n1784), .B(n1391), .Z(out[1150]) );
  XNOR U2227 ( .A(in[956]), .B(n3596), .Z(n1788) );
  NAND U2228 ( .A(n1607), .B(n1392), .Z(n1393) );
  XNOR U2229 ( .A(n1788), .B(n1393), .Z(out[1151]) );
  XNOR U2230 ( .A(n1395), .B(n1394), .Z(n3936) );
  XNOR U2231 ( .A(in[1004]), .B(n3936), .Z(n4629) );
  NAND U2232 ( .A(n1609), .B(n1396), .Z(n1397) );
  XNOR U2233 ( .A(n4629), .B(n1397), .Z(out[1152]) );
  XNOR U2234 ( .A(n1399), .B(n1398), .Z(n3938) );
  XNOR U2235 ( .A(in[1005]), .B(n3938), .Z(n4633) );
  NAND U2236 ( .A(n1611), .B(n1400), .Z(n1401) );
  XNOR U2237 ( .A(n4633), .B(n1401), .Z(out[1153]) );
  XNOR U2238 ( .A(n1403), .B(n1402), .Z(n3940) );
  XNOR U2239 ( .A(in[1006]), .B(n3940), .Z(n4637) );
  NAND U2240 ( .A(n1613), .B(n1404), .Z(n1405) );
  XNOR U2241 ( .A(n4637), .B(n1405), .Z(out[1154]) );
  XNOR U2242 ( .A(n1407), .B(n1406), .Z(n3942) );
  XNOR U2243 ( .A(in[1007]), .B(n3942), .Z(n4641) );
  NAND U2244 ( .A(n1615), .B(n1408), .Z(n1409) );
  XNOR U2245 ( .A(n4641), .B(n1409), .Z(out[1155]) );
  XNOR U2246 ( .A(n1411), .B(n1410), .Z(n3948) );
  XNOR U2247 ( .A(in[1008]), .B(n3948), .Z(n4645) );
  NAND U2248 ( .A(n1618), .B(n1412), .Z(n1413) );
  XNOR U2249 ( .A(n4645), .B(n1413), .Z(out[1156]) );
  XNOR U2250 ( .A(n1415), .B(n1414), .Z(n3950) );
  XNOR U2251 ( .A(in[1009]), .B(n3950), .Z(n4649) );
  NAND U2252 ( .A(n1620), .B(n1416), .Z(n1417) );
  XNOR U2253 ( .A(n4649), .B(n1417), .Z(out[1157]) );
  XNOR U2254 ( .A(n1419), .B(n1418), .Z(n3952) );
  XNOR U2255 ( .A(in[1010]), .B(n3952), .Z(n4653) );
  NAND U2256 ( .A(n1622), .B(n1420), .Z(n1421) );
  XNOR U2257 ( .A(n4653), .B(n1421), .Z(out[1158]) );
  XNOR U2258 ( .A(n1423), .B(n1422), .Z(n3954) );
  XNOR U2259 ( .A(in[1011]), .B(n3954), .Z(n4657) );
  NAND U2260 ( .A(n1624), .B(n1424), .Z(n1425) );
  XNOR U2261 ( .A(n4657), .B(n1425), .Z(out[1159]) );
  XOR U2262 ( .A(in[586]), .B(n3656), .Z(n2582) );
  XOR U2263 ( .A(in[241]), .B(n3757), .Z(n3117) );
  XNOR U2264 ( .A(in[1461]), .B(n3794), .Z(n3114) );
  NAND U2265 ( .A(n3117), .B(n3114), .Z(n1426) );
  XNOR U2266 ( .A(n2582), .B(n1426), .Z(out[115]) );
  XNOR U2267 ( .A(n1428), .B(n1427), .Z(n3956) );
  XNOR U2268 ( .A(in[1012]), .B(n3956), .Z(n4661) );
  NAND U2269 ( .A(n1626), .B(n1429), .Z(n1430) );
  XNOR U2270 ( .A(n4661), .B(n1430), .Z(out[1160]) );
  XNOR U2271 ( .A(n1432), .B(n1431), .Z(n3958) );
  XNOR U2272 ( .A(in[1013]), .B(n3958), .Z(n4665) );
  NAND U2273 ( .A(n1628), .B(n1433), .Z(n1434) );
  XNOR U2274 ( .A(n4665), .B(n1434), .Z(out[1161]) );
  XNOR U2275 ( .A(n1436), .B(n1435), .Z(n3960) );
  XNOR U2276 ( .A(in[1014]), .B(n3960), .Z(n4673) );
  NAND U2277 ( .A(n1630), .B(n1437), .Z(n1438) );
  XNOR U2278 ( .A(n4673), .B(n1438), .Z(out[1162]) );
  XNOR U2279 ( .A(n1440), .B(n1439), .Z(n3962) );
  XNOR U2280 ( .A(in[1015]), .B(n3962), .Z(n4677) );
  NAND U2281 ( .A(n1632), .B(n1441), .Z(n1442) );
  XNOR U2282 ( .A(n4677), .B(n1442), .Z(out[1163]) );
  XNOR U2283 ( .A(n1444), .B(n1443), .Z(n3818) );
  XNOR U2284 ( .A(in[1016]), .B(n3818), .Z(n4681) );
  NAND U2285 ( .A(n1634), .B(n1445), .Z(n1446) );
  XNOR U2286 ( .A(n4681), .B(n1446), .Z(out[1164]) );
  XNOR U2287 ( .A(n1448), .B(n1447), .Z(n3820) );
  XNOR U2288 ( .A(in[1017]), .B(n3820), .Z(n4685) );
  NAND U2289 ( .A(n1636), .B(n1449), .Z(n1450) );
  XNOR U2290 ( .A(n4685), .B(n1450), .Z(out[1165]) );
  XNOR U2291 ( .A(n1452), .B(n1451), .Z(n3822) );
  XNOR U2292 ( .A(in[1018]), .B(n3822), .Z(n4689) );
  NAND U2293 ( .A(n1639), .B(n1453), .Z(n1454) );
  XNOR U2294 ( .A(n4689), .B(n1454), .Z(out[1166]) );
  XNOR U2295 ( .A(n1456), .B(n1455), .Z(n3824) );
  XNOR U2296 ( .A(in[1019]), .B(n3824), .Z(n4693) );
  NAND U2297 ( .A(n1641), .B(n1457), .Z(n1458) );
  XNOR U2298 ( .A(n4693), .B(n1458), .Z(out[1167]) );
  XOR U2299 ( .A(n1460), .B(n1459), .Z(n3826) );
  XNOR U2300 ( .A(in[1020]), .B(n3826), .Z(n4697) );
  NAND U2301 ( .A(n1643), .B(n1461), .Z(n1462) );
  XNOR U2302 ( .A(n4697), .B(n1462), .Z(out[1168]) );
  XOR U2303 ( .A(n1464), .B(n1463), .Z(n3828) );
  XNOR U2304 ( .A(in[1021]), .B(n3828), .Z(n4701) );
  NAND U2305 ( .A(n1645), .B(n1465), .Z(n1466) );
  XNOR U2306 ( .A(n4701), .B(n1466), .Z(out[1169]) );
  XOR U2307 ( .A(in[587]), .B(n3660), .Z(n2584) );
  XOR U2308 ( .A(in[242]), .B(n3761), .Z(n3141) );
  XNOR U2309 ( .A(in[1462]), .B(n3804), .Z(n3138) );
  NAND U2310 ( .A(n3141), .B(n3138), .Z(n1467) );
  XNOR U2311 ( .A(n2584), .B(n1467), .Z(out[116]) );
  XOR U2312 ( .A(n1469), .B(n1468), .Z(n3834) );
  XNOR U2313 ( .A(in[1022]), .B(n3834), .Z(n4705) );
  NAND U2314 ( .A(n1647), .B(n1470), .Z(n1471) );
  XNOR U2315 ( .A(n4705), .B(n1471), .Z(out[1170]) );
  XNOR U2316 ( .A(n1473), .B(n1472), .Z(n3836) );
  XNOR U2317 ( .A(in[1023]), .B(n3836), .Z(n4709) );
  NAND U2318 ( .A(n1649), .B(n1474), .Z(n1475) );
  XNOR U2319 ( .A(n4709), .B(n1475), .Z(out[1171]) );
  XOR U2320 ( .A(n1477), .B(n1476), .Z(n3838) );
  XNOR U2321 ( .A(in[960]), .B(n3838), .Z(n4717) );
  NAND U2322 ( .A(n1651), .B(n1478), .Z(n1479) );
  XNOR U2323 ( .A(n4717), .B(n1479), .Z(out[1172]) );
  XOR U2324 ( .A(n1481), .B(n1480), .Z(n3840) );
  XNOR U2325 ( .A(in[961]), .B(n3840), .Z(n4721) );
  NAND U2326 ( .A(n1653), .B(n1482), .Z(n1483) );
  XNOR U2327 ( .A(n4721), .B(n1483), .Z(out[1173]) );
  XOR U2328 ( .A(n1485), .B(n1484), .Z(n3842) );
  XNOR U2329 ( .A(in[962]), .B(n3842), .Z(n4725) );
  NAND U2330 ( .A(n1655), .B(n1486), .Z(n1487) );
  XNOR U2331 ( .A(n4725), .B(n1487), .Z(out[1174]) );
  XOR U2332 ( .A(n1489), .B(n1488), .Z(n3844) );
  XNOR U2333 ( .A(in[963]), .B(n3844), .Z(n4729) );
  NAND U2334 ( .A(n1657), .B(n1490), .Z(n1491) );
  XNOR U2335 ( .A(n4729), .B(n1491), .Z(out[1175]) );
  XOR U2336 ( .A(n1493), .B(n1492), .Z(n3846) );
  XNOR U2337 ( .A(in[964]), .B(n3846), .Z(n4733) );
  NAND U2338 ( .A(n1660), .B(n1494), .Z(n1495) );
  XNOR U2339 ( .A(n4733), .B(n1495), .Z(out[1176]) );
  XOR U2340 ( .A(n1497), .B(n1496), .Z(n3848) );
  XNOR U2341 ( .A(in[965]), .B(n3848), .Z(n4737) );
  NAND U2342 ( .A(n1662), .B(n1498), .Z(n1499) );
  XNOR U2343 ( .A(n4737), .B(n1499), .Z(out[1177]) );
  XOR U2344 ( .A(n1501), .B(n1500), .Z(n3850) );
  XNOR U2345 ( .A(in[966]), .B(n3850), .Z(n4741) );
  NAND U2346 ( .A(n1664), .B(n1502), .Z(n1503) );
  XNOR U2347 ( .A(n4741), .B(n1503), .Z(out[1178]) );
  XOR U2348 ( .A(n1505), .B(n1504), .Z(n3852) );
  XNOR U2349 ( .A(in[967]), .B(n3852), .Z(n4745) );
  NAND U2350 ( .A(n1666), .B(n1506), .Z(n1507) );
  XNOR U2351 ( .A(n4745), .B(n1507), .Z(out[1179]) );
  XOR U2352 ( .A(in[588]), .B(n3668), .Z(n2586) );
  XOR U2353 ( .A(in[243]), .B(n3765), .Z(n3165) );
  XNOR U2354 ( .A(in[1463]), .B(n3808), .Z(n3162) );
  NAND U2355 ( .A(n3165), .B(n3162), .Z(n1508) );
  XNOR U2356 ( .A(n2586), .B(n1508), .Z(out[117]) );
  XOR U2357 ( .A(n1510), .B(n1509), .Z(n3856) );
  XNOR U2358 ( .A(in[968]), .B(n3856), .Z(n4749) );
  NAND U2359 ( .A(n1668), .B(n1511), .Z(n1512) );
  XNOR U2360 ( .A(n4749), .B(n1512), .Z(out[1180]) );
  XOR U2361 ( .A(n1514), .B(n1513), .Z(n3858) );
  XNOR U2362 ( .A(in[969]), .B(n3858), .Z(n4753) );
  NAND U2363 ( .A(n1670), .B(n1515), .Z(n1516) );
  XNOR U2364 ( .A(n4753), .B(n1516), .Z(out[1181]) );
  XNOR U2365 ( .A(n1518), .B(n1517), .Z(n3860) );
  XNOR U2366 ( .A(in[970]), .B(n3860), .Z(n4761) );
  NAND U2367 ( .A(n1672), .B(n1519), .Z(n1520) );
  XNOR U2368 ( .A(n4761), .B(n1520), .Z(out[1182]) );
  XOR U2369 ( .A(n1522), .B(n1521), .Z(n3862) );
  XNOR U2370 ( .A(in[971]), .B(n3862), .Z(n4765) );
  NAND U2371 ( .A(n1674), .B(n1523), .Z(n1524) );
  XNOR U2372 ( .A(n4765), .B(n1524), .Z(out[1183]) );
  XOR U2373 ( .A(n1526), .B(n1525), .Z(n3864) );
  XNOR U2374 ( .A(in[972]), .B(n3864), .Z(n4769) );
  NAND U2375 ( .A(n1676), .B(n1527), .Z(n1528) );
  XNOR U2376 ( .A(n4769), .B(n1528), .Z(out[1184]) );
  XOR U2377 ( .A(n1530), .B(n1529), .Z(n3866) );
  XNOR U2378 ( .A(in[973]), .B(n3866), .Z(n4773) );
  NAND U2379 ( .A(n1678), .B(n1531), .Z(n1532) );
  XNOR U2380 ( .A(n4773), .B(n1532), .Z(out[1185]) );
  XOR U2381 ( .A(n1534), .B(n1533), .Z(n3868) );
  XNOR U2382 ( .A(in[974]), .B(n3868), .Z(n4777) );
  NAND U2383 ( .A(n1681), .B(n1535), .Z(n1536) );
  XNOR U2384 ( .A(n4777), .B(n1536), .Z(out[1186]) );
  XNOR U2385 ( .A(n1538), .B(n1537), .Z(n3870) );
  XNOR U2386 ( .A(in[975]), .B(n3870), .Z(n4781) );
  NAND U2387 ( .A(n1683), .B(n1539), .Z(n1540) );
  XNOR U2388 ( .A(n4781), .B(n1540), .Z(out[1187]) );
  XNOR U2389 ( .A(n1542), .B(n1541), .Z(n3872) );
  XNOR U2390 ( .A(in[976]), .B(n3872), .Z(n4785) );
  NAND U2391 ( .A(n1685), .B(n1543), .Z(n1544) );
  XNOR U2392 ( .A(n4785), .B(n1544), .Z(out[1188]) );
  XOR U2393 ( .A(n1546), .B(n1545), .Z(n3874) );
  XNOR U2394 ( .A(in[977]), .B(n3874), .Z(n4789) );
  NAND U2395 ( .A(n1687), .B(n1547), .Z(n1548) );
  XNOR U2396 ( .A(n4789), .B(n1548), .Z(out[1189]) );
  XOR U2397 ( .A(in[589]), .B(n3672), .Z(n2588) );
  XOR U2398 ( .A(in[244]), .B(n3769), .Z(n3189) );
  XNOR U2399 ( .A(in[1464]), .B(n3812), .Z(n3186) );
  NAND U2400 ( .A(n3189), .B(n3186), .Z(n1549) );
  XNOR U2401 ( .A(n2588), .B(n1549), .Z(out[118]) );
  XOR U2402 ( .A(n1551), .B(n1550), .Z(n3878) );
  XNOR U2403 ( .A(in[978]), .B(n3878), .Z(n4793) );
  NAND U2404 ( .A(n1689), .B(n1552), .Z(n1553) );
  XNOR U2405 ( .A(n4793), .B(n1553), .Z(out[1190]) );
  XNOR U2406 ( .A(n1555), .B(n1554), .Z(n3880) );
  XNOR U2407 ( .A(in[979]), .B(n3880), .Z(n4797) );
  NAND U2408 ( .A(n1691), .B(n1556), .Z(n1557) );
  XNOR U2409 ( .A(n4797), .B(n1557), .Z(out[1191]) );
  OR U2410 ( .A(n1694), .B(n1558), .Z(n1559) );
  XNOR U2411 ( .A(n1693), .B(n1559), .Z(out[1192]) );
  OR U2412 ( .A(n1698), .B(n1560), .Z(n1561) );
  XNOR U2413 ( .A(n1697), .B(n1561), .Z(out[1193]) );
  OR U2414 ( .A(n1702), .B(n1562), .Z(n1563) );
  XNOR U2415 ( .A(n1701), .B(n1563), .Z(out[1194]) );
  OR U2416 ( .A(n1706), .B(n1564), .Z(n1565) );
  XNOR U2417 ( .A(n1705), .B(n1565), .Z(out[1195]) );
  OR U2418 ( .A(n1711), .B(n1566), .Z(n1567) );
  XNOR U2419 ( .A(n1710), .B(n1567), .Z(out[1196]) );
  OR U2420 ( .A(n1715), .B(n1568), .Z(n1569) );
  XNOR U2421 ( .A(n1714), .B(n1569), .Z(out[1197]) );
  OR U2422 ( .A(n1719), .B(n1570), .Z(n1571) );
  XNOR U2423 ( .A(n1718), .B(n1571), .Z(out[1198]) );
  OR U2424 ( .A(n1723), .B(n1572), .Z(n1573) );
  XNOR U2425 ( .A(n1722), .B(n1573), .Z(out[1199]) );
  XOR U2426 ( .A(in[590]), .B(n3676), .Z(n2590) );
  XOR U2427 ( .A(in[245]), .B(n3773), .Z(n3213) );
  XNOR U2428 ( .A(in[1465]), .B(n3816), .Z(n3210) );
  NAND U2429 ( .A(n3213), .B(n3210), .Z(n1574) );
  XNOR U2430 ( .A(n2590), .B(n1574), .Z(out[119]) );
  XOR U2431 ( .A(in[201]), .B(n3581), .Z(n3945) );
  XNOR U2432 ( .A(in[1421]), .B(n3618), .Z(n3944) );
  XOR U2433 ( .A(in[1044]), .B(n4123), .Z(n2635) );
  NAND U2434 ( .A(n3944), .B(n2635), .Z(n1575) );
  XNOR U2435 ( .A(n3945), .B(n1575), .Z(out[11]) );
  OR U2436 ( .A(n1727), .B(n1576), .Z(n1577) );
  XNOR U2437 ( .A(n1726), .B(n1577), .Z(out[1200]) );
  OR U2438 ( .A(n1731), .B(n1578), .Z(n1579) );
  XNOR U2439 ( .A(n1730), .B(n1579), .Z(out[1201]) );
  OR U2440 ( .A(n1735), .B(n1580), .Z(n1581) );
  XNOR U2441 ( .A(n1734), .B(n1581), .Z(out[1202]) );
  OR U2442 ( .A(n1739), .B(n1582), .Z(n1583) );
  XNOR U2443 ( .A(n1738), .B(n1583), .Z(out[1203]) );
  OR U2444 ( .A(n1743), .B(n1584), .Z(n1585) );
  XNOR U2445 ( .A(n1742), .B(n1585), .Z(out[1204]) );
  OR U2446 ( .A(n1747), .B(n1586), .Z(n1587) );
  XNOR U2447 ( .A(n1746), .B(n1587), .Z(out[1205]) );
  OR U2448 ( .A(n1752), .B(n1588), .Z(n1589) );
  XNOR U2449 ( .A(n1751), .B(n1589), .Z(out[1206]) );
  OR U2450 ( .A(n1756), .B(n1590), .Z(n1591) );
  XNOR U2451 ( .A(n1755), .B(n1591), .Z(out[1207]) );
  OR U2452 ( .A(n1760), .B(n1592), .Z(n1593) );
  XNOR U2453 ( .A(n1759), .B(n1593), .Z(out[1208]) );
  OR U2454 ( .A(n1764), .B(n1594), .Z(n1595) );
  XNOR U2455 ( .A(n1763), .B(n1595), .Z(out[1209]) );
  XOR U2456 ( .A(in[591]), .B(n3680), .Z(n2592) );
  XOR U2457 ( .A(in[246]), .B(n3777), .Z(n3237) );
  XNOR U2458 ( .A(in[1466]), .B(n3538), .Z(n3234) );
  NAND U2459 ( .A(n3237), .B(n3234), .Z(n1596) );
  XNOR U2460 ( .A(n2592), .B(n1596), .Z(out[120]) );
  OR U2461 ( .A(n1768), .B(n1597), .Z(n1598) );
  XNOR U2462 ( .A(n1767), .B(n1598), .Z(out[1210]) );
  OR U2463 ( .A(n1772), .B(n1599), .Z(n1600) );
  XNOR U2464 ( .A(n1771), .B(n1600), .Z(out[1211]) );
  OR U2465 ( .A(n1776), .B(n1601), .Z(n1602) );
  XNOR U2466 ( .A(n1775), .B(n1602), .Z(out[1212]) );
  OR U2467 ( .A(n1780), .B(n1603), .Z(n1604) );
  XNOR U2468 ( .A(n1779), .B(n1604), .Z(out[1213]) );
  OR U2469 ( .A(n1784), .B(n1605), .Z(n1606) );
  XNOR U2470 ( .A(n1783), .B(n1606), .Z(out[1214]) );
  OR U2471 ( .A(n1788), .B(n1607), .Z(n1608) );
  XNOR U2472 ( .A(n1787), .B(n1608), .Z(out[1215]) );
  OR U2473 ( .A(n4629), .B(n1609), .Z(n1610) );
  XNOR U2474 ( .A(n4628), .B(n1610), .Z(out[1216]) );
  OR U2475 ( .A(n4633), .B(n1611), .Z(n1612) );
  XNOR U2476 ( .A(n4632), .B(n1612), .Z(out[1217]) );
  OR U2477 ( .A(n4637), .B(n1613), .Z(n1614) );
  XNOR U2478 ( .A(n4636), .B(n1614), .Z(out[1218]) );
  OR U2479 ( .A(n4641), .B(n1615), .Z(n1616) );
  XNOR U2480 ( .A(n4640), .B(n1616), .Z(out[1219]) );
  XOR U2481 ( .A(in[592]), .B(n3684), .Z(n2594) );
  XOR U2482 ( .A(in[247]), .B(n3781), .Z(n3269) );
  XNOR U2483 ( .A(in[1467]), .B(n3542), .Z(n3266) );
  NAND U2484 ( .A(n3269), .B(n3266), .Z(n1617) );
  XNOR U2485 ( .A(n2594), .B(n1617), .Z(out[121]) );
  OR U2486 ( .A(n4645), .B(n1618), .Z(n1619) );
  XNOR U2487 ( .A(n4644), .B(n1619), .Z(out[1220]) );
  OR U2488 ( .A(n4649), .B(n1620), .Z(n1621) );
  XNOR U2489 ( .A(n4648), .B(n1621), .Z(out[1221]) );
  OR U2490 ( .A(n4653), .B(n1622), .Z(n1623) );
  XNOR U2491 ( .A(n4652), .B(n1623), .Z(out[1222]) );
  OR U2492 ( .A(n4657), .B(n1624), .Z(n1625) );
  XNOR U2493 ( .A(n4656), .B(n1625), .Z(out[1223]) );
  OR U2494 ( .A(n4661), .B(n1626), .Z(n1627) );
  XNOR U2495 ( .A(n4660), .B(n1627), .Z(out[1224]) );
  OR U2496 ( .A(n4665), .B(n1628), .Z(n1629) );
  XNOR U2497 ( .A(n4664), .B(n1629), .Z(out[1225]) );
  OR U2498 ( .A(n4673), .B(n1630), .Z(n1631) );
  XNOR U2499 ( .A(n4672), .B(n1631), .Z(out[1226]) );
  OR U2500 ( .A(n4677), .B(n1632), .Z(n1633) );
  XNOR U2501 ( .A(n4676), .B(n1633), .Z(out[1227]) );
  OR U2502 ( .A(n4681), .B(n1634), .Z(n1635) );
  XNOR U2503 ( .A(n4680), .B(n1635), .Z(out[1228]) );
  OR U2504 ( .A(n4685), .B(n1636), .Z(n1637) );
  XNOR U2505 ( .A(n4684), .B(n1637), .Z(out[1229]) );
  XOR U2506 ( .A(in[593]), .B(n3688), .Z(n2597) );
  XOR U2507 ( .A(in[248]), .B(n3785), .Z(n3313) );
  XNOR U2508 ( .A(in[1468]), .B(n3546), .Z(n3310) );
  NAND U2509 ( .A(n3313), .B(n3310), .Z(n1638) );
  XNOR U2510 ( .A(n2597), .B(n1638), .Z(out[122]) );
  OR U2511 ( .A(n4689), .B(n1639), .Z(n1640) );
  XNOR U2512 ( .A(n4688), .B(n1640), .Z(out[1230]) );
  OR U2513 ( .A(n4693), .B(n1641), .Z(n1642) );
  XNOR U2514 ( .A(n4692), .B(n1642), .Z(out[1231]) );
  OR U2515 ( .A(n4697), .B(n1643), .Z(n1644) );
  XNOR U2516 ( .A(n4696), .B(n1644), .Z(out[1232]) );
  OR U2517 ( .A(n4701), .B(n1645), .Z(n1646) );
  XNOR U2518 ( .A(n4700), .B(n1646), .Z(out[1233]) );
  OR U2519 ( .A(n4705), .B(n1647), .Z(n1648) );
  XNOR U2520 ( .A(n4704), .B(n1648), .Z(out[1234]) );
  OR U2521 ( .A(n4709), .B(n1649), .Z(n1650) );
  XNOR U2522 ( .A(n4708), .B(n1650), .Z(out[1235]) );
  OR U2523 ( .A(n4717), .B(n1651), .Z(n1652) );
  XNOR U2524 ( .A(n4716), .B(n1652), .Z(out[1236]) );
  OR U2525 ( .A(n4721), .B(n1653), .Z(n1654) );
  XNOR U2526 ( .A(n4720), .B(n1654), .Z(out[1237]) );
  OR U2527 ( .A(n4725), .B(n1655), .Z(n1656) );
  XNOR U2528 ( .A(n4724), .B(n1656), .Z(out[1238]) );
  OR U2529 ( .A(n4729), .B(n1657), .Z(n1658) );
  XNOR U2530 ( .A(n4728), .B(n1658), .Z(out[1239]) );
  XOR U2531 ( .A(in[594]), .B(n3692), .Z(n2599) );
  XOR U2532 ( .A(in[249]), .B(n3789), .Z(n3357) );
  XNOR U2533 ( .A(in[1469]), .B(n3550), .Z(n3354) );
  NAND U2534 ( .A(n3357), .B(n3354), .Z(n1659) );
  XNOR U2535 ( .A(n2599), .B(n1659), .Z(out[123]) );
  OR U2536 ( .A(n4733), .B(n1660), .Z(n1661) );
  XNOR U2537 ( .A(n4732), .B(n1661), .Z(out[1240]) );
  OR U2538 ( .A(n4737), .B(n1662), .Z(n1663) );
  XNOR U2539 ( .A(n4736), .B(n1663), .Z(out[1241]) );
  OR U2540 ( .A(n4741), .B(n1664), .Z(n1665) );
  XNOR U2541 ( .A(n4740), .B(n1665), .Z(out[1242]) );
  OR U2542 ( .A(n4745), .B(n1666), .Z(n1667) );
  XNOR U2543 ( .A(n4744), .B(n1667), .Z(out[1243]) );
  OR U2544 ( .A(n4749), .B(n1668), .Z(n1669) );
  XNOR U2545 ( .A(n4748), .B(n1669), .Z(out[1244]) );
  OR U2546 ( .A(n4753), .B(n1670), .Z(n1671) );
  XNOR U2547 ( .A(n4752), .B(n1671), .Z(out[1245]) );
  OR U2548 ( .A(n4761), .B(n1672), .Z(n1673) );
  XNOR U2549 ( .A(n4760), .B(n1673), .Z(out[1246]) );
  OR U2550 ( .A(n4765), .B(n1674), .Z(n1675) );
  XNOR U2551 ( .A(n4764), .B(n1675), .Z(out[1247]) );
  OR U2552 ( .A(n4769), .B(n1676), .Z(n1677) );
  XNOR U2553 ( .A(n4768), .B(n1677), .Z(out[1248]) );
  OR U2554 ( .A(n4773), .B(n1678), .Z(n1679) );
  XNOR U2555 ( .A(n4772), .B(n1679), .Z(out[1249]) );
  XOR U2556 ( .A(in[595]), .B(n3696), .Z(n2601) );
  XOR U2557 ( .A(in[250]), .B(n3793), .Z(n3403) );
  XNOR U2558 ( .A(in[1470]), .B(n3554), .Z(n3400) );
  NAND U2559 ( .A(n3403), .B(n3400), .Z(n1680) );
  XNOR U2560 ( .A(n2601), .B(n1680), .Z(out[124]) );
  OR U2561 ( .A(n4777), .B(n1681), .Z(n1682) );
  XNOR U2562 ( .A(n4776), .B(n1682), .Z(out[1250]) );
  OR U2563 ( .A(n4781), .B(n1683), .Z(n1684) );
  XNOR U2564 ( .A(n4780), .B(n1684), .Z(out[1251]) );
  OR U2565 ( .A(n4785), .B(n1685), .Z(n1686) );
  XNOR U2566 ( .A(n4784), .B(n1686), .Z(out[1252]) );
  OR U2567 ( .A(n4789), .B(n1687), .Z(n1688) );
  XNOR U2568 ( .A(n4788), .B(n1688), .Z(out[1253]) );
  OR U2569 ( .A(n4793), .B(n1689), .Z(n1690) );
  XNOR U2570 ( .A(n4792), .B(n1690), .Z(out[1254]) );
  OR U2571 ( .A(n4797), .B(n1691), .Z(n1692) );
  XNOR U2572 ( .A(n4796), .B(n1692), .Z(out[1255]) );
  ANDN U2573 ( .B(n1694), .A(n1693), .Z(n1695) );
  XNOR U2574 ( .A(n1696), .B(n1695), .Z(out[1256]) );
  ANDN U2575 ( .B(n1698), .A(n1697), .Z(n1699) );
  XNOR U2576 ( .A(n1700), .B(n1699), .Z(out[1257]) );
  ANDN U2577 ( .B(n1702), .A(n1701), .Z(n1703) );
  XNOR U2578 ( .A(n1704), .B(n1703), .Z(out[1258]) );
  ANDN U2579 ( .B(n1706), .A(n1705), .Z(n1707) );
  XNOR U2580 ( .A(n1708), .B(n1707), .Z(out[1259]) );
  XOR U2581 ( .A(in[596]), .B(n3700), .Z(n2603) );
  XNOR U2582 ( .A(in[251]), .B(n3803), .Z(n3447) );
  XNOR U2583 ( .A(in[1471]), .B(n3558), .Z(n3444) );
  NAND U2584 ( .A(n3447), .B(n3444), .Z(n1709) );
  XNOR U2585 ( .A(n2603), .B(n1709), .Z(out[125]) );
  ANDN U2586 ( .B(n1711), .A(n1710), .Z(n1712) );
  XNOR U2587 ( .A(n1713), .B(n1712), .Z(out[1260]) );
  ANDN U2588 ( .B(n1715), .A(n1714), .Z(n1716) );
  XNOR U2589 ( .A(n1717), .B(n1716), .Z(out[1261]) );
  ANDN U2590 ( .B(n1719), .A(n1718), .Z(n1720) );
  XNOR U2591 ( .A(n1721), .B(n1720), .Z(out[1262]) );
  ANDN U2592 ( .B(n1723), .A(n1722), .Z(n1724) );
  XNOR U2593 ( .A(n1725), .B(n1724), .Z(out[1263]) );
  ANDN U2594 ( .B(n1727), .A(n1726), .Z(n1728) );
  XNOR U2595 ( .A(n1729), .B(n1728), .Z(out[1264]) );
  ANDN U2596 ( .B(n1731), .A(n1730), .Z(n1732) );
  XNOR U2597 ( .A(n1733), .B(n1732), .Z(out[1265]) );
  ANDN U2598 ( .B(n1735), .A(n1734), .Z(n1736) );
  XNOR U2599 ( .A(n1737), .B(n1736), .Z(out[1266]) );
  ANDN U2600 ( .B(n1739), .A(n1738), .Z(n1740) );
  XNOR U2601 ( .A(n1741), .B(n1740), .Z(out[1267]) );
  ANDN U2602 ( .B(n1743), .A(n1742), .Z(n1744) );
  XNOR U2603 ( .A(n1745), .B(n1744), .Z(out[1268]) );
  ANDN U2604 ( .B(n1747), .A(n1746), .Z(n1748) );
  XNOR U2605 ( .A(n1749), .B(n1748), .Z(out[1269]) );
  XOR U2606 ( .A(in[597]), .B(n3704), .Z(n2605) );
  XNOR U2607 ( .A(in[252]), .B(n3807), .Z(n3491) );
  XNOR U2608 ( .A(in[1408]), .B(n3562), .Z(n3488) );
  NAND U2609 ( .A(n3491), .B(n3488), .Z(n1750) );
  XNOR U2610 ( .A(n2605), .B(n1750), .Z(out[126]) );
  ANDN U2611 ( .B(n1752), .A(n1751), .Z(n1753) );
  XNOR U2612 ( .A(n1754), .B(n1753), .Z(out[1270]) );
  ANDN U2613 ( .B(n1756), .A(n1755), .Z(n1757) );
  XNOR U2614 ( .A(n1758), .B(n1757), .Z(out[1271]) );
  ANDN U2615 ( .B(n1760), .A(n1759), .Z(n1761) );
  XNOR U2616 ( .A(n1762), .B(n1761), .Z(out[1272]) );
  ANDN U2617 ( .B(n1764), .A(n1763), .Z(n1765) );
  XNOR U2618 ( .A(n1766), .B(n1765), .Z(out[1273]) );
  ANDN U2619 ( .B(n1768), .A(n1767), .Z(n1769) );
  XNOR U2620 ( .A(n1770), .B(n1769), .Z(out[1274]) );
  ANDN U2621 ( .B(n1772), .A(n1771), .Z(n1773) );
  XNOR U2622 ( .A(n1774), .B(n1773), .Z(out[1275]) );
  ANDN U2623 ( .B(n1776), .A(n1775), .Z(n1777) );
  XNOR U2624 ( .A(n1778), .B(n1777), .Z(out[1276]) );
  ANDN U2625 ( .B(n1780), .A(n1779), .Z(n1781) );
  XNOR U2626 ( .A(n1782), .B(n1781), .Z(out[1277]) );
  ANDN U2627 ( .B(n1784), .A(n1783), .Z(n1785) );
  XNOR U2628 ( .A(n1786), .B(n1785), .Z(out[1278]) );
  ANDN U2629 ( .B(n1788), .A(n1787), .Z(n1789) );
  XNOR U2630 ( .A(n1790), .B(n1789), .Z(out[1279]) );
  XOR U2631 ( .A(in[598]), .B(n3712), .Z(n2607) );
  XNOR U2632 ( .A(in[253]), .B(n3811), .Z(n3535) );
  XNOR U2633 ( .A(in[1409]), .B(n3566), .Z(n3532) );
  NAND U2634 ( .A(n3535), .B(n3532), .Z(n1791) );
  XNOR U2635 ( .A(n2607), .B(n1791), .Z(out[127]) );
  XNOR U2636 ( .A(in[50]), .B(n3952), .Z(n1934) );
  XOR U2637 ( .A(in[1536]), .B(n3612), .Z(n2206) );
  XNOR U2638 ( .A(in[1172]), .B(n3629), .Z(n2204) );
  NAND U2639 ( .A(n2206), .B(n2204), .Z(n1792) );
  XNOR U2640 ( .A(n1934), .B(n1792), .Z(out[1280]) );
  XNOR U2641 ( .A(in[51]), .B(n3954), .Z(n1936) );
  XOR U2642 ( .A(in[1537]), .B(n3616), .Z(n2211) );
  XNOR U2643 ( .A(in[1173]), .B(n3633), .Z(n2209) );
  NAND U2644 ( .A(n2211), .B(n2209), .Z(n1793) );
  XNOR U2645 ( .A(n1936), .B(n1793), .Z(out[1281]) );
  XNOR U2646 ( .A(in[52]), .B(n3956), .Z(n1939) );
  XOR U2647 ( .A(in[1538]), .B(n3624), .Z(n2217) );
  XNOR U2648 ( .A(in[1174]), .B(n3637), .Z(n2214) );
  NAND U2649 ( .A(n2217), .B(n2214), .Z(n1794) );
  XNOR U2650 ( .A(n1939), .B(n1794), .Z(out[1282]) );
  XNOR U2651 ( .A(in[53]), .B(n3958), .Z(n1941) );
  XOR U2652 ( .A(in[1539]), .B(n3628), .Z(n2220) );
  XNOR U2653 ( .A(in[1175]), .B(n3641), .Z(n2218) );
  NAND U2654 ( .A(n2220), .B(n2218), .Z(n1795) );
  XNOR U2655 ( .A(n1941), .B(n1795), .Z(out[1283]) );
  XNOR U2656 ( .A(in[54]), .B(n3960), .Z(n1943) );
  XNOR U2657 ( .A(in[1540]), .B(n3632), .Z(n2227) );
  XNOR U2658 ( .A(in[1176]), .B(n3645), .Z(n2224) );
  NAND U2659 ( .A(n2227), .B(n2224), .Z(n1796) );
  XNOR U2660 ( .A(n1943), .B(n1796), .Z(out[1284]) );
  XNOR U2661 ( .A(in[55]), .B(n3962), .Z(n1945) );
  XNOR U2662 ( .A(in[1541]), .B(n3636), .Z(n2231) );
  XNOR U2663 ( .A(in[1177]), .B(n3649), .Z(n2228) );
  NAND U2664 ( .A(n2231), .B(n2228), .Z(n1797) );
  XNOR U2665 ( .A(n1945), .B(n1797), .Z(out[1285]) );
  XNOR U2666 ( .A(in[56]), .B(n3818), .Z(n1947) );
  XNOR U2667 ( .A(in[1542]), .B(n3640), .Z(n2235) );
  XNOR U2668 ( .A(in[1178]), .B(n3653), .Z(n2232) );
  NAND U2669 ( .A(n2235), .B(n2232), .Z(n1798) );
  XNOR U2670 ( .A(n1947), .B(n1798), .Z(out[1286]) );
  XNOR U2671 ( .A(in[57]), .B(n3820), .Z(n1949) );
  XNOR U2672 ( .A(in[1543]), .B(n3644), .Z(n2238) );
  XNOR U2673 ( .A(in[1179]), .B(n3657), .Z(n2236) );
  NAND U2674 ( .A(n2238), .B(n2236), .Z(n1799) );
  XNOR U2675 ( .A(n1949), .B(n1799), .Z(out[1287]) );
  XNOR U2676 ( .A(in[58]), .B(n3822), .Z(n1951) );
  XNOR U2677 ( .A(in[1544]), .B(n3648), .Z(n2244) );
  XNOR U2678 ( .A(in[1180]), .B(n3661), .Z(n2241) );
  NAND U2679 ( .A(n2244), .B(n2241), .Z(n1800) );
  XNOR U2680 ( .A(n1951), .B(n1800), .Z(out[1288]) );
  XNOR U2681 ( .A(in[59]), .B(n3824), .Z(n1953) );
  XNOR U2682 ( .A(in[1545]), .B(n3652), .Z(n2248) );
  XNOR U2683 ( .A(in[1181]), .B(n3669), .Z(n2245) );
  NAND U2684 ( .A(n2248), .B(n2245), .Z(n1801) );
  XNOR U2685 ( .A(n1953), .B(n1801), .Z(out[1289]) );
  XNOR U2686 ( .A(in[665]), .B(n3892), .Z(n2610) );
  XNOR U2687 ( .A(in[599]), .B(n3716), .Z(n3579) );
  NAND U2688 ( .A(n3579), .B(n3577), .Z(n1802) );
  XNOR U2689 ( .A(n2610), .B(n1802), .Z(out[128]) );
  XNOR U2690 ( .A(in[60]), .B(n3826), .Z(n1955) );
  XNOR U2691 ( .A(in[1546]), .B(n3656), .Z(n2252) );
  XNOR U2692 ( .A(in[1182]), .B(n3673), .Z(n2249) );
  NAND U2693 ( .A(n2252), .B(n2249), .Z(n1803) );
  XNOR U2694 ( .A(n1955), .B(n1803), .Z(out[1290]) );
  XNOR U2695 ( .A(in[61]), .B(n3828), .Z(n1957) );
  XNOR U2696 ( .A(in[1547]), .B(n3660), .Z(n2256) );
  XNOR U2697 ( .A(in[1183]), .B(n3677), .Z(n2253) );
  NAND U2698 ( .A(n2256), .B(n2253), .Z(n1804) );
  XNOR U2699 ( .A(n1957), .B(n1804), .Z(out[1291]) );
  XNOR U2700 ( .A(in[62]), .B(n3834), .Z(n1960) );
  XNOR U2701 ( .A(in[1548]), .B(n3668), .Z(n2260) );
  XNOR U2702 ( .A(in[1184]), .B(n3681), .Z(n2257) );
  NAND U2703 ( .A(n2260), .B(n2257), .Z(n1805) );
  XNOR U2704 ( .A(n1960), .B(n1805), .Z(out[1292]) );
  XNOR U2705 ( .A(in[63]), .B(n3836), .Z(n1962) );
  XNOR U2706 ( .A(in[1549]), .B(n3672), .Z(n2264) );
  XNOR U2707 ( .A(in[1185]), .B(n3685), .Z(n2261) );
  NAND U2708 ( .A(n2264), .B(n2261), .Z(n1806) );
  XNOR U2709 ( .A(n1962), .B(n1806), .Z(out[1293]) );
  XNOR U2710 ( .A(in[0]), .B(n3838), .Z(n1964) );
  XNOR U2711 ( .A(in[1550]), .B(n3676), .Z(n2269) );
  XOR U2712 ( .A(n3689), .B(in[1186]), .Z(n2266) );
  NAND U2713 ( .A(n2269), .B(n2266), .Z(n1807) );
  XNOR U2714 ( .A(n1964), .B(n1807), .Z(out[1294]) );
  XNOR U2715 ( .A(in[1]), .B(n3840), .Z(n1966) );
  XNOR U2716 ( .A(in[1551]), .B(n3680), .Z(n2272) );
  XOR U2717 ( .A(n3693), .B(in[1187]), .Z(n2270) );
  NAND U2718 ( .A(n2272), .B(n2270), .Z(n1808) );
  XNOR U2719 ( .A(n1966), .B(n1808), .Z(out[1295]) );
  XNOR U2720 ( .A(in[2]), .B(n3842), .Z(n1968) );
  XNOR U2721 ( .A(in[1552]), .B(n3684), .Z(n2278) );
  XOR U2722 ( .A(n3697), .B(in[1188]), .Z(n2275) );
  NAND U2723 ( .A(n2278), .B(n2275), .Z(n1809) );
  XNOR U2724 ( .A(n1968), .B(n1809), .Z(out[1296]) );
  XNOR U2725 ( .A(in[3]), .B(n3844), .Z(n1970) );
  XNOR U2726 ( .A(in[1553]), .B(n3688), .Z(n2282) );
  XOR U2727 ( .A(n3701), .B(in[1189]), .Z(n2279) );
  NAND U2728 ( .A(n2282), .B(n2279), .Z(n1810) );
  XNOR U2729 ( .A(n1970), .B(n1810), .Z(out[1297]) );
  XNOR U2730 ( .A(in[4]), .B(n3846), .Z(n1972) );
  XNOR U2731 ( .A(in[1554]), .B(n3692), .Z(n2286) );
  XNOR U2732 ( .A(in[1190]), .B(n3705), .Z(n2283) );
  NAND U2733 ( .A(n2286), .B(n2283), .Z(n1811) );
  XNOR U2734 ( .A(n1972), .B(n1811), .Z(out[1298]) );
  XNOR U2735 ( .A(in[5]), .B(n3848), .Z(n1974) );
  XNOR U2736 ( .A(in[1555]), .B(n3696), .Z(n2290) );
  XNOR U2737 ( .A(in[1191]), .B(n3713), .Z(n2287) );
  NAND U2738 ( .A(n2290), .B(n2287), .Z(n1812) );
  XNOR U2739 ( .A(n1974), .B(n1812), .Z(out[1299]) );
  XNOR U2740 ( .A(in[666]), .B(n3894), .Z(n2612) );
  XNOR U2741 ( .A(in[600]), .B(n3720), .Z(n3623) );
  XOR U2742 ( .A(in[255]), .B(n3537), .Z(n3621) );
  NAND U2743 ( .A(n3623), .B(n3621), .Z(n1813) );
  XNOR U2744 ( .A(n2612), .B(n1813), .Z(out[129]) );
  XOR U2745 ( .A(in[202]), .B(n3585), .Z(n3971) );
  XNOR U2746 ( .A(in[1422]), .B(n3626), .Z(n3970) );
  XOR U2747 ( .A(in[1045]), .B(n4126), .Z(n2638) );
  NAND U2748 ( .A(n3970), .B(n2638), .Z(n1814) );
  XNOR U2749 ( .A(n3971), .B(n1814), .Z(out[12]) );
  XNOR U2750 ( .A(in[6]), .B(n3850), .Z(n1976) );
  XNOR U2751 ( .A(in[1556]), .B(n3700), .Z(n2294) );
  XNOR U2752 ( .A(in[1192]), .B(n3717), .Z(n2291) );
  NAND U2753 ( .A(n2294), .B(n2291), .Z(n1815) );
  XNOR U2754 ( .A(n1976), .B(n1815), .Z(out[1300]) );
  XNOR U2755 ( .A(in[7]), .B(n3852), .Z(n1978) );
  XNOR U2756 ( .A(in[1557]), .B(n3704), .Z(n2298) );
  XNOR U2757 ( .A(in[1193]), .B(n3721), .Z(n2295) );
  NAND U2758 ( .A(n2298), .B(n2295), .Z(n1816) );
  XNOR U2759 ( .A(n1978), .B(n1816), .Z(out[1301]) );
  XNOR U2760 ( .A(in[8]), .B(n3856), .Z(n1981) );
  XNOR U2761 ( .A(in[1558]), .B(n3712), .Z(n2302) );
  XNOR U2762 ( .A(in[1194]), .B(n3725), .Z(n2299) );
  NAND U2763 ( .A(n2302), .B(n2299), .Z(n1817) );
  XNOR U2764 ( .A(n1981), .B(n1817), .Z(out[1302]) );
  XNOR U2765 ( .A(in[9]), .B(n3858), .Z(n1983) );
  XNOR U2766 ( .A(in[1559]), .B(n3716), .Z(n2306) );
  XNOR U2767 ( .A(in[1195]), .B(n3729), .Z(n2303) );
  NAND U2768 ( .A(n2306), .B(n2303), .Z(n1818) );
  XNOR U2769 ( .A(n1983), .B(n1818), .Z(out[1303]) );
  XNOR U2770 ( .A(in[10]), .B(n3860), .Z(n1985) );
  XNOR U2771 ( .A(in[1560]), .B(n3720), .Z(n2311) );
  XNOR U2772 ( .A(in[1196]), .B(n3733), .Z(n2308) );
  NAND U2773 ( .A(n2311), .B(n2308), .Z(n1819) );
  XNOR U2774 ( .A(n1985), .B(n1819), .Z(out[1304]) );
  XNOR U2775 ( .A(in[11]), .B(n3862), .Z(n1987) );
  XNOR U2776 ( .A(in[1561]), .B(n3724), .Z(n2315) );
  XNOR U2777 ( .A(in[1197]), .B(n3737), .Z(n2312) );
  NAND U2778 ( .A(n2315), .B(n2312), .Z(n1820) );
  XNOR U2779 ( .A(n1987), .B(n1820), .Z(out[1305]) );
  XNOR U2780 ( .A(in[12]), .B(n3864), .Z(n1989) );
  XNOR U2781 ( .A(in[1562]), .B(n3728), .Z(n2319) );
  XNOR U2782 ( .A(in[1198]), .B(n3741), .Z(n2316) );
  NAND U2783 ( .A(n2319), .B(n2316), .Z(n1821) );
  XNOR U2784 ( .A(n1989), .B(n1821), .Z(out[1306]) );
  XNOR U2785 ( .A(in[13]), .B(n3866), .Z(n1991) );
  XNOR U2786 ( .A(in[1563]), .B(n3732), .Z(n2323) );
  XNOR U2787 ( .A(in[1199]), .B(n3745), .Z(n2320) );
  NAND U2788 ( .A(n2323), .B(n2320), .Z(n1822) );
  XNOR U2789 ( .A(n1991), .B(n1822), .Z(out[1307]) );
  XNOR U2790 ( .A(in[14]), .B(n3868), .Z(n1993) );
  XNOR U2791 ( .A(in[1564]), .B(n3736), .Z(n2327) );
  XNOR U2792 ( .A(in[1200]), .B(n3749), .Z(n2324) );
  NAND U2793 ( .A(n2327), .B(n2324), .Z(n1823) );
  XNOR U2794 ( .A(n1993), .B(n1823), .Z(out[1308]) );
  XNOR U2795 ( .A(in[15]), .B(n3870), .Z(n1995) );
  XNOR U2796 ( .A(in[1565]), .B(n3740), .Z(n2331) );
  XNOR U2797 ( .A(in[1201]), .B(n3757), .Z(n2328) );
  NAND U2798 ( .A(n2331), .B(n2328), .Z(n1824) );
  XNOR U2799 ( .A(n1995), .B(n1824), .Z(out[1309]) );
  XNOR U2800 ( .A(in[667]), .B(n3896), .Z(n2615) );
  XNOR U2801 ( .A(in[601]), .B(n3724), .Z(n3667) );
  XOR U2802 ( .A(in[192]), .B(n3541), .Z(n3664) );
  NAND U2803 ( .A(n3667), .B(n3664), .Z(n1825) );
  XNOR U2804 ( .A(n2615), .B(n1825), .Z(out[130]) );
  XNOR U2805 ( .A(in[16]), .B(n3872), .Z(n1997) );
  XNOR U2806 ( .A(in[1566]), .B(n3744), .Z(n2335) );
  XNOR U2807 ( .A(in[1202]), .B(n3761), .Z(n2332) );
  NAND U2808 ( .A(n2335), .B(n2332), .Z(n1826) );
  XNOR U2809 ( .A(n1997), .B(n1826), .Z(out[1310]) );
  XNOR U2810 ( .A(in[17]), .B(n3874), .Z(n1999) );
  XNOR U2811 ( .A(in[1567]), .B(n3748), .Z(n2338) );
  XNOR U2812 ( .A(in[1203]), .B(n3765), .Z(n2336) );
  NAND U2813 ( .A(n2338), .B(n2336), .Z(n1827) );
  XNOR U2814 ( .A(n1999), .B(n1827), .Z(out[1311]) );
  XNOR U2815 ( .A(in[18]), .B(n3878), .Z(n2002) );
  XNOR U2816 ( .A(in[1568]), .B(n3756), .Z(n2344) );
  XNOR U2817 ( .A(in[1204]), .B(n3769), .Z(n2341) );
  NAND U2818 ( .A(n2344), .B(n2341), .Z(n1828) );
  XNOR U2819 ( .A(n2002), .B(n1828), .Z(out[1312]) );
  XNOR U2820 ( .A(in[19]), .B(n3880), .Z(n2004) );
  XNOR U2821 ( .A(in[1569]), .B(n3760), .Z(n2348) );
  XNOR U2822 ( .A(in[1205]), .B(n3773), .Z(n2345) );
  NAND U2823 ( .A(n2348), .B(n2345), .Z(n1829) );
  XNOR U2824 ( .A(n2004), .B(n1829), .Z(out[1313]) );
  XNOR U2825 ( .A(in[20]), .B(n3882), .Z(n2006) );
  XNOR U2826 ( .A(in[1570]), .B(n3764), .Z(n2353) );
  XNOR U2827 ( .A(in[1206]), .B(n3777), .Z(n2350) );
  NAND U2828 ( .A(n2353), .B(n2350), .Z(n1830) );
  XNOR U2829 ( .A(n2006), .B(n1830), .Z(out[1314]) );
  XNOR U2830 ( .A(in[21]), .B(n3884), .Z(n2008) );
  XNOR U2831 ( .A(in[1571]), .B(n3768), .Z(n2357) );
  XNOR U2832 ( .A(in[1207]), .B(n3781), .Z(n2354) );
  NAND U2833 ( .A(n2357), .B(n2354), .Z(n1831) );
  XNOR U2834 ( .A(n2008), .B(n1831), .Z(out[1315]) );
  XNOR U2835 ( .A(in[22]), .B(n3886), .Z(n2010) );
  XNOR U2836 ( .A(in[1572]), .B(n3772), .Z(n2361) );
  XNOR U2837 ( .A(in[1208]), .B(n3785), .Z(n2358) );
  NAND U2838 ( .A(n2361), .B(n2358), .Z(n1832) );
  XNOR U2839 ( .A(n2010), .B(n1832), .Z(out[1316]) );
  XNOR U2840 ( .A(in[23]), .B(n3888), .Z(n2012) );
  XOR U2841 ( .A(in[1573]), .B(n3776), .Z(n2365) );
  XNOR U2842 ( .A(in[1209]), .B(n3789), .Z(n2362) );
  NAND U2843 ( .A(n2365), .B(n2362), .Z(n1833) );
  XNOR U2844 ( .A(n2012), .B(n1833), .Z(out[1317]) );
  XNOR U2845 ( .A(in[24]), .B(n3890), .Z(n2014) );
  XOR U2846 ( .A(in[1574]), .B(n3780), .Z(n2369) );
  XNOR U2847 ( .A(in[1210]), .B(n3793), .Z(n2366) );
  NAND U2848 ( .A(n2369), .B(n2366), .Z(n1834) );
  XNOR U2849 ( .A(n2014), .B(n1834), .Z(out[1318]) );
  XNOR U2850 ( .A(in[25]), .B(n3892), .Z(n2016) );
  XOR U2851 ( .A(in[1575]), .B(n3784), .Z(n2373) );
  XOR U2852 ( .A(in[1211]), .B(n3803), .Z(n2370) );
  NAND U2853 ( .A(n2373), .B(n2370), .Z(n1835) );
  XNOR U2854 ( .A(n2016), .B(n1835), .Z(out[1319]) );
  XNOR U2855 ( .A(in[668]), .B(n3900), .Z(n2617) );
  XNOR U2856 ( .A(in[602]), .B(n3728), .Z(n3711) );
  XOR U2857 ( .A(in[193]), .B(n3545), .Z(n3708) );
  NAND U2858 ( .A(n3711), .B(n3708), .Z(n1836) );
  XNOR U2859 ( .A(n2617), .B(n1836), .Z(out[131]) );
  XNOR U2860 ( .A(in[26]), .B(n3894), .Z(n2018) );
  XOR U2861 ( .A(in[1576]), .B(n3788), .Z(n2377) );
  XOR U2862 ( .A(in[1212]), .B(n3807), .Z(n2374) );
  NAND U2863 ( .A(n2377), .B(n2374), .Z(n1837) );
  XNOR U2864 ( .A(n2018), .B(n1837), .Z(out[1320]) );
  XNOR U2865 ( .A(in[27]), .B(n3896), .Z(n2020) );
  XOR U2866 ( .A(in[1577]), .B(n3792), .Z(n2381) );
  XOR U2867 ( .A(in[1213]), .B(n3811), .Z(n2378) );
  NAND U2868 ( .A(n2381), .B(n2378), .Z(n1838) );
  XNOR U2869 ( .A(n2020), .B(n1838), .Z(out[1321]) );
  XNOR U2870 ( .A(in[28]), .B(n3900), .Z(n2023) );
  XOR U2871 ( .A(in[1578]), .B(n3802), .Z(n2385) );
  XNOR U2872 ( .A(in[1214]), .B(n3815), .Z(n2382) );
  NAND U2873 ( .A(n2385), .B(n2382), .Z(n1839) );
  XNOR U2874 ( .A(n2023), .B(n1839), .Z(out[1322]) );
  XNOR U2875 ( .A(in[29]), .B(n3902), .Z(n2025) );
  XOR U2876 ( .A(in[1579]), .B(n3806), .Z(n2389) );
  XOR U2877 ( .A(in[1215]), .B(n3537), .Z(n2386) );
  NAND U2878 ( .A(n2389), .B(n2386), .Z(n1840) );
  XNOR U2879 ( .A(n2025), .B(n1840), .Z(out[1323]) );
  XNOR U2880 ( .A(in[30]), .B(n3904), .Z(n2027) );
  XOR U2881 ( .A(in[1580]), .B(n3810), .Z(n2394) );
  XOR U2882 ( .A(in[1152]), .B(n3541), .Z(n2391) );
  NAND U2883 ( .A(n2394), .B(n2391), .Z(n1841) );
  XNOR U2884 ( .A(n2027), .B(n1841), .Z(out[1324]) );
  XNOR U2885 ( .A(in[31]), .B(n3906), .Z(n2029) );
  XOR U2886 ( .A(in[1581]), .B(n3814), .Z(n2398) );
  XOR U2887 ( .A(in[1153]), .B(n3545), .Z(n2395) );
  NAND U2888 ( .A(n2398), .B(n2395), .Z(n1842) );
  XNOR U2889 ( .A(n2029), .B(n1842), .Z(out[1325]) );
  XNOR U2890 ( .A(in[32]), .B(n3908), .Z(n2031) );
  XOR U2891 ( .A(in[1582]), .B(n3536), .Z(n2402) );
  XOR U2892 ( .A(in[1154]), .B(n3549), .Z(n2399) );
  NAND U2893 ( .A(n2402), .B(n2399), .Z(n1843) );
  XNOR U2894 ( .A(n2031), .B(n1843), .Z(out[1326]) );
  XNOR U2895 ( .A(in[33]), .B(n3910), .Z(n2033) );
  XOR U2896 ( .A(in[1583]), .B(n3540), .Z(n2406) );
  XOR U2897 ( .A(in[1155]), .B(n3553), .Z(n2403) );
  NAND U2898 ( .A(n2406), .B(n2403), .Z(n1844) );
  XNOR U2899 ( .A(n2033), .B(n1844), .Z(out[1327]) );
  XNOR U2900 ( .A(in[34]), .B(n3912), .Z(n2035) );
  XOR U2901 ( .A(in[1584]), .B(n3544), .Z(n2410) );
  XOR U2902 ( .A(in[1156]), .B(n3557), .Z(n2407) );
  NAND U2903 ( .A(n2410), .B(n2407), .Z(n1845) );
  XNOR U2904 ( .A(n2035), .B(n1845), .Z(out[1328]) );
  XNOR U2905 ( .A(in[35]), .B(n3914), .Z(n2037) );
  XOR U2906 ( .A(in[1585]), .B(n3548), .Z(n2414) );
  XOR U2907 ( .A(in[1157]), .B(n3561), .Z(n2411) );
  NAND U2908 ( .A(n2414), .B(n2411), .Z(n1846) );
  XNOR U2909 ( .A(n2037), .B(n1846), .Z(out[1329]) );
  XNOR U2910 ( .A(in[669]), .B(n3902), .Z(n2620) );
  XNOR U2911 ( .A(in[603]), .B(n3732), .Z(n3755) );
  XOR U2912 ( .A(in[194]), .B(n3549), .Z(n3752) );
  NAND U2913 ( .A(n3755), .B(n3752), .Z(n1847) );
  XNOR U2914 ( .A(n2620), .B(n1847), .Z(out[132]) );
  XNOR U2915 ( .A(in[36]), .B(n3916), .Z(n2039) );
  XOR U2916 ( .A(in[1586]), .B(n3552), .Z(n2418) );
  XOR U2917 ( .A(in[1158]), .B(n3565), .Z(n2415) );
  NAND U2918 ( .A(n2418), .B(n2415), .Z(n1848) );
  XNOR U2919 ( .A(n2039), .B(n1848), .Z(out[1330]) );
  XNOR U2920 ( .A(in[37]), .B(n3918), .Z(n2041) );
  XOR U2921 ( .A(in[1587]), .B(n3556), .Z(n2422) );
  XOR U2922 ( .A(in[1159]), .B(n3569), .Z(n2419) );
  NAND U2923 ( .A(n2422), .B(n2419), .Z(n1849) );
  XNOR U2924 ( .A(n2041), .B(n1849), .Z(out[1331]) );
  XNOR U2925 ( .A(in[38]), .B(n3924), .Z(n2044) );
  XOR U2926 ( .A(in[1588]), .B(n3560), .Z(n2426) );
  XOR U2927 ( .A(in[1160]), .B(n3573), .Z(n2423) );
  NAND U2928 ( .A(n2426), .B(n2423), .Z(n1850) );
  XNOR U2929 ( .A(n2044), .B(n1850), .Z(out[1332]) );
  XNOR U2930 ( .A(in[39]), .B(n3926), .Z(n2046) );
  XOR U2931 ( .A(in[1589]), .B(n3564), .Z(n2430) );
  XOR U2932 ( .A(in[1161]), .B(n3581), .Z(n2427) );
  NAND U2933 ( .A(n2430), .B(n2427), .Z(n1851) );
  XNOR U2934 ( .A(n2046), .B(n1851), .Z(out[1333]) );
  XNOR U2935 ( .A(in[40]), .B(n3928), .Z(n2048) );
  XOR U2936 ( .A(in[1590]), .B(n3568), .Z(n2435) );
  XOR U2937 ( .A(in[1162]), .B(n3585), .Z(n2432) );
  NAND U2938 ( .A(n2435), .B(n2432), .Z(n1852) );
  XNOR U2939 ( .A(n2048), .B(n1852), .Z(out[1334]) );
  XNOR U2940 ( .A(in[41]), .B(n3930), .Z(n2050) );
  XOR U2941 ( .A(in[1591]), .B(n3572), .Z(n2439) );
  XOR U2942 ( .A(in[1163]), .B(n3589), .Z(n2436) );
  NAND U2943 ( .A(n2439), .B(n2436), .Z(n1853) );
  XNOR U2944 ( .A(n2050), .B(n1853), .Z(out[1335]) );
  XNOR U2945 ( .A(in[42]), .B(n3932), .Z(n2052) );
  XOR U2946 ( .A(in[1592]), .B(n3580), .Z(n2443) );
  XOR U2947 ( .A(in[1164]), .B(n3593), .Z(n2440) );
  NAND U2948 ( .A(n2443), .B(n2440), .Z(n1854) );
  XNOR U2949 ( .A(n2052), .B(n1854), .Z(out[1336]) );
  XNOR U2950 ( .A(in[43]), .B(n3934), .Z(n2054) );
  XOR U2951 ( .A(in[1593]), .B(n3584), .Z(n2447) );
  XOR U2952 ( .A(in[1165]), .B(n3597), .Z(n2444) );
  NAND U2953 ( .A(n2447), .B(n2444), .Z(n1855) );
  XNOR U2954 ( .A(n2054), .B(n1855), .Z(out[1337]) );
  XNOR U2955 ( .A(in[44]), .B(n3936), .Z(n2056) );
  XOR U2956 ( .A(in[1594]), .B(n3588), .Z(n2451) );
  XOR U2957 ( .A(in[1166]), .B(n3601), .Z(n2448) );
  NAND U2958 ( .A(n2451), .B(n2448), .Z(n1856) );
  XNOR U2959 ( .A(n2056), .B(n1856), .Z(out[1338]) );
  XNOR U2960 ( .A(in[45]), .B(n3938), .Z(n2058) );
  XOR U2961 ( .A(in[1595]), .B(n3592), .Z(n2455) );
  XOR U2962 ( .A(in[1167]), .B(n3605), .Z(n2452) );
  NAND U2963 ( .A(n2455), .B(n2452), .Z(n1857) );
  XNOR U2964 ( .A(n2058), .B(n1857), .Z(out[1339]) );
  XNOR U2965 ( .A(in[670]), .B(n3904), .Z(n2622) );
  XNOR U2966 ( .A(in[604]), .B(n3736), .Z(n3799) );
  XOR U2967 ( .A(in[195]), .B(n3553), .Z(n3796) );
  NAND U2968 ( .A(n3799), .B(n3796), .Z(n1858) );
  XNOR U2969 ( .A(n2622), .B(n1858), .Z(out[133]) );
  XNOR U2970 ( .A(in[46]), .B(n3940), .Z(n2060) );
  XOR U2971 ( .A(in[1596]), .B(n3596), .Z(n2459) );
  XOR U2972 ( .A(in[1168]), .B(n3609), .Z(n2456) );
  NAND U2973 ( .A(n2459), .B(n2456), .Z(n1859) );
  XNOR U2974 ( .A(n2060), .B(n1859), .Z(out[1340]) );
  XNOR U2975 ( .A(in[47]), .B(n3942), .Z(n2062) );
  XOR U2976 ( .A(in[1597]), .B(n3600), .Z(n2463) );
  XOR U2977 ( .A(in[1169]), .B(n3613), .Z(n2460) );
  NAND U2978 ( .A(n2463), .B(n2460), .Z(n1860) );
  XNOR U2979 ( .A(n2062), .B(n1860), .Z(out[1341]) );
  XNOR U2980 ( .A(in[48]), .B(n3948), .Z(n2065) );
  XOR U2981 ( .A(in[1598]), .B(n3604), .Z(n2467) );
  XOR U2982 ( .A(in[1170]), .B(n3617), .Z(n2464) );
  NAND U2983 ( .A(n2467), .B(n2464), .Z(n1861) );
  XNOR U2984 ( .A(n2065), .B(n1861), .Z(out[1342]) );
  XNOR U2985 ( .A(in[49]), .B(n3950), .Z(n2067) );
  XOR U2986 ( .A(in[1599]), .B(n3608), .Z(n2470) );
  XNOR U2987 ( .A(in[1171]), .B(n3625), .Z(n2468) );
  NAND U2988 ( .A(n2470), .B(n2468), .Z(n1862) );
  XNOR U2989 ( .A(n2067), .B(n1862), .Z(out[1343]) );
  XOR U2990 ( .A(in[427]), .B(n3980), .Z(n2069) );
  NOR U2991 ( .A(n1934), .B(n2206), .Z(n1863) );
  XNOR U2992 ( .A(n2069), .B(n1863), .Z(out[1344]) );
  XOR U2993 ( .A(in[428]), .B(n3983), .Z(n2071) );
  NOR U2994 ( .A(n1936), .B(n2211), .Z(n1864) );
  XNOR U2995 ( .A(n2071), .B(n1864), .Z(out[1345]) );
  XOR U2996 ( .A(in[429]), .B(n3986), .Z(n2073) );
  NOR U2997 ( .A(n1939), .B(n2217), .Z(n1865) );
  XNOR U2998 ( .A(n2073), .B(n1865), .Z(out[1346]) );
  XOR U2999 ( .A(in[430]), .B(n3989), .Z(n2075) );
  NOR U3000 ( .A(n1941), .B(n2220), .Z(n1866) );
  XNOR U3001 ( .A(n2075), .B(n1866), .Z(out[1347]) );
  XOR U3002 ( .A(in[431]), .B(n3992), .Z(n2077) );
  NOR U3003 ( .A(n1943), .B(n2227), .Z(n1867) );
  XNOR U3004 ( .A(n2077), .B(n1867), .Z(out[1348]) );
  XOR U3005 ( .A(in[432]), .B(n3995), .Z(n2079) );
  NOR U3006 ( .A(n1945), .B(n2231), .Z(n1868) );
  XNOR U3007 ( .A(n2079), .B(n1868), .Z(out[1349]) );
  XNOR U3008 ( .A(in[671]), .B(n3906), .Z(n2624) );
  XNOR U3009 ( .A(in[605]), .B(n3740), .Z(n3833) );
  XOR U3010 ( .A(in[196]), .B(n3557), .Z(n3830) );
  NAND U3011 ( .A(n3833), .B(n3830), .Z(n1869) );
  XNOR U3012 ( .A(n2624), .B(n1869), .Z(out[134]) );
  XOR U3013 ( .A(in[433]), .B(n3998), .Z(n2081) );
  NOR U3014 ( .A(n1947), .B(n2235), .Z(n1870) );
  XNOR U3015 ( .A(n2081), .B(n1870), .Z(out[1350]) );
  XOR U3016 ( .A(in[434]), .B(n4001), .Z(n2083) );
  NOR U3017 ( .A(n1949), .B(n2238), .Z(n1871) );
  XNOR U3018 ( .A(n2083), .B(n1871), .Z(out[1351]) );
  XOR U3019 ( .A(in[435]), .B(n4008), .Z(n2086) );
  NOR U3020 ( .A(n1951), .B(n2244), .Z(n1872) );
  XNOR U3021 ( .A(n2086), .B(n1872), .Z(out[1352]) );
  XOR U3022 ( .A(in[436]), .B(n4011), .Z(n2088) );
  NOR U3023 ( .A(n1953), .B(n2248), .Z(n1873) );
  XNOR U3024 ( .A(n2088), .B(n1873), .Z(out[1353]) );
  XOR U3025 ( .A(in[437]), .B(n4014), .Z(n2090) );
  NOR U3026 ( .A(n1955), .B(n2252), .Z(n1874) );
  XNOR U3027 ( .A(n2090), .B(n1874), .Z(out[1354]) );
  XOR U3028 ( .A(in[438]), .B(n4017), .Z(n2092) );
  NOR U3029 ( .A(n1957), .B(n2256), .Z(n1875) );
  XNOR U3030 ( .A(n2092), .B(n1875), .Z(out[1355]) );
  XOR U3031 ( .A(in[439]), .B(n4020), .Z(n2094) );
  NOR U3032 ( .A(n1960), .B(n2260), .Z(n1876) );
  XNOR U3033 ( .A(n2094), .B(n1876), .Z(out[1356]) );
  XOR U3034 ( .A(in[440]), .B(n4023), .Z(n2096) );
  NOR U3035 ( .A(n1962), .B(n2264), .Z(n1877) );
  XNOR U3036 ( .A(n2096), .B(n1877), .Z(out[1357]) );
  XOR U3037 ( .A(in[441]), .B(n4026), .Z(n2098) );
  NOR U3038 ( .A(n1964), .B(n2269), .Z(n1878) );
  XNOR U3039 ( .A(n2098), .B(n1878), .Z(out[1358]) );
  XOR U3040 ( .A(in[442]), .B(n4029), .Z(n2100) );
  NOR U3041 ( .A(n1966), .B(n2272), .Z(n1879) );
  XNOR U3042 ( .A(n2100), .B(n1879), .Z(out[1359]) );
  XNOR U3043 ( .A(in[672]), .B(n3908), .Z(n2626) );
  XNOR U3044 ( .A(in[606]), .B(n3744), .Z(n3855) );
  XOR U3045 ( .A(in[197]), .B(n3561), .Z(n4079) );
  NAND U3046 ( .A(n3855), .B(n4079), .Z(n1880) );
  XNOR U3047 ( .A(n2626), .B(n1880), .Z(out[135]) );
  XOR U3048 ( .A(in[443]), .B(n4032), .Z(n2102) );
  NOR U3049 ( .A(n1968), .B(n2278), .Z(n1881) );
  XNOR U3050 ( .A(n2102), .B(n1881), .Z(out[1360]) );
  XOR U3051 ( .A(in[444]), .B(n4035), .Z(n2104) );
  NOR U3052 ( .A(n1970), .B(n2282), .Z(n1882) );
  XNOR U3053 ( .A(n2104), .B(n1882), .Z(out[1361]) );
  XOR U3054 ( .A(in[445]), .B(n4042), .Z(n2107) );
  NOR U3055 ( .A(n1972), .B(n2286), .Z(n1883) );
  XNOR U3056 ( .A(n2107), .B(n1883), .Z(out[1362]) );
  XOR U3057 ( .A(in[446]), .B(n4045), .Z(n2109) );
  NOR U3058 ( .A(n1974), .B(n2290), .Z(n1884) );
  XNOR U3059 ( .A(n2109), .B(n1884), .Z(out[1363]) );
  XOR U3060 ( .A(in[447]), .B(n4048), .Z(n2111) );
  NOR U3061 ( .A(n1976), .B(n2294), .Z(n1885) );
  XNOR U3062 ( .A(n2111), .B(n1885), .Z(out[1364]) );
  XOR U3063 ( .A(in[384]), .B(n4051), .Z(n2113) );
  NOR U3064 ( .A(n1978), .B(n2298), .Z(n1886) );
  XNOR U3065 ( .A(n2113), .B(n1886), .Z(out[1365]) );
  XOR U3066 ( .A(in[385]), .B(n4054), .Z(n2115) );
  NOR U3067 ( .A(n1981), .B(n2302), .Z(n1887) );
  XNOR U3068 ( .A(n2115), .B(n1887), .Z(out[1366]) );
  XOR U3069 ( .A(in[386]), .B(n4057), .Z(n2117) );
  NOR U3070 ( .A(n1983), .B(n2306), .Z(n1888) );
  XNOR U3071 ( .A(n2117), .B(n1888), .Z(out[1367]) );
  XOR U3072 ( .A(in[387]), .B(n4060), .Z(n2119) );
  NOR U3073 ( .A(n1985), .B(n2311), .Z(n1889) );
  XNOR U3074 ( .A(n2119), .B(n1889), .Z(out[1368]) );
  XOR U3075 ( .A(in[388]), .B(n4063), .Z(n2121) );
  NOR U3076 ( .A(n1987), .B(n2315), .Z(n1890) );
  XNOR U3077 ( .A(n2121), .B(n1890), .Z(out[1369]) );
  XNOR U3078 ( .A(in[673]), .B(n3910), .Z(n2628) );
  XNOR U3079 ( .A(in[607]), .B(n3748), .Z(n3877) );
  XOR U3080 ( .A(in[198]), .B(n3565), .Z(n4363) );
  NAND U3081 ( .A(n3877), .B(n4363), .Z(n1891) );
  XNOR U3082 ( .A(n2628), .B(n1891), .Z(out[136]) );
  XOR U3083 ( .A(in[389]), .B(n4066), .Z(n2123) );
  NOR U3084 ( .A(n1989), .B(n2319), .Z(n1892) );
  XNOR U3085 ( .A(n2123), .B(n1892), .Z(out[1370]) );
  XOR U3086 ( .A(in[390]), .B(n4069), .Z(n2125) );
  NOR U3087 ( .A(n1991), .B(n2323), .Z(n1893) );
  XNOR U3088 ( .A(n2125), .B(n1893), .Z(out[1371]) );
  XOR U3089 ( .A(in[391]), .B(n4080), .Z(n2129) );
  NOR U3090 ( .A(n1993), .B(n2327), .Z(n1894) );
  XNOR U3091 ( .A(n2129), .B(n1894), .Z(out[1372]) );
  XOR U3092 ( .A(in[392]), .B(n4083), .Z(n2131) );
  NOR U3093 ( .A(n1995), .B(n2331), .Z(n1895) );
  XNOR U3094 ( .A(n2131), .B(n1895), .Z(out[1373]) );
  XOR U3095 ( .A(in[393]), .B(n4086), .Z(n2133) );
  NOR U3096 ( .A(n1997), .B(n2335), .Z(n1896) );
  XNOR U3097 ( .A(n2133), .B(n1896), .Z(out[1374]) );
  XOR U3098 ( .A(in[394]), .B(n4089), .Z(n2135) );
  NOR U3099 ( .A(n1999), .B(n2338), .Z(n1897) );
  XNOR U3100 ( .A(n2135), .B(n1897), .Z(out[1375]) );
  XOR U3101 ( .A(in[395]), .B(n4092), .Z(n2137) );
  NOR U3102 ( .A(n2002), .B(n2344), .Z(n1898) );
  XNOR U3103 ( .A(n2137), .B(n1898), .Z(out[1376]) );
  XNOR U3104 ( .A(n4095), .B(in[396]), .Z(n2139) );
  NOR U3105 ( .A(n2004), .B(n2348), .Z(n1899) );
  XNOR U3106 ( .A(n2139), .B(n1899), .Z(out[1377]) );
  XNOR U3107 ( .A(n4098), .B(in[397]), .Z(n2141) );
  NOR U3108 ( .A(n2006), .B(n2353), .Z(n1900) );
  XNOR U3109 ( .A(n2141), .B(n1900), .Z(out[1378]) );
  XNOR U3110 ( .A(n4101), .B(in[398]), .Z(n2143) );
  NOR U3111 ( .A(n2008), .B(n2357), .Z(n1901) );
  XNOR U3112 ( .A(n2143), .B(n1901), .Z(out[1379]) );
  XNOR U3113 ( .A(in[674]), .B(n3912), .Z(n2630) );
  XNOR U3114 ( .A(in[608]), .B(n3756), .Z(n3899) );
  XOR U3115 ( .A(in[199]), .B(n3569), .Z(n4807) );
  NAND U3116 ( .A(n3899), .B(n4807), .Z(n1902) );
  XNOR U3117 ( .A(n2630), .B(n1902), .Z(out[137]) );
  XNOR U3118 ( .A(n4104), .B(in[399]), .Z(n2145) );
  NOR U3119 ( .A(n2010), .B(n2361), .Z(n1903) );
  XNOR U3120 ( .A(n2145), .B(n1903), .Z(out[1380]) );
  XNOR U3121 ( .A(n4107), .B(in[400]), .Z(n2147) );
  NOR U3122 ( .A(n2012), .B(n2365), .Z(n1904) );
  XNOR U3123 ( .A(n2147), .B(n1904), .Z(out[1381]) );
  XNOR U3124 ( .A(n4114), .B(in[401]), .Z(n2150) );
  NOR U3125 ( .A(n2014), .B(n2369), .Z(n1905) );
  XNOR U3126 ( .A(n2150), .B(n1905), .Z(out[1382]) );
  XNOR U3127 ( .A(n4117), .B(in[402]), .Z(n2152) );
  NOR U3128 ( .A(n2016), .B(n2373), .Z(n1906) );
  XNOR U3129 ( .A(n2152), .B(n1906), .Z(out[1383]) );
  XNOR U3130 ( .A(n4120), .B(in[403]), .Z(n2154) );
  NOR U3131 ( .A(n2018), .B(n2377), .Z(n1907) );
  XNOR U3132 ( .A(n2154), .B(n1907), .Z(out[1384]) );
  XNOR U3133 ( .A(in[404]), .B(n4123), .Z(n2156) );
  NOR U3134 ( .A(n2020), .B(n2381), .Z(n1908) );
  XNOR U3135 ( .A(n2156), .B(n1908), .Z(out[1385]) );
  XNOR U3136 ( .A(in[405]), .B(n4126), .Z(n2158) );
  NOR U3137 ( .A(n2023), .B(n2385), .Z(n1909) );
  XNOR U3138 ( .A(n2158), .B(n1909), .Z(out[1386]) );
  XNOR U3139 ( .A(in[406]), .B(n4129), .Z(n2160) );
  NOR U3140 ( .A(n2025), .B(n2389), .Z(n1910) );
  XNOR U3141 ( .A(n2160), .B(n1910), .Z(out[1387]) );
  XNOR U3142 ( .A(in[407]), .B(n4132), .Z(n2162) );
  NOR U3143 ( .A(n2027), .B(n2394), .Z(n1911) );
  XNOR U3144 ( .A(n2162), .B(n1911), .Z(out[1388]) );
  XNOR U3145 ( .A(in[408]), .B(n4135), .Z(n2164) );
  NOR U3146 ( .A(n2029), .B(n2398), .Z(n1912) );
  XNOR U3147 ( .A(n2164), .B(n1912), .Z(out[1389]) );
  XNOR U3148 ( .A(in[675]), .B(n3914), .Z(n2633) );
  XNOR U3149 ( .A(in[609]), .B(n3760), .Z(n3923) );
  NAND U3150 ( .A(n3923), .B(n3921), .Z(n1913) );
  XNOR U3151 ( .A(n2633), .B(n1913), .Z(out[138]) );
  XNOR U3152 ( .A(in[409]), .B(n4138), .Z(n2166) );
  NOR U3153 ( .A(n2031), .B(n2402), .Z(n1914) );
  XNOR U3154 ( .A(n2166), .B(n1914), .Z(out[1390]) );
  XNOR U3155 ( .A(in[410]), .B(n4141), .Z(n2168) );
  NOR U3156 ( .A(n2033), .B(n2406), .Z(n1915) );
  XNOR U3157 ( .A(n2168), .B(n1915), .Z(out[1391]) );
  XNOR U3158 ( .A(in[411]), .B(n4148), .Z(n2171) );
  NOR U3159 ( .A(n2035), .B(n2410), .Z(n1916) );
  XNOR U3160 ( .A(n2171), .B(n1916), .Z(out[1392]) );
  XNOR U3161 ( .A(in[412]), .B(n4151), .Z(n2173) );
  NOR U3162 ( .A(n2037), .B(n2414), .Z(n1917) );
  XNOR U3163 ( .A(n2173), .B(n1917), .Z(out[1393]) );
  XNOR U3164 ( .A(in[413]), .B(n4154), .Z(n2175) );
  NOR U3165 ( .A(n2039), .B(n2418), .Z(n1918) );
  XNOR U3166 ( .A(n2175), .B(n1918), .Z(out[1394]) );
  XNOR U3167 ( .A(in[414]), .B(n4157), .Z(n2177) );
  NOR U3168 ( .A(n2041), .B(n2422), .Z(n1919) );
  XNOR U3169 ( .A(n2177), .B(n1919), .Z(out[1395]) );
  XNOR U3170 ( .A(in[415]), .B(n4160), .Z(n2179) );
  NOR U3171 ( .A(n2044), .B(n2426), .Z(n1920) );
  XNOR U3172 ( .A(n2179), .B(n1920), .Z(out[1396]) );
  XNOR U3173 ( .A(in[416]), .B(n4163), .Z(n2181) );
  NOR U3174 ( .A(n2046), .B(n2430), .Z(n1921) );
  XNOR U3175 ( .A(n2181), .B(n1921), .Z(out[1397]) );
  XNOR U3176 ( .A(in[417]), .B(n4166), .Z(n2183) );
  NOR U3177 ( .A(n2048), .B(n2435), .Z(n1922) );
  XNOR U3178 ( .A(n2183), .B(n1922), .Z(out[1398]) );
  XNOR U3179 ( .A(in[418]), .B(n4169), .Z(n2185) );
  NOR U3180 ( .A(n2050), .B(n2439), .Z(n1923) );
  XNOR U3181 ( .A(n2185), .B(n1923), .Z(out[1399]) );
  XNOR U3182 ( .A(in[676]), .B(n3916), .Z(n2636) );
  XNOR U3183 ( .A(in[610]), .B(n3764), .Z(n3947) );
  NAND U3184 ( .A(n3947), .B(n3945), .Z(n1924) );
  XNOR U3185 ( .A(n2636), .B(n1924), .Z(out[139]) );
  XOR U3186 ( .A(in[203]), .B(n3589), .Z(n4005) );
  XNOR U3187 ( .A(in[1423]), .B(n3630), .Z(n4004) );
  XOR U3188 ( .A(in[1046]), .B(n4129), .Z(n2641) );
  NAND U3189 ( .A(n4004), .B(n2641), .Z(n1925) );
  XNOR U3190 ( .A(n4005), .B(n1925), .Z(out[13]) );
  XNOR U3191 ( .A(in[419]), .B(n4172), .Z(n2187) );
  NOR U3192 ( .A(n2052), .B(n2443), .Z(n1926) );
  XNOR U3193 ( .A(n2187), .B(n1926), .Z(out[1400]) );
  XOR U3194 ( .A(in[420]), .B(n4175), .Z(n2189) );
  NOR U3195 ( .A(n2054), .B(n2447), .Z(n1927) );
  XNOR U3196 ( .A(n2189), .B(n1927), .Z(out[1401]) );
  XOR U3197 ( .A(in[421]), .B(n4182), .Z(n2192) );
  NOR U3198 ( .A(n2056), .B(n2451), .Z(n1928) );
  XNOR U3199 ( .A(n2192), .B(n1928), .Z(out[1402]) );
  XOR U3200 ( .A(in[422]), .B(n4185), .Z(n2194) );
  NOR U3201 ( .A(n2058), .B(n2455), .Z(n1929) );
  XNOR U3202 ( .A(n2194), .B(n1929), .Z(out[1403]) );
  XOR U3203 ( .A(in[423]), .B(n3964), .Z(n2196) );
  NOR U3204 ( .A(n2060), .B(n2459), .Z(n1930) );
  XNOR U3205 ( .A(n2196), .B(n1930), .Z(out[1404]) );
  XOR U3206 ( .A(in[424]), .B(n3967), .Z(n2198) );
  NOR U3207 ( .A(n2062), .B(n2463), .Z(n1931) );
  XNOR U3208 ( .A(n2198), .B(n1931), .Z(out[1405]) );
  XOR U3209 ( .A(in[425]), .B(n3974), .Z(n2200) );
  NOR U3210 ( .A(n2065), .B(n2467), .Z(n1932) );
  XNOR U3211 ( .A(n2200), .B(n1932), .Z(out[1406]) );
  XOR U3212 ( .A(in[426]), .B(n3977), .Z(n2202) );
  NOR U3213 ( .A(n2067), .B(n2470), .Z(n1933) );
  XNOR U3214 ( .A(n2202), .B(n1933), .Z(out[1407]) );
  XOR U3215 ( .A(in[789]), .B(n3654), .Z(n2205) );
  NAND U3216 ( .A(n2069), .B(n1934), .Z(n1935) );
  XNOR U3217 ( .A(n2205), .B(n1935), .Z(out[1408]) );
  XOR U3218 ( .A(in[790]), .B(n3658), .Z(n2210) );
  NAND U3219 ( .A(n2071), .B(n1936), .Z(n1937) );
  XNOR U3220 ( .A(n2210), .B(n1937), .Z(out[1409]) );
  XNOR U3221 ( .A(in[677]), .B(n3918), .Z(n2639) );
  XNOR U3222 ( .A(in[611]), .B(n3768), .Z(n3973) );
  NAND U3223 ( .A(n3973), .B(n3971), .Z(n1938) );
  XNOR U3224 ( .A(n2639), .B(n1938), .Z(out[140]) );
  XOR U3225 ( .A(in[791]), .B(n3662), .Z(n2215) );
  NAND U3226 ( .A(n2073), .B(n1939), .Z(n1940) );
  XNOR U3227 ( .A(n2215), .B(n1940), .Z(out[1410]) );
  XOR U3228 ( .A(in[792]), .B(n3670), .Z(n2219) );
  NAND U3229 ( .A(n2075), .B(n1941), .Z(n1942) );
  XNOR U3230 ( .A(n2219), .B(n1942), .Z(out[1411]) );
  XOR U3231 ( .A(in[793]), .B(n3674), .Z(n2225) );
  NAND U3232 ( .A(n2077), .B(n1943), .Z(n1944) );
  XNOR U3233 ( .A(n2225), .B(n1944), .Z(out[1412]) );
  XOR U3234 ( .A(in[794]), .B(n3678), .Z(n2229) );
  NAND U3235 ( .A(n2079), .B(n1945), .Z(n1946) );
  XNOR U3236 ( .A(n2229), .B(n1946), .Z(out[1413]) );
  XOR U3237 ( .A(in[795]), .B(n3682), .Z(n2233) );
  NAND U3238 ( .A(n2081), .B(n1947), .Z(n1948) );
  XNOR U3239 ( .A(n2233), .B(n1948), .Z(out[1414]) );
  XOR U3240 ( .A(in[796]), .B(n3686), .Z(n2237) );
  NAND U3241 ( .A(n2083), .B(n1949), .Z(n1950) );
  XNOR U3242 ( .A(n2237), .B(n1950), .Z(out[1415]) );
  XOR U3243 ( .A(in[797]), .B(n3690), .Z(n2242) );
  NAND U3244 ( .A(n2086), .B(n1951), .Z(n1952) );
  XNOR U3245 ( .A(n2242), .B(n1952), .Z(out[1416]) );
  XOR U3246 ( .A(in[798]), .B(n3694), .Z(n2246) );
  NAND U3247 ( .A(n2088), .B(n1953), .Z(n1954) );
  XNOR U3248 ( .A(n2246), .B(n1954), .Z(out[1417]) );
  XOR U3249 ( .A(in[799]), .B(n3698), .Z(n2250) );
  NAND U3250 ( .A(n2090), .B(n1955), .Z(n1956) );
  XNOR U3251 ( .A(n2250), .B(n1956), .Z(out[1418]) );
  XOR U3252 ( .A(in[800]), .B(n3702), .Z(n2254) );
  NAND U3253 ( .A(n2092), .B(n1957), .Z(n1958) );
  XNOR U3254 ( .A(n2254), .B(n1958), .Z(out[1419]) );
  XNOR U3255 ( .A(in[678]), .B(n3924), .Z(n2642) );
  XNOR U3256 ( .A(in[612]), .B(n3772), .Z(n4007) );
  NAND U3257 ( .A(n4007), .B(n4005), .Z(n1959) );
  XNOR U3258 ( .A(n2642), .B(n1959), .Z(out[141]) );
  XOR U3259 ( .A(in[801]), .B(n3706), .Z(n2258) );
  NAND U3260 ( .A(n2094), .B(n1960), .Z(n1961) );
  XNOR U3261 ( .A(n2258), .B(n1961), .Z(out[1420]) );
  XOR U3262 ( .A(in[802]), .B(n3714), .Z(n2262) );
  NAND U3263 ( .A(n2096), .B(n1962), .Z(n1963) );
  XNOR U3264 ( .A(n2262), .B(n1963), .Z(out[1421]) );
  XOR U3265 ( .A(in[803]), .B(n3718), .Z(n2267) );
  NAND U3266 ( .A(n2098), .B(n1964), .Z(n1965) );
  XNOR U3267 ( .A(n2267), .B(n1965), .Z(out[1422]) );
  XOR U3268 ( .A(in[804]), .B(n3722), .Z(n2271) );
  NAND U3269 ( .A(n2100), .B(n1966), .Z(n1967) );
  XNOR U3270 ( .A(n2271), .B(n1967), .Z(out[1423]) );
  XOR U3271 ( .A(in[805]), .B(n3726), .Z(n2276) );
  NAND U3272 ( .A(n2102), .B(n1968), .Z(n1969) );
  XNOR U3273 ( .A(n2276), .B(n1969), .Z(out[1424]) );
  XNOR U3274 ( .A(in[806]), .B(n3730), .Z(n2280) );
  NAND U3275 ( .A(n2104), .B(n1970), .Z(n1971) );
  XNOR U3276 ( .A(n2280), .B(n1971), .Z(out[1425]) );
  XNOR U3277 ( .A(in[807]), .B(n3734), .Z(n2284) );
  NAND U3278 ( .A(n2107), .B(n1972), .Z(n1973) );
  XNOR U3279 ( .A(n2284), .B(n1973), .Z(out[1426]) );
  XNOR U3280 ( .A(in[808]), .B(n3738), .Z(n2288) );
  NAND U3281 ( .A(n2109), .B(n1974), .Z(n1975) );
  XNOR U3282 ( .A(n2288), .B(n1975), .Z(out[1427]) );
  XNOR U3283 ( .A(in[809]), .B(n3742), .Z(n2292) );
  NAND U3284 ( .A(n2111), .B(n1976), .Z(n1977) );
  XNOR U3285 ( .A(n2292), .B(n1977), .Z(out[1428]) );
  XNOR U3286 ( .A(in[810]), .B(n3746), .Z(n2296) );
  NAND U3287 ( .A(n2113), .B(n1978), .Z(n1979) );
  XNOR U3288 ( .A(n2296), .B(n1979), .Z(out[1429]) );
  XNOR U3289 ( .A(in[679]), .B(n3926), .Z(n2646) );
  XOR U3290 ( .A(in[613]), .B(n3776), .Z(n4041) );
  XOR U3291 ( .A(in[204]), .B(n3593), .Z(n4039) );
  NAND U3292 ( .A(n4041), .B(n4039), .Z(n1980) );
  XNOR U3293 ( .A(n2646), .B(n1980), .Z(out[142]) );
  XNOR U3294 ( .A(in[811]), .B(n3750), .Z(n2300) );
  NAND U3295 ( .A(n2115), .B(n1981), .Z(n1982) );
  XNOR U3296 ( .A(n2300), .B(n1982), .Z(out[1430]) );
  XNOR U3297 ( .A(in[812]), .B(n3758), .Z(n2304) );
  NAND U3298 ( .A(n2117), .B(n1983), .Z(n1984) );
  XNOR U3299 ( .A(n2304), .B(n1984), .Z(out[1431]) );
  XNOR U3300 ( .A(in[813]), .B(n3762), .Z(n2309) );
  NAND U3301 ( .A(n2119), .B(n1985), .Z(n1986) );
  XNOR U3302 ( .A(n2309), .B(n1986), .Z(out[1432]) );
  XNOR U3303 ( .A(in[814]), .B(n3766), .Z(n2313) );
  NAND U3304 ( .A(n2121), .B(n1987), .Z(n1988) );
  XNOR U3305 ( .A(n2313), .B(n1988), .Z(out[1433]) );
  XNOR U3306 ( .A(in[815]), .B(n3770), .Z(n2317) );
  NAND U3307 ( .A(n2123), .B(n1989), .Z(n1990) );
  XNOR U3308 ( .A(n2317), .B(n1990), .Z(out[1434]) );
  XNOR U3309 ( .A(in[816]), .B(n3774), .Z(n2321) );
  NAND U3310 ( .A(n2125), .B(n1991), .Z(n1992) );
  XNOR U3311 ( .A(n2321), .B(n1992), .Z(out[1435]) );
  XNOR U3312 ( .A(in[817]), .B(n3778), .Z(n2325) );
  NAND U3313 ( .A(n2129), .B(n1993), .Z(n1994) );
  XNOR U3314 ( .A(n2325), .B(n1994), .Z(out[1436]) );
  XNOR U3315 ( .A(in[818]), .B(n3782), .Z(n2329) );
  NAND U3316 ( .A(n2131), .B(n1995), .Z(n1996) );
  XNOR U3317 ( .A(n2329), .B(n1996), .Z(out[1437]) );
  XNOR U3318 ( .A(in[819]), .B(n3786), .Z(n2333) );
  NAND U3319 ( .A(n2133), .B(n1997), .Z(n1998) );
  XNOR U3320 ( .A(n2333), .B(n1998), .Z(out[1438]) );
  XNOR U3321 ( .A(in[820]), .B(n3790), .Z(n2337) );
  NAND U3322 ( .A(n2135), .B(n1999), .Z(n2000) );
  XNOR U3323 ( .A(n2337), .B(n2000), .Z(out[1439]) );
  XNOR U3324 ( .A(in[680]), .B(n3928), .Z(n2649) );
  XOR U3325 ( .A(in[614]), .B(n3780), .Z(n4075) );
  XOR U3326 ( .A(in[205]), .B(n3597), .Z(n4073) );
  NAND U3327 ( .A(n4075), .B(n4073), .Z(n2001) );
  XNOR U3328 ( .A(n2649), .B(n2001), .Z(out[143]) );
  XNOR U3329 ( .A(in[821]), .B(n3794), .Z(n2342) );
  NAND U3330 ( .A(n2137), .B(n2002), .Z(n2003) );
  XNOR U3331 ( .A(n2342), .B(n2003), .Z(out[1440]) );
  XNOR U3332 ( .A(in[822]), .B(n3804), .Z(n2346) );
  NAND U3333 ( .A(n2139), .B(n2004), .Z(n2005) );
  XNOR U3334 ( .A(n2346), .B(n2005), .Z(out[1441]) );
  XNOR U3335 ( .A(in[823]), .B(n3808), .Z(n2351) );
  NAND U3336 ( .A(n2141), .B(n2006), .Z(n2007) );
  XNOR U3337 ( .A(n2351), .B(n2007), .Z(out[1442]) );
  XNOR U3338 ( .A(in[824]), .B(n3812), .Z(n2355) );
  NAND U3339 ( .A(n2143), .B(n2008), .Z(n2009) );
  XNOR U3340 ( .A(n2355), .B(n2009), .Z(out[1443]) );
  XNOR U3341 ( .A(in[825]), .B(n3816), .Z(n2359) );
  NAND U3342 ( .A(n2145), .B(n2010), .Z(n2011) );
  XNOR U3343 ( .A(n2359), .B(n2011), .Z(out[1444]) );
  XNOR U3344 ( .A(in[826]), .B(n3538), .Z(n2363) );
  NAND U3345 ( .A(n2147), .B(n2012), .Z(n2013) );
  XNOR U3346 ( .A(n2363), .B(n2013), .Z(out[1445]) );
  XNOR U3347 ( .A(in[827]), .B(n3542), .Z(n2367) );
  NAND U3348 ( .A(n2150), .B(n2014), .Z(n2015) );
  XNOR U3349 ( .A(n2367), .B(n2015), .Z(out[1446]) );
  XNOR U3350 ( .A(in[828]), .B(n3546), .Z(n2371) );
  NAND U3351 ( .A(n2152), .B(n2016), .Z(n2017) );
  XNOR U3352 ( .A(n2371), .B(n2017), .Z(out[1447]) );
  XNOR U3353 ( .A(in[829]), .B(n3550), .Z(n2375) );
  NAND U3354 ( .A(n2154), .B(n2018), .Z(n2019) );
  XNOR U3355 ( .A(n2375), .B(n2019), .Z(out[1448]) );
  XNOR U3356 ( .A(in[830]), .B(n3554), .Z(n2379) );
  NAND U3357 ( .A(n2156), .B(n2020), .Z(n2021) );
  XNOR U3358 ( .A(n2379), .B(n2021), .Z(out[1449]) );
  XNOR U3359 ( .A(in[681]), .B(n3930), .Z(n2652) );
  XOR U3360 ( .A(in[615]), .B(n3784), .Z(n4113) );
  XOR U3361 ( .A(in[206]), .B(n3601), .Z(n4111) );
  NAND U3362 ( .A(n4113), .B(n4111), .Z(n2022) );
  XNOR U3363 ( .A(n2652), .B(n2022), .Z(out[144]) );
  XNOR U3364 ( .A(in[831]), .B(n3558), .Z(n2383) );
  NAND U3365 ( .A(n2158), .B(n2023), .Z(n2024) );
  XNOR U3366 ( .A(n2383), .B(n2024), .Z(out[1450]) );
  XNOR U3367 ( .A(in[768]), .B(n3562), .Z(n2387) );
  NAND U3368 ( .A(n2160), .B(n2025), .Z(n2026) );
  XNOR U3369 ( .A(n2387), .B(n2026), .Z(out[1451]) );
  XNOR U3370 ( .A(in[769]), .B(n3566), .Z(n2392) );
  NAND U3371 ( .A(n2162), .B(n2027), .Z(n2028) );
  XNOR U3372 ( .A(n2392), .B(n2028), .Z(out[1452]) );
  XOR U3373 ( .A(n3570), .B(in[770]), .Z(n2396) );
  NAND U3374 ( .A(n2164), .B(n2029), .Z(n2030) );
  XNOR U3375 ( .A(n2396), .B(n2030), .Z(out[1453]) );
  XOR U3376 ( .A(n3574), .B(in[771]), .Z(n2400) );
  NAND U3377 ( .A(n2166), .B(n2031), .Z(n2032) );
  XNOR U3378 ( .A(n2400), .B(n2032), .Z(out[1454]) );
  XOR U3379 ( .A(n3582), .B(in[772]), .Z(n2404) );
  NAND U3380 ( .A(n2168), .B(n2033), .Z(n2034) );
  XNOR U3381 ( .A(n2404), .B(n2034), .Z(out[1455]) );
  XOR U3382 ( .A(n3586), .B(in[773]), .Z(n2408) );
  NAND U3383 ( .A(n2171), .B(n2035), .Z(n2036) );
  XNOR U3384 ( .A(n2408), .B(n2036), .Z(out[1456]) );
  XOR U3385 ( .A(n3590), .B(in[774]), .Z(n2412) );
  NAND U3386 ( .A(n2173), .B(n2037), .Z(n2038) );
  XNOR U3387 ( .A(n2412), .B(n2038), .Z(out[1457]) );
  XOR U3388 ( .A(n3594), .B(in[775]), .Z(n2416) );
  NAND U3389 ( .A(n2175), .B(n2039), .Z(n2040) );
  XNOR U3390 ( .A(n2416), .B(n2040), .Z(out[1458]) );
  XOR U3391 ( .A(n3598), .B(in[776]), .Z(n2420) );
  NAND U3392 ( .A(n2177), .B(n2041), .Z(n2042) );
  XNOR U3393 ( .A(n2420), .B(n2042), .Z(out[1459]) );
  XNOR U3394 ( .A(in[682]), .B(n3932), .Z(n2655) );
  XOR U3395 ( .A(in[616]), .B(n3788), .Z(n4147) );
  XOR U3396 ( .A(in[207]), .B(n3605), .Z(n4145) );
  NAND U3397 ( .A(n4147), .B(n4145), .Z(n2043) );
  XNOR U3398 ( .A(n2655), .B(n2043), .Z(out[145]) );
  XOR U3399 ( .A(in[777]), .B(n3602), .Z(n2424) );
  NAND U3400 ( .A(n2179), .B(n2044), .Z(n2045) );
  XNOR U3401 ( .A(n2424), .B(n2045), .Z(out[1460]) );
  XOR U3402 ( .A(n3606), .B(in[778]), .Z(n2428) );
  NAND U3403 ( .A(n2181), .B(n2046), .Z(n2047) );
  XNOR U3404 ( .A(n2428), .B(n2047), .Z(out[1461]) );
  XOR U3405 ( .A(n3610), .B(in[779]), .Z(n2433) );
  NAND U3406 ( .A(n2183), .B(n2048), .Z(n2049) );
  XNOR U3407 ( .A(n2433), .B(n2049), .Z(out[1462]) );
  XOR U3408 ( .A(in[780]), .B(n3614), .Z(n2437) );
  NAND U3409 ( .A(n2185), .B(n2050), .Z(n2051) );
  XNOR U3410 ( .A(n2437), .B(n2051), .Z(out[1463]) );
  XOR U3411 ( .A(in[781]), .B(n3618), .Z(n2441) );
  NAND U3412 ( .A(n2187), .B(n2052), .Z(n2053) );
  XNOR U3413 ( .A(n2441), .B(n2053), .Z(out[1464]) );
  XOR U3414 ( .A(in[782]), .B(n3626), .Z(n2445) );
  NAND U3415 ( .A(n2189), .B(n2054), .Z(n2055) );
  XNOR U3416 ( .A(n2445), .B(n2055), .Z(out[1465]) );
  XOR U3417 ( .A(in[783]), .B(n3630), .Z(n2449) );
  NAND U3418 ( .A(n2192), .B(n2056), .Z(n2057) );
  XNOR U3419 ( .A(n2449), .B(n2057), .Z(out[1466]) );
  XOR U3420 ( .A(in[784]), .B(n3634), .Z(n2453) );
  NAND U3421 ( .A(n2194), .B(n2058), .Z(n2059) );
  XNOR U3422 ( .A(n2453), .B(n2059), .Z(out[1467]) );
  XOR U3423 ( .A(in[785]), .B(n3638), .Z(n2457) );
  NAND U3424 ( .A(n2196), .B(n2060), .Z(n2061) );
  XNOR U3425 ( .A(n2457), .B(n2061), .Z(out[1468]) );
  XOR U3426 ( .A(in[786]), .B(n3642), .Z(n2461) );
  NAND U3427 ( .A(n2198), .B(n2062), .Z(n2063) );
  XNOR U3428 ( .A(n2461), .B(n2063), .Z(out[1469]) );
  XNOR U3429 ( .A(in[683]), .B(n3934), .Z(n2658) );
  XOR U3430 ( .A(in[617]), .B(n3792), .Z(n4181) );
  XOR U3431 ( .A(in[208]), .B(n3609), .Z(n4179) );
  NAND U3432 ( .A(n4181), .B(n4179), .Z(n2064) );
  XNOR U3433 ( .A(n2658), .B(n2064), .Z(out[146]) );
  XOR U3434 ( .A(in[787]), .B(n3646), .Z(n2465) );
  NAND U3435 ( .A(n2200), .B(n2065), .Z(n2066) );
  XNOR U3436 ( .A(n2465), .B(n2066), .Z(out[1470]) );
  XOR U3437 ( .A(in[788]), .B(n3650), .Z(n2469) );
  NAND U3438 ( .A(n2202), .B(n2067), .Z(n2068) );
  XNOR U3439 ( .A(n2469), .B(n2068), .Z(out[1471]) );
  OR U3440 ( .A(n2205), .B(n2069), .Z(n2070) );
  XNOR U3441 ( .A(n2204), .B(n2070), .Z(out[1472]) );
  OR U3442 ( .A(n2210), .B(n2071), .Z(n2072) );
  XNOR U3443 ( .A(n2209), .B(n2072), .Z(out[1473]) );
  OR U3444 ( .A(n2215), .B(n2073), .Z(n2074) );
  XNOR U3445 ( .A(n2214), .B(n2074), .Z(out[1474]) );
  OR U3446 ( .A(n2219), .B(n2075), .Z(n2076) );
  XNOR U3447 ( .A(n2218), .B(n2076), .Z(out[1475]) );
  OR U3448 ( .A(n2225), .B(n2077), .Z(n2078) );
  XNOR U3449 ( .A(n2224), .B(n2078), .Z(out[1476]) );
  OR U3450 ( .A(n2229), .B(n2079), .Z(n2080) );
  XNOR U3451 ( .A(n2228), .B(n2080), .Z(out[1477]) );
  OR U3452 ( .A(n2233), .B(n2081), .Z(n2082) );
  XNOR U3453 ( .A(n2232), .B(n2082), .Z(out[1478]) );
  OR U3454 ( .A(n2237), .B(n2083), .Z(n2084) );
  XNOR U3455 ( .A(n2236), .B(n2084), .Z(out[1479]) );
  XNOR U3456 ( .A(in[684]), .B(n3936), .Z(n2661) );
  XOR U3457 ( .A(in[618]), .B(n3802), .Z(n4207) );
  XOR U3458 ( .A(in[209]), .B(n3613), .Z(n4205) );
  NAND U3459 ( .A(n4207), .B(n4205), .Z(n2085) );
  XNOR U3460 ( .A(n2661), .B(n2085), .Z(out[147]) );
  OR U3461 ( .A(n2242), .B(n2086), .Z(n2087) );
  XNOR U3462 ( .A(n2241), .B(n2087), .Z(out[1480]) );
  OR U3463 ( .A(n2246), .B(n2088), .Z(n2089) );
  XNOR U3464 ( .A(n2245), .B(n2089), .Z(out[1481]) );
  OR U3465 ( .A(n2250), .B(n2090), .Z(n2091) );
  XNOR U3466 ( .A(n2249), .B(n2091), .Z(out[1482]) );
  OR U3467 ( .A(n2254), .B(n2092), .Z(n2093) );
  XNOR U3468 ( .A(n2253), .B(n2093), .Z(out[1483]) );
  OR U3469 ( .A(n2258), .B(n2094), .Z(n2095) );
  XNOR U3470 ( .A(n2257), .B(n2095), .Z(out[1484]) );
  OR U3471 ( .A(n2262), .B(n2096), .Z(n2097) );
  XNOR U3472 ( .A(n2261), .B(n2097), .Z(out[1485]) );
  OR U3473 ( .A(n2267), .B(n2098), .Z(n2099) );
  XNOR U3474 ( .A(n2266), .B(n2099), .Z(out[1486]) );
  OR U3475 ( .A(n2271), .B(n2100), .Z(n2101) );
  XNOR U3476 ( .A(n2270), .B(n2101), .Z(out[1487]) );
  OR U3477 ( .A(n2276), .B(n2102), .Z(n2103) );
  XNOR U3478 ( .A(n2275), .B(n2103), .Z(out[1488]) );
  OR U3479 ( .A(n2280), .B(n2104), .Z(n2105) );
  XNOR U3480 ( .A(n2279), .B(n2105), .Z(out[1489]) );
  XNOR U3481 ( .A(in[685]), .B(n3938), .Z(n2664) );
  XOR U3482 ( .A(in[619]), .B(n3806), .Z(n4231) );
  XOR U3483 ( .A(in[210]), .B(n3617), .Z(n4229) );
  NAND U3484 ( .A(n4231), .B(n4229), .Z(n2106) );
  XNOR U3485 ( .A(n2664), .B(n2106), .Z(out[148]) );
  OR U3486 ( .A(n2284), .B(n2107), .Z(n2108) );
  XNOR U3487 ( .A(n2283), .B(n2108), .Z(out[1490]) );
  OR U3488 ( .A(n2288), .B(n2109), .Z(n2110) );
  XNOR U3489 ( .A(n2287), .B(n2110), .Z(out[1491]) );
  OR U3490 ( .A(n2292), .B(n2111), .Z(n2112) );
  XNOR U3491 ( .A(n2291), .B(n2112), .Z(out[1492]) );
  OR U3492 ( .A(n2296), .B(n2113), .Z(n2114) );
  XNOR U3493 ( .A(n2295), .B(n2114), .Z(out[1493]) );
  OR U3494 ( .A(n2300), .B(n2115), .Z(n2116) );
  XNOR U3495 ( .A(n2299), .B(n2116), .Z(out[1494]) );
  OR U3496 ( .A(n2304), .B(n2117), .Z(n2118) );
  XNOR U3497 ( .A(n2303), .B(n2118), .Z(out[1495]) );
  OR U3498 ( .A(n2309), .B(n2119), .Z(n2120) );
  XNOR U3499 ( .A(n2308), .B(n2120), .Z(out[1496]) );
  OR U3500 ( .A(n2313), .B(n2121), .Z(n2122) );
  XNOR U3501 ( .A(n2312), .B(n2122), .Z(out[1497]) );
  OR U3502 ( .A(n2317), .B(n2123), .Z(n2124) );
  XNOR U3503 ( .A(n2316), .B(n2124), .Z(out[1498]) );
  OR U3504 ( .A(n2321), .B(n2125), .Z(n2126) );
  XNOR U3505 ( .A(n2320), .B(n2126), .Z(out[1499]) );
  XNOR U3506 ( .A(in[686]), .B(n3940), .Z(n2666) );
  XOR U3507 ( .A(in[620]), .B(n3810), .Z(n4255) );
  XNOR U3508 ( .A(in[211]), .B(n3625), .Z(n4253) );
  NAND U3509 ( .A(n4255), .B(n4253), .Z(n2127) );
  XNOR U3510 ( .A(n2666), .B(n2127), .Z(out[149]) );
  XNOR U3511 ( .A(in[1424]), .B(n3634), .Z(n4038) );
  XOR U3512 ( .A(in[1047]), .B(n4132), .Z(n2645) );
  NAND U3513 ( .A(n4038), .B(n2645), .Z(n2128) );
  XNOR U3514 ( .A(n4039), .B(n2128), .Z(out[14]) );
  OR U3515 ( .A(n2325), .B(n2129), .Z(n2130) );
  XNOR U3516 ( .A(n2324), .B(n2130), .Z(out[1500]) );
  OR U3517 ( .A(n2329), .B(n2131), .Z(n2132) );
  XNOR U3518 ( .A(n2328), .B(n2132), .Z(out[1501]) );
  OR U3519 ( .A(n2333), .B(n2133), .Z(n2134) );
  XNOR U3520 ( .A(n2332), .B(n2134), .Z(out[1502]) );
  OR U3521 ( .A(n2337), .B(n2135), .Z(n2136) );
  XNOR U3522 ( .A(n2336), .B(n2136), .Z(out[1503]) );
  OR U3523 ( .A(n2342), .B(n2137), .Z(n2138) );
  XNOR U3524 ( .A(n2341), .B(n2138), .Z(out[1504]) );
  OR U3525 ( .A(n2346), .B(n2139), .Z(n2140) );
  XNOR U3526 ( .A(n2345), .B(n2140), .Z(out[1505]) );
  OR U3527 ( .A(n2351), .B(n2141), .Z(n2142) );
  XNOR U3528 ( .A(n2350), .B(n2142), .Z(out[1506]) );
  OR U3529 ( .A(n2355), .B(n2143), .Z(n2144) );
  XNOR U3530 ( .A(n2354), .B(n2144), .Z(out[1507]) );
  OR U3531 ( .A(n2359), .B(n2145), .Z(n2146) );
  XNOR U3532 ( .A(n2358), .B(n2146), .Z(out[1508]) );
  OR U3533 ( .A(n2363), .B(n2147), .Z(n2148) );
  XNOR U3534 ( .A(n2362), .B(n2148), .Z(out[1509]) );
  XNOR U3535 ( .A(in[687]), .B(n3942), .Z(n2669) );
  XOR U3536 ( .A(in[621]), .B(n3814), .Z(n4279) );
  XNOR U3537 ( .A(in[212]), .B(n3629), .Z(n4277) );
  NAND U3538 ( .A(n4279), .B(n4277), .Z(n2149) );
  XNOR U3539 ( .A(n2669), .B(n2149), .Z(out[150]) );
  OR U3540 ( .A(n2367), .B(n2150), .Z(n2151) );
  XNOR U3541 ( .A(n2366), .B(n2151), .Z(out[1510]) );
  OR U3542 ( .A(n2371), .B(n2152), .Z(n2153) );
  XNOR U3543 ( .A(n2370), .B(n2153), .Z(out[1511]) );
  OR U3544 ( .A(n2375), .B(n2154), .Z(n2155) );
  XNOR U3545 ( .A(n2374), .B(n2155), .Z(out[1512]) );
  OR U3546 ( .A(n2379), .B(n2156), .Z(n2157) );
  XNOR U3547 ( .A(n2378), .B(n2157), .Z(out[1513]) );
  OR U3548 ( .A(n2383), .B(n2158), .Z(n2159) );
  XNOR U3549 ( .A(n2382), .B(n2159), .Z(out[1514]) );
  OR U3550 ( .A(n2387), .B(n2160), .Z(n2161) );
  XNOR U3551 ( .A(n2386), .B(n2161), .Z(out[1515]) );
  OR U3552 ( .A(n2392), .B(n2162), .Z(n2163) );
  XNOR U3553 ( .A(n2391), .B(n2163), .Z(out[1516]) );
  OR U3554 ( .A(n2396), .B(n2164), .Z(n2165) );
  XNOR U3555 ( .A(n2395), .B(n2165), .Z(out[1517]) );
  OR U3556 ( .A(n2400), .B(n2166), .Z(n2167) );
  XNOR U3557 ( .A(n2399), .B(n2167), .Z(out[1518]) );
  OR U3558 ( .A(n2404), .B(n2168), .Z(n2169) );
  XNOR U3559 ( .A(n2403), .B(n2169), .Z(out[1519]) );
  XNOR U3560 ( .A(in[688]), .B(n3948), .Z(n2672) );
  XOR U3561 ( .A(in[622]), .B(n3536), .Z(n4303) );
  XNOR U3562 ( .A(in[213]), .B(n3633), .Z(n4301) );
  NAND U3563 ( .A(n4303), .B(n4301), .Z(n2170) );
  XNOR U3564 ( .A(n2672), .B(n2170), .Z(out[151]) );
  OR U3565 ( .A(n2408), .B(n2171), .Z(n2172) );
  XNOR U3566 ( .A(n2407), .B(n2172), .Z(out[1520]) );
  OR U3567 ( .A(n2412), .B(n2173), .Z(n2174) );
  XNOR U3568 ( .A(n2411), .B(n2174), .Z(out[1521]) );
  OR U3569 ( .A(n2416), .B(n2175), .Z(n2176) );
  XNOR U3570 ( .A(n2415), .B(n2176), .Z(out[1522]) );
  OR U3571 ( .A(n2420), .B(n2177), .Z(n2178) );
  XNOR U3572 ( .A(n2419), .B(n2178), .Z(out[1523]) );
  OR U3573 ( .A(n2424), .B(n2179), .Z(n2180) );
  XNOR U3574 ( .A(n2423), .B(n2180), .Z(out[1524]) );
  OR U3575 ( .A(n2428), .B(n2181), .Z(n2182) );
  XNOR U3576 ( .A(n2427), .B(n2182), .Z(out[1525]) );
  OR U3577 ( .A(n2433), .B(n2183), .Z(n2184) );
  XNOR U3578 ( .A(n2432), .B(n2184), .Z(out[1526]) );
  OR U3579 ( .A(n2437), .B(n2185), .Z(n2186) );
  XNOR U3580 ( .A(n2436), .B(n2186), .Z(out[1527]) );
  OR U3581 ( .A(n2441), .B(n2187), .Z(n2188) );
  XNOR U3582 ( .A(n2440), .B(n2188), .Z(out[1528]) );
  OR U3583 ( .A(n2445), .B(n2189), .Z(n2190) );
  XNOR U3584 ( .A(n2444), .B(n2190), .Z(out[1529]) );
  XNOR U3585 ( .A(in[689]), .B(n3950), .Z(n2676) );
  XOR U3586 ( .A(in[623]), .B(n3540), .Z(n4327) );
  XNOR U3587 ( .A(in[214]), .B(n3637), .Z(n4325) );
  NAND U3588 ( .A(n4327), .B(n4325), .Z(n2191) );
  XNOR U3589 ( .A(n2676), .B(n2191), .Z(out[152]) );
  OR U3590 ( .A(n2449), .B(n2192), .Z(n2193) );
  XNOR U3591 ( .A(n2448), .B(n2193), .Z(out[1530]) );
  OR U3592 ( .A(n2453), .B(n2194), .Z(n2195) );
  XNOR U3593 ( .A(n2452), .B(n2195), .Z(out[1531]) );
  OR U3594 ( .A(n2457), .B(n2196), .Z(n2197) );
  XNOR U3595 ( .A(n2456), .B(n2197), .Z(out[1532]) );
  OR U3596 ( .A(n2461), .B(n2198), .Z(n2199) );
  XNOR U3597 ( .A(n2460), .B(n2199), .Z(out[1533]) );
  OR U3598 ( .A(n2465), .B(n2200), .Z(n2201) );
  XNOR U3599 ( .A(n2464), .B(n2201), .Z(out[1534]) );
  OR U3600 ( .A(n2469), .B(n2202), .Z(n2203) );
  XNOR U3601 ( .A(n2468), .B(n2203), .Z(out[1535]) );
  ANDN U3602 ( .B(n2205), .A(n2204), .Z(n2208) );
  XOR U3603 ( .A(n2206), .B(round_const[0]), .Z(n2207) );
  XNOR U3604 ( .A(n2208), .B(n2207), .Z(out[1536]) );
  ANDN U3605 ( .B(n2210), .A(n2209), .Z(n2213) );
  XOR U3606 ( .A(n2211), .B(round_const[1]), .Z(n2212) );
  XNOR U3607 ( .A(n2213), .B(n2212), .Z(out[1537]) );
  ANDN U3608 ( .B(n2215), .A(n2214), .Z(n2216) );
  XNOR U3609 ( .A(n2217), .B(n2216), .Z(out[1538]) );
  ANDN U3610 ( .B(n2219), .A(n2218), .Z(n2222) );
  XOR U3611 ( .A(n2220), .B(round_const_3), .Z(n2221) );
  XNOR U3612 ( .A(n2222), .B(n2221), .Z(out[1539]) );
  XNOR U3613 ( .A(in[690]), .B(n3952), .Z(n2679) );
  XOR U3614 ( .A(in[624]), .B(n3544), .Z(n4359) );
  XNOR U3615 ( .A(in[215]), .B(n3641), .Z(n4357) );
  NAND U3616 ( .A(n4359), .B(n4357), .Z(n2223) );
  XNOR U3617 ( .A(n2679), .B(n2223), .Z(out[153]) );
  ANDN U3618 ( .B(n2225), .A(n2224), .Z(n2226) );
  XNOR U3619 ( .A(n2227), .B(n2226), .Z(out[1540]) );
  ANDN U3620 ( .B(n2229), .A(n2228), .Z(n2230) );
  XNOR U3621 ( .A(n2231), .B(n2230), .Z(out[1541]) );
  ANDN U3622 ( .B(n2233), .A(n2232), .Z(n2234) );
  XNOR U3623 ( .A(n2235), .B(n2234), .Z(out[1542]) );
  ANDN U3624 ( .B(n2237), .A(n2236), .Z(n2240) );
  XOR U3625 ( .A(n2238), .B(round_const_7), .Z(n2239) );
  XNOR U3626 ( .A(n2240), .B(n2239), .Z(out[1543]) );
  ANDN U3627 ( .B(n2242), .A(n2241), .Z(n2243) );
  XNOR U3628 ( .A(n2244), .B(n2243), .Z(out[1544]) );
  ANDN U3629 ( .B(n2246), .A(n2245), .Z(n2247) );
  XNOR U3630 ( .A(n2248), .B(n2247), .Z(out[1545]) );
  ANDN U3631 ( .B(n2250), .A(n2249), .Z(n2251) );
  XNOR U3632 ( .A(n2252), .B(n2251), .Z(out[1546]) );
  ANDN U3633 ( .B(n2254), .A(n2253), .Z(n2255) );
  XNOR U3634 ( .A(n2256), .B(n2255), .Z(out[1547]) );
  ANDN U3635 ( .B(n2258), .A(n2257), .Z(n2259) );
  XNOR U3636 ( .A(n2260), .B(n2259), .Z(out[1548]) );
  ANDN U3637 ( .B(n2262), .A(n2261), .Z(n2263) );
  XNOR U3638 ( .A(n2264), .B(n2263), .Z(out[1549]) );
  XNOR U3639 ( .A(in[691]), .B(n3954), .Z(n2682) );
  XOR U3640 ( .A(in[625]), .B(n3548), .Z(n4407) );
  XNOR U3641 ( .A(in[216]), .B(n3645), .Z(n4405) );
  NAND U3642 ( .A(n4407), .B(n4405), .Z(n2265) );
  XNOR U3643 ( .A(n2682), .B(n2265), .Z(out[154]) );
  ANDN U3644 ( .B(n2267), .A(n2266), .Z(n2268) );
  XNOR U3645 ( .A(n2269), .B(n2268), .Z(out[1550]) );
  ANDN U3646 ( .B(n2271), .A(n2270), .Z(n2274) );
  XOR U3647 ( .A(n2272), .B(round_const_15), .Z(n2273) );
  XNOR U3648 ( .A(n2274), .B(n2273), .Z(out[1551]) );
  ANDN U3649 ( .B(n2276), .A(n2275), .Z(n2277) );
  XNOR U3650 ( .A(n2278), .B(n2277), .Z(out[1552]) );
  ANDN U3651 ( .B(n2280), .A(n2279), .Z(n2281) );
  XNOR U3652 ( .A(n2282), .B(n2281), .Z(out[1553]) );
  ANDN U3653 ( .B(n2284), .A(n2283), .Z(n2285) );
  XNOR U3654 ( .A(n2286), .B(n2285), .Z(out[1554]) );
  ANDN U3655 ( .B(n2288), .A(n2287), .Z(n2289) );
  XNOR U3656 ( .A(n2290), .B(n2289), .Z(out[1555]) );
  ANDN U3657 ( .B(n2292), .A(n2291), .Z(n2293) );
  XNOR U3658 ( .A(n2294), .B(n2293), .Z(out[1556]) );
  ANDN U3659 ( .B(n2296), .A(n2295), .Z(n2297) );
  XNOR U3660 ( .A(n2298), .B(n2297), .Z(out[1557]) );
  ANDN U3661 ( .B(n2300), .A(n2299), .Z(n2301) );
  XNOR U3662 ( .A(n2302), .B(n2301), .Z(out[1558]) );
  ANDN U3663 ( .B(n2304), .A(n2303), .Z(n2305) );
  XNOR U3664 ( .A(n2306), .B(n2305), .Z(out[1559]) );
  XNOR U3665 ( .A(in[692]), .B(n3956), .Z(n2685) );
  XOR U3666 ( .A(in[626]), .B(n3552), .Z(n4451) );
  XNOR U3667 ( .A(in[217]), .B(n3649), .Z(n4449) );
  NAND U3668 ( .A(n4451), .B(n4449), .Z(n2307) );
  XNOR U3669 ( .A(n2685), .B(n2307), .Z(out[155]) );
  ANDN U3670 ( .B(n2309), .A(n2308), .Z(n2310) );
  XNOR U3671 ( .A(n2311), .B(n2310), .Z(out[1560]) );
  ANDN U3672 ( .B(n2313), .A(n2312), .Z(n2314) );
  XNOR U3673 ( .A(n2315), .B(n2314), .Z(out[1561]) );
  ANDN U3674 ( .B(n2317), .A(n2316), .Z(n2318) );
  XNOR U3675 ( .A(n2319), .B(n2318), .Z(out[1562]) );
  ANDN U3676 ( .B(n2321), .A(n2320), .Z(n2322) );
  XNOR U3677 ( .A(n2323), .B(n2322), .Z(out[1563]) );
  ANDN U3678 ( .B(n2325), .A(n2324), .Z(n2326) );
  XNOR U3679 ( .A(n2327), .B(n2326), .Z(out[1564]) );
  ANDN U3680 ( .B(n2329), .A(n2328), .Z(n2330) );
  XNOR U3681 ( .A(n2331), .B(n2330), .Z(out[1565]) );
  ANDN U3682 ( .B(n2333), .A(n2332), .Z(n2334) );
  XNOR U3683 ( .A(n2335), .B(n2334), .Z(out[1566]) );
  ANDN U3684 ( .B(n2337), .A(n2336), .Z(n2340) );
  XOR U3685 ( .A(n2338), .B(round_const_31), .Z(n2339) );
  XNOR U3686 ( .A(n2340), .B(n2339), .Z(out[1567]) );
  ANDN U3687 ( .B(n2342), .A(n2341), .Z(n2343) );
  XNOR U3688 ( .A(n2344), .B(n2343), .Z(out[1568]) );
  ANDN U3689 ( .B(n2346), .A(n2345), .Z(n2347) );
  XNOR U3690 ( .A(n2348), .B(n2347), .Z(out[1569]) );
  XNOR U3691 ( .A(in[693]), .B(n3958), .Z(n2688) );
  XOR U3692 ( .A(in[627]), .B(n3556), .Z(n4495) );
  XNOR U3693 ( .A(in[218]), .B(n3653), .Z(n4492) );
  NAND U3694 ( .A(n4495), .B(n4492), .Z(n2349) );
  XNOR U3695 ( .A(n2688), .B(n2349), .Z(out[156]) );
  ANDN U3696 ( .B(n2351), .A(n2350), .Z(n2352) );
  XNOR U3697 ( .A(n2353), .B(n2352), .Z(out[1570]) );
  ANDN U3698 ( .B(n2355), .A(n2354), .Z(n2356) );
  XNOR U3699 ( .A(n2357), .B(n2356), .Z(out[1571]) );
  ANDN U3700 ( .B(n2359), .A(n2358), .Z(n2360) );
  XNOR U3701 ( .A(n2361), .B(n2360), .Z(out[1572]) );
  ANDN U3702 ( .B(n2363), .A(n2362), .Z(n2364) );
  XNOR U3703 ( .A(n2365), .B(n2364), .Z(out[1573]) );
  ANDN U3704 ( .B(n2367), .A(n2366), .Z(n2368) );
  XNOR U3705 ( .A(n2369), .B(n2368), .Z(out[1574]) );
  ANDN U3706 ( .B(n2371), .A(n2370), .Z(n2372) );
  XNOR U3707 ( .A(n2373), .B(n2372), .Z(out[1575]) );
  ANDN U3708 ( .B(n2375), .A(n2374), .Z(n2376) );
  XNOR U3709 ( .A(n2377), .B(n2376), .Z(out[1576]) );
  ANDN U3710 ( .B(n2379), .A(n2378), .Z(n2380) );
  XNOR U3711 ( .A(n2381), .B(n2380), .Z(out[1577]) );
  ANDN U3712 ( .B(n2383), .A(n2382), .Z(n2384) );
  XNOR U3713 ( .A(n2385), .B(n2384), .Z(out[1578]) );
  ANDN U3714 ( .B(n2387), .A(n2386), .Z(n2388) );
  XNOR U3715 ( .A(n2389), .B(n2388), .Z(out[1579]) );
  XNOR U3716 ( .A(in[694]), .B(n3960), .Z(n2690) );
  XOR U3717 ( .A(in[628]), .B(n3560), .Z(n4539) );
  XNOR U3718 ( .A(in[219]), .B(n3657), .Z(n4536) );
  NAND U3719 ( .A(n4539), .B(n4536), .Z(n2390) );
  XNOR U3720 ( .A(n2690), .B(n2390), .Z(out[157]) );
  ANDN U3721 ( .B(n2392), .A(n2391), .Z(n2393) );
  XNOR U3722 ( .A(n2394), .B(n2393), .Z(out[1580]) );
  ANDN U3723 ( .B(n2396), .A(n2395), .Z(n2397) );
  XNOR U3724 ( .A(n2398), .B(n2397), .Z(out[1581]) );
  ANDN U3725 ( .B(n2400), .A(n2399), .Z(n2401) );
  XNOR U3726 ( .A(n2402), .B(n2401), .Z(out[1582]) );
  ANDN U3727 ( .B(n2404), .A(n2403), .Z(n2405) );
  XNOR U3728 ( .A(n2406), .B(n2405), .Z(out[1583]) );
  ANDN U3729 ( .B(n2408), .A(n2407), .Z(n2409) );
  XNOR U3730 ( .A(n2410), .B(n2409), .Z(out[1584]) );
  ANDN U3731 ( .B(n2412), .A(n2411), .Z(n2413) );
  XNOR U3732 ( .A(n2414), .B(n2413), .Z(out[1585]) );
  ANDN U3733 ( .B(n2416), .A(n2415), .Z(n2417) );
  XNOR U3734 ( .A(n2418), .B(n2417), .Z(out[1586]) );
  ANDN U3735 ( .B(n2420), .A(n2419), .Z(n2421) );
  XNOR U3736 ( .A(n2422), .B(n2421), .Z(out[1587]) );
  ANDN U3737 ( .B(n2424), .A(n2423), .Z(n2425) );
  XNOR U3738 ( .A(n2426), .B(n2425), .Z(out[1588]) );
  ANDN U3739 ( .B(n2428), .A(n2427), .Z(n2429) );
  XNOR U3740 ( .A(n2430), .B(n2429), .Z(out[1589]) );
  XNOR U3741 ( .A(in[695]), .B(n3962), .Z(n2692) );
  XOR U3742 ( .A(in[629]), .B(n3564), .Z(n4583) );
  XNOR U3743 ( .A(in[220]), .B(n3661), .Z(n4580) );
  NAND U3744 ( .A(n4583), .B(n4580), .Z(n2431) );
  XNOR U3745 ( .A(n2692), .B(n2431), .Z(out[158]) );
  ANDN U3746 ( .B(n2433), .A(n2432), .Z(n2434) );
  XNOR U3747 ( .A(n2435), .B(n2434), .Z(out[1590]) );
  ANDN U3748 ( .B(n2437), .A(n2436), .Z(n2438) );
  XNOR U3749 ( .A(n2439), .B(n2438), .Z(out[1591]) );
  ANDN U3750 ( .B(n2441), .A(n2440), .Z(n2442) );
  XNOR U3751 ( .A(n2443), .B(n2442), .Z(out[1592]) );
  ANDN U3752 ( .B(n2445), .A(n2444), .Z(n2446) );
  XNOR U3753 ( .A(n2447), .B(n2446), .Z(out[1593]) );
  ANDN U3754 ( .B(n2449), .A(n2448), .Z(n2450) );
  XNOR U3755 ( .A(n2451), .B(n2450), .Z(out[1594]) );
  ANDN U3756 ( .B(n2453), .A(n2452), .Z(n2454) );
  XNOR U3757 ( .A(n2455), .B(n2454), .Z(out[1595]) );
  ANDN U3758 ( .B(n2457), .A(n2456), .Z(n2458) );
  XNOR U3759 ( .A(n2459), .B(n2458), .Z(out[1596]) );
  ANDN U3760 ( .B(n2461), .A(n2460), .Z(n2462) );
  XNOR U3761 ( .A(n2463), .B(n2462), .Z(out[1597]) );
  ANDN U3762 ( .B(n2465), .A(n2464), .Z(n2466) );
  XNOR U3763 ( .A(n2467), .B(n2466), .Z(out[1598]) );
  ANDN U3764 ( .B(n2469), .A(n2468), .Z(n2472) );
  XOR U3765 ( .A(n2470), .B(round_const_63), .Z(n2471) );
  XNOR U3766 ( .A(n2472), .B(n2471), .Z(out[1599]) );
  XNOR U3767 ( .A(in[696]), .B(n3818), .Z(n2694) );
  XOR U3768 ( .A(in[630]), .B(n3568), .Z(n4627) );
  XNOR U3769 ( .A(in[221]), .B(n3669), .Z(n4624) );
  NAND U3770 ( .A(n4627), .B(n4624), .Z(n2473) );
  XNOR U3771 ( .A(n2694), .B(n2473), .Z(out[159]) );
  XNOR U3772 ( .A(in[1425]), .B(n3638), .Z(n4072) );
  XOR U3773 ( .A(in[1048]), .B(n4135), .Z(n2648) );
  NAND U3774 ( .A(n4072), .B(n2648), .Z(n2474) );
  XNOR U3775 ( .A(n4073), .B(n2474), .Z(out[15]) );
  XNOR U3776 ( .A(in[697]), .B(n3820), .Z(n2696) );
  XOR U3777 ( .A(in[631]), .B(n3572), .Z(n4671) );
  XNOR U3778 ( .A(in[222]), .B(n3673), .Z(n4668) );
  NAND U3779 ( .A(n4671), .B(n4668), .Z(n2475) );
  XNOR U3780 ( .A(n2696), .B(n2475), .Z(out[160]) );
  XNOR U3781 ( .A(in[698]), .B(n3822), .Z(n2698) );
  XOR U3782 ( .A(in[632]), .B(n3580), .Z(n4715) );
  XNOR U3783 ( .A(in[223]), .B(n3677), .Z(n4712) );
  NAND U3784 ( .A(n4715), .B(n4712), .Z(n2476) );
  XNOR U3785 ( .A(n2698), .B(n2476), .Z(out[161]) );
  XNOR U3786 ( .A(in[699]), .B(n3824), .Z(n2702) );
  XOR U3787 ( .A(in[633]), .B(n3584), .Z(n4759) );
  XNOR U3788 ( .A(in[224]), .B(n3681), .Z(n4756) );
  NAND U3789 ( .A(n4759), .B(n4756), .Z(n2477) );
  XNOR U3790 ( .A(n2702), .B(n2477), .Z(out[162]) );
  XNOR U3791 ( .A(in[700]), .B(n3826), .Z(n2704) );
  XOR U3792 ( .A(in[634]), .B(n3588), .Z(n4803) );
  XNOR U3793 ( .A(in[225]), .B(n3685), .Z(n4800) );
  NAND U3794 ( .A(n4803), .B(n4800), .Z(n2478) );
  XNOR U3795 ( .A(n2704), .B(n2478), .Z(out[163]) );
  XOR U3796 ( .A(in[701]), .B(n3828), .Z(n2706) );
  NOR U3797 ( .A(n2550), .B(n2831), .Z(n2479) );
  XNOR U3798 ( .A(n2706), .B(n2479), .Z(out[164]) );
  XOR U3799 ( .A(in[702]), .B(n3834), .Z(n2708) );
  NOR U3800 ( .A(n2552), .B(n2845), .Z(n2480) );
  XNOR U3801 ( .A(n2708), .B(n2480), .Z(out[165]) );
  XOR U3802 ( .A(in[703]), .B(n3836), .Z(n2710) );
  NOR U3803 ( .A(n2555), .B(n2859), .Z(n2481) );
  XNOR U3804 ( .A(n2710), .B(n2481), .Z(out[166]) );
  XOR U3805 ( .A(in[640]), .B(n3838), .Z(n2712) );
  NOR U3806 ( .A(n2557), .B(n2873), .Z(n2482) );
  XNOR U3807 ( .A(n2712), .B(n2482), .Z(out[167]) );
  XOR U3808 ( .A(in[641]), .B(n3840), .Z(n2714) );
  NOR U3809 ( .A(n2559), .B(n2889), .Z(n2483) );
  XNOR U3810 ( .A(n2714), .B(n2483), .Z(out[168]) );
  XOR U3811 ( .A(in[642]), .B(n3842), .Z(n2716) );
  NOR U3812 ( .A(n2561), .B(n2903), .Z(n2484) );
  XNOR U3813 ( .A(n2716), .B(n2484), .Z(out[169]) );
  XNOR U3814 ( .A(in[1426]), .B(n3642), .Z(n4110) );
  XOR U3815 ( .A(in[1049]), .B(n4138), .Z(n2651) );
  NAND U3816 ( .A(n4110), .B(n2651), .Z(n2485) );
  XNOR U3817 ( .A(n4111), .B(n2485), .Z(out[16]) );
  XOR U3818 ( .A(in[643]), .B(n3844), .Z(n2718) );
  NOR U3819 ( .A(n2563), .B(n2917), .Z(n2486) );
  XNOR U3820 ( .A(n2718), .B(n2486), .Z(out[170]) );
  XOR U3821 ( .A(in[644]), .B(n3846), .Z(n2720) );
  NOR U3822 ( .A(n2565), .B(n2931), .Z(n2487) );
  XNOR U3823 ( .A(n2720), .B(n2487), .Z(out[171]) );
  XOR U3824 ( .A(in[645]), .B(n3848), .Z(n2726) );
  NOR U3825 ( .A(n2567), .B(n2947), .Z(n2488) );
  XNOR U3826 ( .A(n2726), .B(n2488), .Z(out[172]) );
  XOR U3827 ( .A(in[646]), .B(n3850), .Z(n2728) );
  NOR U3828 ( .A(n2569), .B(n2971), .Z(n2489) );
  XNOR U3829 ( .A(n2728), .B(n2489), .Z(out[173]) );
  XOR U3830 ( .A(in[647]), .B(n3852), .Z(n2730) );
  NOR U3831 ( .A(n2571), .B(n2995), .Z(n2490) );
  XNOR U3832 ( .A(n2730), .B(n2490), .Z(out[174]) );
  XOR U3833 ( .A(in[648]), .B(n3856), .Z(n2732) );
  NOR U3834 ( .A(n2573), .B(n3019), .Z(n2491) );
  XNOR U3835 ( .A(n2732), .B(n2491), .Z(out[175]) );
  XOR U3836 ( .A(in[649]), .B(n3858), .Z(n2734) );
  NOR U3837 ( .A(n2576), .B(n3043), .Z(n2492) );
  XNOR U3838 ( .A(n2734), .B(n2492), .Z(out[176]) );
  XOR U3839 ( .A(in[650]), .B(n3860), .Z(n2736) );
  NOR U3840 ( .A(n2578), .B(n3067), .Z(n2493) );
  XNOR U3841 ( .A(n2736), .B(n2493), .Z(out[177]) );
  XOR U3842 ( .A(in[651]), .B(n3862), .Z(n2738) );
  NOR U3843 ( .A(n2580), .B(n3093), .Z(n2494) );
  XNOR U3844 ( .A(n2738), .B(n2494), .Z(out[178]) );
  XOR U3845 ( .A(in[652]), .B(n3864), .Z(n2740) );
  NOR U3846 ( .A(n2582), .B(n3117), .Z(n2495) );
  XNOR U3847 ( .A(n2740), .B(n2495), .Z(out[179]) );
  XNOR U3848 ( .A(in[1427]), .B(n3646), .Z(n4144) );
  XOR U3849 ( .A(in[1050]), .B(n4141), .Z(n2654) );
  NAND U3850 ( .A(n4144), .B(n2654), .Z(n2496) );
  XNOR U3851 ( .A(n4145), .B(n2496), .Z(out[17]) );
  XOR U3852 ( .A(in[653]), .B(n3866), .Z(n2742) );
  NOR U3853 ( .A(n2584), .B(n3141), .Z(n2497) );
  XNOR U3854 ( .A(n2742), .B(n2497), .Z(out[180]) );
  XOR U3855 ( .A(in[654]), .B(n3868), .Z(n2744) );
  NOR U3856 ( .A(n2586), .B(n3165), .Z(n2498) );
  XNOR U3857 ( .A(n2744), .B(n2498), .Z(out[181]) );
  XOR U3858 ( .A(in[655]), .B(n3870), .Z(n2748) );
  NOR U3859 ( .A(n2588), .B(n3189), .Z(n2499) );
  XNOR U3860 ( .A(n2748), .B(n2499), .Z(out[182]) );
  XOR U3861 ( .A(in[656]), .B(n3872), .Z(n2750) );
  NOR U3862 ( .A(n2590), .B(n3213), .Z(n2500) );
  XNOR U3863 ( .A(n2750), .B(n2500), .Z(out[183]) );
  XOR U3864 ( .A(in[657]), .B(n3874), .Z(n2752) );
  NOR U3865 ( .A(n2592), .B(n3237), .Z(n2501) );
  XNOR U3866 ( .A(n2752), .B(n2501), .Z(out[184]) );
  XOR U3867 ( .A(in[658]), .B(n3878), .Z(n2754) );
  NOR U3868 ( .A(n2594), .B(n3269), .Z(n2502) );
  XNOR U3869 ( .A(n2754), .B(n2502), .Z(out[185]) );
  XOR U3870 ( .A(in[659]), .B(n3880), .Z(n2756) );
  NOR U3871 ( .A(n2597), .B(n3313), .Z(n2503) );
  XNOR U3872 ( .A(n2756), .B(n2503), .Z(out[186]) );
  XOR U3873 ( .A(in[660]), .B(n3882), .Z(n2758) );
  NOR U3874 ( .A(n2599), .B(n3357), .Z(n2504) );
  XNOR U3875 ( .A(n2758), .B(n2504), .Z(out[187]) );
  XOR U3876 ( .A(in[661]), .B(n3884), .Z(n2760) );
  NOR U3877 ( .A(n2601), .B(n3403), .Z(n2505) );
  XNOR U3878 ( .A(n2760), .B(n2505), .Z(out[188]) );
  XOR U3879 ( .A(in[662]), .B(n3886), .Z(n2762) );
  NOR U3880 ( .A(n2603), .B(n3447), .Z(n2506) );
  XNOR U3881 ( .A(n2762), .B(n2506), .Z(out[189]) );
  XNOR U3882 ( .A(in[1428]), .B(n3650), .Z(n4178) );
  XOR U3883 ( .A(in[1051]), .B(n4148), .Z(n2657) );
  NAND U3884 ( .A(n4178), .B(n2657), .Z(n2507) );
  XNOR U3885 ( .A(n4179), .B(n2507), .Z(out[18]) );
  XOR U3886 ( .A(in[663]), .B(n3888), .Z(n2764) );
  NOR U3887 ( .A(n2605), .B(n3491), .Z(n2508) );
  XNOR U3888 ( .A(n2764), .B(n2508), .Z(out[190]) );
  XOR U3889 ( .A(in[664]), .B(n3890), .Z(n2766) );
  NOR U3890 ( .A(n2607), .B(n3535), .Z(n2509) );
  XNOR U3891 ( .A(n2766), .B(n2509), .Z(out[191]) );
  OR U3892 ( .A(n2610), .B(n3579), .Z(n2510) );
  XNOR U3893 ( .A(n2609), .B(n2510), .Z(out[192]) );
  XOR U3894 ( .A(in[1034]), .B(n4089), .Z(n2613) );
  NOR U3895 ( .A(n2612), .B(n3623), .Z(n2511) );
  XNOR U3896 ( .A(n2613), .B(n2511), .Z(out[193]) );
  XOR U3897 ( .A(in[1035]), .B(n4092), .Z(n2724) );
  NOR U3898 ( .A(n2615), .B(n3667), .Z(n2512) );
  XNOR U3899 ( .A(n2724), .B(n2512), .Z(out[194]) );
  XNOR U3900 ( .A(n4095), .B(in[1036]), .Z(n2874) );
  NOR U3901 ( .A(n2617), .B(n3711), .Z(n2513) );
  XNOR U3902 ( .A(n2874), .B(n2513), .Z(out[195]) );
  XNOR U3903 ( .A(n4098), .B(in[1037]), .Z(n3068) );
  NOR U3904 ( .A(n2620), .B(n3755), .Z(n2514) );
  XNOR U3905 ( .A(n3068), .B(n2514), .Z(out[196]) );
  XNOR U3906 ( .A(n4101), .B(in[1038]), .Z(n3358) );
  NOR U3907 ( .A(n2622), .B(n3799), .Z(n2515) );
  XNOR U3908 ( .A(n3358), .B(n2515), .Z(out[197]) );
  XNOR U3909 ( .A(n4104), .B(in[1039]), .Z(n3800) );
  NOR U3910 ( .A(n2624), .B(n3833), .Z(n2516) );
  XNOR U3911 ( .A(n3800), .B(n2516), .Z(out[198]) );
  XNOR U3912 ( .A(n4107), .B(in[1040]), .Z(n4076) );
  NOR U3913 ( .A(n2626), .B(n3855), .Z(n2517) );
  XNOR U3914 ( .A(n4076), .B(n2517), .Z(out[199]) );
  XNOR U3915 ( .A(in[1429]), .B(n3654), .Z(n4204) );
  XOR U3916 ( .A(in[1052]), .B(n4151), .Z(n2660) );
  NAND U3917 ( .A(n4204), .B(n2660), .Z(n2518) );
  XNOR U3918 ( .A(n4205), .B(n2518), .Z(out[19]) );
  XNOR U3919 ( .A(n3574), .B(in[1411]), .Z(n3620) );
  NANDN U3920 ( .A(n2613), .B(n3620), .Z(n2519) );
  XNOR U3921 ( .A(n3621), .B(n2519), .Z(out[1]) );
  XNOR U3922 ( .A(n4114), .B(in[1041]), .Z(n4360) );
  NOR U3923 ( .A(n2628), .B(n3877), .Z(n2520) );
  XNOR U3924 ( .A(n4360), .B(n2520), .Z(out[200]) );
  XNOR U3925 ( .A(n4117), .B(in[1042]), .Z(n4804) );
  NOR U3926 ( .A(n2630), .B(n3899), .Z(n2521) );
  XNOR U3927 ( .A(n4804), .B(n2521), .Z(out[201]) );
  OR U3928 ( .A(n2633), .B(n3923), .Z(n2522) );
  XNOR U3929 ( .A(n2632), .B(n2522), .Z(out[202]) );
  OR U3930 ( .A(n2636), .B(n3947), .Z(n2523) );
  XNOR U3931 ( .A(n2635), .B(n2523), .Z(out[203]) );
  OR U3932 ( .A(n2639), .B(n3973), .Z(n2524) );
  XNOR U3933 ( .A(n2638), .B(n2524), .Z(out[204]) );
  OR U3934 ( .A(n2642), .B(n4007), .Z(n2525) );
  XNOR U3935 ( .A(n2641), .B(n2525), .Z(out[205]) );
  OR U3936 ( .A(n2646), .B(n4041), .Z(n2526) );
  XNOR U3937 ( .A(n2645), .B(n2526), .Z(out[206]) );
  OR U3938 ( .A(n2649), .B(n4075), .Z(n2527) );
  XNOR U3939 ( .A(n2648), .B(n2527), .Z(out[207]) );
  OR U3940 ( .A(n2652), .B(n4113), .Z(n2528) );
  XNOR U3941 ( .A(n2651), .B(n2528), .Z(out[208]) );
  OR U3942 ( .A(n2655), .B(n4147), .Z(n2529) );
  XNOR U3943 ( .A(n2654), .B(n2529), .Z(out[209]) );
  XNOR U3944 ( .A(in[1430]), .B(n3658), .Z(n4228) );
  XOR U3945 ( .A(in[1053]), .B(n4154), .Z(n2663) );
  NAND U3946 ( .A(n4228), .B(n2663), .Z(n2530) );
  XNOR U3947 ( .A(n4229), .B(n2530), .Z(out[20]) );
  OR U3948 ( .A(n2658), .B(n4181), .Z(n2531) );
  XNOR U3949 ( .A(n2657), .B(n2531), .Z(out[210]) );
  OR U3950 ( .A(n2661), .B(n4207), .Z(n2532) );
  XNOR U3951 ( .A(n2660), .B(n2532), .Z(out[211]) );
  OR U3952 ( .A(n2664), .B(n4231), .Z(n2533) );
  XNOR U3953 ( .A(n2663), .B(n2533), .Z(out[212]) );
  XNOR U3954 ( .A(in[1054]), .B(n4157), .Z(n2667) );
  NOR U3955 ( .A(n2666), .B(n4255), .Z(n2534) );
  XNOR U3956 ( .A(n2667), .B(n2534), .Z(out[213]) );
  XNOR U3957 ( .A(in[1055]), .B(n4160), .Z(n2670) );
  NOR U3958 ( .A(n2669), .B(n4279), .Z(n2535) );
  XNOR U3959 ( .A(n2670), .B(n2535), .Z(out[214]) );
  XNOR U3960 ( .A(in[1056]), .B(n4163), .Z(n2673) );
  NOR U3961 ( .A(n2672), .B(n4303), .Z(n2536) );
  XNOR U3962 ( .A(n2673), .B(n2536), .Z(out[215]) );
  XNOR U3963 ( .A(in[1057]), .B(n4166), .Z(n2677) );
  NOR U3964 ( .A(n2676), .B(n4327), .Z(n2537) );
  XNOR U3965 ( .A(n2677), .B(n2537), .Z(out[216]) );
  XNOR U3966 ( .A(in[1058]), .B(n4169), .Z(n2680) );
  NOR U3967 ( .A(n2679), .B(n4359), .Z(n2538) );
  XNOR U3968 ( .A(n2680), .B(n2538), .Z(out[217]) );
  XNOR U3969 ( .A(in[1059]), .B(n4172), .Z(n2683) );
  NOR U3970 ( .A(n2682), .B(n4407), .Z(n2539) );
  XNOR U3971 ( .A(n2683), .B(n2539), .Z(out[218]) );
  XOR U3972 ( .A(in[1060]), .B(n4175), .Z(n2686) );
  NOR U3973 ( .A(n2685), .B(n4451), .Z(n2540) );
  XNOR U3974 ( .A(n2686), .B(n2540), .Z(out[219]) );
  XNOR U3975 ( .A(in[1431]), .B(n3662), .Z(n4252) );
  NANDN U3976 ( .A(n2667), .B(n4252), .Z(n2541) );
  XNOR U3977 ( .A(n4253), .B(n2541), .Z(out[21]) );
  XOR U3978 ( .A(in[1061]), .B(n4182), .Z(n2700) );
  NOR U3979 ( .A(n2688), .B(n4495), .Z(n2542) );
  XNOR U3980 ( .A(n2700), .B(n2542), .Z(out[220]) );
  XOR U3981 ( .A(in[1062]), .B(n4185), .Z(n2722) );
  NOR U3982 ( .A(n2690), .B(n4539), .Z(n2543) );
  XNOR U3983 ( .A(n2722), .B(n2543), .Z(out[221]) );
  XOR U3984 ( .A(in[1063]), .B(n3964), .Z(n2746) );
  NOR U3985 ( .A(n2692), .B(n4583), .Z(n2544) );
  XNOR U3986 ( .A(n2746), .B(n2544), .Z(out[222]) );
  XOR U3987 ( .A(in[1064]), .B(n3967), .Z(n2768) );
  NOR U3988 ( .A(n2694), .B(n4627), .Z(n2545) );
  XNOR U3989 ( .A(n2768), .B(n2545), .Z(out[223]) );
  XOR U3990 ( .A(in[1065]), .B(n3974), .Z(n2780) );
  NOR U3991 ( .A(n2696), .B(n4671), .Z(n2546) );
  XNOR U3992 ( .A(n2780), .B(n2546), .Z(out[224]) );
  XOR U3993 ( .A(in[1066]), .B(n3977), .Z(n2792) );
  NOR U3994 ( .A(n2698), .B(n4715), .Z(n2547) );
  XNOR U3995 ( .A(n2792), .B(n2547), .Z(out[225]) );
  XOR U3996 ( .A(in[1067]), .B(n3980), .Z(n2804) );
  NOR U3997 ( .A(n2702), .B(n4759), .Z(n2548) );
  XNOR U3998 ( .A(n2804), .B(n2548), .Z(out[226]) );
  XOR U3999 ( .A(in[1068]), .B(n3983), .Z(n2816) );
  NOR U4000 ( .A(n2704), .B(n4803), .Z(n2549) );
  XNOR U4001 ( .A(n2816), .B(n2549), .Z(out[227]) );
  XNOR U4002 ( .A(in[1069]), .B(n3986), .Z(n2829) );
  NAND U4003 ( .A(n2706), .B(n2550), .Z(n2551) );
  XNOR U4004 ( .A(n2829), .B(n2551), .Z(out[228]) );
  XNOR U4005 ( .A(in[1070]), .B(n3989), .Z(n2843) );
  NAND U4006 ( .A(n2708), .B(n2552), .Z(n2553) );
  XNOR U4007 ( .A(n2843), .B(n2553), .Z(out[229]) );
  XNOR U4008 ( .A(in[1432]), .B(n3670), .Z(n4276) );
  NANDN U4009 ( .A(n2670), .B(n4276), .Z(n2554) );
  XNOR U4010 ( .A(n4277), .B(n2554), .Z(out[22]) );
  XNOR U4011 ( .A(in[1071]), .B(n3992), .Z(n2857) );
  NAND U4012 ( .A(n2710), .B(n2555), .Z(n2556) );
  XNOR U4013 ( .A(n2857), .B(n2556), .Z(out[230]) );
  XNOR U4014 ( .A(in[1072]), .B(n3995), .Z(n2871) );
  NAND U4015 ( .A(n2712), .B(n2557), .Z(n2558) );
  XNOR U4016 ( .A(n2871), .B(n2558), .Z(out[231]) );
  XNOR U4017 ( .A(in[1073]), .B(n3998), .Z(n2887) );
  NAND U4018 ( .A(n2714), .B(n2559), .Z(n2560) );
  XNOR U4019 ( .A(n2887), .B(n2560), .Z(out[232]) );
  XNOR U4020 ( .A(in[1074]), .B(n4001), .Z(n2901) );
  NAND U4021 ( .A(n2716), .B(n2561), .Z(n2562) );
  XNOR U4022 ( .A(n2901), .B(n2562), .Z(out[233]) );
  XNOR U4023 ( .A(in[1075]), .B(n4008), .Z(n2915) );
  NAND U4024 ( .A(n2718), .B(n2563), .Z(n2564) );
  XNOR U4025 ( .A(n2915), .B(n2564), .Z(out[234]) );
  XNOR U4026 ( .A(in[1076]), .B(n4011), .Z(n2929) );
  NAND U4027 ( .A(n2720), .B(n2565), .Z(n2566) );
  XNOR U4028 ( .A(n2929), .B(n2566), .Z(out[235]) );
  XNOR U4029 ( .A(in[1077]), .B(n4014), .Z(n2945) );
  NAND U4030 ( .A(n2726), .B(n2567), .Z(n2568) );
  XNOR U4031 ( .A(n2945), .B(n2568), .Z(out[236]) );
  XNOR U4032 ( .A(in[1078]), .B(n4017), .Z(n2969) );
  NAND U4033 ( .A(n2728), .B(n2569), .Z(n2570) );
  XNOR U4034 ( .A(n2969), .B(n2570), .Z(out[237]) );
  XNOR U4035 ( .A(in[1079]), .B(n4020), .Z(n2993) );
  NAND U4036 ( .A(n2730), .B(n2571), .Z(n2572) );
  XNOR U4037 ( .A(n2993), .B(n2572), .Z(out[238]) );
  XNOR U4038 ( .A(in[1080]), .B(n4023), .Z(n3017) );
  NAND U4039 ( .A(n2732), .B(n2573), .Z(n2574) );
  XNOR U4040 ( .A(n3017), .B(n2574), .Z(out[239]) );
  XNOR U4041 ( .A(in[1433]), .B(n3674), .Z(n4300) );
  NANDN U4042 ( .A(n2673), .B(n4300), .Z(n2575) );
  XNOR U4043 ( .A(n4301), .B(n2575), .Z(out[23]) );
  XNOR U4044 ( .A(in[1081]), .B(n4026), .Z(n3041) );
  NAND U4045 ( .A(n2734), .B(n2576), .Z(n2577) );
  XNOR U4046 ( .A(n3041), .B(n2577), .Z(out[240]) );
  XNOR U4047 ( .A(in[1082]), .B(n4029), .Z(n3065) );
  NAND U4048 ( .A(n2736), .B(n2578), .Z(n2579) );
  XNOR U4049 ( .A(n3065), .B(n2579), .Z(out[241]) );
  XNOR U4050 ( .A(in[1083]), .B(n4032), .Z(n3091) );
  NAND U4051 ( .A(n2738), .B(n2580), .Z(n2581) );
  XNOR U4052 ( .A(n3091), .B(n2581), .Z(out[242]) );
  XNOR U4053 ( .A(in[1084]), .B(n4035), .Z(n3115) );
  NAND U4054 ( .A(n2740), .B(n2582), .Z(n2583) );
  XNOR U4055 ( .A(n3115), .B(n2583), .Z(out[243]) );
  XNOR U4056 ( .A(in[1085]), .B(n4042), .Z(n3139) );
  NAND U4057 ( .A(n2742), .B(n2584), .Z(n2585) );
  XNOR U4058 ( .A(n3139), .B(n2585), .Z(out[244]) );
  XNOR U4059 ( .A(in[1086]), .B(n4045), .Z(n3163) );
  NAND U4060 ( .A(n2744), .B(n2586), .Z(n2587) );
  XNOR U4061 ( .A(n3163), .B(n2587), .Z(out[245]) );
  XNOR U4062 ( .A(in[1087]), .B(n4048), .Z(n3187) );
  NAND U4063 ( .A(n2748), .B(n2588), .Z(n2589) );
  XNOR U4064 ( .A(n3187), .B(n2589), .Z(out[246]) );
  XNOR U4065 ( .A(in[1024]), .B(n4051), .Z(n3211) );
  NAND U4066 ( .A(n2750), .B(n2590), .Z(n2591) );
  XNOR U4067 ( .A(n3211), .B(n2591), .Z(out[247]) );
  XNOR U4068 ( .A(in[1025]), .B(n4054), .Z(n3235) );
  NAND U4069 ( .A(n2752), .B(n2592), .Z(n2593) );
  XNOR U4070 ( .A(n3235), .B(n2593), .Z(out[248]) );
  XNOR U4071 ( .A(in[1026]), .B(n4057), .Z(n3267) );
  NAND U4072 ( .A(n2754), .B(n2594), .Z(n2595) );
  XNOR U4073 ( .A(n3267), .B(n2595), .Z(out[249]) );
  XNOR U4074 ( .A(in[1434]), .B(n3678), .Z(n4324) );
  NANDN U4075 ( .A(n2677), .B(n4324), .Z(n2596) );
  XNOR U4076 ( .A(n4325), .B(n2596), .Z(out[24]) );
  XNOR U4077 ( .A(in[1027]), .B(n4060), .Z(n3311) );
  NAND U4078 ( .A(n2756), .B(n2597), .Z(n2598) );
  XNOR U4079 ( .A(n3311), .B(n2598), .Z(out[250]) );
  XNOR U4080 ( .A(in[1028]), .B(n4063), .Z(n3355) );
  NAND U4081 ( .A(n2758), .B(n2599), .Z(n2600) );
  XNOR U4082 ( .A(n3355), .B(n2600), .Z(out[251]) );
  XNOR U4083 ( .A(in[1029]), .B(n4066), .Z(n3401) );
  NAND U4084 ( .A(n2760), .B(n2601), .Z(n2602) );
  XNOR U4085 ( .A(n3401), .B(n2602), .Z(out[252]) );
  XNOR U4086 ( .A(in[1030]), .B(n4069), .Z(n3445) );
  NAND U4087 ( .A(n2762), .B(n2603), .Z(n2604) );
  XNOR U4088 ( .A(n3445), .B(n2604), .Z(out[253]) );
  XNOR U4089 ( .A(in[1031]), .B(n4080), .Z(n3489) );
  NAND U4090 ( .A(n2764), .B(n2605), .Z(n2606) );
  XNOR U4091 ( .A(n3489), .B(n2606), .Z(out[254]) );
  XNOR U4092 ( .A(in[1032]), .B(n4083), .Z(n3533) );
  NAND U4093 ( .A(n2766), .B(n2607), .Z(n2608) );
  XNOR U4094 ( .A(n3533), .B(n2608), .Z(out[255]) );
  ANDN U4095 ( .B(n2610), .A(n2609), .Z(n2611) );
  XNOR U4096 ( .A(n3576), .B(n2611), .Z(out[256]) );
  AND U4097 ( .A(n2613), .B(n2612), .Z(n2614) );
  XNOR U4098 ( .A(n3620), .B(n2614), .Z(out[257]) );
  XOR U4099 ( .A(n3582), .B(in[1412]), .Z(n3665) );
  NAND U4100 ( .A(n2724), .B(n2615), .Z(n2616) );
  XNOR U4101 ( .A(n3665), .B(n2616), .Z(out[258]) );
  XOR U4102 ( .A(n3586), .B(in[1413]), .Z(n3709) );
  NAND U4103 ( .A(n2874), .B(n2617), .Z(n2618) );
  XNOR U4104 ( .A(n3709), .B(n2618), .Z(out[259]) );
  XNOR U4105 ( .A(in[1435]), .B(n3682), .Z(n4356) );
  NANDN U4106 ( .A(n2680), .B(n4356), .Z(n2619) );
  XNOR U4107 ( .A(n4357), .B(n2619), .Z(out[25]) );
  XOR U4108 ( .A(n3590), .B(in[1414]), .Z(n3753) );
  NAND U4109 ( .A(n3068), .B(n2620), .Z(n2621) );
  XNOR U4110 ( .A(n3753), .B(n2621), .Z(out[260]) );
  XOR U4111 ( .A(n3594), .B(in[1415]), .Z(n3797) );
  NAND U4112 ( .A(n3358), .B(n2622), .Z(n2623) );
  XNOR U4113 ( .A(n3797), .B(n2623), .Z(out[261]) );
  XOR U4114 ( .A(n3598), .B(in[1416]), .Z(n3831) );
  NAND U4115 ( .A(n3800), .B(n2624), .Z(n2625) );
  XNOR U4116 ( .A(n3831), .B(n2625), .Z(out[262]) );
  XOR U4117 ( .A(in[1417]), .B(n3602), .Z(n4077) );
  NAND U4118 ( .A(n4076), .B(n2626), .Z(n2627) );
  XNOR U4119 ( .A(n4077), .B(n2627), .Z(out[263]) );
  XOR U4120 ( .A(n3606), .B(in[1418]), .Z(n4361) );
  NAND U4121 ( .A(n4360), .B(n2628), .Z(n2629) );
  XNOR U4122 ( .A(n4361), .B(n2629), .Z(out[264]) );
  XOR U4123 ( .A(n3610), .B(in[1419]), .Z(n4805) );
  NAND U4124 ( .A(n4804), .B(n2630), .Z(n2631) );
  XNOR U4125 ( .A(n4805), .B(n2631), .Z(out[265]) );
  ANDN U4126 ( .B(n2633), .A(n2632), .Z(n2634) );
  XNOR U4127 ( .A(n3920), .B(n2634), .Z(out[266]) );
  ANDN U4128 ( .B(n2636), .A(n2635), .Z(n2637) );
  XNOR U4129 ( .A(n3944), .B(n2637), .Z(out[267]) );
  ANDN U4130 ( .B(n2639), .A(n2638), .Z(n2640) );
  XNOR U4131 ( .A(n3970), .B(n2640), .Z(out[268]) );
  ANDN U4132 ( .B(n2642), .A(n2641), .Z(n2643) );
  XNOR U4133 ( .A(n4004), .B(n2643), .Z(out[269]) );
  XNOR U4134 ( .A(in[1436]), .B(n3686), .Z(n4404) );
  NANDN U4135 ( .A(n2683), .B(n4404), .Z(n2644) );
  XNOR U4136 ( .A(n4405), .B(n2644), .Z(out[26]) );
  ANDN U4137 ( .B(n2646), .A(n2645), .Z(n2647) );
  XNOR U4138 ( .A(n4038), .B(n2647), .Z(out[270]) );
  ANDN U4139 ( .B(n2649), .A(n2648), .Z(n2650) );
  XNOR U4140 ( .A(n4072), .B(n2650), .Z(out[271]) );
  ANDN U4141 ( .B(n2652), .A(n2651), .Z(n2653) );
  XNOR U4142 ( .A(n4110), .B(n2653), .Z(out[272]) );
  ANDN U4143 ( .B(n2655), .A(n2654), .Z(n2656) );
  XNOR U4144 ( .A(n4144), .B(n2656), .Z(out[273]) );
  ANDN U4145 ( .B(n2658), .A(n2657), .Z(n2659) );
  XNOR U4146 ( .A(n4178), .B(n2659), .Z(out[274]) );
  ANDN U4147 ( .B(n2661), .A(n2660), .Z(n2662) );
  XNOR U4148 ( .A(n4204), .B(n2662), .Z(out[275]) );
  ANDN U4149 ( .B(n2664), .A(n2663), .Z(n2665) );
  XNOR U4150 ( .A(n4228), .B(n2665), .Z(out[276]) );
  AND U4151 ( .A(n2667), .B(n2666), .Z(n2668) );
  XNOR U4152 ( .A(n4252), .B(n2668), .Z(out[277]) );
  AND U4153 ( .A(n2670), .B(n2669), .Z(n2671) );
  XNOR U4154 ( .A(n4276), .B(n2671), .Z(out[278]) );
  AND U4155 ( .A(n2673), .B(n2672), .Z(n2674) );
  XNOR U4156 ( .A(n4300), .B(n2674), .Z(out[279]) );
  XNOR U4157 ( .A(in[1437]), .B(n3690), .Z(n4448) );
  NANDN U4158 ( .A(n2686), .B(n4448), .Z(n2675) );
  XNOR U4159 ( .A(n4449), .B(n2675), .Z(out[27]) );
  AND U4160 ( .A(n2677), .B(n2676), .Z(n2678) );
  XNOR U4161 ( .A(n4324), .B(n2678), .Z(out[280]) );
  AND U4162 ( .A(n2680), .B(n2679), .Z(n2681) );
  XNOR U4163 ( .A(n4356), .B(n2681), .Z(out[281]) );
  AND U4164 ( .A(n2683), .B(n2682), .Z(n2684) );
  XNOR U4165 ( .A(n4404), .B(n2684), .Z(out[282]) );
  AND U4166 ( .A(n2686), .B(n2685), .Z(n2687) );
  XNOR U4167 ( .A(n4448), .B(n2687), .Z(out[283]) );
  XOR U4168 ( .A(in[1438]), .B(n3694), .Z(n4493) );
  NAND U4169 ( .A(n2700), .B(n2688), .Z(n2689) );
  XNOR U4170 ( .A(n4493), .B(n2689), .Z(out[284]) );
  XOR U4171 ( .A(in[1439]), .B(n3698), .Z(n4537) );
  NAND U4172 ( .A(n2722), .B(n2690), .Z(n2691) );
  XNOR U4173 ( .A(n4537), .B(n2691), .Z(out[285]) );
  XOR U4174 ( .A(in[1440]), .B(n3702), .Z(n4581) );
  NAND U4175 ( .A(n2746), .B(n2692), .Z(n2693) );
  XNOR U4176 ( .A(n4581), .B(n2693), .Z(out[286]) );
  XOR U4177 ( .A(in[1441]), .B(n3706), .Z(n4625) );
  NAND U4178 ( .A(n2768), .B(n2694), .Z(n2695) );
  XNOR U4179 ( .A(n4625), .B(n2695), .Z(out[287]) );
  XOR U4180 ( .A(in[1442]), .B(n3714), .Z(n4669) );
  NAND U4181 ( .A(n2780), .B(n2696), .Z(n2697) );
  XNOR U4182 ( .A(n4669), .B(n2697), .Z(out[288]) );
  XOR U4183 ( .A(in[1443]), .B(n3718), .Z(n4713) );
  NAND U4184 ( .A(n2792), .B(n2698), .Z(n2699) );
  XNOR U4185 ( .A(n4713), .B(n2699), .Z(out[289]) );
  OR U4186 ( .A(n4493), .B(n2700), .Z(n2701) );
  XNOR U4187 ( .A(n4492), .B(n2701), .Z(out[28]) );
  XOR U4188 ( .A(in[1444]), .B(n3722), .Z(n4757) );
  NAND U4189 ( .A(n2804), .B(n2702), .Z(n2703) );
  XNOR U4190 ( .A(n4757), .B(n2703), .Z(out[290]) );
  XOR U4191 ( .A(in[1445]), .B(n3726), .Z(n4801) );
  NAND U4192 ( .A(n2816), .B(n2704), .Z(n2705) );
  XNOR U4193 ( .A(n4801), .B(n2705), .Z(out[291]) );
  OR U4194 ( .A(n2829), .B(n2706), .Z(n2707) );
  XNOR U4195 ( .A(n2828), .B(n2707), .Z(out[292]) );
  OR U4196 ( .A(n2843), .B(n2708), .Z(n2709) );
  XNOR U4197 ( .A(n2842), .B(n2709), .Z(out[293]) );
  OR U4198 ( .A(n2857), .B(n2710), .Z(n2711) );
  XNOR U4199 ( .A(n2856), .B(n2711), .Z(out[294]) );
  OR U4200 ( .A(n2871), .B(n2712), .Z(n2713) );
  XNOR U4201 ( .A(n2870), .B(n2713), .Z(out[295]) );
  OR U4202 ( .A(n2887), .B(n2714), .Z(n2715) );
  XNOR U4203 ( .A(n2886), .B(n2715), .Z(out[296]) );
  OR U4204 ( .A(n2901), .B(n2716), .Z(n2717) );
  XNOR U4205 ( .A(n2900), .B(n2717), .Z(out[297]) );
  OR U4206 ( .A(n2915), .B(n2718), .Z(n2719) );
  XNOR U4207 ( .A(n2914), .B(n2719), .Z(out[298]) );
  OR U4208 ( .A(n2929), .B(n2720), .Z(n2721) );
  XNOR U4209 ( .A(n2928), .B(n2721), .Z(out[299]) );
  OR U4210 ( .A(n4537), .B(n2722), .Z(n2723) );
  XNOR U4211 ( .A(n4536), .B(n2723), .Z(out[29]) );
  OR U4212 ( .A(n3665), .B(n2724), .Z(n2725) );
  XNOR U4213 ( .A(n3664), .B(n2725), .Z(out[2]) );
  OR U4214 ( .A(n2945), .B(n2726), .Z(n2727) );
  XNOR U4215 ( .A(n2944), .B(n2727), .Z(out[300]) );
  OR U4216 ( .A(n2969), .B(n2728), .Z(n2729) );
  XNOR U4217 ( .A(n2968), .B(n2729), .Z(out[301]) );
  OR U4218 ( .A(n2993), .B(n2730), .Z(n2731) );
  XNOR U4219 ( .A(n2992), .B(n2731), .Z(out[302]) );
  OR U4220 ( .A(n3017), .B(n2732), .Z(n2733) );
  XNOR U4221 ( .A(n3016), .B(n2733), .Z(out[303]) );
  OR U4222 ( .A(n3041), .B(n2734), .Z(n2735) );
  XNOR U4223 ( .A(n3040), .B(n2735), .Z(out[304]) );
  OR U4224 ( .A(n3065), .B(n2736), .Z(n2737) );
  XNOR U4225 ( .A(n3064), .B(n2737), .Z(out[305]) );
  OR U4226 ( .A(n3091), .B(n2738), .Z(n2739) );
  XNOR U4227 ( .A(n3090), .B(n2739), .Z(out[306]) );
  OR U4228 ( .A(n3115), .B(n2740), .Z(n2741) );
  XNOR U4229 ( .A(n3114), .B(n2741), .Z(out[307]) );
  OR U4230 ( .A(n3139), .B(n2742), .Z(n2743) );
  XNOR U4231 ( .A(n3138), .B(n2743), .Z(out[308]) );
  OR U4232 ( .A(n3163), .B(n2744), .Z(n2745) );
  XNOR U4233 ( .A(n3162), .B(n2745), .Z(out[309]) );
  OR U4234 ( .A(n4581), .B(n2746), .Z(n2747) );
  XNOR U4235 ( .A(n4580), .B(n2747), .Z(out[30]) );
  OR U4236 ( .A(n3187), .B(n2748), .Z(n2749) );
  XNOR U4237 ( .A(n3186), .B(n2749), .Z(out[310]) );
  OR U4238 ( .A(n3211), .B(n2750), .Z(n2751) );
  XNOR U4239 ( .A(n3210), .B(n2751), .Z(out[311]) );
  OR U4240 ( .A(n3235), .B(n2752), .Z(n2753) );
  XNOR U4241 ( .A(n3234), .B(n2753), .Z(out[312]) );
  OR U4242 ( .A(n3267), .B(n2754), .Z(n2755) );
  XNOR U4243 ( .A(n3266), .B(n2755), .Z(out[313]) );
  OR U4244 ( .A(n3311), .B(n2756), .Z(n2757) );
  XNOR U4245 ( .A(n3310), .B(n2757), .Z(out[314]) );
  OR U4246 ( .A(n3355), .B(n2758), .Z(n2759) );
  XNOR U4247 ( .A(n3354), .B(n2759), .Z(out[315]) );
  OR U4248 ( .A(n3401), .B(n2760), .Z(n2761) );
  XNOR U4249 ( .A(n3400), .B(n2761), .Z(out[316]) );
  OR U4250 ( .A(n3445), .B(n2762), .Z(n2763) );
  XNOR U4251 ( .A(n3444), .B(n2763), .Z(out[317]) );
  OR U4252 ( .A(n3489), .B(n2764), .Z(n2765) );
  XNOR U4253 ( .A(n3488), .B(n2765), .Z(out[318]) );
  OR U4254 ( .A(n3533), .B(n2766), .Z(n2767) );
  XNOR U4255 ( .A(n3532), .B(n2767), .Z(out[319]) );
  OR U4256 ( .A(n4625), .B(n2768), .Z(n2769) );
  XNOR U4257 ( .A(n4624), .B(n2769), .Z(out[31]) );
  XNOR U4258 ( .A(in[72]), .B(n4083), .Z(n2940) );
  XOR U4259 ( .A(in[1317]), .B(n3918), .Z(n3253) );
  XOR U4260 ( .A(in[1244]), .B(n3736), .Z(n3250) );
  NAND U4261 ( .A(n3253), .B(n3250), .Z(n2770) );
  XNOR U4262 ( .A(n2940), .B(n2770), .Z(out[320]) );
  XNOR U4263 ( .A(in[73]), .B(n4086), .Z(n2942) );
  XOR U4264 ( .A(in[1318]), .B(n3924), .Z(n3257) );
  XOR U4265 ( .A(in[1245]), .B(n3740), .Z(n3254) );
  NAND U4266 ( .A(n3257), .B(n3254), .Z(n2771) );
  XNOR U4267 ( .A(n2942), .B(n2771), .Z(out[321]) );
  XNOR U4268 ( .A(in[74]), .B(n4089), .Z(n2948) );
  XOR U4269 ( .A(in[1319]), .B(n3926), .Z(n3261) );
  XOR U4270 ( .A(in[1246]), .B(n3744), .Z(n3258) );
  NAND U4271 ( .A(n3261), .B(n3258), .Z(n2772) );
  XNOR U4272 ( .A(n2948), .B(n2772), .Z(out[322]) );
  XNOR U4273 ( .A(in[75]), .B(n4092), .Z(n2950) );
  XOR U4274 ( .A(in[1320]), .B(n3928), .Z(n3265) );
  XOR U4275 ( .A(in[1247]), .B(n3748), .Z(n3262) );
  NAND U4276 ( .A(n3265), .B(n3262), .Z(n2773) );
  XNOR U4277 ( .A(n2950), .B(n2773), .Z(out[323]) );
  XOR U4278 ( .A(n4095), .B(in[76]), .Z(n2952) );
  XOR U4279 ( .A(in[1321]), .B(n3930), .Z(n3273) );
  XOR U4280 ( .A(in[1248]), .B(n3756), .Z(n3270) );
  NAND U4281 ( .A(n3273), .B(n3270), .Z(n2774) );
  XNOR U4282 ( .A(n2952), .B(n2774), .Z(out[324]) );
  XOR U4283 ( .A(n4098), .B(in[77]), .Z(n2954) );
  XOR U4284 ( .A(in[1322]), .B(n3932), .Z(n3277) );
  XOR U4285 ( .A(in[1249]), .B(n3760), .Z(n3274) );
  NAND U4286 ( .A(n3277), .B(n3274), .Z(n2775) );
  XNOR U4287 ( .A(n2954), .B(n2775), .Z(out[325]) );
  XOR U4288 ( .A(n4101), .B(in[78]), .Z(n2956) );
  XOR U4289 ( .A(in[1323]), .B(n3934), .Z(n3281) );
  XOR U4290 ( .A(in[1250]), .B(n3764), .Z(n3278) );
  NAND U4291 ( .A(n3281), .B(n3278), .Z(n2776) );
  XNOR U4292 ( .A(n2956), .B(n2776), .Z(out[326]) );
  XOR U4293 ( .A(n4104), .B(in[79]), .Z(n2958) );
  XOR U4294 ( .A(in[1324]), .B(n3936), .Z(n3285) );
  XOR U4295 ( .A(in[1251]), .B(n3768), .Z(n3282) );
  NAND U4296 ( .A(n3285), .B(n3282), .Z(n2777) );
  XNOR U4297 ( .A(n2958), .B(n2777), .Z(out[327]) );
  XOR U4298 ( .A(n4107), .B(in[80]), .Z(n2960) );
  XOR U4299 ( .A(in[1325]), .B(n3938), .Z(n3289) );
  XOR U4300 ( .A(in[1252]), .B(n3772), .Z(n3286) );
  NAND U4301 ( .A(n3289), .B(n3286), .Z(n2778) );
  XNOR U4302 ( .A(n2960), .B(n2778), .Z(out[328]) );
  XOR U4303 ( .A(n4114), .B(in[81]), .Z(n2962) );
  XOR U4304 ( .A(in[1326]), .B(n3940), .Z(n3293) );
  XNOR U4305 ( .A(in[1253]), .B(n3776), .Z(n3290) );
  NAND U4306 ( .A(n3293), .B(n3290), .Z(n2779) );
  XNOR U4307 ( .A(n2962), .B(n2779), .Z(out[329]) );
  OR U4308 ( .A(n4669), .B(n2780), .Z(n2781) );
  XNOR U4309 ( .A(n4668), .B(n2781), .Z(out[32]) );
  XOR U4310 ( .A(n4117), .B(in[82]), .Z(n2964) );
  XOR U4311 ( .A(in[1327]), .B(n3942), .Z(n3297) );
  XNOR U4312 ( .A(in[1254]), .B(n3780), .Z(n3294) );
  NAND U4313 ( .A(n3297), .B(n3294), .Z(n2782) );
  XNOR U4314 ( .A(n2964), .B(n2782), .Z(out[330]) );
  XOR U4315 ( .A(n4120), .B(in[83]), .Z(n2966) );
  XOR U4316 ( .A(in[1328]), .B(n3948), .Z(n3301) );
  XNOR U4317 ( .A(in[1255]), .B(n3784), .Z(n3298) );
  NAND U4318 ( .A(n3301), .B(n3298), .Z(n2783) );
  XNOR U4319 ( .A(n2966), .B(n2783), .Z(out[331]) );
  XOR U4320 ( .A(in[84]), .B(n4123), .Z(n2972) );
  XOR U4321 ( .A(in[1329]), .B(n3950), .Z(n3305) );
  XNOR U4322 ( .A(in[1256]), .B(n3788), .Z(n3302) );
  NAND U4323 ( .A(n3305), .B(n3302), .Z(n2784) );
  XNOR U4324 ( .A(n2972), .B(n2784), .Z(out[332]) );
  XOR U4325 ( .A(in[85]), .B(n4126), .Z(n2974) );
  XOR U4326 ( .A(in[1330]), .B(n3952), .Z(n3309) );
  XNOR U4327 ( .A(in[1257]), .B(n3792), .Z(n3306) );
  NAND U4328 ( .A(n3309), .B(n3306), .Z(n2785) );
  XNOR U4329 ( .A(n2974), .B(n2785), .Z(out[333]) );
  XOR U4330 ( .A(in[86]), .B(n4129), .Z(n2976) );
  XOR U4331 ( .A(in[1331]), .B(n3954), .Z(n3317) );
  XNOR U4332 ( .A(in[1258]), .B(n3802), .Z(n3314) );
  NAND U4333 ( .A(n3317), .B(n3314), .Z(n2786) );
  XNOR U4334 ( .A(n2976), .B(n2786), .Z(out[334]) );
  XOR U4335 ( .A(in[87]), .B(n4132), .Z(n2978) );
  XOR U4336 ( .A(in[1332]), .B(n3956), .Z(n3321) );
  XNOR U4337 ( .A(in[1259]), .B(n3806), .Z(n3318) );
  NAND U4338 ( .A(n3321), .B(n3318), .Z(n2787) );
  XNOR U4339 ( .A(n2978), .B(n2787), .Z(out[335]) );
  XOR U4340 ( .A(in[88]), .B(n4135), .Z(n2980) );
  XOR U4341 ( .A(in[1333]), .B(n3958), .Z(n3325) );
  XNOR U4342 ( .A(in[1260]), .B(n3810), .Z(n3322) );
  NAND U4343 ( .A(n3325), .B(n3322), .Z(n2788) );
  XNOR U4344 ( .A(n2980), .B(n2788), .Z(out[336]) );
  XOR U4345 ( .A(in[89]), .B(n4138), .Z(n2982) );
  XOR U4346 ( .A(in[1334]), .B(n3960), .Z(n3329) );
  XNOR U4347 ( .A(in[1261]), .B(n3814), .Z(n3326) );
  NAND U4348 ( .A(n3329), .B(n3326), .Z(n2789) );
  XNOR U4349 ( .A(n2982), .B(n2789), .Z(out[337]) );
  XOR U4350 ( .A(in[90]), .B(n4141), .Z(n2984) );
  XOR U4351 ( .A(in[1335]), .B(n3962), .Z(n3333) );
  XNOR U4352 ( .A(in[1262]), .B(n3536), .Z(n3330) );
  NAND U4353 ( .A(n3333), .B(n3330), .Z(n2790) );
  XNOR U4354 ( .A(n2984), .B(n2790), .Z(out[338]) );
  XOR U4355 ( .A(in[91]), .B(n4148), .Z(n2986) );
  XOR U4356 ( .A(in[1336]), .B(n3818), .Z(n3337) );
  XNOR U4357 ( .A(in[1263]), .B(n3540), .Z(n3334) );
  NAND U4358 ( .A(n3337), .B(n3334), .Z(n2791) );
  XNOR U4359 ( .A(n2986), .B(n2791), .Z(out[339]) );
  OR U4360 ( .A(n4713), .B(n2792), .Z(n2793) );
  XNOR U4361 ( .A(n4712), .B(n2793), .Z(out[33]) );
  XOR U4362 ( .A(in[92]), .B(n4151), .Z(n2988) );
  XOR U4363 ( .A(in[1337]), .B(n3820), .Z(n3341) );
  XNOR U4364 ( .A(in[1264]), .B(n3544), .Z(n3338) );
  NAND U4365 ( .A(n3341), .B(n3338), .Z(n2794) );
  XNOR U4366 ( .A(n2988), .B(n2794), .Z(out[340]) );
  XOR U4367 ( .A(in[93]), .B(n4154), .Z(n2990) );
  XOR U4368 ( .A(in[1338]), .B(n3822), .Z(n3345) );
  XNOR U4369 ( .A(in[1265]), .B(n3548), .Z(n3342) );
  NAND U4370 ( .A(n3345), .B(n3342), .Z(n2795) );
  XNOR U4371 ( .A(n2990), .B(n2795), .Z(out[341]) );
  XOR U4372 ( .A(in[94]), .B(n4157), .Z(n2996) );
  XOR U4373 ( .A(in[1339]), .B(n3824), .Z(n3349) );
  XNOR U4374 ( .A(in[1266]), .B(n3552), .Z(n3346) );
  NAND U4375 ( .A(n3349), .B(n3346), .Z(n2796) );
  XNOR U4376 ( .A(n2996), .B(n2796), .Z(out[342]) );
  XOR U4377 ( .A(in[95]), .B(n4160), .Z(n2998) );
  XOR U4378 ( .A(in[1340]), .B(n3826), .Z(n3353) );
  XNOR U4379 ( .A(in[1267]), .B(n3556), .Z(n3350) );
  NAND U4380 ( .A(n3353), .B(n3350), .Z(n2797) );
  XNOR U4381 ( .A(n2998), .B(n2797), .Z(out[343]) );
  XOR U4382 ( .A(in[96]), .B(n4163), .Z(n3000) );
  XOR U4383 ( .A(in[1341]), .B(n3828), .Z(n3363) );
  XNOR U4384 ( .A(in[1268]), .B(n3560), .Z(n3360) );
  NAND U4385 ( .A(n3363), .B(n3360), .Z(n2798) );
  XNOR U4386 ( .A(n3000), .B(n2798), .Z(out[344]) );
  XOR U4387 ( .A(in[97]), .B(n4166), .Z(n3002) );
  XOR U4388 ( .A(in[1342]), .B(n3834), .Z(n3367) );
  XNOR U4389 ( .A(in[1269]), .B(n3564), .Z(n3364) );
  NAND U4390 ( .A(n3367), .B(n3364), .Z(n2799) );
  XNOR U4391 ( .A(n3002), .B(n2799), .Z(out[345]) );
  XOR U4392 ( .A(in[98]), .B(n4169), .Z(n3004) );
  XOR U4393 ( .A(in[1343]), .B(n3836), .Z(n3371) );
  XNOR U4394 ( .A(in[1270]), .B(n3568), .Z(n3368) );
  NAND U4395 ( .A(n3371), .B(n3368), .Z(n2800) );
  XNOR U4396 ( .A(n3004), .B(n2800), .Z(out[346]) );
  XOR U4397 ( .A(in[99]), .B(n4172), .Z(n3006) );
  XOR U4398 ( .A(in[1280]), .B(n3838), .Z(n3375) );
  XNOR U4399 ( .A(in[1271]), .B(n3572), .Z(n3372) );
  NAND U4400 ( .A(n3375), .B(n3372), .Z(n2801) );
  XNOR U4401 ( .A(n3006), .B(n2801), .Z(out[347]) );
  XNOR U4402 ( .A(in[100]), .B(n4175), .Z(n3008) );
  XOR U4403 ( .A(in[1281]), .B(n3840), .Z(n3379) );
  XNOR U4404 ( .A(in[1272]), .B(n3580), .Z(n3376) );
  NAND U4405 ( .A(n3379), .B(n3376), .Z(n2802) );
  XNOR U4406 ( .A(n3008), .B(n2802), .Z(out[348]) );
  XNOR U4407 ( .A(in[101]), .B(n4182), .Z(n3010) );
  XOR U4408 ( .A(in[1282]), .B(n3842), .Z(n3383) );
  XNOR U4409 ( .A(in[1273]), .B(n3584), .Z(n3380) );
  NAND U4410 ( .A(n3383), .B(n3380), .Z(n2803) );
  XNOR U4411 ( .A(n3010), .B(n2803), .Z(out[349]) );
  OR U4412 ( .A(n4757), .B(n2804), .Z(n2805) );
  XNOR U4413 ( .A(n4756), .B(n2805), .Z(out[34]) );
  XNOR U4414 ( .A(in[102]), .B(n4185), .Z(n3012) );
  XOR U4415 ( .A(in[1283]), .B(n3844), .Z(n3387) );
  XNOR U4416 ( .A(in[1274]), .B(n3588), .Z(n3384) );
  NAND U4417 ( .A(n3387), .B(n3384), .Z(n2806) );
  XNOR U4418 ( .A(n3012), .B(n2806), .Z(out[350]) );
  XNOR U4419 ( .A(in[103]), .B(n3964), .Z(n3014) );
  XOR U4420 ( .A(in[1284]), .B(n3846), .Z(n3391) );
  XNOR U4421 ( .A(in[1275]), .B(n3592), .Z(n3388) );
  NAND U4422 ( .A(n3391), .B(n3388), .Z(n2807) );
  XNOR U4423 ( .A(n3014), .B(n2807), .Z(out[351]) );
  XNOR U4424 ( .A(in[104]), .B(n3967), .Z(n3020) );
  XOR U4425 ( .A(in[1285]), .B(n3848), .Z(n3395) );
  XNOR U4426 ( .A(in[1276]), .B(n3596), .Z(n3392) );
  NAND U4427 ( .A(n3395), .B(n3392), .Z(n2808) );
  XNOR U4428 ( .A(n3020), .B(n2808), .Z(out[352]) );
  XNOR U4429 ( .A(in[105]), .B(n3974), .Z(n3022) );
  XOR U4430 ( .A(in[1286]), .B(n3850), .Z(n3399) );
  XNOR U4431 ( .A(in[1277]), .B(n3600), .Z(n3396) );
  NAND U4432 ( .A(n3399), .B(n3396), .Z(n2809) );
  XNOR U4433 ( .A(n3022), .B(n2809), .Z(out[353]) );
  XNOR U4434 ( .A(in[106]), .B(n3977), .Z(n3024) );
  XOR U4435 ( .A(in[1287]), .B(n3852), .Z(n3407) );
  XNOR U4436 ( .A(in[1278]), .B(n3604), .Z(n3404) );
  NAND U4437 ( .A(n3407), .B(n3404), .Z(n2810) );
  XNOR U4438 ( .A(n3024), .B(n2810), .Z(out[354]) );
  XNOR U4439 ( .A(in[107]), .B(n3980), .Z(n3026) );
  XOR U4440 ( .A(in[1288]), .B(n3856), .Z(n3411) );
  XNOR U4441 ( .A(in[1279]), .B(n3608), .Z(n3408) );
  NAND U4442 ( .A(n3411), .B(n3408), .Z(n2811) );
  XNOR U4443 ( .A(n3026), .B(n2811), .Z(out[355]) );
  XNOR U4444 ( .A(in[108]), .B(n3983), .Z(n3028) );
  XOR U4445 ( .A(in[1289]), .B(n3858), .Z(n3415) );
  XNOR U4446 ( .A(in[1216]), .B(n3612), .Z(n3412) );
  NAND U4447 ( .A(n3415), .B(n3412), .Z(n2812) );
  XNOR U4448 ( .A(n3028), .B(n2812), .Z(out[356]) );
  XNOR U4449 ( .A(in[109]), .B(n3986), .Z(n3030) );
  XOR U4450 ( .A(in[1290]), .B(n3860), .Z(n3419) );
  XNOR U4451 ( .A(in[1217]), .B(n3616), .Z(n3416) );
  NAND U4452 ( .A(n3419), .B(n3416), .Z(n2813) );
  XNOR U4453 ( .A(n3030), .B(n2813), .Z(out[357]) );
  XNOR U4454 ( .A(in[110]), .B(n3989), .Z(n3032) );
  XOR U4455 ( .A(in[1291]), .B(n3862), .Z(n3423) );
  XNOR U4456 ( .A(in[1218]), .B(n3624), .Z(n3420) );
  NAND U4457 ( .A(n3423), .B(n3420), .Z(n2814) );
  XNOR U4458 ( .A(n3032), .B(n2814), .Z(out[358]) );
  XNOR U4459 ( .A(in[111]), .B(n3992), .Z(n3034) );
  XOR U4460 ( .A(in[1292]), .B(n3864), .Z(n3427) );
  XNOR U4461 ( .A(in[1219]), .B(n3628), .Z(n3424) );
  NAND U4462 ( .A(n3427), .B(n3424), .Z(n2815) );
  XNOR U4463 ( .A(n3034), .B(n2815), .Z(out[359]) );
  OR U4464 ( .A(n4801), .B(n2816), .Z(n2817) );
  XNOR U4465 ( .A(n4800), .B(n2817), .Z(out[35]) );
  XNOR U4466 ( .A(in[112]), .B(n3995), .Z(n3036) );
  XOR U4467 ( .A(in[1293]), .B(n3866), .Z(n3431) );
  XOR U4468 ( .A(in[1220]), .B(n3632), .Z(n3428) );
  NAND U4469 ( .A(n3431), .B(n3428), .Z(n2818) );
  XNOR U4470 ( .A(n3036), .B(n2818), .Z(out[360]) );
  XNOR U4471 ( .A(in[113]), .B(n3998), .Z(n3038) );
  XOR U4472 ( .A(in[1294]), .B(n3868), .Z(n3435) );
  XOR U4473 ( .A(in[1221]), .B(n3636), .Z(n3432) );
  NAND U4474 ( .A(n3435), .B(n3432), .Z(n2819) );
  XNOR U4475 ( .A(n3038), .B(n2819), .Z(out[361]) );
  XNOR U4476 ( .A(in[114]), .B(n4001), .Z(n3044) );
  XOR U4477 ( .A(in[1295]), .B(n3870), .Z(n3439) );
  XOR U4478 ( .A(in[1222]), .B(n3640), .Z(n3436) );
  NAND U4479 ( .A(n3439), .B(n3436), .Z(n2820) );
  XNOR U4480 ( .A(n3044), .B(n2820), .Z(out[362]) );
  XNOR U4481 ( .A(in[115]), .B(n4008), .Z(n3046) );
  XOR U4482 ( .A(in[1296]), .B(n3872), .Z(n3443) );
  XOR U4483 ( .A(in[1223]), .B(n3644), .Z(n3440) );
  NAND U4484 ( .A(n3443), .B(n3440), .Z(n2821) );
  XNOR U4485 ( .A(n3046), .B(n2821), .Z(out[363]) );
  XNOR U4486 ( .A(in[116]), .B(n4011), .Z(n3048) );
  XOR U4487 ( .A(in[1297]), .B(n3874), .Z(n3451) );
  XOR U4488 ( .A(in[1224]), .B(n3648), .Z(n3448) );
  NAND U4489 ( .A(n3451), .B(n3448), .Z(n2822) );
  XNOR U4490 ( .A(n3048), .B(n2822), .Z(out[364]) );
  XNOR U4491 ( .A(in[117]), .B(n4014), .Z(n3050) );
  XOR U4492 ( .A(in[1298]), .B(n3878), .Z(n3455) );
  XOR U4493 ( .A(in[1225]), .B(n3652), .Z(n3452) );
  NAND U4494 ( .A(n3455), .B(n3452), .Z(n2823) );
  XNOR U4495 ( .A(n3050), .B(n2823), .Z(out[365]) );
  XNOR U4496 ( .A(in[118]), .B(n4017), .Z(n3052) );
  XOR U4497 ( .A(in[1299]), .B(n3880), .Z(n3459) );
  XOR U4498 ( .A(in[1226]), .B(n3656), .Z(n3456) );
  NAND U4499 ( .A(n3459), .B(n3456), .Z(n2824) );
  XNOR U4500 ( .A(n3052), .B(n2824), .Z(out[366]) );
  XNOR U4501 ( .A(in[119]), .B(n4020), .Z(n3054) );
  XOR U4502 ( .A(in[1300]), .B(n3882), .Z(n3463) );
  XOR U4503 ( .A(in[1227]), .B(n3660), .Z(n3460) );
  NAND U4504 ( .A(n3463), .B(n3460), .Z(n2825) );
  XNOR U4505 ( .A(n3054), .B(n2825), .Z(out[367]) );
  XNOR U4506 ( .A(in[120]), .B(n4023), .Z(n3056) );
  XOR U4507 ( .A(in[1301]), .B(n3884), .Z(n3467) );
  XOR U4508 ( .A(in[1228]), .B(n3668), .Z(n3464) );
  NAND U4509 ( .A(n3467), .B(n3464), .Z(n2826) );
  XNOR U4510 ( .A(n3056), .B(n2826), .Z(out[368]) );
  XNOR U4511 ( .A(in[121]), .B(n4026), .Z(n3058) );
  XOR U4512 ( .A(in[1302]), .B(n3886), .Z(n3471) );
  XOR U4513 ( .A(in[1229]), .B(n3672), .Z(n3468) );
  NAND U4514 ( .A(n3471), .B(n3468), .Z(n2827) );
  XNOR U4515 ( .A(n3058), .B(n2827), .Z(out[369]) );
  ANDN U4516 ( .B(n2829), .A(n2828), .Z(n2830) );
  XNOR U4517 ( .A(n2831), .B(n2830), .Z(out[36]) );
  XNOR U4518 ( .A(in[122]), .B(n4029), .Z(n3060) );
  XOR U4519 ( .A(in[1303]), .B(n3888), .Z(n3475) );
  XOR U4520 ( .A(in[1230]), .B(n3676), .Z(n3472) );
  NAND U4521 ( .A(n3475), .B(n3472), .Z(n2832) );
  XNOR U4522 ( .A(n3060), .B(n2832), .Z(out[370]) );
  XNOR U4523 ( .A(in[123]), .B(n4032), .Z(n3062) );
  XOR U4524 ( .A(in[1304]), .B(n3890), .Z(n3479) );
  XOR U4525 ( .A(in[1231]), .B(n3680), .Z(n3476) );
  NAND U4526 ( .A(n3479), .B(n3476), .Z(n2833) );
  XNOR U4527 ( .A(n3062), .B(n2833), .Z(out[371]) );
  XNOR U4528 ( .A(in[124]), .B(n4035), .Z(n3070) );
  XOR U4529 ( .A(in[1305]), .B(n3892), .Z(n3483) );
  XOR U4530 ( .A(in[1232]), .B(n3684), .Z(n3480) );
  NAND U4531 ( .A(n3483), .B(n3480), .Z(n2834) );
  XNOR U4532 ( .A(n3070), .B(n2834), .Z(out[372]) );
  XNOR U4533 ( .A(in[125]), .B(n4042), .Z(n3072) );
  XOR U4534 ( .A(in[1306]), .B(n3894), .Z(n3487) );
  XOR U4535 ( .A(in[1233]), .B(n3688), .Z(n3484) );
  NAND U4536 ( .A(n3487), .B(n3484), .Z(n2835) );
  XNOR U4537 ( .A(n3072), .B(n2835), .Z(out[373]) );
  XNOR U4538 ( .A(in[126]), .B(n4045), .Z(n3074) );
  XOR U4539 ( .A(in[1307]), .B(n3896), .Z(n3495) );
  XOR U4540 ( .A(in[1234]), .B(n3692), .Z(n3492) );
  NAND U4541 ( .A(n3495), .B(n3492), .Z(n2836) );
  XNOR U4542 ( .A(n3074), .B(n2836), .Z(out[374]) );
  XNOR U4543 ( .A(in[127]), .B(n4048), .Z(n3076) );
  XOR U4544 ( .A(in[1308]), .B(n3900), .Z(n3499) );
  XOR U4545 ( .A(in[1235]), .B(n3696), .Z(n3496) );
  NAND U4546 ( .A(n3499), .B(n3496), .Z(n2837) );
  XNOR U4547 ( .A(n3076), .B(n2837), .Z(out[375]) );
  XNOR U4548 ( .A(in[64]), .B(n4051), .Z(n3078) );
  XOR U4549 ( .A(in[1309]), .B(n3902), .Z(n3503) );
  XOR U4550 ( .A(in[1236]), .B(n3700), .Z(n3500) );
  NAND U4551 ( .A(n3503), .B(n3500), .Z(n2838) );
  XNOR U4552 ( .A(n3078), .B(n2838), .Z(out[376]) );
  XNOR U4553 ( .A(in[65]), .B(n4054), .Z(n3080) );
  XOR U4554 ( .A(in[1310]), .B(n3904), .Z(n3507) );
  XOR U4555 ( .A(in[1237]), .B(n3704), .Z(n3504) );
  NAND U4556 ( .A(n3507), .B(n3504), .Z(n2839) );
  XNOR U4557 ( .A(n3080), .B(n2839), .Z(out[377]) );
  XNOR U4558 ( .A(in[66]), .B(n4057), .Z(n3082) );
  XOR U4559 ( .A(in[1311]), .B(n3906), .Z(n3511) );
  XOR U4560 ( .A(in[1238]), .B(n3712), .Z(n3508) );
  NAND U4561 ( .A(n3511), .B(n3508), .Z(n2840) );
  XNOR U4562 ( .A(n3082), .B(n2840), .Z(out[378]) );
  XNOR U4563 ( .A(in[67]), .B(n4060), .Z(n3084) );
  XOR U4564 ( .A(in[1312]), .B(n3908), .Z(n3515) );
  XOR U4565 ( .A(in[1239]), .B(n3716), .Z(n3512) );
  NAND U4566 ( .A(n3515), .B(n3512), .Z(n2841) );
  XNOR U4567 ( .A(n3084), .B(n2841), .Z(out[379]) );
  ANDN U4568 ( .B(n2843), .A(n2842), .Z(n2844) );
  XNOR U4569 ( .A(n2845), .B(n2844), .Z(out[37]) );
  XNOR U4570 ( .A(in[68]), .B(n4063), .Z(n3086) );
  XOR U4571 ( .A(in[1313]), .B(n3910), .Z(n3519) );
  XOR U4572 ( .A(in[1240]), .B(n3720), .Z(n3516) );
  NAND U4573 ( .A(n3519), .B(n3516), .Z(n2846) );
  XNOR U4574 ( .A(n3086), .B(n2846), .Z(out[380]) );
  XNOR U4575 ( .A(in[69]), .B(n4066), .Z(n3088) );
  XOR U4576 ( .A(in[1314]), .B(n3912), .Z(n3523) );
  XOR U4577 ( .A(in[1241]), .B(n3724), .Z(n3520) );
  NAND U4578 ( .A(n3523), .B(n3520), .Z(n2847) );
  XNOR U4579 ( .A(n3088), .B(n2847), .Z(out[381]) );
  XNOR U4580 ( .A(in[70]), .B(n4069), .Z(n3094) );
  XOR U4581 ( .A(in[1315]), .B(n3914), .Z(n3527) );
  XOR U4582 ( .A(in[1242]), .B(n3728), .Z(n3524) );
  NAND U4583 ( .A(n3527), .B(n3524), .Z(n2848) );
  XNOR U4584 ( .A(n3094), .B(n2848), .Z(out[382]) );
  XNOR U4585 ( .A(in[71]), .B(n4080), .Z(n3096) );
  XOR U4586 ( .A(in[1316]), .B(n3916), .Z(n3531) );
  XOR U4587 ( .A(in[1243]), .B(n3732), .Z(n3528) );
  NAND U4588 ( .A(n3531), .B(n3528), .Z(n2849) );
  XNOR U4589 ( .A(n3096), .B(n2849), .Z(out[383]) );
  XOR U4590 ( .A(in[497]), .B(n3778), .Z(n3098) );
  NOR U4591 ( .A(n2940), .B(n3253), .Z(n2850) );
  XNOR U4592 ( .A(n3098), .B(n2850), .Z(out[384]) );
  XOR U4593 ( .A(in[498]), .B(n3782), .Z(n3100) );
  NOR U4594 ( .A(n2942), .B(n3257), .Z(n2851) );
  XNOR U4595 ( .A(n3100), .B(n2851), .Z(out[385]) );
  XOR U4596 ( .A(in[499]), .B(n3786), .Z(n3102) );
  NOR U4597 ( .A(n2948), .B(n3261), .Z(n2852) );
  XNOR U4598 ( .A(n3102), .B(n2852), .Z(out[386]) );
  XOR U4599 ( .A(in[500]), .B(n3790), .Z(n3104) );
  NOR U4600 ( .A(n2950), .B(n3265), .Z(n2853) );
  XNOR U4601 ( .A(n3104), .B(n2853), .Z(out[387]) );
  XOR U4602 ( .A(in[501]), .B(n3794), .Z(n3106) );
  NOR U4603 ( .A(n2952), .B(n3273), .Z(n2854) );
  XNOR U4604 ( .A(n3106), .B(n2854), .Z(out[388]) );
  XOR U4605 ( .A(in[502]), .B(n3804), .Z(n3108) );
  NOR U4606 ( .A(n2954), .B(n3277), .Z(n2855) );
  XNOR U4607 ( .A(n3108), .B(n2855), .Z(out[389]) );
  ANDN U4608 ( .B(n2857), .A(n2856), .Z(n2858) );
  XNOR U4609 ( .A(n2859), .B(n2858), .Z(out[38]) );
  XOR U4610 ( .A(in[503]), .B(n3808), .Z(n3110) );
  NOR U4611 ( .A(n2956), .B(n3281), .Z(n2860) );
  XNOR U4612 ( .A(n3110), .B(n2860), .Z(out[390]) );
  XOR U4613 ( .A(in[504]), .B(n3812), .Z(n3112) );
  NOR U4614 ( .A(n2958), .B(n3285), .Z(n2861) );
  XNOR U4615 ( .A(n3112), .B(n2861), .Z(out[391]) );
  XOR U4616 ( .A(in[505]), .B(n3816), .Z(n3118) );
  NOR U4617 ( .A(n2960), .B(n3289), .Z(n2862) );
  XNOR U4618 ( .A(n3118), .B(n2862), .Z(out[392]) );
  XOR U4619 ( .A(in[506]), .B(n3538), .Z(n3120) );
  NOR U4620 ( .A(n2962), .B(n3293), .Z(n2863) );
  XNOR U4621 ( .A(n3120), .B(n2863), .Z(out[393]) );
  XOR U4622 ( .A(in[507]), .B(n3542), .Z(n3122) );
  NOR U4623 ( .A(n2964), .B(n3297), .Z(n2864) );
  XNOR U4624 ( .A(n3122), .B(n2864), .Z(out[394]) );
  XOR U4625 ( .A(in[508]), .B(n3546), .Z(n3124) );
  NOR U4626 ( .A(n2966), .B(n3301), .Z(n2865) );
  XNOR U4627 ( .A(n3124), .B(n2865), .Z(out[395]) );
  XOR U4628 ( .A(in[509]), .B(n3550), .Z(n3126) );
  NOR U4629 ( .A(n2972), .B(n3305), .Z(n2866) );
  XNOR U4630 ( .A(n3126), .B(n2866), .Z(out[396]) );
  XOR U4631 ( .A(in[510]), .B(n3554), .Z(n3128) );
  NOR U4632 ( .A(n2974), .B(n3309), .Z(n2867) );
  XNOR U4633 ( .A(n3128), .B(n2867), .Z(out[397]) );
  XOR U4634 ( .A(in[511]), .B(n3558), .Z(n3130) );
  NOR U4635 ( .A(n2976), .B(n3317), .Z(n2868) );
  XNOR U4636 ( .A(n3130), .B(n2868), .Z(out[398]) );
  XOR U4637 ( .A(in[448]), .B(n3562), .Z(n3132) );
  NOR U4638 ( .A(n2978), .B(n3321), .Z(n2869) );
  XNOR U4639 ( .A(n3132), .B(n2869), .Z(out[399]) );
  ANDN U4640 ( .B(n2871), .A(n2870), .Z(n2872) );
  XNOR U4641 ( .A(n2873), .B(n2872), .Z(out[39]) );
  OR U4642 ( .A(n3709), .B(n2874), .Z(n2875) );
  XNOR U4643 ( .A(n3708), .B(n2875), .Z(out[3]) );
  XOR U4644 ( .A(in[449]), .B(n3566), .Z(n3134) );
  NOR U4645 ( .A(n2980), .B(n3325), .Z(n2876) );
  XNOR U4646 ( .A(n3134), .B(n2876), .Z(out[400]) );
  XNOR U4647 ( .A(n3570), .B(in[450]), .Z(n3136) );
  NOR U4648 ( .A(n2982), .B(n3329), .Z(n2877) );
  XNOR U4649 ( .A(n3136), .B(n2877), .Z(out[401]) );
  XNOR U4650 ( .A(n3574), .B(in[451]), .Z(n3142) );
  NOR U4651 ( .A(n2984), .B(n3333), .Z(n2878) );
  XNOR U4652 ( .A(n3142), .B(n2878), .Z(out[402]) );
  XNOR U4653 ( .A(n3582), .B(in[452]), .Z(n3144) );
  NOR U4654 ( .A(n2986), .B(n3337), .Z(n2879) );
  XNOR U4655 ( .A(n3144), .B(n2879), .Z(out[403]) );
  XNOR U4656 ( .A(n3586), .B(in[453]), .Z(n3146) );
  NOR U4657 ( .A(n2988), .B(n3341), .Z(n2880) );
  XNOR U4658 ( .A(n3146), .B(n2880), .Z(out[404]) );
  XNOR U4659 ( .A(n3590), .B(in[454]), .Z(n3148) );
  NOR U4660 ( .A(n2990), .B(n3345), .Z(n2881) );
  XNOR U4661 ( .A(n3148), .B(n2881), .Z(out[405]) );
  XNOR U4662 ( .A(n3594), .B(in[455]), .Z(n3150) );
  NOR U4663 ( .A(n2996), .B(n3349), .Z(n2882) );
  XNOR U4664 ( .A(n3150), .B(n2882), .Z(out[406]) );
  XNOR U4665 ( .A(n3598), .B(in[456]), .Z(n3152) );
  NOR U4666 ( .A(n2998), .B(n3353), .Z(n2883) );
  XNOR U4667 ( .A(n3152), .B(n2883), .Z(out[407]) );
  XNOR U4668 ( .A(in[457]), .B(n3602), .Z(n3154) );
  NOR U4669 ( .A(n3000), .B(n3363), .Z(n2884) );
  XNOR U4670 ( .A(n3154), .B(n2884), .Z(out[408]) );
  XNOR U4671 ( .A(n3606), .B(in[458]), .Z(n3156) );
  NOR U4672 ( .A(n3002), .B(n3367), .Z(n2885) );
  XNOR U4673 ( .A(n3156), .B(n2885), .Z(out[409]) );
  ANDN U4674 ( .B(n2887), .A(n2886), .Z(n2888) );
  XNOR U4675 ( .A(n2889), .B(n2888), .Z(out[40]) );
  XNOR U4676 ( .A(n3610), .B(in[459]), .Z(n3158) );
  NOR U4677 ( .A(n3004), .B(n3371), .Z(n2890) );
  XNOR U4678 ( .A(n3158), .B(n2890), .Z(out[410]) );
  XNOR U4679 ( .A(in[460]), .B(n3614), .Z(n3160) );
  NOR U4680 ( .A(n3006), .B(n3375), .Z(n2891) );
  XNOR U4681 ( .A(n3160), .B(n2891), .Z(out[411]) );
  XNOR U4682 ( .A(in[461]), .B(n3618), .Z(n3166) );
  NOR U4683 ( .A(n3008), .B(n3379), .Z(n2892) );
  XNOR U4684 ( .A(n3166), .B(n2892), .Z(out[412]) );
  XNOR U4685 ( .A(in[462]), .B(n3626), .Z(n3168) );
  NOR U4686 ( .A(n3010), .B(n3383), .Z(n2893) );
  XNOR U4687 ( .A(n3168), .B(n2893), .Z(out[413]) );
  XNOR U4688 ( .A(in[463]), .B(n3630), .Z(n3170) );
  NOR U4689 ( .A(n3012), .B(n3387), .Z(n2894) );
  XNOR U4690 ( .A(n3170), .B(n2894), .Z(out[414]) );
  XNOR U4691 ( .A(in[464]), .B(n3634), .Z(n3172) );
  NOR U4692 ( .A(n3014), .B(n3391), .Z(n2895) );
  XNOR U4693 ( .A(n3172), .B(n2895), .Z(out[415]) );
  XNOR U4694 ( .A(in[465]), .B(n3638), .Z(n3174) );
  NOR U4695 ( .A(n3020), .B(n3395), .Z(n2896) );
  XNOR U4696 ( .A(n3174), .B(n2896), .Z(out[416]) );
  XNOR U4697 ( .A(in[466]), .B(n3642), .Z(n3176) );
  NOR U4698 ( .A(n3022), .B(n3399), .Z(n2897) );
  XNOR U4699 ( .A(n3176), .B(n2897), .Z(out[417]) );
  XNOR U4700 ( .A(in[467]), .B(n3646), .Z(n3178) );
  NOR U4701 ( .A(n3024), .B(n3407), .Z(n2898) );
  XNOR U4702 ( .A(n3178), .B(n2898), .Z(out[418]) );
  XNOR U4703 ( .A(in[468]), .B(n3650), .Z(n3180) );
  NOR U4704 ( .A(n3026), .B(n3411), .Z(n2899) );
  XNOR U4705 ( .A(n3180), .B(n2899), .Z(out[419]) );
  ANDN U4706 ( .B(n2901), .A(n2900), .Z(n2902) );
  XNOR U4707 ( .A(n2903), .B(n2902), .Z(out[41]) );
  XNOR U4708 ( .A(in[469]), .B(n3654), .Z(n3182) );
  NOR U4709 ( .A(n3028), .B(n3415), .Z(n2904) );
  XNOR U4710 ( .A(n3182), .B(n2904), .Z(out[420]) );
  XNOR U4711 ( .A(in[470]), .B(n3658), .Z(n3184) );
  NOR U4712 ( .A(n3030), .B(n3419), .Z(n2905) );
  XNOR U4713 ( .A(n3184), .B(n2905), .Z(out[421]) );
  XNOR U4714 ( .A(in[471]), .B(n3662), .Z(n3190) );
  NOR U4715 ( .A(n3032), .B(n3423), .Z(n2906) );
  XNOR U4716 ( .A(n3190), .B(n2906), .Z(out[422]) );
  XNOR U4717 ( .A(in[472]), .B(n3670), .Z(n3192) );
  NOR U4718 ( .A(n3034), .B(n3427), .Z(n2907) );
  XNOR U4719 ( .A(n3192), .B(n2907), .Z(out[423]) );
  XNOR U4720 ( .A(in[473]), .B(n3674), .Z(n3194) );
  NOR U4721 ( .A(n3036), .B(n3431), .Z(n2908) );
  XNOR U4722 ( .A(n3194), .B(n2908), .Z(out[424]) );
  XNOR U4723 ( .A(in[474]), .B(n3678), .Z(n3196) );
  NOR U4724 ( .A(n3038), .B(n3435), .Z(n2909) );
  XNOR U4725 ( .A(n3196), .B(n2909), .Z(out[425]) );
  XNOR U4726 ( .A(in[475]), .B(n3682), .Z(n3198) );
  NOR U4727 ( .A(n3044), .B(n3439), .Z(n2910) );
  XNOR U4728 ( .A(n3198), .B(n2910), .Z(out[426]) );
  XNOR U4729 ( .A(in[476]), .B(n3686), .Z(n3200) );
  NOR U4730 ( .A(n3046), .B(n3443), .Z(n2911) );
  XNOR U4731 ( .A(n3200), .B(n2911), .Z(out[427]) );
  XNOR U4732 ( .A(in[477]), .B(n3690), .Z(n3202) );
  NOR U4733 ( .A(n3048), .B(n3451), .Z(n2912) );
  XNOR U4734 ( .A(n3202), .B(n2912), .Z(out[428]) );
  XNOR U4735 ( .A(in[478]), .B(n3694), .Z(n3204) );
  NOR U4736 ( .A(n3050), .B(n3455), .Z(n2913) );
  XNOR U4737 ( .A(n3204), .B(n2913), .Z(out[429]) );
  ANDN U4738 ( .B(n2915), .A(n2914), .Z(n2916) );
  XNOR U4739 ( .A(n2917), .B(n2916), .Z(out[42]) );
  XNOR U4740 ( .A(in[479]), .B(n3698), .Z(n3206) );
  NOR U4741 ( .A(n3052), .B(n3459), .Z(n2918) );
  XNOR U4742 ( .A(n3206), .B(n2918), .Z(out[430]) );
  XNOR U4743 ( .A(in[480]), .B(n3702), .Z(n3208) );
  NOR U4744 ( .A(n3054), .B(n3463), .Z(n2919) );
  XNOR U4745 ( .A(n3208), .B(n2919), .Z(out[431]) );
  XNOR U4746 ( .A(in[481]), .B(n3706), .Z(n3214) );
  NOR U4747 ( .A(n3056), .B(n3467), .Z(n2920) );
  XNOR U4748 ( .A(n3214), .B(n2920), .Z(out[432]) );
  XNOR U4749 ( .A(in[482]), .B(n3714), .Z(n3216) );
  NOR U4750 ( .A(n3058), .B(n3471), .Z(n2921) );
  XNOR U4751 ( .A(n3216), .B(n2921), .Z(out[433]) );
  XNOR U4752 ( .A(in[483]), .B(n3718), .Z(n3218) );
  NOR U4753 ( .A(n3060), .B(n3475), .Z(n2922) );
  XNOR U4754 ( .A(n3218), .B(n2922), .Z(out[434]) );
  XNOR U4755 ( .A(in[484]), .B(n3722), .Z(n3220) );
  NOR U4756 ( .A(n3062), .B(n3479), .Z(n2923) );
  XNOR U4757 ( .A(n3220), .B(n2923), .Z(out[435]) );
  XNOR U4758 ( .A(in[485]), .B(n3726), .Z(n3222) );
  NOR U4759 ( .A(n3070), .B(n3483), .Z(n2924) );
  XNOR U4760 ( .A(n3222), .B(n2924), .Z(out[436]) );
  XOR U4761 ( .A(in[486]), .B(n3730), .Z(n3224) );
  NOR U4762 ( .A(n3072), .B(n3487), .Z(n2925) );
  XNOR U4763 ( .A(n3224), .B(n2925), .Z(out[437]) );
  XOR U4764 ( .A(in[487]), .B(n3734), .Z(n3226) );
  NOR U4765 ( .A(n3074), .B(n3495), .Z(n2926) );
  XNOR U4766 ( .A(n3226), .B(n2926), .Z(out[438]) );
  XOR U4767 ( .A(in[488]), .B(n3738), .Z(n3228) );
  NOR U4768 ( .A(n3076), .B(n3499), .Z(n2927) );
  XNOR U4769 ( .A(n3228), .B(n2927), .Z(out[439]) );
  ANDN U4770 ( .B(n2929), .A(n2928), .Z(n2930) );
  XNOR U4771 ( .A(n2931), .B(n2930), .Z(out[43]) );
  XOR U4772 ( .A(in[489]), .B(n3742), .Z(n3230) );
  NOR U4773 ( .A(n3078), .B(n3503), .Z(n2932) );
  XNOR U4774 ( .A(n3230), .B(n2932), .Z(out[440]) );
  XOR U4775 ( .A(in[490]), .B(n3746), .Z(n3232) );
  NOR U4776 ( .A(n3080), .B(n3507), .Z(n2933) );
  XNOR U4777 ( .A(n3232), .B(n2933), .Z(out[441]) );
  XOR U4778 ( .A(in[491]), .B(n3750), .Z(n3238) );
  NOR U4779 ( .A(n3082), .B(n3511), .Z(n2934) );
  XNOR U4780 ( .A(n3238), .B(n2934), .Z(out[442]) );
  XOR U4781 ( .A(in[492]), .B(n3758), .Z(n3240) );
  NOR U4782 ( .A(n3084), .B(n3515), .Z(n2935) );
  XNOR U4783 ( .A(n3240), .B(n2935), .Z(out[443]) );
  XOR U4784 ( .A(in[493]), .B(n3762), .Z(n3242) );
  NOR U4785 ( .A(n3086), .B(n3519), .Z(n2936) );
  XNOR U4786 ( .A(n3242), .B(n2936), .Z(out[444]) );
  XOR U4787 ( .A(in[494]), .B(n3766), .Z(n3244) );
  NOR U4788 ( .A(n3088), .B(n3523), .Z(n2937) );
  XNOR U4789 ( .A(n3244), .B(n2937), .Z(out[445]) );
  XOR U4790 ( .A(in[495]), .B(n3770), .Z(n3246) );
  NOR U4791 ( .A(n3094), .B(n3527), .Z(n2938) );
  XNOR U4792 ( .A(n3246), .B(n2938), .Z(out[446]) );
  XOR U4793 ( .A(in[496]), .B(n3774), .Z(n3248) );
  NOR U4794 ( .A(n3096), .B(n3531), .Z(n2939) );
  XNOR U4795 ( .A(n3248), .B(n2939), .Z(out[447]) );
  XNOR U4796 ( .A(in[886]), .B(n3777), .Z(n3251) );
  NAND U4797 ( .A(n3098), .B(n2940), .Z(n2941) );
  XNOR U4798 ( .A(n3251), .B(n2941), .Z(out[448]) );
  XNOR U4799 ( .A(in[887]), .B(n3781), .Z(n3255) );
  NAND U4800 ( .A(n3100), .B(n2942), .Z(n2943) );
  XNOR U4801 ( .A(n3255), .B(n2943), .Z(out[449]) );
  ANDN U4802 ( .B(n2945), .A(n2944), .Z(n2946) );
  XNOR U4803 ( .A(n2947), .B(n2946), .Z(out[44]) );
  XNOR U4804 ( .A(in[888]), .B(n3785), .Z(n3259) );
  NAND U4805 ( .A(n3102), .B(n2948), .Z(n2949) );
  XNOR U4806 ( .A(n3259), .B(n2949), .Z(out[450]) );
  XNOR U4807 ( .A(in[889]), .B(n3789), .Z(n3263) );
  NAND U4808 ( .A(n3104), .B(n2950), .Z(n2951) );
  XNOR U4809 ( .A(n3263), .B(n2951), .Z(out[451]) );
  XNOR U4810 ( .A(in[890]), .B(n3793), .Z(n3271) );
  NAND U4811 ( .A(n3106), .B(n2952), .Z(n2953) );
  XNOR U4812 ( .A(n3271), .B(n2953), .Z(out[452]) );
  XOR U4813 ( .A(in[891]), .B(n3803), .Z(n3275) );
  NAND U4814 ( .A(n3108), .B(n2954), .Z(n2955) );
  XNOR U4815 ( .A(n3275), .B(n2955), .Z(out[453]) );
  XOR U4816 ( .A(in[892]), .B(n3807), .Z(n3279) );
  NAND U4817 ( .A(n3110), .B(n2956), .Z(n2957) );
  XNOR U4818 ( .A(n3279), .B(n2957), .Z(out[454]) );
  XOR U4819 ( .A(in[893]), .B(n3811), .Z(n3283) );
  NAND U4820 ( .A(n3112), .B(n2958), .Z(n2959) );
  XNOR U4821 ( .A(n3283), .B(n2959), .Z(out[455]) );
  XNOR U4822 ( .A(in[894]), .B(n3815), .Z(n3287) );
  NAND U4823 ( .A(n3118), .B(n2960), .Z(n2961) );
  XNOR U4824 ( .A(n3287), .B(n2961), .Z(out[456]) );
  XOR U4825 ( .A(in[895]), .B(n3537), .Z(n3291) );
  NAND U4826 ( .A(n3120), .B(n2962), .Z(n2963) );
  XNOR U4827 ( .A(n3291), .B(n2963), .Z(out[457]) );
  XOR U4828 ( .A(in[832]), .B(n3541), .Z(n3295) );
  NAND U4829 ( .A(n3122), .B(n2964), .Z(n2965) );
  XNOR U4830 ( .A(n3295), .B(n2965), .Z(out[458]) );
  XOR U4831 ( .A(in[833]), .B(n3545), .Z(n3299) );
  NAND U4832 ( .A(n3124), .B(n2966), .Z(n2967) );
  XNOR U4833 ( .A(n3299), .B(n2967), .Z(out[459]) );
  ANDN U4834 ( .B(n2969), .A(n2968), .Z(n2970) );
  XNOR U4835 ( .A(n2971), .B(n2970), .Z(out[45]) );
  XOR U4836 ( .A(in[834]), .B(n3549), .Z(n3303) );
  NAND U4837 ( .A(n3126), .B(n2972), .Z(n2973) );
  XNOR U4838 ( .A(n3303), .B(n2973), .Z(out[460]) );
  XOR U4839 ( .A(in[835]), .B(n3553), .Z(n3307) );
  NAND U4840 ( .A(n3128), .B(n2974), .Z(n2975) );
  XNOR U4841 ( .A(n3307), .B(n2975), .Z(out[461]) );
  XOR U4842 ( .A(in[836]), .B(n3557), .Z(n3315) );
  NAND U4843 ( .A(n3130), .B(n2976), .Z(n2977) );
  XNOR U4844 ( .A(n3315), .B(n2977), .Z(out[462]) );
  XOR U4845 ( .A(in[837]), .B(n3561), .Z(n3319) );
  NAND U4846 ( .A(n3132), .B(n2978), .Z(n2979) );
  XNOR U4847 ( .A(n3319), .B(n2979), .Z(out[463]) );
  XOR U4848 ( .A(in[838]), .B(n3565), .Z(n3323) );
  NAND U4849 ( .A(n3134), .B(n2980), .Z(n2981) );
  XNOR U4850 ( .A(n3323), .B(n2981), .Z(out[464]) );
  XOR U4851 ( .A(in[839]), .B(n3569), .Z(n3327) );
  NAND U4852 ( .A(n3136), .B(n2982), .Z(n2983) );
  XNOR U4853 ( .A(n3327), .B(n2983), .Z(out[465]) );
  XOR U4854 ( .A(in[840]), .B(n3573), .Z(n3331) );
  NAND U4855 ( .A(n3142), .B(n2984), .Z(n2985) );
  XNOR U4856 ( .A(n3331), .B(n2985), .Z(out[466]) );
  XOR U4857 ( .A(in[841]), .B(n3581), .Z(n3335) );
  NAND U4858 ( .A(n3144), .B(n2986), .Z(n2987) );
  XNOR U4859 ( .A(n3335), .B(n2987), .Z(out[467]) );
  XOR U4860 ( .A(in[842]), .B(n3585), .Z(n3339) );
  NAND U4861 ( .A(n3146), .B(n2988), .Z(n2989) );
  XNOR U4862 ( .A(n3339), .B(n2989), .Z(out[468]) );
  XOR U4863 ( .A(in[843]), .B(n3589), .Z(n3343) );
  NAND U4864 ( .A(n3148), .B(n2990), .Z(n2991) );
  XNOR U4865 ( .A(n3343), .B(n2991), .Z(out[469]) );
  ANDN U4866 ( .B(n2993), .A(n2992), .Z(n2994) );
  XNOR U4867 ( .A(n2995), .B(n2994), .Z(out[46]) );
  XOR U4868 ( .A(in[844]), .B(n3593), .Z(n3347) );
  NAND U4869 ( .A(n3150), .B(n2996), .Z(n2997) );
  XNOR U4870 ( .A(n3347), .B(n2997), .Z(out[470]) );
  XOR U4871 ( .A(in[845]), .B(n3597), .Z(n3351) );
  NAND U4872 ( .A(n3152), .B(n2998), .Z(n2999) );
  XNOR U4873 ( .A(n3351), .B(n2999), .Z(out[471]) );
  XOR U4874 ( .A(in[846]), .B(n3601), .Z(n3361) );
  NAND U4875 ( .A(n3154), .B(n3000), .Z(n3001) );
  XNOR U4876 ( .A(n3361), .B(n3001), .Z(out[472]) );
  XOR U4877 ( .A(in[847]), .B(n3605), .Z(n3365) );
  NAND U4878 ( .A(n3156), .B(n3002), .Z(n3003) );
  XNOR U4879 ( .A(n3365), .B(n3003), .Z(out[473]) );
  XOR U4880 ( .A(in[848]), .B(n3609), .Z(n3369) );
  NAND U4881 ( .A(n3158), .B(n3004), .Z(n3005) );
  XNOR U4882 ( .A(n3369), .B(n3005), .Z(out[474]) );
  XOR U4883 ( .A(in[849]), .B(n3613), .Z(n3373) );
  NAND U4884 ( .A(n3160), .B(n3006), .Z(n3007) );
  XNOR U4885 ( .A(n3373), .B(n3007), .Z(out[475]) );
  XOR U4886 ( .A(in[850]), .B(n3617), .Z(n3377) );
  NAND U4887 ( .A(n3166), .B(n3008), .Z(n3009) );
  XNOR U4888 ( .A(n3377), .B(n3009), .Z(out[476]) );
  XNOR U4889 ( .A(in[851]), .B(n3625), .Z(n3381) );
  NAND U4890 ( .A(n3168), .B(n3010), .Z(n3011) );
  XNOR U4891 ( .A(n3381), .B(n3011), .Z(out[477]) );
  XNOR U4892 ( .A(in[852]), .B(n3629), .Z(n3385) );
  NAND U4893 ( .A(n3170), .B(n3012), .Z(n3013) );
  XNOR U4894 ( .A(n3385), .B(n3013), .Z(out[478]) );
  XNOR U4895 ( .A(in[853]), .B(n3633), .Z(n3389) );
  NAND U4896 ( .A(n3172), .B(n3014), .Z(n3015) );
  XNOR U4897 ( .A(n3389), .B(n3015), .Z(out[479]) );
  ANDN U4898 ( .B(n3017), .A(n3016), .Z(n3018) );
  XNOR U4899 ( .A(n3019), .B(n3018), .Z(out[47]) );
  XNOR U4900 ( .A(in[854]), .B(n3637), .Z(n3393) );
  NAND U4901 ( .A(n3174), .B(n3020), .Z(n3021) );
  XNOR U4902 ( .A(n3393), .B(n3021), .Z(out[480]) );
  XNOR U4903 ( .A(in[855]), .B(n3641), .Z(n3397) );
  NAND U4904 ( .A(n3176), .B(n3022), .Z(n3023) );
  XNOR U4905 ( .A(n3397), .B(n3023), .Z(out[481]) );
  XNOR U4906 ( .A(in[856]), .B(n3645), .Z(n3405) );
  NAND U4907 ( .A(n3178), .B(n3024), .Z(n3025) );
  XNOR U4908 ( .A(n3405), .B(n3025), .Z(out[482]) );
  XNOR U4909 ( .A(in[857]), .B(n3649), .Z(n3409) );
  NAND U4910 ( .A(n3180), .B(n3026), .Z(n3027) );
  XNOR U4911 ( .A(n3409), .B(n3027), .Z(out[483]) );
  XNOR U4912 ( .A(in[858]), .B(n3653), .Z(n3413) );
  NAND U4913 ( .A(n3182), .B(n3028), .Z(n3029) );
  XNOR U4914 ( .A(n3413), .B(n3029), .Z(out[484]) );
  XNOR U4915 ( .A(in[859]), .B(n3657), .Z(n3417) );
  NAND U4916 ( .A(n3184), .B(n3030), .Z(n3031) );
  XNOR U4917 ( .A(n3417), .B(n3031), .Z(out[485]) );
  XNOR U4918 ( .A(in[860]), .B(n3661), .Z(n3421) );
  NAND U4919 ( .A(n3190), .B(n3032), .Z(n3033) );
  XNOR U4920 ( .A(n3421), .B(n3033), .Z(out[486]) );
  XNOR U4921 ( .A(in[861]), .B(n3669), .Z(n3425) );
  NAND U4922 ( .A(n3192), .B(n3034), .Z(n3035) );
  XNOR U4923 ( .A(n3425), .B(n3035), .Z(out[487]) );
  XNOR U4924 ( .A(in[862]), .B(n3673), .Z(n3429) );
  NAND U4925 ( .A(n3194), .B(n3036), .Z(n3037) );
  XNOR U4926 ( .A(n3429), .B(n3037), .Z(out[488]) );
  XNOR U4927 ( .A(in[863]), .B(n3677), .Z(n3433) );
  NAND U4928 ( .A(n3196), .B(n3038), .Z(n3039) );
  XNOR U4929 ( .A(n3433), .B(n3039), .Z(out[489]) );
  ANDN U4930 ( .B(n3041), .A(n3040), .Z(n3042) );
  XNOR U4931 ( .A(n3043), .B(n3042), .Z(out[48]) );
  XNOR U4932 ( .A(in[864]), .B(n3681), .Z(n3437) );
  NAND U4933 ( .A(n3198), .B(n3044), .Z(n3045) );
  XNOR U4934 ( .A(n3437), .B(n3045), .Z(out[490]) );
  XNOR U4935 ( .A(in[865]), .B(n3685), .Z(n3441) );
  NAND U4936 ( .A(n3200), .B(n3046), .Z(n3047) );
  XNOR U4937 ( .A(n3441), .B(n3047), .Z(out[491]) );
  XOR U4938 ( .A(n3689), .B(in[866]), .Z(n3449) );
  NAND U4939 ( .A(n3202), .B(n3048), .Z(n3049) );
  XNOR U4940 ( .A(n3449), .B(n3049), .Z(out[492]) );
  XOR U4941 ( .A(n3693), .B(in[867]), .Z(n3453) );
  NAND U4942 ( .A(n3204), .B(n3050), .Z(n3051) );
  XNOR U4943 ( .A(n3453), .B(n3051), .Z(out[493]) );
  XOR U4944 ( .A(n3697), .B(in[868]), .Z(n3457) );
  NAND U4945 ( .A(n3206), .B(n3052), .Z(n3053) );
  XNOR U4946 ( .A(n3457), .B(n3053), .Z(out[494]) );
  XOR U4947 ( .A(n3701), .B(in[869]), .Z(n3461) );
  NAND U4948 ( .A(n3208), .B(n3054), .Z(n3055) );
  XNOR U4949 ( .A(n3461), .B(n3055), .Z(out[495]) );
  XNOR U4950 ( .A(in[870]), .B(n3705), .Z(n3465) );
  NAND U4951 ( .A(n3214), .B(n3056), .Z(n3057) );
  XNOR U4952 ( .A(n3465), .B(n3057), .Z(out[496]) );
  XNOR U4953 ( .A(in[871]), .B(n3713), .Z(n3469) );
  NAND U4954 ( .A(n3216), .B(n3058), .Z(n3059) );
  XNOR U4955 ( .A(n3469), .B(n3059), .Z(out[497]) );
  XNOR U4956 ( .A(in[872]), .B(n3717), .Z(n3473) );
  NAND U4957 ( .A(n3218), .B(n3060), .Z(n3061) );
  XNOR U4958 ( .A(n3473), .B(n3061), .Z(out[498]) );
  XNOR U4959 ( .A(in[873]), .B(n3721), .Z(n3477) );
  NAND U4960 ( .A(n3220), .B(n3062), .Z(n3063) );
  XNOR U4961 ( .A(n3477), .B(n3063), .Z(out[499]) );
  ANDN U4962 ( .B(n3065), .A(n3064), .Z(n3066) );
  XNOR U4963 ( .A(n3067), .B(n3066), .Z(out[49]) );
  OR U4964 ( .A(n3753), .B(n3068), .Z(n3069) );
  XNOR U4965 ( .A(n3752), .B(n3069), .Z(out[4]) );
  XNOR U4966 ( .A(in[874]), .B(n3725), .Z(n3481) );
  NAND U4967 ( .A(n3222), .B(n3070), .Z(n3071) );
  XNOR U4968 ( .A(n3481), .B(n3071), .Z(out[500]) );
  XNOR U4969 ( .A(in[875]), .B(n3729), .Z(n3485) );
  NAND U4970 ( .A(n3224), .B(n3072), .Z(n3073) );
  XNOR U4971 ( .A(n3485), .B(n3073), .Z(out[501]) );
  XNOR U4972 ( .A(in[876]), .B(n3733), .Z(n3493) );
  NAND U4973 ( .A(n3226), .B(n3074), .Z(n3075) );
  XNOR U4974 ( .A(n3493), .B(n3075), .Z(out[502]) );
  XNOR U4975 ( .A(in[877]), .B(n3737), .Z(n3497) );
  NAND U4976 ( .A(n3228), .B(n3076), .Z(n3077) );
  XNOR U4977 ( .A(n3497), .B(n3077), .Z(out[503]) );
  XNOR U4978 ( .A(in[878]), .B(n3741), .Z(n3501) );
  NAND U4979 ( .A(n3230), .B(n3078), .Z(n3079) );
  XNOR U4980 ( .A(n3501), .B(n3079), .Z(out[504]) );
  XNOR U4981 ( .A(in[879]), .B(n3745), .Z(n3505) );
  NAND U4982 ( .A(n3232), .B(n3080), .Z(n3081) );
  XNOR U4983 ( .A(n3505), .B(n3081), .Z(out[505]) );
  XNOR U4984 ( .A(in[880]), .B(n3749), .Z(n3509) );
  NAND U4985 ( .A(n3238), .B(n3082), .Z(n3083) );
  XNOR U4986 ( .A(n3509), .B(n3083), .Z(out[506]) );
  XNOR U4987 ( .A(in[881]), .B(n3757), .Z(n3513) );
  NAND U4988 ( .A(n3240), .B(n3084), .Z(n3085) );
  XNOR U4989 ( .A(n3513), .B(n3085), .Z(out[507]) );
  XNOR U4990 ( .A(in[882]), .B(n3761), .Z(n3517) );
  NAND U4991 ( .A(n3242), .B(n3086), .Z(n3087) );
  XNOR U4992 ( .A(n3517), .B(n3087), .Z(out[508]) );
  XNOR U4993 ( .A(in[883]), .B(n3765), .Z(n3521) );
  NAND U4994 ( .A(n3244), .B(n3088), .Z(n3089) );
  XNOR U4995 ( .A(n3521), .B(n3089), .Z(out[509]) );
  ANDN U4996 ( .B(n3091), .A(n3090), .Z(n3092) );
  XNOR U4997 ( .A(n3093), .B(n3092), .Z(out[50]) );
  XNOR U4998 ( .A(in[884]), .B(n3769), .Z(n3525) );
  NAND U4999 ( .A(n3246), .B(n3094), .Z(n3095) );
  XNOR U5000 ( .A(n3525), .B(n3095), .Z(out[510]) );
  XNOR U5001 ( .A(in[885]), .B(n3773), .Z(n3529) );
  NAND U5002 ( .A(n3248), .B(n3096), .Z(n3097) );
  XNOR U5003 ( .A(n3529), .B(n3097), .Z(out[511]) );
  OR U5004 ( .A(n3251), .B(n3098), .Z(n3099) );
  XNOR U5005 ( .A(n3250), .B(n3099), .Z(out[512]) );
  OR U5006 ( .A(n3255), .B(n3100), .Z(n3101) );
  XNOR U5007 ( .A(n3254), .B(n3101), .Z(out[513]) );
  OR U5008 ( .A(n3259), .B(n3102), .Z(n3103) );
  XNOR U5009 ( .A(n3258), .B(n3103), .Z(out[514]) );
  OR U5010 ( .A(n3263), .B(n3104), .Z(n3105) );
  XNOR U5011 ( .A(n3262), .B(n3105), .Z(out[515]) );
  OR U5012 ( .A(n3271), .B(n3106), .Z(n3107) );
  XNOR U5013 ( .A(n3270), .B(n3107), .Z(out[516]) );
  OR U5014 ( .A(n3275), .B(n3108), .Z(n3109) );
  XNOR U5015 ( .A(n3274), .B(n3109), .Z(out[517]) );
  OR U5016 ( .A(n3279), .B(n3110), .Z(n3111) );
  XNOR U5017 ( .A(n3278), .B(n3111), .Z(out[518]) );
  OR U5018 ( .A(n3283), .B(n3112), .Z(n3113) );
  XNOR U5019 ( .A(n3282), .B(n3113), .Z(out[519]) );
  ANDN U5020 ( .B(n3115), .A(n3114), .Z(n3116) );
  XNOR U5021 ( .A(n3117), .B(n3116), .Z(out[51]) );
  OR U5022 ( .A(n3287), .B(n3118), .Z(n3119) );
  XNOR U5023 ( .A(n3286), .B(n3119), .Z(out[520]) );
  OR U5024 ( .A(n3291), .B(n3120), .Z(n3121) );
  XNOR U5025 ( .A(n3290), .B(n3121), .Z(out[521]) );
  OR U5026 ( .A(n3295), .B(n3122), .Z(n3123) );
  XNOR U5027 ( .A(n3294), .B(n3123), .Z(out[522]) );
  OR U5028 ( .A(n3299), .B(n3124), .Z(n3125) );
  XNOR U5029 ( .A(n3298), .B(n3125), .Z(out[523]) );
  OR U5030 ( .A(n3303), .B(n3126), .Z(n3127) );
  XNOR U5031 ( .A(n3302), .B(n3127), .Z(out[524]) );
  OR U5032 ( .A(n3307), .B(n3128), .Z(n3129) );
  XNOR U5033 ( .A(n3306), .B(n3129), .Z(out[525]) );
  OR U5034 ( .A(n3315), .B(n3130), .Z(n3131) );
  XNOR U5035 ( .A(n3314), .B(n3131), .Z(out[526]) );
  OR U5036 ( .A(n3319), .B(n3132), .Z(n3133) );
  XNOR U5037 ( .A(n3318), .B(n3133), .Z(out[527]) );
  OR U5038 ( .A(n3323), .B(n3134), .Z(n3135) );
  XNOR U5039 ( .A(n3322), .B(n3135), .Z(out[528]) );
  OR U5040 ( .A(n3327), .B(n3136), .Z(n3137) );
  XNOR U5041 ( .A(n3326), .B(n3137), .Z(out[529]) );
  ANDN U5042 ( .B(n3139), .A(n3138), .Z(n3140) );
  XNOR U5043 ( .A(n3141), .B(n3140), .Z(out[52]) );
  OR U5044 ( .A(n3331), .B(n3142), .Z(n3143) );
  XNOR U5045 ( .A(n3330), .B(n3143), .Z(out[530]) );
  OR U5046 ( .A(n3335), .B(n3144), .Z(n3145) );
  XNOR U5047 ( .A(n3334), .B(n3145), .Z(out[531]) );
  OR U5048 ( .A(n3339), .B(n3146), .Z(n3147) );
  XNOR U5049 ( .A(n3338), .B(n3147), .Z(out[532]) );
  OR U5050 ( .A(n3343), .B(n3148), .Z(n3149) );
  XNOR U5051 ( .A(n3342), .B(n3149), .Z(out[533]) );
  OR U5052 ( .A(n3347), .B(n3150), .Z(n3151) );
  XNOR U5053 ( .A(n3346), .B(n3151), .Z(out[534]) );
  OR U5054 ( .A(n3351), .B(n3152), .Z(n3153) );
  XNOR U5055 ( .A(n3350), .B(n3153), .Z(out[535]) );
  OR U5056 ( .A(n3361), .B(n3154), .Z(n3155) );
  XNOR U5057 ( .A(n3360), .B(n3155), .Z(out[536]) );
  OR U5058 ( .A(n3365), .B(n3156), .Z(n3157) );
  XNOR U5059 ( .A(n3364), .B(n3157), .Z(out[537]) );
  OR U5060 ( .A(n3369), .B(n3158), .Z(n3159) );
  XNOR U5061 ( .A(n3368), .B(n3159), .Z(out[538]) );
  OR U5062 ( .A(n3373), .B(n3160), .Z(n3161) );
  XNOR U5063 ( .A(n3372), .B(n3161), .Z(out[539]) );
  ANDN U5064 ( .B(n3163), .A(n3162), .Z(n3164) );
  XNOR U5065 ( .A(n3165), .B(n3164), .Z(out[53]) );
  OR U5066 ( .A(n3377), .B(n3166), .Z(n3167) );
  XNOR U5067 ( .A(n3376), .B(n3167), .Z(out[540]) );
  OR U5068 ( .A(n3381), .B(n3168), .Z(n3169) );
  XNOR U5069 ( .A(n3380), .B(n3169), .Z(out[541]) );
  OR U5070 ( .A(n3385), .B(n3170), .Z(n3171) );
  XNOR U5071 ( .A(n3384), .B(n3171), .Z(out[542]) );
  OR U5072 ( .A(n3389), .B(n3172), .Z(n3173) );
  XNOR U5073 ( .A(n3388), .B(n3173), .Z(out[543]) );
  OR U5074 ( .A(n3393), .B(n3174), .Z(n3175) );
  XNOR U5075 ( .A(n3392), .B(n3175), .Z(out[544]) );
  OR U5076 ( .A(n3397), .B(n3176), .Z(n3177) );
  XNOR U5077 ( .A(n3396), .B(n3177), .Z(out[545]) );
  OR U5078 ( .A(n3405), .B(n3178), .Z(n3179) );
  XNOR U5079 ( .A(n3404), .B(n3179), .Z(out[546]) );
  OR U5080 ( .A(n3409), .B(n3180), .Z(n3181) );
  XNOR U5081 ( .A(n3408), .B(n3181), .Z(out[547]) );
  OR U5082 ( .A(n3413), .B(n3182), .Z(n3183) );
  XNOR U5083 ( .A(n3412), .B(n3183), .Z(out[548]) );
  OR U5084 ( .A(n3417), .B(n3184), .Z(n3185) );
  XNOR U5085 ( .A(n3416), .B(n3185), .Z(out[549]) );
  ANDN U5086 ( .B(n3187), .A(n3186), .Z(n3188) );
  XNOR U5087 ( .A(n3189), .B(n3188), .Z(out[54]) );
  OR U5088 ( .A(n3421), .B(n3190), .Z(n3191) );
  XNOR U5089 ( .A(n3420), .B(n3191), .Z(out[550]) );
  OR U5090 ( .A(n3425), .B(n3192), .Z(n3193) );
  XNOR U5091 ( .A(n3424), .B(n3193), .Z(out[551]) );
  OR U5092 ( .A(n3429), .B(n3194), .Z(n3195) );
  XNOR U5093 ( .A(n3428), .B(n3195), .Z(out[552]) );
  OR U5094 ( .A(n3433), .B(n3196), .Z(n3197) );
  XNOR U5095 ( .A(n3432), .B(n3197), .Z(out[553]) );
  OR U5096 ( .A(n3437), .B(n3198), .Z(n3199) );
  XNOR U5097 ( .A(n3436), .B(n3199), .Z(out[554]) );
  OR U5098 ( .A(n3441), .B(n3200), .Z(n3201) );
  XNOR U5099 ( .A(n3440), .B(n3201), .Z(out[555]) );
  OR U5100 ( .A(n3449), .B(n3202), .Z(n3203) );
  XNOR U5101 ( .A(n3448), .B(n3203), .Z(out[556]) );
  OR U5102 ( .A(n3453), .B(n3204), .Z(n3205) );
  XNOR U5103 ( .A(n3452), .B(n3205), .Z(out[557]) );
  OR U5104 ( .A(n3457), .B(n3206), .Z(n3207) );
  XNOR U5105 ( .A(n3456), .B(n3207), .Z(out[558]) );
  OR U5106 ( .A(n3461), .B(n3208), .Z(n3209) );
  XNOR U5107 ( .A(n3460), .B(n3209), .Z(out[559]) );
  ANDN U5108 ( .B(n3211), .A(n3210), .Z(n3212) );
  XNOR U5109 ( .A(n3213), .B(n3212), .Z(out[55]) );
  OR U5110 ( .A(n3465), .B(n3214), .Z(n3215) );
  XNOR U5111 ( .A(n3464), .B(n3215), .Z(out[560]) );
  OR U5112 ( .A(n3469), .B(n3216), .Z(n3217) );
  XNOR U5113 ( .A(n3468), .B(n3217), .Z(out[561]) );
  OR U5114 ( .A(n3473), .B(n3218), .Z(n3219) );
  XNOR U5115 ( .A(n3472), .B(n3219), .Z(out[562]) );
  OR U5116 ( .A(n3477), .B(n3220), .Z(n3221) );
  XNOR U5117 ( .A(n3476), .B(n3221), .Z(out[563]) );
  OR U5118 ( .A(n3481), .B(n3222), .Z(n3223) );
  XNOR U5119 ( .A(n3480), .B(n3223), .Z(out[564]) );
  OR U5120 ( .A(n3485), .B(n3224), .Z(n3225) );
  XNOR U5121 ( .A(n3484), .B(n3225), .Z(out[565]) );
  OR U5122 ( .A(n3493), .B(n3226), .Z(n3227) );
  XNOR U5123 ( .A(n3492), .B(n3227), .Z(out[566]) );
  OR U5124 ( .A(n3497), .B(n3228), .Z(n3229) );
  XNOR U5125 ( .A(n3496), .B(n3229), .Z(out[567]) );
  OR U5126 ( .A(n3501), .B(n3230), .Z(n3231) );
  XNOR U5127 ( .A(n3500), .B(n3231), .Z(out[568]) );
  OR U5128 ( .A(n3505), .B(n3232), .Z(n3233) );
  XNOR U5129 ( .A(n3504), .B(n3233), .Z(out[569]) );
  ANDN U5130 ( .B(n3235), .A(n3234), .Z(n3236) );
  XNOR U5131 ( .A(n3237), .B(n3236), .Z(out[56]) );
  OR U5132 ( .A(n3509), .B(n3238), .Z(n3239) );
  XNOR U5133 ( .A(n3508), .B(n3239), .Z(out[570]) );
  OR U5134 ( .A(n3513), .B(n3240), .Z(n3241) );
  XNOR U5135 ( .A(n3512), .B(n3241), .Z(out[571]) );
  OR U5136 ( .A(n3517), .B(n3242), .Z(n3243) );
  XNOR U5137 ( .A(n3516), .B(n3243), .Z(out[572]) );
  OR U5138 ( .A(n3521), .B(n3244), .Z(n3245) );
  XNOR U5139 ( .A(n3520), .B(n3245), .Z(out[573]) );
  OR U5140 ( .A(n3525), .B(n3246), .Z(n3247) );
  XNOR U5141 ( .A(n3524), .B(n3247), .Z(out[574]) );
  OR U5142 ( .A(n3529), .B(n3248), .Z(n3249) );
  XNOR U5143 ( .A(n3528), .B(n3249), .Z(out[575]) );
  ANDN U5144 ( .B(n3251), .A(n3250), .Z(n3252) );
  XNOR U5145 ( .A(n3253), .B(n3252), .Z(out[576]) );
  ANDN U5146 ( .B(n3255), .A(n3254), .Z(n3256) );
  XNOR U5147 ( .A(n3257), .B(n3256), .Z(out[577]) );
  ANDN U5148 ( .B(n3259), .A(n3258), .Z(n3260) );
  XNOR U5149 ( .A(n3261), .B(n3260), .Z(out[578]) );
  ANDN U5150 ( .B(n3263), .A(n3262), .Z(n3264) );
  XNOR U5151 ( .A(n3265), .B(n3264), .Z(out[579]) );
  ANDN U5152 ( .B(n3267), .A(n3266), .Z(n3268) );
  XNOR U5153 ( .A(n3269), .B(n3268), .Z(out[57]) );
  ANDN U5154 ( .B(n3271), .A(n3270), .Z(n3272) );
  XNOR U5155 ( .A(n3273), .B(n3272), .Z(out[580]) );
  ANDN U5156 ( .B(n3275), .A(n3274), .Z(n3276) );
  XNOR U5157 ( .A(n3277), .B(n3276), .Z(out[581]) );
  ANDN U5158 ( .B(n3279), .A(n3278), .Z(n3280) );
  XNOR U5159 ( .A(n3281), .B(n3280), .Z(out[582]) );
  ANDN U5160 ( .B(n3283), .A(n3282), .Z(n3284) );
  XNOR U5161 ( .A(n3285), .B(n3284), .Z(out[583]) );
  ANDN U5162 ( .B(n3287), .A(n3286), .Z(n3288) );
  XNOR U5163 ( .A(n3289), .B(n3288), .Z(out[584]) );
  ANDN U5164 ( .B(n3291), .A(n3290), .Z(n3292) );
  XNOR U5165 ( .A(n3293), .B(n3292), .Z(out[585]) );
  ANDN U5166 ( .B(n3295), .A(n3294), .Z(n3296) );
  XNOR U5167 ( .A(n3297), .B(n3296), .Z(out[586]) );
  ANDN U5168 ( .B(n3299), .A(n3298), .Z(n3300) );
  XNOR U5169 ( .A(n3301), .B(n3300), .Z(out[587]) );
  ANDN U5170 ( .B(n3303), .A(n3302), .Z(n3304) );
  XNOR U5171 ( .A(n3305), .B(n3304), .Z(out[588]) );
  ANDN U5172 ( .B(n3307), .A(n3306), .Z(n3308) );
  XNOR U5173 ( .A(n3309), .B(n3308), .Z(out[589]) );
  ANDN U5174 ( .B(n3311), .A(n3310), .Z(n3312) );
  XNOR U5175 ( .A(n3313), .B(n3312), .Z(out[58]) );
  ANDN U5176 ( .B(n3315), .A(n3314), .Z(n3316) );
  XNOR U5177 ( .A(n3317), .B(n3316), .Z(out[590]) );
  ANDN U5178 ( .B(n3319), .A(n3318), .Z(n3320) );
  XNOR U5179 ( .A(n3321), .B(n3320), .Z(out[591]) );
  ANDN U5180 ( .B(n3323), .A(n3322), .Z(n3324) );
  XNOR U5181 ( .A(n3325), .B(n3324), .Z(out[592]) );
  ANDN U5182 ( .B(n3327), .A(n3326), .Z(n3328) );
  XNOR U5183 ( .A(n3329), .B(n3328), .Z(out[593]) );
  ANDN U5184 ( .B(n3331), .A(n3330), .Z(n3332) );
  XNOR U5185 ( .A(n3333), .B(n3332), .Z(out[594]) );
  ANDN U5186 ( .B(n3335), .A(n3334), .Z(n3336) );
  XNOR U5187 ( .A(n3337), .B(n3336), .Z(out[595]) );
  ANDN U5188 ( .B(n3339), .A(n3338), .Z(n3340) );
  XNOR U5189 ( .A(n3341), .B(n3340), .Z(out[596]) );
  ANDN U5190 ( .B(n3343), .A(n3342), .Z(n3344) );
  XNOR U5191 ( .A(n3345), .B(n3344), .Z(out[597]) );
  ANDN U5192 ( .B(n3347), .A(n3346), .Z(n3348) );
  XNOR U5193 ( .A(n3349), .B(n3348), .Z(out[598]) );
  ANDN U5194 ( .B(n3351), .A(n3350), .Z(n3352) );
  XNOR U5195 ( .A(n3353), .B(n3352), .Z(out[599]) );
  ANDN U5196 ( .B(n3355), .A(n3354), .Z(n3356) );
  XNOR U5197 ( .A(n3357), .B(n3356), .Z(out[59]) );
  OR U5198 ( .A(n3797), .B(n3358), .Z(n3359) );
  XNOR U5199 ( .A(n3796), .B(n3359), .Z(out[5]) );
  ANDN U5200 ( .B(n3361), .A(n3360), .Z(n3362) );
  XNOR U5201 ( .A(n3363), .B(n3362), .Z(out[600]) );
  ANDN U5202 ( .B(n3365), .A(n3364), .Z(n3366) );
  XNOR U5203 ( .A(n3367), .B(n3366), .Z(out[601]) );
  ANDN U5204 ( .B(n3369), .A(n3368), .Z(n3370) );
  XNOR U5205 ( .A(n3371), .B(n3370), .Z(out[602]) );
  ANDN U5206 ( .B(n3373), .A(n3372), .Z(n3374) );
  XNOR U5207 ( .A(n3375), .B(n3374), .Z(out[603]) );
  ANDN U5208 ( .B(n3377), .A(n3376), .Z(n3378) );
  XNOR U5209 ( .A(n3379), .B(n3378), .Z(out[604]) );
  ANDN U5210 ( .B(n3381), .A(n3380), .Z(n3382) );
  XNOR U5211 ( .A(n3383), .B(n3382), .Z(out[605]) );
  ANDN U5212 ( .B(n3385), .A(n3384), .Z(n3386) );
  XNOR U5213 ( .A(n3387), .B(n3386), .Z(out[606]) );
  ANDN U5214 ( .B(n3389), .A(n3388), .Z(n3390) );
  XNOR U5215 ( .A(n3391), .B(n3390), .Z(out[607]) );
  ANDN U5216 ( .B(n3393), .A(n3392), .Z(n3394) );
  XNOR U5217 ( .A(n3395), .B(n3394), .Z(out[608]) );
  ANDN U5218 ( .B(n3397), .A(n3396), .Z(n3398) );
  XNOR U5219 ( .A(n3399), .B(n3398), .Z(out[609]) );
  ANDN U5220 ( .B(n3401), .A(n3400), .Z(n3402) );
  XNOR U5221 ( .A(n3403), .B(n3402), .Z(out[60]) );
  ANDN U5222 ( .B(n3405), .A(n3404), .Z(n3406) );
  XNOR U5223 ( .A(n3407), .B(n3406), .Z(out[610]) );
  ANDN U5224 ( .B(n3409), .A(n3408), .Z(n3410) );
  XNOR U5225 ( .A(n3411), .B(n3410), .Z(out[611]) );
  ANDN U5226 ( .B(n3413), .A(n3412), .Z(n3414) );
  XNOR U5227 ( .A(n3415), .B(n3414), .Z(out[612]) );
  ANDN U5228 ( .B(n3417), .A(n3416), .Z(n3418) );
  XNOR U5229 ( .A(n3419), .B(n3418), .Z(out[613]) );
  ANDN U5230 ( .B(n3421), .A(n3420), .Z(n3422) );
  XNOR U5231 ( .A(n3423), .B(n3422), .Z(out[614]) );
  ANDN U5232 ( .B(n3425), .A(n3424), .Z(n3426) );
  XNOR U5233 ( .A(n3427), .B(n3426), .Z(out[615]) );
  ANDN U5234 ( .B(n3429), .A(n3428), .Z(n3430) );
  XNOR U5235 ( .A(n3431), .B(n3430), .Z(out[616]) );
  ANDN U5236 ( .B(n3433), .A(n3432), .Z(n3434) );
  XNOR U5237 ( .A(n3435), .B(n3434), .Z(out[617]) );
  ANDN U5238 ( .B(n3437), .A(n3436), .Z(n3438) );
  XNOR U5239 ( .A(n3439), .B(n3438), .Z(out[618]) );
  ANDN U5240 ( .B(n3441), .A(n3440), .Z(n3442) );
  XNOR U5241 ( .A(n3443), .B(n3442), .Z(out[619]) );
  ANDN U5242 ( .B(n3445), .A(n3444), .Z(n3446) );
  XNOR U5243 ( .A(n3447), .B(n3446), .Z(out[61]) );
  ANDN U5244 ( .B(n3449), .A(n3448), .Z(n3450) );
  XNOR U5245 ( .A(n3451), .B(n3450), .Z(out[620]) );
  ANDN U5246 ( .B(n3453), .A(n3452), .Z(n3454) );
  XNOR U5247 ( .A(n3455), .B(n3454), .Z(out[621]) );
  ANDN U5248 ( .B(n3457), .A(n3456), .Z(n3458) );
  XNOR U5249 ( .A(n3459), .B(n3458), .Z(out[622]) );
  ANDN U5250 ( .B(n3461), .A(n3460), .Z(n3462) );
  XNOR U5251 ( .A(n3463), .B(n3462), .Z(out[623]) );
  ANDN U5252 ( .B(n3465), .A(n3464), .Z(n3466) );
  XNOR U5253 ( .A(n3467), .B(n3466), .Z(out[624]) );
  ANDN U5254 ( .B(n3469), .A(n3468), .Z(n3470) );
  XNOR U5255 ( .A(n3471), .B(n3470), .Z(out[625]) );
  ANDN U5256 ( .B(n3473), .A(n3472), .Z(n3474) );
  XNOR U5257 ( .A(n3475), .B(n3474), .Z(out[626]) );
  ANDN U5258 ( .B(n3477), .A(n3476), .Z(n3478) );
  XNOR U5259 ( .A(n3479), .B(n3478), .Z(out[627]) );
  ANDN U5260 ( .B(n3481), .A(n3480), .Z(n3482) );
  XNOR U5261 ( .A(n3483), .B(n3482), .Z(out[628]) );
  ANDN U5262 ( .B(n3485), .A(n3484), .Z(n3486) );
  XNOR U5263 ( .A(n3487), .B(n3486), .Z(out[629]) );
  ANDN U5264 ( .B(n3489), .A(n3488), .Z(n3490) );
  XNOR U5265 ( .A(n3491), .B(n3490), .Z(out[62]) );
  ANDN U5266 ( .B(n3493), .A(n3492), .Z(n3494) );
  XNOR U5267 ( .A(n3495), .B(n3494), .Z(out[630]) );
  ANDN U5268 ( .B(n3497), .A(n3496), .Z(n3498) );
  XNOR U5269 ( .A(n3499), .B(n3498), .Z(out[631]) );
  ANDN U5270 ( .B(n3501), .A(n3500), .Z(n3502) );
  XNOR U5271 ( .A(n3503), .B(n3502), .Z(out[632]) );
  ANDN U5272 ( .B(n3505), .A(n3504), .Z(n3506) );
  XNOR U5273 ( .A(n3507), .B(n3506), .Z(out[633]) );
  ANDN U5274 ( .B(n3509), .A(n3508), .Z(n3510) );
  XNOR U5275 ( .A(n3511), .B(n3510), .Z(out[634]) );
  ANDN U5276 ( .B(n3513), .A(n3512), .Z(n3514) );
  XNOR U5277 ( .A(n3515), .B(n3514), .Z(out[635]) );
  ANDN U5278 ( .B(n3517), .A(n3516), .Z(n3518) );
  XNOR U5279 ( .A(n3519), .B(n3518), .Z(out[636]) );
  ANDN U5280 ( .B(n3521), .A(n3520), .Z(n3522) );
  XNOR U5281 ( .A(n3523), .B(n3522), .Z(out[637]) );
  ANDN U5282 ( .B(n3525), .A(n3524), .Z(n3526) );
  XNOR U5283 ( .A(n3527), .B(n3526), .Z(out[638]) );
  ANDN U5284 ( .B(n3529), .A(n3528), .Z(n3530) );
  XNOR U5285 ( .A(n3531), .B(n3530), .Z(out[639]) );
  ANDN U5286 ( .B(n3533), .A(n3532), .Z(n3534) );
  XNOR U5287 ( .A(n3535), .B(n3534), .Z(out[63]) );
  XNOR U5288 ( .A(in[302]), .B(n3536), .Z(n3965) );
  XNOR U5289 ( .A(in[1535]), .B(n3537), .Z(n4343) );
  XNOR U5290 ( .A(in[1146]), .B(n3538), .Z(n4340) );
  NAND U5291 ( .A(n4343), .B(n4340), .Z(n3539) );
  XNOR U5292 ( .A(n3965), .B(n3539), .Z(out[640]) );
  XNOR U5293 ( .A(in[303]), .B(n3540), .Z(n3968) );
  XNOR U5294 ( .A(in[1472]), .B(n3541), .Z(n4347) );
  XNOR U5295 ( .A(in[1147]), .B(n3542), .Z(n4344) );
  NAND U5296 ( .A(n4347), .B(n4344), .Z(n3543) );
  XNOR U5297 ( .A(n3968), .B(n3543), .Z(out[641]) );
  XNOR U5298 ( .A(in[304]), .B(n3544), .Z(n3975) );
  XNOR U5299 ( .A(in[1473]), .B(n3545), .Z(n4351) );
  XNOR U5300 ( .A(in[1148]), .B(n3546), .Z(n4348) );
  NAND U5301 ( .A(n4351), .B(n4348), .Z(n3547) );
  XNOR U5302 ( .A(n3975), .B(n3547), .Z(out[642]) );
  XNOR U5303 ( .A(in[305]), .B(n3548), .Z(n3978) );
  XNOR U5304 ( .A(in[1474]), .B(n3549), .Z(n4355) );
  XNOR U5305 ( .A(in[1149]), .B(n3550), .Z(n4352) );
  NAND U5306 ( .A(n4355), .B(n4352), .Z(n3551) );
  XNOR U5307 ( .A(n3978), .B(n3551), .Z(out[643]) );
  XNOR U5308 ( .A(in[306]), .B(n3552), .Z(n3981) );
  XNOR U5309 ( .A(in[1475]), .B(n3553), .Z(n4367) );
  XNOR U5310 ( .A(in[1150]), .B(n3554), .Z(n4364) );
  NAND U5311 ( .A(n4367), .B(n4364), .Z(n3555) );
  XNOR U5312 ( .A(n3981), .B(n3555), .Z(out[644]) );
  XNOR U5313 ( .A(in[307]), .B(n3556), .Z(n3984) );
  XNOR U5314 ( .A(in[1476]), .B(n3557), .Z(n4371) );
  XNOR U5315 ( .A(in[1151]), .B(n3558), .Z(n4368) );
  NAND U5316 ( .A(n4371), .B(n4368), .Z(n3559) );
  XNOR U5317 ( .A(n3984), .B(n3559), .Z(out[645]) );
  XNOR U5318 ( .A(in[308]), .B(n3560), .Z(n3987) );
  XNOR U5319 ( .A(in[1477]), .B(n3561), .Z(n4375) );
  XNOR U5320 ( .A(in[1088]), .B(n3562), .Z(n4372) );
  NAND U5321 ( .A(n4375), .B(n4372), .Z(n3563) );
  XNOR U5322 ( .A(n3987), .B(n3563), .Z(out[646]) );
  XNOR U5323 ( .A(in[309]), .B(n3564), .Z(n3990) );
  XNOR U5324 ( .A(in[1478]), .B(n3565), .Z(n4379) );
  XNOR U5325 ( .A(in[1089]), .B(n3566), .Z(n4376) );
  NAND U5326 ( .A(n4379), .B(n4376), .Z(n3567) );
  XNOR U5327 ( .A(n3990), .B(n3567), .Z(out[647]) );
  XNOR U5328 ( .A(in[310]), .B(n3568), .Z(n3993) );
  XNOR U5329 ( .A(in[1479]), .B(n3569), .Z(n4383) );
  XOR U5330 ( .A(n3570), .B(in[1090]), .Z(n4380) );
  NAND U5331 ( .A(n4383), .B(n4380), .Z(n3571) );
  XNOR U5332 ( .A(n3993), .B(n3571), .Z(out[648]) );
  XNOR U5333 ( .A(in[311]), .B(n3572), .Z(n3996) );
  XNOR U5334 ( .A(in[1480]), .B(n3573), .Z(n4387) );
  XOR U5335 ( .A(n3574), .B(in[1091]), .Z(n4384) );
  NAND U5336 ( .A(n4387), .B(n4384), .Z(n3575) );
  XNOR U5337 ( .A(n3996), .B(n3575), .Z(out[649]) );
  NOR U5338 ( .A(n3577), .B(n3576), .Z(n3578) );
  XNOR U5339 ( .A(n3579), .B(n3578), .Z(out[64]) );
  XNOR U5340 ( .A(in[312]), .B(n3580), .Z(n3999) );
  XNOR U5341 ( .A(in[1481]), .B(n3581), .Z(n4391) );
  XOR U5342 ( .A(n3582), .B(in[1092]), .Z(n4388) );
  NAND U5343 ( .A(n4391), .B(n4388), .Z(n3583) );
  XNOR U5344 ( .A(n3999), .B(n3583), .Z(out[650]) );
  XNOR U5345 ( .A(in[313]), .B(n3584), .Z(n4002) );
  XNOR U5346 ( .A(in[1482]), .B(n3585), .Z(n4395) );
  XOR U5347 ( .A(n3586), .B(in[1093]), .Z(n4392) );
  NAND U5348 ( .A(n4395), .B(n4392), .Z(n3587) );
  XNOR U5349 ( .A(n4002), .B(n3587), .Z(out[651]) );
  XNOR U5350 ( .A(in[314]), .B(n3588), .Z(n4009) );
  XNOR U5351 ( .A(in[1483]), .B(n3589), .Z(n4399) );
  XOR U5352 ( .A(n3590), .B(in[1094]), .Z(n4396) );
  NAND U5353 ( .A(n4399), .B(n4396), .Z(n3591) );
  XNOR U5354 ( .A(n4009), .B(n3591), .Z(out[652]) );
  XNOR U5355 ( .A(in[315]), .B(n3592), .Z(n4012) );
  XNOR U5356 ( .A(in[1484]), .B(n3593), .Z(n4403) );
  XOR U5357 ( .A(n3594), .B(in[1095]), .Z(n4400) );
  NAND U5358 ( .A(n4403), .B(n4400), .Z(n3595) );
  XNOR U5359 ( .A(n4012), .B(n3595), .Z(out[653]) );
  XNOR U5360 ( .A(in[316]), .B(n3596), .Z(n4015) );
  XNOR U5361 ( .A(in[1485]), .B(n3597), .Z(n4411) );
  XOR U5362 ( .A(n3598), .B(in[1096]), .Z(n4408) );
  NAND U5363 ( .A(n4411), .B(n4408), .Z(n3599) );
  XNOR U5364 ( .A(n4015), .B(n3599), .Z(out[654]) );
  XNOR U5365 ( .A(in[317]), .B(n3600), .Z(n4018) );
  XNOR U5366 ( .A(in[1486]), .B(n3601), .Z(n4415) );
  XOR U5367 ( .A(in[1097]), .B(n3602), .Z(n4412) );
  NAND U5368 ( .A(n4415), .B(n4412), .Z(n3603) );
  XNOR U5369 ( .A(n4018), .B(n3603), .Z(out[655]) );
  XNOR U5370 ( .A(in[318]), .B(n3604), .Z(n4021) );
  XNOR U5371 ( .A(in[1487]), .B(n3605), .Z(n4419) );
  XOR U5372 ( .A(n3606), .B(in[1098]), .Z(n4416) );
  NAND U5373 ( .A(n4419), .B(n4416), .Z(n3607) );
  XNOR U5374 ( .A(n4021), .B(n3607), .Z(out[656]) );
  XNOR U5375 ( .A(in[319]), .B(n3608), .Z(n4024) );
  XNOR U5376 ( .A(in[1488]), .B(n3609), .Z(n4423) );
  XOR U5377 ( .A(n3610), .B(in[1099]), .Z(n4420) );
  NAND U5378 ( .A(n4423), .B(n4420), .Z(n3611) );
  XNOR U5379 ( .A(n4024), .B(n3611), .Z(out[657]) );
  XNOR U5380 ( .A(in[256]), .B(n3612), .Z(n4027) );
  XNOR U5381 ( .A(in[1489]), .B(n3613), .Z(n4427) );
  XOR U5382 ( .A(in[1100]), .B(n3614), .Z(n4424) );
  NAND U5383 ( .A(n4427), .B(n4424), .Z(n3615) );
  XNOR U5384 ( .A(n4027), .B(n3615), .Z(out[658]) );
  XNOR U5385 ( .A(in[257]), .B(n3616), .Z(n4030) );
  XNOR U5386 ( .A(in[1490]), .B(n3617), .Z(n4431) );
  XOR U5387 ( .A(in[1101]), .B(n3618), .Z(n4428) );
  NAND U5388 ( .A(n4431), .B(n4428), .Z(n3619) );
  XNOR U5389 ( .A(n4030), .B(n3619), .Z(out[659]) );
  NOR U5390 ( .A(n3621), .B(n3620), .Z(n3622) );
  XNOR U5391 ( .A(n3623), .B(n3622), .Z(out[65]) );
  XNOR U5392 ( .A(in[258]), .B(n3624), .Z(n4033) );
  XOR U5393 ( .A(in[1491]), .B(n3625), .Z(n4435) );
  XOR U5394 ( .A(in[1102]), .B(n3626), .Z(n4432) );
  NAND U5395 ( .A(n4435), .B(n4432), .Z(n3627) );
  XNOR U5396 ( .A(n4033), .B(n3627), .Z(out[660]) );
  XNOR U5397 ( .A(in[259]), .B(n3628), .Z(n4036) );
  XOR U5398 ( .A(in[1492]), .B(n3629), .Z(n4439) );
  XOR U5399 ( .A(in[1103]), .B(n3630), .Z(n4436) );
  NAND U5400 ( .A(n4439), .B(n4436), .Z(n3631) );
  XNOR U5401 ( .A(n4036), .B(n3631), .Z(out[661]) );
  XOR U5402 ( .A(in[260]), .B(n3632), .Z(n4043) );
  XOR U5403 ( .A(in[1493]), .B(n3633), .Z(n4443) );
  XOR U5404 ( .A(in[1104]), .B(n3634), .Z(n4440) );
  NAND U5405 ( .A(n4443), .B(n4440), .Z(n3635) );
  XNOR U5406 ( .A(n4043), .B(n3635), .Z(out[662]) );
  XOR U5407 ( .A(in[261]), .B(n3636), .Z(n4046) );
  XOR U5408 ( .A(in[1494]), .B(n3637), .Z(n4447) );
  XOR U5409 ( .A(in[1105]), .B(n3638), .Z(n4444) );
  NAND U5410 ( .A(n4447), .B(n4444), .Z(n3639) );
  XNOR U5411 ( .A(n4046), .B(n3639), .Z(out[663]) );
  XOR U5412 ( .A(in[262]), .B(n3640), .Z(n4049) );
  XOR U5413 ( .A(in[1495]), .B(n3641), .Z(n4455) );
  XOR U5414 ( .A(in[1106]), .B(n3642), .Z(n4452) );
  NAND U5415 ( .A(n4455), .B(n4452), .Z(n3643) );
  XNOR U5416 ( .A(n4049), .B(n3643), .Z(out[664]) );
  XOR U5417 ( .A(in[263]), .B(n3644), .Z(n4052) );
  XOR U5418 ( .A(in[1496]), .B(n3645), .Z(n4459) );
  XOR U5419 ( .A(in[1107]), .B(n3646), .Z(n4456) );
  NAND U5420 ( .A(n4459), .B(n4456), .Z(n3647) );
  XNOR U5421 ( .A(n4052), .B(n3647), .Z(out[665]) );
  XOR U5422 ( .A(in[264]), .B(n3648), .Z(n4055) );
  XOR U5423 ( .A(in[1497]), .B(n3649), .Z(n4463) );
  XOR U5424 ( .A(in[1108]), .B(n3650), .Z(n4460) );
  NAND U5425 ( .A(n4463), .B(n4460), .Z(n3651) );
  XNOR U5426 ( .A(n4055), .B(n3651), .Z(out[666]) );
  XOR U5427 ( .A(in[265]), .B(n3652), .Z(n4058) );
  XOR U5428 ( .A(in[1498]), .B(n3653), .Z(n4467) );
  XOR U5429 ( .A(in[1109]), .B(n3654), .Z(n4464) );
  NAND U5430 ( .A(n4467), .B(n4464), .Z(n3655) );
  XNOR U5431 ( .A(n4058), .B(n3655), .Z(out[667]) );
  XOR U5432 ( .A(in[266]), .B(n3656), .Z(n4061) );
  XOR U5433 ( .A(in[1499]), .B(n3657), .Z(n4471) );
  XOR U5434 ( .A(in[1110]), .B(n3658), .Z(n4468) );
  NAND U5435 ( .A(n4471), .B(n4468), .Z(n3659) );
  XNOR U5436 ( .A(n4061), .B(n3659), .Z(out[668]) );
  XOR U5437 ( .A(in[267]), .B(n3660), .Z(n4064) );
  XOR U5438 ( .A(in[1500]), .B(n3661), .Z(n4475) );
  XOR U5439 ( .A(in[1111]), .B(n3662), .Z(n4472) );
  NAND U5440 ( .A(n4475), .B(n4472), .Z(n3663) );
  XNOR U5441 ( .A(n4064), .B(n3663), .Z(out[669]) );
  ANDN U5442 ( .B(n3665), .A(n3664), .Z(n3666) );
  XNOR U5443 ( .A(n3667), .B(n3666), .Z(out[66]) );
  XOR U5444 ( .A(in[268]), .B(n3668), .Z(n4067) );
  XOR U5445 ( .A(in[1501]), .B(n3669), .Z(n4479) );
  XOR U5446 ( .A(in[1112]), .B(n3670), .Z(n4476) );
  NAND U5447 ( .A(n4479), .B(n4476), .Z(n3671) );
  XNOR U5448 ( .A(n4067), .B(n3671), .Z(out[670]) );
  XOR U5449 ( .A(in[269]), .B(n3672), .Z(n4070) );
  XOR U5450 ( .A(in[1502]), .B(n3673), .Z(n4483) );
  XOR U5451 ( .A(in[1113]), .B(n3674), .Z(n4480) );
  NAND U5452 ( .A(n4483), .B(n4480), .Z(n3675) );
  XNOR U5453 ( .A(n4070), .B(n3675), .Z(out[671]) );
  XOR U5454 ( .A(in[270]), .B(n3676), .Z(n4081) );
  XOR U5455 ( .A(in[1503]), .B(n3677), .Z(n4487) );
  XOR U5456 ( .A(in[1114]), .B(n3678), .Z(n4484) );
  NAND U5457 ( .A(n4487), .B(n4484), .Z(n3679) );
  XNOR U5458 ( .A(n4081), .B(n3679), .Z(out[672]) );
  XOR U5459 ( .A(in[271]), .B(n3680), .Z(n4084) );
  XOR U5460 ( .A(in[1504]), .B(n3681), .Z(n4491) );
  XOR U5461 ( .A(in[1115]), .B(n3682), .Z(n4488) );
  NAND U5462 ( .A(n4491), .B(n4488), .Z(n3683) );
  XNOR U5463 ( .A(n4084), .B(n3683), .Z(out[673]) );
  XOR U5464 ( .A(in[272]), .B(n3684), .Z(n4087) );
  XOR U5465 ( .A(in[1505]), .B(n3685), .Z(n4499) );
  XOR U5466 ( .A(in[1116]), .B(n3686), .Z(n4496) );
  NAND U5467 ( .A(n4499), .B(n4496), .Z(n3687) );
  XNOR U5468 ( .A(n4087), .B(n3687), .Z(out[674]) );
  XOR U5469 ( .A(in[273]), .B(n3688), .Z(n4090) );
  XNOR U5470 ( .A(n3689), .B(in[1506]), .Z(n4503) );
  XOR U5471 ( .A(in[1117]), .B(n3690), .Z(n4500) );
  NAND U5472 ( .A(n4503), .B(n4500), .Z(n3691) );
  XNOR U5473 ( .A(n4090), .B(n3691), .Z(out[675]) );
  XOR U5474 ( .A(in[274]), .B(n3692), .Z(n4093) );
  XNOR U5475 ( .A(n3693), .B(in[1507]), .Z(n4507) );
  XOR U5476 ( .A(in[1118]), .B(n3694), .Z(n4504) );
  NAND U5477 ( .A(n4507), .B(n4504), .Z(n3695) );
  XNOR U5478 ( .A(n4093), .B(n3695), .Z(out[676]) );
  XOR U5479 ( .A(in[275]), .B(n3696), .Z(n4096) );
  XNOR U5480 ( .A(n3697), .B(in[1508]), .Z(n4511) );
  XOR U5481 ( .A(in[1119]), .B(n3698), .Z(n4508) );
  NAND U5482 ( .A(n4511), .B(n4508), .Z(n3699) );
  XNOR U5483 ( .A(n4096), .B(n3699), .Z(out[677]) );
  XOR U5484 ( .A(in[276]), .B(n3700), .Z(n4099) );
  XNOR U5485 ( .A(n3701), .B(in[1509]), .Z(n4515) );
  XOR U5486 ( .A(in[1120]), .B(n3702), .Z(n4512) );
  NAND U5487 ( .A(n4515), .B(n4512), .Z(n3703) );
  XNOR U5488 ( .A(n4099), .B(n3703), .Z(out[678]) );
  XOR U5489 ( .A(in[277]), .B(n3704), .Z(n4102) );
  XOR U5490 ( .A(in[1510]), .B(n3705), .Z(n4519) );
  XOR U5491 ( .A(in[1121]), .B(n3706), .Z(n4516) );
  NAND U5492 ( .A(n4519), .B(n4516), .Z(n3707) );
  XNOR U5493 ( .A(n4102), .B(n3707), .Z(out[679]) );
  ANDN U5494 ( .B(n3709), .A(n3708), .Z(n3710) );
  XNOR U5495 ( .A(n3711), .B(n3710), .Z(out[67]) );
  XOR U5496 ( .A(in[278]), .B(n3712), .Z(n4105) );
  XOR U5497 ( .A(in[1511]), .B(n3713), .Z(n4523) );
  XOR U5498 ( .A(in[1122]), .B(n3714), .Z(n4520) );
  NAND U5499 ( .A(n4523), .B(n4520), .Z(n3715) );
  XNOR U5500 ( .A(n4105), .B(n3715), .Z(out[680]) );
  XOR U5501 ( .A(in[279]), .B(n3716), .Z(n4108) );
  XOR U5502 ( .A(in[1512]), .B(n3717), .Z(n4527) );
  XOR U5503 ( .A(in[1123]), .B(n3718), .Z(n4524) );
  NAND U5504 ( .A(n4527), .B(n4524), .Z(n3719) );
  XNOR U5505 ( .A(n4108), .B(n3719), .Z(out[681]) );
  XOR U5506 ( .A(in[280]), .B(n3720), .Z(n4115) );
  XOR U5507 ( .A(in[1513]), .B(n3721), .Z(n4531) );
  XOR U5508 ( .A(in[1124]), .B(n3722), .Z(n4528) );
  NAND U5509 ( .A(n4531), .B(n4528), .Z(n3723) );
  XNOR U5510 ( .A(n4115), .B(n3723), .Z(out[682]) );
  XOR U5511 ( .A(in[281]), .B(n3724), .Z(n4118) );
  XOR U5512 ( .A(in[1514]), .B(n3725), .Z(n4535) );
  XOR U5513 ( .A(in[1125]), .B(n3726), .Z(n4532) );
  NAND U5514 ( .A(n4535), .B(n4532), .Z(n3727) );
  XNOR U5515 ( .A(n4118), .B(n3727), .Z(out[683]) );
  XOR U5516 ( .A(in[282]), .B(n3728), .Z(n4121) );
  XOR U5517 ( .A(in[1515]), .B(n3729), .Z(n4543) );
  XNOR U5518 ( .A(in[1126]), .B(n3730), .Z(n4540) );
  NAND U5519 ( .A(n4543), .B(n4540), .Z(n3731) );
  XNOR U5520 ( .A(n4121), .B(n3731), .Z(out[684]) );
  XOR U5521 ( .A(in[283]), .B(n3732), .Z(n4124) );
  XOR U5522 ( .A(in[1516]), .B(n3733), .Z(n4547) );
  XNOR U5523 ( .A(in[1127]), .B(n3734), .Z(n4544) );
  NAND U5524 ( .A(n4547), .B(n4544), .Z(n3735) );
  XNOR U5525 ( .A(n4124), .B(n3735), .Z(out[685]) );
  XOR U5526 ( .A(in[284]), .B(n3736), .Z(n4127) );
  XOR U5527 ( .A(in[1517]), .B(n3737), .Z(n4551) );
  XNOR U5528 ( .A(in[1128]), .B(n3738), .Z(n4548) );
  NAND U5529 ( .A(n4551), .B(n4548), .Z(n3739) );
  XNOR U5530 ( .A(n4127), .B(n3739), .Z(out[686]) );
  XOR U5531 ( .A(in[285]), .B(n3740), .Z(n4130) );
  XOR U5532 ( .A(in[1518]), .B(n3741), .Z(n4555) );
  XNOR U5533 ( .A(in[1129]), .B(n3742), .Z(n4552) );
  NAND U5534 ( .A(n4555), .B(n4552), .Z(n3743) );
  XNOR U5535 ( .A(n4130), .B(n3743), .Z(out[687]) );
  XOR U5536 ( .A(in[286]), .B(n3744), .Z(n4133) );
  XOR U5537 ( .A(in[1519]), .B(n3745), .Z(n4559) );
  XNOR U5538 ( .A(in[1130]), .B(n3746), .Z(n4556) );
  NAND U5539 ( .A(n4559), .B(n4556), .Z(n3747) );
  XNOR U5540 ( .A(n4133), .B(n3747), .Z(out[688]) );
  XOR U5541 ( .A(in[287]), .B(n3748), .Z(n4136) );
  XOR U5542 ( .A(in[1520]), .B(n3749), .Z(n4563) );
  XNOR U5543 ( .A(in[1131]), .B(n3750), .Z(n4560) );
  NAND U5544 ( .A(n4563), .B(n4560), .Z(n3751) );
  XNOR U5545 ( .A(n4136), .B(n3751), .Z(out[689]) );
  ANDN U5546 ( .B(n3753), .A(n3752), .Z(n3754) );
  XNOR U5547 ( .A(n3755), .B(n3754), .Z(out[68]) );
  XOR U5548 ( .A(in[288]), .B(n3756), .Z(n4139) );
  XOR U5549 ( .A(in[1521]), .B(n3757), .Z(n4567) );
  XNOR U5550 ( .A(in[1132]), .B(n3758), .Z(n4564) );
  NAND U5551 ( .A(n4567), .B(n4564), .Z(n3759) );
  XNOR U5552 ( .A(n4139), .B(n3759), .Z(out[690]) );
  XOR U5553 ( .A(in[289]), .B(n3760), .Z(n4142) );
  XOR U5554 ( .A(in[1522]), .B(n3761), .Z(n4571) );
  XNOR U5555 ( .A(in[1133]), .B(n3762), .Z(n4568) );
  NAND U5556 ( .A(n4571), .B(n4568), .Z(n3763) );
  XNOR U5557 ( .A(n4142), .B(n3763), .Z(out[691]) );
  XOR U5558 ( .A(in[290]), .B(n3764), .Z(n4149) );
  XOR U5559 ( .A(in[1523]), .B(n3765), .Z(n4575) );
  XNOR U5560 ( .A(in[1134]), .B(n3766), .Z(n4572) );
  NAND U5561 ( .A(n4575), .B(n4572), .Z(n3767) );
  XNOR U5562 ( .A(n4149), .B(n3767), .Z(out[692]) );
  XOR U5563 ( .A(in[291]), .B(n3768), .Z(n4152) );
  XOR U5564 ( .A(in[1524]), .B(n3769), .Z(n4579) );
  XNOR U5565 ( .A(in[1135]), .B(n3770), .Z(n4576) );
  NAND U5566 ( .A(n4579), .B(n4576), .Z(n3771) );
  XNOR U5567 ( .A(n4152), .B(n3771), .Z(out[693]) );
  XOR U5568 ( .A(in[292]), .B(n3772), .Z(n4155) );
  XOR U5569 ( .A(in[1525]), .B(n3773), .Z(n4587) );
  XNOR U5570 ( .A(in[1136]), .B(n3774), .Z(n4584) );
  NAND U5571 ( .A(n4587), .B(n4584), .Z(n3775) );
  XNOR U5572 ( .A(n4155), .B(n3775), .Z(out[694]) );
  XNOR U5573 ( .A(in[293]), .B(n3776), .Z(n4158) );
  XOR U5574 ( .A(in[1526]), .B(n3777), .Z(n4591) );
  XNOR U5575 ( .A(in[1137]), .B(n3778), .Z(n4588) );
  NAND U5576 ( .A(n4591), .B(n4588), .Z(n3779) );
  XNOR U5577 ( .A(n4158), .B(n3779), .Z(out[695]) );
  XNOR U5578 ( .A(in[294]), .B(n3780), .Z(n4161) );
  XOR U5579 ( .A(in[1527]), .B(n3781), .Z(n4595) );
  XNOR U5580 ( .A(in[1138]), .B(n3782), .Z(n4592) );
  NAND U5581 ( .A(n4595), .B(n4592), .Z(n3783) );
  XNOR U5582 ( .A(n4161), .B(n3783), .Z(out[696]) );
  XNOR U5583 ( .A(in[295]), .B(n3784), .Z(n4164) );
  XOR U5584 ( .A(in[1528]), .B(n3785), .Z(n4599) );
  XNOR U5585 ( .A(in[1139]), .B(n3786), .Z(n4596) );
  NAND U5586 ( .A(n4599), .B(n4596), .Z(n3787) );
  XNOR U5587 ( .A(n4164), .B(n3787), .Z(out[697]) );
  XNOR U5588 ( .A(in[296]), .B(n3788), .Z(n4167) );
  XOR U5589 ( .A(in[1529]), .B(n3789), .Z(n4603) );
  XNOR U5590 ( .A(in[1140]), .B(n3790), .Z(n4600) );
  NAND U5591 ( .A(n4603), .B(n4600), .Z(n3791) );
  XNOR U5592 ( .A(n4167), .B(n3791), .Z(out[698]) );
  XNOR U5593 ( .A(in[297]), .B(n3792), .Z(n4170) );
  XOR U5594 ( .A(in[1530]), .B(n3793), .Z(n4607) );
  XNOR U5595 ( .A(in[1141]), .B(n3794), .Z(n4604) );
  NAND U5596 ( .A(n4607), .B(n4604), .Z(n3795) );
  XNOR U5597 ( .A(n4170), .B(n3795), .Z(out[699]) );
  ANDN U5598 ( .B(n3797), .A(n3796), .Z(n3798) );
  XNOR U5599 ( .A(n3799), .B(n3798), .Z(out[69]) );
  OR U5600 ( .A(n3831), .B(n3800), .Z(n3801) );
  XNOR U5601 ( .A(n3830), .B(n3801), .Z(out[6]) );
  XNOR U5602 ( .A(in[298]), .B(n3802), .Z(n4173) );
  XNOR U5603 ( .A(in[1531]), .B(n3803), .Z(n4611) );
  XNOR U5604 ( .A(in[1142]), .B(n3804), .Z(n4608) );
  NAND U5605 ( .A(n4611), .B(n4608), .Z(n3805) );
  XNOR U5606 ( .A(n4173), .B(n3805), .Z(out[700]) );
  XNOR U5607 ( .A(in[299]), .B(n3806), .Z(n4176) );
  XNOR U5608 ( .A(in[1532]), .B(n3807), .Z(n4615) );
  XNOR U5609 ( .A(in[1143]), .B(n3808), .Z(n4612) );
  NAND U5610 ( .A(n4615), .B(n4612), .Z(n3809) );
  XNOR U5611 ( .A(n4176), .B(n3809), .Z(out[701]) );
  XNOR U5612 ( .A(in[300]), .B(n3810), .Z(n4183) );
  XNOR U5613 ( .A(in[1533]), .B(n3811), .Z(n4619) );
  XNOR U5614 ( .A(in[1144]), .B(n3812), .Z(n4616) );
  NAND U5615 ( .A(n4619), .B(n4616), .Z(n3813) );
  XNOR U5616 ( .A(n4183), .B(n3813), .Z(out[702]) );
  XNOR U5617 ( .A(in[301]), .B(n3814), .Z(n4186) );
  XOR U5618 ( .A(in[1534]), .B(n3815), .Z(n4623) );
  XNOR U5619 ( .A(in[1145]), .B(n3816), .Z(n4620) );
  NAND U5620 ( .A(n4623), .B(n4620), .Z(n3817) );
  XNOR U5621 ( .A(n4186), .B(n3817), .Z(out[703]) );
  XOR U5622 ( .A(in[376]), .B(n3818), .Z(n4188) );
  NOR U5623 ( .A(n3965), .B(n4343), .Z(n3819) );
  XNOR U5624 ( .A(n4188), .B(n3819), .Z(out[704]) );
  XOR U5625 ( .A(in[377]), .B(n3820), .Z(n4190) );
  NOR U5626 ( .A(n3968), .B(n4347), .Z(n3821) );
  XNOR U5627 ( .A(n4190), .B(n3821), .Z(out[705]) );
  XOR U5628 ( .A(in[378]), .B(n3822), .Z(n4192) );
  NOR U5629 ( .A(n3975), .B(n4351), .Z(n3823) );
  XNOR U5630 ( .A(n4192), .B(n3823), .Z(out[706]) );
  XOR U5631 ( .A(in[379]), .B(n3824), .Z(n4194) );
  NOR U5632 ( .A(n3978), .B(n4355), .Z(n3825) );
  XNOR U5633 ( .A(n4194), .B(n3825), .Z(out[707]) );
  XOR U5634 ( .A(in[380]), .B(n3826), .Z(n4196) );
  NOR U5635 ( .A(n3981), .B(n4367), .Z(n3827) );
  XNOR U5636 ( .A(n4196), .B(n3827), .Z(out[708]) );
  XOR U5637 ( .A(in[381]), .B(n3828), .Z(n4198) );
  NOR U5638 ( .A(n3984), .B(n4371), .Z(n3829) );
  XNOR U5639 ( .A(n4198), .B(n3829), .Z(out[709]) );
  ANDN U5640 ( .B(n3831), .A(n3830), .Z(n3832) );
  XNOR U5641 ( .A(n3833), .B(n3832), .Z(out[70]) );
  XOR U5642 ( .A(in[382]), .B(n3834), .Z(n4200) );
  NOR U5643 ( .A(n3987), .B(n4375), .Z(n3835) );
  XNOR U5644 ( .A(n4200), .B(n3835), .Z(out[710]) );
  XOR U5645 ( .A(in[383]), .B(n3836), .Z(n4202) );
  NOR U5646 ( .A(n3990), .B(n4379), .Z(n3837) );
  XNOR U5647 ( .A(n4202), .B(n3837), .Z(out[711]) );
  XOR U5648 ( .A(in[320]), .B(n3838), .Z(n4208) );
  NOR U5649 ( .A(n3993), .B(n4383), .Z(n3839) );
  XNOR U5650 ( .A(n4208), .B(n3839), .Z(out[712]) );
  XOR U5651 ( .A(in[321]), .B(n3840), .Z(n4210) );
  NOR U5652 ( .A(n3996), .B(n4387), .Z(n3841) );
  XNOR U5653 ( .A(n4210), .B(n3841), .Z(out[713]) );
  XOR U5654 ( .A(in[322]), .B(n3842), .Z(n4212) );
  NOR U5655 ( .A(n3999), .B(n4391), .Z(n3843) );
  XNOR U5656 ( .A(n4212), .B(n3843), .Z(out[714]) );
  XOR U5657 ( .A(in[323]), .B(n3844), .Z(n4214) );
  NOR U5658 ( .A(n4002), .B(n4395), .Z(n3845) );
  XNOR U5659 ( .A(n4214), .B(n3845), .Z(out[715]) );
  XOR U5660 ( .A(in[324]), .B(n3846), .Z(n4216) );
  NOR U5661 ( .A(n4009), .B(n4399), .Z(n3847) );
  XNOR U5662 ( .A(n4216), .B(n3847), .Z(out[716]) );
  XOR U5663 ( .A(in[325]), .B(n3848), .Z(n4218) );
  NOR U5664 ( .A(n4012), .B(n4403), .Z(n3849) );
  XNOR U5665 ( .A(n4218), .B(n3849), .Z(out[717]) );
  XOR U5666 ( .A(in[326]), .B(n3850), .Z(n4220) );
  NOR U5667 ( .A(n4015), .B(n4411), .Z(n3851) );
  XNOR U5668 ( .A(n4220), .B(n3851), .Z(out[718]) );
  XOR U5669 ( .A(in[327]), .B(n3852), .Z(n4222) );
  NOR U5670 ( .A(n4018), .B(n4415), .Z(n3853) );
  XNOR U5671 ( .A(n4222), .B(n3853), .Z(out[719]) );
  ANDN U5672 ( .B(n4077), .A(n4079), .Z(n3854) );
  XNOR U5673 ( .A(n3855), .B(n3854), .Z(out[71]) );
  XOR U5674 ( .A(in[328]), .B(n3856), .Z(n4224) );
  NOR U5675 ( .A(n4021), .B(n4419), .Z(n3857) );
  XNOR U5676 ( .A(n4224), .B(n3857), .Z(out[720]) );
  XOR U5677 ( .A(in[329]), .B(n3858), .Z(n4226) );
  NOR U5678 ( .A(n4024), .B(n4423), .Z(n3859) );
  XNOR U5679 ( .A(n4226), .B(n3859), .Z(out[721]) );
  XOR U5680 ( .A(in[330]), .B(n3860), .Z(n4232) );
  NOR U5681 ( .A(n4027), .B(n4427), .Z(n3861) );
  XNOR U5682 ( .A(n4232), .B(n3861), .Z(out[722]) );
  XOR U5683 ( .A(in[331]), .B(n3862), .Z(n4234) );
  NOR U5684 ( .A(n4030), .B(n4431), .Z(n3863) );
  XNOR U5685 ( .A(n4234), .B(n3863), .Z(out[723]) );
  XOR U5686 ( .A(in[332]), .B(n3864), .Z(n4236) );
  NOR U5687 ( .A(n4033), .B(n4435), .Z(n3865) );
  XNOR U5688 ( .A(n4236), .B(n3865), .Z(out[724]) );
  XOR U5689 ( .A(in[333]), .B(n3866), .Z(n4238) );
  NOR U5690 ( .A(n4036), .B(n4439), .Z(n3867) );
  XNOR U5691 ( .A(n4238), .B(n3867), .Z(out[725]) );
  XOR U5692 ( .A(in[334]), .B(n3868), .Z(n4240) );
  NOR U5693 ( .A(n4043), .B(n4443), .Z(n3869) );
  XNOR U5694 ( .A(n4240), .B(n3869), .Z(out[726]) );
  XOR U5695 ( .A(in[335]), .B(n3870), .Z(n4242) );
  NOR U5696 ( .A(n4046), .B(n4447), .Z(n3871) );
  XNOR U5697 ( .A(n4242), .B(n3871), .Z(out[727]) );
  XOR U5698 ( .A(in[336]), .B(n3872), .Z(n4244) );
  NOR U5699 ( .A(n4049), .B(n4455), .Z(n3873) );
  XNOR U5700 ( .A(n4244), .B(n3873), .Z(out[728]) );
  XOR U5701 ( .A(in[337]), .B(n3874), .Z(n4246) );
  NOR U5702 ( .A(n4052), .B(n4459), .Z(n3875) );
  XNOR U5703 ( .A(n4246), .B(n3875), .Z(out[729]) );
  ANDN U5704 ( .B(n4361), .A(n4363), .Z(n3876) );
  XNOR U5705 ( .A(n3877), .B(n3876), .Z(out[72]) );
  XOR U5706 ( .A(in[338]), .B(n3878), .Z(n4248) );
  NOR U5707 ( .A(n4055), .B(n4463), .Z(n3879) );
  XNOR U5708 ( .A(n4248), .B(n3879), .Z(out[730]) );
  XOR U5709 ( .A(in[339]), .B(n3880), .Z(n4250) );
  NOR U5710 ( .A(n4058), .B(n4467), .Z(n3881) );
  XNOR U5711 ( .A(n4250), .B(n3881), .Z(out[731]) );
  XOR U5712 ( .A(in[340]), .B(n3882), .Z(n4256) );
  NOR U5713 ( .A(n4061), .B(n4471), .Z(n3883) );
  XNOR U5714 ( .A(n4256), .B(n3883), .Z(out[732]) );
  XOR U5715 ( .A(in[341]), .B(n3884), .Z(n4258) );
  NOR U5716 ( .A(n4064), .B(n4475), .Z(n3885) );
  XNOR U5717 ( .A(n4258), .B(n3885), .Z(out[733]) );
  XOR U5718 ( .A(in[342]), .B(n3886), .Z(n4260) );
  NOR U5719 ( .A(n4067), .B(n4479), .Z(n3887) );
  XNOR U5720 ( .A(n4260), .B(n3887), .Z(out[734]) );
  XOR U5721 ( .A(in[343]), .B(n3888), .Z(n4262) );
  NOR U5722 ( .A(n4070), .B(n4483), .Z(n3889) );
  XNOR U5723 ( .A(n4262), .B(n3889), .Z(out[735]) );
  XOR U5724 ( .A(in[344]), .B(n3890), .Z(n4264) );
  NOR U5725 ( .A(n4081), .B(n4487), .Z(n3891) );
  XNOR U5726 ( .A(n4264), .B(n3891), .Z(out[736]) );
  XOR U5727 ( .A(in[345]), .B(n3892), .Z(n4266) );
  NOR U5728 ( .A(n4084), .B(n4491), .Z(n3893) );
  XNOR U5729 ( .A(n4266), .B(n3893), .Z(out[737]) );
  XOR U5730 ( .A(in[346]), .B(n3894), .Z(n4268) );
  NOR U5731 ( .A(n4087), .B(n4499), .Z(n3895) );
  XNOR U5732 ( .A(n4268), .B(n3895), .Z(out[738]) );
  XOR U5733 ( .A(in[347]), .B(n3896), .Z(n4270) );
  NOR U5734 ( .A(n4090), .B(n4503), .Z(n3897) );
  XNOR U5735 ( .A(n4270), .B(n3897), .Z(out[739]) );
  ANDN U5736 ( .B(n4805), .A(n4807), .Z(n3898) );
  XNOR U5737 ( .A(n3899), .B(n3898), .Z(out[73]) );
  XOR U5738 ( .A(in[348]), .B(n3900), .Z(n4272) );
  NOR U5739 ( .A(n4093), .B(n4507), .Z(n3901) );
  XNOR U5740 ( .A(n4272), .B(n3901), .Z(out[740]) );
  XOR U5741 ( .A(in[349]), .B(n3902), .Z(n4274) );
  NOR U5742 ( .A(n4096), .B(n4511), .Z(n3903) );
  XNOR U5743 ( .A(n4274), .B(n3903), .Z(out[741]) );
  XOR U5744 ( .A(in[350]), .B(n3904), .Z(n4280) );
  NOR U5745 ( .A(n4099), .B(n4515), .Z(n3905) );
  XNOR U5746 ( .A(n4280), .B(n3905), .Z(out[742]) );
  XOR U5747 ( .A(in[351]), .B(n3906), .Z(n4282) );
  NOR U5748 ( .A(n4102), .B(n4519), .Z(n3907) );
  XNOR U5749 ( .A(n4282), .B(n3907), .Z(out[743]) );
  XOR U5750 ( .A(in[352]), .B(n3908), .Z(n4284) );
  NOR U5751 ( .A(n4105), .B(n4523), .Z(n3909) );
  XNOR U5752 ( .A(n4284), .B(n3909), .Z(out[744]) );
  XOR U5753 ( .A(in[353]), .B(n3910), .Z(n4286) );
  NOR U5754 ( .A(n4108), .B(n4527), .Z(n3911) );
  XNOR U5755 ( .A(n4286), .B(n3911), .Z(out[745]) );
  XOR U5756 ( .A(in[354]), .B(n3912), .Z(n4288) );
  NOR U5757 ( .A(n4115), .B(n4531), .Z(n3913) );
  XNOR U5758 ( .A(n4288), .B(n3913), .Z(out[746]) );
  XOR U5759 ( .A(in[355]), .B(n3914), .Z(n4290) );
  NOR U5760 ( .A(n4118), .B(n4535), .Z(n3915) );
  XNOR U5761 ( .A(n4290), .B(n3915), .Z(out[747]) );
  XOR U5762 ( .A(in[356]), .B(n3916), .Z(n4292) );
  NOR U5763 ( .A(n4121), .B(n4543), .Z(n3917) );
  XNOR U5764 ( .A(n4292), .B(n3917), .Z(out[748]) );
  XOR U5765 ( .A(in[357]), .B(n3918), .Z(n4294) );
  NOR U5766 ( .A(n4124), .B(n4547), .Z(n3919) );
  XNOR U5767 ( .A(n4294), .B(n3919), .Z(out[749]) );
  NOR U5768 ( .A(n3921), .B(n3920), .Z(n3922) );
  XNOR U5769 ( .A(n3923), .B(n3922), .Z(out[74]) );
  XOR U5770 ( .A(in[358]), .B(n3924), .Z(n4296) );
  NOR U5771 ( .A(n4127), .B(n4551), .Z(n3925) );
  XNOR U5772 ( .A(n4296), .B(n3925), .Z(out[750]) );
  XOR U5773 ( .A(in[359]), .B(n3926), .Z(n4298) );
  NOR U5774 ( .A(n4130), .B(n4555), .Z(n3927) );
  XNOR U5775 ( .A(n4298), .B(n3927), .Z(out[751]) );
  XOR U5776 ( .A(in[360]), .B(n3928), .Z(n4304) );
  NOR U5777 ( .A(n4133), .B(n4559), .Z(n3929) );
  XNOR U5778 ( .A(n4304), .B(n3929), .Z(out[752]) );
  XOR U5779 ( .A(in[361]), .B(n3930), .Z(n4306) );
  NOR U5780 ( .A(n4136), .B(n4563), .Z(n3931) );
  XNOR U5781 ( .A(n4306), .B(n3931), .Z(out[753]) );
  XOR U5782 ( .A(in[362]), .B(n3932), .Z(n4308) );
  NOR U5783 ( .A(n4139), .B(n4567), .Z(n3933) );
  XNOR U5784 ( .A(n4308), .B(n3933), .Z(out[754]) );
  XOR U5785 ( .A(in[363]), .B(n3934), .Z(n4310) );
  NOR U5786 ( .A(n4142), .B(n4571), .Z(n3935) );
  XNOR U5787 ( .A(n4310), .B(n3935), .Z(out[755]) );
  XOR U5788 ( .A(in[364]), .B(n3936), .Z(n4312) );
  NOR U5789 ( .A(n4149), .B(n4575), .Z(n3937) );
  XNOR U5790 ( .A(n4312), .B(n3937), .Z(out[756]) );
  XOR U5791 ( .A(in[365]), .B(n3938), .Z(n4314) );
  NOR U5792 ( .A(n4152), .B(n4579), .Z(n3939) );
  XNOR U5793 ( .A(n4314), .B(n3939), .Z(out[757]) );
  XOR U5794 ( .A(in[366]), .B(n3940), .Z(n4316) );
  NOR U5795 ( .A(n4155), .B(n4587), .Z(n3941) );
  XNOR U5796 ( .A(n4316), .B(n3941), .Z(out[758]) );
  XOR U5797 ( .A(in[367]), .B(n3942), .Z(n4318) );
  NOR U5798 ( .A(n4158), .B(n4591), .Z(n3943) );
  XNOR U5799 ( .A(n4318), .B(n3943), .Z(out[759]) );
  NOR U5800 ( .A(n3945), .B(n3944), .Z(n3946) );
  XNOR U5801 ( .A(n3947), .B(n3946), .Z(out[75]) );
  XOR U5802 ( .A(in[368]), .B(n3948), .Z(n4320) );
  NOR U5803 ( .A(n4161), .B(n4595), .Z(n3949) );
  XNOR U5804 ( .A(n4320), .B(n3949), .Z(out[760]) );
  XOR U5805 ( .A(in[369]), .B(n3950), .Z(n4322) );
  NOR U5806 ( .A(n4164), .B(n4599), .Z(n3951) );
  XNOR U5807 ( .A(n4322), .B(n3951), .Z(out[761]) );
  XOR U5808 ( .A(in[370]), .B(n3952), .Z(n4328) );
  NOR U5809 ( .A(n4167), .B(n4603), .Z(n3953) );
  XNOR U5810 ( .A(n4328), .B(n3953), .Z(out[762]) );
  XOR U5811 ( .A(in[371]), .B(n3954), .Z(n4330) );
  NOR U5812 ( .A(n4170), .B(n4607), .Z(n3955) );
  XNOR U5813 ( .A(n4330), .B(n3955), .Z(out[763]) );
  XOR U5814 ( .A(in[372]), .B(n3956), .Z(n4332) );
  NOR U5815 ( .A(n4173), .B(n4611), .Z(n3957) );
  XNOR U5816 ( .A(n4332), .B(n3957), .Z(out[764]) );
  XOR U5817 ( .A(in[373]), .B(n3958), .Z(n4334) );
  NOR U5818 ( .A(n4176), .B(n4615), .Z(n3959) );
  XNOR U5819 ( .A(n4334), .B(n3959), .Z(out[765]) );
  XOR U5820 ( .A(in[374]), .B(n3960), .Z(n4336) );
  NOR U5821 ( .A(n4183), .B(n4619), .Z(n3961) );
  XNOR U5822 ( .A(n4336), .B(n3961), .Z(out[766]) );
  XOR U5823 ( .A(in[375]), .B(n3962), .Z(n4338) );
  NOR U5824 ( .A(n4186), .B(n4623), .Z(n3963) );
  XNOR U5825 ( .A(n4338), .B(n3963), .Z(out[767]) );
  XNOR U5826 ( .A(in[743]), .B(n3964), .Z(n4341) );
  NAND U5827 ( .A(n4188), .B(n3965), .Z(n3966) );
  XNOR U5828 ( .A(n4341), .B(n3966), .Z(out[768]) );
  XNOR U5829 ( .A(in[744]), .B(n3967), .Z(n4345) );
  NAND U5830 ( .A(n4190), .B(n3968), .Z(n3969) );
  XNOR U5831 ( .A(n4345), .B(n3969), .Z(out[769]) );
  NOR U5832 ( .A(n3971), .B(n3970), .Z(n3972) );
  XNOR U5833 ( .A(n3973), .B(n3972), .Z(out[76]) );
  XNOR U5834 ( .A(in[745]), .B(n3974), .Z(n4349) );
  NAND U5835 ( .A(n4192), .B(n3975), .Z(n3976) );
  XNOR U5836 ( .A(n4349), .B(n3976), .Z(out[770]) );
  XNOR U5837 ( .A(in[746]), .B(n3977), .Z(n4353) );
  NAND U5838 ( .A(n4194), .B(n3978), .Z(n3979) );
  XNOR U5839 ( .A(n4353), .B(n3979), .Z(out[771]) );
  XNOR U5840 ( .A(in[747]), .B(n3980), .Z(n4365) );
  NAND U5841 ( .A(n4196), .B(n3981), .Z(n3982) );
  XNOR U5842 ( .A(n4365), .B(n3982), .Z(out[772]) );
  XNOR U5843 ( .A(in[748]), .B(n3983), .Z(n4369) );
  NAND U5844 ( .A(n4198), .B(n3984), .Z(n3985) );
  XNOR U5845 ( .A(n4369), .B(n3985), .Z(out[773]) );
  XNOR U5846 ( .A(in[749]), .B(n3986), .Z(n4373) );
  NAND U5847 ( .A(n4200), .B(n3987), .Z(n3988) );
  XNOR U5848 ( .A(n4373), .B(n3988), .Z(out[774]) );
  XNOR U5849 ( .A(in[750]), .B(n3989), .Z(n4377) );
  NAND U5850 ( .A(n4202), .B(n3990), .Z(n3991) );
  XNOR U5851 ( .A(n4377), .B(n3991), .Z(out[775]) );
  XNOR U5852 ( .A(in[751]), .B(n3992), .Z(n4381) );
  NAND U5853 ( .A(n4208), .B(n3993), .Z(n3994) );
  XNOR U5854 ( .A(n4381), .B(n3994), .Z(out[776]) );
  XNOR U5855 ( .A(in[752]), .B(n3995), .Z(n4385) );
  NAND U5856 ( .A(n4210), .B(n3996), .Z(n3997) );
  XNOR U5857 ( .A(n4385), .B(n3997), .Z(out[777]) );
  XNOR U5858 ( .A(in[753]), .B(n3998), .Z(n4389) );
  NAND U5859 ( .A(n4212), .B(n3999), .Z(n4000) );
  XNOR U5860 ( .A(n4389), .B(n4000), .Z(out[778]) );
  XNOR U5861 ( .A(in[754]), .B(n4001), .Z(n4393) );
  NAND U5862 ( .A(n4214), .B(n4002), .Z(n4003) );
  XNOR U5863 ( .A(n4393), .B(n4003), .Z(out[779]) );
  NOR U5864 ( .A(n4005), .B(n4004), .Z(n4006) );
  XNOR U5865 ( .A(n4007), .B(n4006), .Z(out[77]) );
  XNOR U5866 ( .A(in[755]), .B(n4008), .Z(n4397) );
  NAND U5867 ( .A(n4216), .B(n4009), .Z(n4010) );
  XNOR U5868 ( .A(n4397), .B(n4010), .Z(out[780]) );
  XNOR U5869 ( .A(in[756]), .B(n4011), .Z(n4401) );
  NAND U5870 ( .A(n4218), .B(n4012), .Z(n4013) );
  XNOR U5871 ( .A(n4401), .B(n4013), .Z(out[781]) );
  XNOR U5872 ( .A(in[757]), .B(n4014), .Z(n4409) );
  NAND U5873 ( .A(n4220), .B(n4015), .Z(n4016) );
  XNOR U5874 ( .A(n4409), .B(n4016), .Z(out[782]) );
  XNOR U5875 ( .A(in[758]), .B(n4017), .Z(n4413) );
  NAND U5876 ( .A(n4222), .B(n4018), .Z(n4019) );
  XNOR U5877 ( .A(n4413), .B(n4019), .Z(out[783]) );
  XNOR U5878 ( .A(in[759]), .B(n4020), .Z(n4417) );
  NAND U5879 ( .A(n4224), .B(n4021), .Z(n4022) );
  XNOR U5880 ( .A(n4417), .B(n4022), .Z(out[784]) );
  XNOR U5881 ( .A(in[760]), .B(n4023), .Z(n4421) );
  NAND U5882 ( .A(n4226), .B(n4024), .Z(n4025) );
  XNOR U5883 ( .A(n4421), .B(n4025), .Z(out[785]) );
  XNOR U5884 ( .A(in[761]), .B(n4026), .Z(n4425) );
  NAND U5885 ( .A(n4232), .B(n4027), .Z(n4028) );
  XNOR U5886 ( .A(n4425), .B(n4028), .Z(out[786]) );
  XNOR U5887 ( .A(in[762]), .B(n4029), .Z(n4429) );
  NAND U5888 ( .A(n4234), .B(n4030), .Z(n4031) );
  XNOR U5889 ( .A(n4429), .B(n4031), .Z(out[787]) );
  XNOR U5890 ( .A(in[763]), .B(n4032), .Z(n4433) );
  NAND U5891 ( .A(n4236), .B(n4033), .Z(n4034) );
  XNOR U5892 ( .A(n4433), .B(n4034), .Z(out[788]) );
  XNOR U5893 ( .A(in[764]), .B(n4035), .Z(n4437) );
  NAND U5894 ( .A(n4238), .B(n4036), .Z(n4037) );
  XNOR U5895 ( .A(n4437), .B(n4037), .Z(out[789]) );
  NOR U5896 ( .A(n4039), .B(n4038), .Z(n4040) );
  XNOR U5897 ( .A(n4041), .B(n4040), .Z(out[78]) );
  XNOR U5898 ( .A(in[765]), .B(n4042), .Z(n4441) );
  NAND U5899 ( .A(n4240), .B(n4043), .Z(n4044) );
  XNOR U5900 ( .A(n4441), .B(n4044), .Z(out[790]) );
  XNOR U5901 ( .A(in[766]), .B(n4045), .Z(n4445) );
  NAND U5902 ( .A(n4242), .B(n4046), .Z(n4047) );
  XNOR U5903 ( .A(n4445), .B(n4047), .Z(out[791]) );
  XNOR U5904 ( .A(in[767]), .B(n4048), .Z(n4453) );
  NAND U5905 ( .A(n4244), .B(n4049), .Z(n4050) );
  XNOR U5906 ( .A(n4453), .B(n4050), .Z(out[792]) );
  XNOR U5907 ( .A(in[704]), .B(n4051), .Z(n4457) );
  NAND U5908 ( .A(n4246), .B(n4052), .Z(n4053) );
  XNOR U5909 ( .A(n4457), .B(n4053), .Z(out[793]) );
  XNOR U5910 ( .A(in[705]), .B(n4054), .Z(n4461) );
  NAND U5911 ( .A(n4248), .B(n4055), .Z(n4056) );
  XNOR U5912 ( .A(n4461), .B(n4056), .Z(out[794]) );
  XNOR U5913 ( .A(in[706]), .B(n4057), .Z(n4465) );
  NAND U5914 ( .A(n4250), .B(n4058), .Z(n4059) );
  XNOR U5915 ( .A(n4465), .B(n4059), .Z(out[795]) );
  XNOR U5916 ( .A(in[707]), .B(n4060), .Z(n4469) );
  NAND U5917 ( .A(n4256), .B(n4061), .Z(n4062) );
  XNOR U5918 ( .A(n4469), .B(n4062), .Z(out[796]) );
  XNOR U5919 ( .A(in[708]), .B(n4063), .Z(n4473) );
  NAND U5920 ( .A(n4258), .B(n4064), .Z(n4065) );
  XNOR U5921 ( .A(n4473), .B(n4065), .Z(out[797]) );
  XNOR U5922 ( .A(in[709]), .B(n4066), .Z(n4477) );
  NAND U5923 ( .A(n4260), .B(n4067), .Z(n4068) );
  XNOR U5924 ( .A(n4477), .B(n4068), .Z(out[798]) );
  XNOR U5925 ( .A(in[710]), .B(n4069), .Z(n4481) );
  NAND U5926 ( .A(n4262), .B(n4070), .Z(n4071) );
  XNOR U5927 ( .A(n4481), .B(n4071), .Z(out[799]) );
  NOR U5928 ( .A(n4073), .B(n4072), .Z(n4074) );
  XNOR U5929 ( .A(n4075), .B(n4074), .Z(out[79]) );
  OR U5930 ( .A(n4077), .B(n4076), .Z(n4078) );
  XNOR U5931 ( .A(n4079), .B(n4078), .Z(out[7]) );
  XNOR U5932 ( .A(in[711]), .B(n4080), .Z(n4485) );
  NAND U5933 ( .A(n4264), .B(n4081), .Z(n4082) );
  XNOR U5934 ( .A(n4485), .B(n4082), .Z(out[800]) );
  XNOR U5935 ( .A(in[712]), .B(n4083), .Z(n4489) );
  NAND U5936 ( .A(n4266), .B(n4084), .Z(n4085) );
  XNOR U5937 ( .A(n4489), .B(n4085), .Z(out[801]) );
  XNOR U5938 ( .A(in[713]), .B(n4086), .Z(n4497) );
  NAND U5939 ( .A(n4268), .B(n4087), .Z(n4088) );
  XNOR U5940 ( .A(n4497), .B(n4088), .Z(out[802]) );
  XNOR U5941 ( .A(in[714]), .B(n4089), .Z(n4501) );
  NAND U5942 ( .A(n4270), .B(n4090), .Z(n4091) );
  XNOR U5943 ( .A(n4501), .B(n4091), .Z(out[803]) );
  XNOR U5944 ( .A(in[715]), .B(n4092), .Z(n4505) );
  NAND U5945 ( .A(n4272), .B(n4093), .Z(n4094) );
  XNOR U5946 ( .A(n4505), .B(n4094), .Z(out[804]) );
  XOR U5947 ( .A(n4095), .B(in[716]), .Z(n4509) );
  NAND U5948 ( .A(n4274), .B(n4096), .Z(n4097) );
  XNOR U5949 ( .A(n4509), .B(n4097), .Z(out[805]) );
  XOR U5950 ( .A(n4098), .B(in[717]), .Z(n4513) );
  NAND U5951 ( .A(n4280), .B(n4099), .Z(n4100) );
  XNOR U5952 ( .A(n4513), .B(n4100), .Z(out[806]) );
  XOR U5953 ( .A(n4101), .B(in[718]), .Z(n4517) );
  NAND U5954 ( .A(n4282), .B(n4102), .Z(n4103) );
  XNOR U5955 ( .A(n4517), .B(n4103), .Z(out[807]) );
  XOR U5956 ( .A(n4104), .B(in[719]), .Z(n4521) );
  NAND U5957 ( .A(n4284), .B(n4105), .Z(n4106) );
  XNOR U5958 ( .A(n4521), .B(n4106), .Z(out[808]) );
  XOR U5959 ( .A(n4107), .B(in[720]), .Z(n4525) );
  NAND U5960 ( .A(n4286), .B(n4108), .Z(n4109) );
  XNOR U5961 ( .A(n4525), .B(n4109), .Z(out[809]) );
  NOR U5962 ( .A(n4111), .B(n4110), .Z(n4112) );
  XNOR U5963 ( .A(n4113), .B(n4112), .Z(out[80]) );
  XOR U5964 ( .A(n4114), .B(in[721]), .Z(n4529) );
  NAND U5965 ( .A(n4288), .B(n4115), .Z(n4116) );
  XNOR U5966 ( .A(n4529), .B(n4116), .Z(out[810]) );
  XOR U5967 ( .A(n4117), .B(in[722]), .Z(n4533) );
  NAND U5968 ( .A(n4290), .B(n4118), .Z(n4119) );
  XNOR U5969 ( .A(n4533), .B(n4119), .Z(out[811]) );
  XOR U5970 ( .A(n4120), .B(in[723]), .Z(n4541) );
  NAND U5971 ( .A(n4292), .B(n4121), .Z(n4122) );
  XNOR U5972 ( .A(n4541), .B(n4122), .Z(out[812]) );
  XOR U5973 ( .A(in[724]), .B(n4123), .Z(n4545) );
  NAND U5974 ( .A(n4294), .B(n4124), .Z(n4125) );
  XNOR U5975 ( .A(n4545), .B(n4125), .Z(out[813]) );
  XOR U5976 ( .A(in[725]), .B(n4126), .Z(n4549) );
  NAND U5977 ( .A(n4296), .B(n4127), .Z(n4128) );
  XNOR U5978 ( .A(n4549), .B(n4128), .Z(out[814]) );
  XOR U5979 ( .A(in[726]), .B(n4129), .Z(n4553) );
  NAND U5980 ( .A(n4298), .B(n4130), .Z(n4131) );
  XNOR U5981 ( .A(n4553), .B(n4131), .Z(out[815]) );
  XOR U5982 ( .A(in[727]), .B(n4132), .Z(n4557) );
  NAND U5983 ( .A(n4304), .B(n4133), .Z(n4134) );
  XNOR U5984 ( .A(n4557), .B(n4134), .Z(out[816]) );
  XOR U5985 ( .A(in[728]), .B(n4135), .Z(n4561) );
  NAND U5986 ( .A(n4306), .B(n4136), .Z(n4137) );
  XNOR U5987 ( .A(n4561), .B(n4137), .Z(out[817]) );
  XOR U5988 ( .A(in[729]), .B(n4138), .Z(n4565) );
  NAND U5989 ( .A(n4308), .B(n4139), .Z(n4140) );
  XNOR U5990 ( .A(n4565), .B(n4140), .Z(out[818]) );
  XOR U5991 ( .A(in[730]), .B(n4141), .Z(n4569) );
  NAND U5992 ( .A(n4310), .B(n4142), .Z(n4143) );
  XNOR U5993 ( .A(n4569), .B(n4143), .Z(out[819]) );
  NOR U5994 ( .A(n4145), .B(n4144), .Z(n4146) );
  XNOR U5995 ( .A(n4147), .B(n4146), .Z(out[81]) );
  XOR U5996 ( .A(in[731]), .B(n4148), .Z(n4573) );
  NAND U5997 ( .A(n4312), .B(n4149), .Z(n4150) );
  XNOR U5998 ( .A(n4573), .B(n4150), .Z(out[820]) );
  XOR U5999 ( .A(in[732]), .B(n4151), .Z(n4577) );
  NAND U6000 ( .A(n4314), .B(n4152), .Z(n4153) );
  XNOR U6001 ( .A(n4577), .B(n4153), .Z(out[821]) );
  XOR U6002 ( .A(in[733]), .B(n4154), .Z(n4585) );
  NAND U6003 ( .A(n4316), .B(n4155), .Z(n4156) );
  XNOR U6004 ( .A(n4585), .B(n4156), .Z(out[822]) );
  XOR U6005 ( .A(in[734]), .B(n4157), .Z(n4589) );
  NAND U6006 ( .A(n4318), .B(n4158), .Z(n4159) );
  XNOR U6007 ( .A(n4589), .B(n4159), .Z(out[823]) );
  XOR U6008 ( .A(in[735]), .B(n4160), .Z(n4593) );
  NAND U6009 ( .A(n4320), .B(n4161), .Z(n4162) );
  XNOR U6010 ( .A(n4593), .B(n4162), .Z(out[824]) );
  XOR U6011 ( .A(in[736]), .B(n4163), .Z(n4597) );
  NAND U6012 ( .A(n4322), .B(n4164), .Z(n4165) );
  XNOR U6013 ( .A(n4597), .B(n4165), .Z(out[825]) );
  XOR U6014 ( .A(in[737]), .B(n4166), .Z(n4601) );
  NAND U6015 ( .A(n4328), .B(n4167), .Z(n4168) );
  XNOR U6016 ( .A(n4601), .B(n4168), .Z(out[826]) );
  XOR U6017 ( .A(in[738]), .B(n4169), .Z(n4605) );
  NAND U6018 ( .A(n4330), .B(n4170), .Z(n4171) );
  XNOR U6019 ( .A(n4605), .B(n4171), .Z(out[827]) );
  XOR U6020 ( .A(in[739]), .B(n4172), .Z(n4609) );
  NAND U6021 ( .A(n4332), .B(n4173), .Z(n4174) );
  XNOR U6022 ( .A(n4609), .B(n4174), .Z(out[828]) );
  XNOR U6023 ( .A(in[740]), .B(n4175), .Z(n4613) );
  NAND U6024 ( .A(n4334), .B(n4176), .Z(n4177) );
  XNOR U6025 ( .A(n4613), .B(n4177), .Z(out[829]) );
  NOR U6026 ( .A(n4179), .B(n4178), .Z(n4180) );
  XNOR U6027 ( .A(n4181), .B(n4180), .Z(out[82]) );
  XNOR U6028 ( .A(in[741]), .B(n4182), .Z(n4617) );
  NAND U6029 ( .A(n4336), .B(n4183), .Z(n4184) );
  XNOR U6030 ( .A(n4617), .B(n4184), .Z(out[830]) );
  XNOR U6031 ( .A(in[742]), .B(n4185), .Z(n4621) );
  NAND U6032 ( .A(n4338), .B(n4186), .Z(n4187) );
  XNOR U6033 ( .A(n4621), .B(n4187), .Z(out[831]) );
  OR U6034 ( .A(n4341), .B(n4188), .Z(n4189) );
  XNOR U6035 ( .A(n4340), .B(n4189), .Z(out[832]) );
  OR U6036 ( .A(n4345), .B(n4190), .Z(n4191) );
  XNOR U6037 ( .A(n4344), .B(n4191), .Z(out[833]) );
  OR U6038 ( .A(n4349), .B(n4192), .Z(n4193) );
  XNOR U6039 ( .A(n4348), .B(n4193), .Z(out[834]) );
  OR U6040 ( .A(n4353), .B(n4194), .Z(n4195) );
  XNOR U6041 ( .A(n4352), .B(n4195), .Z(out[835]) );
  OR U6042 ( .A(n4365), .B(n4196), .Z(n4197) );
  XNOR U6043 ( .A(n4364), .B(n4197), .Z(out[836]) );
  OR U6044 ( .A(n4369), .B(n4198), .Z(n4199) );
  XNOR U6045 ( .A(n4368), .B(n4199), .Z(out[837]) );
  OR U6046 ( .A(n4373), .B(n4200), .Z(n4201) );
  XNOR U6047 ( .A(n4372), .B(n4201), .Z(out[838]) );
  OR U6048 ( .A(n4377), .B(n4202), .Z(n4203) );
  XNOR U6049 ( .A(n4376), .B(n4203), .Z(out[839]) );
  NOR U6050 ( .A(n4205), .B(n4204), .Z(n4206) );
  XNOR U6051 ( .A(n4207), .B(n4206), .Z(out[83]) );
  OR U6052 ( .A(n4381), .B(n4208), .Z(n4209) );
  XNOR U6053 ( .A(n4380), .B(n4209), .Z(out[840]) );
  OR U6054 ( .A(n4385), .B(n4210), .Z(n4211) );
  XNOR U6055 ( .A(n4384), .B(n4211), .Z(out[841]) );
  OR U6056 ( .A(n4389), .B(n4212), .Z(n4213) );
  XNOR U6057 ( .A(n4388), .B(n4213), .Z(out[842]) );
  OR U6058 ( .A(n4393), .B(n4214), .Z(n4215) );
  XNOR U6059 ( .A(n4392), .B(n4215), .Z(out[843]) );
  OR U6060 ( .A(n4397), .B(n4216), .Z(n4217) );
  XNOR U6061 ( .A(n4396), .B(n4217), .Z(out[844]) );
  OR U6062 ( .A(n4401), .B(n4218), .Z(n4219) );
  XNOR U6063 ( .A(n4400), .B(n4219), .Z(out[845]) );
  OR U6064 ( .A(n4409), .B(n4220), .Z(n4221) );
  XNOR U6065 ( .A(n4408), .B(n4221), .Z(out[846]) );
  OR U6066 ( .A(n4413), .B(n4222), .Z(n4223) );
  XNOR U6067 ( .A(n4412), .B(n4223), .Z(out[847]) );
  OR U6068 ( .A(n4417), .B(n4224), .Z(n4225) );
  XNOR U6069 ( .A(n4416), .B(n4225), .Z(out[848]) );
  OR U6070 ( .A(n4421), .B(n4226), .Z(n4227) );
  XNOR U6071 ( .A(n4420), .B(n4227), .Z(out[849]) );
  NOR U6072 ( .A(n4229), .B(n4228), .Z(n4230) );
  XNOR U6073 ( .A(n4231), .B(n4230), .Z(out[84]) );
  OR U6074 ( .A(n4425), .B(n4232), .Z(n4233) );
  XNOR U6075 ( .A(n4424), .B(n4233), .Z(out[850]) );
  OR U6076 ( .A(n4429), .B(n4234), .Z(n4235) );
  XNOR U6077 ( .A(n4428), .B(n4235), .Z(out[851]) );
  OR U6078 ( .A(n4433), .B(n4236), .Z(n4237) );
  XNOR U6079 ( .A(n4432), .B(n4237), .Z(out[852]) );
  OR U6080 ( .A(n4437), .B(n4238), .Z(n4239) );
  XNOR U6081 ( .A(n4436), .B(n4239), .Z(out[853]) );
  OR U6082 ( .A(n4441), .B(n4240), .Z(n4241) );
  XNOR U6083 ( .A(n4440), .B(n4241), .Z(out[854]) );
  OR U6084 ( .A(n4445), .B(n4242), .Z(n4243) );
  XNOR U6085 ( .A(n4444), .B(n4243), .Z(out[855]) );
  OR U6086 ( .A(n4453), .B(n4244), .Z(n4245) );
  XNOR U6087 ( .A(n4452), .B(n4245), .Z(out[856]) );
  OR U6088 ( .A(n4457), .B(n4246), .Z(n4247) );
  XNOR U6089 ( .A(n4456), .B(n4247), .Z(out[857]) );
  OR U6090 ( .A(n4461), .B(n4248), .Z(n4249) );
  XNOR U6091 ( .A(n4460), .B(n4249), .Z(out[858]) );
  OR U6092 ( .A(n4465), .B(n4250), .Z(n4251) );
  XNOR U6093 ( .A(n4464), .B(n4251), .Z(out[859]) );
  NOR U6094 ( .A(n4253), .B(n4252), .Z(n4254) );
  XNOR U6095 ( .A(n4255), .B(n4254), .Z(out[85]) );
  OR U6096 ( .A(n4469), .B(n4256), .Z(n4257) );
  XNOR U6097 ( .A(n4468), .B(n4257), .Z(out[860]) );
  OR U6098 ( .A(n4473), .B(n4258), .Z(n4259) );
  XNOR U6099 ( .A(n4472), .B(n4259), .Z(out[861]) );
  OR U6100 ( .A(n4477), .B(n4260), .Z(n4261) );
  XNOR U6101 ( .A(n4476), .B(n4261), .Z(out[862]) );
  OR U6102 ( .A(n4481), .B(n4262), .Z(n4263) );
  XNOR U6103 ( .A(n4480), .B(n4263), .Z(out[863]) );
  OR U6104 ( .A(n4485), .B(n4264), .Z(n4265) );
  XNOR U6105 ( .A(n4484), .B(n4265), .Z(out[864]) );
  OR U6106 ( .A(n4489), .B(n4266), .Z(n4267) );
  XNOR U6107 ( .A(n4488), .B(n4267), .Z(out[865]) );
  OR U6108 ( .A(n4497), .B(n4268), .Z(n4269) );
  XNOR U6109 ( .A(n4496), .B(n4269), .Z(out[866]) );
  OR U6110 ( .A(n4501), .B(n4270), .Z(n4271) );
  XNOR U6111 ( .A(n4500), .B(n4271), .Z(out[867]) );
  OR U6112 ( .A(n4505), .B(n4272), .Z(n4273) );
  XNOR U6113 ( .A(n4504), .B(n4273), .Z(out[868]) );
  OR U6114 ( .A(n4509), .B(n4274), .Z(n4275) );
  XNOR U6115 ( .A(n4508), .B(n4275), .Z(out[869]) );
  NOR U6116 ( .A(n4277), .B(n4276), .Z(n4278) );
  XNOR U6117 ( .A(n4279), .B(n4278), .Z(out[86]) );
  OR U6118 ( .A(n4513), .B(n4280), .Z(n4281) );
  XNOR U6119 ( .A(n4512), .B(n4281), .Z(out[870]) );
  OR U6120 ( .A(n4517), .B(n4282), .Z(n4283) );
  XNOR U6121 ( .A(n4516), .B(n4283), .Z(out[871]) );
  OR U6122 ( .A(n4521), .B(n4284), .Z(n4285) );
  XNOR U6123 ( .A(n4520), .B(n4285), .Z(out[872]) );
  OR U6124 ( .A(n4525), .B(n4286), .Z(n4287) );
  XNOR U6125 ( .A(n4524), .B(n4287), .Z(out[873]) );
  OR U6126 ( .A(n4529), .B(n4288), .Z(n4289) );
  XNOR U6127 ( .A(n4528), .B(n4289), .Z(out[874]) );
  OR U6128 ( .A(n4533), .B(n4290), .Z(n4291) );
  XNOR U6129 ( .A(n4532), .B(n4291), .Z(out[875]) );
  OR U6130 ( .A(n4541), .B(n4292), .Z(n4293) );
  XNOR U6131 ( .A(n4540), .B(n4293), .Z(out[876]) );
  OR U6132 ( .A(n4545), .B(n4294), .Z(n4295) );
  XNOR U6133 ( .A(n4544), .B(n4295), .Z(out[877]) );
  OR U6134 ( .A(n4549), .B(n4296), .Z(n4297) );
  XNOR U6135 ( .A(n4548), .B(n4297), .Z(out[878]) );
  OR U6136 ( .A(n4553), .B(n4298), .Z(n4299) );
  XNOR U6137 ( .A(n4552), .B(n4299), .Z(out[879]) );
  NOR U6138 ( .A(n4301), .B(n4300), .Z(n4302) );
  XNOR U6139 ( .A(n4303), .B(n4302), .Z(out[87]) );
  OR U6140 ( .A(n4557), .B(n4304), .Z(n4305) );
  XNOR U6141 ( .A(n4556), .B(n4305), .Z(out[880]) );
  OR U6142 ( .A(n4561), .B(n4306), .Z(n4307) );
  XNOR U6143 ( .A(n4560), .B(n4307), .Z(out[881]) );
  OR U6144 ( .A(n4565), .B(n4308), .Z(n4309) );
  XNOR U6145 ( .A(n4564), .B(n4309), .Z(out[882]) );
  OR U6146 ( .A(n4569), .B(n4310), .Z(n4311) );
  XNOR U6147 ( .A(n4568), .B(n4311), .Z(out[883]) );
  OR U6148 ( .A(n4573), .B(n4312), .Z(n4313) );
  XNOR U6149 ( .A(n4572), .B(n4313), .Z(out[884]) );
  OR U6150 ( .A(n4577), .B(n4314), .Z(n4315) );
  XNOR U6151 ( .A(n4576), .B(n4315), .Z(out[885]) );
  OR U6152 ( .A(n4585), .B(n4316), .Z(n4317) );
  XNOR U6153 ( .A(n4584), .B(n4317), .Z(out[886]) );
  OR U6154 ( .A(n4589), .B(n4318), .Z(n4319) );
  XNOR U6155 ( .A(n4588), .B(n4319), .Z(out[887]) );
  OR U6156 ( .A(n4593), .B(n4320), .Z(n4321) );
  XNOR U6157 ( .A(n4592), .B(n4321), .Z(out[888]) );
  OR U6158 ( .A(n4597), .B(n4322), .Z(n4323) );
  XNOR U6159 ( .A(n4596), .B(n4323), .Z(out[889]) );
  NOR U6160 ( .A(n4325), .B(n4324), .Z(n4326) );
  XNOR U6161 ( .A(n4327), .B(n4326), .Z(out[88]) );
  OR U6162 ( .A(n4601), .B(n4328), .Z(n4329) );
  XNOR U6163 ( .A(n4600), .B(n4329), .Z(out[890]) );
  OR U6164 ( .A(n4605), .B(n4330), .Z(n4331) );
  XNOR U6165 ( .A(n4604), .B(n4331), .Z(out[891]) );
  OR U6166 ( .A(n4609), .B(n4332), .Z(n4333) );
  XNOR U6167 ( .A(n4608), .B(n4333), .Z(out[892]) );
  OR U6168 ( .A(n4613), .B(n4334), .Z(n4335) );
  XNOR U6169 ( .A(n4612), .B(n4335), .Z(out[893]) );
  OR U6170 ( .A(n4617), .B(n4336), .Z(n4337) );
  XNOR U6171 ( .A(n4616), .B(n4337), .Z(out[894]) );
  OR U6172 ( .A(n4621), .B(n4338), .Z(n4339) );
  XNOR U6173 ( .A(n4620), .B(n4339), .Z(out[895]) );
  ANDN U6174 ( .B(n4341), .A(n4340), .Z(n4342) );
  XNOR U6175 ( .A(n4343), .B(n4342), .Z(out[896]) );
  ANDN U6176 ( .B(n4345), .A(n4344), .Z(n4346) );
  XNOR U6177 ( .A(n4347), .B(n4346), .Z(out[897]) );
  ANDN U6178 ( .B(n4349), .A(n4348), .Z(n4350) );
  XNOR U6179 ( .A(n4351), .B(n4350), .Z(out[898]) );
  ANDN U6180 ( .B(n4353), .A(n4352), .Z(n4354) );
  XNOR U6181 ( .A(n4355), .B(n4354), .Z(out[899]) );
  NOR U6182 ( .A(n4357), .B(n4356), .Z(n4358) );
  XNOR U6183 ( .A(n4359), .B(n4358), .Z(out[89]) );
  OR U6184 ( .A(n4361), .B(n4360), .Z(n4362) );
  XNOR U6185 ( .A(n4363), .B(n4362), .Z(out[8]) );
  ANDN U6186 ( .B(n4365), .A(n4364), .Z(n4366) );
  XNOR U6187 ( .A(n4367), .B(n4366), .Z(out[900]) );
  ANDN U6188 ( .B(n4369), .A(n4368), .Z(n4370) );
  XNOR U6189 ( .A(n4371), .B(n4370), .Z(out[901]) );
  ANDN U6190 ( .B(n4373), .A(n4372), .Z(n4374) );
  XNOR U6191 ( .A(n4375), .B(n4374), .Z(out[902]) );
  ANDN U6192 ( .B(n4377), .A(n4376), .Z(n4378) );
  XNOR U6193 ( .A(n4379), .B(n4378), .Z(out[903]) );
  ANDN U6194 ( .B(n4381), .A(n4380), .Z(n4382) );
  XNOR U6195 ( .A(n4383), .B(n4382), .Z(out[904]) );
  ANDN U6196 ( .B(n4385), .A(n4384), .Z(n4386) );
  XNOR U6197 ( .A(n4387), .B(n4386), .Z(out[905]) );
  ANDN U6198 ( .B(n4389), .A(n4388), .Z(n4390) );
  XNOR U6199 ( .A(n4391), .B(n4390), .Z(out[906]) );
  ANDN U6200 ( .B(n4393), .A(n4392), .Z(n4394) );
  XNOR U6201 ( .A(n4395), .B(n4394), .Z(out[907]) );
  ANDN U6202 ( .B(n4397), .A(n4396), .Z(n4398) );
  XNOR U6203 ( .A(n4399), .B(n4398), .Z(out[908]) );
  ANDN U6204 ( .B(n4401), .A(n4400), .Z(n4402) );
  XNOR U6205 ( .A(n4403), .B(n4402), .Z(out[909]) );
  NOR U6206 ( .A(n4405), .B(n4404), .Z(n4406) );
  XNOR U6207 ( .A(n4407), .B(n4406), .Z(out[90]) );
  ANDN U6208 ( .B(n4409), .A(n4408), .Z(n4410) );
  XNOR U6209 ( .A(n4411), .B(n4410), .Z(out[910]) );
  ANDN U6210 ( .B(n4413), .A(n4412), .Z(n4414) );
  XNOR U6211 ( .A(n4415), .B(n4414), .Z(out[911]) );
  ANDN U6212 ( .B(n4417), .A(n4416), .Z(n4418) );
  XNOR U6213 ( .A(n4419), .B(n4418), .Z(out[912]) );
  ANDN U6214 ( .B(n4421), .A(n4420), .Z(n4422) );
  XNOR U6215 ( .A(n4423), .B(n4422), .Z(out[913]) );
  ANDN U6216 ( .B(n4425), .A(n4424), .Z(n4426) );
  XNOR U6217 ( .A(n4427), .B(n4426), .Z(out[914]) );
  ANDN U6218 ( .B(n4429), .A(n4428), .Z(n4430) );
  XNOR U6219 ( .A(n4431), .B(n4430), .Z(out[915]) );
  ANDN U6220 ( .B(n4433), .A(n4432), .Z(n4434) );
  XNOR U6221 ( .A(n4435), .B(n4434), .Z(out[916]) );
  ANDN U6222 ( .B(n4437), .A(n4436), .Z(n4438) );
  XNOR U6223 ( .A(n4439), .B(n4438), .Z(out[917]) );
  ANDN U6224 ( .B(n4441), .A(n4440), .Z(n4442) );
  XNOR U6225 ( .A(n4443), .B(n4442), .Z(out[918]) );
  ANDN U6226 ( .B(n4445), .A(n4444), .Z(n4446) );
  XNOR U6227 ( .A(n4447), .B(n4446), .Z(out[919]) );
  NOR U6228 ( .A(n4449), .B(n4448), .Z(n4450) );
  XNOR U6229 ( .A(n4451), .B(n4450), .Z(out[91]) );
  ANDN U6230 ( .B(n4453), .A(n4452), .Z(n4454) );
  XNOR U6231 ( .A(n4455), .B(n4454), .Z(out[920]) );
  ANDN U6232 ( .B(n4457), .A(n4456), .Z(n4458) );
  XNOR U6233 ( .A(n4459), .B(n4458), .Z(out[921]) );
  ANDN U6234 ( .B(n4461), .A(n4460), .Z(n4462) );
  XNOR U6235 ( .A(n4463), .B(n4462), .Z(out[922]) );
  ANDN U6236 ( .B(n4465), .A(n4464), .Z(n4466) );
  XNOR U6237 ( .A(n4467), .B(n4466), .Z(out[923]) );
  ANDN U6238 ( .B(n4469), .A(n4468), .Z(n4470) );
  XNOR U6239 ( .A(n4471), .B(n4470), .Z(out[924]) );
  ANDN U6240 ( .B(n4473), .A(n4472), .Z(n4474) );
  XNOR U6241 ( .A(n4475), .B(n4474), .Z(out[925]) );
  ANDN U6242 ( .B(n4477), .A(n4476), .Z(n4478) );
  XNOR U6243 ( .A(n4479), .B(n4478), .Z(out[926]) );
  ANDN U6244 ( .B(n4481), .A(n4480), .Z(n4482) );
  XNOR U6245 ( .A(n4483), .B(n4482), .Z(out[927]) );
  ANDN U6246 ( .B(n4485), .A(n4484), .Z(n4486) );
  XNOR U6247 ( .A(n4487), .B(n4486), .Z(out[928]) );
  ANDN U6248 ( .B(n4489), .A(n4488), .Z(n4490) );
  XNOR U6249 ( .A(n4491), .B(n4490), .Z(out[929]) );
  ANDN U6250 ( .B(n4493), .A(n4492), .Z(n4494) );
  XNOR U6251 ( .A(n4495), .B(n4494), .Z(out[92]) );
  ANDN U6252 ( .B(n4497), .A(n4496), .Z(n4498) );
  XNOR U6253 ( .A(n4499), .B(n4498), .Z(out[930]) );
  ANDN U6254 ( .B(n4501), .A(n4500), .Z(n4502) );
  XNOR U6255 ( .A(n4503), .B(n4502), .Z(out[931]) );
  ANDN U6256 ( .B(n4505), .A(n4504), .Z(n4506) );
  XNOR U6257 ( .A(n4507), .B(n4506), .Z(out[932]) );
  ANDN U6258 ( .B(n4509), .A(n4508), .Z(n4510) );
  XNOR U6259 ( .A(n4511), .B(n4510), .Z(out[933]) );
  ANDN U6260 ( .B(n4513), .A(n4512), .Z(n4514) );
  XNOR U6261 ( .A(n4515), .B(n4514), .Z(out[934]) );
  ANDN U6262 ( .B(n4517), .A(n4516), .Z(n4518) );
  XNOR U6263 ( .A(n4519), .B(n4518), .Z(out[935]) );
  ANDN U6264 ( .B(n4521), .A(n4520), .Z(n4522) );
  XNOR U6265 ( .A(n4523), .B(n4522), .Z(out[936]) );
  ANDN U6266 ( .B(n4525), .A(n4524), .Z(n4526) );
  XNOR U6267 ( .A(n4527), .B(n4526), .Z(out[937]) );
  ANDN U6268 ( .B(n4529), .A(n4528), .Z(n4530) );
  XNOR U6269 ( .A(n4531), .B(n4530), .Z(out[938]) );
  ANDN U6270 ( .B(n4533), .A(n4532), .Z(n4534) );
  XNOR U6271 ( .A(n4535), .B(n4534), .Z(out[939]) );
  ANDN U6272 ( .B(n4537), .A(n4536), .Z(n4538) );
  XNOR U6273 ( .A(n4539), .B(n4538), .Z(out[93]) );
  ANDN U6274 ( .B(n4541), .A(n4540), .Z(n4542) );
  XNOR U6275 ( .A(n4543), .B(n4542), .Z(out[940]) );
  ANDN U6276 ( .B(n4545), .A(n4544), .Z(n4546) );
  XNOR U6277 ( .A(n4547), .B(n4546), .Z(out[941]) );
  ANDN U6278 ( .B(n4549), .A(n4548), .Z(n4550) );
  XNOR U6279 ( .A(n4551), .B(n4550), .Z(out[942]) );
  ANDN U6280 ( .B(n4553), .A(n4552), .Z(n4554) );
  XNOR U6281 ( .A(n4555), .B(n4554), .Z(out[943]) );
  ANDN U6282 ( .B(n4557), .A(n4556), .Z(n4558) );
  XNOR U6283 ( .A(n4559), .B(n4558), .Z(out[944]) );
  ANDN U6284 ( .B(n4561), .A(n4560), .Z(n4562) );
  XNOR U6285 ( .A(n4563), .B(n4562), .Z(out[945]) );
  ANDN U6286 ( .B(n4565), .A(n4564), .Z(n4566) );
  XNOR U6287 ( .A(n4567), .B(n4566), .Z(out[946]) );
  ANDN U6288 ( .B(n4569), .A(n4568), .Z(n4570) );
  XNOR U6289 ( .A(n4571), .B(n4570), .Z(out[947]) );
  ANDN U6290 ( .B(n4573), .A(n4572), .Z(n4574) );
  XNOR U6291 ( .A(n4575), .B(n4574), .Z(out[948]) );
  ANDN U6292 ( .B(n4577), .A(n4576), .Z(n4578) );
  XNOR U6293 ( .A(n4579), .B(n4578), .Z(out[949]) );
  ANDN U6294 ( .B(n4581), .A(n4580), .Z(n4582) );
  XNOR U6295 ( .A(n4583), .B(n4582), .Z(out[94]) );
  ANDN U6296 ( .B(n4585), .A(n4584), .Z(n4586) );
  XNOR U6297 ( .A(n4587), .B(n4586), .Z(out[950]) );
  ANDN U6298 ( .B(n4589), .A(n4588), .Z(n4590) );
  XNOR U6299 ( .A(n4591), .B(n4590), .Z(out[951]) );
  ANDN U6300 ( .B(n4593), .A(n4592), .Z(n4594) );
  XNOR U6301 ( .A(n4595), .B(n4594), .Z(out[952]) );
  ANDN U6302 ( .B(n4597), .A(n4596), .Z(n4598) );
  XNOR U6303 ( .A(n4599), .B(n4598), .Z(out[953]) );
  ANDN U6304 ( .B(n4601), .A(n4600), .Z(n4602) );
  XNOR U6305 ( .A(n4603), .B(n4602), .Z(out[954]) );
  ANDN U6306 ( .B(n4605), .A(n4604), .Z(n4606) );
  XNOR U6307 ( .A(n4607), .B(n4606), .Z(out[955]) );
  ANDN U6308 ( .B(n4609), .A(n4608), .Z(n4610) );
  XNOR U6309 ( .A(n4611), .B(n4610), .Z(out[956]) );
  ANDN U6310 ( .B(n4613), .A(n4612), .Z(n4614) );
  XNOR U6311 ( .A(n4615), .B(n4614), .Z(out[957]) );
  ANDN U6312 ( .B(n4617), .A(n4616), .Z(n4618) );
  XNOR U6313 ( .A(n4619), .B(n4618), .Z(out[958]) );
  ANDN U6314 ( .B(n4621), .A(n4620), .Z(n4622) );
  XNOR U6315 ( .A(n4623), .B(n4622), .Z(out[959]) );
  ANDN U6316 ( .B(n4625), .A(n4624), .Z(n4626) );
  XNOR U6317 ( .A(n4627), .B(n4626), .Z(out[95]) );
  ANDN U6318 ( .B(n4629), .A(n4628), .Z(n4630) );
  XNOR U6319 ( .A(n4631), .B(n4630), .Z(out[960]) );
  ANDN U6320 ( .B(n4633), .A(n4632), .Z(n4634) );
  XNOR U6321 ( .A(n4635), .B(n4634), .Z(out[961]) );
  ANDN U6322 ( .B(n4637), .A(n4636), .Z(n4638) );
  XNOR U6323 ( .A(n4639), .B(n4638), .Z(out[962]) );
  ANDN U6324 ( .B(n4641), .A(n4640), .Z(n4642) );
  XNOR U6325 ( .A(n4643), .B(n4642), .Z(out[963]) );
  ANDN U6326 ( .B(n4645), .A(n4644), .Z(n4646) );
  XNOR U6327 ( .A(n4647), .B(n4646), .Z(out[964]) );
  ANDN U6328 ( .B(n4649), .A(n4648), .Z(n4650) );
  XNOR U6329 ( .A(n4651), .B(n4650), .Z(out[965]) );
  ANDN U6330 ( .B(n4653), .A(n4652), .Z(n4654) );
  XNOR U6331 ( .A(n4655), .B(n4654), .Z(out[966]) );
  ANDN U6332 ( .B(n4657), .A(n4656), .Z(n4658) );
  XNOR U6333 ( .A(n4659), .B(n4658), .Z(out[967]) );
  ANDN U6334 ( .B(n4661), .A(n4660), .Z(n4662) );
  XNOR U6335 ( .A(n4663), .B(n4662), .Z(out[968]) );
  ANDN U6336 ( .B(n4665), .A(n4664), .Z(n4666) );
  XNOR U6337 ( .A(n4667), .B(n4666), .Z(out[969]) );
  ANDN U6338 ( .B(n4669), .A(n4668), .Z(n4670) );
  XNOR U6339 ( .A(n4671), .B(n4670), .Z(out[96]) );
  ANDN U6340 ( .B(n4673), .A(n4672), .Z(n4674) );
  XNOR U6341 ( .A(n4675), .B(n4674), .Z(out[970]) );
  ANDN U6342 ( .B(n4677), .A(n4676), .Z(n4678) );
  XNOR U6343 ( .A(n4679), .B(n4678), .Z(out[971]) );
  ANDN U6344 ( .B(n4681), .A(n4680), .Z(n4682) );
  XNOR U6345 ( .A(n4683), .B(n4682), .Z(out[972]) );
  ANDN U6346 ( .B(n4685), .A(n4684), .Z(n4686) );
  XNOR U6347 ( .A(n4687), .B(n4686), .Z(out[973]) );
  ANDN U6348 ( .B(n4689), .A(n4688), .Z(n4690) );
  XNOR U6349 ( .A(n4691), .B(n4690), .Z(out[974]) );
  ANDN U6350 ( .B(n4693), .A(n4692), .Z(n4694) );
  XNOR U6351 ( .A(n4695), .B(n4694), .Z(out[975]) );
  ANDN U6352 ( .B(n4697), .A(n4696), .Z(n4698) );
  XNOR U6353 ( .A(n4699), .B(n4698), .Z(out[976]) );
  ANDN U6354 ( .B(n4701), .A(n4700), .Z(n4702) );
  XNOR U6355 ( .A(n4703), .B(n4702), .Z(out[977]) );
  ANDN U6356 ( .B(n4705), .A(n4704), .Z(n4706) );
  XNOR U6357 ( .A(n4707), .B(n4706), .Z(out[978]) );
  ANDN U6358 ( .B(n4709), .A(n4708), .Z(n4710) );
  XNOR U6359 ( .A(n4711), .B(n4710), .Z(out[979]) );
  ANDN U6360 ( .B(n4713), .A(n4712), .Z(n4714) );
  XNOR U6361 ( .A(n4715), .B(n4714), .Z(out[97]) );
  ANDN U6362 ( .B(n4717), .A(n4716), .Z(n4718) );
  XNOR U6363 ( .A(n4719), .B(n4718), .Z(out[980]) );
  ANDN U6364 ( .B(n4721), .A(n4720), .Z(n4722) );
  XNOR U6365 ( .A(n4723), .B(n4722), .Z(out[981]) );
  ANDN U6366 ( .B(n4725), .A(n4724), .Z(n4726) );
  XNOR U6367 ( .A(n4727), .B(n4726), .Z(out[982]) );
  ANDN U6368 ( .B(n4729), .A(n4728), .Z(n4730) );
  XNOR U6369 ( .A(n4731), .B(n4730), .Z(out[983]) );
  ANDN U6370 ( .B(n4733), .A(n4732), .Z(n4734) );
  XNOR U6371 ( .A(n4735), .B(n4734), .Z(out[984]) );
  ANDN U6372 ( .B(n4737), .A(n4736), .Z(n4738) );
  XNOR U6373 ( .A(n4739), .B(n4738), .Z(out[985]) );
  ANDN U6374 ( .B(n4741), .A(n4740), .Z(n4742) );
  XNOR U6375 ( .A(n4743), .B(n4742), .Z(out[986]) );
  ANDN U6376 ( .B(n4745), .A(n4744), .Z(n4746) );
  XNOR U6377 ( .A(n4747), .B(n4746), .Z(out[987]) );
  ANDN U6378 ( .B(n4749), .A(n4748), .Z(n4750) );
  XNOR U6379 ( .A(n4751), .B(n4750), .Z(out[988]) );
  ANDN U6380 ( .B(n4753), .A(n4752), .Z(n4754) );
  XNOR U6381 ( .A(n4755), .B(n4754), .Z(out[989]) );
  ANDN U6382 ( .B(n4757), .A(n4756), .Z(n4758) );
  XNOR U6383 ( .A(n4759), .B(n4758), .Z(out[98]) );
  ANDN U6384 ( .B(n4761), .A(n4760), .Z(n4762) );
  XNOR U6385 ( .A(n4763), .B(n4762), .Z(out[990]) );
  ANDN U6386 ( .B(n4765), .A(n4764), .Z(n4766) );
  XNOR U6387 ( .A(n4767), .B(n4766), .Z(out[991]) );
  ANDN U6388 ( .B(n4769), .A(n4768), .Z(n4770) );
  XNOR U6389 ( .A(n4771), .B(n4770), .Z(out[992]) );
  ANDN U6390 ( .B(n4773), .A(n4772), .Z(n4774) );
  XNOR U6391 ( .A(n4775), .B(n4774), .Z(out[993]) );
  ANDN U6392 ( .B(n4777), .A(n4776), .Z(n4778) );
  XNOR U6393 ( .A(n4779), .B(n4778), .Z(out[994]) );
  ANDN U6394 ( .B(n4781), .A(n4780), .Z(n4782) );
  XNOR U6395 ( .A(n4783), .B(n4782), .Z(out[995]) );
  ANDN U6396 ( .B(n4785), .A(n4784), .Z(n4786) );
  XNOR U6397 ( .A(n4787), .B(n4786), .Z(out[996]) );
  ANDN U6398 ( .B(n4789), .A(n4788), .Z(n4790) );
  XNOR U6399 ( .A(n4791), .B(n4790), .Z(out[997]) );
  ANDN U6400 ( .B(n4793), .A(n4792), .Z(n4794) );
  XNOR U6401 ( .A(n4795), .B(n4794), .Z(out[998]) );
  ANDN U6402 ( .B(n4797), .A(n4796), .Z(n4798) );
  XNOR U6403 ( .A(n4799), .B(n4798), .Z(out[999]) );
  ANDN U6404 ( .B(n4801), .A(n4800), .Z(n4802) );
  XNOR U6405 ( .A(n4803), .B(n4802), .Z(out[99]) );
  OR U6406 ( .A(n4805), .B(n4804), .Z(n4806) );
  XNOR U6407 ( .A(n4807), .B(n4806), .Z(out[9]) );
endmodule


module round_3 ( in, round_const, out );
  input [1599:0] in;
  input [63:0] round_const;
  output [1599:0] out;
  wire   round_const_63, round_const_31, round_const_15, round_const_3, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806;
  assign round_const_63 = round_const[63];
  assign round_const_31 = round_const[31];
  assign round_const_15 = round_const[15];
  assign round_const_3 = round_const[3];

  XOR U1 ( .A(in[1469]), .B(in[509]), .Z(n2) );
  XNOR U2 ( .A(in[829]), .B(in[189]), .Z(n1) );
  XNOR U3 ( .A(n2), .B(n1), .Z(n3) );
  XOR U4 ( .A(in[1149]), .B(n3), .Z(n872) );
  XOR U5 ( .A(in[1598]), .B(in[638]), .Z(n5) );
  XNOR U6 ( .A(in[958]), .B(in[318]), .Z(n4) );
  XNOR U7 ( .A(n5), .B(n4), .Z(n6) );
  XOR U8 ( .A(in[1278]), .B(n6), .Z(n1473) );
  XNOR U9 ( .A(n872), .B(n1473), .Z(n3814) );
  XNOR U10 ( .A(in[254]), .B(n3814), .Z(n3576) );
  XOR U11 ( .A(in[1345]), .B(in[65]), .Z(n8) );
  XNOR U12 ( .A(in[1025]), .B(in[385]), .Z(n7) );
  XNOR U13 ( .A(n8), .B(n7), .Z(n9) );
  XOR U14 ( .A(in[705]), .B(n9), .Z(n1481) );
  XOR U15 ( .A(in[1474]), .B(in[514]), .Z(n11) );
  XNOR U16 ( .A(in[834]), .B(in[194]), .Z(n10) );
  XNOR U17 ( .A(n11), .B(n10), .Z(n12) );
  XNOR U18 ( .A(in[1154]), .B(n12), .Z(n1188) );
  XNOR U19 ( .A(n1481), .B(n1188), .Z(n3569) );
  XNOR U20 ( .A(in[1410]), .B(n3569), .Z(n3575) );
  XOR U21 ( .A(in[328]), .B(in[8]), .Z(n14) );
  XNOR U22 ( .A(in[968]), .B(in[648]), .Z(n13) );
  XNOR U23 ( .A(n14), .B(n13), .Z(n15) );
  XOR U24 ( .A(in[1288]), .B(n15), .Z(n1209) );
  XOR U25 ( .A(in[137]), .B(in[457]), .Z(n17) );
  XNOR U26 ( .A(in[777]), .B(in[1417]), .Z(n16) );
  XNOR U27 ( .A(n17), .B(n16), .Z(n18) );
  XOR U28 ( .A(in[1097]), .B(n18), .Z(n1141) );
  XNOR U29 ( .A(n1209), .B(n1141), .Z(n4085) );
  XNOR U30 ( .A(in[1033]), .B(n4085), .Z(n2608) );
  NAND U31 ( .A(n3575), .B(n2608), .Z(n19) );
  XNOR U32 ( .A(n3576), .B(n19), .Z(out[0]) );
  XOR U33 ( .A(in[1515]), .B(in[555]), .Z(n21) );
  XNOR U34 ( .A(in[875]), .B(in[235]), .Z(n20) );
  XNOR U35 ( .A(n21), .B(n20), .Z(n22) );
  XOR U36 ( .A(in[1195]), .B(n22), .Z(n1329) );
  XOR U37 ( .A(in[1386]), .B(in[106]), .Z(n24) );
  XNOR U38 ( .A(in[1066]), .B(in[746]), .Z(n23) );
  XNOR U39 ( .A(n24), .B(n23), .Z(n25) );
  XOR U40 ( .A(in[426]), .B(n25), .Z(n475) );
  XNOR U41 ( .A(n1329), .B(n475), .Z(n3749) );
  XNOR U42 ( .A(in[171]), .B(n3749), .Z(n1301) );
  XOR U43 ( .A(in[971]), .B(in[1291]), .Z(n27) );
  XNOR U44 ( .A(in[11]), .B(in[331]), .Z(n26) );
  XNOR U45 ( .A(n27), .B(n26), .Z(n28) );
  XOR U46 ( .A(in[651]), .B(n28), .Z(n1220) );
  XOR U47 ( .A(in[140]), .B(in[460]), .Z(n30) );
  XNOR U48 ( .A(in[1100]), .B(in[1420]), .Z(n29) );
  XNOR U49 ( .A(n30), .B(n29), .Z(n31) );
  XNOR U50 ( .A(in[780]), .B(n31), .Z(n1159) );
  XNOR U51 ( .A(n1220), .B(n1159), .Z(n4094) );
  XNOR U52 ( .A(in[1356]), .B(n4094), .Z(n1696) );
  XOR U53 ( .A(in[1364]), .B(in[724]), .Z(n33) );
  XNOR U54 ( .A(in[84]), .B(in[404]), .Z(n32) );
  XNOR U55 ( .A(n33), .B(n32), .Z(n34) );
  XOR U56 ( .A(in[1044]), .B(n34), .Z(n777) );
  XOR U57 ( .A(in[1555]), .B(in[595]), .Z(n36) );
  XNOR U58 ( .A(in[915]), .B(in[275]), .Z(n35) );
  XNOR U59 ( .A(n36), .B(n35), .Z(n37) );
  XOR U60 ( .A(in[1235]), .B(n37), .Z(n489) );
  XNOR U61 ( .A(n777), .B(n489), .Z(n3881) );
  XNOR U62 ( .A(in[980]), .B(n3881), .Z(n1693) );
  NAND U63 ( .A(n1696), .B(n1693), .Z(n38) );
  XNOR U64 ( .A(n1301), .B(n38), .Z(out[1000]) );
  XOR U65 ( .A(in[1387]), .B(in[107]), .Z(n40) );
  XNOR U66 ( .A(in[1067]), .B(in[747]), .Z(n39) );
  XNOR U67 ( .A(n40), .B(n39), .Z(n41) );
  XOR U68 ( .A(in[427]), .B(n41), .Z(n486) );
  XOR U69 ( .A(in[1516]), .B(in[556]), .Z(n43) );
  XNOR U70 ( .A(in[876]), .B(in[236]), .Z(n42) );
  XNOR U71 ( .A(n43), .B(n42), .Z(n44) );
  XOR U72 ( .A(in[1196]), .B(n44), .Z(n1333) );
  XNOR U73 ( .A(n486), .B(n1333), .Z(n3757) );
  XNOR U74 ( .A(in[172]), .B(n3757), .Z(n1305) );
  XOR U75 ( .A(in[972]), .B(in[12]), .Z(n46) );
  XNOR U76 ( .A(in[1292]), .B(in[332]), .Z(n45) );
  XNOR U77 ( .A(n46), .B(n45), .Z(n47) );
  XOR U78 ( .A(in[652]), .B(n47), .Z(n1223) );
  XOR U79 ( .A(in[141]), .B(in[461]), .Z(n49) );
  XNOR U80 ( .A(in[1101]), .B(in[1421]), .Z(n48) );
  XNOR U81 ( .A(n49), .B(n48), .Z(n50) );
  XNOR U82 ( .A(in[781]), .B(n50), .Z(n1164) );
  XNOR U83 ( .A(n1223), .B(n1164), .Z(n4097) );
  XNOR U84 ( .A(in[1357]), .B(n4097), .Z(n1700) );
  XOR U85 ( .A(in[1365]), .B(in[725]), .Z(n52) );
  XNOR U86 ( .A(in[85]), .B(in[405]), .Z(n51) );
  XNOR U87 ( .A(n52), .B(n51), .Z(n53) );
  XOR U88 ( .A(in[1045]), .B(n53), .Z(n790) );
  XOR U89 ( .A(in[1556]), .B(in[596]), .Z(n55) );
  XNOR U90 ( .A(in[916]), .B(in[276]), .Z(n54) );
  XNOR U91 ( .A(n55), .B(n54), .Z(n56) );
  XOR U92 ( .A(in[1236]), .B(n56), .Z(n504) );
  XNOR U93 ( .A(n790), .B(n504), .Z(n3883) );
  XNOR U94 ( .A(in[981]), .B(n3883), .Z(n1697) );
  NAND U95 ( .A(n1700), .B(n1697), .Z(n57) );
  XNOR U96 ( .A(n1305), .B(n57), .Z(out[1001]) );
  XOR U97 ( .A(in[1388]), .B(in[108]), .Z(n59) );
  XNOR U98 ( .A(in[1068]), .B(in[748]), .Z(n58) );
  XNOR U99 ( .A(n59), .B(n58), .Z(n60) );
  XOR U100 ( .A(in[428]), .B(n60), .Z(n1395) );
  XOR U101 ( .A(in[1517]), .B(in[557]), .Z(n62) );
  XNOR U102 ( .A(in[877]), .B(in[237]), .Z(n61) );
  XNOR U103 ( .A(n62), .B(n61), .Z(n63) );
  XOR U104 ( .A(in[1197]), .B(n63), .Z(n1337) );
  XNOR U105 ( .A(n1395), .B(n1337), .Z(n3761) );
  XNOR U106 ( .A(in[173]), .B(n3761), .Z(n1310) );
  XOR U107 ( .A(in[142]), .B(in[1422]), .Z(n65) );
  XNOR U108 ( .A(in[1102]), .B(in[782]), .Z(n64) );
  XNOR U109 ( .A(n65), .B(n64), .Z(n66) );
  XOR U110 ( .A(in[462]), .B(n66), .Z(n1169) );
  XOR U111 ( .A(in[973]), .B(in[13]), .Z(n68) );
  XNOR U112 ( .A(in[1293]), .B(in[333]), .Z(n67) );
  XNOR U113 ( .A(n68), .B(n67), .Z(n69) );
  XNOR U114 ( .A(in[653]), .B(n69), .Z(n1226) );
  XNOR U115 ( .A(n1169), .B(n1226), .Z(n4100) );
  XNOR U116 ( .A(in[1358]), .B(n4100), .Z(n1704) );
  XOR U117 ( .A(in[1366]), .B(in[726]), .Z(n71) );
  XNOR U118 ( .A(in[86]), .B(in[406]), .Z(n70) );
  XNOR U119 ( .A(n71), .B(n70), .Z(n72) );
  XOR U120 ( .A(in[1046]), .B(n72), .Z(n803) );
  XOR U121 ( .A(in[1557]), .B(in[597]), .Z(n74) );
  XNOR U122 ( .A(in[917]), .B(in[277]), .Z(n73) );
  XNOR U123 ( .A(n74), .B(n73), .Z(n75) );
  XOR U124 ( .A(in[1237]), .B(n75), .Z(n519) );
  XNOR U125 ( .A(n803), .B(n519), .Z(n3885) );
  XNOR U126 ( .A(in[982]), .B(n3885), .Z(n1701) );
  NAND U127 ( .A(n1704), .B(n1701), .Z(n76) );
  XNOR U128 ( .A(n1310), .B(n76), .Z(out[1002]) );
  XOR U129 ( .A(in[1389]), .B(in[109]), .Z(n78) );
  XNOR U130 ( .A(in[1069]), .B(in[749]), .Z(n77) );
  XNOR U131 ( .A(n78), .B(n77), .Z(n79) );
  XOR U132 ( .A(in[429]), .B(n79), .Z(n1399) );
  XOR U133 ( .A(in[1518]), .B(in[558]), .Z(n81) );
  XNOR U134 ( .A(in[878]), .B(in[238]), .Z(n80) );
  XNOR U135 ( .A(n81), .B(n80), .Z(n82) );
  XOR U136 ( .A(in[1198]), .B(n82), .Z(n1341) );
  XNOR U137 ( .A(n1399), .B(n1341), .Z(n3765) );
  XNOR U138 ( .A(in[174]), .B(n3765), .Z(n1314) );
  XOR U139 ( .A(in[143]), .B(in[1423]), .Z(n84) );
  XNOR U140 ( .A(in[1103]), .B(in[783]), .Z(n83) );
  XNOR U141 ( .A(n84), .B(n83), .Z(n85) );
  XOR U142 ( .A(in[463]), .B(n85), .Z(n1174) );
  XOR U143 ( .A(in[974]), .B(in[14]), .Z(n87) );
  XNOR U144 ( .A(in[1294]), .B(in[334]), .Z(n86) );
  XNOR U145 ( .A(n87), .B(n86), .Z(n88) );
  XNOR U146 ( .A(in[654]), .B(n88), .Z(n1229) );
  XNOR U147 ( .A(n1174), .B(n1229), .Z(n4103) );
  XNOR U148 ( .A(in[1359]), .B(n4103), .Z(n1708) );
  XOR U149 ( .A(in[1367]), .B(in[727]), .Z(n90) );
  XNOR U150 ( .A(in[87]), .B(in[407]), .Z(n89) );
  XNOR U151 ( .A(n90), .B(n89), .Z(n91) );
  XOR U152 ( .A(in[1047]), .B(n91), .Z(n816) );
  XOR U153 ( .A(in[1558]), .B(in[598]), .Z(n93) );
  XNOR U154 ( .A(in[918]), .B(in[278]), .Z(n92) );
  XNOR U155 ( .A(n93), .B(n92), .Z(n94) );
  XOR U156 ( .A(in[1238]), .B(n94), .Z(n534) );
  XNOR U157 ( .A(n816), .B(n534), .Z(n3887) );
  XNOR U158 ( .A(in[983]), .B(n3887), .Z(n1705) );
  NAND U159 ( .A(n1708), .B(n1705), .Z(n95) );
  XNOR U160 ( .A(n1314), .B(n95), .Z(out[1003]) );
  XOR U161 ( .A(in[1390]), .B(in[110]), .Z(n97) );
  XNOR U162 ( .A(in[1070]), .B(in[750]), .Z(n96) );
  XNOR U163 ( .A(n97), .B(n96), .Z(n98) );
  XOR U164 ( .A(in[430]), .B(n98), .Z(n1403) );
  XOR U165 ( .A(in[1519]), .B(in[559]), .Z(n100) );
  XNOR U166 ( .A(in[879]), .B(in[239]), .Z(n99) );
  XNOR U167 ( .A(n100), .B(n99), .Z(n101) );
  XOR U168 ( .A(in[1199]), .B(n101), .Z(n1345) );
  XNOR U169 ( .A(n1403), .B(n1345), .Z(n3769) );
  XNOR U170 ( .A(in[175]), .B(n3769), .Z(n1318) );
  XOR U171 ( .A(in[144]), .B(in[1424]), .Z(n103) );
  XNOR U172 ( .A(in[1104]), .B(in[784]), .Z(n102) );
  XNOR U173 ( .A(n103), .B(n102), .Z(n104) );
  XOR U174 ( .A(in[464]), .B(n104), .Z(n1179) );
  XOR U175 ( .A(in[975]), .B(in[15]), .Z(n106) );
  XNOR U176 ( .A(in[1295]), .B(in[335]), .Z(n105) );
  XNOR U177 ( .A(n106), .B(n105), .Z(n107) );
  XNOR U178 ( .A(in[655]), .B(n107), .Z(n1232) );
  XNOR U179 ( .A(n1179), .B(n1232), .Z(n4106) );
  XNOR U180 ( .A(in[1360]), .B(n4106), .Z(n1713) );
  XOR U181 ( .A(in[1368]), .B(in[728]), .Z(n109) );
  XNOR U182 ( .A(in[88]), .B(in[408]), .Z(n108) );
  XNOR U183 ( .A(n109), .B(n108), .Z(n110) );
  XOR U184 ( .A(in[1048]), .B(n110), .Z(n829) );
  XOR U185 ( .A(in[1559]), .B(in[599]), .Z(n112) );
  XNOR U186 ( .A(in[919]), .B(in[279]), .Z(n111) );
  XNOR U187 ( .A(n112), .B(n111), .Z(n113) );
  XOR U188 ( .A(in[1239]), .B(n113), .Z(n549) );
  XNOR U189 ( .A(n829), .B(n549), .Z(n3889) );
  XNOR U190 ( .A(in[984]), .B(n3889), .Z(n1710) );
  NAND U191 ( .A(n1713), .B(n1710), .Z(n114) );
  XNOR U192 ( .A(n1318), .B(n114), .Z(out[1004]) );
  XOR U193 ( .A(in[1391]), .B(in[111]), .Z(n116) );
  XNOR U194 ( .A(in[1071]), .B(in[751]), .Z(n115) );
  XNOR U195 ( .A(n116), .B(n115), .Z(n117) );
  XOR U196 ( .A(in[431]), .B(n117), .Z(n1407) );
  XOR U197 ( .A(in[1520]), .B(in[560]), .Z(n119) );
  XNOR U198 ( .A(in[880]), .B(in[240]), .Z(n118) );
  XNOR U199 ( .A(n119), .B(n118), .Z(n120) );
  XOR U200 ( .A(in[1200]), .B(n120), .Z(n1350) );
  XNOR U201 ( .A(n1407), .B(n1350), .Z(n3773) );
  XNOR U202 ( .A(in[176]), .B(n3773), .Z(n1322) );
  XOR U203 ( .A(in[145]), .B(in[1425]), .Z(n122) );
  XNOR U204 ( .A(in[1105]), .B(in[785]), .Z(n121) );
  XNOR U205 ( .A(n122), .B(n121), .Z(n123) );
  XOR U206 ( .A(in[465]), .B(n123), .Z(n1184) );
  XOR U207 ( .A(in[976]), .B(in[16]), .Z(n125) );
  XNOR U208 ( .A(in[1296]), .B(in[336]), .Z(n124) );
  XNOR U209 ( .A(n125), .B(n124), .Z(n126) );
  XNOR U210 ( .A(in[656]), .B(n126), .Z(n1235) );
  XNOR U211 ( .A(n1184), .B(n1235), .Z(n4113) );
  XNOR U212 ( .A(in[1361]), .B(n4113), .Z(n1717) );
  XOR U213 ( .A(in[1369]), .B(in[729]), .Z(n128) );
  XNOR U214 ( .A(in[89]), .B(in[409]), .Z(n127) );
  XNOR U215 ( .A(n128), .B(n127), .Z(n129) );
  XOR U216 ( .A(in[1049]), .B(n129), .Z(n842) );
  XOR U217 ( .A(in[1560]), .B(in[600]), .Z(n131) );
  XNOR U218 ( .A(in[920]), .B(in[280]), .Z(n130) );
  XNOR U219 ( .A(n131), .B(n130), .Z(n132) );
  XOR U220 ( .A(in[1240]), .B(n132), .Z(n564) );
  XNOR U221 ( .A(n842), .B(n564), .Z(n3891) );
  XNOR U222 ( .A(in[985]), .B(n3891), .Z(n1714) );
  NAND U223 ( .A(n1717), .B(n1714), .Z(n133) );
  XNOR U224 ( .A(n1322), .B(n133), .Z(out[1005]) );
  XOR U225 ( .A(in[1392]), .B(in[112]), .Z(n135) );
  XNOR U226 ( .A(in[1072]), .B(in[752]), .Z(n134) );
  XNOR U227 ( .A(n135), .B(n134), .Z(n136) );
  XOR U228 ( .A(in[432]), .B(n136), .Z(n1411) );
  XOR U229 ( .A(in[1521]), .B(in[561]), .Z(n138) );
  XNOR U230 ( .A(in[881]), .B(in[241]), .Z(n137) );
  XNOR U231 ( .A(n138), .B(n137), .Z(n139) );
  XOR U232 ( .A(in[1201]), .B(n139), .Z(n1354) );
  XNOR U233 ( .A(n1411), .B(n1354), .Z(n3777) );
  XNOR U234 ( .A(in[177]), .B(n3777), .Z(n1326) );
  XOR U235 ( .A(in[17]), .B(in[657]), .Z(n141) );
  XNOR U236 ( .A(in[977]), .B(in[337]), .Z(n140) );
  XNOR U237 ( .A(n141), .B(n140), .Z(n142) );
  XOR U238 ( .A(in[1297]), .B(n142), .Z(n1238) );
  XOR U239 ( .A(in[1426]), .B(in[466]), .Z(n144) );
  XNOR U240 ( .A(in[786]), .B(in[146]), .Z(n143) );
  XNOR U241 ( .A(n144), .B(n143), .Z(n145) );
  XNOR U242 ( .A(in[1106]), .B(n145), .Z(n488) );
  XNOR U243 ( .A(n1238), .B(n488), .Z(n4116) );
  XNOR U244 ( .A(n4116), .B(in[1362]), .Z(n1721) );
  XOR U245 ( .A(in[1370]), .B(in[730]), .Z(n147) );
  XNOR U246 ( .A(in[90]), .B(in[410]), .Z(n146) );
  XNOR U247 ( .A(n147), .B(n146), .Z(n148) );
  XOR U248 ( .A(in[1050]), .B(n148), .Z(n857) );
  XOR U249 ( .A(in[1561]), .B(in[601]), .Z(n150) );
  XNOR U250 ( .A(in[921]), .B(in[281]), .Z(n149) );
  XNOR U251 ( .A(n150), .B(n149), .Z(n151) );
  XOR U252 ( .A(in[1241]), .B(n151), .Z(n590) );
  XNOR U253 ( .A(n857), .B(n590), .Z(n3893) );
  XNOR U254 ( .A(in[986]), .B(n3893), .Z(n1718) );
  NAND U255 ( .A(n1721), .B(n1718), .Z(n152) );
  XNOR U256 ( .A(n1326), .B(n152), .Z(out[1006]) );
  XOR U257 ( .A(in[1393]), .B(in[113]), .Z(n154) );
  XNOR U258 ( .A(in[1073]), .B(in[753]), .Z(n153) );
  XNOR U259 ( .A(n154), .B(n153), .Z(n155) );
  XOR U260 ( .A(in[433]), .B(n155), .Z(n1415) );
  XOR U261 ( .A(in[1522]), .B(in[562]), .Z(n157) );
  XNOR U262 ( .A(in[882]), .B(in[242]), .Z(n156) );
  XNOR U263 ( .A(n157), .B(n156), .Z(n158) );
  XOR U264 ( .A(in[1202]), .B(n158), .Z(n1358) );
  XNOR U265 ( .A(n1415), .B(n1358), .Z(n3781) );
  XNOR U266 ( .A(in[178]), .B(n3781), .Z(n1330) );
  XOR U267 ( .A(in[147]), .B(in[1427]), .Z(n160) );
  XNOR U268 ( .A(in[1107]), .B(in[787]), .Z(n159) );
  XNOR U269 ( .A(n160), .B(n159), .Z(n161) );
  XOR U270 ( .A(in[467]), .B(n161), .Z(n503) );
  XOR U271 ( .A(in[978]), .B(in[18]), .Z(n163) );
  XNOR U272 ( .A(in[1298]), .B(in[338]), .Z(n162) );
  XNOR U273 ( .A(n163), .B(n162), .Z(n164) );
  XNOR U274 ( .A(in[658]), .B(n164), .Z(n1241) );
  XNOR U275 ( .A(n503), .B(n1241), .Z(n4119) );
  XNOR U276 ( .A(in[1363]), .B(n4119), .Z(n1725) );
  XOR U277 ( .A(in[1371]), .B(in[731]), .Z(n166) );
  XNOR U278 ( .A(in[91]), .B(in[411]), .Z(n165) );
  XNOR U279 ( .A(n166), .B(n165), .Z(n167) );
  XOR U280 ( .A(in[1051]), .B(n167), .Z(n870) );
  XOR U281 ( .A(in[1562]), .B(in[602]), .Z(n169) );
  XNOR U282 ( .A(in[922]), .B(in[282]), .Z(n168) );
  XNOR U283 ( .A(n169), .B(n168), .Z(n170) );
  XOR U284 ( .A(in[1242]), .B(n170), .Z(n605) );
  XNOR U285 ( .A(n870), .B(n605), .Z(n3895) );
  XNOR U286 ( .A(in[987]), .B(n3895), .Z(n1722) );
  NAND U287 ( .A(n1725), .B(n1722), .Z(n171) );
  XNOR U288 ( .A(n1330), .B(n171), .Z(out[1007]) );
  XOR U289 ( .A(in[1394]), .B(in[114]), .Z(n173) );
  XNOR U290 ( .A(in[1074]), .B(in[754]), .Z(n172) );
  XNOR U291 ( .A(n173), .B(n172), .Z(n174) );
  XOR U292 ( .A(in[434]), .B(n174), .Z(n1419) );
  XOR U293 ( .A(in[1523]), .B(in[563]), .Z(n176) );
  XNOR U294 ( .A(in[883]), .B(in[243]), .Z(n175) );
  XNOR U295 ( .A(n176), .B(n175), .Z(n177) );
  XOR U296 ( .A(in[1203]), .B(n177), .Z(n1362) );
  XNOR U297 ( .A(n1419), .B(n1362), .Z(n3785) );
  XNOR U298 ( .A(in[179]), .B(n3785), .Z(n1334) );
  XOR U299 ( .A(in[979]), .B(in[19]), .Z(n179) );
  XNOR U300 ( .A(in[1299]), .B(in[339]), .Z(n178) );
  XNOR U301 ( .A(n179), .B(n178), .Z(n180) );
  XOR U302 ( .A(in[659]), .B(n180), .Z(n1245) );
  XOR U303 ( .A(in[148]), .B(in[1428]), .Z(n182) );
  XNOR U304 ( .A(in[1108]), .B(in[788]), .Z(n181) );
  XNOR U305 ( .A(n182), .B(n181), .Z(n183) );
  XNOR U306 ( .A(in[468]), .B(n183), .Z(n518) );
  XNOR U307 ( .A(n1245), .B(n518), .Z(n4122) );
  XNOR U308 ( .A(in[1364]), .B(n4122), .Z(n1729) );
  XOR U309 ( .A(in[1372]), .B(in[732]), .Z(n185) );
  XNOR U310 ( .A(in[92]), .B(in[412]), .Z(n184) );
  XNOR U311 ( .A(n185), .B(n184), .Z(n186) );
  XOR U312 ( .A(in[1052]), .B(n186), .Z(n890) );
  XOR U313 ( .A(in[1563]), .B(in[603]), .Z(n188) );
  XNOR U314 ( .A(in[923]), .B(in[283]), .Z(n187) );
  XNOR U315 ( .A(n188), .B(n187), .Z(n189) );
  XOR U316 ( .A(in[1243]), .B(n189), .Z(n620) );
  XNOR U317 ( .A(n890), .B(n620), .Z(n3899) );
  XNOR U318 ( .A(in[988]), .B(n3899), .Z(n1726) );
  NAND U319 ( .A(n1729), .B(n1726), .Z(n190) );
  XNOR U320 ( .A(n1334), .B(n190), .Z(out[1008]) );
  XOR U321 ( .A(in[1395]), .B(in[115]), .Z(n192) );
  XNOR U322 ( .A(in[1075]), .B(in[755]), .Z(n191) );
  XNOR U323 ( .A(n192), .B(n191), .Z(n193) );
  XOR U324 ( .A(in[435]), .B(n193), .Z(n1423) );
  XOR U325 ( .A(in[1524]), .B(in[564]), .Z(n195) );
  XNOR U326 ( .A(in[884]), .B(in[244]), .Z(n194) );
  XNOR U327 ( .A(n195), .B(n194), .Z(n196) );
  XOR U328 ( .A(in[1204]), .B(n196), .Z(n1366) );
  XNOR U329 ( .A(n1423), .B(n1366), .Z(n3789) );
  XNOR U330 ( .A(in[180]), .B(n3789), .Z(n1338) );
  XOR U331 ( .A(in[340]), .B(in[660]), .Z(n198) );
  XNOR U332 ( .A(in[20]), .B(in[1300]), .Z(n197) );
  XNOR U333 ( .A(n198), .B(n197), .Z(n199) );
  XOR U334 ( .A(in[980]), .B(n199), .Z(n1248) );
  XOR U335 ( .A(in[149]), .B(in[1429]), .Z(n201) );
  XNOR U336 ( .A(in[1109]), .B(in[789]), .Z(n200) );
  XNOR U337 ( .A(n201), .B(n200), .Z(n202) );
  XNOR U338 ( .A(in[469]), .B(n202), .Z(n533) );
  XNOR U339 ( .A(n1248), .B(n533), .Z(n4125) );
  XNOR U340 ( .A(in[1365]), .B(n4125), .Z(n1733) );
  XOR U341 ( .A(in[1373]), .B(in[733]), .Z(n204) );
  XNOR U342 ( .A(in[93]), .B(in[413]), .Z(n203) );
  XNOR U343 ( .A(n204), .B(n203), .Z(n205) );
  XOR U344 ( .A(in[1053]), .B(n205), .Z(n903) );
  XOR U345 ( .A(in[1564]), .B(in[604]), .Z(n207) );
  XNOR U346 ( .A(in[924]), .B(in[284]), .Z(n206) );
  XNOR U347 ( .A(n207), .B(n206), .Z(n208) );
  XOR U348 ( .A(in[1244]), .B(n208), .Z(n635) );
  XNOR U349 ( .A(n903), .B(n635), .Z(n3901) );
  XNOR U350 ( .A(in[989]), .B(n3901), .Z(n1730) );
  NAND U351 ( .A(n1733), .B(n1730), .Z(n209) );
  XNOR U352 ( .A(n1338), .B(n209), .Z(out[1009]) );
  XOR U353 ( .A(in[1339]), .B(in[59]), .Z(n211) );
  XNOR U354 ( .A(in[699]), .B(in[379]), .Z(n210) );
  XNOR U355 ( .A(n211), .B(n210), .Z(n212) );
  XOR U356 ( .A(in[1019]), .B(n212), .Z(n861) );
  XOR U357 ( .A(in[1530]), .B(in[570]), .Z(n214) );
  XNOR U358 ( .A(in[1210]), .B(in[250]), .Z(n213) );
  XNOR U359 ( .A(n214), .B(n213), .Z(n215) );
  XOR U360 ( .A(in[890]), .B(n215), .Z(n327) );
  XNOR U361 ( .A(n861), .B(n327), .Z(n3591) );
  XNOR U362 ( .A(in[635]), .B(n3591), .Z(n2549) );
  XOR U363 ( .A(in[161]), .B(in[1441]), .Z(n217) );
  XNOR U364 ( .A(in[801]), .B(in[1121]), .Z(n216) );
  XNOR U365 ( .A(n217), .B(n216), .Z(n218) );
  XOR U366 ( .A(in[481]), .B(n218), .Z(n454) );
  XOR U367 ( .A(in[1570]), .B(in[610]), .Z(n220) );
  XNOR U368 ( .A(in[930]), .B(in[290]), .Z(n219) );
  XNOR U369 ( .A(n220), .B(n219), .Z(n221) );
  XNOR U370 ( .A(in[1250]), .B(n221), .Z(n337) );
  XNOR U371 ( .A(n454), .B(n337), .Z(n3688) );
  XNOR U372 ( .A(in[226]), .B(n3688), .Z(n2830) );
  XOR U373 ( .A(in[1061]), .B(in[421]), .Z(n223) );
  XNOR U374 ( .A(in[741]), .B(in[1381]), .Z(n222) );
  XNOR U375 ( .A(n223), .B(n222), .Z(n224) );
  XOR U376 ( .A(in[101]), .B(n224), .Z(n373) );
  XOR U377 ( .A(in[1510]), .B(in[550]), .Z(n226) );
  XNOR U378 ( .A(in[870]), .B(in[230]), .Z(n225) );
  XNOR U379 ( .A(n226), .B(n225), .Z(n227) );
  XOR U380 ( .A(in[1190]), .B(n227), .Z(n1309) );
  XNOR U381 ( .A(n373), .B(n1309), .Z(n3729) );
  XNOR U382 ( .A(in[1446]), .B(n3729), .Z(n2827) );
  NAND U383 ( .A(n2830), .B(n2827), .Z(n228) );
  XNOR U384 ( .A(n2549), .B(n228), .Z(out[100]) );
  XOR U385 ( .A(in[1396]), .B(in[116]), .Z(n230) );
  XNOR U386 ( .A(in[1076]), .B(in[756]), .Z(n229) );
  XNOR U387 ( .A(n230), .B(n229), .Z(n231) );
  XOR U388 ( .A(in[436]), .B(n231), .Z(n1428) );
  XOR U389 ( .A(in[1525]), .B(in[565]), .Z(n233) );
  XNOR U390 ( .A(in[885]), .B(in[245]), .Z(n232) );
  XNOR U391 ( .A(n233), .B(n232), .Z(n234) );
  XOR U392 ( .A(in[1205]), .B(n234), .Z(n1370) );
  XNOR U393 ( .A(n1428), .B(n1370), .Z(n3793) );
  XNOR U394 ( .A(in[181]), .B(n3793), .Z(n1342) );
  XOR U395 ( .A(in[341]), .B(in[661]), .Z(n236) );
  XNOR U396 ( .A(in[21]), .B(in[1301]), .Z(n235) );
  XNOR U397 ( .A(n236), .B(n235), .Z(n237) );
  XOR U398 ( .A(in[981]), .B(n237), .Z(n1251) );
  XOR U399 ( .A(in[150]), .B(in[1430]), .Z(n239) );
  XNOR U400 ( .A(in[1110]), .B(in[790]), .Z(n238) );
  XNOR U401 ( .A(n239), .B(n238), .Z(n240) );
  XNOR U402 ( .A(in[470]), .B(n240), .Z(n548) );
  XNOR U403 ( .A(n1251), .B(n548), .Z(n4128) );
  XNOR U404 ( .A(in[1366]), .B(n4128), .Z(n1737) );
  XOR U405 ( .A(in[1374]), .B(in[734]), .Z(n242) );
  XNOR U406 ( .A(in[94]), .B(in[414]), .Z(n241) );
  XNOR U407 ( .A(n242), .B(n241), .Z(n243) );
  XOR U408 ( .A(in[1054]), .B(n243), .Z(n916) );
  XOR U409 ( .A(in[1565]), .B(in[605]), .Z(n245) );
  XNOR U410 ( .A(in[925]), .B(in[285]), .Z(n244) );
  XNOR U411 ( .A(n245), .B(n244), .Z(n246) );
  XOR U412 ( .A(in[1245]), .B(n246), .Z(n650) );
  XNOR U413 ( .A(n916), .B(n650), .Z(n3903) );
  XNOR U414 ( .A(in[990]), .B(n3903), .Z(n1734) );
  NAND U415 ( .A(n1737), .B(n1734), .Z(n247) );
  XNOR U416 ( .A(n1342), .B(n247), .Z(out[1010]) );
  XOR U417 ( .A(in[1526]), .B(in[566]), .Z(n249) );
  XNOR U418 ( .A(in[886]), .B(in[246]), .Z(n248) );
  XNOR U419 ( .A(n249), .B(n248), .Z(n250) );
  XOR U420 ( .A(in[1206]), .B(n250), .Z(n1374) );
  XOR U421 ( .A(in[1397]), .B(in[117]), .Z(n252) );
  XNOR U422 ( .A(in[1077]), .B(in[757]), .Z(n251) );
  XNOR U423 ( .A(n252), .B(n251), .Z(n253) );
  XOR U424 ( .A(in[437]), .B(n253), .Z(n1432) );
  XNOR U425 ( .A(n1374), .B(n1432), .Z(n3803) );
  XNOR U426 ( .A(in[182]), .B(n3803), .Z(n1346) );
  XOR U427 ( .A(in[342]), .B(in[662]), .Z(n255) );
  XNOR U428 ( .A(in[22]), .B(in[1302]), .Z(n254) );
  XNOR U429 ( .A(n255), .B(n254), .Z(n256) );
  XOR U430 ( .A(in[982]), .B(n256), .Z(n1254) );
  XOR U431 ( .A(in[151]), .B(in[1431]), .Z(n258) );
  XNOR U432 ( .A(in[1111]), .B(in[791]), .Z(n257) );
  XNOR U433 ( .A(n258), .B(n257), .Z(n259) );
  XNOR U434 ( .A(in[471]), .B(n259), .Z(n563) );
  XNOR U435 ( .A(n1254), .B(n563), .Z(n4131) );
  XNOR U436 ( .A(in[1367]), .B(n4131), .Z(n1741) );
  XOR U437 ( .A(in[1375]), .B(in[735]), .Z(n261) );
  XNOR U438 ( .A(in[95]), .B(in[415]), .Z(n260) );
  XNOR U439 ( .A(n261), .B(n260), .Z(n262) );
  XOR U440 ( .A(in[1055]), .B(n262), .Z(n929) );
  XOR U441 ( .A(in[1566]), .B(in[606]), .Z(n264) );
  XNOR U442 ( .A(in[926]), .B(in[286]), .Z(n263) );
  XNOR U443 ( .A(n264), .B(n263), .Z(n265) );
  XOR U444 ( .A(in[1246]), .B(n265), .Z(n665) );
  XNOR U445 ( .A(n929), .B(n665), .Z(n3905) );
  XNOR U446 ( .A(in[991]), .B(n3905), .Z(n1738) );
  NAND U447 ( .A(n1741), .B(n1738), .Z(n266) );
  XNOR U448 ( .A(n1346), .B(n266), .Z(out[1011]) );
  XOR U449 ( .A(in[1527]), .B(in[567]), .Z(n268) );
  XNOR U450 ( .A(in[887]), .B(in[247]), .Z(n267) );
  XNOR U451 ( .A(n268), .B(n267), .Z(n269) );
  XOR U452 ( .A(in[1207]), .B(n269), .Z(n1378) );
  XOR U453 ( .A(in[1398]), .B(in[118]), .Z(n271) );
  XNOR U454 ( .A(in[1078]), .B(in[758]), .Z(n270) );
  XNOR U455 ( .A(n271), .B(n270), .Z(n272) );
  XOR U456 ( .A(in[438]), .B(n272), .Z(n1436) );
  XNOR U457 ( .A(n1378), .B(n1436), .Z(n3807) );
  XNOR U458 ( .A(in[183]), .B(n3807), .Z(n1351) );
  XOR U459 ( .A(in[152]), .B(in[1432]), .Z(n274) );
  XNOR U460 ( .A(in[1112]), .B(in[792]), .Z(n273) );
  XNOR U461 ( .A(n274), .B(n273), .Z(n275) );
  XOR U462 ( .A(in[472]), .B(n275), .Z(n589) );
  XOR U463 ( .A(in[343]), .B(in[663]), .Z(n277) );
  XNOR U464 ( .A(in[23]), .B(in[1303]), .Z(n276) );
  XNOR U465 ( .A(n277), .B(n276), .Z(n278) );
  XNOR U466 ( .A(in[983]), .B(n278), .Z(n1257) );
  XNOR U467 ( .A(n589), .B(n1257), .Z(n4134) );
  XNOR U468 ( .A(in[1368]), .B(n4134), .Z(n1745) );
  XOR U469 ( .A(in[1376]), .B(in[736]), .Z(n280) );
  XNOR U470 ( .A(in[96]), .B(in[416]), .Z(n279) );
  XNOR U471 ( .A(n280), .B(n279), .Z(n281) );
  XOR U472 ( .A(in[1056]), .B(n281), .Z(n944) );
  XOR U473 ( .A(in[1567]), .B(in[607]), .Z(n283) );
  XNOR U474 ( .A(in[927]), .B(in[287]), .Z(n282) );
  XNOR U475 ( .A(n283), .B(n282), .Z(n284) );
  XOR U476 ( .A(in[1247]), .B(n284), .Z(n680) );
  XNOR U477 ( .A(n944), .B(n680), .Z(n3907) );
  XNOR U478 ( .A(in[992]), .B(n3907), .Z(n1742) );
  NAND U479 ( .A(n1745), .B(n1742), .Z(n285) );
  XNOR U480 ( .A(n1351), .B(n285), .Z(out[1012]) );
  XOR U481 ( .A(in[1528]), .B(in[568]), .Z(n287) );
  XNOR U482 ( .A(in[888]), .B(in[248]), .Z(n286) );
  XNOR U483 ( .A(n287), .B(n286), .Z(n288) );
  XOR U484 ( .A(in[1208]), .B(n288), .Z(n1382) );
  XOR U485 ( .A(in[1399]), .B(in[119]), .Z(n290) );
  XNOR U486 ( .A(in[1079]), .B(in[759]), .Z(n289) );
  XNOR U487 ( .A(n290), .B(n289), .Z(n291) );
  XOR U488 ( .A(in[439]), .B(n291), .Z(n1440) );
  XNOR U489 ( .A(n1382), .B(n1440), .Z(n3811) );
  XNOR U490 ( .A(in[184]), .B(n3811), .Z(n1355) );
  XOR U491 ( .A(in[153]), .B(in[1433]), .Z(n293) );
  XNOR U492 ( .A(in[1113]), .B(in[793]), .Z(n292) );
  XNOR U493 ( .A(n293), .B(n292), .Z(n294) );
  XOR U494 ( .A(in[473]), .B(n294), .Z(n604) );
  XOR U495 ( .A(in[344]), .B(in[664]), .Z(n296) );
  XNOR U496 ( .A(in[24]), .B(in[1304]), .Z(n295) );
  XNOR U497 ( .A(n296), .B(n295), .Z(n297) );
  XNOR U498 ( .A(in[984]), .B(n297), .Z(n1260) );
  XNOR U499 ( .A(n604), .B(n1260), .Z(n4137) );
  XNOR U500 ( .A(in[1369]), .B(n4137), .Z(n1749) );
  XOR U501 ( .A(in[1377]), .B(in[737]), .Z(n299) );
  XNOR U502 ( .A(in[97]), .B(in[417]), .Z(n298) );
  XNOR U503 ( .A(n299), .B(n298), .Z(n300) );
  XOR U504 ( .A(in[1057]), .B(n300), .Z(n959) );
  XOR U505 ( .A(in[1568]), .B(in[608]), .Z(n302) );
  XNOR U506 ( .A(in[928]), .B(in[288]), .Z(n301) );
  XNOR U507 ( .A(n302), .B(n301), .Z(n303) );
  XOR U508 ( .A(in[1248]), .B(n303), .Z(n695) );
  XNOR U509 ( .A(n959), .B(n695), .Z(n3909) );
  XNOR U510 ( .A(in[993]), .B(n3909), .Z(n1746) );
  NAND U511 ( .A(n1749), .B(n1746), .Z(n304) );
  XNOR U512 ( .A(n1355), .B(n304), .Z(out[1013]) );
  XOR U513 ( .A(in[1529]), .B(in[569]), .Z(n306) );
  XNOR U514 ( .A(in[889]), .B(in[249]), .Z(n305) );
  XNOR U515 ( .A(n306), .B(n305), .Z(n307) );
  XOR U516 ( .A(in[1209]), .B(n307), .Z(n1386) );
  XOR U517 ( .A(in[1400]), .B(in[120]), .Z(n309) );
  XNOR U518 ( .A(in[1080]), .B(in[760]), .Z(n308) );
  XNOR U519 ( .A(n309), .B(n308), .Z(n310) );
  XOR U520 ( .A(in[440]), .B(n310), .Z(n1444) );
  XNOR U521 ( .A(n1386), .B(n1444), .Z(n3815) );
  XNOR U522 ( .A(in[185]), .B(n3815), .Z(n1359) );
  XOR U523 ( .A(in[345]), .B(in[665]), .Z(n312) );
  XNOR U524 ( .A(in[25]), .B(in[1305]), .Z(n311) );
  XNOR U525 ( .A(n312), .B(n311), .Z(n313) );
  XOR U526 ( .A(in[985]), .B(n313), .Z(n1263) );
  XOR U527 ( .A(in[154]), .B(in[1434]), .Z(n315) );
  XNOR U528 ( .A(in[1114]), .B(in[794]), .Z(n314) );
  XNOR U529 ( .A(n315), .B(n314), .Z(n316) );
  XNOR U530 ( .A(in[474]), .B(n316), .Z(n619) );
  XNOR U531 ( .A(n1263), .B(n619), .Z(n4140) );
  XNOR U532 ( .A(in[1370]), .B(n4140), .Z(n1754) );
  XOR U533 ( .A(in[1569]), .B(in[609]), .Z(n318) );
  XNOR U534 ( .A(in[929]), .B(in[289]), .Z(n317) );
  XNOR U535 ( .A(n318), .B(n317), .Z(n319) );
  XOR U536 ( .A(in[1249]), .B(n319), .Z(n710) );
  XOR U537 ( .A(in[1378]), .B(in[738]), .Z(n321) );
  XNOR U538 ( .A(in[98]), .B(in[418]), .Z(n320) );
  XNOR U539 ( .A(n321), .B(n320), .Z(n322) );
  XOR U540 ( .A(in[1058]), .B(n322), .Z(n974) );
  XNOR U541 ( .A(n710), .B(n974), .Z(n3911) );
  XNOR U542 ( .A(in[994]), .B(n3911), .Z(n1751) );
  NAND U543 ( .A(n1754), .B(n1751), .Z(n323) );
  XNOR U544 ( .A(n1359), .B(n323), .Z(out[1014]) );
  XOR U545 ( .A(in[1401]), .B(in[121]), .Z(n325) );
  XNOR U546 ( .A(in[1081]), .B(in[761]), .Z(n324) );
  XNOR U547 ( .A(n325), .B(n324), .Z(n326) );
  XOR U548 ( .A(in[441]), .B(n326), .Z(n1448) );
  XNOR U549 ( .A(n327), .B(n1448), .Z(n3537) );
  XNOR U550 ( .A(in[186]), .B(n3537), .Z(n1363) );
  XOR U551 ( .A(in[155]), .B(in[1435]), .Z(n329) );
  XNOR U552 ( .A(in[1115]), .B(in[795]), .Z(n328) );
  XNOR U553 ( .A(n329), .B(n328), .Z(n330) );
  XOR U554 ( .A(in[475]), .B(n330), .Z(n634) );
  XOR U555 ( .A(in[346]), .B(in[666]), .Z(n332) );
  XNOR U556 ( .A(in[26]), .B(in[1306]), .Z(n331) );
  XNOR U557 ( .A(n332), .B(n331), .Z(n333) );
  XNOR U558 ( .A(in[986]), .B(n333), .Z(n1266) );
  XNOR U559 ( .A(n634), .B(n1266), .Z(n4147) );
  XNOR U560 ( .A(in[1371]), .B(n4147), .Z(n1758) );
  XOR U561 ( .A(in[1379]), .B(in[739]), .Z(n335) );
  XNOR U562 ( .A(in[99]), .B(in[419]), .Z(n334) );
  XNOR U563 ( .A(n335), .B(n334), .Z(n336) );
  XNOR U564 ( .A(in[1059]), .B(n336), .Z(n989) );
  XNOR U565 ( .A(n337), .B(n989), .Z(n3913) );
  XNOR U566 ( .A(in[995]), .B(n3913), .Z(n1755) );
  NAND U567 ( .A(n1758), .B(n1755), .Z(n338) );
  XNOR U568 ( .A(n1363), .B(n338), .Z(out[1015]) );
  XOR U569 ( .A(in[1402]), .B(in[122]), .Z(n340) );
  XNOR U570 ( .A(in[1082]), .B(in[762]), .Z(n339) );
  XNOR U571 ( .A(n340), .B(n339), .Z(n341) );
  XOR U572 ( .A(in[442]), .B(n341), .Z(n1452) );
  XOR U573 ( .A(in[1531]), .B(in[571]), .Z(n343) );
  XNOR U574 ( .A(in[1211]), .B(in[251]), .Z(n342) );
  XNOR U575 ( .A(n343), .B(n342), .Z(n344) );
  XOR U576 ( .A(in[891]), .B(n344), .Z(n416) );
  XNOR U577 ( .A(n1452), .B(n416), .Z(n3541) );
  XNOR U578 ( .A(in[187]), .B(n3541), .Z(n1367) );
  XOR U579 ( .A(in[156]), .B(in[1436]), .Z(n346) );
  XNOR U580 ( .A(in[1116]), .B(in[796]), .Z(n345) );
  XNOR U581 ( .A(n346), .B(n345), .Z(n347) );
  XOR U582 ( .A(in[476]), .B(n347), .Z(n649) );
  XOR U583 ( .A(in[347]), .B(in[667]), .Z(n349) );
  XNOR U584 ( .A(in[27]), .B(in[1307]), .Z(n348) );
  XNOR U585 ( .A(n349), .B(n348), .Z(n350) );
  XNOR U586 ( .A(in[987]), .B(n350), .Z(n1269) );
  XNOR U587 ( .A(n649), .B(n1269), .Z(n4150) );
  XNOR U588 ( .A(in[1372]), .B(n4150), .Z(n1762) );
  XOR U589 ( .A(in[1060]), .B(in[420]), .Z(n352) );
  XNOR U590 ( .A(in[740]), .B(in[1380]), .Z(n351) );
  XNOR U591 ( .A(n352), .B(n351), .Z(n353) );
  XOR U592 ( .A(in[100]), .B(n353), .Z(n1004) );
  XOR U593 ( .A(in[1571]), .B(in[611]), .Z(n355) );
  XNOR U594 ( .A(in[931]), .B(in[291]), .Z(n354) );
  XNOR U595 ( .A(n355), .B(n354), .Z(n356) );
  XOR U596 ( .A(in[1251]), .B(n356), .Z(n420) );
  XNOR U597 ( .A(n1004), .B(n420), .Z(n3915) );
  XNOR U598 ( .A(in[996]), .B(n3915), .Z(n1759) );
  NAND U599 ( .A(n1762), .B(n1759), .Z(n357) );
  XNOR U600 ( .A(n1367), .B(n357), .Z(out[1016]) );
  XOR U601 ( .A(in[1403]), .B(in[123]), .Z(n359) );
  XNOR U602 ( .A(in[1083]), .B(in[763]), .Z(n358) );
  XNOR U603 ( .A(n359), .B(n358), .Z(n360) );
  XOR U604 ( .A(in[443]), .B(n360), .Z(n1456) );
  XOR U605 ( .A(in[1532]), .B(in[572]), .Z(n362) );
  XNOR U606 ( .A(in[1212]), .B(in[252]), .Z(n361) );
  XNOR U607 ( .A(n362), .B(n361), .Z(n363) );
  XOR U608 ( .A(in[892]), .B(n363), .Z(n581) );
  XNOR U609 ( .A(n1456), .B(n581), .Z(n3545) );
  XNOR U610 ( .A(in[188]), .B(n3545), .Z(n1371) );
  XOR U611 ( .A(in[157]), .B(in[1437]), .Z(n365) );
  XNOR U612 ( .A(in[1117]), .B(in[797]), .Z(n364) );
  XNOR U613 ( .A(n365), .B(n364), .Z(n366) );
  XOR U614 ( .A(in[477]), .B(n366), .Z(n664) );
  XOR U615 ( .A(in[348]), .B(in[668]), .Z(n368) );
  XNOR U616 ( .A(in[28]), .B(in[1308]), .Z(n367) );
  XNOR U617 ( .A(n368), .B(n367), .Z(n369) );
  XNOR U618 ( .A(in[988]), .B(n369), .Z(n1272) );
  XNOR U619 ( .A(n664), .B(n1272), .Z(n4153) );
  XNOR U620 ( .A(in[1373]), .B(n4153), .Z(n1766) );
  XOR U621 ( .A(in[1572]), .B(in[612]), .Z(n371) );
  XNOR U622 ( .A(in[932]), .B(in[292]), .Z(n370) );
  XNOR U623 ( .A(n371), .B(n370), .Z(n372) );
  XOR U624 ( .A(in[1252]), .B(n372), .Z(n583) );
  XNOR U625 ( .A(n373), .B(n583), .Z(n3917) );
  XNOR U626 ( .A(in[997]), .B(n3917), .Z(n1763) );
  NAND U627 ( .A(n1766), .B(n1763), .Z(n374) );
  XNOR U628 ( .A(n1371), .B(n374), .Z(out[1017]) );
  XOR U629 ( .A(in[1404]), .B(in[124]), .Z(n376) );
  XNOR U630 ( .A(in[1084]), .B(in[764]), .Z(n375) );
  XNOR U631 ( .A(n376), .B(n375), .Z(n377) );
  XOR U632 ( .A(in[444]), .B(n377), .Z(n1460) );
  XOR U633 ( .A(in[1533]), .B(in[573]), .Z(n379) );
  XNOR U634 ( .A(in[1213]), .B(in[253]), .Z(n378) );
  XNOR U635 ( .A(n379), .B(n378), .Z(n380) );
  XOR U636 ( .A(in[893]), .B(n380), .Z(n740) );
  XNOR U637 ( .A(n1460), .B(n740), .Z(n3549) );
  XNOR U638 ( .A(in[189]), .B(n3549), .Z(n1375) );
  XOR U639 ( .A(in[158]), .B(in[1438]), .Z(n382) );
  XNOR U640 ( .A(in[1118]), .B(in[798]), .Z(n381) );
  XNOR U641 ( .A(n382), .B(n381), .Z(n383) );
  XOR U642 ( .A(in[478]), .B(n383), .Z(n679) );
  XOR U643 ( .A(in[349]), .B(in[669]), .Z(n385) );
  XNOR U644 ( .A(in[29]), .B(in[1309]), .Z(n384) );
  XNOR U645 ( .A(n385), .B(n384), .Z(n386) );
  XNOR U646 ( .A(in[989]), .B(n386), .Z(n1276) );
  XNOR U647 ( .A(n679), .B(n1276), .Z(n4156) );
  XNOR U648 ( .A(in[1374]), .B(n4156), .Z(n1770) );
  XOR U649 ( .A(in[1062]), .B(in[422]), .Z(n388) );
  XNOR U650 ( .A(in[742]), .B(in[1382]), .Z(n387) );
  XNOR U651 ( .A(n388), .B(n387), .Z(n389) );
  XOR U652 ( .A(in[102]), .B(n389), .Z(n424) );
  XOR U653 ( .A(in[1573]), .B(in[613]), .Z(n391) );
  XNOR U654 ( .A(in[933]), .B(in[293]), .Z(n390) );
  XNOR U655 ( .A(n391), .B(n390), .Z(n392) );
  XOR U656 ( .A(in[1253]), .B(n392), .Z(n742) );
  XNOR U657 ( .A(n424), .B(n742), .Z(n3923) );
  XNOR U658 ( .A(in[998]), .B(n3923), .Z(n1767) );
  NAND U659 ( .A(n1770), .B(n1767), .Z(n393) );
  XNOR U660 ( .A(n1375), .B(n393), .Z(out[1018]) );
  XOR U661 ( .A(in[1405]), .B(in[125]), .Z(n395) );
  XNOR U662 ( .A(in[1085]), .B(in[765]), .Z(n394) );
  XNOR U663 ( .A(n395), .B(n394), .Z(n396) );
  XOR U664 ( .A(in[445]), .B(n396), .Z(n1464) );
  XOR U665 ( .A(in[1534]), .B(in[894]), .Z(n398) );
  XNOR U666 ( .A(in[574]), .B(in[1214]), .Z(n397) );
  XNOR U667 ( .A(n398), .B(n397), .Z(n399) );
  XOR U668 ( .A(in[254]), .B(n399), .Z(n877) );
  XNOR U669 ( .A(n1464), .B(n877), .Z(n3553) );
  XNOR U670 ( .A(in[190]), .B(n3553), .Z(n1379) );
  XOR U671 ( .A(in[1439]), .B(in[479]), .Z(n401) );
  XNOR U672 ( .A(in[799]), .B(in[159]), .Z(n400) );
  XNOR U673 ( .A(n401), .B(n400), .Z(n402) );
  XOR U674 ( .A(in[1119]), .B(n402), .Z(n694) );
  XOR U675 ( .A(in[350]), .B(in[670]), .Z(n404) );
  XNOR U676 ( .A(in[30]), .B(in[1310]), .Z(n403) );
  XNOR U677 ( .A(n404), .B(n403), .Z(n405) );
  XNOR U678 ( .A(in[990]), .B(n405), .Z(n1279) );
  XNOR U679 ( .A(n694), .B(n1279), .Z(n4159) );
  XNOR U680 ( .A(in[1375]), .B(n4159), .Z(n1774) );
  XOR U681 ( .A(in[1063]), .B(in[423]), .Z(n407) );
  XNOR U682 ( .A(in[743]), .B(in[1383]), .Z(n406) );
  XNOR U683 ( .A(n407), .B(n406), .Z(n408) );
  XOR U684 ( .A(in[103]), .B(n408), .Z(n587) );
  XOR U685 ( .A(in[1574]), .B(in[614]), .Z(n410) );
  XNOR U686 ( .A(in[934]), .B(in[294]), .Z(n409) );
  XNOR U687 ( .A(n410), .B(n409), .Z(n411) );
  XOR U688 ( .A(in[1254]), .B(n411), .Z(n786) );
  XNOR U689 ( .A(n587), .B(n786), .Z(n3925) );
  XNOR U690 ( .A(in[999]), .B(n3925), .Z(n1771) );
  NAND U691 ( .A(n1774), .B(n1771), .Z(n412) );
  XNOR U692 ( .A(n1379), .B(n412), .Z(out[1019]) );
  XOR U693 ( .A(in[1340]), .B(in[60]), .Z(n414) );
  XNOR U694 ( .A(in[700]), .B(in[380]), .Z(n413) );
  XNOR U695 ( .A(n414), .B(n413), .Z(n415) );
  XOR U696 ( .A(in[1020]), .B(n415), .Z(n871) );
  XNOR U697 ( .A(n416), .B(n871), .Z(n3595) );
  XNOR U698 ( .A(in[636]), .B(n3595), .Z(n2551) );
  XOR U699 ( .A(in[162]), .B(in[1442]), .Z(n418) );
  XNOR U700 ( .A(in[802]), .B(in[1122]), .Z(n417) );
  XNOR U701 ( .A(n418), .B(n417), .Z(n419) );
  XNOR U702 ( .A(in[482]), .B(n419), .Z(n471) );
  XNOR U703 ( .A(n420), .B(n471), .Z(n3692) );
  XNOR U704 ( .A(in[227]), .B(n3692), .Z(n2844) );
  XOR U705 ( .A(in[1511]), .B(in[551]), .Z(n422) );
  XNOR U706 ( .A(in[871]), .B(in[231]), .Z(n421) );
  XNOR U707 ( .A(n422), .B(n421), .Z(n423) );
  XOR U708 ( .A(in[1191]), .B(n423), .Z(n1313) );
  XNOR U709 ( .A(n424), .B(n1313), .Z(n3733) );
  XNOR U710 ( .A(in[1447]), .B(n3733), .Z(n2841) );
  NAND U711 ( .A(n2844), .B(n2841), .Z(n425) );
  XNOR U712 ( .A(n2551), .B(n425), .Z(out[101]) );
  XOR U713 ( .A(in[1406]), .B(in[126]), .Z(n427) );
  XNOR U714 ( .A(in[1086]), .B(in[766]), .Z(n426) );
  XNOR U715 ( .A(n427), .B(n426), .Z(n428) );
  XOR U716 ( .A(in[446]), .B(n428), .Z(n1469) );
  XOR U717 ( .A(in[1535]), .B(in[575]), .Z(n430) );
  XNOR U718 ( .A(in[895]), .B(in[255]), .Z(n429) );
  XNOR U719 ( .A(n430), .B(n429), .Z(n431) );
  XOR U720 ( .A(in[1215]), .B(n431), .Z(n1024) );
  XNOR U721 ( .A(n1469), .B(n1024), .Z(n3557) );
  XNOR U722 ( .A(in[191]), .B(n3557), .Z(n1383) );
  XOR U723 ( .A(in[1440]), .B(in[480]), .Z(n433) );
  XNOR U724 ( .A(in[800]), .B(in[160]), .Z(n432) );
  XNOR U725 ( .A(n433), .B(n432), .Z(n434) );
  XOR U726 ( .A(in[1120]), .B(n434), .Z(n709) );
  XOR U727 ( .A(in[351]), .B(in[671]), .Z(n436) );
  XNOR U728 ( .A(in[31]), .B(in[1311]), .Z(n435) );
  XNOR U729 ( .A(n436), .B(n435), .Z(n437) );
  XNOR U730 ( .A(in[991]), .B(n437), .Z(n1282) );
  XNOR U731 ( .A(n709), .B(n1282), .Z(n4162) );
  XNOR U732 ( .A(in[1376]), .B(n4162), .Z(n1778) );
  XOR U733 ( .A(in[1064]), .B(in[424]), .Z(n439) );
  XNOR U734 ( .A(in[744]), .B(in[1384]), .Z(n438) );
  XNOR U735 ( .A(n439), .B(n438), .Z(n440) );
  XOR U736 ( .A(in[104]), .B(n440), .Z(n746) );
  XOR U737 ( .A(in[1575]), .B(in[615]), .Z(n442) );
  XNOR U738 ( .A(in[935]), .B(in[295]), .Z(n441) );
  XNOR U739 ( .A(n442), .B(n441), .Z(n443) );
  XOR U740 ( .A(in[1255]), .B(n443), .Z(n799) );
  XNOR U741 ( .A(n746), .B(n799), .Z(n3927) );
  XNOR U742 ( .A(in[1000]), .B(n3927), .Z(n1775) );
  NAND U743 ( .A(n1778), .B(n1775), .Z(n444) );
  XNOR U744 ( .A(n1383), .B(n444), .Z(out[1020]) );
  XOR U745 ( .A(in[1407]), .B(in[127]), .Z(n446) );
  XNOR U746 ( .A(in[1087]), .B(in[767]), .Z(n445) );
  XNOR U747 ( .A(n446), .B(n445), .Z(n447) );
  XOR U748 ( .A(in[447]), .B(n447), .Z(n1472) );
  XOR U749 ( .A(in[1472]), .B(in[512]), .Z(n449) );
  XNOR U750 ( .A(in[832]), .B(in[192]), .Z(n448) );
  XNOR U751 ( .A(n449), .B(n448), .Z(n450) );
  XOR U752 ( .A(in[1152]), .B(n450), .Z(n1091) );
  XNOR U753 ( .A(n1472), .B(n1091), .Z(n3561) );
  XNOR U754 ( .A(in[128]), .B(n3561), .Z(n1387) );
  XOR U755 ( .A(in[352]), .B(in[672]), .Z(n452) );
  XNOR U756 ( .A(in[32]), .B(in[1312]), .Z(n451) );
  XNOR U757 ( .A(n452), .B(n451), .Z(n453) );
  XNOR U758 ( .A(in[992]), .B(n453), .Z(n1285) );
  XNOR U759 ( .A(n454), .B(n1285), .Z(n4165) );
  XNOR U760 ( .A(in[1377]), .B(n4165), .Z(n1782) );
  XOR U761 ( .A(in[1065]), .B(in[425]), .Z(n456) );
  XNOR U762 ( .A(in[745]), .B(in[1385]), .Z(n455) );
  XNOR U763 ( .A(n456), .B(n455), .Z(n457) );
  XOR U764 ( .A(in[105]), .B(n457), .Z(n881) );
  XOR U765 ( .A(in[1576]), .B(in[616]), .Z(n459) );
  XNOR U766 ( .A(in[936]), .B(in[296]), .Z(n458) );
  XNOR U767 ( .A(n459), .B(n458), .Z(n460) );
  XOR U768 ( .A(in[1256]), .B(n460), .Z(n812) );
  XNOR U769 ( .A(n881), .B(n812), .Z(n3929) );
  XNOR U770 ( .A(in[1001]), .B(n3929), .Z(n1779) );
  NAND U771 ( .A(n1782), .B(n1779), .Z(n461) );
  XNOR U772 ( .A(n1387), .B(n461), .Z(out[1021]) );
  XOR U773 ( .A(in[1344]), .B(in[64]), .Z(n463) );
  XNOR U774 ( .A(in[1024]), .B(in[384]), .Z(n462) );
  XNOR U775 ( .A(n463), .B(n462), .Z(n464) );
  XOR U776 ( .A(in[704]), .B(n464), .Z(n1477) );
  XOR U777 ( .A(in[1473]), .B(in[513]), .Z(n466) );
  XNOR U778 ( .A(in[833]), .B(in[193]), .Z(n465) );
  XNOR U779 ( .A(n466), .B(n465), .Z(n467) );
  XOR U780 ( .A(in[1153]), .B(n467), .Z(n1144) );
  XNOR U781 ( .A(n1477), .B(n1144), .Z(n3565) );
  XNOR U782 ( .A(in[129]), .B(n3565), .Z(n1390) );
  XOR U783 ( .A(in[353]), .B(in[673]), .Z(n469) );
  XNOR U784 ( .A(in[33]), .B(in[1313]), .Z(n468) );
  XNOR U785 ( .A(n469), .B(n468), .Z(n470) );
  XOR U786 ( .A(in[993]), .B(n470), .Z(n1288) );
  XNOR U787 ( .A(n1288), .B(n471), .Z(n4168) );
  XNOR U788 ( .A(in[1378]), .B(n4168), .Z(n1786) );
  XOR U789 ( .A(in[1577]), .B(in[617]), .Z(n473) );
  XNOR U790 ( .A(in[937]), .B(in[297]), .Z(n472) );
  XNOR U791 ( .A(n473), .B(n472), .Z(n474) );
  XOR U792 ( .A(in[1257]), .B(n474), .Z(n825) );
  XNOR U793 ( .A(n475), .B(n825), .Z(n3931) );
  XNOR U794 ( .A(in[1002]), .B(n3931), .Z(n1783) );
  NAND U795 ( .A(n1786), .B(n1783), .Z(n476) );
  XNOR U796 ( .A(n1390), .B(n476), .Z(out[1022]) );
  XOR U797 ( .A(n3569), .B(in[130]), .Z(n1392) );
  XOR U798 ( .A(in[163]), .B(in[1443]), .Z(n478) );
  XNOR U799 ( .A(in[803]), .B(in[1123]), .Z(n477) );
  XNOR U800 ( .A(n478), .B(n477), .Z(n479) );
  XOR U801 ( .A(in[483]), .B(n479), .Z(n582) );
  XOR U802 ( .A(in[354]), .B(in[674]), .Z(n481) );
  XNOR U803 ( .A(in[34]), .B(in[1314]), .Z(n480) );
  XNOR U804 ( .A(n481), .B(n480), .Z(n482) );
  XNOR U805 ( .A(in[994]), .B(n482), .Z(n1291) );
  XNOR U806 ( .A(n582), .B(n1291), .Z(n4171) );
  XNOR U807 ( .A(in[1379]), .B(n4171), .Z(n1790) );
  XOR U808 ( .A(in[1578]), .B(in[618]), .Z(n484) );
  XNOR U809 ( .A(in[938]), .B(in[298]), .Z(n483) );
  XNOR U810 ( .A(n484), .B(n483), .Z(n485) );
  XOR U811 ( .A(in[1258]), .B(n485), .Z(n838) );
  XNOR U812 ( .A(n486), .B(n838), .Z(n3933) );
  XNOR U813 ( .A(in[1003]), .B(n3933), .Z(n1787) );
  NAND U814 ( .A(n1790), .B(n1787), .Z(n487) );
  XNOR U815 ( .A(n1392), .B(n487), .Z(out[1023]) );
  XOR U816 ( .A(n489), .B(n488), .Z(n3624) );
  XNOR U817 ( .A(in[531]), .B(n3624), .Z(n1396) );
  XOR U818 ( .A(in[1346]), .B(in[66]), .Z(n491) );
  XNOR U819 ( .A(in[1026]), .B(in[386]), .Z(n490) );
  XNOR U820 ( .A(n491), .B(n490), .Z(n492) );
  XOR U821 ( .A(in[706]), .B(n492), .Z(n1485) );
  XOR U822 ( .A(in[1475]), .B(in[515]), .Z(n494) );
  XNOR U823 ( .A(in[835]), .B(in[195]), .Z(n493) );
  XNOR U824 ( .A(n494), .B(n493), .Z(n495) );
  XNOR U825 ( .A(in[1155]), .B(n495), .Z(n1196) );
  XNOR U826 ( .A(n1485), .B(n1196), .Z(n3573) );
  XNOR U827 ( .A(in[131]), .B(n3573), .Z(n4630) );
  XOR U828 ( .A(in[35]), .B(in[675]), .Z(n497) );
  XNOR U829 ( .A(in[355]), .B(in[1315]), .Z(n496) );
  XNOR U830 ( .A(n497), .B(n496), .Z(n498) );
  XOR U831 ( .A(in[995]), .B(n498), .Z(n1294) );
  XOR U832 ( .A(in[164]), .B(in[1444]), .Z(n500) );
  XNOR U833 ( .A(in[804]), .B(in[1124]), .Z(n499) );
  XNOR U834 ( .A(n500), .B(n499), .Z(n501) );
  XOR U835 ( .A(in[484]), .B(n501), .Z(n741) );
  XNOR U836 ( .A(n1294), .B(n741), .Z(n4174) );
  XNOR U837 ( .A(in[1380]), .B(n4174), .Z(n4627) );
  NAND U838 ( .A(n4630), .B(n4627), .Z(n502) );
  XNOR U839 ( .A(n1396), .B(n502), .Z(out[1024]) );
  XNOR U840 ( .A(n504), .B(n503), .Z(n3628) );
  XNOR U841 ( .A(in[532]), .B(n3628), .Z(n1400) );
  XOR U842 ( .A(in[1347]), .B(in[67]), .Z(n506) );
  XNOR U843 ( .A(in[1027]), .B(in[387]), .Z(n505) );
  XNOR U844 ( .A(n506), .B(n505), .Z(n507) );
  XOR U845 ( .A(in[707]), .B(n507), .Z(n1489) );
  XOR U846 ( .A(in[1476]), .B(in[516]), .Z(n509) );
  XNOR U847 ( .A(in[836]), .B(in[196]), .Z(n508) );
  XNOR U848 ( .A(n509), .B(n508), .Z(n510) );
  XNOR U849 ( .A(in[1156]), .B(n510), .Z(n1199) );
  XNOR U850 ( .A(n1489), .B(n1199), .Z(n3581) );
  XNOR U851 ( .A(in[132]), .B(n3581), .Z(n4634) );
  XOR U852 ( .A(in[1445]), .B(in[165]), .Z(n512) );
  XNOR U853 ( .A(in[805]), .B(in[1125]), .Z(n511) );
  XNOR U854 ( .A(n512), .B(n511), .Z(n513) );
  XOR U855 ( .A(in[485]), .B(n513), .Z(n785) );
  XOR U856 ( .A(in[36]), .B(in[676]), .Z(n515) );
  XNOR U857 ( .A(in[356]), .B(in[1316]), .Z(n514) );
  XNOR U858 ( .A(n515), .B(n514), .Z(n516) );
  XOR U859 ( .A(in[996]), .B(n516), .Z(n1297) );
  XNOR U860 ( .A(n785), .B(n1297), .Z(n4181) );
  XNOR U861 ( .A(in[1381]), .B(n4181), .Z(n4631) );
  NAND U862 ( .A(n4634), .B(n4631), .Z(n517) );
  XNOR U863 ( .A(n1400), .B(n517), .Z(out[1025]) );
  XOR U864 ( .A(n519), .B(n518), .Z(n3632) );
  XNOR U865 ( .A(in[533]), .B(n3632), .Z(n1404) );
  XOR U866 ( .A(in[1348]), .B(in[68]), .Z(n521) );
  XNOR U867 ( .A(in[1028]), .B(in[388]), .Z(n520) );
  XNOR U868 ( .A(n521), .B(n520), .Z(n522) );
  XOR U869 ( .A(in[708]), .B(n522), .Z(n1493) );
  XOR U870 ( .A(in[1477]), .B(in[517]), .Z(n524) );
  XNOR U871 ( .A(in[837]), .B(in[197]), .Z(n523) );
  XNOR U872 ( .A(n524), .B(n523), .Z(n525) );
  XNOR U873 ( .A(in[1157]), .B(n525), .Z(n1202) );
  XNOR U874 ( .A(n1493), .B(n1202), .Z(n3585) );
  XNOR U875 ( .A(in[133]), .B(n3585), .Z(n4638) );
  XOR U876 ( .A(in[37]), .B(in[677]), .Z(n527) );
  XNOR U877 ( .A(in[357]), .B(in[1317]), .Z(n526) );
  XNOR U878 ( .A(n527), .B(n526), .Z(n528) );
  XOR U879 ( .A(in[997]), .B(n528), .Z(n1300) );
  XOR U880 ( .A(in[166]), .B(in[806]), .Z(n530) );
  XNOR U881 ( .A(in[1126]), .B(in[486]), .Z(n529) );
  XNOR U882 ( .A(n530), .B(n529), .Z(n531) );
  XOR U883 ( .A(in[1446]), .B(n531), .Z(n798) );
  XNOR U884 ( .A(n1300), .B(n798), .Z(n4184) );
  XNOR U885 ( .A(in[1382]), .B(n4184), .Z(n4635) );
  NAND U886 ( .A(n4638), .B(n4635), .Z(n532) );
  XNOR U887 ( .A(n1404), .B(n532), .Z(out[1026]) );
  XOR U888 ( .A(n534), .B(n533), .Z(n3636) );
  XNOR U889 ( .A(in[534]), .B(n3636), .Z(n1408) );
  XOR U890 ( .A(in[1349]), .B(in[69]), .Z(n536) );
  XNOR U891 ( .A(in[1029]), .B(in[389]), .Z(n535) );
  XNOR U892 ( .A(n536), .B(n535), .Z(n537) );
  XOR U893 ( .A(in[709]), .B(n537), .Z(n1497) );
  XOR U894 ( .A(in[1478]), .B(in[518]), .Z(n539) );
  XNOR U895 ( .A(in[838]), .B(in[198]), .Z(n538) );
  XNOR U896 ( .A(n539), .B(n538), .Z(n540) );
  XNOR U897 ( .A(in[1158]), .B(n540), .Z(n1205) );
  XNOR U898 ( .A(n1497), .B(n1205), .Z(n3589) );
  XNOR U899 ( .A(in[134]), .B(n3589), .Z(n4642) );
  XOR U900 ( .A(in[167]), .B(in[807]), .Z(n542) );
  XNOR U901 ( .A(in[1127]), .B(in[487]), .Z(n541) );
  XNOR U902 ( .A(n542), .B(n541), .Z(n543) );
  XOR U903 ( .A(in[1447]), .B(n543), .Z(n811) );
  XOR U904 ( .A(in[38]), .B(in[678]), .Z(n545) );
  XNOR U905 ( .A(in[358]), .B(in[1318]), .Z(n544) );
  XNOR U906 ( .A(n545), .B(n544), .Z(n546) );
  XOR U907 ( .A(in[998]), .B(n546), .Z(n1304) );
  XNOR U908 ( .A(n811), .B(n1304), .Z(n3963) );
  XNOR U909 ( .A(in[1383]), .B(n3963), .Z(n4639) );
  NAND U910 ( .A(n4642), .B(n4639), .Z(n547) );
  XNOR U911 ( .A(n1408), .B(n547), .Z(out[1027]) );
  XOR U912 ( .A(n549), .B(n548), .Z(n3640) );
  XNOR U913 ( .A(in[535]), .B(n3640), .Z(n1412) );
  XOR U914 ( .A(in[1350]), .B(in[70]), .Z(n551) );
  XNOR U915 ( .A(in[1030]), .B(in[390]), .Z(n550) );
  XNOR U916 ( .A(n551), .B(n550), .Z(n552) );
  XOR U917 ( .A(in[710]), .B(n552), .Z(n1501) );
  XOR U918 ( .A(in[199]), .B(in[1479]), .Z(n554) );
  XNOR U919 ( .A(in[1159]), .B(in[839]), .Z(n553) );
  XNOR U920 ( .A(n554), .B(n553), .Z(n555) );
  XNOR U921 ( .A(in[519]), .B(n555), .Z(n1208) );
  XNOR U922 ( .A(n1501), .B(n1208), .Z(n3593) );
  XNOR U923 ( .A(in[135]), .B(n3593), .Z(n4646) );
  XOR U924 ( .A(in[39]), .B(in[679]), .Z(n557) );
  XNOR U925 ( .A(in[359]), .B(in[1319]), .Z(n556) );
  XNOR U926 ( .A(n557), .B(n556), .Z(n558) );
  XOR U927 ( .A(in[999]), .B(n558), .Z(n1308) );
  XOR U928 ( .A(in[168]), .B(in[1448]), .Z(n560) );
  XNOR U929 ( .A(in[1128]), .B(in[808]), .Z(n559) );
  XNOR U930 ( .A(n560), .B(n559), .Z(n561) );
  XOR U931 ( .A(in[488]), .B(n561), .Z(n824) );
  XNOR U932 ( .A(n1308), .B(n824), .Z(n3966) );
  XNOR U933 ( .A(in[1384]), .B(n3966), .Z(n4643) );
  NAND U934 ( .A(n4646), .B(n4643), .Z(n562) );
  XNOR U935 ( .A(n1412), .B(n562), .Z(out[1028]) );
  XOR U936 ( .A(n564), .B(n563), .Z(n3644) );
  XNOR U937 ( .A(in[536]), .B(n3644), .Z(n1416) );
  XOR U938 ( .A(in[1351]), .B(in[711]), .Z(n566) );
  XNOR U939 ( .A(in[1031]), .B(in[391]), .Z(n565) );
  XNOR U940 ( .A(n566), .B(n565), .Z(n567) );
  XOR U941 ( .A(in[71]), .B(n567), .Z(n1505) );
  XOR U942 ( .A(in[1480]), .B(in[520]), .Z(n569) );
  XNOR U943 ( .A(in[840]), .B(in[200]), .Z(n568) );
  XNOR U944 ( .A(n569), .B(n568), .Z(n570) );
  XNOR U945 ( .A(in[1160]), .B(n570), .Z(n1213) );
  XNOR U946 ( .A(n1505), .B(n1213), .Z(n3597) );
  XNOR U947 ( .A(in[136]), .B(n3597), .Z(n4650) );
  XOR U948 ( .A(in[169]), .B(in[1449]), .Z(n572) );
  XNOR U949 ( .A(in[1129]), .B(in[809]), .Z(n571) );
  XNOR U950 ( .A(n572), .B(n571), .Z(n573) );
  XOR U951 ( .A(in[489]), .B(n573), .Z(n837) );
  XOR U952 ( .A(in[680]), .B(in[1320]), .Z(n575) );
  XNOR U953 ( .A(in[40]), .B(in[360]), .Z(n574) );
  XNOR U954 ( .A(n575), .B(n574), .Z(n576) );
  XOR U955 ( .A(in[1000]), .B(n576), .Z(n1312) );
  XNOR U956 ( .A(n837), .B(n1312), .Z(n3973) );
  XNOR U957 ( .A(in[1385]), .B(n3973), .Z(n4647) );
  NAND U958 ( .A(n4650), .B(n4647), .Z(n577) );
  XNOR U959 ( .A(n1416), .B(n577), .Z(out[1029]) );
  XOR U960 ( .A(in[1341]), .B(in[61]), .Z(n579) );
  XNOR U961 ( .A(in[701]), .B(in[381]), .Z(n578) );
  XNOR U962 ( .A(n579), .B(n578), .Z(n580) );
  XOR U963 ( .A(in[1021]), .B(n580), .Z(n894) );
  XNOR U964 ( .A(n581), .B(n894), .Z(n3599) );
  XNOR U965 ( .A(in[637]), .B(n3599), .Z(n2554) );
  XOR U966 ( .A(n583), .B(n582), .Z(n3696) );
  XNOR U967 ( .A(in[228]), .B(n3696), .Z(n2858) );
  XOR U968 ( .A(in[1512]), .B(in[552]), .Z(n585) );
  XNOR U969 ( .A(in[872]), .B(in[232]), .Z(n584) );
  XNOR U970 ( .A(n585), .B(n584), .Z(n586) );
  XOR U971 ( .A(in[1192]), .B(n586), .Z(n1317) );
  XNOR U972 ( .A(n587), .B(n1317), .Z(n3737) );
  XNOR U973 ( .A(in[1448]), .B(n3737), .Z(n2855) );
  NAND U974 ( .A(n2858), .B(n2855), .Z(n588) );
  XNOR U975 ( .A(n2554), .B(n588), .Z(out[102]) );
  XNOR U976 ( .A(n590), .B(n589), .Z(n3648) );
  XNOR U977 ( .A(in[537]), .B(n3648), .Z(n1420) );
  XOR U978 ( .A(in[1352]), .B(in[712]), .Z(n592) );
  XNOR U979 ( .A(in[1032]), .B(in[392]), .Z(n591) );
  XNOR U980 ( .A(n592), .B(n591), .Z(n593) );
  XOR U981 ( .A(in[72]), .B(n593), .Z(n1510) );
  XOR U982 ( .A(in[1481]), .B(in[521]), .Z(n595) );
  XNOR U983 ( .A(in[841]), .B(in[201]), .Z(n594) );
  XNOR U984 ( .A(n595), .B(n594), .Z(n596) );
  XNOR U985 ( .A(in[1161]), .B(n596), .Z(n1216) );
  XNOR U986 ( .A(n1510), .B(n1216), .Z(n3601) );
  XNOR U987 ( .A(in[137]), .B(n3601), .Z(n4654) );
  XOR U988 ( .A(in[170]), .B(in[1450]), .Z(n598) );
  XNOR U989 ( .A(in[1130]), .B(in[810]), .Z(n597) );
  XNOR U990 ( .A(n598), .B(n597), .Z(n599) );
  XOR U991 ( .A(in[490]), .B(n599), .Z(n853) );
  XOR U992 ( .A(in[681]), .B(in[1321]), .Z(n601) );
  XNOR U993 ( .A(in[41]), .B(in[361]), .Z(n600) );
  XNOR U994 ( .A(n601), .B(n600), .Z(n602) );
  XOR U995 ( .A(in[1001]), .B(n602), .Z(n1316) );
  XNOR U996 ( .A(n853), .B(n1316), .Z(n3976) );
  XNOR U997 ( .A(in[1386]), .B(n3976), .Z(n4651) );
  NAND U998 ( .A(n4654), .B(n4651), .Z(n603) );
  XNOR U999 ( .A(n1420), .B(n603), .Z(out[1030]) );
  XNOR U1000 ( .A(n605), .B(n604), .Z(n3652) );
  XNOR U1001 ( .A(in[538]), .B(n3652), .Z(n1424) );
  XOR U1002 ( .A(in[1353]), .B(in[393]), .Z(n607) );
  XNOR U1003 ( .A(in[713]), .B(in[73]), .Z(n606) );
  XNOR U1004 ( .A(n607), .B(n606), .Z(n608) );
  XOR U1005 ( .A(in[1033]), .B(n608), .Z(n1514) );
  XOR U1006 ( .A(in[1482]), .B(in[522]), .Z(n610) );
  XNOR U1007 ( .A(in[842]), .B(in[202]), .Z(n609) );
  XNOR U1008 ( .A(n610), .B(n609), .Z(n611) );
  XNOR U1009 ( .A(in[1162]), .B(n611), .Z(n1219) );
  XNOR U1010 ( .A(n1514), .B(n1219), .Z(n3605) );
  XNOR U1011 ( .A(in[138]), .B(n3605), .Z(n4658) );
  XOR U1012 ( .A(in[682]), .B(in[1322]), .Z(n613) );
  XNOR U1013 ( .A(in[42]), .B(in[362]), .Z(n612) );
  XNOR U1014 ( .A(n613), .B(n612), .Z(n614) );
  XOR U1015 ( .A(in[1002]), .B(n614), .Z(n1321) );
  XOR U1016 ( .A(in[811]), .B(in[491]), .Z(n616) );
  XNOR U1017 ( .A(in[1451]), .B(in[1131]), .Z(n615) );
  XNOR U1018 ( .A(n616), .B(n615), .Z(n617) );
  XOR U1019 ( .A(in[171]), .B(n617), .Z(n866) );
  XNOR U1020 ( .A(n1321), .B(n866), .Z(n3979) );
  XNOR U1021 ( .A(in[1387]), .B(n3979), .Z(n4655) );
  NAND U1022 ( .A(n4658), .B(n4655), .Z(n618) );
  XNOR U1023 ( .A(n1424), .B(n618), .Z(out[1031]) );
  XOR U1024 ( .A(n620), .B(n619), .Z(n3656) );
  XNOR U1025 ( .A(in[539]), .B(n3656), .Z(n1429) );
  XOR U1026 ( .A(in[1354]), .B(in[714]), .Z(n622) );
  XNOR U1027 ( .A(in[74]), .B(in[394]), .Z(n621) );
  XNOR U1028 ( .A(n622), .B(n621), .Z(n623) );
  XOR U1029 ( .A(in[1034]), .B(n623), .Z(n1518) );
  XOR U1030 ( .A(in[1483]), .B(in[523]), .Z(n625) );
  XNOR U1031 ( .A(in[843]), .B(in[203]), .Z(n624) );
  XNOR U1032 ( .A(n625), .B(n624), .Z(n626) );
  XNOR U1033 ( .A(in[1163]), .B(n626), .Z(n1222) );
  XNOR U1034 ( .A(n1518), .B(n1222), .Z(n3609) );
  XNOR U1035 ( .A(n3609), .B(in[139]), .Z(n4662) );
  XOR U1036 ( .A(in[812]), .B(in[492]), .Z(n628) );
  XNOR U1037 ( .A(in[1452]), .B(in[1132]), .Z(n627) );
  XNOR U1038 ( .A(n628), .B(n627), .Z(n629) );
  XOR U1039 ( .A(in[172]), .B(n629), .Z(n886) );
  XOR U1040 ( .A(in[683]), .B(in[1323]), .Z(n631) );
  XNOR U1041 ( .A(in[43]), .B(in[363]), .Z(n630) );
  XNOR U1042 ( .A(n631), .B(n630), .Z(n632) );
  XOR U1043 ( .A(in[1003]), .B(n632), .Z(n1325) );
  XNOR U1044 ( .A(n886), .B(n1325), .Z(n3982) );
  XNOR U1045 ( .A(in[1388]), .B(n3982), .Z(n4659) );
  NAND U1046 ( .A(n4662), .B(n4659), .Z(n633) );
  XNOR U1047 ( .A(n1429), .B(n633), .Z(out[1032]) );
  XNOR U1048 ( .A(n635), .B(n634), .Z(n3660) );
  XNOR U1049 ( .A(in[540]), .B(n3660), .Z(n1433) );
  XOR U1050 ( .A(in[1355]), .B(in[715]), .Z(n637) );
  XNOR U1051 ( .A(in[1035]), .B(in[395]), .Z(n636) );
  XNOR U1052 ( .A(n637), .B(n636), .Z(n638) );
  XOR U1053 ( .A(in[75]), .B(n638), .Z(n1522) );
  XOR U1054 ( .A(in[1484]), .B(in[524]), .Z(n640) );
  XNOR U1055 ( .A(in[844]), .B(in[204]), .Z(n639) );
  XNOR U1056 ( .A(n640), .B(n639), .Z(n641) );
  XNOR U1057 ( .A(in[1164]), .B(n641), .Z(n1225) );
  XNOR U1058 ( .A(n1522), .B(n1225), .Z(n3613) );
  XNOR U1059 ( .A(in[140]), .B(n3613), .Z(n4666) );
  XOR U1060 ( .A(in[813]), .B(in[493]), .Z(n643) );
  XNOR U1061 ( .A(in[1453]), .B(in[1133]), .Z(n642) );
  XNOR U1062 ( .A(n643), .B(n642), .Z(n644) );
  XOR U1063 ( .A(in[173]), .B(n644), .Z(n899) );
  XOR U1064 ( .A(in[1324]), .B(in[44]), .Z(n646) );
  XNOR U1065 ( .A(in[684]), .B(in[364]), .Z(n645) );
  XNOR U1066 ( .A(n646), .B(n645), .Z(n647) );
  XOR U1067 ( .A(in[1004]), .B(n647), .Z(n1328) );
  XNOR U1068 ( .A(n899), .B(n1328), .Z(n3985) );
  XNOR U1069 ( .A(in[1389]), .B(n3985), .Z(n4663) );
  NAND U1070 ( .A(n4666), .B(n4663), .Z(n648) );
  XNOR U1071 ( .A(n1433), .B(n648), .Z(out[1033]) );
  XNOR U1072 ( .A(n650), .B(n649), .Z(n3668) );
  XNOR U1073 ( .A(in[541]), .B(n3668), .Z(n1437) );
  XOR U1074 ( .A(in[76]), .B(in[1036]), .Z(n652) );
  XNOR U1075 ( .A(in[716]), .B(in[396]), .Z(n651) );
  XNOR U1076 ( .A(n652), .B(n651), .Z(n653) );
  XOR U1077 ( .A(in[1356]), .B(n653), .Z(n1526) );
  XOR U1078 ( .A(in[1485]), .B(in[525]), .Z(n655) );
  XNOR U1079 ( .A(in[845]), .B(in[205]), .Z(n654) );
  XNOR U1080 ( .A(n655), .B(n654), .Z(n656) );
  XNOR U1081 ( .A(in[1165]), .B(n656), .Z(n1228) );
  XNOR U1082 ( .A(n1526), .B(n1228), .Z(n3617) );
  XNOR U1083 ( .A(in[141]), .B(n3617), .Z(n4674) );
  XOR U1084 ( .A(in[814]), .B(in[494]), .Z(n658) );
  XNOR U1085 ( .A(in[1454]), .B(in[1134]), .Z(n657) );
  XNOR U1086 ( .A(n658), .B(n657), .Z(n659) );
  XOR U1087 ( .A(in[174]), .B(n659), .Z(n912) );
  XOR U1088 ( .A(in[1325]), .B(in[45]), .Z(n661) );
  XNOR U1089 ( .A(in[685]), .B(in[365]), .Z(n660) );
  XNOR U1090 ( .A(n661), .B(n660), .Z(n662) );
  XOR U1091 ( .A(in[1005]), .B(n662), .Z(n1332) );
  XNOR U1092 ( .A(n912), .B(n1332), .Z(n3988) );
  XNOR U1093 ( .A(in[1390]), .B(n3988), .Z(n4671) );
  NAND U1094 ( .A(n4674), .B(n4671), .Z(n663) );
  XNOR U1095 ( .A(n1437), .B(n663), .Z(out[1034]) );
  XNOR U1096 ( .A(n665), .B(n664), .Z(n3672) );
  XNOR U1097 ( .A(in[542]), .B(n3672), .Z(n1441) );
  XOR U1098 ( .A(in[77]), .B(in[1037]), .Z(n667) );
  XNOR U1099 ( .A(in[717]), .B(in[397]), .Z(n666) );
  XNOR U1100 ( .A(n667), .B(n666), .Z(n668) );
  XOR U1101 ( .A(in[1357]), .B(n668), .Z(n1530) );
  XOR U1102 ( .A(in[1486]), .B(in[526]), .Z(n670) );
  XNOR U1103 ( .A(in[846]), .B(in[206]), .Z(n669) );
  XNOR U1104 ( .A(n670), .B(n669), .Z(n671) );
  XNOR U1105 ( .A(in[1166]), .B(n671), .Z(n1231) );
  XNOR U1106 ( .A(n1530), .B(n1231), .Z(n3625) );
  XNOR U1107 ( .A(in[142]), .B(n3625), .Z(n4678) );
  XOR U1108 ( .A(in[815]), .B(in[495]), .Z(n673) );
  XNOR U1109 ( .A(in[1455]), .B(in[1135]), .Z(n672) );
  XNOR U1110 ( .A(n673), .B(n672), .Z(n674) );
  XOR U1111 ( .A(in[175]), .B(n674), .Z(n925) );
  XOR U1112 ( .A(in[1326]), .B(in[46]), .Z(n676) );
  XNOR U1113 ( .A(in[686]), .B(in[366]), .Z(n675) );
  XNOR U1114 ( .A(n676), .B(n675), .Z(n677) );
  XOR U1115 ( .A(in[1006]), .B(n677), .Z(n1336) );
  XNOR U1116 ( .A(n925), .B(n1336), .Z(n3991) );
  XNOR U1117 ( .A(in[1391]), .B(n3991), .Z(n4675) );
  NAND U1118 ( .A(n4678), .B(n4675), .Z(n678) );
  XNOR U1119 ( .A(n1441), .B(n678), .Z(out[1035]) );
  XNOR U1120 ( .A(n680), .B(n679), .Z(n3676) );
  XNOR U1121 ( .A(in[543]), .B(n3676), .Z(n1445) );
  XOR U1122 ( .A(in[78]), .B(in[1038]), .Z(n682) );
  XNOR U1123 ( .A(in[718]), .B(in[398]), .Z(n681) );
  XNOR U1124 ( .A(n682), .B(n681), .Z(n683) );
  XOR U1125 ( .A(in[1358]), .B(n683), .Z(n1534) );
  XOR U1126 ( .A(in[1487]), .B(in[527]), .Z(n685) );
  XNOR U1127 ( .A(in[847]), .B(in[207]), .Z(n684) );
  XNOR U1128 ( .A(n685), .B(n684), .Z(n686) );
  XNOR U1129 ( .A(in[1167]), .B(n686), .Z(n1234) );
  XNOR U1130 ( .A(n1534), .B(n1234), .Z(n3629) );
  XNOR U1131 ( .A(in[143]), .B(n3629), .Z(n4682) );
  XOR U1132 ( .A(in[1327]), .B(in[47]), .Z(n688) );
  XNOR U1133 ( .A(in[687]), .B(in[367]), .Z(n687) );
  XNOR U1134 ( .A(n688), .B(n687), .Z(n689) );
  XOR U1135 ( .A(in[1007]), .B(n689), .Z(n1340) );
  XOR U1136 ( .A(in[816]), .B(in[496]), .Z(n691) );
  XNOR U1137 ( .A(in[1456]), .B(in[1136]), .Z(n690) );
  XNOR U1138 ( .A(n691), .B(n690), .Z(n692) );
  XOR U1139 ( .A(in[176]), .B(n692), .Z(n940) );
  XNOR U1140 ( .A(n1340), .B(n940), .Z(n3994) );
  XNOR U1141 ( .A(in[1392]), .B(n3994), .Z(n4679) );
  NAND U1142 ( .A(n4682), .B(n4679), .Z(n693) );
  XNOR U1143 ( .A(n1445), .B(n693), .Z(out[1036]) );
  XNOR U1144 ( .A(n695), .B(n694), .Z(n3680) );
  XNOR U1145 ( .A(in[544]), .B(n3680), .Z(n1449) );
  XOR U1146 ( .A(in[79]), .B(in[1039]), .Z(n697) );
  XNOR U1147 ( .A(in[719]), .B(in[399]), .Z(n696) );
  XNOR U1148 ( .A(n697), .B(n696), .Z(n698) );
  XOR U1149 ( .A(in[1359]), .B(n698), .Z(n1538) );
  XOR U1150 ( .A(in[1488]), .B(in[528]), .Z(n700) );
  XNOR U1151 ( .A(in[848]), .B(in[208]), .Z(n699) );
  XNOR U1152 ( .A(n700), .B(n699), .Z(n701) );
  XNOR U1153 ( .A(in[1168]), .B(n701), .Z(n1237) );
  XNOR U1154 ( .A(n1538), .B(n1237), .Z(n3633) );
  XNOR U1155 ( .A(in[144]), .B(n3633), .Z(n4686) );
  XOR U1156 ( .A(in[1328]), .B(in[48]), .Z(n703) );
  XNOR U1157 ( .A(in[688]), .B(in[368]), .Z(n702) );
  XNOR U1158 ( .A(n703), .B(n702), .Z(n704) );
  XOR U1159 ( .A(in[1008]), .B(n704), .Z(n1344) );
  XOR U1160 ( .A(in[817]), .B(in[497]), .Z(n706) );
  XNOR U1161 ( .A(in[1457]), .B(in[1137]), .Z(n705) );
  XNOR U1162 ( .A(n706), .B(n705), .Z(n707) );
  XOR U1163 ( .A(in[177]), .B(n707), .Z(n955) );
  XNOR U1164 ( .A(n1344), .B(n955), .Z(n3997) );
  XNOR U1165 ( .A(in[1393]), .B(n3997), .Z(n4683) );
  NAND U1166 ( .A(n4686), .B(n4683), .Z(n708) );
  XNOR U1167 ( .A(n1449), .B(n708), .Z(out[1037]) );
  XNOR U1168 ( .A(n710), .B(n709), .Z(n3684) );
  XNOR U1169 ( .A(in[545]), .B(n3684), .Z(n1453) );
  XOR U1170 ( .A(in[80]), .B(in[1040]), .Z(n712) );
  XNOR U1171 ( .A(in[720]), .B(in[400]), .Z(n711) );
  XNOR U1172 ( .A(n712), .B(n711), .Z(n713) );
  XOR U1173 ( .A(in[1360]), .B(n713), .Z(n1542) );
  XOR U1174 ( .A(in[1489]), .B(in[529]), .Z(n715) );
  XNOR U1175 ( .A(in[849]), .B(in[209]), .Z(n714) );
  XNOR U1176 ( .A(n715), .B(n714), .Z(n716) );
  XNOR U1177 ( .A(in[1169]), .B(n716), .Z(n1240) );
  XNOR U1178 ( .A(n1542), .B(n1240), .Z(n3637) );
  XNOR U1179 ( .A(in[145]), .B(n3637), .Z(n4690) );
  XOR U1180 ( .A(in[818]), .B(in[498]), .Z(n718) );
  XNOR U1181 ( .A(in[1458]), .B(in[1138]), .Z(n717) );
  XNOR U1182 ( .A(n718), .B(n717), .Z(n719) );
  XOR U1183 ( .A(in[178]), .B(n719), .Z(n970) );
  XOR U1184 ( .A(in[1329]), .B(in[49]), .Z(n721) );
  XNOR U1185 ( .A(in[689]), .B(in[369]), .Z(n720) );
  XNOR U1186 ( .A(n721), .B(n720), .Z(n722) );
  XOR U1187 ( .A(in[1009]), .B(n722), .Z(n1349) );
  XNOR U1188 ( .A(n970), .B(n1349), .Z(n4000) );
  XNOR U1189 ( .A(in[1394]), .B(n4000), .Z(n4687) );
  NAND U1190 ( .A(n4690), .B(n4687), .Z(n723) );
  XNOR U1191 ( .A(n1453), .B(n723), .Z(out[1038]) );
  XOR U1192 ( .A(n3688), .B(in[546]), .Z(n1457) );
  XOR U1193 ( .A(in[81]), .B(in[1041]), .Z(n725) );
  XNOR U1194 ( .A(in[721]), .B(in[401]), .Z(n724) );
  XNOR U1195 ( .A(n725), .B(n724), .Z(n726) );
  XOR U1196 ( .A(in[1361]), .B(n726), .Z(n1546) );
  XOR U1197 ( .A(in[1490]), .B(in[530]), .Z(n728) );
  XNOR U1198 ( .A(in[850]), .B(in[210]), .Z(n727) );
  XNOR U1199 ( .A(n728), .B(n727), .Z(n729) );
  XNOR U1200 ( .A(in[1170]), .B(n729), .Z(n1244) );
  XNOR U1201 ( .A(n1546), .B(n1244), .Z(n3641) );
  XNOR U1202 ( .A(in[146]), .B(n3641), .Z(n4694) );
  XOR U1203 ( .A(in[1330]), .B(in[50]), .Z(n731) );
  XNOR U1204 ( .A(in[690]), .B(in[370]), .Z(n730) );
  XNOR U1205 ( .A(n731), .B(n730), .Z(n732) );
  XOR U1206 ( .A(in[1010]), .B(n732), .Z(n1353) );
  XOR U1207 ( .A(in[819]), .B(in[499]), .Z(n734) );
  XNOR U1208 ( .A(in[1459]), .B(in[1139]), .Z(n733) );
  XNOR U1209 ( .A(n734), .B(n733), .Z(n735) );
  XOR U1210 ( .A(in[179]), .B(n735), .Z(n985) );
  XNOR U1211 ( .A(n1353), .B(n985), .Z(n4007) );
  XNOR U1212 ( .A(in[1395]), .B(n4007), .Z(n4691) );
  NAND U1213 ( .A(n4694), .B(n4691), .Z(n736) );
  XNOR U1214 ( .A(n1457), .B(n736), .Z(out[1039]) );
  XOR U1215 ( .A(in[1342]), .B(in[62]), .Z(n738) );
  XNOR U1216 ( .A(in[702]), .B(in[382]), .Z(n737) );
  XNOR U1217 ( .A(n738), .B(n737), .Z(n739) );
  XOR U1218 ( .A(in[1022]), .B(n739), .Z(n907) );
  XNOR U1219 ( .A(n740), .B(n907), .Z(n3603) );
  XNOR U1220 ( .A(in[638]), .B(n3603), .Z(n2556) );
  XOR U1221 ( .A(n742), .B(n741), .Z(n3700) );
  XNOR U1222 ( .A(in[229]), .B(n3700), .Z(n2872) );
  XOR U1223 ( .A(in[1513]), .B(in[553]), .Z(n744) );
  XNOR U1224 ( .A(in[873]), .B(in[233]), .Z(n743) );
  XNOR U1225 ( .A(n744), .B(n743), .Z(n745) );
  XOR U1226 ( .A(in[1193]), .B(n745), .Z(n1320) );
  XNOR U1227 ( .A(n746), .B(n1320), .Z(n3741) );
  XNOR U1228 ( .A(in[1449]), .B(n3741), .Z(n2869) );
  NAND U1229 ( .A(n2872), .B(n2869), .Z(n747) );
  XNOR U1230 ( .A(n2556), .B(n747), .Z(out[103]) );
  XOR U1231 ( .A(n3692), .B(in[547]), .Z(n1461) );
  XOR U1232 ( .A(in[1042]), .B(in[402]), .Z(n749) );
  XNOR U1233 ( .A(in[722]), .B(in[82]), .Z(n748) );
  XNOR U1234 ( .A(n749), .B(n748), .Z(n750) );
  XOR U1235 ( .A(in[1362]), .B(n750), .Z(n1551) );
  XOR U1236 ( .A(in[851]), .B(in[1171]), .Z(n752) );
  XNOR U1237 ( .A(in[1491]), .B(in[211]), .Z(n751) );
  XNOR U1238 ( .A(n752), .B(n751), .Z(n753) );
  XNOR U1239 ( .A(in[531]), .B(n753), .Z(n1247) );
  XNOR U1240 ( .A(n1551), .B(n1247), .Z(n3645) );
  XNOR U1241 ( .A(in[147]), .B(n3645), .Z(n4698) );
  XOR U1242 ( .A(in[820]), .B(in[500]), .Z(n755) );
  XNOR U1243 ( .A(in[1460]), .B(in[1140]), .Z(n754) );
  XNOR U1244 ( .A(n755), .B(n754), .Z(n756) );
  XOR U1245 ( .A(in[180]), .B(n756), .Z(n1000) );
  XOR U1246 ( .A(in[1331]), .B(in[51]), .Z(n758) );
  XNOR U1247 ( .A(in[691]), .B(in[371]), .Z(n757) );
  XNOR U1248 ( .A(n758), .B(n757), .Z(n759) );
  XOR U1249 ( .A(in[1011]), .B(n759), .Z(n1357) );
  XNOR U1250 ( .A(n1000), .B(n1357), .Z(n4010) );
  XNOR U1251 ( .A(in[1396]), .B(n4010), .Z(n4695) );
  NAND U1252 ( .A(n4698), .B(n4695), .Z(n760) );
  XNOR U1253 ( .A(n1461), .B(n760), .Z(out[1040]) );
  XOR U1254 ( .A(n3696), .B(in[548]), .Z(n1465) );
  XOR U1255 ( .A(in[83]), .B(in[1043]), .Z(n762) );
  XNOR U1256 ( .A(in[723]), .B(in[403]), .Z(n761) );
  XNOR U1257 ( .A(n762), .B(n761), .Z(n763) );
  XOR U1258 ( .A(in[1363]), .B(n763), .Z(n1555) );
  XOR U1259 ( .A(in[852]), .B(in[1172]), .Z(n765) );
  XNOR U1260 ( .A(in[1492]), .B(in[212]), .Z(n764) );
  XNOR U1261 ( .A(n765), .B(n764), .Z(n766) );
  XNOR U1262 ( .A(in[532]), .B(n766), .Z(n1250) );
  XNOR U1263 ( .A(n1555), .B(n1250), .Z(n3649) );
  XNOR U1264 ( .A(in[148]), .B(n3649), .Z(n4702) );
  XOR U1265 ( .A(in[821]), .B(in[501]), .Z(n768) );
  XNOR U1266 ( .A(in[1461]), .B(in[1141]), .Z(n767) );
  XNOR U1267 ( .A(n768), .B(n767), .Z(n769) );
  XOR U1268 ( .A(in[181]), .B(n769), .Z(n1015) );
  XOR U1269 ( .A(in[1332]), .B(in[52]), .Z(n771) );
  XNOR U1270 ( .A(in[692]), .B(in[372]), .Z(n770) );
  XNOR U1271 ( .A(n771), .B(n770), .Z(n772) );
  XOR U1272 ( .A(in[1012]), .B(n772), .Z(n1361) );
  XNOR U1273 ( .A(n1015), .B(n1361), .Z(n4013) );
  XNOR U1274 ( .A(in[1397]), .B(n4013), .Z(n4699) );
  NAND U1275 ( .A(n4702), .B(n4699), .Z(n773) );
  XNOR U1276 ( .A(n1465), .B(n773), .Z(out[1041]) );
  XOR U1277 ( .A(n3700), .B(in[549]), .Z(n1470) );
  XOR U1278 ( .A(in[853]), .B(in[1173]), .Z(n775) );
  XNOR U1279 ( .A(in[1493]), .B(in[213]), .Z(n774) );
  XNOR U1280 ( .A(n775), .B(n774), .Z(n776) );
  XNOR U1281 ( .A(in[533]), .B(n776), .Z(n1253) );
  XNOR U1282 ( .A(n777), .B(n1253), .Z(n3653) );
  XNOR U1283 ( .A(in[149]), .B(n3653), .Z(n4706) );
  XOR U1284 ( .A(in[822]), .B(in[502]), .Z(n779) );
  XNOR U1285 ( .A(in[1462]), .B(in[1142]), .Z(n778) );
  XNOR U1286 ( .A(n779), .B(n778), .Z(n780) );
  XOR U1287 ( .A(in[182]), .B(n780), .Z(n1029) );
  XOR U1288 ( .A(in[1333]), .B(in[53]), .Z(n782) );
  XNOR U1289 ( .A(in[693]), .B(in[373]), .Z(n781) );
  XNOR U1290 ( .A(n782), .B(n781), .Z(n783) );
  XOR U1291 ( .A(in[1013]), .B(n783), .Z(n1365) );
  XNOR U1292 ( .A(n1029), .B(n1365), .Z(n4016) );
  XNOR U1293 ( .A(in[1398]), .B(n4016), .Z(n4703) );
  NAND U1294 ( .A(n4706), .B(n4703), .Z(n784) );
  XNOR U1295 ( .A(n1470), .B(n784), .Z(out[1042]) );
  XNOR U1296 ( .A(n786), .B(n785), .Z(n3704) );
  XNOR U1297 ( .A(in[550]), .B(n3704), .Z(n1474) );
  XOR U1298 ( .A(in[854]), .B(in[1174]), .Z(n788) );
  XNOR U1299 ( .A(in[1494]), .B(in[214]), .Z(n787) );
  XNOR U1300 ( .A(n788), .B(n787), .Z(n789) );
  XNOR U1301 ( .A(in[534]), .B(n789), .Z(n1256) );
  XNOR U1302 ( .A(n790), .B(n1256), .Z(n3657) );
  XNOR U1303 ( .A(in[150]), .B(n3657), .Z(n4710) );
  XOR U1304 ( .A(in[823]), .B(in[503]), .Z(n792) );
  XNOR U1305 ( .A(in[1463]), .B(in[1143]), .Z(n791) );
  XNOR U1306 ( .A(n792), .B(n791), .Z(n793) );
  XOR U1307 ( .A(in[183]), .B(n793), .Z(n1040) );
  XOR U1308 ( .A(in[1334]), .B(in[54]), .Z(n795) );
  XNOR U1309 ( .A(in[694]), .B(in[374]), .Z(n794) );
  XNOR U1310 ( .A(n795), .B(n794), .Z(n796) );
  XOR U1311 ( .A(in[1014]), .B(n796), .Z(n1369) );
  XNOR U1312 ( .A(n1040), .B(n1369), .Z(n4019) );
  XNOR U1313 ( .A(in[1399]), .B(n4019), .Z(n4707) );
  NAND U1314 ( .A(n4710), .B(n4707), .Z(n797) );
  XNOR U1315 ( .A(n1474), .B(n797), .Z(out[1043]) );
  XNOR U1316 ( .A(n799), .B(n798), .Z(n3712) );
  XNOR U1317 ( .A(in[551]), .B(n3712), .Z(n1478) );
  XOR U1318 ( .A(in[855]), .B(in[1175]), .Z(n801) );
  XNOR U1319 ( .A(in[1495]), .B(in[215]), .Z(n800) );
  XNOR U1320 ( .A(n801), .B(n800), .Z(n802) );
  XNOR U1321 ( .A(in[535]), .B(n802), .Z(n1259) );
  XNOR U1322 ( .A(n803), .B(n1259), .Z(n3661) );
  XNOR U1323 ( .A(in[151]), .B(n3661), .Z(n4718) );
  XOR U1324 ( .A(in[824]), .B(in[504]), .Z(n805) );
  XNOR U1325 ( .A(in[1464]), .B(in[1144]), .Z(n804) );
  XNOR U1326 ( .A(n805), .B(n804), .Z(n806) );
  XOR U1327 ( .A(in[184]), .B(n806), .Z(n1045) );
  XOR U1328 ( .A(in[1335]), .B(in[55]), .Z(n808) );
  XNOR U1329 ( .A(in[695]), .B(in[375]), .Z(n807) );
  XNOR U1330 ( .A(n808), .B(n807), .Z(n809) );
  XOR U1331 ( .A(in[1015]), .B(n809), .Z(n1373) );
  XNOR U1332 ( .A(n1045), .B(n1373), .Z(n4022) );
  XNOR U1333 ( .A(in[1400]), .B(n4022), .Z(n4715) );
  NAND U1334 ( .A(n4718), .B(n4715), .Z(n810) );
  XNOR U1335 ( .A(n1478), .B(n810), .Z(out[1044]) );
  XNOR U1336 ( .A(n812), .B(n811), .Z(n3716) );
  XNOR U1337 ( .A(in[552]), .B(n3716), .Z(n1482) );
  XOR U1338 ( .A(in[856]), .B(in[1176]), .Z(n814) );
  XNOR U1339 ( .A(in[1496]), .B(in[216]), .Z(n813) );
  XNOR U1340 ( .A(n814), .B(n813), .Z(n815) );
  XNOR U1341 ( .A(in[536]), .B(n815), .Z(n1262) );
  XNOR U1342 ( .A(n816), .B(n1262), .Z(n3669) );
  XNOR U1343 ( .A(in[152]), .B(n3669), .Z(n4722) );
  XOR U1344 ( .A(in[825]), .B(in[505]), .Z(n818) );
  XNOR U1345 ( .A(in[1465]), .B(in[1145]), .Z(n817) );
  XNOR U1346 ( .A(n818), .B(n817), .Z(n819) );
  XOR U1347 ( .A(in[185]), .B(n819), .Z(n1056) );
  XOR U1348 ( .A(in[1336]), .B(in[56]), .Z(n821) );
  XNOR U1349 ( .A(in[696]), .B(in[376]), .Z(n820) );
  XNOR U1350 ( .A(n821), .B(n820), .Z(n822) );
  XOR U1351 ( .A(in[1016]), .B(n822), .Z(n1377) );
  XNOR U1352 ( .A(n1056), .B(n1377), .Z(n4025) );
  XNOR U1353 ( .A(in[1401]), .B(n4025), .Z(n4719) );
  NAND U1354 ( .A(n4722), .B(n4719), .Z(n823) );
  XNOR U1355 ( .A(n1482), .B(n823), .Z(out[1045]) );
  XNOR U1356 ( .A(n825), .B(n824), .Z(n3720) );
  XNOR U1357 ( .A(in[553]), .B(n3720), .Z(n1486) );
  XOR U1358 ( .A(in[857]), .B(in[1177]), .Z(n827) );
  XNOR U1359 ( .A(in[1497]), .B(in[217]), .Z(n826) );
  XNOR U1360 ( .A(n827), .B(n826), .Z(n828) );
  XNOR U1361 ( .A(in[537]), .B(n828), .Z(n1265) );
  XNOR U1362 ( .A(n829), .B(n1265), .Z(n3673) );
  XNOR U1363 ( .A(in[153]), .B(n3673), .Z(n4726) );
  XOR U1364 ( .A(in[1337]), .B(in[57]), .Z(n831) );
  XNOR U1365 ( .A(in[697]), .B(in[377]), .Z(n830) );
  XNOR U1366 ( .A(n831), .B(n830), .Z(n832) );
  XOR U1367 ( .A(in[1017]), .B(n832), .Z(n1381) );
  XOR U1368 ( .A(in[826]), .B(in[506]), .Z(n834) );
  XNOR U1369 ( .A(in[1466]), .B(in[1146]), .Z(n833) );
  XNOR U1370 ( .A(n834), .B(n833), .Z(n835) );
  XOR U1371 ( .A(in[186]), .B(n835), .Z(n1067) );
  XNOR U1372 ( .A(n1381), .B(n1067), .Z(n4028) );
  XNOR U1373 ( .A(in[1402]), .B(n4028), .Z(n4723) );
  NAND U1374 ( .A(n4726), .B(n4723), .Z(n836) );
  XNOR U1375 ( .A(n1486), .B(n836), .Z(out[1046]) );
  XNOR U1376 ( .A(n838), .B(n837), .Z(n3724) );
  XNOR U1377 ( .A(in[554]), .B(n3724), .Z(n1490) );
  XOR U1378 ( .A(in[858]), .B(in[1178]), .Z(n840) );
  XNOR U1379 ( .A(in[1498]), .B(in[218]), .Z(n839) );
  XNOR U1380 ( .A(n840), .B(n839), .Z(n841) );
  XNOR U1381 ( .A(in[538]), .B(n841), .Z(n1268) );
  XNOR U1382 ( .A(n842), .B(n1268), .Z(n3677) );
  XNOR U1383 ( .A(in[154]), .B(n3677), .Z(n4730) );
  XOR U1384 ( .A(in[1338]), .B(in[58]), .Z(n844) );
  XNOR U1385 ( .A(in[698]), .B(in[378]), .Z(n843) );
  XNOR U1386 ( .A(n844), .B(n843), .Z(n845) );
  XOR U1387 ( .A(in[1018]), .B(n845), .Z(n1385) );
  XOR U1388 ( .A(in[827]), .B(in[507]), .Z(n847) );
  XNOR U1389 ( .A(in[1467]), .B(in[1147]), .Z(n846) );
  XNOR U1390 ( .A(n847), .B(n846), .Z(n848) );
  XOR U1391 ( .A(in[187]), .B(n848), .Z(n1072) );
  XNOR U1392 ( .A(n1385), .B(n1072), .Z(n4031) );
  XNOR U1393 ( .A(in[1403]), .B(n4031), .Z(n4727) );
  NAND U1394 ( .A(n4730), .B(n4727), .Z(n849) );
  XNOR U1395 ( .A(n1490), .B(n849), .Z(out[1047]) );
  XOR U1396 ( .A(in[1579]), .B(in[619]), .Z(n851) );
  XNOR U1397 ( .A(in[939]), .B(in[299]), .Z(n850) );
  XNOR U1398 ( .A(n851), .B(n850), .Z(n852) );
  XOR U1399 ( .A(in[1259]), .B(n852), .Z(n1394) );
  XNOR U1400 ( .A(n853), .B(n1394), .Z(n3728) );
  XNOR U1401 ( .A(in[555]), .B(n3728), .Z(n1494) );
  XOR U1402 ( .A(in[859]), .B(in[1179]), .Z(n855) );
  XNOR U1403 ( .A(in[1499]), .B(in[219]), .Z(n854) );
  XNOR U1404 ( .A(n855), .B(n854), .Z(n856) );
  XNOR U1405 ( .A(in[539]), .B(n856), .Z(n1271) );
  XNOR U1406 ( .A(n857), .B(n1271), .Z(n3681) );
  XNOR U1407 ( .A(in[155]), .B(n3681), .Z(n4734) );
  XOR U1408 ( .A(in[828]), .B(in[508]), .Z(n859) );
  XNOR U1409 ( .A(in[1468]), .B(in[1148]), .Z(n858) );
  XNOR U1410 ( .A(n859), .B(n858), .Z(n860) );
  XOR U1411 ( .A(in[188]), .B(n860), .Z(n1077) );
  XNOR U1412 ( .A(n861), .B(n1077), .Z(n4034) );
  XNOR U1413 ( .A(in[1404]), .B(n4034), .Z(n4731) );
  NAND U1414 ( .A(n4734), .B(n4731), .Z(n862) );
  XNOR U1415 ( .A(n1494), .B(n862), .Z(out[1048]) );
  XOR U1416 ( .A(in[1580]), .B(in[620]), .Z(n864) );
  XNOR U1417 ( .A(in[940]), .B(in[300]), .Z(n863) );
  XNOR U1418 ( .A(n864), .B(n863), .Z(n865) );
  XOR U1419 ( .A(in[1260]), .B(n865), .Z(n1398) );
  XNOR U1420 ( .A(n866), .B(n1398), .Z(n3732) );
  XNOR U1421 ( .A(in[556]), .B(n3732), .Z(n1498) );
  XOR U1422 ( .A(in[860]), .B(in[1180]), .Z(n868) );
  XNOR U1423 ( .A(in[1500]), .B(in[220]), .Z(n867) );
  XNOR U1424 ( .A(n868), .B(n867), .Z(n869) );
  XNOR U1425 ( .A(in[540]), .B(n869), .Z(n1275) );
  XNOR U1426 ( .A(n870), .B(n1275), .Z(n3685) );
  XNOR U1427 ( .A(in[156]), .B(n3685), .Z(n4738) );
  XNOR U1428 ( .A(n872), .B(n871), .Z(n4041) );
  XNOR U1429 ( .A(in[1405]), .B(n4041), .Z(n4735) );
  NAND U1430 ( .A(n4738), .B(n4735), .Z(n873) );
  XNOR U1431 ( .A(n1498), .B(n873), .Z(out[1049]) );
  XOR U1432 ( .A(in[1343]), .B(in[63]), .Z(n875) );
  XNOR U1433 ( .A(in[703]), .B(in[383]), .Z(n874) );
  XNOR U1434 ( .A(n875), .B(n874), .Z(n876) );
  XOR U1435 ( .A(in[1023]), .B(n876), .Z(n920) );
  XNOR U1436 ( .A(n877), .B(n920), .Z(n3607) );
  XNOR U1437 ( .A(in[639]), .B(n3607), .Z(n2558) );
  XOR U1438 ( .A(in[230]), .B(n3704), .Z(n2888) );
  XOR U1439 ( .A(in[874]), .B(in[1194]), .Z(n879) );
  XNOR U1440 ( .A(in[1514]), .B(in[234]), .Z(n878) );
  XNOR U1441 ( .A(n879), .B(n878), .Z(n880) );
  XOR U1442 ( .A(in[554]), .B(n880), .Z(n1324) );
  XNOR U1443 ( .A(n881), .B(n1324), .Z(n3745) );
  XNOR U1444 ( .A(in[1450]), .B(n3745), .Z(n2885) );
  NAND U1445 ( .A(n2888), .B(n2885), .Z(n882) );
  XNOR U1446 ( .A(n2558), .B(n882), .Z(out[104]) );
  XOR U1447 ( .A(in[1581]), .B(in[621]), .Z(n884) );
  XNOR U1448 ( .A(in[941]), .B(in[301]), .Z(n883) );
  XNOR U1449 ( .A(n884), .B(n883), .Z(n885) );
  XOR U1450 ( .A(in[1261]), .B(n885), .Z(n1402) );
  XNOR U1451 ( .A(n886), .B(n1402), .Z(n3736) );
  XNOR U1452 ( .A(in[557]), .B(n3736), .Z(n1502) );
  XOR U1453 ( .A(in[861]), .B(in[1181]), .Z(n888) );
  XNOR U1454 ( .A(in[1501]), .B(in[221]), .Z(n887) );
  XNOR U1455 ( .A(n888), .B(n887), .Z(n889) );
  XNOR U1456 ( .A(in[541]), .B(n889), .Z(n1278) );
  XNOR U1457 ( .A(n890), .B(n1278), .Z(n3689) );
  XNOR U1458 ( .A(in[157]), .B(n3689), .Z(n4742) );
  XOR U1459 ( .A(in[830]), .B(in[510]), .Z(n892) );
  XNOR U1460 ( .A(in[1470]), .B(in[1150]), .Z(n891) );
  XNOR U1461 ( .A(n892), .B(n891), .Z(n893) );
  XOR U1462 ( .A(in[190]), .B(n893), .Z(n1083) );
  XNOR U1463 ( .A(n894), .B(n1083), .Z(n4044) );
  XNOR U1464 ( .A(in[1406]), .B(n4044), .Z(n4739) );
  NAND U1465 ( .A(n4742), .B(n4739), .Z(n895) );
  XNOR U1466 ( .A(n1502), .B(n895), .Z(out[1050]) );
  XOR U1467 ( .A(in[1582]), .B(in[622]), .Z(n897) );
  XNOR U1468 ( .A(in[942]), .B(in[302]), .Z(n896) );
  XNOR U1469 ( .A(n897), .B(n896), .Z(n898) );
  XOR U1470 ( .A(in[1262]), .B(n898), .Z(n1406) );
  XNOR U1471 ( .A(n899), .B(n1406), .Z(n3740) );
  XNOR U1472 ( .A(in[558]), .B(n3740), .Z(n1506) );
  XOR U1473 ( .A(in[862]), .B(in[1182]), .Z(n901) );
  XNOR U1474 ( .A(in[1502]), .B(in[222]), .Z(n900) );
  XNOR U1475 ( .A(n901), .B(n900), .Z(n902) );
  XNOR U1476 ( .A(in[542]), .B(n902), .Z(n1281) );
  XNOR U1477 ( .A(n903), .B(n1281), .Z(n3693) );
  XNOR U1478 ( .A(in[158]), .B(n3693), .Z(n4746) );
  XOR U1479 ( .A(in[831]), .B(in[511]), .Z(n905) );
  XNOR U1480 ( .A(in[1471]), .B(in[1151]), .Z(n904) );
  XNOR U1481 ( .A(n905), .B(n904), .Z(n906) );
  XOR U1482 ( .A(in[191]), .B(n906), .Z(n1088) );
  XNOR U1483 ( .A(n907), .B(n1088), .Z(n4047) );
  XNOR U1484 ( .A(in[1407]), .B(n4047), .Z(n4743) );
  NAND U1485 ( .A(n4746), .B(n4743), .Z(n908) );
  XNOR U1486 ( .A(n1506), .B(n908), .Z(out[1051]) );
  XOR U1487 ( .A(in[1583]), .B(in[623]), .Z(n910) );
  XNOR U1488 ( .A(in[943]), .B(in[303]), .Z(n909) );
  XNOR U1489 ( .A(n910), .B(n909), .Z(n911) );
  XOR U1490 ( .A(in[1263]), .B(n911), .Z(n1410) );
  XNOR U1491 ( .A(n912), .B(n1410), .Z(n3744) );
  XNOR U1492 ( .A(in[559]), .B(n3744), .Z(n1511) );
  XOR U1493 ( .A(in[863]), .B(in[1183]), .Z(n914) );
  XNOR U1494 ( .A(in[1503]), .B(in[223]), .Z(n913) );
  XNOR U1495 ( .A(n914), .B(n913), .Z(n915) );
  XNOR U1496 ( .A(in[543]), .B(n915), .Z(n1284) );
  XNOR U1497 ( .A(n916), .B(n1284), .Z(n3697) );
  XNOR U1498 ( .A(in[159]), .B(n3697), .Z(n4750) );
  XOR U1499 ( .A(in[768]), .B(in[1088]), .Z(n918) );
  XNOR U1500 ( .A(in[448]), .B(in[1408]), .Z(n917) );
  XNOR U1501 ( .A(n918), .B(n917), .Z(n919) );
  XOR U1502 ( .A(in[128]), .B(n919), .Z(n1096) );
  XNOR U1503 ( .A(n920), .B(n1096), .Z(n4050) );
  XNOR U1504 ( .A(in[1344]), .B(n4050), .Z(n4747) );
  NAND U1505 ( .A(n4750), .B(n4747), .Z(n921) );
  XNOR U1506 ( .A(n1511), .B(n921), .Z(out[1052]) );
  XOR U1507 ( .A(in[1584]), .B(in[624]), .Z(n923) );
  XNOR U1508 ( .A(in[944]), .B(in[304]), .Z(n922) );
  XNOR U1509 ( .A(n923), .B(n922), .Z(n924) );
  XOR U1510 ( .A(in[1264]), .B(n924), .Z(n1414) );
  XNOR U1511 ( .A(n925), .B(n1414), .Z(n3748) );
  XNOR U1512 ( .A(in[560]), .B(n3748), .Z(n1515) );
  XOR U1513 ( .A(in[224]), .B(in[864]), .Z(n927) );
  XNOR U1514 ( .A(in[1184]), .B(in[1504]), .Z(n926) );
  XNOR U1515 ( .A(n927), .B(n926), .Z(n928) );
  XNOR U1516 ( .A(in[544]), .B(n928), .Z(n1287) );
  XNOR U1517 ( .A(n929), .B(n1287), .Z(n3701) );
  XNOR U1518 ( .A(in[160]), .B(n3701), .Z(n4754) );
  XOR U1519 ( .A(in[1280]), .B(in[640]), .Z(n931) );
  XNOR U1520 ( .A(in[960]), .B(in[320]), .Z(n930) );
  XNOR U1521 ( .A(n931), .B(n930), .Z(n932) );
  XOR U1522 ( .A(in[0]), .B(n932), .Z(n1023) );
  XOR U1523 ( .A(in[769]), .B(in[1089]), .Z(n934) );
  XNOR U1524 ( .A(in[449]), .B(in[1409]), .Z(n933) );
  XNOR U1525 ( .A(n934), .B(n933), .Z(n935) );
  XOR U1526 ( .A(in[129]), .B(n935), .Z(n1101) );
  XNOR U1527 ( .A(n1023), .B(n1101), .Z(n4053) );
  XNOR U1528 ( .A(in[1345]), .B(n4053), .Z(n4751) );
  NAND U1529 ( .A(n4754), .B(n4751), .Z(n936) );
  XNOR U1530 ( .A(n1515), .B(n936), .Z(out[1053]) );
  XOR U1531 ( .A(in[1585]), .B(in[625]), .Z(n938) );
  XNOR U1532 ( .A(in[945]), .B(in[305]), .Z(n937) );
  XNOR U1533 ( .A(n938), .B(n937), .Z(n939) );
  XOR U1534 ( .A(in[1265]), .B(n939), .Z(n1418) );
  XNOR U1535 ( .A(n940), .B(n1418), .Z(n3756) );
  XNOR U1536 ( .A(in[561]), .B(n3756), .Z(n1519) );
  XOR U1537 ( .A(in[225]), .B(in[865]), .Z(n942) );
  XNOR U1538 ( .A(in[1185]), .B(in[1505]), .Z(n941) );
  XNOR U1539 ( .A(n942), .B(n941), .Z(n943) );
  XNOR U1540 ( .A(in[545]), .B(n943), .Z(n1290) );
  XNOR U1541 ( .A(n944), .B(n1290), .Z(n3705) );
  XNOR U1542 ( .A(in[161]), .B(n3705), .Z(n4762) );
  XOR U1543 ( .A(in[1]), .B(in[641]), .Z(n946) );
  XNOR U1544 ( .A(in[961]), .B(in[321]), .Z(n945) );
  XNOR U1545 ( .A(n946), .B(n945), .Z(n947) );
  XOR U1546 ( .A(in[1281]), .B(n947), .Z(n1090) );
  XOR U1547 ( .A(in[1090]), .B(in[450]), .Z(n949) );
  XNOR U1548 ( .A(in[130]), .B(in[770]), .Z(n948) );
  XNOR U1549 ( .A(n949), .B(n948), .Z(n950) );
  XOR U1550 ( .A(in[1410]), .B(n950), .Z(n1106) );
  XNOR U1551 ( .A(n1090), .B(n1106), .Z(n4056) );
  XNOR U1552 ( .A(in[1346]), .B(n4056), .Z(n4759) );
  NAND U1553 ( .A(n4762), .B(n4759), .Z(n951) );
  XNOR U1554 ( .A(n1519), .B(n951), .Z(out[1054]) );
  XOR U1555 ( .A(in[1586]), .B(in[626]), .Z(n953) );
  XNOR U1556 ( .A(in[946]), .B(in[306]), .Z(n952) );
  XNOR U1557 ( .A(n953), .B(n952), .Z(n954) );
  XOR U1558 ( .A(in[1266]), .B(n954), .Z(n1422) );
  XNOR U1559 ( .A(n955), .B(n1422), .Z(n3760) );
  XNOR U1560 ( .A(in[562]), .B(n3760), .Z(n1523) );
  XOR U1561 ( .A(in[1186]), .B(in[1506]), .Z(n957) );
  XNOR U1562 ( .A(in[546]), .B(in[866]), .Z(n956) );
  XNOR U1563 ( .A(n957), .B(n956), .Z(n958) );
  XNOR U1564 ( .A(in[226]), .B(n958), .Z(n1293) );
  XNOR U1565 ( .A(n959), .B(n1293), .Z(n3713) );
  XNOR U1566 ( .A(in[162]), .B(n3713), .Z(n4766) );
  XOR U1567 ( .A(in[2]), .B(in[642]), .Z(n961) );
  XNOR U1568 ( .A(in[962]), .B(in[322]), .Z(n960) );
  XNOR U1569 ( .A(n961), .B(n960), .Z(n962) );
  XOR U1570 ( .A(in[1282]), .B(n962), .Z(n1143) );
  XOR U1571 ( .A(in[771]), .B(in[1091]), .Z(n964) );
  XNOR U1572 ( .A(in[451]), .B(in[1411]), .Z(n963) );
  XNOR U1573 ( .A(n964), .B(n963), .Z(n965) );
  XOR U1574 ( .A(in[131]), .B(n965), .Z(n1111) );
  XNOR U1575 ( .A(n1143), .B(n1111), .Z(n4059) );
  XNOR U1576 ( .A(in[1347]), .B(n4059), .Z(n4763) );
  NAND U1577 ( .A(n4766), .B(n4763), .Z(n966) );
  XNOR U1578 ( .A(n1523), .B(n966), .Z(out[1055]) );
  XOR U1579 ( .A(in[1587]), .B(in[627]), .Z(n968) );
  XNOR U1580 ( .A(in[947]), .B(in[307]), .Z(n967) );
  XNOR U1581 ( .A(n968), .B(n967), .Z(n969) );
  XOR U1582 ( .A(in[1267]), .B(n969), .Z(n1427) );
  XNOR U1583 ( .A(n970), .B(n1427), .Z(n3764) );
  XNOR U1584 ( .A(in[563]), .B(n3764), .Z(n1527) );
  XOR U1585 ( .A(in[1187]), .B(in[1507]), .Z(n972) );
  XNOR U1586 ( .A(in[547]), .B(in[867]), .Z(n971) );
  XNOR U1587 ( .A(n972), .B(n971), .Z(n973) );
  XNOR U1588 ( .A(in[227]), .B(n973), .Z(n1296) );
  XNOR U1589 ( .A(n974), .B(n1296), .Z(n3717) );
  XNOR U1590 ( .A(in[163]), .B(n3717), .Z(n4770) );
  XOR U1591 ( .A(in[772]), .B(in[1092]), .Z(n976) );
  XNOR U1592 ( .A(in[452]), .B(in[1412]), .Z(n975) );
  XNOR U1593 ( .A(n976), .B(n975), .Z(n977) );
  XOR U1594 ( .A(in[132]), .B(n977), .Z(n1116) );
  XOR U1595 ( .A(in[323]), .B(in[643]), .Z(n979) );
  XNOR U1596 ( .A(in[963]), .B(in[3]), .Z(n978) );
  XNOR U1597 ( .A(n979), .B(n978), .Z(n980) );
  XOR U1598 ( .A(in[1283]), .B(n980), .Z(n1189) );
  XNOR U1599 ( .A(n1116), .B(n1189), .Z(n4062) );
  XNOR U1600 ( .A(in[1348]), .B(n4062), .Z(n4767) );
  NAND U1601 ( .A(n4770), .B(n4767), .Z(n981) );
  XNOR U1602 ( .A(n1527), .B(n981), .Z(out[1056]) );
  XOR U1603 ( .A(in[1588]), .B(in[628]), .Z(n983) );
  XNOR U1604 ( .A(in[948]), .B(in[308]), .Z(n982) );
  XNOR U1605 ( .A(n983), .B(n982), .Z(n984) );
  XOR U1606 ( .A(in[1268]), .B(n984), .Z(n1431) );
  XNOR U1607 ( .A(n985), .B(n1431), .Z(n3768) );
  XNOR U1608 ( .A(in[564]), .B(n3768), .Z(n1531) );
  XOR U1609 ( .A(in[1188]), .B(in[1508]), .Z(n987) );
  XNOR U1610 ( .A(in[548]), .B(in[868]), .Z(n986) );
  XNOR U1611 ( .A(n987), .B(n986), .Z(n988) );
  XOR U1612 ( .A(in[228]), .B(n988), .Z(n1299) );
  XNOR U1613 ( .A(n1299), .B(n989), .Z(n3721) );
  XNOR U1614 ( .A(in[164]), .B(n3721), .Z(n4774) );
  XOR U1615 ( .A(in[773]), .B(in[1093]), .Z(n991) );
  XNOR U1616 ( .A(in[453]), .B(in[1413]), .Z(n990) );
  XNOR U1617 ( .A(n991), .B(n990), .Z(n992) );
  XOR U1618 ( .A(in[133]), .B(n992), .Z(n1121) );
  XOR U1619 ( .A(in[324]), .B(in[644]), .Z(n994) );
  XNOR U1620 ( .A(in[964]), .B(in[4]), .Z(n993) );
  XNOR U1621 ( .A(n994), .B(n993), .Z(n995) );
  XOR U1622 ( .A(in[1284]), .B(n995), .Z(n1197) );
  XNOR U1623 ( .A(n1121), .B(n1197), .Z(n4065) );
  XNOR U1624 ( .A(in[1349]), .B(n4065), .Z(n4771) );
  NAND U1625 ( .A(n4774), .B(n4771), .Z(n996) );
  XNOR U1626 ( .A(n1531), .B(n996), .Z(out[1057]) );
  XOR U1627 ( .A(in[1589]), .B(in[629]), .Z(n998) );
  XNOR U1628 ( .A(in[949]), .B(in[309]), .Z(n997) );
  XNOR U1629 ( .A(n998), .B(n997), .Z(n999) );
  XOR U1630 ( .A(in[1269]), .B(n999), .Z(n1435) );
  XNOR U1631 ( .A(n1000), .B(n1435), .Z(n3772) );
  XNOR U1632 ( .A(in[565]), .B(n3772), .Z(n1535) );
  XOR U1633 ( .A(in[1189]), .B(in[1509]), .Z(n1002) );
  XNOR U1634 ( .A(in[549]), .B(in[869]), .Z(n1001) );
  XNOR U1635 ( .A(n1002), .B(n1001), .Z(n1003) );
  XNOR U1636 ( .A(in[229]), .B(n1003), .Z(n1303) );
  XNOR U1637 ( .A(n1004), .B(n1303), .Z(n3725) );
  XNOR U1638 ( .A(in[165]), .B(n3725), .Z(n4778) );
  XOR U1639 ( .A(in[774]), .B(in[1094]), .Z(n1006) );
  XNOR U1640 ( .A(in[454]), .B(in[1414]), .Z(n1005) );
  XNOR U1641 ( .A(n1006), .B(n1005), .Z(n1007) );
  XOR U1642 ( .A(in[134]), .B(n1007), .Z(n1126) );
  XOR U1643 ( .A(in[325]), .B(in[645]), .Z(n1009) );
  XNOR U1644 ( .A(in[965]), .B(in[5]), .Z(n1008) );
  XNOR U1645 ( .A(n1009), .B(n1008), .Z(n1010) );
  XOR U1646 ( .A(in[1285]), .B(n1010), .Z(n1200) );
  XNOR U1647 ( .A(n1126), .B(n1200), .Z(n4068) );
  XNOR U1648 ( .A(in[1350]), .B(n4068), .Z(n4775) );
  NAND U1649 ( .A(n4778), .B(n4775), .Z(n1011) );
  XNOR U1650 ( .A(n1535), .B(n1011), .Z(out[1058]) );
  XOR U1651 ( .A(in[1590]), .B(in[630]), .Z(n1013) );
  XNOR U1652 ( .A(in[950]), .B(in[310]), .Z(n1012) );
  XNOR U1653 ( .A(n1013), .B(n1012), .Z(n1014) );
  XOR U1654 ( .A(in[1270]), .B(n1014), .Z(n1439) );
  XNOR U1655 ( .A(n1015), .B(n1439), .Z(n3776) );
  XNOR U1656 ( .A(in[566]), .B(n3776), .Z(n1539) );
  XOR U1657 ( .A(in[166]), .B(n3729), .Z(n4782) );
  XOR U1658 ( .A(in[326]), .B(in[6]), .Z(n1017) );
  XNOR U1659 ( .A(in[966]), .B(in[646]), .Z(n1016) );
  XNOR U1660 ( .A(n1017), .B(n1016), .Z(n1018) );
  XOR U1661 ( .A(in[1286]), .B(n1018), .Z(n1203) );
  XOR U1662 ( .A(in[775]), .B(in[1095]), .Z(n1020) );
  XNOR U1663 ( .A(in[455]), .B(in[1415]), .Z(n1019) );
  XNOR U1664 ( .A(n1020), .B(n1019), .Z(n1021) );
  XOR U1665 ( .A(in[135]), .B(n1021), .Z(n1131) );
  XNOR U1666 ( .A(n1203), .B(n1131), .Z(n4079) );
  XNOR U1667 ( .A(in[1351]), .B(n4079), .Z(n4779) );
  NAND U1668 ( .A(n4782), .B(n4779), .Z(n1022) );
  XNOR U1669 ( .A(n1539), .B(n1022), .Z(out[1059]) );
  XNOR U1670 ( .A(n1024), .B(n1023), .Z(n3611) );
  XNOR U1671 ( .A(in[576]), .B(n3611), .Z(n2560) );
  XOR U1672 ( .A(in[231]), .B(n3712), .Z(n2902) );
  XNOR U1673 ( .A(in[1451]), .B(n3749), .Z(n2899) );
  NAND U1674 ( .A(n2902), .B(n2899), .Z(n1025) );
  XNOR U1675 ( .A(n2560), .B(n1025), .Z(out[105]) );
  XOR U1676 ( .A(in[1591]), .B(in[631]), .Z(n1027) );
  XNOR U1677 ( .A(in[951]), .B(in[311]), .Z(n1026) );
  XNOR U1678 ( .A(n1027), .B(n1026), .Z(n1028) );
  XOR U1679 ( .A(in[1271]), .B(n1028), .Z(n1443) );
  XNOR U1680 ( .A(n1029), .B(n1443), .Z(n3780) );
  XNOR U1681 ( .A(in[567]), .B(n3780), .Z(n1543) );
  XOR U1682 ( .A(in[167]), .B(n3733), .Z(n4786) );
  XOR U1683 ( .A(in[327]), .B(in[7]), .Z(n1031) );
  XNOR U1684 ( .A(in[967]), .B(in[647]), .Z(n1030) );
  XNOR U1685 ( .A(n1031), .B(n1030), .Z(n1032) );
  XOR U1686 ( .A(in[1287]), .B(n1032), .Z(n1206) );
  XOR U1687 ( .A(in[776]), .B(in[1096]), .Z(n1034) );
  XNOR U1688 ( .A(in[456]), .B(in[1416]), .Z(n1033) );
  XNOR U1689 ( .A(n1034), .B(n1033), .Z(n1035) );
  XOR U1690 ( .A(in[136]), .B(n1035), .Z(n1136) );
  XNOR U1691 ( .A(n1206), .B(n1136), .Z(n4082) );
  XNOR U1692 ( .A(in[1352]), .B(n4082), .Z(n4783) );
  NAND U1693 ( .A(n4786), .B(n4783), .Z(n1036) );
  XNOR U1694 ( .A(n1543), .B(n1036), .Z(out[1060]) );
  XOR U1695 ( .A(in[632]), .B(in[1592]), .Z(n1038) );
  XNOR U1696 ( .A(in[1272]), .B(in[312]), .Z(n1037) );
  XNOR U1697 ( .A(n1038), .B(n1037), .Z(n1039) );
  XOR U1698 ( .A(in[952]), .B(n1039), .Z(n1447) );
  XNOR U1699 ( .A(n1040), .B(n1447), .Z(n3784) );
  XNOR U1700 ( .A(in[568]), .B(n3784), .Z(n1547) );
  XOR U1701 ( .A(in[168]), .B(n3737), .Z(n4790) );
  XNOR U1702 ( .A(in[1353]), .B(n4085), .Z(n4787) );
  NAND U1703 ( .A(n4790), .B(n4787), .Z(n1041) );
  XNOR U1704 ( .A(n1547), .B(n1041), .Z(out[1061]) );
  XOR U1705 ( .A(in[633]), .B(in[1593]), .Z(n1043) );
  XNOR U1706 ( .A(in[1273]), .B(in[313]), .Z(n1042) );
  XNOR U1707 ( .A(n1043), .B(n1042), .Z(n1044) );
  XOR U1708 ( .A(in[953]), .B(n1044), .Z(n1451) );
  XNOR U1709 ( .A(n1045), .B(n1451), .Z(n3788) );
  XNOR U1710 ( .A(in[569]), .B(n3788), .Z(n1552) );
  XOR U1711 ( .A(in[169]), .B(n3741), .Z(n4794) );
  XOR U1712 ( .A(in[778]), .B(in[1098]), .Z(n1047) );
  XNOR U1713 ( .A(in[458]), .B(in[1418]), .Z(n1046) );
  XNOR U1714 ( .A(n1047), .B(n1046), .Z(n1048) );
  XOR U1715 ( .A(in[138]), .B(n1048), .Z(n1149) );
  XOR U1716 ( .A(in[329]), .B(in[969]), .Z(n1050) );
  XNOR U1717 ( .A(in[9]), .B(in[649]), .Z(n1049) );
  XNOR U1718 ( .A(n1050), .B(n1049), .Z(n1051) );
  XOR U1719 ( .A(in[1289]), .B(n1051), .Z(n1214) );
  XNOR U1720 ( .A(n1149), .B(n1214), .Z(n4088) );
  XNOR U1721 ( .A(in[1354]), .B(n4088), .Z(n4791) );
  NAND U1722 ( .A(n4794), .B(n4791), .Z(n1052) );
  XNOR U1723 ( .A(n1552), .B(n1052), .Z(out[1062]) );
  XOR U1724 ( .A(in[634]), .B(in[1594]), .Z(n1054) );
  XNOR U1725 ( .A(in[1274]), .B(in[314]), .Z(n1053) );
  XNOR U1726 ( .A(n1054), .B(n1053), .Z(n1055) );
  XOR U1727 ( .A(in[954]), .B(n1055), .Z(n1455) );
  XNOR U1728 ( .A(n1056), .B(n1455), .Z(n3792) );
  XNOR U1729 ( .A(in[570]), .B(n3792), .Z(n1556) );
  XOR U1730 ( .A(in[170]), .B(n3745), .Z(n4798) );
  XOR U1731 ( .A(in[1290]), .B(in[650]), .Z(n1058) );
  XNOR U1732 ( .A(in[970]), .B(in[330]), .Z(n1057) );
  XNOR U1733 ( .A(n1058), .B(n1057), .Z(n1059) );
  XOR U1734 ( .A(in[10]), .B(n1059), .Z(n1217) );
  XOR U1735 ( .A(in[1419]), .B(in[779]), .Z(n1061) );
  XNOR U1736 ( .A(in[1099]), .B(in[459]), .Z(n1060) );
  XNOR U1737 ( .A(n1061), .B(n1060), .Z(n1062) );
  XOR U1738 ( .A(in[139]), .B(n1062), .Z(n1154) );
  XNOR U1739 ( .A(n1217), .B(n1154), .Z(n4091) );
  XNOR U1740 ( .A(in[1355]), .B(n4091), .Z(n4795) );
  NAND U1741 ( .A(n4798), .B(n4795), .Z(n1063) );
  XNOR U1742 ( .A(n1556), .B(n1063), .Z(out[1063]) );
  XOR U1743 ( .A(in[955]), .B(in[1275]), .Z(n1065) );
  XNOR U1744 ( .A(in[1595]), .B(in[315]), .Z(n1064) );
  XNOR U1745 ( .A(n1065), .B(n1064), .Z(n1066) );
  XNOR U1746 ( .A(in[635]), .B(n1066), .Z(n1459) );
  XNOR U1747 ( .A(n1067), .B(n1459), .Z(n3802) );
  XNOR U1748 ( .A(in[571]), .B(n3802), .Z(n1558) );
  NOR U1749 ( .A(n1301), .B(n1696), .Z(n1068) );
  XNOR U1750 ( .A(n1558), .B(n1068), .Z(out[1064]) );
  XOR U1751 ( .A(in[956]), .B(in[1276]), .Z(n1070) );
  XNOR U1752 ( .A(in[1596]), .B(in[316]), .Z(n1069) );
  XNOR U1753 ( .A(n1070), .B(n1069), .Z(n1071) );
  XNOR U1754 ( .A(in[636]), .B(n1071), .Z(n1463) );
  XNOR U1755 ( .A(n1072), .B(n1463), .Z(n3806) );
  XNOR U1756 ( .A(in[572]), .B(n3806), .Z(n1560) );
  NOR U1757 ( .A(n1305), .B(n1700), .Z(n1073) );
  XNOR U1758 ( .A(n1560), .B(n1073), .Z(out[1065]) );
  XOR U1759 ( .A(in[957]), .B(in[1277]), .Z(n1075) );
  XNOR U1760 ( .A(in[1597]), .B(in[317]), .Z(n1074) );
  XNOR U1761 ( .A(n1075), .B(n1074), .Z(n1076) );
  XNOR U1762 ( .A(in[637]), .B(n1076), .Z(n1468) );
  XNOR U1763 ( .A(n1077), .B(n1468), .Z(n3810) );
  XNOR U1764 ( .A(in[573]), .B(n3810), .Z(n1562) );
  NOR U1765 ( .A(n1310), .B(n1704), .Z(n1078) );
  XNOR U1766 ( .A(n1562), .B(n1078), .Z(out[1066]) );
  XOR U1767 ( .A(in[574]), .B(n3814), .Z(n1564) );
  NOR U1768 ( .A(n1314), .B(n1708), .Z(n1079) );
  XNOR U1769 ( .A(n1564), .B(n1079), .Z(out[1067]) );
  XOR U1770 ( .A(in[959]), .B(in[1279]), .Z(n1081) );
  XNOR U1771 ( .A(in[1599]), .B(in[319]), .Z(n1080) );
  XNOR U1772 ( .A(n1081), .B(n1080), .Z(n1082) );
  XNOR U1773 ( .A(in[639]), .B(n1082), .Z(n1476) );
  XNOR U1774 ( .A(n1083), .B(n1476), .Z(n3536) );
  XNOR U1775 ( .A(in[575]), .B(n3536), .Z(n1566) );
  NOR U1776 ( .A(n1318), .B(n1713), .Z(n1084) );
  XNOR U1777 ( .A(n1566), .B(n1084), .Z(out[1068]) );
  XOR U1778 ( .A(in[896]), .B(in[1216]), .Z(n1086) );
  XNOR U1779 ( .A(in[1536]), .B(in[256]), .Z(n1085) );
  XNOR U1780 ( .A(n1086), .B(n1085), .Z(n1087) );
  XNOR U1781 ( .A(in[576]), .B(n1087), .Z(n1480) );
  XNOR U1782 ( .A(n1088), .B(n1480), .Z(n3540) );
  XNOR U1783 ( .A(in[512]), .B(n3540), .Z(n1568) );
  NOR U1784 ( .A(n1322), .B(n1717), .Z(n1089) );
  XNOR U1785 ( .A(n1568), .B(n1089), .Z(out[1069]) );
  XNOR U1786 ( .A(n1091), .B(n1090), .Z(n3615) );
  XNOR U1787 ( .A(in[577]), .B(n3615), .Z(n2562) );
  XOR U1788 ( .A(in[232]), .B(n3716), .Z(n2916) );
  XNOR U1789 ( .A(in[1452]), .B(n3757), .Z(n2913) );
  NAND U1790 ( .A(n2916), .B(n2913), .Z(n1092) );
  XNOR U1791 ( .A(n2562), .B(n1092), .Z(out[106]) );
  XOR U1792 ( .A(in[897]), .B(in[1217]), .Z(n1094) );
  XNOR U1793 ( .A(in[1537]), .B(in[257]), .Z(n1093) );
  XNOR U1794 ( .A(n1094), .B(n1093), .Z(n1095) );
  XNOR U1795 ( .A(in[577]), .B(n1095), .Z(n1484) );
  XNOR U1796 ( .A(n1096), .B(n1484), .Z(n3544) );
  XNOR U1797 ( .A(in[513]), .B(n3544), .Z(n1570) );
  NOR U1798 ( .A(n1326), .B(n1721), .Z(n1097) );
  XNOR U1799 ( .A(n1570), .B(n1097), .Z(out[1070]) );
  XOR U1800 ( .A(in[1538]), .B(in[578]), .Z(n1099) );
  XNOR U1801 ( .A(in[898]), .B(in[258]), .Z(n1098) );
  XNOR U1802 ( .A(n1099), .B(n1098), .Z(n1100) );
  XNOR U1803 ( .A(in[1218]), .B(n1100), .Z(n1488) );
  XNOR U1804 ( .A(n1101), .B(n1488), .Z(n3548) );
  XNOR U1805 ( .A(in[514]), .B(n3548), .Z(n1572) );
  NOR U1806 ( .A(n1330), .B(n1725), .Z(n1102) );
  XNOR U1807 ( .A(n1572), .B(n1102), .Z(out[1071]) );
  XOR U1808 ( .A(in[1539]), .B(in[579]), .Z(n1104) );
  XNOR U1809 ( .A(in[899]), .B(in[259]), .Z(n1103) );
  XNOR U1810 ( .A(n1104), .B(n1103), .Z(n1105) );
  XNOR U1811 ( .A(in[1219]), .B(n1105), .Z(n1492) );
  XNOR U1812 ( .A(n1106), .B(n1492), .Z(n3552) );
  XNOR U1813 ( .A(in[515]), .B(n3552), .Z(n1576) );
  NOR U1814 ( .A(n1334), .B(n1729), .Z(n1107) );
  XNOR U1815 ( .A(n1576), .B(n1107), .Z(out[1072]) );
  XOR U1816 ( .A(in[1540]), .B(in[580]), .Z(n1109) );
  XNOR U1817 ( .A(in[900]), .B(in[260]), .Z(n1108) );
  XNOR U1818 ( .A(n1109), .B(n1108), .Z(n1110) );
  XNOR U1819 ( .A(in[1220]), .B(n1110), .Z(n1496) );
  XNOR U1820 ( .A(n1111), .B(n1496), .Z(n3556) );
  XNOR U1821 ( .A(in[516]), .B(n3556), .Z(n1578) );
  NOR U1822 ( .A(n1338), .B(n1733), .Z(n1112) );
  XNOR U1823 ( .A(n1578), .B(n1112), .Z(out[1073]) );
  XOR U1824 ( .A(in[1541]), .B(in[581]), .Z(n1114) );
  XNOR U1825 ( .A(in[901]), .B(in[261]), .Z(n1113) );
  XNOR U1826 ( .A(n1114), .B(n1113), .Z(n1115) );
  XNOR U1827 ( .A(in[1221]), .B(n1115), .Z(n1500) );
  XNOR U1828 ( .A(n1116), .B(n1500), .Z(n3560) );
  XNOR U1829 ( .A(in[517]), .B(n3560), .Z(n1580) );
  NOR U1830 ( .A(n1342), .B(n1737), .Z(n1117) );
  XNOR U1831 ( .A(n1580), .B(n1117), .Z(out[1074]) );
  XOR U1832 ( .A(in[1542]), .B(in[582]), .Z(n1119) );
  XNOR U1833 ( .A(in[902]), .B(in[262]), .Z(n1118) );
  XNOR U1834 ( .A(n1119), .B(n1118), .Z(n1120) );
  XNOR U1835 ( .A(in[1222]), .B(n1120), .Z(n1504) );
  XNOR U1836 ( .A(n1121), .B(n1504), .Z(n3564) );
  XNOR U1837 ( .A(in[518]), .B(n3564), .Z(n1582) );
  NOR U1838 ( .A(n1346), .B(n1741), .Z(n1122) );
  XNOR U1839 ( .A(n1582), .B(n1122), .Z(out[1075]) );
  XOR U1840 ( .A(in[1543]), .B(in[583]), .Z(n1124) );
  XNOR U1841 ( .A(in[903]), .B(in[263]), .Z(n1123) );
  XNOR U1842 ( .A(n1124), .B(n1123), .Z(n1125) );
  XNOR U1843 ( .A(in[1223]), .B(n1125), .Z(n1509) );
  XNOR U1844 ( .A(n1126), .B(n1509), .Z(n3568) );
  XNOR U1845 ( .A(in[519]), .B(n3568), .Z(n1584) );
  NOR U1846 ( .A(n1351), .B(n1745), .Z(n1127) );
  XNOR U1847 ( .A(n1584), .B(n1127), .Z(out[1076]) );
  XOR U1848 ( .A(in[1544]), .B(in[584]), .Z(n1129) );
  XNOR U1849 ( .A(in[904]), .B(in[264]), .Z(n1128) );
  XNOR U1850 ( .A(n1129), .B(n1128), .Z(n1130) );
  XNOR U1851 ( .A(in[1224]), .B(n1130), .Z(n1513) );
  XNOR U1852 ( .A(n1131), .B(n1513), .Z(n3572) );
  XNOR U1853 ( .A(in[520]), .B(n3572), .Z(n1586) );
  NOR U1854 ( .A(n1355), .B(n1749), .Z(n1132) );
  XNOR U1855 ( .A(n1586), .B(n1132), .Z(out[1077]) );
  XOR U1856 ( .A(in[1545]), .B(in[585]), .Z(n1134) );
  XNOR U1857 ( .A(in[905]), .B(in[265]), .Z(n1133) );
  XNOR U1858 ( .A(n1134), .B(n1133), .Z(n1135) );
  XNOR U1859 ( .A(in[1225]), .B(n1135), .Z(n1517) );
  XNOR U1860 ( .A(n1136), .B(n1517), .Z(n3580) );
  XNOR U1861 ( .A(in[521]), .B(n3580), .Z(n1588) );
  NOR U1862 ( .A(n1359), .B(n1754), .Z(n1137) );
  XNOR U1863 ( .A(n1588), .B(n1137), .Z(out[1078]) );
  XOR U1864 ( .A(in[1546]), .B(in[586]), .Z(n1139) );
  XNOR U1865 ( .A(in[906]), .B(in[266]), .Z(n1138) );
  XNOR U1866 ( .A(n1139), .B(n1138), .Z(n1140) );
  XNOR U1867 ( .A(in[1226]), .B(n1140), .Z(n1521) );
  XNOR U1868 ( .A(n1141), .B(n1521), .Z(n3584) );
  XNOR U1869 ( .A(in[522]), .B(n3584), .Z(n1590) );
  NOR U1870 ( .A(n1363), .B(n1758), .Z(n1142) );
  XNOR U1871 ( .A(n1590), .B(n1142), .Z(out[1079]) );
  XNOR U1872 ( .A(n1144), .B(n1143), .Z(n3623) );
  XNOR U1873 ( .A(in[578]), .B(n3623), .Z(n2564) );
  XOR U1874 ( .A(in[233]), .B(n3720), .Z(n2930) );
  XNOR U1875 ( .A(in[1453]), .B(n3761), .Z(n2927) );
  NAND U1876 ( .A(n2930), .B(n2927), .Z(n1145) );
  XNOR U1877 ( .A(n2564), .B(n1145), .Z(out[107]) );
  XOR U1878 ( .A(in[1547]), .B(in[587]), .Z(n1147) );
  XNOR U1879 ( .A(in[907]), .B(in[267]), .Z(n1146) );
  XNOR U1880 ( .A(n1147), .B(n1146), .Z(n1148) );
  XNOR U1881 ( .A(in[1227]), .B(n1148), .Z(n1525) );
  XNOR U1882 ( .A(n1149), .B(n1525), .Z(n3588) );
  XNOR U1883 ( .A(in[523]), .B(n3588), .Z(n1592) );
  NOR U1884 ( .A(n1367), .B(n1762), .Z(n1150) );
  XNOR U1885 ( .A(n1592), .B(n1150), .Z(out[1080]) );
  XOR U1886 ( .A(in[1548]), .B(in[588]), .Z(n1152) );
  XNOR U1887 ( .A(in[908]), .B(in[268]), .Z(n1151) );
  XNOR U1888 ( .A(n1152), .B(n1151), .Z(n1153) );
  XNOR U1889 ( .A(in[1228]), .B(n1153), .Z(n1529) );
  XNOR U1890 ( .A(n1154), .B(n1529), .Z(n3592) );
  XNOR U1891 ( .A(in[524]), .B(n3592), .Z(n1594) );
  NOR U1892 ( .A(n1371), .B(n1766), .Z(n1155) );
  XNOR U1893 ( .A(n1594), .B(n1155), .Z(out[1081]) );
  XOR U1894 ( .A(in[1549]), .B(in[589]), .Z(n1157) );
  XNOR U1895 ( .A(in[909]), .B(in[269]), .Z(n1156) );
  XNOR U1896 ( .A(n1157), .B(n1156), .Z(n1158) );
  XOR U1897 ( .A(in[1229]), .B(n1158), .Z(n1533) );
  XNOR U1898 ( .A(n1533), .B(n1159), .Z(n3596) );
  XNOR U1899 ( .A(in[525]), .B(n3596), .Z(n1597) );
  NOR U1900 ( .A(n1375), .B(n1770), .Z(n1160) );
  XNOR U1901 ( .A(n1597), .B(n1160), .Z(out[1082]) );
  XOR U1902 ( .A(in[1550]), .B(in[590]), .Z(n1162) );
  XNOR U1903 ( .A(in[910]), .B(in[270]), .Z(n1161) );
  XNOR U1904 ( .A(n1162), .B(n1161), .Z(n1163) );
  XOR U1905 ( .A(in[1230]), .B(n1163), .Z(n1537) );
  XNOR U1906 ( .A(n1537), .B(n1164), .Z(n3600) );
  XNOR U1907 ( .A(in[526]), .B(n3600), .Z(n1599) );
  NOR U1908 ( .A(n1379), .B(n1774), .Z(n1165) );
  XNOR U1909 ( .A(n1599), .B(n1165), .Z(out[1083]) );
  XOR U1910 ( .A(in[1551]), .B(in[591]), .Z(n1167) );
  XNOR U1911 ( .A(in[911]), .B(in[271]), .Z(n1166) );
  XNOR U1912 ( .A(n1167), .B(n1166), .Z(n1168) );
  XNOR U1913 ( .A(in[1231]), .B(n1168), .Z(n1541) );
  XNOR U1914 ( .A(n1169), .B(n1541), .Z(n3604) );
  XNOR U1915 ( .A(in[527]), .B(n3604), .Z(n1601) );
  NOR U1916 ( .A(n1383), .B(n1778), .Z(n1170) );
  XNOR U1917 ( .A(n1601), .B(n1170), .Z(out[1084]) );
  XOR U1918 ( .A(in[1552]), .B(in[592]), .Z(n1172) );
  XNOR U1919 ( .A(in[912]), .B(in[272]), .Z(n1171) );
  XNOR U1920 ( .A(n1172), .B(n1171), .Z(n1173) );
  XNOR U1921 ( .A(in[1232]), .B(n1173), .Z(n1545) );
  XNOR U1922 ( .A(n1174), .B(n1545), .Z(n3608) );
  XNOR U1923 ( .A(in[528]), .B(n3608), .Z(n1603) );
  NOR U1924 ( .A(n1387), .B(n1782), .Z(n1175) );
  XNOR U1925 ( .A(n1603), .B(n1175), .Z(out[1085]) );
  XOR U1926 ( .A(in[1553]), .B(in[593]), .Z(n1177) );
  XNOR U1927 ( .A(in[913]), .B(in[273]), .Z(n1176) );
  XNOR U1928 ( .A(n1177), .B(n1176), .Z(n1178) );
  XNOR U1929 ( .A(in[1233]), .B(n1178), .Z(n1550) );
  XNOR U1930 ( .A(n1179), .B(n1550), .Z(n3612) );
  XNOR U1931 ( .A(in[529]), .B(n3612), .Z(n1605) );
  NOR U1932 ( .A(n1390), .B(n1786), .Z(n1180) );
  XNOR U1933 ( .A(n1605), .B(n1180), .Z(out[1086]) );
  XOR U1934 ( .A(in[1554]), .B(in[594]), .Z(n1182) );
  XNOR U1935 ( .A(in[914]), .B(in[274]), .Z(n1181) );
  XNOR U1936 ( .A(n1182), .B(n1181), .Z(n1183) );
  XNOR U1937 ( .A(in[1234]), .B(n1183), .Z(n1554) );
  XNOR U1938 ( .A(n1184), .B(n1554), .Z(n3616) );
  XNOR U1939 ( .A(in[530]), .B(n3616), .Z(n1607) );
  NOR U1940 ( .A(n1392), .B(n1790), .Z(n1185) );
  XNOR U1941 ( .A(n1607), .B(n1185), .Z(out[1087]) );
  XOR U1942 ( .A(in[957]), .B(n3599), .Z(n1609) );
  NOR U1943 ( .A(n1396), .B(n4630), .Z(n1186) );
  XNOR U1944 ( .A(n1609), .B(n1186), .Z(out[1088]) );
  XOR U1945 ( .A(in[958]), .B(n3603), .Z(n1611) );
  NOR U1946 ( .A(n1400), .B(n4634), .Z(n1187) );
  XNOR U1947 ( .A(n1611), .B(n1187), .Z(out[1089]) );
  XOR U1948 ( .A(n1189), .B(n1188), .Z(n3627) );
  XNOR U1949 ( .A(in[579]), .B(n3627), .Z(n2566) );
  XOR U1950 ( .A(in[234]), .B(n3724), .Z(n2946) );
  XNOR U1951 ( .A(in[1454]), .B(n3765), .Z(n2943) );
  NAND U1952 ( .A(n2946), .B(n2943), .Z(n1190) );
  XNOR U1953 ( .A(n2566), .B(n1190), .Z(out[108]) );
  XOR U1954 ( .A(in[959]), .B(n3607), .Z(n1613) );
  NOR U1955 ( .A(n1404), .B(n4638), .Z(n1191) );
  XNOR U1956 ( .A(n1613), .B(n1191), .Z(out[1090]) );
  XOR U1957 ( .A(in[896]), .B(n3611), .Z(n1615) );
  NOR U1958 ( .A(n1408), .B(n4642), .Z(n1192) );
  XNOR U1959 ( .A(n1615), .B(n1192), .Z(out[1091]) );
  XOR U1960 ( .A(in[897]), .B(n3615), .Z(n1618) );
  NOR U1961 ( .A(n1412), .B(n4646), .Z(n1193) );
  XNOR U1962 ( .A(n1618), .B(n1193), .Z(out[1092]) );
  XOR U1963 ( .A(in[898]), .B(n3623), .Z(n1620) );
  NOR U1964 ( .A(n1416), .B(n4650), .Z(n1194) );
  XNOR U1965 ( .A(n1620), .B(n1194), .Z(out[1093]) );
  XOR U1966 ( .A(in[899]), .B(n3627), .Z(n1622) );
  NOR U1967 ( .A(n1420), .B(n4654), .Z(n1195) );
  XNOR U1968 ( .A(n1622), .B(n1195), .Z(out[1094]) );
  XNOR U1969 ( .A(n1197), .B(n1196), .Z(n3631) );
  XNOR U1970 ( .A(in[900]), .B(n3631), .Z(n1624) );
  NOR U1971 ( .A(n1424), .B(n4658), .Z(n1198) );
  XNOR U1972 ( .A(n1624), .B(n1198), .Z(out[1095]) );
  XNOR U1973 ( .A(n1200), .B(n1199), .Z(n3635) );
  XNOR U1974 ( .A(in[901]), .B(n3635), .Z(n1626) );
  NOR U1975 ( .A(n1429), .B(n4662), .Z(n1201) );
  XNOR U1976 ( .A(n1626), .B(n1201), .Z(out[1096]) );
  XNOR U1977 ( .A(n1203), .B(n1202), .Z(n3639) );
  XNOR U1978 ( .A(in[902]), .B(n3639), .Z(n1628) );
  NOR U1979 ( .A(n1433), .B(n4666), .Z(n1204) );
  XNOR U1980 ( .A(n1628), .B(n1204), .Z(out[1097]) );
  XNOR U1981 ( .A(n1206), .B(n1205), .Z(n3643) );
  XNOR U1982 ( .A(in[903]), .B(n3643), .Z(n1630) );
  NOR U1983 ( .A(n1437), .B(n4674), .Z(n1207) );
  XNOR U1984 ( .A(n1630), .B(n1207), .Z(out[1098]) );
  XNOR U1985 ( .A(n1209), .B(n1208), .Z(n3647) );
  XNOR U1986 ( .A(in[904]), .B(n3647), .Z(n1632) );
  NOR U1987 ( .A(n1441), .B(n4678), .Z(n1210) );
  XNOR U1988 ( .A(n1632), .B(n1210), .Z(out[1099]) );
  XOR U1989 ( .A(in[580]), .B(n3631), .Z(n2568) );
  XOR U1990 ( .A(in[235]), .B(n3728), .Z(n2970) );
  XNOR U1991 ( .A(in[1455]), .B(n3769), .Z(n2967) );
  NAND U1992 ( .A(n2970), .B(n2967), .Z(n1211) );
  XNOR U1993 ( .A(n2568), .B(n1211), .Z(out[109]) );
  XOR U1994 ( .A(in[200]), .B(n3572), .Z(n3920) );
  XNOR U1995 ( .A(in[1420]), .B(n3613), .Z(n3919) );
  XOR U1996 ( .A(n4119), .B(in[1043]), .Z(n2631) );
  NAND U1997 ( .A(n3919), .B(n2631), .Z(n1212) );
  XNOR U1998 ( .A(n3920), .B(n1212), .Z(out[10]) );
  XNOR U1999 ( .A(n1214), .B(n1213), .Z(n3651) );
  XNOR U2000 ( .A(in[905]), .B(n3651), .Z(n1634) );
  NOR U2001 ( .A(n1445), .B(n4682), .Z(n1215) );
  XNOR U2002 ( .A(n1634), .B(n1215), .Z(out[1100]) );
  XNOR U2003 ( .A(n1217), .B(n1216), .Z(n3655) );
  XNOR U2004 ( .A(in[906]), .B(n3655), .Z(n1636) );
  NOR U2005 ( .A(n1449), .B(n4686), .Z(n1218) );
  XNOR U2006 ( .A(n1636), .B(n1218), .Z(out[1101]) );
  XNOR U2007 ( .A(n1220), .B(n1219), .Z(n3659) );
  XNOR U2008 ( .A(in[907]), .B(n3659), .Z(n1639) );
  NOR U2009 ( .A(n1453), .B(n4690), .Z(n1221) );
  XNOR U2010 ( .A(n1639), .B(n1221), .Z(out[1102]) );
  XNOR U2011 ( .A(n1223), .B(n1222), .Z(n3667) );
  XNOR U2012 ( .A(in[908]), .B(n3667), .Z(n1641) );
  NOR U2013 ( .A(n1457), .B(n4694), .Z(n1224) );
  XNOR U2014 ( .A(n1641), .B(n1224), .Z(out[1103]) );
  XOR U2015 ( .A(n1226), .B(n1225), .Z(n3671) );
  XNOR U2016 ( .A(in[909]), .B(n3671), .Z(n1643) );
  NOR U2017 ( .A(n1461), .B(n4698), .Z(n1227) );
  XNOR U2018 ( .A(n1643), .B(n1227), .Z(out[1104]) );
  XOR U2019 ( .A(n1229), .B(n1228), .Z(n3675) );
  XNOR U2020 ( .A(in[910]), .B(n3675), .Z(n1645) );
  NOR U2021 ( .A(n1465), .B(n4702), .Z(n1230) );
  XNOR U2022 ( .A(n1645), .B(n1230), .Z(out[1105]) );
  XOR U2023 ( .A(n1232), .B(n1231), .Z(n3679) );
  XNOR U2024 ( .A(in[911]), .B(n3679), .Z(n1647) );
  NOR U2025 ( .A(n1470), .B(n4706), .Z(n1233) );
  XNOR U2026 ( .A(n1647), .B(n1233), .Z(out[1106]) );
  XOR U2027 ( .A(n1235), .B(n1234), .Z(n3683) );
  XNOR U2028 ( .A(in[912]), .B(n3683), .Z(n1649) );
  NOR U2029 ( .A(n1474), .B(n4710), .Z(n1236) );
  XNOR U2030 ( .A(n1649), .B(n1236), .Z(out[1107]) );
  XNOR U2031 ( .A(n1238), .B(n1237), .Z(n3687) );
  XNOR U2032 ( .A(in[913]), .B(n3687), .Z(n1651) );
  NOR U2033 ( .A(n1478), .B(n4718), .Z(n1239) );
  XNOR U2034 ( .A(n1651), .B(n1239), .Z(out[1108]) );
  XOR U2035 ( .A(n1241), .B(n1240), .Z(n3691) );
  XNOR U2036 ( .A(in[914]), .B(n3691), .Z(n1653) );
  NOR U2037 ( .A(n1482), .B(n4722), .Z(n1242) );
  XNOR U2038 ( .A(n1653), .B(n1242), .Z(out[1109]) );
  XOR U2039 ( .A(in[581]), .B(n3635), .Z(n2570) );
  XOR U2040 ( .A(in[236]), .B(n3732), .Z(n2994) );
  XNOR U2041 ( .A(in[1456]), .B(n3773), .Z(n2991) );
  NAND U2042 ( .A(n2994), .B(n2991), .Z(n1243) );
  XNOR U2043 ( .A(n2570), .B(n1243), .Z(out[110]) );
  XNOR U2044 ( .A(n1245), .B(n1244), .Z(n3695) );
  XNOR U2045 ( .A(in[915]), .B(n3695), .Z(n1655) );
  NOR U2046 ( .A(n1486), .B(n4726), .Z(n1246) );
  XNOR U2047 ( .A(n1655), .B(n1246), .Z(out[1110]) );
  XNOR U2048 ( .A(n1248), .B(n1247), .Z(n3699) );
  XNOR U2049 ( .A(in[916]), .B(n3699), .Z(n1657) );
  NOR U2050 ( .A(n1490), .B(n4730), .Z(n1249) );
  XNOR U2051 ( .A(n1657), .B(n1249), .Z(out[1111]) );
  XNOR U2052 ( .A(n1251), .B(n1250), .Z(n3703) );
  XNOR U2053 ( .A(in[917]), .B(n3703), .Z(n1660) );
  NOR U2054 ( .A(n1494), .B(n4734), .Z(n1252) );
  XNOR U2055 ( .A(n1660), .B(n1252), .Z(out[1112]) );
  XNOR U2056 ( .A(n1254), .B(n1253), .Z(n3711) );
  XNOR U2057 ( .A(in[918]), .B(n3711), .Z(n1662) );
  NOR U2058 ( .A(n1498), .B(n4738), .Z(n1255) );
  XNOR U2059 ( .A(n1662), .B(n1255), .Z(out[1113]) );
  XOR U2060 ( .A(n1257), .B(n1256), .Z(n3715) );
  XNOR U2061 ( .A(in[919]), .B(n3715), .Z(n1664) );
  NOR U2062 ( .A(n1502), .B(n4742), .Z(n1258) );
  XNOR U2063 ( .A(n1664), .B(n1258), .Z(out[1114]) );
  XOR U2064 ( .A(n1260), .B(n1259), .Z(n3719) );
  XNOR U2065 ( .A(in[920]), .B(n3719), .Z(n1666) );
  NOR U2066 ( .A(n1506), .B(n4746), .Z(n1261) );
  XNOR U2067 ( .A(n1666), .B(n1261), .Z(out[1115]) );
  XNOR U2068 ( .A(n1263), .B(n1262), .Z(n3723) );
  XNOR U2069 ( .A(in[921]), .B(n3723), .Z(n1668) );
  NOR U2070 ( .A(n1511), .B(n4750), .Z(n1264) );
  XNOR U2071 ( .A(n1668), .B(n1264), .Z(out[1116]) );
  XOR U2072 ( .A(n1266), .B(n1265), .Z(n3727) );
  XNOR U2073 ( .A(in[922]), .B(n3727), .Z(n1670) );
  NOR U2074 ( .A(n1515), .B(n4754), .Z(n1267) );
  XNOR U2075 ( .A(n1670), .B(n1267), .Z(out[1117]) );
  XOR U2076 ( .A(n1269), .B(n1268), .Z(n3731) );
  XNOR U2077 ( .A(in[923]), .B(n3731), .Z(n1672) );
  NOR U2078 ( .A(n1519), .B(n4762), .Z(n1270) );
  XNOR U2079 ( .A(n1672), .B(n1270), .Z(out[1118]) );
  XOR U2080 ( .A(n1272), .B(n1271), .Z(n3735) );
  XNOR U2081 ( .A(in[924]), .B(n3735), .Z(n1674) );
  NOR U2082 ( .A(n1523), .B(n4766), .Z(n1273) );
  XNOR U2083 ( .A(n1674), .B(n1273), .Z(out[1119]) );
  XOR U2084 ( .A(in[582]), .B(n3639), .Z(n2572) );
  XOR U2085 ( .A(in[237]), .B(n3736), .Z(n3018) );
  XNOR U2086 ( .A(in[1457]), .B(n3777), .Z(n3015) );
  NAND U2087 ( .A(n3018), .B(n3015), .Z(n1274) );
  XNOR U2088 ( .A(n2572), .B(n1274), .Z(out[111]) );
  XOR U2089 ( .A(n1276), .B(n1275), .Z(n3739) );
  XNOR U2090 ( .A(in[925]), .B(n3739), .Z(n1676) );
  NOR U2091 ( .A(n1527), .B(n4770), .Z(n1277) );
  XNOR U2092 ( .A(n1676), .B(n1277), .Z(out[1120]) );
  XOR U2093 ( .A(n1279), .B(n1278), .Z(n3743) );
  XNOR U2094 ( .A(in[926]), .B(n3743), .Z(n1678) );
  NOR U2095 ( .A(n1531), .B(n4774), .Z(n1280) );
  XNOR U2096 ( .A(n1678), .B(n1280), .Z(out[1121]) );
  XOR U2097 ( .A(n1282), .B(n1281), .Z(n3747) );
  XNOR U2098 ( .A(in[927]), .B(n3747), .Z(n1681) );
  NOR U2099 ( .A(n1535), .B(n4778), .Z(n1283) );
  XNOR U2100 ( .A(n1681), .B(n1283), .Z(out[1122]) );
  XOR U2101 ( .A(n1285), .B(n1284), .Z(n3755) );
  XNOR U2102 ( .A(in[928]), .B(n3755), .Z(n1683) );
  NOR U2103 ( .A(n1539), .B(n4782), .Z(n1286) );
  XNOR U2104 ( .A(n1683), .B(n1286), .Z(out[1123]) );
  XNOR U2105 ( .A(n1288), .B(n1287), .Z(n3759) );
  XNOR U2106 ( .A(in[929]), .B(n3759), .Z(n1685) );
  NOR U2107 ( .A(n1543), .B(n4786), .Z(n1289) );
  XNOR U2108 ( .A(n1685), .B(n1289), .Z(out[1124]) );
  XOR U2109 ( .A(n1291), .B(n1290), .Z(n3763) );
  XNOR U2110 ( .A(in[930]), .B(n3763), .Z(n1687) );
  NOR U2111 ( .A(n1547), .B(n4790), .Z(n1292) );
  XNOR U2112 ( .A(n1687), .B(n1292), .Z(out[1125]) );
  XNOR U2113 ( .A(n1294), .B(n1293), .Z(n3767) );
  XNOR U2114 ( .A(in[931]), .B(n3767), .Z(n1689) );
  NOR U2115 ( .A(n1552), .B(n4794), .Z(n1295) );
  XNOR U2116 ( .A(n1689), .B(n1295), .Z(out[1126]) );
  XNOR U2117 ( .A(n1297), .B(n1296), .Z(n3771) );
  XNOR U2118 ( .A(in[932]), .B(n3771), .Z(n1691) );
  NOR U2119 ( .A(n1556), .B(n4798), .Z(n1298) );
  XNOR U2120 ( .A(n1691), .B(n1298), .Z(out[1127]) );
  XNOR U2121 ( .A(n1300), .B(n1299), .Z(n3775) );
  XNOR U2122 ( .A(in[933]), .B(n3775), .Z(n1694) );
  NAND U2123 ( .A(n1558), .B(n1301), .Z(n1302) );
  XNOR U2124 ( .A(n1694), .B(n1302), .Z(out[1128]) );
  XOR U2125 ( .A(n1304), .B(n1303), .Z(n3779) );
  XNOR U2126 ( .A(in[934]), .B(n3779), .Z(n1698) );
  NAND U2127 ( .A(n1560), .B(n1305), .Z(n1306) );
  XNOR U2128 ( .A(n1698), .B(n1306), .Z(out[1129]) );
  XOR U2129 ( .A(in[583]), .B(n3643), .Z(n2575) );
  XOR U2130 ( .A(in[238]), .B(n3740), .Z(n3042) );
  XNOR U2131 ( .A(in[1458]), .B(n3781), .Z(n3039) );
  NAND U2132 ( .A(n3042), .B(n3039), .Z(n1307) );
  XNOR U2133 ( .A(n2575), .B(n1307), .Z(out[112]) );
  XNOR U2134 ( .A(n1309), .B(n1308), .Z(n3783) );
  XNOR U2135 ( .A(in[935]), .B(n3783), .Z(n1702) );
  NAND U2136 ( .A(n1562), .B(n1310), .Z(n1311) );
  XNOR U2137 ( .A(n1702), .B(n1311), .Z(out[1130]) );
  XNOR U2138 ( .A(n1313), .B(n1312), .Z(n3787) );
  XNOR U2139 ( .A(in[936]), .B(n3787), .Z(n1706) );
  NAND U2140 ( .A(n1564), .B(n1314), .Z(n1315) );
  XNOR U2141 ( .A(n1706), .B(n1315), .Z(out[1131]) );
  XNOR U2142 ( .A(n1317), .B(n1316), .Z(n3791) );
  XNOR U2143 ( .A(in[937]), .B(n3791), .Z(n1711) );
  NAND U2144 ( .A(n1566), .B(n1318), .Z(n1319) );
  XNOR U2145 ( .A(n1711), .B(n1319), .Z(out[1132]) );
  XNOR U2146 ( .A(n1321), .B(n1320), .Z(n3801) );
  XNOR U2147 ( .A(in[938]), .B(n3801), .Z(n1715) );
  NAND U2148 ( .A(n1568), .B(n1322), .Z(n1323) );
  XNOR U2149 ( .A(n1715), .B(n1323), .Z(out[1133]) );
  XNOR U2150 ( .A(n1325), .B(n1324), .Z(n3805) );
  XNOR U2151 ( .A(in[939]), .B(n3805), .Z(n1719) );
  NAND U2152 ( .A(n1570), .B(n1326), .Z(n1327) );
  XNOR U2153 ( .A(n1719), .B(n1327), .Z(out[1134]) );
  XNOR U2154 ( .A(n1329), .B(n1328), .Z(n3809) );
  XNOR U2155 ( .A(in[940]), .B(n3809), .Z(n1723) );
  NAND U2156 ( .A(n1572), .B(n1330), .Z(n1331) );
  XNOR U2157 ( .A(n1723), .B(n1331), .Z(out[1135]) );
  XNOR U2158 ( .A(n1333), .B(n1332), .Z(n3813) );
  XNOR U2159 ( .A(in[941]), .B(n3813), .Z(n1727) );
  NAND U2160 ( .A(n1576), .B(n1334), .Z(n1335) );
  XNOR U2161 ( .A(n1727), .B(n1335), .Z(out[1136]) );
  XNOR U2162 ( .A(n1337), .B(n1336), .Z(n3535) );
  XNOR U2163 ( .A(in[942]), .B(n3535), .Z(n1731) );
  NAND U2164 ( .A(n1578), .B(n1338), .Z(n1339) );
  XNOR U2165 ( .A(n1731), .B(n1339), .Z(out[1137]) );
  XNOR U2166 ( .A(n1341), .B(n1340), .Z(n3539) );
  XNOR U2167 ( .A(in[943]), .B(n3539), .Z(n1735) );
  NAND U2168 ( .A(n1580), .B(n1342), .Z(n1343) );
  XNOR U2169 ( .A(n1735), .B(n1343), .Z(out[1138]) );
  XNOR U2170 ( .A(n1345), .B(n1344), .Z(n3543) );
  XNOR U2171 ( .A(in[944]), .B(n3543), .Z(n1739) );
  NAND U2172 ( .A(n1582), .B(n1346), .Z(n1347) );
  XNOR U2173 ( .A(n1739), .B(n1347), .Z(out[1139]) );
  XOR U2174 ( .A(in[584]), .B(n3647), .Z(n2577) );
  XOR U2175 ( .A(in[239]), .B(n3744), .Z(n3066) );
  XNOR U2176 ( .A(in[1459]), .B(n3785), .Z(n3063) );
  NAND U2177 ( .A(n3066), .B(n3063), .Z(n1348) );
  XNOR U2178 ( .A(n2577), .B(n1348), .Z(out[113]) );
  XNOR U2179 ( .A(n1350), .B(n1349), .Z(n3547) );
  XNOR U2180 ( .A(in[945]), .B(n3547), .Z(n1743) );
  NAND U2181 ( .A(n1584), .B(n1351), .Z(n1352) );
  XNOR U2182 ( .A(n1743), .B(n1352), .Z(out[1140]) );
  XNOR U2183 ( .A(n1354), .B(n1353), .Z(n3551) );
  XNOR U2184 ( .A(in[946]), .B(n3551), .Z(n1747) );
  NAND U2185 ( .A(n1586), .B(n1355), .Z(n1356) );
  XNOR U2186 ( .A(n1747), .B(n1356), .Z(out[1141]) );
  XNOR U2187 ( .A(n1358), .B(n1357), .Z(n3555) );
  XNOR U2188 ( .A(in[947]), .B(n3555), .Z(n1752) );
  NAND U2189 ( .A(n1588), .B(n1359), .Z(n1360) );
  XNOR U2190 ( .A(n1752), .B(n1360), .Z(out[1142]) );
  XNOR U2191 ( .A(n1362), .B(n1361), .Z(n3559) );
  XNOR U2192 ( .A(in[948]), .B(n3559), .Z(n1756) );
  NAND U2193 ( .A(n1590), .B(n1363), .Z(n1364) );
  XNOR U2194 ( .A(n1756), .B(n1364), .Z(out[1143]) );
  XNOR U2195 ( .A(n1366), .B(n1365), .Z(n3563) );
  XNOR U2196 ( .A(in[949]), .B(n3563), .Z(n1760) );
  NAND U2197 ( .A(n1592), .B(n1367), .Z(n1368) );
  XNOR U2198 ( .A(n1760), .B(n1368), .Z(out[1144]) );
  XNOR U2199 ( .A(n1370), .B(n1369), .Z(n3567) );
  XNOR U2200 ( .A(in[950]), .B(n3567), .Z(n1764) );
  NAND U2201 ( .A(n1594), .B(n1371), .Z(n1372) );
  XNOR U2202 ( .A(n1764), .B(n1372), .Z(out[1145]) );
  XNOR U2203 ( .A(n1374), .B(n1373), .Z(n3571) );
  XNOR U2204 ( .A(in[951]), .B(n3571), .Z(n1768) );
  NAND U2205 ( .A(n1597), .B(n1375), .Z(n1376) );
  XNOR U2206 ( .A(n1768), .B(n1376), .Z(out[1146]) );
  XNOR U2207 ( .A(n1378), .B(n1377), .Z(n3579) );
  XNOR U2208 ( .A(in[952]), .B(n3579), .Z(n1772) );
  NAND U2209 ( .A(n1599), .B(n1379), .Z(n1380) );
  XNOR U2210 ( .A(n1772), .B(n1380), .Z(out[1147]) );
  XNOR U2211 ( .A(n1382), .B(n1381), .Z(n3583) );
  XNOR U2212 ( .A(in[953]), .B(n3583), .Z(n1776) );
  NAND U2213 ( .A(n1601), .B(n1383), .Z(n1384) );
  XNOR U2214 ( .A(n1776), .B(n1384), .Z(out[1148]) );
  XNOR U2215 ( .A(n1386), .B(n1385), .Z(n3587) );
  XNOR U2216 ( .A(in[954]), .B(n3587), .Z(n1780) );
  NAND U2217 ( .A(n1603), .B(n1387), .Z(n1388) );
  XNOR U2218 ( .A(n1780), .B(n1388), .Z(out[1149]) );
  XOR U2219 ( .A(in[585]), .B(n3651), .Z(n2579) );
  XOR U2220 ( .A(in[240]), .B(n3748), .Z(n3092) );
  XNOR U2221 ( .A(in[1460]), .B(n3789), .Z(n3089) );
  NAND U2222 ( .A(n3092), .B(n3089), .Z(n1389) );
  XNOR U2223 ( .A(n2579), .B(n1389), .Z(out[114]) );
  XNOR U2224 ( .A(in[955]), .B(n3591), .Z(n1784) );
  NAND U2225 ( .A(n1605), .B(n1390), .Z(n1391) );
  XNOR U2226 ( .A(n1784), .B(n1391), .Z(out[1150]) );
  XNOR U2227 ( .A(in[956]), .B(n3595), .Z(n1788) );
  NAND U2228 ( .A(n1607), .B(n1392), .Z(n1393) );
  XNOR U2229 ( .A(n1788), .B(n1393), .Z(out[1151]) );
  XNOR U2230 ( .A(n1395), .B(n1394), .Z(n3935) );
  XNOR U2231 ( .A(in[1004]), .B(n3935), .Z(n4628) );
  NAND U2232 ( .A(n1609), .B(n1396), .Z(n1397) );
  XNOR U2233 ( .A(n4628), .B(n1397), .Z(out[1152]) );
  XNOR U2234 ( .A(n1399), .B(n1398), .Z(n3937) );
  XNOR U2235 ( .A(in[1005]), .B(n3937), .Z(n4632) );
  NAND U2236 ( .A(n1611), .B(n1400), .Z(n1401) );
  XNOR U2237 ( .A(n4632), .B(n1401), .Z(out[1153]) );
  XNOR U2238 ( .A(n1403), .B(n1402), .Z(n3939) );
  XNOR U2239 ( .A(in[1006]), .B(n3939), .Z(n4636) );
  NAND U2240 ( .A(n1613), .B(n1404), .Z(n1405) );
  XNOR U2241 ( .A(n4636), .B(n1405), .Z(out[1154]) );
  XNOR U2242 ( .A(n1407), .B(n1406), .Z(n3941) );
  XNOR U2243 ( .A(in[1007]), .B(n3941), .Z(n4640) );
  NAND U2244 ( .A(n1615), .B(n1408), .Z(n1409) );
  XNOR U2245 ( .A(n4640), .B(n1409), .Z(out[1155]) );
  XNOR U2246 ( .A(n1411), .B(n1410), .Z(n3947) );
  XNOR U2247 ( .A(in[1008]), .B(n3947), .Z(n4644) );
  NAND U2248 ( .A(n1618), .B(n1412), .Z(n1413) );
  XNOR U2249 ( .A(n4644), .B(n1413), .Z(out[1156]) );
  XNOR U2250 ( .A(n1415), .B(n1414), .Z(n3949) );
  XNOR U2251 ( .A(in[1009]), .B(n3949), .Z(n4648) );
  NAND U2252 ( .A(n1620), .B(n1416), .Z(n1417) );
  XNOR U2253 ( .A(n4648), .B(n1417), .Z(out[1157]) );
  XNOR U2254 ( .A(n1419), .B(n1418), .Z(n3951) );
  XNOR U2255 ( .A(in[1010]), .B(n3951), .Z(n4652) );
  NAND U2256 ( .A(n1622), .B(n1420), .Z(n1421) );
  XNOR U2257 ( .A(n4652), .B(n1421), .Z(out[1158]) );
  XNOR U2258 ( .A(n1423), .B(n1422), .Z(n3953) );
  XNOR U2259 ( .A(in[1011]), .B(n3953), .Z(n4656) );
  NAND U2260 ( .A(n1624), .B(n1424), .Z(n1425) );
  XNOR U2261 ( .A(n4656), .B(n1425), .Z(out[1159]) );
  XOR U2262 ( .A(in[586]), .B(n3655), .Z(n2581) );
  XOR U2263 ( .A(in[241]), .B(n3756), .Z(n3116) );
  XNOR U2264 ( .A(in[1461]), .B(n3793), .Z(n3113) );
  NAND U2265 ( .A(n3116), .B(n3113), .Z(n1426) );
  XNOR U2266 ( .A(n2581), .B(n1426), .Z(out[115]) );
  XNOR U2267 ( .A(n1428), .B(n1427), .Z(n3955) );
  XNOR U2268 ( .A(in[1012]), .B(n3955), .Z(n4660) );
  NAND U2269 ( .A(n1626), .B(n1429), .Z(n1430) );
  XNOR U2270 ( .A(n4660), .B(n1430), .Z(out[1160]) );
  XNOR U2271 ( .A(n1432), .B(n1431), .Z(n3957) );
  XNOR U2272 ( .A(in[1013]), .B(n3957), .Z(n4664) );
  NAND U2273 ( .A(n1628), .B(n1433), .Z(n1434) );
  XNOR U2274 ( .A(n4664), .B(n1434), .Z(out[1161]) );
  XNOR U2275 ( .A(n1436), .B(n1435), .Z(n3959) );
  XNOR U2276 ( .A(in[1014]), .B(n3959), .Z(n4672) );
  NAND U2277 ( .A(n1630), .B(n1437), .Z(n1438) );
  XNOR U2278 ( .A(n4672), .B(n1438), .Z(out[1162]) );
  XNOR U2279 ( .A(n1440), .B(n1439), .Z(n3961) );
  XNOR U2280 ( .A(in[1015]), .B(n3961), .Z(n4676) );
  NAND U2281 ( .A(n1632), .B(n1441), .Z(n1442) );
  XNOR U2282 ( .A(n4676), .B(n1442), .Z(out[1163]) );
  XNOR U2283 ( .A(n1444), .B(n1443), .Z(n3817) );
  XNOR U2284 ( .A(in[1016]), .B(n3817), .Z(n4680) );
  NAND U2285 ( .A(n1634), .B(n1445), .Z(n1446) );
  XNOR U2286 ( .A(n4680), .B(n1446), .Z(out[1164]) );
  XNOR U2287 ( .A(n1448), .B(n1447), .Z(n3819) );
  XNOR U2288 ( .A(in[1017]), .B(n3819), .Z(n4684) );
  NAND U2289 ( .A(n1636), .B(n1449), .Z(n1450) );
  XNOR U2290 ( .A(n4684), .B(n1450), .Z(out[1165]) );
  XNOR U2291 ( .A(n1452), .B(n1451), .Z(n3821) );
  XNOR U2292 ( .A(in[1018]), .B(n3821), .Z(n4688) );
  NAND U2293 ( .A(n1639), .B(n1453), .Z(n1454) );
  XNOR U2294 ( .A(n4688), .B(n1454), .Z(out[1166]) );
  XNOR U2295 ( .A(n1456), .B(n1455), .Z(n3823) );
  XNOR U2296 ( .A(in[1019]), .B(n3823), .Z(n4692) );
  NAND U2297 ( .A(n1641), .B(n1457), .Z(n1458) );
  XNOR U2298 ( .A(n4692), .B(n1458), .Z(out[1167]) );
  XOR U2299 ( .A(n1460), .B(n1459), .Z(n3825) );
  XNOR U2300 ( .A(in[1020]), .B(n3825), .Z(n4696) );
  NAND U2301 ( .A(n1643), .B(n1461), .Z(n1462) );
  XNOR U2302 ( .A(n4696), .B(n1462), .Z(out[1168]) );
  XOR U2303 ( .A(n1464), .B(n1463), .Z(n3827) );
  XNOR U2304 ( .A(in[1021]), .B(n3827), .Z(n4700) );
  NAND U2305 ( .A(n1645), .B(n1465), .Z(n1466) );
  XNOR U2306 ( .A(n4700), .B(n1466), .Z(out[1169]) );
  XOR U2307 ( .A(in[587]), .B(n3659), .Z(n2583) );
  XOR U2308 ( .A(in[242]), .B(n3760), .Z(n3140) );
  XNOR U2309 ( .A(in[1462]), .B(n3803), .Z(n3137) );
  NAND U2310 ( .A(n3140), .B(n3137), .Z(n1467) );
  XNOR U2311 ( .A(n2583), .B(n1467), .Z(out[116]) );
  XOR U2312 ( .A(n1469), .B(n1468), .Z(n3833) );
  XNOR U2313 ( .A(in[1022]), .B(n3833), .Z(n4704) );
  NAND U2314 ( .A(n1647), .B(n1470), .Z(n1471) );
  XNOR U2315 ( .A(n4704), .B(n1471), .Z(out[1170]) );
  XNOR U2316 ( .A(n1473), .B(n1472), .Z(n3835) );
  XNOR U2317 ( .A(in[1023]), .B(n3835), .Z(n4708) );
  NAND U2318 ( .A(n1649), .B(n1474), .Z(n1475) );
  XNOR U2319 ( .A(n4708), .B(n1475), .Z(out[1171]) );
  XOR U2320 ( .A(n1477), .B(n1476), .Z(n3837) );
  XNOR U2321 ( .A(in[960]), .B(n3837), .Z(n4716) );
  NAND U2322 ( .A(n1651), .B(n1478), .Z(n1479) );
  XNOR U2323 ( .A(n4716), .B(n1479), .Z(out[1172]) );
  XOR U2324 ( .A(n1481), .B(n1480), .Z(n3839) );
  XNOR U2325 ( .A(in[961]), .B(n3839), .Z(n4720) );
  NAND U2326 ( .A(n1653), .B(n1482), .Z(n1483) );
  XNOR U2327 ( .A(n4720), .B(n1483), .Z(out[1173]) );
  XOR U2328 ( .A(n1485), .B(n1484), .Z(n3841) );
  XNOR U2329 ( .A(in[962]), .B(n3841), .Z(n4724) );
  NAND U2330 ( .A(n1655), .B(n1486), .Z(n1487) );
  XNOR U2331 ( .A(n4724), .B(n1487), .Z(out[1174]) );
  XOR U2332 ( .A(n1489), .B(n1488), .Z(n3843) );
  XNOR U2333 ( .A(in[963]), .B(n3843), .Z(n4728) );
  NAND U2334 ( .A(n1657), .B(n1490), .Z(n1491) );
  XNOR U2335 ( .A(n4728), .B(n1491), .Z(out[1175]) );
  XOR U2336 ( .A(n1493), .B(n1492), .Z(n3845) );
  XNOR U2337 ( .A(in[964]), .B(n3845), .Z(n4732) );
  NAND U2338 ( .A(n1660), .B(n1494), .Z(n1495) );
  XNOR U2339 ( .A(n4732), .B(n1495), .Z(out[1176]) );
  XOR U2340 ( .A(n1497), .B(n1496), .Z(n3847) );
  XNOR U2341 ( .A(in[965]), .B(n3847), .Z(n4736) );
  NAND U2342 ( .A(n1662), .B(n1498), .Z(n1499) );
  XNOR U2343 ( .A(n4736), .B(n1499), .Z(out[1177]) );
  XOR U2344 ( .A(n1501), .B(n1500), .Z(n3849) );
  XNOR U2345 ( .A(in[966]), .B(n3849), .Z(n4740) );
  NAND U2346 ( .A(n1664), .B(n1502), .Z(n1503) );
  XNOR U2347 ( .A(n4740), .B(n1503), .Z(out[1178]) );
  XOR U2348 ( .A(n1505), .B(n1504), .Z(n3851) );
  XNOR U2349 ( .A(in[967]), .B(n3851), .Z(n4744) );
  NAND U2350 ( .A(n1666), .B(n1506), .Z(n1507) );
  XNOR U2351 ( .A(n4744), .B(n1507), .Z(out[1179]) );
  XOR U2352 ( .A(in[588]), .B(n3667), .Z(n2585) );
  XOR U2353 ( .A(in[243]), .B(n3764), .Z(n3164) );
  XNOR U2354 ( .A(in[1463]), .B(n3807), .Z(n3161) );
  NAND U2355 ( .A(n3164), .B(n3161), .Z(n1508) );
  XNOR U2356 ( .A(n2585), .B(n1508), .Z(out[117]) );
  XOR U2357 ( .A(n1510), .B(n1509), .Z(n3855) );
  XNOR U2358 ( .A(in[968]), .B(n3855), .Z(n4748) );
  NAND U2359 ( .A(n1668), .B(n1511), .Z(n1512) );
  XNOR U2360 ( .A(n4748), .B(n1512), .Z(out[1180]) );
  XOR U2361 ( .A(n1514), .B(n1513), .Z(n3857) );
  XNOR U2362 ( .A(in[969]), .B(n3857), .Z(n4752) );
  NAND U2363 ( .A(n1670), .B(n1515), .Z(n1516) );
  XNOR U2364 ( .A(n4752), .B(n1516), .Z(out[1181]) );
  XOR U2365 ( .A(n1518), .B(n1517), .Z(n3859) );
  XNOR U2366 ( .A(in[970]), .B(n3859), .Z(n4760) );
  NAND U2367 ( .A(n1672), .B(n1519), .Z(n1520) );
  XNOR U2368 ( .A(n4760), .B(n1520), .Z(out[1182]) );
  XOR U2369 ( .A(n1522), .B(n1521), .Z(n3861) );
  XNOR U2370 ( .A(in[971]), .B(n3861), .Z(n4764) );
  NAND U2371 ( .A(n1674), .B(n1523), .Z(n1524) );
  XNOR U2372 ( .A(n4764), .B(n1524), .Z(out[1183]) );
  XOR U2373 ( .A(n1526), .B(n1525), .Z(n3863) );
  XNOR U2374 ( .A(in[972]), .B(n3863), .Z(n4768) );
  NAND U2375 ( .A(n1676), .B(n1527), .Z(n1528) );
  XNOR U2376 ( .A(n4768), .B(n1528), .Z(out[1184]) );
  XOR U2377 ( .A(n1530), .B(n1529), .Z(n3865) );
  XNOR U2378 ( .A(in[973]), .B(n3865), .Z(n4772) );
  NAND U2379 ( .A(n1678), .B(n1531), .Z(n1532) );
  XNOR U2380 ( .A(n4772), .B(n1532), .Z(out[1185]) );
  XNOR U2381 ( .A(n1534), .B(n1533), .Z(n3867) );
  XNOR U2382 ( .A(in[974]), .B(n3867), .Z(n4776) );
  NAND U2383 ( .A(n1681), .B(n1535), .Z(n1536) );
  XNOR U2384 ( .A(n4776), .B(n1536), .Z(out[1186]) );
  XNOR U2385 ( .A(n1538), .B(n1537), .Z(n3869) );
  XNOR U2386 ( .A(in[975]), .B(n3869), .Z(n4780) );
  NAND U2387 ( .A(n1683), .B(n1539), .Z(n1540) );
  XNOR U2388 ( .A(n4780), .B(n1540), .Z(out[1187]) );
  XOR U2389 ( .A(n1542), .B(n1541), .Z(n3871) );
  XNOR U2390 ( .A(in[976]), .B(n3871), .Z(n4784) );
  NAND U2391 ( .A(n1685), .B(n1543), .Z(n1544) );
  XNOR U2392 ( .A(n4784), .B(n1544), .Z(out[1188]) );
  XOR U2393 ( .A(n1546), .B(n1545), .Z(n3873) );
  XNOR U2394 ( .A(in[977]), .B(n3873), .Z(n4788) );
  NAND U2395 ( .A(n1687), .B(n1547), .Z(n1548) );
  XNOR U2396 ( .A(n4788), .B(n1548), .Z(out[1189]) );
  XOR U2397 ( .A(in[589]), .B(n3671), .Z(n2587) );
  XOR U2398 ( .A(in[244]), .B(n3768), .Z(n3188) );
  XNOR U2399 ( .A(in[1464]), .B(n3811), .Z(n3185) );
  NAND U2400 ( .A(n3188), .B(n3185), .Z(n1549) );
  XNOR U2401 ( .A(n2587), .B(n1549), .Z(out[118]) );
  XOR U2402 ( .A(n1551), .B(n1550), .Z(n3877) );
  XNOR U2403 ( .A(in[978]), .B(n3877), .Z(n4792) );
  NAND U2404 ( .A(n1689), .B(n1552), .Z(n1553) );
  XNOR U2405 ( .A(n4792), .B(n1553), .Z(out[1190]) );
  XOR U2406 ( .A(n1555), .B(n1554), .Z(n3879) );
  XNOR U2407 ( .A(in[979]), .B(n3879), .Z(n4796) );
  NAND U2408 ( .A(n1691), .B(n1556), .Z(n1557) );
  XNOR U2409 ( .A(n4796), .B(n1557), .Z(out[1191]) );
  OR U2410 ( .A(n1694), .B(n1558), .Z(n1559) );
  XNOR U2411 ( .A(n1693), .B(n1559), .Z(out[1192]) );
  OR U2412 ( .A(n1698), .B(n1560), .Z(n1561) );
  XNOR U2413 ( .A(n1697), .B(n1561), .Z(out[1193]) );
  OR U2414 ( .A(n1702), .B(n1562), .Z(n1563) );
  XNOR U2415 ( .A(n1701), .B(n1563), .Z(out[1194]) );
  OR U2416 ( .A(n1706), .B(n1564), .Z(n1565) );
  XNOR U2417 ( .A(n1705), .B(n1565), .Z(out[1195]) );
  OR U2418 ( .A(n1711), .B(n1566), .Z(n1567) );
  XNOR U2419 ( .A(n1710), .B(n1567), .Z(out[1196]) );
  OR U2420 ( .A(n1715), .B(n1568), .Z(n1569) );
  XNOR U2421 ( .A(n1714), .B(n1569), .Z(out[1197]) );
  OR U2422 ( .A(n1719), .B(n1570), .Z(n1571) );
  XNOR U2423 ( .A(n1718), .B(n1571), .Z(out[1198]) );
  OR U2424 ( .A(n1723), .B(n1572), .Z(n1573) );
  XNOR U2425 ( .A(n1722), .B(n1573), .Z(out[1199]) );
  XOR U2426 ( .A(in[590]), .B(n3675), .Z(n2589) );
  XOR U2427 ( .A(in[245]), .B(n3772), .Z(n3212) );
  XNOR U2428 ( .A(in[1465]), .B(n3815), .Z(n3209) );
  NAND U2429 ( .A(n3212), .B(n3209), .Z(n1574) );
  XNOR U2430 ( .A(n2589), .B(n1574), .Z(out[119]) );
  XOR U2431 ( .A(in[201]), .B(n3580), .Z(n3944) );
  XNOR U2432 ( .A(in[1421]), .B(n3617), .Z(n3943) );
  XOR U2433 ( .A(in[1044]), .B(n4122), .Z(n2634) );
  NAND U2434 ( .A(n3943), .B(n2634), .Z(n1575) );
  XNOR U2435 ( .A(n3944), .B(n1575), .Z(out[11]) );
  OR U2436 ( .A(n1727), .B(n1576), .Z(n1577) );
  XNOR U2437 ( .A(n1726), .B(n1577), .Z(out[1200]) );
  OR U2438 ( .A(n1731), .B(n1578), .Z(n1579) );
  XNOR U2439 ( .A(n1730), .B(n1579), .Z(out[1201]) );
  OR U2440 ( .A(n1735), .B(n1580), .Z(n1581) );
  XNOR U2441 ( .A(n1734), .B(n1581), .Z(out[1202]) );
  OR U2442 ( .A(n1739), .B(n1582), .Z(n1583) );
  XNOR U2443 ( .A(n1738), .B(n1583), .Z(out[1203]) );
  OR U2444 ( .A(n1743), .B(n1584), .Z(n1585) );
  XNOR U2445 ( .A(n1742), .B(n1585), .Z(out[1204]) );
  OR U2446 ( .A(n1747), .B(n1586), .Z(n1587) );
  XNOR U2447 ( .A(n1746), .B(n1587), .Z(out[1205]) );
  OR U2448 ( .A(n1752), .B(n1588), .Z(n1589) );
  XNOR U2449 ( .A(n1751), .B(n1589), .Z(out[1206]) );
  OR U2450 ( .A(n1756), .B(n1590), .Z(n1591) );
  XNOR U2451 ( .A(n1755), .B(n1591), .Z(out[1207]) );
  OR U2452 ( .A(n1760), .B(n1592), .Z(n1593) );
  XNOR U2453 ( .A(n1759), .B(n1593), .Z(out[1208]) );
  OR U2454 ( .A(n1764), .B(n1594), .Z(n1595) );
  XNOR U2455 ( .A(n1763), .B(n1595), .Z(out[1209]) );
  XOR U2456 ( .A(in[591]), .B(n3679), .Z(n2591) );
  XOR U2457 ( .A(in[246]), .B(n3776), .Z(n3236) );
  XNOR U2458 ( .A(in[1466]), .B(n3537), .Z(n3233) );
  NAND U2459 ( .A(n3236), .B(n3233), .Z(n1596) );
  XNOR U2460 ( .A(n2591), .B(n1596), .Z(out[120]) );
  OR U2461 ( .A(n1768), .B(n1597), .Z(n1598) );
  XNOR U2462 ( .A(n1767), .B(n1598), .Z(out[1210]) );
  OR U2463 ( .A(n1772), .B(n1599), .Z(n1600) );
  XNOR U2464 ( .A(n1771), .B(n1600), .Z(out[1211]) );
  OR U2465 ( .A(n1776), .B(n1601), .Z(n1602) );
  XNOR U2466 ( .A(n1775), .B(n1602), .Z(out[1212]) );
  OR U2467 ( .A(n1780), .B(n1603), .Z(n1604) );
  XNOR U2468 ( .A(n1779), .B(n1604), .Z(out[1213]) );
  OR U2469 ( .A(n1784), .B(n1605), .Z(n1606) );
  XNOR U2470 ( .A(n1783), .B(n1606), .Z(out[1214]) );
  OR U2471 ( .A(n1788), .B(n1607), .Z(n1608) );
  XNOR U2472 ( .A(n1787), .B(n1608), .Z(out[1215]) );
  OR U2473 ( .A(n4628), .B(n1609), .Z(n1610) );
  XNOR U2474 ( .A(n4627), .B(n1610), .Z(out[1216]) );
  OR U2475 ( .A(n4632), .B(n1611), .Z(n1612) );
  XNOR U2476 ( .A(n4631), .B(n1612), .Z(out[1217]) );
  OR U2477 ( .A(n4636), .B(n1613), .Z(n1614) );
  XNOR U2478 ( .A(n4635), .B(n1614), .Z(out[1218]) );
  OR U2479 ( .A(n4640), .B(n1615), .Z(n1616) );
  XNOR U2480 ( .A(n4639), .B(n1616), .Z(out[1219]) );
  XOR U2481 ( .A(in[592]), .B(n3683), .Z(n2593) );
  XOR U2482 ( .A(in[247]), .B(n3780), .Z(n3268) );
  XNOR U2483 ( .A(in[1467]), .B(n3541), .Z(n3265) );
  NAND U2484 ( .A(n3268), .B(n3265), .Z(n1617) );
  XNOR U2485 ( .A(n2593), .B(n1617), .Z(out[121]) );
  OR U2486 ( .A(n4644), .B(n1618), .Z(n1619) );
  XNOR U2487 ( .A(n4643), .B(n1619), .Z(out[1220]) );
  OR U2488 ( .A(n4648), .B(n1620), .Z(n1621) );
  XNOR U2489 ( .A(n4647), .B(n1621), .Z(out[1221]) );
  OR U2490 ( .A(n4652), .B(n1622), .Z(n1623) );
  XNOR U2491 ( .A(n4651), .B(n1623), .Z(out[1222]) );
  OR U2492 ( .A(n4656), .B(n1624), .Z(n1625) );
  XNOR U2493 ( .A(n4655), .B(n1625), .Z(out[1223]) );
  OR U2494 ( .A(n4660), .B(n1626), .Z(n1627) );
  XNOR U2495 ( .A(n4659), .B(n1627), .Z(out[1224]) );
  OR U2496 ( .A(n4664), .B(n1628), .Z(n1629) );
  XNOR U2497 ( .A(n4663), .B(n1629), .Z(out[1225]) );
  OR U2498 ( .A(n4672), .B(n1630), .Z(n1631) );
  XNOR U2499 ( .A(n4671), .B(n1631), .Z(out[1226]) );
  OR U2500 ( .A(n4676), .B(n1632), .Z(n1633) );
  XNOR U2501 ( .A(n4675), .B(n1633), .Z(out[1227]) );
  OR U2502 ( .A(n4680), .B(n1634), .Z(n1635) );
  XNOR U2503 ( .A(n4679), .B(n1635), .Z(out[1228]) );
  OR U2504 ( .A(n4684), .B(n1636), .Z(n1637) );
  XNOR U2505 ( .A(n4683), .B(n1637), .Z(out[1229]) );
  XOR U2506 ( .A(in[593]), .B(n3687), .Z(n2596) );
  XOR U2507 ( .A(in[248]), .B(n3784), .Z(n3312) );
  XNOR U2508 ( .A(in[1468]), .B(n3545), .Z(n3309) );
  NAND U2509 ( .A(n3312), .B(n3309), .Z(n1638) );
  XNOR U2510 ( .A(n2596), .B(n1638), .Z(out[122]) );
  OR U2511 ( .A(n4688), .B(n1639), .Z(n1640) );
  XNOR U2512 ( .A(n4687), .B(n1640), .Z(out[1230]) );
  OR U2513 ( .A(n4692), .B(n1641), .Z(n1642) );
  XNOR U2514 ( .A(n4691), .B(n1642), .Z(out[1231]) );
  OR U2515 ( .A(n4696), .B(n1643), .Z(n1644) );
  XNOR U2516 ( .A(n4695), .B(n1644), .Z(out[1232]) );
  OR U2517 ( .A(n4700), .B(n1645), .Z(n1646) );
  XNOR U2518 ( .A(n4699), .B(n1646), .Z(out[1233]) );
  OR U2519 ( .A(n4704), .B(n1647), .Z(n1648) );
  XNOR U2520 ( .A(n4703), .B(n1648), .Z(out[1234]) );
  OR U2521 ( .A(n4708), .B(n1649), .Z(n1650) );
  XNOR U2522 ( .A(n4707), .B(n1650), .Z(out[1235]) );
  OR U2523 ( .A(n4716), .B(n1651), .Z(n1652) );
  XNOR U2524 ( .A(n4715), .B(n1652), .Z(out[1236]) );
  OR U2525 ( .A(n4720), .B(n1653), .Z(n1654) );
  XNOR U2526 ( .A(n4719), .B(n1654), .Z(out[1237]) );
  OR U2527 ( .A(n4724), .B(n1655), .Z(n1656) );
  XNOR U2528 ( .A(n4723), .B(n1656), .Z(out[1238]) );
  OR U2529 ( .A(n4728), .B(n1657), .Z(n1658) );
  XNOR U2530 ( .A(n4727), .B(n1658), .Z(out[1239]) );
  XOR U2531 ( .A(in[594]), .B(n3691), .Z(n2598) );
  XOR U2532 ( .A(in[249]), .B(n3788), .Z(n3356) );
  XNOR U2533 ( .A(in[1469]), .B(n3549), .Z(n3353) );
  NAND U2534 ( .A(n3356), .B(n3353), .Z(n1659) );
  XNOR U2535 ( .A(n2598), .B(n1659), .Z(out[123]) );
  OR U2536 ( .A(n4732), .B(n1660), .Z(n1661) );
  XNOR U2537 ( .A(n4731), .B(n1661), .Z(out[1240]) );
  OR U2538 ( .A(n4736), .B(n1662), .Z(n1663) );
  XNOR U2539 ( .A(n4735), .B(n1663), .Z(out[1241]) );
  OR U2540 ( .A(n4740), .B(n1664), .Z(n1665) );
  XNOR U2541 ( .A(n4739), .B(n1665), .Z(out[1242]) );
  OR U2542 ( .A(n4744), .B(n1666), .Z(n1667) );
  XNOR U2543 ( .A(n4743), .B(n1667), .Z(out[1243]) );
  OR U2544 ( .A(n4748), .B(n1668), .Z(n1669) );
  XNOR U2545 ( .A(n4747), .B(n1669), .Z(out[1244]) );
  OR U2546 ( .A(n4752), .B(n1670), .Z(n1671) );
  XNOR U2547 ( .A(n4751), .B(n1671), .Z(out[1245]) );
  OR U2548 ( .A(n4760), .B(n1672), .Z(n1673) );
  XNOR U2549 ( .A(n4759), .B(n1673), .Z(out[1246]) );
  OR U2550 ( .A(n4764), .B(n1674), .Z(n1675) );
  XNOR U2551 ( .A(n4763), .B(n1675), .Z(out[1247]) );
  OR U2552 ( .A(n4768), .B(n1676), .Z(n1677) );
  XNOR U2553 ( .A(n4767), .B(n1677), .Z(out[1248]) );
  OR U2554 ( .A(n4772), .B(n1678), .Z(n1679) );
  XNOR U2555 ( .A(n4771), .B(n1679), .Z(out[1249]) );
  XOR U2556 ( .A(in[595]), .B(n3695), .Z(n2600) );
  XOR U2557 ( .A(in[250]), .B(n3792), .Z(n3402) );
  XNOR U2558 ( .A(in[1470]), .B(n3553), .Z(n3399) );
  NAND U2559 ( .A(n3402), .B(n3399), .Z(n1680) );
  XNOR U2560 ( .A(n2600), .B(n1680), .Z(out[124]) );
  OR U2561 ( .A(n4776), .B(n1681), .Z(n1682) );
  XNOR U2562 ( .A(n4775), .B(n1682), .Z(out[1250]) );
  OR U2563 ( .A(n4780), .B(n1683), .Z(n1684) );
  XNOR U2564 ( .A(n4779), .B(n1684), .Z(out[1251]) );
  OR U2565 ( .A(n4784), .B(n1685), .Z(n1686) );
  XNOR U2566 ( .A(n4783), .B(n1686), .Z(out[1252]) );
  OR U2567 ( .A(n4788), .B(n1687), .Z(n1688) );
  XNOR U2568 ( .A(n4787), .B(n1688), .Z(out[1253]) );
  OR U2569 ( .A(n4792), .B(n1689), .Z(n1690) );
  XNOR U2570 ( .A(n4791), .B(n1690), .Z(out[1254]) );
  OR U2571 ( .A(n4796), .B(n1691), .Z(n1692) );
  XNOR U2572 ( .A(n4795), .B(n1692), .Z(out[1255]) );
  ANDN U2573 ( .B(n1694), .A(n1693), .Z(n1695) );
  XNOR U2574 ( .A(n1696), .B(n1695), .Z(out[1256]) );
  ANDN U2575 ( .B(n1698), .A(n1697), .Z(n1699) );
  XNOR U2576 ( .A(n1700), .B(n1699), .Z(out[1257]) );
  ANDN U2577 ( .B(n1702), .A(n1701), .Z(n1703) );
  XNOR U2578 ( .A(n1704), .B(n1703), .Z(out[1258]) );
  ANDN U2579 ( .B(n1706), .A(n1705), .Z(n1707) );
  XNOR U2580 ( .A(n1708), .B(n1707), .Z(out[1259]) );
  XOR U2581 ( .A(in[596]), .B(n3699), .Z(n2602) );
  XNOR U2582 ( .A(in[251]), .B(n3802), .Z(n3446) );
  XNOR U2583 ( .A(in[1471]), .B(n3557), .Z(n3443) );
  NAND U2584 ( .A(n3446), .B(n3443), .Z(n1709) );
  XNOR U2585 ( .A(n2602), .B(n1709), .Z(out[125]) );
  ANDN U2586 ( .B(n1711), .A(n1710), .Z(n1712) );
  XNOR U2587 ( .A(n1713), .B(n1712), .Z(out[1260]) );
  ANDN U2588 ( .B(n1715), .A(n1714), .Z(n1716) );
  XNOR U2589 ( .A(n1717), .B(n1716), .Z(out[1261]) );
  ANDN U2590 ( .B(n1719), .A(n1718), .Z(n1720) );
  XNOR U2591 ( .A(n1721), .B(n1720), .Z(out[1262]) );
  ANDN U2592 ( .B(n1723), .A(n1722), .Z(n1724) );
  XNOR U2593 ( .A(n1725), .B(n1724), .Z(out[1263]) );
  ANDN U2594 ( .B(n1727), .A(n1726), .Z(n1728) );
  XNOR U2595 ( .A(n1729), .B(n1728), .Z(out[1264]) );
  ANDN U2596 ( .B(n1731), .A(n1730), .Z(n1732) );
  XNOR U2597 ( .A(n1733), .B(n1732), .Z(out[1265]) );
  ANDN U2598 ( .B(n1735), .A(n1734), .Z(n1736) );
  XNOR U2599 ( .A(n1737), .B(n1736), .Z(out[1266]) );
  ANDN U2600 ( .B(n1739), .A(n1738), .Z(n1740) );
  XNOR U2601 ( .A(n1741), .B(n1740), .Z(out[1267]) );
  ANDN U2602 ( .B(n1743), .A(n1742), .Z(n1744) );
  XNOR U2603 ( .A(n1745), .B(n1744), .Z(out[1268]) );
  ANDN U2604 ( .B(n1747), .A(n1746), .Z(n1748) );
  XNOR U2605 ( .A(n1749), .B(n1748), .Z(out[1269]) );
  XOR U2606 ( .A(in[597]), .B(n3703), .Z(n2604) );
  XNOR U2607 ( .A(in[252]), .B(n3806), .Z(n3490) );
  XNOR U2608 ( .A(in[1408]), .B(n3561), .Z(n3487) );
  NAND U2609 ( .A(n3490), .B(n3487), .Z(n1750) );
  XNOR U2610 ( .A(n2604), .B(n1750), .Z(out[126]) );
  ANDN U2611 ( .B(n1752), .A(n1751), .Z(n1753) );
  XNOR U2612 ( .A(n1754), .B(n1753), .Z(out[1270]) );
  ANDN U2613 ( .B(n1756), .A(n1755), .Z(n1757) );
  XNOR U2614 ( .A(n1758), .B(n1757), .Z(out[1271]) );
  ANDN U2615 ( .B(n1760), .A(n1759), .Z(n1761) );
  XNOR U2616 ( .A(n1762), .B(n1761), .Z(out[1272]) );
  ANDN U2617 ( .B(n1764), .A(n1763), .Z(n1765) );
  XNOR U2618 ( .A(n1766), .B(n1765), .Z(out[1273]) );
  ANDN U2619 ( .B(n1768), .A(n1767), .Z(n1769) );
  XNOR U2620 ( .A(n1770), .B(n1769), .Z(out[1274]) );
  ANDN U2621 ( .B(n1772), .A(n1771), .Z(n1773) );
  XNOR U2622 ( .A(n1774), .B(n1773), .Z(out[1275]) );
  ANDN U2623 ( .B(n1776), .A(n1775), .Z(n1777) );
  XNOR U2624 ( .A(n1778), .B(n1777), .Z(out[1276]) );
  ANDN U2625 ( .B(n1780), .A(n1779), .Z(n1781) );
  XNOR U2626 ( .A(n1782), .B(n1781), .Z(out[1277]) );
  ANDN U2627 ( .B(n1784), .A(n1783), .Z(n1785) );
  XNOR U2628 ( .A(n1786), .B(n1785), .Z(out[1278]) );
  ANDN U2629 ( .B(n1788), .A(n1787), .Z(n1789) );
  XNOR U2630 ( .A(n1790), .B(n1789), .Z(out[1279]) );
  XOR U2631 ( .A(in[598]), .B(n3711), .Z(n2606) );
  XNOR U2632 ( .A(in[253]), .B(n3810), .Z(n3534) );
  XNOR U2633 ( .A(in[1409]), .B(n3565), .Z(n3531) );
  NAND U2634 ( .A(n3534), .B(n3531), .Z(n1791) );
  XNOR U2635 ( .A(n2606), .B(n1791), .Z(out[127]) );
  XNOR U2636 ( .A(in[50]), .B(n3951), .Z(n1934) );
  XOR U2637 ( .A(in[1536]), .B(n3611), .Z(n2206) );
  XNOR U2638 ( .A(in[1172]), .B(n3628), .Z(n2204) );
  NAND U2639 ( .A(n2206), .B(n2204), .Z(n1792) );
  XNOR U2640 ( .A(n1934), .B(n1792), .Z(out[1280]) );
  XNOR U2641 ( .A(in[51]), .B(n3953), .Z(n1936) );
  XOR U2642 ( .A(in[1537]), .B(n3615), .Z(n2211) );
  XNOR U2643 ( .A(in[1173]), .B(n3632), .Z(n2209) );
  NAND U2644 ( .A(n2211), .B(n2209), .Z(n1793) );
  XNOR U2645 ( .A(n1936), .B(n1793), .Z(out[1281]) );
  XNOR U2646 ( .A(in[52]), .B(n3955), .Z(n1939) );
  XOR U2647 ( .A(in[1538]), .B(n3623), .Z(n2217) );
  XNOR U2648 ( .A(in[1174]), .B(n3636), .Z(n2214) );
  NAND U2649 ( .A(n2217), .B(n2214), .Z(n1794) );
  XNOR U2650 ( .A(n1939), .B(n1794), .Z(out[1282]) );
  XNOR U2651 ( .A(in[53]), .B(n3957), .Z(n1941) );
  XOR U2652 ( .A(in[1539]), .B(n3627), .Z(n2220) );
  XNOR U2653 ( .A(in[1175]), .B(n3640), .Z(n2218) );
  NAND U2654 ( .A(n2220), .B(n2218), .Z(n1795) );
  XNOR U2655 ( .A(n1941), .B(n1795), .Z(out[1283]) );
  XNOR U2656 ( .A(in[54]), .B(n3959), .Z(n1943) );
  XNOR U2657 ( .A(in[1540]), .B(n3631), .Z(n2227) );
  XNOR U2658 ( .A(in[1176]), .B(n3644), .Z(n2224) );
  NAND U2659 ( .A(n2227), .B(n2224), .Z(n1796) );
  XNOR U2660 ( .A(n1943), .B(n1796), .Z(out[1284]) );
  XNOR U2661 ( .A(in[55]), .B(n3961), .Z(n1945) );
  XNOR U2662 ( .A(in[1541]), .B(n3635), .Z(n2231) );
  XNOR U2663 ( .A(in[1177]), .B(n3648), .Z(n2228) );
  NAND U2664 ( .A(n2231), .B(n2228), .Z(n1797) );
  XNOR U2665 ( .A(n1945), .B(n1797), .Z(out[1285]) );
  XNOR U2666 ( .A(in[56]), .B(n3817), .Z(n1947) );
  XNOR U2667 ( .A(in[1542]), .B(n3639), .Z(n2235) );
  XNOR U2668 ( .A(in[1178]), .B(n3652), .Z(n2232) );
  NAND U2669 ( .A(n2235), .B(n2232), .Z(n1798) );
  XNOR U2670 ( .A(n1947), .B(n1798), .Z(out[1286]) );
  XNOR U2671 ( .A(in[57]), .B(n3819), .Z(n1949) );
  XNOR U2672 ( .A(in[1543]), .B(n3643), .Z(n2239) );
  XNOR U2673 ( .A(in[1179]), .B(n3656), .Z(n2236) );
  NAND U2674 ( .A(n2239), .B(n2236), .Z(n1799) );
  XNOR U2675 ( .A(n1949), .B(n1799), .Z(out[1287]) );
  XNOR U2676 ( .A(in[58]), .B(n3821), .Z(n1951) );
  XNOR U2677 ( .A(in[1544]), .B(n3647), .Z(n2243) );
  XNOR U2678 ( .A(in[1180]), .B(n3660), .Z(n2240) );
  NAND U2679 ( .A(n2243), .B(n2240), .Z(n1800) );
  XNOR U2680 ( .A(n1951), .B(n1800), .Z(out[1288]) );
  XNOR U2681 ( .A(in[59]), .B(n3823), .Z(n1953) );
  XNOR U2682 ( .A(in[1545]), .B(n3651), .Z(n2247) );
  XNOR U2683 ( .A(in[1181]), .B(n3668), .Z(n2244) );
  NAND U2684 ( .A(n2247), .B(n2244), .Z(n1801) );
  XNOR U2685 ( .A(n1953), .B(n1801), .Z(out[1289]) );
  XNOR U2686 ( .A(in[665]), .B(n3891), .Z(n2609) );
  XNOR U2687 ( .A(in[599]), .B(n3715), .Z(n3578) );
  NAND U2688 ( .A(n3578), .B(n3576), .Z(n1802) );
  XNOR U2689 ( .A(n2609), .B(n1802), .Z(out[128]) );
  XNOR U2690 ( .A(in[60]), .B(n3825), .Z(n1955) );
  XNOR U2691 ( .A(in[1546]), .B(n3655), .Z(n2251) );
  XNOR U2692 ( .A(in[1182]), .B(n3672), .Z(n2248) );
  NAND U2693 ( .A(n2251), .B(n2248), .Z(n1803) );
  XNOR U2694 ( .A(n1955), .B(n1803), .Z(out[1290]) );
  XNOR U2695 ( .A(in[61]), .B(n3827), .Z(n1957) );
  XNOR U2696 ( .A(in[1547]), .B(n3659), .Z(n2255) );
  XNOR U2697 ( .A(in[1183]), .B(n3676), .Z(n2252) );
  NAND U2698 ( .A(n2255), .B(n2252), .Z(n1804) );
  XNOR U2699 ( .A(n1957), .B(n1804), .Z(out[1291]) );
  XNOR U2700 ( .A(in[62]), .B(n3833), .Z(n1960) );
  XNOR U2701 ( .A(in[1548]), .B(n3667), .Z(n2259) );
  XNOR U2702 ( .A(in[1184]), .B(n3680), .Z(n2256) );
  NAND U2703 ( .A(n2259), .B(n2256), .Z(n1805) );
  XNOR U2704 ( .A(n1960), .B(n1805), .Z(out[1292]) );
  XNOR U2705 ( .A(in[63]), .B(n3835), .Z(n1962) );
  XNOR U2706 ( .A(in[1549]), .B(n3671), .Z(n2263) );
  XNOR U2707 ( .A(in[1185]), .B(n3684), .Z(n2260) );
  NAND U2708 ( .A(n2263), .B(n2260), .Z(n1806) );
  XNOR U2709 ( .A(n1962), .B(n1806), .Z(out[1293]) );
  XNOR U2710 ( .A(in[0]), .B(n3837), .Z(n1964) );
  XNOR U2711 ( .A(in[1550]), .B(n3675), .Z(n2268) );
  XOR U2712 ( .A(n3688), .B(in[1186]), .Z(n2265) );
  NAND U2713 ( .A(n2268), .B(n2265), .Z(n1807) );
  XNOR U2714 ( .A(n1964), .B(n1807), .Z(out[1294]) );
  XNOR U2715 ( .A(in[1]), .B(n3839), .Z(n1966) );
  XNOR U2716 ( .A(in[1551]), .B(n3679), .Z(n2271) );
  XOR U2717 ( .A(n3692), .B(in[1187]), .Z(n2269) );
  NAND U2718 ( .A(n2271), .B(n2269), .Z(n1808) );
  XNOR U2719 ( .A(n1966), .B(n1808), .Z(out[1295]) );
  XNOR U2720 ( .A(in[2]), .B(n3841), .Z(n1968) );
  XNOR U2721 ( .A(in[1552]), .B(n3683), .Z(n2277) );
  XOR U2722 ( .A(n3696), .B(in[1188]), .Z(n2274) );
  NAND U2723 ( .A(n2277), .B(n2274), .Z(n1809) );
  XNOR U2724 ( .A(n1968), .B(n1809), .Z(out[1296]) );
  XNOR U2725 ( .A(in[3]), .B(n3843), .Z(n1970) );
  XNOR U2726 ( .A(in[1553]), .B(n3687), .Z(n2281) );
  XOR U2727 ( .A(n3700), .B(in[1189]), .Z(n2278) );
  NAND U2728 ( .A(n2281), .B(n2278), .Z(n1810) );
  XNOR U2729 ( .A(n1970), .B(n1810), .Z(out[1297]) );
  XNOR U2730 ( .A(in[4]), .B(n3845), .Z(n1972) );
  XNOR U2731 ( .A(in[1554]), .B(n3691), .Z(n2285) );
  XNOR U2732 ( .A(in[1190]), .B(n3704), .Z(n2282) );
  NAND U2733 ( .A(n2285), .B(n2282), .Z(n1811) );
  XNOR U2734 ( .A(n1972), .B(n1811), .Z(out[1298]) );
  XNOR U2735 ( .A(in[5]), .B(n3847), .Z(n1974) );
  XNOR U2736 ( .A(in[1555]), .B(n3695), .Z(n2289) );
  XNOR U2737 ( .A(in[1191]), .B(n3712), .Z(n2286) );
  NAND U2738 ( .A(n2289), .B(n2286), .Z(n1812) );
  XNOR U2739 ( .A(n1974), .B(n1812), .Z(out[1299]) );
  XNOR U2740 ( .A(in[666]), .B(n3893), .Z(n2611) );
  XNOR U2741 ( .A(in[600]), .B(n3719), .Z(n3622) );
  XOR U2742 ( .A(in[255]), .B(n3536), .Z(n3620) );
  NAND U2743 ( .A(n3622), .B(n3620), .Z(n1813) );
  XNOR U2744 ( .A(n2611), .B(n1813), .Z(out[129]) );
  XOR U2745 ( .A(in[202]), .B(n3584), .Z(n3970) );
  XNOR U2746 ( .A(in[1422]), .B(n3625), .Z(n3969) );
  XOR U2747 ( .A(in[1045]), .B(n4125), .Z(n2637) );
  NAND U2748 ( .A(n3969), .B(n2637), .Z(n1814) );
  XNOR U2749 ( .A(n3970), .B(n1814), .Z(out[12]) );
  XNOR U2750 ( .A(in[6]), .B(n3849), .Z(n1976) );
  XNOR U2751 ( .A(in[1556]), .B(n3699), .Z(n2293) );
  XNOR U2752 ( .A(in[1192]), .B(n3716), .Z(n2290) );
  NAND U2753 ( .A(n2293), .B(n2290), .Z(n1815) );
  XNOR U2754 ( .A(n1976), .B(n1815), .Z(out[1300]) );
  XNOR U2755 ( .A(in[7]), .B(n3851), .Z(n1978) );
  XNOR U2756 ( .A(in[1557]), .B(n3703), .Z(n2297) );
  XNOR U2757 ( .A(in[1193]), .B(n3720), .Z(n2294) );
  NAND U2758 ( .A(n2297), .B(n2294), .Z(n1816) );
  XNOR U2759 ( .A(n1978), .B(n1816), .Z(out[1301]) );
  XNOR U2760 ( .A(in[8]), .B(n3855), .Z(n1981) );
  XNOR U2761 ( .A(in[1558]), .B(n3711), .Z(n2301) );
  XNOR U2762 ( .A(in[1194]), .B(n3724), .Z(n2298) );
  NAND U2763 ( .A(n2301), .B(n2298), .Z(n1817) );
  XNOR U2764 ( .A(n1981), .B(n1817), .Z(out[1302]) );
  XNOR U2765 ( .A(in[9]), .B(n3857), .Z(n1983) );
  XNOR U2766 ( .A(in[1559]), .B(n3715), .Z(n2305) );
  XNOR U2767 ( .A(in[1195]), .B(n3728), .Z(n2302) );
  NAND U2768 ( .A(n2305), .B(n2302), .Z(n1818) );
  XNOR U2769 ( .A(n1983), .B(n1818), .Z(out[1303]) );
  XNOR U2770 ( .A(in[10]), .B(n3859), .Z(n1985) );
  XNOR U2771 ( .A(in[1560]), .B(n3719), .Z(n2310) );
  XNOR U2772 ( .A(in[1196]), .B(n3732), .Z(n2307) );
  NAND U2773 ( .A(n2310), .B(n2307), .Z(n1819) );
  XNOR U2774 ( .A(n1985), .B(n1819), .Z(out[1304]) );
  XNOR U2775 ( .A(in[11]), .B(n3861), .Z(n1987) );
  XNOR U2776 ( .A(in[1561]), .B(n3723), .Z(n2314) );
  XNOR U2777 ( .A(in[1197]), .B(n3736), .Z(n2311) );
  NAND U2778 ( .A(n2314), .B(n2311), .Z(n1820) );
  XNOR U2779 ( .A(n1987), .B(n1820), .Z(out[1305]) );
  XNOR U2780 ( .A(in[12]), .B(n3863), .Z(n1989) );
  XNOR U2781 ( .A(in[1562]), .B(n3727), .Z(n2318) );
  XNOR U2782 ( .A(in[1198]), .B(n3740), .Z(n2315) );
  NAND U2783 ( .A(n2318), .B(n2315), .Z(n1821) );
  XNOR U2784 ( .A(n1989), .B(n1821), .Z(out[1306]) );
  XNOR U2785 ( .A(in[13]), .B(n3865), .Z(n1991) );
  XNOR U2786 ( .A(in[1563]), .B(n3731), .Z(n2322) );
  XNOR U2787 ( .A(in[1199]), .B(n3744), .Z(n2319) );
  NAND U2788 ( .A(n2322), .B(n2319), .Z(n1822) );
  XNOR U2789 ( .A(n1991), .B(n1822), .Z(out[1307]) );
  XNOR U2790 ( .A(in[14]), .B(n3867), .Z(n1993) );
  XNOR U2791 ( .A(in[1564]), .B(n3735), .Z(n2326) );
  XNOR U2792 ( .A(in[1200]), .B(n3748), .Z(n2323) );
  NAND U2793 ( .A(n2326), .B(n2323), .Z(n1823) );
  XNOR U2794 ( .A(n1993), .B(n1823), .Z(out[1308]) );
  XNOR U2795 ( .A(in[15]), .B(n3869), .Z(n1995) );
  XNOR U2796 ( .A(in[1565]), .B(n3739), .Z(n2330) );
  XNOR U2797 ( .A(in[1201]), .B(n3756), .Z(n2327) );
  NAND U2798 ( .A(n2330), .B(n2327), .Z(n1824) );
  XNOR U2799 ( .A(n1995), .B(n1824), .Z(out[1309]) );
  XNOR U2800 ( .A(in[667]), .B(n3895), .Z(n2614) );
  XNOR U2801 ( .A(in[601]), .B(n3723), .Z(n3666) );
  XOR U2802 ( .A(in[192]), .B(n3540), .Z(n3663) );
  NAND U2803 ( .A(n3666), .B(n3663), .Z(n1825) );
  XNOR U2804 ( .A(n2614), .B(n1825), .Z(out[130]) );
  XNOR U2805 ( .A(in[16]), .B(n3871), .Z(n1997) );
  XNOR U2806 ( .A(in[1566]), .B(n3743), .Z(n2334) );
  XNOR U2807 ( .A(in[1202]), .B(n3760), .Z(n2331) );
  NAND U2808 ( .A(n2334), .B(n2331), .Z(n1826) );
  XNOR U2809 ( .A(n1997), .B(n1826), .Z(out[1310]) );
  XNOR U2810 ( .A(in[17]), .B(n3873), .Z(n1999) );
  XNOR U2811 ( .A(in[1567]), .B(n3747), .Z(n2337) );
  XNOR U2812 ( .A(in[1203]), .B(n3764), .Z(n2335) );
  NAND U2813 ( .A(n2337), .B(n2335), .Z(n1827) );
  XNOR U2814 ( .A(n1999), .B(n1827), .Z(out[1311]) );
  XNOR U2815 ( .A(in[18]), .B(n3877), .Z(n2002) );
  XNOR U2816 ( .A(in[1568]), .B(n3755), .Z(n2343) );
  XNOR U2817 ( .A(in[1204]), .B(n3768), .Z(n2340) );
  NAND U2818 ( .A(n2343), .B(n2340), .Z(n1828) );
  XNOR U2819 ( .A(n2002), .B(n1828), .Z(out[1312]) );
  XNOR U2820 ( .A(in[19]), .B(n3879), .Z(n2004) );
  XNOR U2821 ( .A(in[1569]), .B(n3759), .Z(n2347) );
  XNOR U2822 ( .A(in[1205]), .B(n3772), .Z(n2344) );
  NAND U2823 ( .A(n2347), .B(n2344), .Z(n1829) );
  XNOR U2824 ( .A(n2004), .B(n1829), .Z(out[1313]) );
  XNOR U2825 ( .A(in[20]), .B(n3881), .Z(n2006) );
  XNOR U2826 ( .A(in[1570]), .B(n3763), .Z(n2352) );
  XNOR U2827 ( .A(in[1206]), .B(n3776), .Z(n2349) );
  NAND U2828 ( .A(n2352), .B(n2349), .Z(n1830) );
  XNOR U2829 ( .A(n2006), .B(n1830), .Z(out[1314]) );
  XNOR U2830 ( .A(in[21]), .B(n3883), .Z(n2008) );
  XNOR U2831 ( .A(in[1571]), .B(n3767), .Z(n2356) );
  XNOR U2832 ( .A(in[1207]), .B(n3780), .Z(n2353) );
  NAND U2833 ( .A(n2356), .B(n2353), .Z(n1831) );
  XNOR U2834 ( .A(n2008), .B(n1831), .Z(out[1315]) );
  XNOR U2835 ( .A(in[22]), .B(n3885), .Z(n2010) );
  XNOR U2836 ( .A(in[1572]), .B(n3771), .Z(n2360) );
  XNOR U2837 ( .A(in[1208]), .B(n3784), .Z(n2357) );
  NAND U2838 ( .A(n2360), .B(n2357), .Z(n1832) );
  XNOR U2839 ( .A(n2010), .B(n1832), .Z(out[1316]) );
  XNOR U2840 ( .A(in[23]), .B(n3887), .Z(n2012) );
  XOR U2841 ( .A(in[1573]), .B(n3775), .Z(n2364) );
  XNOR U2842 ( .A(in[1209]), .B(n3788), .Z(n2361) );
  NAND U2843 ( .A(n2364), .B(n2361), .Z(n1833) );
  XNOR U2844 ( .A(n2012), .B(n1833), .Z(out[1317]) );
  XNOR U2845 ( .A(in[24]), .B(n3889), .Z(n2014) );
  XOR U2846 ( .A(in[1574]), .B(n3779), .Z(n2368) );
  XNOR U2847 ( .A(in[1210]), .B(n3792), .Z(n2365) );
  NAND U2848 ( .A(n2368), .B(n2365), .Z(n1834) );
  XNOR U2849 ( .A(n2014), .B(n1834), .Z(out[1318]) );
  XNOR U2850 ( .A(in[25]), .B(n3891), .Z(n2016) );
  XOR U2851 ( .A(in[1575]), .B(n3783), .Z(n2372) );
  XOR U2852 ( .A(in[1211]), .B(n3802), .Z(n2369) );
  NAND U2853 ( .A(n2372), .B(n2369), .Z(n1835) );
  XNOR U2854 ( .A(n2016), .B(n1835), .Z(out[1319]) );
  XNOR U2855 ( .A(in[668]), .B(n3899), .Z(n2616) );
  XNOR U2856 ( .A(in[602]), .B(n3727), .Z(n3710) );
  XOR U2857 ( .A(in[193]), .B(n3544), .Z(n3707) );
  NAND U2858 ( .A(n3710), .B(n3707), .Z(n1836) );
  XNOR U2859 ( .A(n2616), .B(n1836), .Z(out[131]) );
  XNOR U2860 ( .A(in[26]), .B(n3893), .Z(n2018) );
  XOR U2861 ( .A(in[1576]), .B(n3787), .Z(n2376) );
  XOR U2862 ( .A(in[1212]), .B(n3806), .Z(n2373) );
  NAND U2863 ( .A(n2376), .B(n2373), .Z(n1837) );
  XNOR U2864 ( .A(n2018), .B(n1837), .Z(out[1320]) );
  XNOR U2865 ( .A(in[27]), .B(n3895), .Z(n2020) );
  XOR U2866 ( .A(in[1577]), .B(n3791), .Z(n2380) );
  XOR U2867 ( .A(in[1213]), .B(n3810), .Z(n2377) );
  NAND U2868 ( .A(n2380), .B(n2377), .Z(n1838) );
  XNOR U2869 ( .A(n2020), .B(n1838), .Z(out[1321]) );
  XNOR U2870 ( .A(in[28]), .B(n3899), .Z(n2023) );
  XOR U2871 ( .A(in[1578]), .B(n3801), .Z(n2384) );
  XNOR U2872 ( .A(in[1214]), .B(n3814), .Z(n2381) );
  NAND U2873 ( .A(n2384), .B(n2381), .Z(n1839) );
  XNOR U2874 ( .A(n2023), .B(n1839), .Z(out[1322]) );
  XNOR U2875 ( .A(in[29]), .B(n3901), .Z(n2025) );
  XOR U2876 ( .A(in[1579]), .B(n3805), .Z(n2388) );
  XOR U2877 ( .A(in[1215]), .B(n3536), .Z(n2385) );
  NAND U2878 ( .A(n2388), .B(n2385), .Z(n1840) );
  XNOR U2879 ( .A(n2025), .B(n1840), .Z(out[1323]) );
  XNOR U2880 ( .A(in[30]), .B(n3903), .Z(n2027) );
  XOR U2881 ( .A(in[1580]), .B(n3809), .Z(n2393) );
  XOR U2882 ( .A(in[1152]), .B(n3540), .Z(n2390) );
  NAND U2883 ( .A(n2393), .B(n2390), .Z(n1841) );
  XNOR U2884 ( .A(n2027), .B(n1841), .Z(out[1324]) );
  XNOR U2885 ( .A(in[31]), .B(n3905), .Z(n2029) );
  XOR U2886 ( .A(in[1581]), .B(n3813), .Z(n2397) );
  XOR U2887 ( .A(in[1153]), .B(n3544), .Z(n2394) );
  NAND U2888 ( .A(n2397), .B(n2394), .Z(n1842) );
  XNOR U2889 ( .A(n2029), .B(n1842), .Z(out[1325]) );
  XNOR U2890 ( .A(in[32]), .B(n3907), .Z(n2031) );
  XOR U2891 ( .A(in[1582]), .B(n3535), .Z(n2401) );
  XOR U2892 ( .A(in[1154]), .B(n3548), .Z(n2398) );
  NAND U2893 ( .A(n2401), .B(n2398), .Z(n1843) );
  XNOR U2894 ( .A(n2031), .B(n1843), .Z(out[1326]) );
  XNOR U2895 ( .A(in[33]), .B(n3909), .Z(n2033) );
  XOR U2896 ( .A(in[1583]), .B(n3539), .Z(n2405) );
  XOR U2897 ( .A(in[1155]), .B(n3552), .Z(n2402) );
  NAND U2898 ( .A(n2405), .B(n2402), .Z(n1844) );
  XNOR U2899 ( .A(n2033), .B(n1844), .Z(out[1327]) );
  XNOR U2900 ( .A(in[34]), .B(n3911), .Z(n2035) );
  XOR U2901 ( .A(in[1584]), .B(n3543), .Z(n2409) );
  XOR U2902 ( .A(in[1156]), .B(n3556), .Z(n2406) );
  NAND U2903 ( .A(n2409), .B(n2406), .Z(n1845) );
  XNOR U2904 ( .A(n2035), .B(n1845), .Z(out[1328]) );
  XNOR U2905 ( .A(in[35]), .B(n3913), .Z(n2037) );
  XOR U2906 ( .A(in[1585]), .B(n3547), .Z(n2413) );
  XOR U2907 ( .A(in[1157]), .B(n3560), .Z(n2410) );
  NAND U2908 ( .A(n2413), .B(n2410), .Z(n1846) );
  XNOR U2909 ( .A(n2037), .B(n1846), .Z(out[1329]) );
  XNOR U2910 ( .A(in[669]), .B(n3901), .Z(n2619) );
  XNOR U2911 ( .A(in[603]), .B(n3731), .Z(n3754) );
  XOR U2912 ( .A(in[194]), .B(n3548), .Z(n3751) );
  NAND U2913 ( .A(n3754), .B(n3751), .Z(n1847) );
  XNOR U2914 ( .A(n2619), .B(n1847), .Z(out[132]) );
  XNOR U2915 ( .A(in[36]), .B(n3915), .Z(n2039) );
  XOR U2916 ( .A(in[1586]), .B(n3551), .Z(n2417) );
  XOR U2917 ( .A(in[1158]), .B(n3564), .Z(n2414) );
  NAND U2918 ( .A(n2417), .B(n2414), .Z(n1848) );
  XNOR U2919 ( .A(n2039), .B(n1848), .Z(out[1330]) );
  XNOR U2920 ( .A(in[37]), .B(n3917), .Z(n2041) );
  XOR U2921 ( .A(in[1587]), .B(n3555), .Z(n2421) );
  XOR U2922 ( .A(in[1159]), .B(n3568), .Z(n2418) );
  NAND U2923 ( .A(n2421), .B(n2418), .Z(n1849) );
  XNOR U2924 ( .A(n2041), .B(n1849), .Z(out[1331]) );
  XNOR U2925 ( .A(in[38]), .B(n3923), .Z(n2044) );
  XOR U2926 ( .A(in[1588]), .B(n3559), .Z(n2425) );
  XOR U2927 ( .A(in[1160]), .B(n3572), .Z(n2422) );
  NAND U2928 ( .A(n2425), .B(n2422), .Z(n1850) );
  XNOR U2929 ( .A(n2044), .B(n1850), .Z(out[1332]) );
  XNOR U2930 ( .A(in[39]), .B(n3925), .Z(n2046) );
  XOR U2931 ( .A(in[1589]), .B(n3563), .Z(n2429) );
  XOR U2932 ( .A(in[1161]), .B(n3580), .Z(n2426) );
  NAND U2933 ( .A(n2429), .B(n2426), .Z(n1851) );
  XNOR U2934 ( .A(n2046), .B(n1851), .Z(out[1333]) );
  XNOR U2935 ( .A(in[40]), .B(n3927), .Z(n2048) );
  XOR U2936 ( .A(in[1590]), .B(n3567), .Z(n2434) );
  XOR U2937 ( .A(in[1162]), .B(n3584), .Z(n2431) );
  NAND U2938 ( .A(n2434), .B(n2431), .Z(n1852) );
  XNOR U2939 ( .A(n2048), .B(n1852), .Z(out[1334]) );
  XNOR U2940 ( .A(in[41]), .B(n3929), .Z(n2050) );
  XOR U2941 ( .A(in[1591]), .B(n3571), .Z(n2438) );
  XOR U2942 ( .A(in[1163]), .B(n3588), .Z(n2435) );
  NAND U2943 ( .A(n2438), .B(n2435), .Z(n1853) );
  XNOR U2944 ( .A(n2050), .B(n1853), .Z(out[1335]) );
  XNOR U2945 ( .A(in[42]), .B(n3931), .Z(n2052) );
  XOR U2946 ( .A(in[1592]), .B(n3579), .Z(n2442) );
  XOR U2947 ( .A(in[1164]), .B(n3592), .Z(n2439) );
  NAND U2948 ( .A(n2442), .B(n2439), .Z(n1854) );
  XNOR U2949 ( .A(n2052), .B(n1854), .Z(out[1336]) );
  XNOR U2950 ( .A(in[43]), .B(n3933), .Z(n2054) );
  XOR U2951 ( .A(in[1593]), .B(n3583), .Z(n2446) );
  XOR U2952 ( .A(in[1165]), .B(n3596), .Z(n2443) );
  NAND U2953 ( .A(n2446), .B(n2443), .Z(n1855) );
  XNOR U2954 ( .A(n2054), .B(n1855), .Z(out[1337]) );
  XNOR U2955 ( .A(in[44]), .B(n3935), .Z(n2056) );
  XOR U2956 ( .A(in[1594]), .B(n3587), .Z(n2450) );
  XOR U2957 ( .A(in[1166]), .B(n3600), .Z(n2447) );
  NAND U2958 ( .A(n2450), .B(n2447), .Z(n1856) );
  XNOR U2959 ( .A(n2056), .B(n1856), .Z(out[1338]) );
  XNOR U2960 ( .A(in[45]), .B(n3937), .Z(n2058) );
  XOR U2961 ( .A(in[1595]), .B(n3591), .Z(n2454) );
  XOR U2962 ( .A(in[1167]), .B(n3604), .Z(n2451) );
  NAND U2963 ( .A(n2454), .B(n2451), .Z(n1857) );
  XNOR U2964 ( .A(n2058), .B(n1857), .Z(out[1339]) );
  XNOR U2965 ( .A(in[670]), .B(n3903), .Z(n2621) );
  XNOR U2966 ( .A(in[604]), .B(n3735), .Z(n3798) );
  XOR U2967 ( .A(in[195]), .B(n3552), .Z(n3795) );
  NAND U2968 ( .A(n3798), .B(n3795), .Z(n1858) );
  XNOR U2969 ( .A(n2621), .B(n1858), .Z(out[133]) );
  XNOR U2970 ( .A(in[46]), .B(n3939), .Z(n2060) );
  XOR U2971 ( .A(in[1596]), .B(n3595), .Z(n2458) );
  XOR U2972 ( .A(in[1168]), .B(n3608), .Z(n2455) );
  NAND U2973 ( .A(n2458), .B(n2455), .Z(n1859) );
  XNOR U2974 ( .A(n2060), .B(n1859), .Z(out[1340]) );
  XNOR U2975 ( .A(in[47]), .B(n3941), .Z(n2062) );
  XOR U2976 ( .A(in[1597]), .B(n3599), .Z(n2462) );
  XOR U2977 ( .A(in[1169]), .B(n3612), .Z(n2459) );
  NAND U2978 ( .A(n2462), .B(n2459), .Z(n1860) );
  XNOR U2979 ( .A(n2062), .B(n1860), .Z(out[1341]) );
  XNOR U2980 ( .A(in[48]), .B(n3947), .Z(n2065) );
  XOR U2981 ( .A(in[1598]), .B(n3603), .Z(n2466) );
  XOR U2982 ( .A(in[1170]), .B(n3616), .Z(n2463) );
  NAND U2983 ( .A(n2466), .B(n2463), .Z(n1861) );
  XNOR U2984 ( .A(n2065), .B(n1861), .Z(out[1342]) );
  XNOR U2985 ( .A(in[49]), .B(n3949), .Z(n2067) );
  XOR U2986 ( .A(in[1599]), .B(n3607), .Z(n2469) );
  XNOR U2987 ( .A(in[1171]), .B(n3624), .Z(n2467) );
  NAND U2988 ( .A(n2469), .B(n2467), .Z(n1862) );
  XNOR U2989 ( .A(n2067), .B(n1862), .Z(out[1343]) );
  XOR U2990 ( .A(in[427]), .B(n3979), .Z(n2069) );
  NOR U2991 ( .A(n1934), .B(n2206), .Z(n1863) );
  XNOR U2992 ( .A(n2069), .B(n1863), .Z(out[1344]) );
  XOR U2993 ( .A(in[428]), .B(n3982), .Z(n2071) );
  NOR U2994 ( .A(n1936), .B(n2211), .Z(n1864) );
  XNOR U2995 ( .A(n2071), .B(n1864), .Z(out[1345]) );
  XOR U2996 ( .A(in[429]), .B(n3985), .Z(n2073) );
  NOR U2997 ( .A(n1939), .B(n2217), .Z(n1865) );
  XNOR U2998 ( .A(n2073), .B(n1865), .Z(out[1346]) );
  XOR U2999 ( .A(in[430]), .B(n3988), .Z(n2075) );
  NOR U3000 ( .A(n1941), .B(n2220), .Z(n1866) );
  XNOR U3001 ( .A(n2075), .B(n1866), .Z(out[1347]) );
  XOR U3002 ( .A(in[431]), .B(n3991), .Z(n2077) );
  NOR U3003 ( .A(n1943), .B(n2227), .Z(n1867) );
  XNOR U3004 ( .A(n2077), .B(n1867), .Z(out[1348]) );
  XOR U3005 ( .A(in[432]), .B(n3994), .Z(n2079) );
  NOR U3006 ( .A(n1945), .B(n2231), .Z(n1868) );
  XNOR U3007 ( .A(n2079), .B(n1868), .Z(out[1349]) );
  XNOR U3008 ( .A(in[671]), .B(n3905), .Z(n2623) );
  XNOR U3009 ( .A(in[605]), .B(n3739), .Z(n3832) );
  XOR U3010 ( .A(in[196]), .B(n3556), .Z(n3829) );
  NAND U3011 ( .A(n3832), .B(n3829), .Z(n1869) );
  XNOR U3012 ( .A(n2623), .B(n1869), .Z(out[134]) );
  XOR U3013 ( .A(in[433]), .B(n3997), .Z(n2081) );
  NOR U3014 ( .A(n1947), .B(n2235), .Z(n1870) );
  XNOR U3015 ( .A(n2081), .B(n1870), .Z(out[1350]) );
  XOR U3016 ( .A(in[434]), .B(n4000), .Z(n2083) );
  NOR U3017 ( .A(n1949), .B(n2239), .Z(n1871) );
  XNOR U3018 ( .A(n2083), .B(n1871), .Z(out[1351]) );
  XOR U3019 ( .A(in[435]), .B(n4007), .Z(n2086) );
  NOR U3020 ( .A(n1951), .B(n2243), .Z(n1872) );
  XNOR U3021 ( .A(n2086), .B(n1872), .Z(out[1352]) );
  XOR U3022 ( .A(in[436]), .B(n4010), .Z(n2088) );
  NOR U3023 ( .A(n1953), .B(n2247), .Z(n1873) );
  XNOR U3024 ( .A(n2088), .B(n1873), .Z(out[1353]) );
  XOR U3025 ( .A(in[437]), .B(n4013), .Z(n2090) );
  NOR U3026 ( .A(n1955), .B(n2251), .Z(n1874) );
  XNOR U3027 ( .A(n2090), .B(n1874), .Z(out[1354]) );
  XOR U3028 ( .A(in[438]), .B(n4016), .Z(n2092) );
  NOR U3029 ( .A(n1957), .B(n2255), .Z(n1875) );
  XNOR U3030 ( .A(n2092), .B(n1875), .Z(out[1355]) );
  XOR U3031 ( .A(in[439]), .B(n4019), .Z(n2094) );
  NOR U3032 ( .A(n1960), .B(n2259), .Z(n1876) );
  XNOR U3033 ( .A(n2094), .B(n1876), .Z(out[1356]) );
  XOR U3034 ( .A(in[440]), .B(n4022), .Z(n2096) );
  NOR U3035 ( .A(n1962), .B(n2263), .Z(n1877) );
  XNOR U3036 ( .A(n2096), .B(n1877), .Z(out[1357]) );
  XOR U3037 ( .A(in[441]), .B(n4025), .Z(n2098) );
  NOR U3038 ( .A(n1964), .B(n2268), .Z(n1878) );
  XNOR U3039 ( .A(n2098), .B(n1878), .Z(out[1358]) );
  XOR U3040 ( .A(in[442]), .B(n4028), .Z(n2100) );
  NOR U3041 ( .A(n1966), .B(n2271), .Z(n1879) );
  XNOR U3042 ( .A(n2100), .B(n1879), .Z(out[1359]) );
  XNOR U3043 ( .A(in[672]), .B(n3907), .Z(n2625) );
  XNOR U3044 ( .A(in[606]), .B(n3743), .Z(n3854) );
  XOR U3045 ( .A(in[197]), .B(n3560), .Z(n4078) );
  NAND U3046 ( .A(n3854), .B(n4078), .Z(n1880) );
  XNOR U3047 ( .A(n2625), .B(n1880), .Z(out[135]) );
  XOR U3048 ( .A(in[443]), .B(n4031), .Z(n2102) );
  NOR U3049 ( .A(n1968), .B(n2277), .Z(n1881) );
  XNOR U3050 ( .A(n2102), .B(n1881), .Z(out[1360]) );
  XOR U3051 ( .A(in[444]), .B(n4034), .Z(n2104) );
  NOR U3052 ( .A(n1970), .B(n2281), .Z(n1882) );
  XNOR U3053 ( .A(n2104), .B(n1882), .Z(out[1361]) );
  XOR U3054 ( .A(in[445]), .B(n4041), .Z(n2107) );
  NOR U3055 ( .A(n1972), .B(n2285), .Z(n1883) );
  XNOR U3056 ( .A(n2107), .B(n1883), .Z(out[1362]) );
  XOR U3057 ( .A(in[446]), .B(n4044), .Z(n2109) );
  NOR U3058 ( .A(n1974), .B(n2289), .Z(n1884) );
  XNOR U3059 ( .A(n2109), .B(n1884), .Z(out[1363]) );
  XOR U3060 ( .A(in[447]), .B(n4047), .Z(n2111) );
  NOR U3061 ( .A(n1976), .B(n2293), .Z(n1885) );
  XNOR U3062 ( .A(n2111), .B(n1885), .Z(out[1364]) );
  XOR U3063 ( .A(in[384]), .B(n4050), .Z(n2113) );
  NOR U3064 ( .A(n1978), .B(n2297), .Z(n1886) );
  XNOR U3065 ( .A(n2113), .B(n1886), .Z(out[1365]) );
  XOR U3066 ( .A(in[385]), .B(n4053), .Z(n2115) );
  NOR U3067 ( .A(n1981), .B(n2301), .Z(n1887) );
  XNOR U3068 ( .A(n2115), .B(n1887), .Z(out[1366]) );
  XOR U3069 ( .A(in[386]), .B(n4056), .Z(n2117) );
  NOR U3070 ( .A(n1983), .B(n2305), .Z(n1888) );
  XNOR U3071 ( .A(n2117), .B(n1888), .Z(out[1367]) );
  XOR U3072 ( .A(in[387]), .B(n4059), .Z(n2119) );
  NOR U3073 ( .A(n1985), .B(n2310), .Z(n1889) );
  XNOR U3074 ( .A(n2119), .B(n1889), .Z(out[1368]) );
  XOR U3075 ( .A(in[388]), .B(n4062), .Z(n2121) );
  NOR U3076 ( .A(n1987), .B(n2314), .Z(n1890) );
  XNOR U3077 ( .A(n2121), .B(n1890), .Z(out[1369]) );
  XNOR U3078 ( .A(in[673]), .B(n3909), .Z(n2627) );
  XNOR U3079 ( .A(in[607]), .B(n3747), .Z(n3876) );
  XOR U3080 ( .A(in[198]), .B(n3564), .Z(n4362) );
  NAND U3081 ( .A(n3876), .B(n4362), .Z(n1891) );
  XNOR U3082 ( .A(n2627), .B(n1891), .Z(out[136]) );
  XOR U3083 ( .A(in[389]), .B(n4065), .Z(n2123) );
  NOR U3084 ( .A(n1989), .B(n2318), .Z(n1892) );
  XNOR U3085 ( .A(n2123), .B(n1892), .Z(out[1370]) );
  XOR U3086 ( .A(in[390]), .B(n4068), .Z(n2125) );
  NOR U3087 ( .A(n1991), .B(n2322), .Z(n1893) );
  XNOR U3088 ( .A(n2125), .B(n1893), .Z(out[1371]) );
  XOR U3089 ( .A(in[391]), .B(n4079), .Z(n2129) );
  NOR U3090 ( .A(n1993), .B(n2326), .Z(n1894) );
  XNOR U3091 ( .A(n2129), .B(n1894), .Z(out[1372]) );
  XOR U3092 ( .A(in[392]), .B(n4082), .Z(n2131) );
  NOR U3093 ( .A(n1995), .B(n2330), .Z(n1895) );
  XNOR U3094 ( .A(n2131), .B(n1895), .Z(out[1373]) );
  XOR U3095 ( .A(in[393]), .B(n4085), .Z(n2133) );
  NOR U3096 ( .A(n1997), .B(n2334), .Z(n1896) );
  XNOR U3097 ( .A(n2133), .B(n1896), .Z(out[1374]) );
  XOR U3098 ( .A(in[394]), .B(n4088), .Z(n2135) );
  NOR U3099 ( .A(n1999), .B(n2337), .Z(n1897) );
  XNOR U3100 ( .A(n2135), .B(n1897), .Z(out[1375]) );
  XOR U3101 ( .A(in[395]), .B(n4091), .Z(n2137) );
  NOR U3102 ( .A(n2002), .B(n2343), .Z(n1898) );
  XNOR U3103 ( .A(n2137), .B(n1898), .Z(out[1376]) );
  XNOR U3104 ( .A(n4094), .B(in[396]), .Z(n2139) );
  NOR U3105 ( .A(n2004), .B(n2347), .Z(n1899) );
  XNOR U3106 ( .A(n2139), .B(n1899), .Z(out[1377]) );
  XNOR U3107 ( .A(n4097), .B(in[397]), .Z(n2141) );
  NOR U3108 ( .A(n2006), .B(n2352), .Z(n1900) );
  XNOR U3109 ( .A(n2141), .B(n1900), .Z(out[1378]) );
  XNOR U3110 ( .A(n4100), .B(in[398]), .Z(n2143) );
  NOR U3111 ( .A(n2008), .B(n2356), .Z(n1901) );
  XNOR U3112 ( .A(n2143), .B(n1901), .Z(out[1379]) );
  XNOR U3113 ( .A(in[674]), .B(n3911), .Z(n2629) );
  XNOR U3114 ( .A(in[608]), .B(n3755), .Z(n3898) );
  XOR U3115 ( .A(in[199]), .B(n3568), .Z(n4806) );
  NAND U3116 ( .A(n3898), .B(n4806), .Z(n1902) );
  XNOR U3117 ( .A(n2629), .B(n1902), .Z(out[137]) );
  XNOR U3118 ( .A(n4103), .B(in[399]), .Z(n2145) );
  NOR U3119 ( .A(n2010), .B(n2360), .Z(n1903) );
  XNOR U3120 ( .A(n2145), .B(n1903), .Z(out[1380]) );
  XNOR U3121 ( .A(n4106), .B(in[400]), .Z(n2147) );
  NOR U3122 ( .A(n2012), .B(n2364), .Z(n1904) );
  XNOR U3123 ( .A(n2147), .B(n1904), .Z(out[1381]) );
  XNOR U3124 ( .A(n4113), .B(in[401]), .Z(n2150) );
  NOR U3125 ( .A(n2014), .B(n2368), .Z(n1905) );
  XNOR U3126 ( .A(n2150), .B(n1905), .Z(out[1382]) );
  XNOR U3127 ( .A(n4116), .B(in[402]), .Z(n2152) );
  NOR U3128 ( .A(n2016), .B(n2372), .Z(n1906) );
  XNOR U3129 ( .A(n2152), .B(n1906), .Z(out[1383]) );
  XNOR U3130 ( .A(n4119), .B(in[403]), .Z(n2154) );
  NOR U3131 ( .A(n2018), .B(n2376), .Z(n1907) );
  XNOR U3132 ( .A(n2154), .B(n1907), .Z(out[1384]) );
  XNOR U3133 ( .A(in[404]), .B(n4122), .Z(n2156) );
  NOR U3134 ( .A(n2020), .B(n2380), .Z(n1908) );
  XNOR U3135 ( .A(n2156), .B(n1908), .Z(out[1385]) );
  XNOR U3136 ( .A(in[405]), .B(n4125), .Z(n2158) );
  NOR U3137 ( .A(n2023), .B(n2384), .Z(n1909) );
  XNOR U3138 ( .A(n2158), .B(n1909), .Z(out[1386]) );
  XNOR U3139 ( .A(in[406]), .B(n4128), .Z(n2160) );
  NOR U3140 ( .A(n2025), .B(n2388), .Z(n1910) );
  XNOR U3141 ( .A(n2160), .B(n1910), .Z(out[1387]) );
  XNOR U3142 ( .A(in[407]), .B(n4131), .Z(n2162) );
  NOR U3143 ( .A(n2027), .B(n2393), .Z(n1911) );
  XNOR U3144 ( .A(n2162), .B(n1911), .Z(out[1388]) );
  XNOR U3145 ( .A(in[408]), .B(n4134), .Z(n2164) );
  NOR U3146 ( .A(n2029), .B(n2397), .Z(n1912) );
  XNOR U3147 ( .A(n2164), .B(n1912), .Z(out[1389]) );
  XNOR U3148 ( .A(in[675]), .B(n3913), .Z(n2632) );
  XNOR U3149 ( .A(in[609]), .B(n3759), .Z(n3922) );
  NAND U3150 ( .A(n3922), .B(n3920), .Z(n1913) );
  XNOR U3151 ( .A(n2632), .B(n1913), .Z(out[138]) );
  XNOR U3152 ( .A(in[409]), .B(n4137), .Z(n2166) );
  NOR U3153 ( .A(n2031), .B(n2401), .Z(n1914) );
  XNOR U3154 ( .A(n2166), .B(n1914), .Z(out[1390]) );
  XNOR U3155 ( .A(in[410]), .B(n4140), .Z(n2168) );
  NOR U3156 ( .A(n2033), .B(n2405), .Z(n1915) );
  XNOR U3157 ( .A(n2168), .B(n1915), .Z(out[1391]) );
  XNOR U3158 ( .A(in[411]), .B(n4147), .Z(n2171) );
  NOR U3159 ( .A(n2035), .B(n2409), .Z(n1916) );
  XNOR U3160 ( .A(n2171), .B(n1916), .Z(out[1392]) );
  XNOR U3161 ( .A(in[412]), .B(n4150), .Z(n2173) );
  NOR U3162 ( .A(n2037), .B(n2413), .Z(n1917) );
  XNOR U3163 ( .A(n2173), .B(n1917), .Z(out[1393]) );
  XNOR U3164 ( .A(in[413]), .B(n4153), .Z(n2175) );
  NOR U3165 ( .A(n2039), .B(n2417), .Z(n1918) );
  XNOR U3166 ( .A(n2175), .B(n1918), .Z(out[1394]) );
  XNOR U3167 ( .A(in[414]), .B(n4156), .Z(n2177) );
  NOR U3168 ( .A(n2041), .B(n2421), .Z(n1919) );
  XNOR U3169 ( .A(n2177), .B(n1919), .Z(out[1395]) );
  XNOR U3170 ( .A(in[415]), .B(n4159), .Z(n2179) );
  NOR U3171 ( .A(n2044), .B(n2425), .Z(n1920) );
  XNOR U3172 ( .A(n2179), .B(n1920), .Z(out[1396]) );
  XNOR U3173 ( .A(in[416]), .B(n4162), .Z(n2181) );
  NOR U3174 ( .A(n2046), .B(n2429), .Z(n1921) );
  XNOR U3175 ( .A(n2181), .B(n1921), .Z(out[1397]) );
  XNOR U3176 ( .A(in[417]), .B(n4165), .Z(n2183) );
  NOR U3177 ( .A(n2048), .B(n2434), .Z(n1922) );
  XNOR U3178 ( .A(n2183), .B(n1922), .Z(out[1398]) );
  XNOR U3179 ( .A(in[418]), .B(n4168), .Z(n2185) );
  NOR U3180 ( .A(n2050), .B(n2438), .Z(n1923) );
  XNOR U3181 ( .A(n2185), .B(n1923), .Z(out[1399]) );
  XNOR U3182 ( .A(in[676]), .B(n3915), .Z(n2635) );
  XNOR U3183 ( .A(in[610]), .B(n3763), .Z(n3946) );
  NAND U3184 ( .A(n3946), .B(n3944), .Z(n1924) );
  XNOR U3185 ( .A(n2635), .B(n1924), .Z(out[139]) );
  XOR U3186 ( .A(in[203]), .B(n3588), .Z(n4004) );
  XNOR U3187 ( .A(in[1423]), .B(n3629), .Z(n4003) );
  XOR U3188 ( .A(in[1046]), .B(n4128), .Z(n2640) );
  NAND U3189 ( .A(n4003), .B(n2640), .Z(n1925) );
  XNOR U3190 ( .A(n4004), .B(n1925), .Z(out[13]) );
  XNOR U3191 ( .A(in[419]), .B(n4171), .Z(n2187) );
  NOR U3192 ( .A(n2052), .B(n2442), .Z(n1926) );
  XNOR U3193 ( .A(n2187), .B(n1926), .Z(out[1400]) );
  XOR U3194 ( .A(in[420]), .B(n4174), .Z(n2189) );
  NOR U3195 ( .A(n2054), .B(n2446), .Z(n1927) );
  XNOR U3196 ( .A(n2189), .B(n1927), .Z(out[1401]) );
  XOR U3197 ( .A(in[421]), .B(n4181), .Z(n2192) );
  NOR U3198 ( .A(n2056), .B(n2450), .Z(n1928) );
  XNOR U3199 ( .A(n2192), .B(n1928), .Z(out[1402]) );
  XOR U3200 ( .A(in[422]), .B(n4184), .Z(n2194) );
  NOR U3201 ( .A(n2058), .B(n2454), .Z(n1929) );
  XNOR U3202 ( .A(n2194), .B(n1929), .Z(out[1403]) );
  XOR U3203 ( .A(in[423]), .B(n3963), .Z(n2196) );
  NOR U3204 ( .A(n2060), .B(n2458), .Z(n1930) );
  XNOR U3205 ( .A(n2196), .B(n1930), .Z(out[1404]) );
  XOR U3206 ( .A(in[424]), .B(n3966), .Z(n2198) );
  NOR U3207 ( .A(n2062), .B(n2462), .Z(n1931) );
  XNOR U3208 ( .A(n2198), .B(n1931), .Z(out[1405]) );
  XOR U3209 ( .A(in[425]), .B(n3973), .Z(n2200) );
  NOR U3210 ( .A(n2065), .B(n2466), .Z(n1932) );
  XNOR U3211 ( .A(n2200), .B(n1932), .Z(out[1406]) );
  XOR U3212 ( .A(in[426]), .B(n3976), .Z(n2202) );
  NOR U3213 ( .A(n2067), .B(n2469), .Z(n1933) );
  XNOR U3214 ( .A(n2202), .B(n1933), .Z(out[1407]) );
  XOR U3215 ( .A(in[789]), .B(n3653), .Z(n2205) );
  NAND U3216 ( .A(n2069), .B(n1934), .Z(n1935) );
  XNOR U3217 ( .A(n2205), .B(n1935), .Z(out[1408]) );
  XOR U3218 ( .A(in[790]), .B(n3657), .Z(n2210) );
  NAND U3219 ( .A(n2071), .B(n1936), .Z(n1937) );
  XNOR U3220 ( .A(n2210), .B(n1937), .Z(out[1409]) );
  XNOR U3221 ( .A(in[677]), .B(n3917), .Z(n2638) );
  XNOR U3222 ( .A(in[611]), .B(n3767), .Z(n3972) );
  NAND U3223 ( .A(n3972), .B(n3970), .Z(n1938) );
  XNOR U3224 ( .A(n2638), .B(n1938), .Z(out[140]) );
  XOR U3225 ( .A(in[791]), .B(n3661), .Z(n2215) );
  NAND U3226 ( .A(n2073), .B(n1939), .Z(n1940) );
  XNOR U3227 ( .A(n2215), .B(n1940), .Z(out[1410]) );
  XOR U3228 ( .A(in[792]), .B(n3669), .Z(n2219) );
  NAND U3229 ( .A(n2075), .B(n1941), .Z(n1942) );
  XNOR U3230 ( .A(n2219), .B(n1942), .Z(out[1411]) );
  XOR U3231 ( .A(in[793]), .B(n3673), .Z(n2225) );
  NAND U3232 ( .A(n2077), .B(n1943), .Z(n1944) );
  XNOR U3233 ( .A(n2225), .B(n1944), .Z(out[1412]) );
  XOR U3234 ( .A(in[794]), .B(n3677), .Z(n2229) );
  NAND U3235 ( .A(n2079), .B(n1945), .Z(n1946) );
  XNOR U3236 ( .A(n2229), .B(n1946), .Z(out[1413]) );
  XOR U3237 ( .A(in[795]), .B(n3681), .Z(n2233) );
  NAND U3238 ( .A(n2081), .B(n1947), .Z(n1948) );
  XNOR U3239 ( .A(n2233), .B(n1948), .Z(out[1414]) );
  XOR U3240 ( .A(in[796]), .B(n3685), .Z(n2237) );
  NAND U3241 ( .A(n2083), .B(n1949), .Z(n1950) );
  XNOR U3242 ( .A(n2237), .B(n1950), .Z(out[1415]) );
  XOR U3243 ( .A(in[797]), .B(n3689), .Z(n2241) );
  NAND U3244 ( .A(n2086), .B(n1951), .Z(n1952) );
  XNOR U3245 ( .A(n2241), .B(n1952), .Z(out[1416]) );
  XOR U3246 ( .A(in[798]), .B(n3693), .Z(n2245) );
  NAND U3247 ( .A(n2088), .B(n1953), .Z(n1954) );
  XNOR U3248 ( .A(n2245), .B(n1954), .Z(out[1417]) );
  XOR U3249 ( .A(in[799]), .B(n3697), .Z(n2249) );
  NAND U3250 ( .A(n2090), .B(n1955), .Z(n1956) );
  XNOR U3251 ( .A(n2249), .B(n1956), .Z(out[1418]) );
  XOR U3252 ( .A(in[800]), .B(n3701), .Z(n2253) );
  NAND U3253 ( .A(n2092), .B(n1957), .Z(n1958) );
  XNOR U3254 ( .A(n2253), .B(n1958), .Z(out[1419]) );
  XNOR U3255 ( .A(in[678]), .B(n3923), .Z(n2641) );
  XNOR U3256 ( .A(in[612]), .B(n3771), .Z(n4006) );
  NAND U3257 ( .A(n4006), .B(n4004), .Z(n1959) );
  XNOR U3258 ( .A(n2641), .B(n1959), .Z(out[141]) );
  XOR U3259 ( .A(in[801]), .B(n3705), .Z(n2257) );
  NAND U3260 ( .A(n2094), .B(n1960), .Z(n1961) );
  XNOR U3261 ( .A(n2257), .B(n1961), .Z(out[1420]) );
  XOR U3262 ( .A(in[802]), .B(n3713), .Z(n2261) );
  NAND U3263 ( .A(n2096), .B(n1962), .Z(n1963) );
  XNOR U3264 ( .A(n2261), .B(n1963), .Z(out[1421]) );
  XOR U3265 ( .A(in[803]), .B(n3717), .Z(n2266) );
  NAND U3266 ( .A(n2098), .B(n1964), .Z(n1965) );
  XNOR U3267 ( .A(n2266), .B(n1965), .Z(out[1422]) );
  XOR U3268 ( .A(in[804]), .B(n3721), .Z(n2270) );
  NAND U3269 ( .A(n2100), .B(n1966), .Z(n1967) );
  XNOR U3270 ( .A(n2270), .B(n1967), .Z(out[1423]) );
  XOR U3271 ( .A(in[805]), .B(n3725), .Z(n2275) );
  NAND U3272 ( .A(n2102), .B(n1968), .Z(n1969) );
  XNOR U3273 ( .A(n2275), .B(n1969), .Z(out[1424]) );
  XNOR U3274 ( .A(in[806]), .B(n3729), .Z(n2279) );
  NAND U3275 ( .A(n2104), .B(n1970), .Z(n1971) );
  XNOR U3276 ( .A(n2279), .B(n1971), .Z(out[1425]) );
  XNOR U3277 ( .A(in[807]), .B(n3733), .Z(n2283) );
  NAND U3278 ( .A(n2107), .B(n1972), .Z(n1973) );
  XNOR U3279 ( .A(n2283), .B(n1973), .Z(out[1426]) );
  XNOR U3280 ( .A(in[808]), .B(n3737), .Z(n2287) );
  NAND U3281 ( .A(n2109), .B(n1974), .Z(n1975) );
  XNOR U3282 ( .A(n2287), .B(n1975), .Z(out[1427]) );
  XNOR U3283 ( .A(in[809]), .B(n3741), .Z(n2291) );
  NAND U3284 ( .A(n2111), .B(n1976), .Z(n1977) );
  XNOR U3285 ( .A(n2291), .B(n1977), .Z(out[1428]) );
  XNOR U3286 ( .A(in[810]), .B(n3745), .Z(n2295) );
  NAND U3287 ( .A(n2113), .B(n1978), .Z(n1979) );
  XNOR U3288 ( .A(n2295), .B(n1979), .Z(out[1429]) );
  XNOR U3289 ( .A(in[679]), .B(n3925), .Z(n2645) );
  XOR U3290 ( .A(in[613]), .B(n3775), .Z(n4040) );
  XOR U3291 ( .A(in[204]), .B(n3592), .Z(n4038) );
  NAND U3292 ( .A(n4040), .B(n4038), .Z(n1980) );
  XNOR U3293 ( .A(n2645), .B(n1980), .Z(out[142]) );
  XNOR U3294 ( .A(in[811]), .B(n3749), .Z(n2299) );
  NAND U3295 ( .A(n2115), .B(n1981), .Z(n1982) );
  XNOR U3296 ( .A(n2299), .B(n1982), .Z(out[1430]) );
  XNOR U3297 ( .A(in[812]), .B(n3757), .Z(n2303) );
  NAND U3298 ( .A(n2117), .B(n1983), .Z(n1984) );
  XNOR U3299 ( .A(n2303), .B(n1984), .Z(out[1431]) );
  XNOR U3300 ( .A(in[813]), .B(n3761), .Z(n2308) );
  NAND U3301 ( .A(n2119), .B(n1985), .Z(n1986) );
  XNOR U3302 ( .A(n2308), .B(n1986), .Z(out[1432]) );
  XNOR U3303 ( .A(in[814]), .B(n3765), .Z(n2312) );
  NAND U3304 ( .A(n2121), .B(n1987), .Z(n1988) );
  XNOR U3305 ( .A(n2312), .B(n1988), .Z(out[1433]) );
  XNOR U3306 ( .A(in[815]), .B(n3769), .Z(n2316) );
  NAND U3307 ( .A(n2123), .B(n1989), .Z(n1990) );
  XNOR U3308 ( .A(n2316), .B(n1990), .Z(out[1434]) );
  XNOR U3309 ( .A(in[816]), .B(n3773), .Z(n2320) );
  NAND U3310 ( .A(n2125), .B(n1991), .Z(n1992) );
  XNOR U3311 ( .A(n2320), .B(n1992), .Z(out[1435]) );
  XNOR U3312 ( .A(in[817]), .B(n3777), .Z(n2324) );
  NAND U3313 ( .A(n2129), .B(n1993), .Z(n1994) );
  XNOR U3314 ( .A(n2324), .B(n1994), .Z(out[1436]) );
  XNOR U3315 ( .A(in[818]), .B(n3781), .Z(n2328) );
  NAND U3316 ( .A(n2131), .B(n1995), .Z(n1996) );
  XNOR U3317 ( .A(n2328), .B(n1996), .Z(out[1437]) );
  XNOR U3318 ( .A(in[819]), .B(n3785), .Z(n2332) );
  NAND U3319 ( .A(n2133), .B(n1997), .Z(n1998) );
  XNOR U3320 ( .A(n2332), .B(n1998), .Z(out[1438]) );
  XNOR U3321 ( .A(in[820]), .B(n3789), .Z(n2336) );
  NAND U3322 ( .A(n2135), .B(n1999), .Z(n2000) );
  XNOR U3323 ( .A(n2336), .B(n2000), .Z(out[1439]) );
  XNOR U3324 ( .A(in[680]), .B(n3927), .Z(n2648) );
  XOR U3325 ( .A(in[614]), .B(n3779), .Z(n4074) );
  XOR U3326 ( .A(in[205]), .B(n3596), .Z(n4072) );
  NAND U3327 ( .A(n4074), .B(n4072), .Z(n2001) );
  XNOR U3328 ( .A(n2648), .B(n2001), .Z(out[143]) );
  XNOR U3329 ( .A(in[821]), .B(n3793), .Z(n2341) );
  NAND U3330 ( .A(n2137), .B(n2002), .Z(n2003) );
  XNOR U3331 ( .A(n2341), .B(n2003), .Z(out[1440]) );
  XNOR U3332 ( .A(in[822]), .B(n3803), .Z(n2345) );
  NAND U3333 ( .A(n2139), .B(n2004), .Z(n2005) );
  XNOR U3334 ( .A(n2345), .B(n2005), .Z(out[1441]) );
  XNOR U3335 ( .A(in[823]), .B(n3807), .Z(n2350) );
  NAND U3336 ( .A(n2141), .B(n2006), .Z(n2007) );
  XNOR U3337 ( .A(n2350), .B(n2007), .Z(out[1442]) );
  XNOR U3338 ( .A(in[824]), .B(n3811), .Z(n2354) );
  NAND U3339 ( .A(n2143), .B(n2008), .Z(n2009) );
  XNOR U3340 ( .A(n2354), .B(n2009), .Z(out[1443]) );
  XNOR U3341 ( .A(in[825]), .B(n3815), .Z(n2358) );
  NAND U3342 ( .A(n2145), .B(n2010), .Z(n2011) );
  XNOR U3343 ( .A(n2358), .B(n2011), .Z(out[1444]) );
  XNOR U3344 ( .A(in[826]), .B(n3537), .Z(n2362) );
  NAND U3345 ( .A(n2147), .B(n2012), .Z(n2013) );
  XNOR U3346 ( .A(n2362), .B(n2013), .Z(out[1445]) );
  XNOR U3347 ( .A(in[827]), .B(n3541), .Z(n2366) );
  NAND U3348 ( .A(n2150), .B(n2014), .Z(n2015) );
  XNOR U3349 ( .A(n2366), .B(n2015), .Z(out[1446]) );
  XNOR U3350 ( .A(in[828]), .B(n3545), .Z(n2370) );
  NAND U3351 ( .A(n2152), .B(n2016), .Z(n2017) );
  XNOR U3352 ( .A(n2370), .B(n2017), .Z(out[1447]) );
  XNOR U3353 ( .A(in[829]), .B(n3549), .Z(n2374) );
  NAND U3354 ( .A(n2154), .B(n2018), .Z(n2019) );
  XNOR U3355 ( .A(n2374), .B(n2019), .Z(out[1448]) );
  XNOR U3356 ( .A(in[830]), .B(n3553), .Z(n2378) );
  NAND U3357 ( .A(n2156), .B(n2020), .Z(n2021) );
  XNOR U3358 ( .A(n2378), .B(n2021), .Z(out[1449]) );
  XNOR U3359 ( .A(in[681]), .B(n3929), .Z(n2651) );
  XOR U3360 ( .A(in[615]), .B(n3783), .Z(n4112) );
  XOR U3361 ( .A(in[206]), .B(n3600), .Z(n4110) );
  NAND U3362 ( .A(n4112), .B(n4110), .Z(n2022) );
  XNOR U3363 ( .A(n2651), .B(n2022), .Z(out[144]) );
  XNOR U3364 ( .A(in[831]), .B(n3557), .Z(n2382) );
  NAND U3365 ( .A(n2158), .B(n2023), .Z(n2024) );
  XNOR U3366 ( .A(n2382), .B(n2024), .Z(out[1450]) );
  XNOR U3367 ( .A(in[768]), .B(n3561), .Z(n2386) );
  NAND U3368 ( .A(n2160), .B(n2025), .Z(n2026) );
  XNOR U3369 ( .A(n2386), .B(n2026), .Z(out[1451]) );
  XNOR U3370 ( .A(in[769]), .B(n3565), .Z(n2391) );
  NAND U3371 ( .A(n2162), .B(n2027), .Z(n2028) );
  XNOR U3372 ( .A(n2391), .B(n2028), .Z(out[1452]) );
  XOR U3373 ( .A(n3569), .B(in[770]), .Z(n2395) );
  NAND U3374 ( .A(n2164), .B(n2029), .Z(n2030) );
  XNOR U3375 ( .A(n2395), .B(n2030), .Z(out[1453]) );
  XOR U3376 ( .A(n3573), .B(in[771]), .Z(n2399) );
  NAND U3377 ( .A(n2166), .B(n2031), .Z(n2032) );
  XNOR U3378 ( .A(n2399), .B(n2032), .Z(out[1454]) );
  XOR U3379 ( .A(n3581), .B(in[772]), .Z(n2403) );
  NAND U3380 ( .A(n2168), .B(n2033), .Z(n2034) );
  XNOR U3381 ( .A(n2403), .B(n2034), .Z(out[1455]) );
  XOR U3382 ( .A(n3585), .B(in[773]), .Z(n2407) );
  NAND U3383 ( .A(n2171), .B(n2035), .Z(n2036) );
  XNOR U3384 ( .A(n2407), .B(n2036), .Z(out[1456]) );
  XOR U3385 ( .A(n3589), .B(in[774]), .Z(n2411) );
  NAND U3386 ( .A(n2173), .B(n2037), .Z(n2038) );
  XNOR U3387 ( .A(n2411), .B(n2038), .Z(out[1457]) );
  XOR U3388 ( .A(n3593), .B(in[775]), .Z(n2415) );
  NAND U3389 ( .A(n2175), .B(n2039), .Z(n2040) );
  XNOR U3390 ( .A(n2415), .B(n2040), .Z(out[1458]) );
  XOR U3391 ( .A(n3597), .B(in[776]), .Z(n2419) );
  NAND U3392 ( .A(n2177), .B(n2041), .Z(n2042) );
  XNOR U3393 ( .A(n2419), .B(n2042), .Z(out[1459]) );
  XNOR U3394 ( .A(in[682]), .B(n3931), .Z(n2654) );
  XOR U3395 ( .A(in[616]), .B(n3787), .Z(n4146) );
  XOR U3396 ( .A(in[207]), .B(n3604), .Z(n4144) );
  NAND U3397 ( .A(n4146), .B(n4144), .Z(n2043) );
  XNOR U3398 ( .A(n2654), .B(n2043), .Z(out[145]) );
  XOR U3399 ( .A(in[777]), .B(n3601), .Z(n2423) );
  NAND U3400 ( .A(n2179), .B(n2044), .Z(n2045) );
  XNOR U3401 ( .A(n2423), .B(n2045), .Z(out[1460]) );
  XOR U3402 ( .A(n3605), .B(in[778]), .Z(n2427) );
  NAND U3403 ( .A(n2181), .B(n2046), .Z(n2047) );
  XNOR U3404 ( .A(n2427), .B(n2047), .Z(out[1461]) );
  XOR U3405 ( .A(n3609), .B(in[779]), .Z(n2432) );
  NAND U3406 ( .A(n2183), .B(n2048), .Z(n2049) );
  XNOR U3407 ( .A(n2432), .B(n2049), .Z(out[1462]) );
  XOR U3408 ( .A(in[780]), .B(n3613), .Z(n2436) );
  NAND U3409 ( .A(n2185), .B(n2050), .Z(n2051) );
  XNOR U3410 ( .A(n2436), .B(n2051), .Z(out[1463]) );
  XOR U3411 ( .A(in[781]), .B(n3617), .Z(n2440) );
  NAND U3412 ( .A(n2187), .B(n2052), .Z(n2053) );
  XNOR U3413 ( .A(n2440), .B(n2053), .Z(out[1464]) );
  XOR U3414 ( .A(in[782]), .B(n3625), .Z(n2444) );
  NAND U3415 ( .A(n2189), .B(n2054), .Z(n2055) );
  XNOR U3416 ( .A(n2444), .B(n2055), .Z(out[1465]) );
  XOR U3417 ( .A(in[783]), .B(n3629), .Z(n2448) );
  NAND U3418 ( .A(n2192), .B(n2056), .Z(n2057) );
  XNOR U3419 ( .A(n2448), .B(n2057), .Z(out[1466]) );
  XOR U3420 ( .A(in[784]), .B(n3633), .Z(n2452) );
  NAND U3421 ( .A(n2194), .B(n2058), .Z(n2059) );
  XNOR U3422 ( .A(n2452), .B(n2059), .Z(out[1467]) );
  XOR U3423 ( .A(in[785]), .B(n3637), .Z(n2456) );
  NAND U3424 ( .A(n2196), .B(n2060), .Z(n2061) );
  XNOR U3425 ( .A(n2456), .B(n2061), .Z(out[1468]) );
  XOR U3426 ( .A(in[786]), .B(n3641), .Z(n2460) );
  NAND U3427 ( .A(n2198), .B(n2062), .Z(n2063) );
  XNOR U3428 ( .A(n2460), .B(n2063), .Z(out[1469]) );
  XNOR U3429 ( .A(in[683]), .B(n3933), .Z(n2657) );
  XOR U3430 ( .A(in[617]), .B(n3791), .Z(n4180) );
  XOR U3431 ( .A(in[208]), .B(n3608), .Z(n4178) );
  NAND U3432 ( .A(n4180), .B(n4178), .Z(n2064) );
  XNOR U3433 ( .A(n2657), .B(n2064), .Z(out[146]) );
  XOR U3434 ( .A(in[787]), .B(n3645), .Z(n2464) );
  NAND U3435 ( .A(n2200), .B(n2065), .Z(n2066) );
  XNOR U3436 ( .A(n2464), .B(n2066), .Z(out[1470]) );
  XOR U3437 ( .A(in[788]), .B(n3649), .Z(n2468) );
  NAND U3438 ( .A(n2202), .B(n2067), .Z(n2068) );
  XNOR U3439 ( .A(n2468), .B(n2068), .Z(out[1471]) );
  OR U3440 ( .A(n2205), .B(n2069), .Z(n2070) );
  XNOR U3441 ( .A(n2204), .B(n2070), .Z(out[1472]) );
  OR U3442 ( .A(n2210), .B(n2071), .Z(n2072) );
  XNOR U3443 ( .A(n2209), .B(n2072), .Z(out[1473]) );
  OR U3444 ( .A(n2215), .B(n2073), .Z(n2074) );
  XNOR U3445 ( .A(n2214), .B(n2074), .Z(out[1474]) );
  OR U3446 ( .A(n2219), .B(n2075), .Z(n2076) );
  XNOR U3447 ( .A(n2218), .B(n2076), .Z(out[1475]) );
  OR U3448 ( .A(n2225), .B(n2077), .Z(n2078) );
  XNOR U3449 ( .A(n2224), .B(n2078), .Z(out[1476]) );
  OR U3450 ( .A(n2229), .B(n2079), .Z(n2080) );
  XNOR U3451 ( .A(n2228), .B(n2080), .Z(out[1477]) );
  OR U3452 ( .A(n2233), .B(n2081), .Z(n2082) );
  XNOR U3453 ( .A(n2232), .B(n2082), .Z(out[1478]) );
  OR U3454 ( .A(n2237), .B(n2083), .Z(n2084) );
  XNOR U3455 ( .A(n2236), .B(n2084), .Z(out[1479]) );
  XNOR U3456 ( .A(in[684]), .B(n3935), .Z(n2660) );
  XOR U3457 ( .A(in[618]), .B(n3801), .Z(n4206) );
  XOR U3458 ( .A(in[209]), .B(n3612), .Z(n4204) );
  NAND U3459 ( .A(n4206), .B(n4204), .Z(n2085) );
  XNOR U3460 ( .A(n2660), .B(n2085), .Z(out[147]) );
  OR U3461 ( .A(n2241), .B(n2086), .Z(n2087) );
  XNOR U3462 ( .A(n2240), .B(n2087), .Z(out[1480]) );
  OR U3463 ( .A(n2245), .B(n2088), .Z(n2089) );
  XNOR U3464 ( .A(n2244), .B(n2089), .Z(out[1481]) );
  OR U3465 ( .A(n2249), .B(n2090), .Z(n2091) );
  XNOR U3466 ( .A(n2248), .B(n2091), .Z(out[1482]) );
  OR U3467 ( .A(n2253), .B(n2092), .Z(n2093) );
  XNOR U3468 ( .A(n2252), .B(n2093), .Z(out[1483]) );
  OR U3469 ( .A(n2257), .B(n2094), .Z(n2095) );
  XNOR U3470 ( .A(n2256), .B(n2095), .Z(out[1484]) );
  OR U3471 ( .A(n2261), .B(n2096), .Z(n2097) );
  XNOR U3472 ( .A(n2260), .B(n2097), .Z(out[1485]) );
  OR U3473 ( .A(n2266), .B(n2098), .Z(n2099) );
  XNOR U3474 ( .A(n2265), .B(n2099), .Z(out[1486]) );
  OR U3475 ( .A(n2270), .B(n2100), .Z(n2101) );
  XNOR U3476 ( .A(n2269), .B(n2101), .Z(out[1487]) );
  OR U3477 ( .A(n2275), .B(n2102), .Z(n2103) );
  XNOR U3478 ( .A(n2274), .B(n2103), .Z(out[1488]) );
  OR U3479 ( .A(n2279), .B(n2104), .Z(n2105) );
  XNOR U3480 ( .A(n2278), .B(n2105), .Z(out[1489]) );
  XNOR U3481 ( .A(in[685]), .B(n3937), .Z(n2663) );
  XOR U3482 ( .A(in[619]), .B(n3805), .Z(n4230) );
  XOR U3483 ( .A(in[210]), .B(n3616), .Z(n4228) );
  NAND U3484 ( .A(n4230), .B(n4228), .Z(n2106) );
  XNOR U3485 ( .A(n2663), .B(n2106), .Z(out[148]) );
  OR U3486 ( .A(n2283), .B(n2107), .Z(n2108) );
  XNOR U3487 ( .A(n2282), .B(n2108), .Z(out[1490]) );
  OR U3488 ( .A(n2287), .B(n2109), .Z(n2110) );
  XNOR U3489 ( .A(n2286), .B(n2110), .Z(out[1491]) );
  OR U3490 ( .A(n2291), .B(n2111), .Z(n2112) );
  XNOR U3491 ( .A(n2290), .B(n2112), .Z(out[1492]) );
  OR U3492 ( .A(n2295), .B(n2113), .Z(n2114) );
  XNOR U3493 ( .A(n2294), .B(n2114), .Z(out[1493]) );
  OR U3494 ( .A(n2299), .B(n2115), .Z(n2116) );
  XNOR U3495 ( .A(n2298), .B(n2116), .Z(out[1494]) );
  OR U3496 ( .A(n2303), .B(n2117), .Z(n2118) );
  XNOR U3497 ( .A(n2302), .B(n2118), .Z(out[1495]) );
  OR U3498 ( .A(n2308), .B(n2119), .Z(n2120) );
  XNOR U3499 ( .A(n2307), .B(n2120), .Z(out[1496]) );
  OR U3500 ( .A(n2312), .B(n2121), .Z(n2122) );
  XNOR U3501 ( .A(n2311), .B(n2122), .Z(out[1497]) );
  OR U3502 ( .A(n2316), .B(n2123), .Z(n2124) );
  XNOR U3503 ( .A(n2315), .B(n2124), .Z(out[1498]) );
  OR U3504 ( .A(n2320), .B(n2125), .Z(n2126) );
  XNOR U3505 ( .A(n2319), .B(n2126), .Z(out[1499]) );
  XNOR U3506 ( .A(in[686]), .B(n3939), .Z(n2665) );
  XOR U3507 ( .A(in[620]), .B(n3809), .Z(n4254) );
  XNOR U3508 ( .A(in[211]), .B(n3624), .Z(n4252) );
  NAND U3509 ( .A(n4254), .B(n4252), .Z(n2127) );
  XNOR U3510 ( .A(n2665), .B(n2127), .Z(out[149]) );
  XNOR U3511 ( .A(in[1424]), .B(n3633), .Z(n4037) );
  XOR U3512 ( .A(in[1047]), .B(n4131), .Z(n2644) );
  NAND U3513 ( .A(n4037), .B(n2644), .Z(n2128) );
  XNOR U3514 ( .A(n4038), .B(n2128), .Z(out[14]) );
  OR U3515 ( .A(n2324), .B(n2129), .Z(n2130) );
  XNOR U3516 ( .A(n2323), .B(n2130), .Z(out[1500]) );
  OR U3517 ( .A(n2328), .B(n2131), .Z(n2132) );
  XNOR U3518 ( .A(n2327), .B(n2132), .Z(out[1501]) );
  OR U3519 ( .A(n2332), .B(n2133), .Z(n2134) );
  XNOR U3520 ( .A(n2331), .B(n2134), .Z(out[1502]) );
  OR U3521 ( .A(n2336), .B(n2135), .Z(n2136) );
  XNOR U3522 ( .A(n2335), .B(n2136), .Z(out[1503]) );
  OR U3523 ( .A(n2341), .B(n2137), .Z(n2138) );
  XNOR U3524 ( .A(n2340), .B(n2138), .Z(out[1504]) );
  OR U3525 ( .A(n2345), .B(n2139), .Z(n2140) );
  XNOR U3526 ( .A(n2344), .B(n2140), .Z(out[1505]) );
  OR U3527 ( .A(n2350), .B(n2141), .Z(n2142) );
  XNOR U3528 ( .A(n2349), .B(n2142), .Z(out[1506]) );
  OR U3529 ( .A(n2354), .B(n2143), .Z(n2144) );
  XNOR U3530 ( .A(n2353), .B(n2144), .Z(out[1507]) );
  OR U3531 ( .A(n2358), .B(n2145), .Z(n2146) );
  XNOR U3532 ( .A(n2357), .B(n2146), .Z(out[1508]) );
  OR U3533 ( .A(n2362), .B(n2147), .Z(n2148) );
  XNOR U3534 ( .A(n2361), .B(n2148), .Z(out[1509]) );
  XNOR U3535 ( .A(in[687]), .B(n3941), .Z(n2668) );
  XOR U3536 ( .A(in[621]), .B(n3813), .Z(n4278) );
  XNOR U3537 ( .A(in[212]), .B(n3628), .Z(n4276) );
  NAND U3538 ( .A(n4278), .B(n4276), .Z(n2149) );
  XNOR U3539 ( .A(n2668), .B(n2149), .Z(out[150]) );
  OR U3540 ( .A(n2366), .B(n2150), .Z(n2151) );
  XNOR U3541 ( .A(n2365), .B(n2151), .Z(out[1510]) );
  OR U3542 ( .A(n2370), .B(n2152), .Z(n2153) );
  XNOR U3543 ( .A(n2369), .B(n2153), .Z(out[1511]) );
  OR U3544 ( .A(n2374), .B(n2154), .Z(n2155) );
  XNOR U3545 ( .A(n2373), .B(n2155), .Z(out[1512]) );
  OR U3546 ( .A(n2378), .B(n2156), .Z(n2157) );
  XNOR U3547 ( .A(n2377), .B(n2157), .Z(out[1513]) );
  OR U3548 ( .A(n2382), .B(n2158), .Z(n2159) );
  XNOR U3549 ( .A(n2381), .B(n2159), .Z(out[1514]) );
  OR U3550 ( .A(n2386), .B(n2160), .Z(n2161) );
  XNOR U3551 ( .A(n2385), .B(n2161), .Z(out[1515]) );
  OR U3552 ( .A(n2391), .B(n2162), .Z(n2163) );
  XNOR U3553 ( .A(n2390), .B(n2163), .Z(out[1516]) );
  OR U3554 ( .A(n2395), .B(n2164), .Z(n2165) );
  XNOR U3555 ( .A(n2394), .B(n2165), .Z(out[1517]) );
  OR U3556 ( .A(n2399), .B(n2166), .Z(n2167) );
  XNOR U3557 ( .A(n2398), .B(n2167), .Z(out[1518]) );
  OR U3558 ( .A(n2403), .B(n2168), .Z(n2169) );
  XNOR U3559 ( .A(n2402), .B(n2169), .Z(out[1519]) );
  XNOR U3560 ( .A(in[688]), .B(n3947), .Z(n2671) );
  XOR U3561 ( .A(in[622]), .B(n3535), .Z(n4302) );
  XNOR U3562 ( .A(in[213]), .B(n3632), .Z(n4300) );
  NAND U3563 ( .A(n4302), .B(n4300), .Z(n2170) );
  XNOR U3564 ( .A(n2671), .B(n2170), .Z(out[151]) );
  OR U3565 ( .A(n2407), .B(n2171), .Z(n2172) );
  XNOR U3566 ( .A(n2406), .B(n2172), .Z(out[1520]) );
  OR U3567 ( .A(n2411), .B(n2173), .Z(n2174) );
  XNOR U3568 ( .A(n2410), .B(n2174), .Z(out[1521]) );
  OR U3569 ( .A(n2415), .B(n2175), .Z(n2176) );
  XNOR U3570 ( .A(n2414), .B(n2176), .Z(out[1522]) );
  OR U3571 ( .A(n2419), .B(n2177), .Z(n2178) );
  XNOR U3572 ( .A(n2418), .B(n2178), .Z(out[1523]) );
  OR U3573 ( .A(n2423), .B(n2179), .Z(n2180) );
  XNOR U3574 ( .A(n2422), .B(n2180), .Z(out[1524]) );
  OR U3575 ( .A(n2427), .B(n2181), .Z(n2182) );
  XNOR U3576 ( .A(n2426), .B(n2182), .Z(out[1525]) );
  OR U3577 ( .A(n2432), .B(n2183), .Z(n2184) );
  XNOR U3578 ( .A(n2431), .B(n2184), .Z(out[1526]) );
  OR U3579 ( .A(n2436), .B(n2185), .Z(n2186) );
  XNOR U3580 ( .A(n2435), .B(n2186), .Z(out[1527]) );
  OR U3581 ( .A(n2440), .B(n2187), .Z(n2188) );
  XNOR U3582 ( .A(n2439), .B(n2188), .Z(out[1528]) );
  OR U3583 ( .A(n2444), .B(n2189), .Z(n2190) );
  XNOR U3584 ( .A(n2443), .B(n2190), .Z(out[1529]) );
  XNOR U3585 ( .A(in[689]), .B(n3949), .Z(n2675) );
  XOR U3586 ( .A(in[623]), .B(n3539), .Z(n4326) );
  XNOR U3587 ( .A(in[214]), .B(n3636), .Z(n4324) );
  NAND U3588 ( .A(n4326), .B(n4324), .Z(n2191) );
  XNOR U3589 ( .A(n2675), .B(n2191), .Z(out[152]) );
  OR U3590 ( .A(n2448), .B(n2192), .Z(n2193) );
  XNOR U3591 ( .A(n2447), .B(n2193), .Z(out[1530]) );
  OR U3592 ( .A(n2452), .B(n2194), .Z(n2195) );
  XNOR U3593 ( .A(n2451), .B(n2195), .Z(out[1531]) );
  OR U3594 ( .A(n2456), .B(n2196), .Z(n2197) );
  XNOR U3595 ( .A(n2455), .B(n2197), .Z(out[1532]) );
  OR U3596 ( .A(n2460), .B(n2198), .Z(n2199) );
  XNOR U3597 ( .A(n2459), .B(n2199), .Z(out[1533]) );
  OR U3598 ( .A(n2464), .B(n2200), .Z(n2201) );
  XNOR U3599 ( .A(n2463), .B(n2201), .Z(out[1534]) );
  OR U3600 ( .A(n2468), .B(n2202), .Z(n2203) );
  XNOR U3601 ( .A(n2467), .B(n2203), .Z(out[1535]) );
  ANDN U3602 ( .B(n2205), .A(n2204), .Z(n2208) );
  XOR U3603 ( .A(n2206), .B(round_const[0]), .Z(n2207) );
  XNOR U3604 ( .A(n2208), .B(n2207), .Z(out[1536]) );
  ANDN U3605 ( .B(n2210), .A(n2209), .Z(n2213) );
  XOR U3606 ( .A(n2211), .B(round_const[1]), .Z(n2212) );
  XNOR U3607 ( .A(n2213), .B(n2212), .Z(out[1537]) );
  ANDN U3608 ( .B(n2215), .A(n2214), .Z(n2216) );
  XNOR U3609 ( .A(n2217), .B(n2216), .Z(out[1538]) );
  ANDN U3610 ( .B(n2219), .A(n2218), .Z(n2222) );
  XOR U3611 ( .A(n2220), .B(round_const_3), .Z(n2221) );
  XNOR U3612 ( .A(n2222), .B(n2221), .Z(out[1539]) );
  XNOR U3613 ( .A(in[690]), .B(n3951), .Z(n2678) );
  XOR U3614 ( .A(in[624]), .B(n3543), .Z(n4358) );
  XNOR U3615 ( .A(in[215]), .B(n3640), .Z(n4356) );
  NAND U3616 ( .A(n4358), .B(n4356), .Z(n2223) );
  XNOR U3617 ( .A(n2678), .B(n2223), .Z(out[153]) );
  ANDN U3618 ( .B(n2225), .A(n2224), .Z(n2226) );
  XNOR U3619 ( .A(n2227), .B(n2226), .Z(out[1540]) );
  ANDN U3620 ( .B(n2229), .A(n2228), .Z(n2230) );
  XNOR U3621 ( .A(n2231), .B(n2230), .Z(out[1541]) );
  ANDN U3622 ( .B(n2233), .A(n2232), .Z(n2234) );
  XNOR U3623 ( .A(n2235), .B(n2234), .Z(out[1542]) );
  ANDN U3624 ( .B(n2237), .A(n2236), .Z(n2238) );
  XNOR U3625 ( .A(n2239), .B(n2238), .Z(out[1543]) );
  ANDN U3626 ( .B(n2241), .A(n2240), .Z(n2242) );
  XNOR U3627 ( .A(n2243), .B(n2242), .Z(out[1544]) );
  ANDN U3628 ( .B(n2245), .A(n2244), .Z(n2246) );
  XNOR U3629 ( .A(n2247), .B(n2246), .Z(out[1545]) );
  ANDN U3630 ( .B(n2249), .A(n2248), .Z(n2250) );
  XNOR U3631 ( .A(n2251), .B(n2250), .Z(out[1546]) );
  ANDN U3632 ( .B(n2253), .A(n2252), .Z(n2254) );
  XNOR U3633 ( .A(n2255), .B(n2254), .Z(out[1547]) );
  ANDN U3634 ( .B(n2257), .A(n2256), .Z(n2258) );
  XNOR U3635 ( .A(n2259), .B(n2258), .Z(out[1548]) );
  ANDN U3636 ( .B(n2261), .A(n2260), .Z(n2262) );
  XNOR U3637 ( .A(n2263), .B(n2262), .Z(out[1549]) );
  XNOR U3638 ( .A(in[691]), .B(n3953), .Z(n2681) );
  XOR U3639 ( .A(in[625]), .B(n3547), .Z(n4406) );
  XNOR U3640 ( .A(in[216]), .B(n3644), .Z(n4404) );
  NAND U3641 ( .A(n4406), .B(n4404), .Z(n2264) );
  XNOR U3642 ( .A(n2681), .B(n2264), .Z(out[154]) );
  ANDN U3643 ( .B(n2266), .A(n2265), .Z(n2267) );
  XNOR U3644 ( .A(n2268), .B(n2267), .Z(out[1550]) );
  ANDN U3645 ( .B(n2270), .A(n2269), .Z(n2273) );
  XOR U3646 ( .A(n2271), .B(round_const_15), .Z(n2272) );
  XNOR U3647 ( .A(n2273), .B(n2272), .Z(out[1551]) );
  ANDN U3648 ( .B(n2275), .A(n2274), .Z(n2276) );
  XNOR U3649 ( .A(n2277), .B(n2276), .Z(out[1552]) );
  ANDN U3650 ( .B(n2279), .A(n2278), .Z(n2280) );
  XNOR U3651 ( .A(n2281), .B(n2280), .Z(out[1553]) );
  ANDN U3652 ( .B(n2283), .A(n2282), .Z(n2284) );
  XNOR U3653 ( .A(n2285), .B(n2284), .Z(out[1554]) );
  ANDN U3654 ( .B(n2287), .A(n2286), .Z(n2288) );
  XNOR U3655 ( .A(n2289), .B(n2288), .Z(out[1555]) );
  ANDN U3656 ( .B(n2291), .A(n2290), .Z(n2292) );
  XNOR U3657 ( .A(n2293), .B(n2292), .Z(out[1556]) );
  ANDN U3658 ( .B(n2295), .A(n2294), .Z(n2296) );
  XNOR U3659 ( .A(n2297), .B(n2296), .Z(out[1557]) );
  ANDN U3660 ( .B(n2299), .A(n2298), .Z(n2300) );
  XNOR U3661 ( .A(n2301), .B(n2300), .Z(out[1558]) );
  ANDN U3662 ( .B(n2303), .A(n2302), .Z(n2304) );
  XNOR U3663 ( .A(n2305), .B(n2304), .Z(out[1559]) );
  XNOR U3664 ( .A(in[692]), .B(n3955), .Z(n2684) );
  XOR U3665 ( .A(in[626]), .B(n3551), .Z(n4450) );
  XNOR U3666 ( .A(in[217]), .B(n3648), .Z(n4448) );
  NAND U3667 ( .A(n4450), .B(n4448), .Z(n2306) );
  XNOR U3668 ( .A(n2684), .B(n2306), .Z(out[155]) );
  ANDN U3669 ( .B(n2308), .A(n2307), .Z(n2309) );
  XNOR U3670 ( .A(n2310), .B(n2309), .Z(out[1560]) );
  ANDN U3671 ( .B(n2312), .A(n2311), .Z(n2313) );
  XNOR U3672 ( .A(n2314), .B(n2313), .Z(out[1561]) );
  ANDN U3673 ( .B(n2316), .A(n2315), .Z(n2317) );
  XNOR U3674 ( .A(n2318), .B(n2317), .Z(out[1562]) );
  ANDN U3675 ( .B(n2320), .A(n2319), .Z(n2321) );
  XNOR U3676 ( .A(n2322), .B(n2321), .Z(out[1563]) );
  ANDN U3677 ( .B(n2324), .A(n2323), .Z(n2325) );
  XNOR U3678 ( .A(n2326), .B(n2325), .Z(out[1564]) );
  ANDN U3679 ( .B(n2328), .A(n2327), .Z(n2329) );
  XNOR U3680 ( .A(n2330), .B(n2329), .Z(out[1565]) );
  ANDN U3681 ( .B(n2332), .A(n2331), .Z(n2333) );
  XNOR U3682 ( .A(n2334), .B(n2333), .Z(out[1566]) );
  ANDN U3683 ( .B(n2336), .A(n2335), .Z(n2339) );
  XOR U3684 ( .A(n2337), .B(round_const_31), .Z(n2338) );
  XNOR U3685 ( .A(n2339), .B(n2338), .Z(out[1567]) );
  ANDN U3686 ( .B(n2341), .A(n2340), .Z(n2342) );
  XNOR U3687 ( .A(n2343), .B(n2342), .Z(out[1568]) );
  ANDN U3688 ( .B(n2345), .A(n2344), .Z(n2346) );
  XNOR U3689 ( .A(n2347), .B(n2346), .Z(out[1569]) );
  XNOR U3690 ( .A(in[693]), .B(n3957), .Z(n2687) );
  XOR U3691 ( .A(in[627]), .B(n3555), .Z(n4494) );
  XNOR U3692 ( .A(in[218]), .B(n3652), .Z(n4491) );
  NAND U3693 ( .A(n4494), .B(n4491), .Z(n2348) );
  XNOR U3694 ( .A(n2687), .B(n2348), .Z(out[156]) );
  ANDN U3695 ( .B(n2350), .A(n2349), .Z(n2351) );
  XNOR U3696 ( .A(n2352), .B(n2351), .Z(out[1570]) );
  ANDN U3697 ( .B(n2354), .A(n2353), .Z(n2355) );
  XNOR U3698 ( .A(n2356), .B(n2355), .Z(out[1571]) );
  ANDN U3699 ( .B(n2358), .A(n2357), .Z(n2359) );
  XNOR U3700 ( .A(n2360), .B(n2359), .Z(out[1572]) );
  ANDN U3701 ( .B(n2362), .A(n2361), .Z(n2363) );
  XNOR U3702 ( .A(n2364), .B(n2363), .Z(out[1573]) );
  ANDN U3703 ( .B(n2366), .A(n2365), .Z(n2367) );
  XNOR U3704 ( .A(n2368), .B(n2367), .Z(out[1574]) );
  ANDN U3705 ( .B(n2370), .A(n2369), .Z(n2371) );
  XNOR U3706 ( .A(n2372), .B(n2371), .Z(out[1575]) );
  ANDN U3707 ( .B(n2374), .A(n2373), .Z(n2375) );
  XNOR U3708 ( .A(n2376), .B(n2375), .Z(out[1576]) );
  ANDN U3709 ( .B(n2378), .A(n2377), .Z(n2379) );
  XNOR U3710 ( .A(n2380), .B(n2379), .Z(out[1577]) );
  ANDN U3711 ( .B(n2382), .A(n2381), .Z(n2383) );
  XNOR U3712 ( .A(n2384), .B(n2383), .Z(out[1578]) );
  ANDN U3713 ( .B(n2386), .A(n2385), .Z(n2387) );
  XNOR U3714 ( .A(n2388), .B(n2387), .Z(out[1579]) );
  XNOR U3715 ( .A(in[694]), .B(n3959), .Z(n2689) );
  XOR U3716 ( .A(in[628]), .B(n3559), .Z(n4538) );
  XNOR U3717 ( .A(in[219]), .B(n3656), .Z(n4535) );
  NAND U3718 ( .A(n4538), .B(n4535), .Z(n2389) );
  XNOR U3719 ( .A(n2689), .B(n2389), .Z(out[157]) );
  ANDN U3720 ( .B(n2391), .A(n2390), .Z(n2392) );
  XNOR U3721 ( .A(n2393), .B(n2392), .Z(out[1580]) );
  ANDN U3722 ( .B(n2395), .A(n2394), .Z(n2396) );
  XNOR U3723 ( .A(n2397), .B(n2396), .Z(out[1581]) );
  ANDN U3724 ( .B(n2399), .A(n2398), .Z(n2400) );
  XNOR U3725 ( .A(n2401), .B(n2400), .Z(out[1582]) );
  ANDN U3726 ( .B(n2403), .A(n2402), .Z(n2404) );
  XNOR U3727 ( .A(n2405), .B(n2404), .Z(out[1583]) );
  ANDN U3728 ( .B(n2407), .A(n2406), .Z(n2408) );
  XNOR U3729 ( .A(n2409), .B(n2408), .Z(out[1584]) );
  ANDN U3730 ( .B(n2411), .A(n2410), .Z(n2412) );
  XNOR U3731 ( .A(n2413), .B(n2412), .Z(out[1585]) );
  ANDN U3732 ( .B(n2415), .A(n2414), .Z(n2416) );
  XNOR U3733 ( .A(n2417), .B(n2416), .Z(out[1586]) );
  ANDN U3734 ( .B(n2419), .A(n2418), .Z(n2420) );
  XNOR U3735 ( .A(n2421), .B(n2420), .Z(out[1587]) );
  ANDN U3736 ( .B(n2423), .A(n2422), .Z(n2424) );
  XNOR U3737 ( .A(n2425), .B(n2424), .Z(out[1588]) );
  ANDN U3738 ( .B(n2427), .A(n2426), .Z(n2428) );
  XNOR U3739 ( .A(n2429), .B(n2428), .Z(out[1589]) );
  XNOR U3740 ( .A(in[695]), .B(n3961), .Z(n2691) );
  XOR U3741 ( .A(in[629]), .B(n3563), .Z(n4582) );
  XNOR U3742 ( .A(in[220]), .B(n3660), .Z(n4579) );
  NAND U3743 ( .A(n4582), .B(n4579), .Z(n2430) );
  XNOR U3744 ( .A(n2691), .B(n2430), .Z(out[158]) );
  ANDN U3745 ( .B(n2432), .A(n2431), .Z(n2433) );
  XNOR U3746 ( .A(n2434), .B(n2433), .Z(out[1590]) );
  ANDN U3747 ( .B(n2436), .A(n2435), .Z(n2437) );
  XNOR U3748 ( .A(n2438), .B(n2437), .Z(out[1591]) );
  ANDN U3749 ( .B(n2440), .A(n2439), .Z(n2441) );
  XNOR U3750 ( .A(n2442), .B(n2441), .Z(out[1592]) );
  ANDN U3751 ( .B(n2444), .A(n2443), .Z(n2445) );
  XNOR U3752 ( .A(n2446), .B(n2445), .Z(out[1593]) );
  ANDN U3753 ( .B(n2448), .A(n2447), .Z(n2449) );
  XNOR U3754 ( .A(n2450), .B(n2449), .Z(out[1594]) );
  ANDN U3755 ( .B(n2452), .A(n2451), .Z(n2453) );
  XNOR U3756 ( .A(n2454), .B(n2453), .Z(out[1595]) );
  ANDN U3757 ( .B(n2456), .A(n2455), .Z(n2457) );
  XNOR U3758 ( .A(n2458), .B(n2457), .Z(out[1596]) );
  ANDN U3759 ( .B(n2460), .A(n2459), .Z(n2461) );
  XNOR U3760 ( .A(n2462), .B(n2461), .Z(out[1597]) );
  ANDN U3761 ( .B(n2464), .A(n2463), .Z(n2465) );
  XNOR U3762 ( .A(n2466), .B(n2465), .Z(out[1598]) );
  ANDN U3763 ( .B(n2468), .A(n2467), .Z(n2471) );
  XOR U3764 ( .A(n2469), .B(round_const_63), .Z(n2470) );
  XNOR U3765 ( .A(n2471), .B(n2470), .Z(out[1599]) );
  XNOR U3766 ( .A(in[696]), .B(n3817), .Z(n2693) );
  XOR U3767 ( .A(in[630]), .B(n3567), .Z(n4626) );
  XNOR U3768 ( .A(in[221]), .B(n3668), .Z(n4623) );
  NAND U3769 ( .A(n4626), .B(n4623), .Z(n2472) );
  XNOR U3770 ( .A(n2693), .B(n2472), .Z(out[159]) );
  XNOR U3771 ( .A(in[1425]), .B(n3637), .Z(n4071) );
  XOR U3772 ( .A(in[1048]), .B(n4134), .Z(n2647) );
  NAND U3773 ( .A(n4071), .B(n2647), .Z(n2473) );
  XNOR U3774 ( .A(n4072), .B(n2473), .Z(out[15]) );
  XNOR U3775 ( .A(in[697]), .B(n3819), .Z(n2695) );
  XOR U3776 ( .A(in[631]), .B(n3571), .Z(n4670) );
  XNOR U3777 ( .A(in[222]), .B(n3672), .Z(n4667) );
  NAND U3778 ( .A(n4670), .B(n4667), .Z(n2474) );
  XNOR U3779 ( .A(n2695), .B(n2474), .Z(out[160]) );
  XNOR U3780 ( .A(in[698]), .B(n3821), .Z(n2697) );
  XOR U3781 ( .A(in[632]), .B(n3579), .Z(n4714) );
  XNOR U3782 ( .A(in[223]), .B(n3676), .Z(n4711) );
  NAND U3783 ( .A(n4714), .B(n4711), .Z(n2475) );
  XNOR U3784 ( .A(n2697), .B(n2475), .Z(out[161]) );
  XNOR U3785 ( .A(in[699]), .B(n3823), .Z(n2701) );
  XOR U3786 ( .A(in[633]), .B(n3583), .Z(n4758) );
  XNOR U3787 ( .A(in[224]), .B(n3680), .Z(n4755) );
  NAND U3788 ( .A(n4758), .B(n4755), .Z(n2476) );
  XNOR U3789 ( .A(n2701), .B(n2476), .Z(out[162]) );
  XNOR U3790 ( .A(in[700]), .B(n3825), .Z(n2703) );
  XOR U3791 ( .A(in[634]), .B(n3587), .Z(n4802) );
  XNOR U3792 ( .A(in[225]), .B(n3684), .Z(n4799) );
  NAND U3793 ( .A(n4802), .B(n4799), .Z(n2477) );
  XNOR U3794 ( .A(n2703), .B(n2477), .Z(out[163]) );
  XOR U3795 ( .A(in[701]), .B(n3827), .Z(n2705) );
  NOR U3796 ( .A(n2549), .B(n2830), .Z(n2478) );
  XNOR U3797 ( .A(n2705), .B(n2478), .Z(out[164]) );
  XOR U3798 ( .A(in[702]), .B(n3833), .Z(n2707) );
  NOR U3799 ( .A(n2551), .B(n2844), .Z(n2479) );
  XNOR U3800 ( .A(n2707), .B(n2479), .Z(out[165]) );
  XOR U3801 ( .A(in[703]), .B(n3835), .Z(n2709) );
  NOR U3802 ( .A(n2554), .B(n2858), .Z(n2480) );
  XNOR U3803 ( .A(n2709), .B(n2480), .Z(out[166]) );
  XOR U3804 ( .A(in[640]), .B(n3837), .Z(n2711) );
  NOR U3805 ( .A(n2556), .B(n2872), .Z(n2481) );
  XNOR U3806 ( .A(n2711), .B(n2481), .Z(out[167]) );
  XOR U3807 ( .A(in[641]), .B(n3839), .Z(n2713) );
  NOR U3808 ( .A(n2558), .B(n2888), .Z(n2482) );
  XNOR U3809 ( .A(n2713), .B(n2482), .Z(out[168]) );
  XOR U3810 ( .A(in[642]), .B(n3841), .Z(n2715) );
  NOR U3811 ( .A(n2560), .B(n2902), .Z(n2483) );
  XNOR U3812 ( .A(n2715), .B(n2483), .Z(out[169]) );
  XNOR U3813 ( .A(in[1426]), .B(n3641), .Z(n4109) );
  XOR U3814 ( .A(in[1049]), .B(n4137), .Z(n2650) );
  NAND U3815 ( .A(n4109), .B(n2650), .Z(n2484) );
  XNOR U3816 ( .A(n4110), .B(n2484), .Z(out[16]) );
  XOR U3817 ( .A(in[643]), .B(n3843), .Z(n2717) );
  NOR U3818 ( .A(n2562), .B(n2916), .Z(n2485) );
  XNOR U3819 ( .A(n2717), .B(n2485), .Z(out[170]) );
  XOR U3820 ( .A(in[644]), .B(n3845), .Z(n2719) );
  NOR U3821 ( .A(n2564), .B(n2930), .Z(n2486) );
  XNOR U3822 ( .A(n2719), .B(n2486), .Z(out[171]) );
  XOR U3823 ( .A(in[645]), .B(n3847), .Z(n2725) );
  NOR U3824 ( .A(n2566), .B(n2946), .Z(n2487) );
  XNOR U3825 ( .A(n2725), .B(n2487), .Z(out[172]) );
  XOR U3826 ( .A(in[646]), .B(n3849), .Z(n2727) );
  NOR U3827 ( .A(n2568), .B(n2970), .Z(n2488) );
  XNOR U3828 ( .A(n2727), .B(n2488), .Z(out[173]) );
  XOR U3829 ( .A(in[647]), .B(n3851), .Z(n2729) );
  NOR U3830 ( .A(n2570), .B(n2994), .Z(n2489) );
  XNOR U3831 ( .A(n2729), .B(n2489), .Z(out[174]) );
  XOR U3832 ( .A(in[648]), .B(n3855), .Z(n2731) );
  NOR U3833 ( .A(n2572), .B(n3018), .Z(n2490) );
  XNOR U3834 ( .A(n2731), .B(n2490), .Z(out[175]) );
  XOR U3835 ( .A(in[649]), .B(n3857), .Z(n2733) );
  NOR U3836 ( .A(n2575), .B(n3042), .Z(n2491) );
  XNOR U3837 ( .A(n2733), .B(n2491), .Z(out[176]) );
  XOR U3838 ( .A(in[650]), .B(n3859), .Z(n2735) );
  NOR U3839 ( .A(n2577), .B(n3066), .Z(n2492) );
  XNOR U3840 ( .A(n2735), .B(n2492), .Z(out[177]) );
  XOR U3841 ( .A(in[651]), .B(n3861), .Z(n2737) );
  NOR U3842 ( .A(n2579), .B(n3092), .Z(n2493) );
  XNOR U3843 ( .A(n2737), .B(n2493), .Z(out[178]) );
  XOR U3844 ( .A(in[652]), .B(n3863), .Z(n2739) );
  NOR U3845 ( .A(n2581), .B(n3116), .Z(n2494) );
  XNOR U3846 ( .A(n2739), .B(n2494), .Z(out[179]) );
  XNOR U3847 ( .A(in[1427]), .B(n3645), .Z(n4143) );
  XOR U3848 ( .A(in[1050]), .B(n4140), .Z(n2653) );
  NAND U3849 ( .A(n4143), .B(n2653), .Z(n2495) );
  XNOR U3850 ( .A(n4144), .B(n2495), .Z(out[17]) );
  XOR U3851 ( .A(in[653]), .B(n3865), .Z(n2741) );
  NOR U3852 ( .A(n2583), .B(n3140), .Z(n2496) );
  XNOR U3853 ( .A(n2741), .B(n2496), .Z(out[180]) );
  XOR U3854 ( .A(in[654]), .B(n3867), .Z(n2743) );
  NOR U3855 ( .A(n2585), .B(n3164), .Z(n2497) );
  XNOR U3856 ( .A(n2743), .B(n2497), .Z(out[181]) );
  XOR U3857 ( .A(in[655]), .B(n3869), .Z(n2747) );
  NOR U3858 ( .A(n2587), .B(n3188), .Z(n2498) );
  XNOR U3859 ( .A(n2747), .B(n2498), .Z(out[182]) );
  XOR U3860 ( .A(in[656]), .B(n3871), .Z(n2749) );
  NOR U3861 ( .A(n2589), .B(n3212), .Z(n2499) );
  XNOR U3862 ( .A(n2749), .B(n2499), .Z(out[183]) );
  XOR U3863 ( .A(in[657]), .B(n3873), .Z(n2751) );
  NOR U3864 ( .A(n2591), .B(n3236), .Z(n2500) );
  XNOR U3865 ( .A(n2751), .B(n2500), .Z(out[184]) );
  XOR U3866 ( .A(in[658]), .B(n3877), .Z(n2753) );
  NOR U3867 ( .A(n2593), .B(n3268), .Z(n2501) );
  XNOR U3868 ( .A(n2753), .B(n2501), .Z(out[185]) );
  XOR U3869 ( .A(in[659]), .B(n3879), .Z(n2755) );
  NOR U3870 ( .A(n2596), .B(n3312), .Z(n2502) );
  XNOR U3871 ( .A(n2755), .B(n2502), .Z(out[186]) );
  XOR U3872 ( .A(in[660]), .B(n3881), .Z(n2757) );
  NOR U3873 ( .A(n2598), .B(n3356), .Z(n2503) );
  XNOR U3874 ( .A(n2757), .B(n2503), .Z(out[187]) );
  XOR U3875 ( .A(in[661]), .B(n3883), .Z(n2759) );
  NOR U3876 ( .A(n2600), .B(n3402), .Z(n2504) );
  XNOR U3877 ( .A(n2759), .B(n2504), .Z(out[188]) );
  XOR U3878 ( .A(in[662]), .B(n3885), .Z(n2761) );
  NOR U3879 ( .A(n2602), .B(n3446), .Z(n2505) );
  XNOR U3880 ( .A(n2761), .B(n2505), .Z(out[189]) );
  XNOR U3881 ( .A(in[1428]), .B(n3649), .Z(n4177) );
  XOR U3882 ( .A(in[1051]), .B(n4147), .Z(n2656) );
  NAND U3883 ( .A(n4177), .B(n2656), .Z(n2506) );
  XNOR U3884 ( .A(n4178), .B(n2506), .Z(out[18]) );
  XOR U3885 ( .A(in[663]), .B(n3887), .Z(n2763) );
  NOR U3886 ( .A(n2604), .B(n3490), .Z(n2507) );
  XNOR U3887 ( .A(n2763), .B(n2507), .Z(out[190]) );
  XOR U3888 ( .A(in[664]), .B(n3889), .Z(n2765) );
  NOR U3889 ( .A(n2606), .B(n3534), .Z(n2508) );
  XNOR U3890 ( .A(n2765), .B(n2508), .Z(out[191]) );
  OR U3891 ( .A(n2609), .B(n3578), .Z(n2509) );
  XNOR U3892 ( .A(n2608), .B(n2509), .Z(out[192]) );
  XOR U3893 ( .A(in[1034]), .B(n4088), .Z(n2612) );
  NOR U3894 ( .A(n2611), .B(n3622), .Z(n2510) );
  XNOR U3895 ( .A(n2612), .B(n2510), .Z(out[193]) );
  XOR U3896 ( .A(in[1035]), .B(n4091), .Z(n2723) );
  NOR U3897 ( .A(n2614), .B(n3666), .Z(n2511) );
  XNOR U3898 ( .A(n2723), .B(n2511), .Z(out[194]) );
  XNOR U3899 ( .A(n4094), .B(in[1036]), .Z(n2873) );
  NOR U3900 ( .A(n2616), .B(n3710), .Z(n2512) );
  XNOR U3901 ( .A(n2873), .B(n2512), .Z(out[195]) );
  XNOR U3902 ( .A(n4097), .B(in[1037]), .Z(n3067) );
  NOR U3903 ( .A(n2619), .B(n3754), .Z(n2513) );
  XNOR U3904 ( .A(n3067), .B(n2513), .Z(out[196]) );
  XNOR U3905 ( .A(n4100), .B(in[1038]), .Z(n3357) );
  NOR U3906 ( .A(n2621), .B(n3798), .Z(n2514) );
  XNOR U3907 ( .A(n3357), .B(n2514), .Z(out[197]) );
  XNOR U3908 ( .A(n4103), .B(in[1039]), .Z(n3799) );
  NOR U3909 ( .A(n2623), .B(n3832), .Z(n2515) );
  XNOR U3910 ( .A(n3799), .B(n2515), .Z(out[198]) );
  XNOR U3911 ( .A(n4106), .B(in[1040]), .Z(n4075) );
  NOR U3912 ( .A(n2625), .B(n3854), .Z(n2516) );
  XNOR U3913 ( .A(n4075), .B(n2516), .Z(out[199]) );
  XNOR U3914 ( .A(in[1429]), .B(n3653), .Z(n4203) );
  XOR U3915 ( .A(in[1052]), .B(n4150), .Z(n2659) );
  NAND U3916 ( .A(n4203), .B(n2659), .Z(n2517) );
  XNOR U3917 ( .A(n4204), .B(n2517), .Z(out[19]) );
  XNOR U3918 ( .A(n3573), .B(in[1411]), .Z(n3619) );
  NANDN U3919 ( .A(n2612), .B(n3619), .Z(n2518) );
  XNOR U3920 ( .A(n3620), .B(n2518), .Z(out[1]) );
  XNOR U3921 ( .A(n4113), .B(in[1041]), .Z(n4359) );
  NOR U3922 ( .A(n2627), .B(n3876), .Z(n2519) );
  XNOR U3923 ( .A(n4359), .B(n2519), .Z(out[200]) );
  XNOR U3924 ( .A(n4116), .B(in[1042]), .Z(n4803) );
  NOR U3925 ( .A(n2629), .B(n3898), .Z(n2520) );
  XNOR U3926 ( .A(n4803), .B(n2520), .Z(out[201]) );
  OR U3927 ( .A(n2632), .B(n3922), .Z(n2521) );
  XNOR U3928 ( .A(n2631), .B(n2521), .Z(out[202]) );
  OR U3929 ( .A(n2635), .B(n3946), .Z(n2522) );
  XNOR U3930 ( .A(n2634), .B(n2522), .Z(out[203]) );
  OR U3931 ( .A(n2638), .B(n3972), .Z(n2523) );
  XNOR U3932 ( .A(n2637), .B(n2523), .Z(out[204]) );
  OR U3933 ( .A(n2641), .B(n4006), .Z(n2524) );
  XNOR U3934 ( .A(n2640), .B(n2524), .Z(out[205]) );
  OR U3935 ( .A(n2645), .B(n4040), .Z(n2525) );
  XNOR U3936 ( .A(n2644), .B(n2525), .Z(out[206]) );
  OR U3937 ( .A(n2648), .B(n4074), .Z(n2526) );
  XNOR U3938 ( .A(n2647), .B(n2526), .Z(out[207]) );
  OR U3939 ( .A(n2651), .B(n4112), .Z(n2527) );
  XNOR U3940 ( .A(n2650), .B(n2527), .Z(out[208]) );
  OR U3941 ( .A(n2654), .B(n4146), .Z(n2528) );
  XNOR U3942 ( .A(n2653), .B(n2528), .Z(out[209]) );
  XNOR U3943 ( .A(in[1430]), .B(n3657), .Z(n4227) );
  XOR U3944 ( .A(in[1053]), .B(n4153), .Z(n2662) );
  NAND U3945 ( .A(n4227), .B(n2662), .Z(n2529) );
  XNOR U3946 ( .A(n4228), .B(n2529), .Z(out[20]) );
  OR U3947 ( .A(n2657), .B(n4180), .Z(n2530) );
  XNOR U3948 ( .A(n2656), .B(n2530), .Z(out[210]) );
  OR U3949 ( .A(n2660), .B(n4206), .Z(n2531) );
  XNOR U3950 ( .A(n2659), .B(n2531), .Z(out[211]) );
  OR U3951 ( .A(n2663), .B(n4230), .Z(n2532) );
  XNOR U3952 ( .A(n2662), .B(n2532), .Z(out[212]) );
  XNOR U3953 ( .A(in[1054]), .B(n4156), .Z(n2666) );
  NOR U3954 ( .A(n2665), .B(n4254), .Z(n2533) );
  XNOR U3955 ( .A(n2666), .B(n2533), .Z(out[213]) );
  XNOR U3956 ( .A(in[1055]), .B(n4159), .Z(n2669) );
  NOR U3957 ( .A(n2668), .B(n4278), .Z(n2534) );
  XNOR U3958 ( .A(n2669), .B(n2534), .Z(out[214]) );
  XNOR U3959 ( .A(in[1056]), .B(n4162), .Z(n2672) );
  NOR U3960 ( .A(n2671), .B(n4302), .Z(n2535) );
  XNOR U3961 ( .A(n2672), .B(n2535), .Z(out[215]) );
  XNOR U3962 ( .A(in[1057]), .B(n4165), .Z(n2676) );
  NOR U3963 ( .A(n2675), .B(n4326), .Z(n2536) );
  XNOR U3964 ( .A(n2676), .B(n2536), .Z(out[216]) );
  XNOR U3965 ( .A(in[1058]), .B(n4168), .Z(n2679) );
  NOR U3966 ( .A(n2678), .B(n4358), .Z(n2537) );
  XNOR U3967 ( .A(n2679), .B(n2537), .Z(out[217]) );
  XNOR U3968 ( .A(in[1059]), .B(n4171), .Z(n2682) );
  NOR U3969 ( .A(n2681), .B(n4406), .Z(n2538) );
  XNOR U3970 ( .A(n2682), .B(n2538), .Z(out[218]) );
  XOR U3971 ( .A(in[1060]), .B(n4174), .Z(n2685) );
  NOR U3972 ( .A(n2684), .B(n4450), .Z(n2539) );
  XNOR U3973 ( .A(n2685), .B(n2539), .Z(out[219]) );
  XNOR U3974 ( .A(in[1431]), .B(n3661), .Z(n4251) );
  NANDN U3975 ( .A(n2666), .B(n4251), .Z(n2540) );
  XNOR U3976 ( .A(n4252), .B(n2540), .Z(out[21]) );
  XOR U3977 ( .A(in[1061]), .B(n4181), .Z(n2699) );
  NOR U3978 ( .A(n2687), .B(n4494), .Z(n2541) );
  XNOR U3979 ( .A(n2699), .B(n2541), .Z(out[220]) );
  XOR U3980 ( .A(in[1062]), .B(n4184), .Z(n2721) );
  NOR U3981 ( .A(n2689), .B(n4538), .Z(n2542) );
  XNOR U3982 ( .A(n2721), .B(n2542), .Z(out[221]) );
  XOR U3983 ( .A(in[1063]), .B(n3963), .Z(n2745) );
  NOR U3984 ( .A(n2691), .B(n4582), .Z(n2543) );
  XNOR U3985 ( .A(n2745), .B(n2543), .Z(out[222]) );
  XOR U3986 ( .A(in[1064]), .B(n3966), .Z(n2767) );
  NOR U3987 ( .A(n2693), .B(n4626), .Z(n2544) );
  XNOR U3988 ( .A(n2767), .B(n2544), .Z(out[223]) );
  XOR U3989 ( .A(in[1065]), .B(n3973), .Z(n2779) );
  NOR U3990 ( .A(n2695), .B(n4670), .Z(n2545) );
  XNOR U3991 ( .A(n2779), .B(n2545), .Z(out[224]) );
  XOR U3992 ( .A(in[1066]), .B(n3976), .Z(n2791) );
  NOR U3993 ( .A(n2697), .B(n4714), .Z(n2546) );
  XNOR U3994 ( .A(n2791), .B(n2546), .Z(out[225]) );
  XOR U3995 ( .A(in[1067]), .B(n3979), .Z(n2803) );
  NOR U3996 ( .A(n2701), .B(n4758), .Z(n2547) );
  XNOR U3997 ( .A(n2803), .B(n2547), .Z(out[226]) );
  XOR U3998 ( .A(in[1068]), .B(n3982), .Z(n2815) );
  NOR U3999 ( .A(n2703), .B(n4802), .Z(n2548) );
  XNOR U4000 ( .A(n2815), .B(n2548), .Z(out[227]) );
  XNOR U4001 ( .A(in[1069]), .B(n3985), .Z(n2828) );
  NAND U4002 ( .A(n2705), .B(n2549), .Z(n2550) );
  XNOR U4003 ( .A(n2828), .B(n2550), .Z(out[228]) );
  XNOR U4004 ( .A(in[1070]), .B(n3988), .Z(n2842) );
  NAND U4005 ( .A(n2707), .B(n2551), .Z(n2552) );
  XNOR U4006 ( .A(n2842), .B(n2552), .Z(out[229]) );
  XNOR U4007 ( .A(in[1432]), .B(n3669), .Z(n4275) );
  NANDN U4008 ( .A(n2669), .B(n4275), .Z(n2553) );
  XNOR U4009 ( .A(n4276), .B(n2553), .Z(out[22]) );
  XNOR U4010 ( .A(in[1071]), .B(n3991), .Z(n2856) );
  NAND U4011 ( .A(n2709), .B(n2554), .Z(n2555) );
  XNOR U4012 ( .A(n2856), .B(n2555), .Z(out[230]) );
  XNOR U4013 ( .A(in[1072]), .B(n3994), .Z(n2870) );
  NAND U4014 ( .A(n2711), .B(n2556), .Z(n2557) );
  XNOR U4015 ( .A(n2870), .B(n2557), .Z(out[231]) );
  XNOR U4016 ( .A(in[1073]), .B(n3997), .Z(n2886) );
  NAND U4017 ( .A(n2713), .B(n2558), .Z(n2559) );
  XNOR U4018 ( .A(n2886), .B(n2559), .Z(out[232]) );
  XNOR U4019 ( .A(in[1074]), .B(n4000), .Z(n2900) );
  NAND U4020 ( .A(n2715), .B(n2560), .Z(n2561) );
  XNOR U4021 ( .A(n2900), .B(n2561), .Z(out[233]) );
  XNOR U4022 ( .A(in[1075]), .B(n4007), .Z(n2914) );
  NAND U4023 ( .A(n2717), .B(n2562), .Z(n2563) );
  XNOR U4024 ( .A(n2914), .B(n2563), .Z(out[234]) );
  XNOR U4025 ( .A(in[1076]), .B(n4010), .Z(n2928) );
  NAND U4026 ( .A(n2719), .B(n2564), .Z(n2565) );
  XNOR U4027 ( .A(n2928), .B(n2565), .Z(out[235]) );
  XNOR U4028 ( .A(in[1077]), .B(n4013), .Z(n2944) );
  NAND U4029 ( .A(n2725), .B(n2566), .Z(n2567) );
  XNOR U4030 ( .A(n2944), .B(n2567), .Z(out[236]) );
  XNOR U4031 ( .A(in[1078]), .B(n4016), .Z(n2968) );
  NAND U4032 ( .A(n2727), .B(n2568), .Z(n2569) );
  XNOR U4033 ( .A(n2968), .B(n2569), .Z(out[237]) );
  XNOR U4034 ( .A(in[1079]), .B(n4019), .Z(n2992) );
  NAND U4035 ( .A(n2729), .B(n2570), .Z(n2571) );
  XNOR U4036 ( .A(n2992), .B(n2571), .Z(out[238]) );
  XNOR U4037 ( .A(in[1080]), .B(n4022), .Z(n3016) );
  NAND U4038 ( .A(n2731), .B(n2572), .Z(n2573) );
  XNOR U4039 ( .A(n3016), .B(n2573), .Z(out[239]) );
  XNOR U4040 ( .A(in[1433]), .B(n3673), .Z(n4299) );
  NANDN U4041 ( .A(n2672), .B(n4299), .Z(n2574) );
  XNOR U4042 ( .A(n4300), .B(n2574), .Z(out[23]) );
  XNOR U4043 ( .A(in[1081]), .B(n4025), .Z(n3040) );
  NAND U4044 ( .A(n2733), .B(n2575), .Z(n2576) );
  XNOR U4045 ( .A(n3040), .B(n2576), .Z(out[240]) );
  XNOR U4046 ( .A(in[1082]), .B(n4028), .Z(n3064) );
  NAND U4047 ( .A(n2735), .B(n2577), .Z(n2578) );
  XNOR U4048 ( .A(n3064), .B(n2578), .Z(out[241]) );
  XNOR U4049 ( .A(in[1083]), .B(n4031), .Z(n3090) );
  NAND U4050 ( .A(n2737), .B(n2579), .Z(n2580) );
  XNOR U4051 ( .A(n3090), .B(n2580), .Z(out[242]) );
  XNOR U4052 ( .A(in[1084]), .B(n4034), .Z(n3114) );
  NAND U4053 ( .A(n2739), .B(n2581), .Z(n2582) );
  XNOR U4054 ( .A(n3114), .B(n2582), .Z(out[243]) );
  XNOR U4055 ( .A(in[1085]), .B(n4041), .Z(n3138) );
  NAND U4056 ( .A(n2741), .B(n2583), .Z(n2584) );
  XNOR U4057 ( .A(n3138), .B(n2584), .Z(out[244]) );
  XNOR U4058 ( .A(in[1086]), .B(n4044), .Z(n3162) );
  NAND U4059 ( .A(n2743), .B(n2585), .Z(n2586) );
  XNOR U4060 ( .A(n3162), .B(n2586), .Z(out[245]) );
  XNOR U4061 ( .A(in[1087]), .B(n4047), .Z(n3186) );
  NAND U4062 ( .A(n2747), .B(n2587), .Z(n2588) );
  XNOR U4063 ( .A(n3186), .B(n2588), .Z(out[246]) );
  XNOR U4064 ( .A(in[1024]), .B(n4050), .Z(n3210) );
  NAND U4065 ( .A(n2749), .B(n2589), .Z(n2590) );
  XNOR U4066 ( .A(n3210), .B(n2590), .Z(out[247]) );
  XNOR U4067 ( .A(in[1025]), .B(n4053), .Z(n3234) );
  NAND U4068 ( .A(n2751), .B(n2591), .Z(n2592) );
  XNOR U4069 ( .A(n3234), .B(n2592), .Z(out[248]) );
  XNOR U4070 ( .A(in[1026]), .B(n4056), .Z(n3266) );
  NAND U4071 ( .A(n2753), .B(n2593), .Z(n2594) );
  XNOR U4072 ( .A(n3266), .B(n2594), .Z(out[249]) );
  XNOR U4073 ( .A(in[1434]), .B(n3677), .Z(n4323) );
  NANDN U4074 ( .A(n2676), .B(n4323), .Z(n2595) );
  XNOR U4075 ( .A(n4324), .B(n2595), .Z(out[24]) );
  XNOR U4076 ( .A(in[1027]), .B(n4059), .Z(n3310) );
  NAND U4077 ( .A(n2755), .B(n2596), .Z(n2597) );
  XNOR U4078 ( .A(n3310), .B(n2597), .Z(out[250]) );
  XNOR U4079 ( .A(in[1028]), .B(n4062), .Z(n3354) );
  NAND U4080 ( .A(n2757), .B(n2598), .Z(n2599) );
  XNOR U4081 ( .A(n3354), .B(n2599), .Z(out[251]) );
  XNOR U4082 ( .A(in[1029]), .B(n4065), .Z(n3400) );
  NAND U4083 ( .A(n2759), .B(n2600), .Z(n2601) );
  XNOR U4084 ( .A(n3400), .B(n2601), .Z(out[252]) );
  XNOR U4085 ( .A(in[1030]), .B(n4068), .Z(n3444) );
  NAND U4086 ( .A(n2761), .B(n2602), .Z(n2603) );
  XNOR U4087 ( .A(n3444), .B(n2603), .Z(out[253]) );
  XNOR U4088 ( .A(in[1031]), .B(n4079), .Z(n3488) );
  NAND U4089 ( .A(n2763), .B(n2604), .Z(n2605) );
  XNOR U4090 ( .A(n3488), .B(n2605), .Z(out[254]) );
  XNOR U4091 ( .A(in[1032]), .B(n4082), .Z(n3532) );
  NAND U4092 ( .A(n2765), .B(n2606), .Z(n2607) );
  XNOR U4093 ( .A(n3532), .B(n2607), .Z(out[255]) );
  ANDN U4094 ( .B(n2609), .A(n2608), .Z(n2610) );
  XNOR U4095 ( .A(n3575), .B(n2610), .Z(out[256]) );
  AND U4096 ( .A(n2612), .B(n2611), .Z(n2613) );
  XNOR U4097 ( .A(n3619), .B(n2613), .Z(out[257]) );
  XOR U4098 ( .A(n3581), .B(in[1412]), .Z(n3664) );
  NAND U4099 ( .A(n2723), .B(n2614), .Z(n2615) );
  XNOR U4100 ( .A(n3664), .B(n2615), .Z(out[258]) );
  XOR U4101 ( .A(n3585), .B(in[1413]), .Z(n3708) );
  NAND U4102 ( .A(n2873), .B(n2616), .Z(n2617) );
  XNOR U4103 ( .A(n3708), .B(n2617), .Z(out[259]) );
  XNOR U4104 ( .A(in[1435]), .B(n3681), .Z(n4355) );
  NANDN U4105 ( .A(n2679), .B(n4355), .Z(n2618) );
  XNOR U4106 ( .A(n4356), .B(n2618), .Z(out[25]) );
  XOR U4107 ( .A(n3589), .B(in[1414]), .Z(n3752) );
  NAND U4108 ( .A(n3067), .B(n2619), .Z(n2620) );
  XNOR U4109 ( .A(n3752), .B(n2620), .Z(out[260]) );
  XOR U4110 ( .A(n3593), .B(in[1415]), .Z(n3796) );
  NAND U4111 ( .A(n3357), .B(n2621), .Z(n2622) );
  XNOR U4112 ( .A(n3796), .B(n2622), .Z(out[261]) );
  XOR U4113 ( .A(n3597), .B(in[1416]), .Z(n3830) );
  NAND U4114 ( .A(n3799), .B(n2623), .Z(n2624) );
  XNOR U4115 ( .A(n3830), .B(n2624), .Z(out[262]) );
  XOR U4116 ( .A(in[1417]), .B(n3601), .Z(n4076) );
  NAND U4117 ( .A(n4075), .B(n2625), .Z(n2626) );
  XNOR U4118 ( .A(n4076), .B(n2626), .Z(out[263]) );
  XOR U4119 ( .A(n3605), .B(in[1418]), .Z(n4360) );
  NAND U4120 ( .A(n4359), .B(n2627), .Z(n2628) );
  XNOR U4121 ( .A(n4360), .B(n2628), .Z(out[264]) );
  XOR U4122 ( .A(n3609), .B(in[1419]), .Z(n4804) );
  NAND U4123 ( .A(n4803), .B(n2629), .Z(n2630) );
  XNOR U4124 ( .A(n4804), .B(n2630), .Z(out[265]) );
  ANDN U4125 ( .B(n2632), .A(n2631), .Z(n2633) );
  XNOR U4126 ( .A(n3919), .B(n2633), .Z(out[266]) );
  ANDN U4127 ( .B(n2635), .A(n2634), .Z(n2636) );
  XNOR U4128 ( .A(n3943), .B(n2636), .Z(out[267]) );
  ANDN U4129 ( .B(n2638), .A(n2637), .Z(n2639) );
  XNOR U4130 ( .A(n3969), .B(n2639), .Z(out[268]) );
  ANDN U4131 ( .B(n2641), .A(n2640), .Z(n2642) );
  XNOR U4132 ( .A(n4003), .B(n2642), .Z(out[269]) );
  XNOR U4133 ( .A(in[1436]), .B(n3685), .Z(n4403) );
  NANDN U4134 ( .A(n2682), .B(n4403), .Z(n2643) );
  XNOR U4135 ( .A(n4404), .B(n2643), .Z(out[26]) );
  ANDN U4136 ( .B(n2645), .A(n2644), .Z(n2646) );
  XNOR U4137 ( .A(n4037), .B(n2646), .Z(out[270]) );
  ANDN U4138 ( .B(n2648), .A(n2647), .Z(n2649) );
  XNOR U4139 ( .A(n4071), .B(n2649), .Z(out[271]) );
  ANDN U4140 ( .B(n2651), .A(n2650), .Z(n2652) );
  XNOR U4141 ( .A(n4109), .B(n2652), .Z(out[272]) );
  ANDN U4142 ( .B(n2654), .A(n2653), .Z(n2655) );
  XNOR U4143 ( .A(n4143), .B(n2655), .Z(out[273]) );
  ANDN U4144 ( .B(n2657), .A(n2656), .Z(n2658) );
  XNOR U4145 ( .A(n4177), .B(n2658), .Z(out[274]) );
  ANDN U4146 ( .B(n2660), .A(n2659), .Z(n2661) );
  XNOR U4147 ( .A(n4203), .B(n2661), .Z(out[275]) );
  ANDN U4148 ( .B(n2663), .A(n2662), .Z(n2664) );
  XNOR U4149 ( .A(n4227), .B(n2664), .Z(out[276]) );
  AND U4150 ( .A(n2666), .B(n2665), .Z(n2667) );
  XNOR U4151 ( .A(n4251), .B(n2667), .Z(out[277]) );
  AND U4152 ( .A(n2669), .B(n2668), .Z(n2670) );
  XNOR U4153 ( .A(n4275), .B(n2670), .Z(out[278]) );
  AND U4154 ( .A(n2672), .B(n2671), .Z(n2673) );
  XNOR U4155 ( .A(n4299), .B(n2673), .Z(out[279]) );
  XNOR U4156 ( .A(in[1437]), .B(n3689), .Z(n4447) );
  NANDN U4157 ( .A(n2685), .B(n4447), .Z(n2674) );
  XNOR U4158 ( .A(n4448), .B(n2674), .Z(out[27]) );
  AND U4159 ( .A(n2676), .B(n2675), .Z(n2677) );
  XNOR U4160 ( .A(n4323), .B(n2677), .Z(out[280]) );
  AND U4161 ( .A(n2679), .B(n2678), .Z(n2680) );
  XNOR U4162 ( .A(n4355), .B(n2680), .Z(out[281]) );
  AND U4163 ( .A(n2682), .B(n2681), .Z(n2683) );
  XNOR U4164 ( .A(n4403), .B(n2683), .Z(out[282]) );
  AND U4165 ( .A(n2685), .B(n2684), .Z(n2686) );
  XNOR U4166 ( .A(n4447), .B(n2686), .Z(out[283]) );
  XOR U4167 ( .A(in[1438]), .B(n3693), .Z(n4492) );
  NAND U4168 ( .A(n2699), .B(n2687), .Z(n2688) );
  XNOR U4169 ( .A(n4492), .B(n2688), .Z(out[284]) );
  XOR U4170 ( .A(in[1439]), .B(n3697), .Z(n4536) );
  NAND U4171 ( .A(n2721), .B(n2689), .Z(n2690) );
  XNOR U4172 ( .A(n4536), .B(n2690), .Z(out[285]) );
  XOR U4173 ( .A(in[1440]), .B(n3701), .Z(n4580) );
  NAND U4174 ( .A(n2745), .B(n2691), .Z(n2692) );
  XNOR U4175 ( .A(n4580), .B(n2692), .Z(out[286]) );
  XOR U4176 ( .A(in[1441]), .B(n3705), .Z(n4624) );
  NAND U4177 ( .A(n2767), .B(n2693), .Z(n2694) );
  XNOR U4178 ( .A(n4624), .B(n2694), .Z(out[287]) );
  XOR U4179 ( .A(in[1442]), .B(n3713), .Z(n4668) );
  NAND U4180 ( .A(n2779), .B(n2695), .Z(n2696) );
  XNOR U4181 ( .A(n4668), .B(n2696), .Z(out[288]) );
  XOR U4182 ( .A(in[1443]), .B(n3717), .Z(n4712) );
  NAND U4183 ( .A(n2791), .B(n2697), .Z(n2698) );
  XNOR U4184 ( .A(n4712), .B(n2698), .Z(out[289]) );
  OR U4185 ( .A(n4492), .B(n2699), .Z(n2700) );
  XNOR U4186 ( .A(n4491), .B(n2700), .Z(out[28]) );
  XOR U4187 ( .A(in[1444]), .B(n3721), .Z(n4756) );
  NAND U4188 ( .A(n2803), .B(n2701), .Z(n2702) );
  XNOR U4189 ( .A(n4756), .B(n2702), .Z(out[290]) );
  XOR U4190 ( .A(in[1445]), .B(n3725), .Z(n4800) );
  NAND U4191 ( .A(n2815), .B(n2703), .Z(n2704) );
  XNOR U4192 ( .A(n4800), .B(n2704), .Z(out[291]) );
  OR U4193 ( .A(n2828), .B(n2705), .Z(n2706) );
  XNOR U4194 ( .A(n2827), .B(n2706), .Z(out[292]) );
  OR U4195 ( .A(n2842), .B(n2707), .Z(n2708) );
  XNOR U4196 ( .A(n2841), .B(n2708), .Z(out[293]) );
  OR U4197 ( .A(n2856), .B(n2709), .Z(n2710) );
  XNOR U4198 ( .A(n2855), .B(n2710), .Z(out[294]) );
  OR U4199 ( .A(n2870), .B(n2711), .Z(n2712) );
  XNOR U4200 ( .A(n2869), .B(n2712), .Z(out[295]) );
  OR U4201 ( .A(n2886), .B(n2713), .Z(n2714) );
  XNOR U4202 ( .A(n2885), .B(n2714), .Z(out[296]) );
  OR U4203 ( .A(n2900), .B(n2715), .Z(n2716) );
  XNOR U4204 ( .A(n2899), .B(n2716), .Z(out[297]) );
  OR U4205 ( .A(n2914), .B(n2717), .Z(n2718) );
  XNOR U4206 ( .A(n2913), .B(n2718), .Z(out[298]) );
  OR U4207 ( .A(n2928), .B(n2719), .Z(n2720) );
  XNOR U4208 ( .A(n2927), .B(n2720), .Z(out[299]) );
  OR U4209 ( .A(n4536), .B(n2721), .Z(n2722) );
  XNOR U4210 ( .A(n4535), .B(n2722), .Z(out[29]) );
  OR U4211 ( .A(n3664), .B(n2723), .Z(n2724) );
  XNOR U4212 ( .A(n3663), .B(n2724), .Z(out[2]) );
  OR U4213 ( .A(n2944), .B(n2725), .Z(n2726) );
  XNOR U4214 ( .A(n2943), .B(n2726), .Z(out[300]) );
  OR U4215 ( .A(n2968), .B(n2727), .Z(n2728) );
  XNOR U4216 ( .A(n2967), .B(n2728), .Z(out[301]) );
  OR U4217 ( .A(n2992), .B(n2729), .Z(n2730) );
  XNOR U4218 ( .A(n2991), .B(n2730), .Z(out[302]) );
  OR U4219 ( .A(n3016), .B(n2731), .Z(n2732) );
  XNOR U4220 ( .A(n3015), .B(n2732), .Z(out[303]) );
  OR U4221 ( .A(n3040), .B(n2733), .Z(n2734) );
  XNOR U4222 ( .A(n3039), .B(n2734), .Z(out[304]) );
  OR U4223 ( .A(n3064), .B(n2735), .Z(n2736) );
  XNOR U4224 ( .A(n3063), .B(n2736), .Z(out[305]) );
  OR U4225 ( .A(n3090), .B(n2737), .Z(n2738) );
  XNOR U4226 ( .A(n3089), .B(n2738), .Z(out[306]) );
  OR U4227 ( .A(n3114), .B(n2739), .Z(n2740) );
  XNOR U4228 ( .A(n3113), .B(n2740), .Z(out[307]) );
  OR U4229 ( .A(n3138), .B(n2741), .Z(n2742) );
  XNOR U4230 ( .A(n3137), .B(n2742), .Z(out[308]) );
  OR U4231 ( .A(n3162), .B(n2743), .Z(n2744) );
  XNOR U4232 ( .A(n3161), .B(n2744), .Z(out[309]) );
  OR U4233 ( .A(n4580), .B(n2745), .Z(n2746) );
  XNOR U4234 ( .A(n4579), .B(n2746), .Z(out[30]) );
  OR U4235 ( .A(n3186), .B(n2747), .Z(n2748) );
  XNOR U4236 ( .A(n3185), .B(n2748), .Z(out[310]) );
  OR U4237 ( .A(n3210), .B(n2749), .Z(n2750) );
  XNOR U4238 ( .A(n3209), .B(n2750), .Z(out[311]) );
  OR U4239 ( .A(n3234), .B(n2751), .Z(n2752) );
  XNOR U4240 ( .A(n3233), .B(n2752), .Z(out[312]) );
  OR U4241 ( .A(n3266), .B(n2753), .Z(n2754) );
  XNOR U4242 ( .A(n3265), .B(n2754), .Z(out[313]) );
  OR U4243 ( .A(n3310), .B(n2755), .Z(n2756) );
  XNOR U4244 ( .A(n3309), .B(n2756), .Z(out[314]) );
  OR U4245 ( .A(n3354), .B(n2757), .Z(n2758) );
  XNOR U4246 ( .A(n3353), .B(n2758), .Z(out[315]) );
  OR U4247 ( .A(n3400), .B(n2759), .Z(n2760) );
  XNOR U4248 ( .A(n3399), .B(n2760), .Z(out[316]) );
  OR U4249 ( .A(n3444), .B(n2761), .Z(n2762) );
  XNOR U4250 ( .A(n3443), .B(n2762), .Z(out[317]) );
  OR U4251 ( .A(n3488), .B(n2763), .Z(n2764) );
  XNOR U4252 ( .A(n3487), .B(n2764), .Z(out[318]) );
  OR U4253 ( .A(n3532), .B(n2765), .Z(n2766) );
  XNOR U4254 ( .A(n3531), .B(n2766), .Z(out[319]) );
  OR U4255 ( .A(n4624), .B(n2767), .Z(n2768) );
  XNOR U4256 ( .A(n4623), .B(n2768), .Z(out[31]) );
  XNOR U4257 ( .A(in[72]), .B(n4082), .Z(n2939) );
  XOR U4258 ( .A(in[1317]), .B(n3917), .Z(n3252) );
  XOR U4259 ( .A(in[1244]), .B(n3735), .Z(n3249) );
  NAND U4260 ( .A(n3252), .B(n3249), .Z(n2769) );
  XNOR U4261 ( .A(n2939), .B(n2769), .Z(out[320]) );
  XNOR U4262 ( .A(in[73]), .B(n4085), .Z(n2941) );
  XOR U4263 ( .A(in[1318]), .B(n3923), .Z(n3256) );
  XOR U4264 ( .A(in[1245]), .B(n3739), .Z(n3253) );
  NAND U4265 ( .A(n3256), .B(n3253), .Z(n2770) );
  XNOR U4266 ( .A(n2941), .B(n2770), .Z(out[321]) );
  XNOR U4267 ( .A(in[74]), .B(n4088), .Z(n2947) );
  XOR U4268 ( .A(in[1319]), .B(n3925), .Z(n3260) );
  XOR U4269 ( .A(in[1246]), .B(n3743), .Z(n3257) );
  NAND U4270 ( .A(n3260), .B(n3257), .Z(n2771) );
  XNOR U4271 ( .A(n2947), .B(n2771), .Z(out[322]) );
  XNOR U4272 ( .A(in[75]), .B(n4091), .Z(n2949) );
  XOR U4273 ( .A(in[1320]), .B(n3927), .Z(n3264) );
  XOR U4274 ( .A(in[1247]), .B(n3747), .Z(n3261) );
  NAND U4275 ( .A(n3264), .B(n3261), .Z(n2772) );
  XNOR U4276 ( .A(n2949), .B(n2772), .Z(out[323]) );
  XOR U4277 ( .A(n4094), .B(in[76]), .Z(n2951) );
  XOR U4278 ( .A(in[1321]), .B(n3929), .Z(n3272) );
  XOR U4279 ( .A(in[1248]), .B(n3755), .Z(n3269) );
  NAND U4280 ( .A(n3272), .B(n3269), .Z(n2773) );
  XNOR U4281 ( .A(n2951), .B(n2773), .Z(out[324]) );
  XOR U4282 ( .A(n4097), .B(in[77]), .Z(n2953) );
  XOR U4283 ( .A(in[1322]), .B(n3931), .Z(n3276) );
  XOR U4284 ( .A(in[1249]), .B(n3759), .Z(n3273) );
  NAND U4285 ( .A(n3276), .B(n3273), .Z(n2774) );
  XNOR U4286 ( .A(n2953), .B(n2774), .Z(out[325]) );
  XOR U4287 ( .A(n4100), .B(in[78]), .Z(n2955) );
  XOR U4288 ( .A(in[1323]), .B(n3933), .Z(n3280) );
  XOR U4289 ( .A(in[1250]), .B(n3763), .Z(n3277) );
  NAND U4290 ( .A(n3280), .B(n3277), .Z(n2775) );
  XNOR U4291 ( .A(n2955), .B(n2775), .Z(out[326]) );
  XOR U4292 ( .A(n4103), .B(in[79]), .Z(n2957) );
  XOR U4293 ( .A(in[1324]), .B(n3935), .Z(n3284) );
  XOR U4294 ( .A(in[1251]), .B(n3767), .Z(n3281) );
  NAND U4295 ( .A(n3284), .B(n3281), .Z(n2776) );
  XNOR U4296 ( .A(n2957), .B(n2776), .Z(out[327]) );
  XOR U4297 ( .A(n4106), .B(in[80]), .Z(n2959) );
  XOR U4298 ( .A(in[1325]), .B(n3937), .Z(n3288) );
  XOR U4299 ( .A(in[1252]), .B(n3771), .Z(n3285) );
  NAND U4300 ( .A(n3288), .B(n3285), .Z(n2777) );
  XNOR U4301 ( .A(n2959), .B(n2777), .Z(out[328]) );
  XOR U4302 ( .A(n4113), .B(in[81]), .Z(n2961) );
  XOR U4303 ( .A(in[1326]), .B(n3939), .Z(n3292) );
  XNOR U4304 ( .A(in[1253]), .B(n3775), .Z(n3289) );
  NAND U4305 ( .A(n3292), .B(n3289), .Z(n2778) );
  XNOR U4306 ( .A(n2961), .B(n2778), .Z(out[329]) );
  OR U4307 ( .A(n4668), .B(n2779), .Z(n2780) );
  XNOR U4308 ( .A(n4667), .B(n2780), .Z(out[32]) );
  XOR U4309 ( .A(n4116), .B(in[82]), .Z(n2963) );
  XOR U4310 ( .A(in[1327]), .B(n3941), .Z(n3296) );
  XNOR U4311 ( .A(in[1254]), .B(n3779), .Z(n3293) );
  NAND U4312 ( .A(n3296), .B(n3293), .Z(n2781) );
  XNOR U4313 ( .A(n2963), .B(n2781), .Z(out[330]) );
  XOR U4314 ( .A(n4119), .B(in[83]), .Z(n2965) );
  XOR U4315 ( .A(in[1328]), .B(n3947), .Z(n3300) );
  XNOR U4316 ( .A(in[1255]), .B(n3783), .Z(n3297) );
  NAND U4317 ( .A(n3300), .B(n3297), .Z(n2782) );
  XNOR U4318 ( .A(n2965), .B(n2782), .Z(out[331]) );
  XOR U4319 ( .A(in[84]), .B(n4122), .Z(n2971) );
  XOR U4320 ( .A(in[1329]), .B(n3949), .Z(n3304) );
  XNOR U4321 ( .A(in[1256]), .B(n3787), .Z(n3301) );
  NAND U4322 ( .A(n3304), .B(n3301), .Z(n2783) );
  XNOR U4323 ( .A(n2971), .B(n2783), .Z(out[332]) );
  XOR U4324 ( .A(in[85]), .B(n4125), .Z(n2973) );
  XOR U4325 ( .A(in[1330]), .B(n3951), .Z(n3308) );
  XNOR U4326 ( .A(in[1257]), .B(n3791), .Z(n3305) );
  NAND U4327 ( .A(n3308), .B(n3305), .Z(n2784) );
  XNOR U4328 ( .A(n2973), .B(n2784), .Z(out[333]) );
  XOR U4329 ( .A(in[86]), .B(n4128), .Z(n2975) );
  XOR U4330 ( .A(in[1331]), .B(n3953), .Z(n3316) );
  XNOR U4331 ( .A(in[1258]), .B(n3801), .Z(n3313) );
  NAND U4332 ( .A(n3316), .B(n3313), .Z(n2785) );
  XNOR U4333 ( .A(n2975), .B(n2785), .Z(out[334]) );
  XOR U4334 ( .A(in[87]), .B(n4131), .Z(n2977) );
  XOR U4335 ( .A(in[1332]), .B(n3955), .Z(n3320) );
  XNOR U4336 ( .A(in[1259]), .B(n3805), .Z(n3317) );
  NAND U4337 ( .A(n3320), .B(n3317), .Z(n2786) );
  XNOR U4338 ( .A(n2977), .B(n2786), .Z(out[335]) );
  XOR U4339 ( .A(in[88]), .B(n4134), .Z(n2979) );
  XOR U4340 ( .A(in[1333]), .B(n3957), .Z(n3324) );
  XNOR U4341 ( .A(in[1260]), .B(n3809), .Z(n3321) );
  NAND U4342 ( .A(n3324), .B(n3321), .Z(n2787) );
  XNOR U4343 ( .A(n2979), .B(n2787), .Z(out[336]) );
  XOR U4344 ( .A(in[89]), .B(n4137), .Z(n2981) );
  XOR U4345 ( .A(in[1334]), .B(n3959), .Z(n3328) );
  XNOR U4346 ( .A(in[1261]), .B(n3813), .Z(n3325) );
  NAND U4347 ( .A(n3328), .B(n3325), .Z(n2788) );
  XNOR U4348 ( .A(n2981), .B(n2788), .Z(out[337]) );
  XOR U4349 ( .A(in[90]), .B(n4140), .Z(n2983) );
  XOR U4350 ( .A(in[1335]), .B(n3961), .Z(n3332) );
  XNOR U4351 ( .A(in[1262]), .B(n3535), .Z(n3329) );
  NAND U4352 ( .A(n3332), .B(n3329), .Z(n2789) );
  XNOR U4353 ( .A(n2983), .B(n2789), .Z(out[338]) );
  XOR U4354 ( .A(in[91]), .B(n4147), .Z(n2985) );
  XOR U4355 ( .A(in[1336]), .B(n3817), .Z(n3336) );
  XNOR U4356 ( .A(in[1263]), .B(n3539), .Z(n3333) );
  NAND U4357 ( .A(n3336), .B(n3333), .Z(n2790) );
  XNOR U4358 ( .A(n2985), .B(n2790), .Z(out[339]) );
  OR U4359 ( .A(n4712), .B(n2791), .Z(n2792) );
  XNOR U4360 ( .A(n4711), .B(n2792), .Z(out[33]) );
  XOR U4361 ( .A(in[92]), .B(n4150), .Z(n2987) );
  XOR U4362 ( .A(in[1337]), .B(n3819), .Z(n3340) );
  XNOR U4363 ( .A(in[1264]), .B(n3543), .Z(n3337) );
  NAND U4364 ( .A(n3340), .B(n3337), .Z(n2793) );
  XNOR U4365 ( .A(n2987), .B(n2793), .Z(out[340]) );
  XOR U4366 ( .A(in[93]), .B(n4153), .Z(n2989) );
  XOR U4367 ( .A(in[1338]), .B(n3821), .Z(n3344) );
  XNOR U4368 ( .A(in[1265]), .B(n3547), .Z(n3341) );
  NAND U4369 ( .A(n3344), .B(n3341), .Z(n2794) );
  XNOR U4370 ( .A(n2989), .B(n2794), .Z(out[341]) );
  XOR U4371 ( .A(in[94]), .B(n4156), .Z(n2995) );
  XOR U4372 ( .A(in[1339]), .B(n3823), .Z(n3348) );
  XNOR U4373 ( .A(in[1266]), .B(n3551), .Z(n3345) );
  NAND U4374 ( .A(n3348), .B(n3345), .Z(n2795) );
  XNOR U4375 ( .A(n2995), .B(n2795), .Z(out[342]) );
  XOR U4376 ( .A(in[95]), .B(n4159), .Z(n2997) );
  XOR U4377 ( .A(in[1340]), .B(n3825), .Z(n3352) );
  XNOR U4378 ( .A(in[1267]), .B(n3555), .Z(n3349) );
  NAND U4379 ( .A(n3352), .B(n3349), .Z(n2796) );
  XNOR U4380 ( .A(n2997), .B(n2796), .Z(out[343]) );
  XOR U4381 ( .A(in[96]), .B(n4162), .Z(n2999) );
  XOR U4382 ( .A(in[1341]), .B(n3827), .Z(n3362) );
  XNOR U4383 ( .A(in[1268]), .B(n3559), .Z(n3359) );
  NAND U4384 ( .A(n3362), .B(n3359), .Z(n2797) );
  XNOR U4385 ( .A(n2999), .B(n2797), .Z(out[344]) );
  XOR U4386 ( .A(in[97]), .B(n4165), .Z(n3001) );
  XOR U4387 ( .A(in[1342]), .B(n3833), .Z(n3366) );
  XNOR U4388 ( .A(in[1269]), .B(n3563), .Z(n3363) );
  NAND U4389 ( .A(n3366), .B(n3363), .Z(n2798) );
  XNOR U4390 ( .A(n3001), .B(n2798), .Z(out[345]) );
  XOR U4391 ( .A(in[98]), .B(n4168), .Z(n3003) );
  XOR U4392 ( .A(in[1343]), .B(n3835), .Z(n3370) );
  XNOR U4393 ( .A(in[1270]), .B(n3567), .Z(n3367) );
  NAND U4394 ( .A(n3370), .B(n3367), .Z(n2799) );
  XNOR U4395 ( .A(n3003), .B(n2799), .Z(out[346]) );
  XOR U4396 ( .A(in[99]), .B(n4171), .Z(n3005) );
  XOR U4397 ( .A(in[1280]), .B(n3837), .Z(n3374) );
  XNOR U4398 ( .A(in[1271]), .B(n3571), .Z(n3371) );
  NAND U4399 ( .A(n3374), .B(n3371), .Z(n2800) );
  XNOR U4400 ( .A(n3005), .B(n2800), .Z(out[347]) );
  XNOR U4401 ( .A(in[100]), .B(n4174), .Z(n3007) );
  XOR U4402 ( .A(in[1281]), .B(n3839), .Z(n3378) );
  XNOR U4403 ( .A(in[1272]), .B(n3579), .Z(n3375) );
  NAND U4404 ( .A(n3378), .B(n3375), .Z(n2801) );
  XNOR U4405 ( .A(n3007), .B(n2801), .Z(out[348]) );
  XNOR U4406 ( .A(in[101]), .B(n4181), .Z(n3009) );
  XOR U4407 ( .A(in[1282]), .B(n3841), .Z(n3382) );
  XNOR U4408 ( .A(in[1273]), .B(n3583), .Z(n3379) );
  NAND U4409 ( .A(n3382), .B(n3379), .Z(n2802) );
  XNOR U4410 ( .A(n3009), .B(n2802), .Z(out[349]) );
  OR U4411 ( .A(n4756), .B(n2803), .Z(n2804) );
  XNOR U4412 ( .A(n4755), .B(n2804), .Z(out[34]) );
  XNOR U4413 ( .A(in[102]), .B(n4184), .Z(n3011) );
  XOR U4414 ( .A(in[1283]), .B(n3843), .Z(n3386) );
  XNOR U4415 ( .A(in[1274]), .B(n3587), .Z(n3383) );
  NAND U4416 ( .A(n3386), .B(n3383), .Z(n2805) );
  XNOR U4417 ( .A(n3011), .B(n2805), .Z(out[350]) );
  XNOR U4418 ( .A(in[103]), .B(n3963), .Z(n3013) );
  XOR U4419 ( .A(in[1284]), .B(n3845), .Z(n3390) );
  XNOR U4420 ( .A(in[1275]), .B(n3591), .Z(n3387) );
  NAND U4421 ( .A(n3390), .B(n3387), .Z(n2806) );
  XNOR U4422 ( .A(n3013), .B(n2806), .Z(out[351]) );
  XNOR U4423 ( .A(in[104]), .B(n3966), .Z(n3019) );
  XOR U4424 ( .A(in[1285]), .B(n3847), .Z(n3394) );
  XNOR U4425 ( .A(in[1276]), .B(n3595), .Z(n3391) );
  NAND U4426 ( .A(n3394), .B(n3391), .Z(n2807) );
  XNOR U4427 ( .A(n3019), .B(n2807), .Z(out[352]) );
  XNOR U4428 ( .A(in[105]), .B(n3973), .Z(n3021) );
  XOR U4429 ( .A(in[1286]), .B(n3849), .Z(n3398) );
  XNOR U4430 ( .A(in[1277]), .B(n3599), .Z(n3395) );
  NAND U4431 ( .A(n3398), .B(n3395), .Z(n2808) );
  XNOR U4432 ( .A(n3021), .B(n2808), .Z(out[353]) );
  XNOR U4433 ( .A(in[106]), .B(n3976), .Z(n3023) );
  XOR U4434 ( .A(in[1287]), .B(n3851), .Z(n3406) );
  XNOR U4435 ( .A(in[1278]), .B(n3603), .Z(n3403) );
  NAND U4436 ( .A(n3406), .B(n3403), .Z(n2809) );
  XNOR U4437 ( .A(n3023), .B(n2809), .Z(out[354]) );
  XNOR U4438 ( .A(in[107]), .B(n3979), .Z(n3025) );
  XOR U4439 ( .A(in[1288]), .B(n3855), .Z(n3410) );
  XNOR U4440 ( .A(in[1279]), .B(n3607), .Z(n3407) );
  NAND U4441 ( .A(n3410), .B(n3407), .Z(n2810) );
  XNOR U4442 ( .A(n3025), .B(n2810), .Z(out[355]) );
  XNOR U4443 ( .A(in[108]), .B(n3982), .Z(n3027) );
  XOR U4444 ( .A(in[1289]), .B(n3857), .Z(n3414) );
  XNOR U4445 ( .A(in[1216]), .B(n3611), .Z(n3411) );
  NAND U4446 ( .A(n3414), .B(n3411), .Z(n2811) );
  XNOR U4447 ( .A(n3027), .B(n2811), .Z(out[356]) );
  XNOR U4448 ( .A(in[109]), .B(n3985), .Z(n3029) );
  XOR U4449 ( .A(in[1290]), .B(n3859), .Z(n3418) );
  XNOR U4450 ( .A(in[1217]), .B(n3615), .Z(n3415) );
  NAND U4451 ( .A(n3418), .B(n3415), .Z(n2812) );
  XNOR U4452 ( .A(n3029), .B(n2812), .Z(out[357]) );
  XNOR U4453 ( .A(in[110]), .B(n3988), .Z(n3031) );
  XOR U4454 ( .A(in[1291]), .B(n3861), .Z(n3422) );
  XNOR U4455 ( .A(in[1218]), .B(n3623), .Z(n3419) );
  NAND U4456 ( .A(n3422), .B(n3419), .Z(n2813) );
  XNOR U4457 ( .A(n3031), .B(n2813), .Z(out[358]) );
  XNOR U4458 ( .A(in[111]), .B(n3991), .Z(n3033) );
  XOR U4459 ( .A(in[1292]), .B(n3863), .Z(n3426) );
  XNOR U4460 ( .A(in[1219]), .B(n3627), .Z(n3423) );
  NAND U4461 ( .A(n3426), .B(n3423), .Z(n2814) );
  XNOR U4462 ( .A(n3033), .B(n2814), .Z(out[359]) );
  OR U4463 ( .A(n4800), .B(n2815), .Z(n2816) );
  XNOR U4464 ( .A(n4799), .B(n2816), .Z(out[35]) );
  XNOR U4465 ( .A(in[112]), .B(n3994), .Z(n3035) );
  XOR U4466 ( .A(in[1293]), .B(n3865), .Z(n3430) );
  XOR U4467 ( .A(in[1220]), .B(n3631), .Z(n3427) );
  NAND U4468 ( .A(n3430), .B(n3427), .Z(n2817) );
  XNOR U4469 ( .A(n3035), .B(n2817), .Z(out[360]) );
  XNOR U4470 ( .A(in[113]), .B(n3997), .Z(n3037) );
  XOR U4471 ( .A(in[1294]), .B(n3867), .Z(n3434) );
  XOR U4472 ( .A(in[1221]), .B(n3635), .Z(n3431) );
  NAND U4473 ( .A(n3434), .B(n3431), .Z(n2818) );
  XNOR U4474 ( .A(n3037), .B(n2818), .Z(out[361]) );
  XNOR U4475 ( .A(in[114]), .B(n4000), .Z(n3043) );
  XOR U4476 ( .A(in[1295]), .B(n3869), .Z(n3438) );
  XOR U4477 ( .A(in[1222]), .B(n3639), .Z(n3435) );
  NAND U4478 ( .A(n3438), .B(n3435), .Z(n2819) );
  XNOR U4479 ( .A(n3043), .B(n2819), .Z(out[362]) );
  XNOR U4480 ( .A(in[115]), .B(n4007), .Z(n3045) );
  XOR U4481 ( .A(in[1296]), .B(n3871), .Z(n3442) );
  XOR U4482 ( .A(in[1223]), .B(n3643), .Z(n3439) );
  NAND U4483 ( .A(n3442), .B(n3439), .Z(n2820) );
  XNOR U4484 ( .A(n3045), .B(n2820), .Z(out[363]) );
  XNOR U4485 ( .A(in[116]), .B(n4010), .Z(n3047) );
  XOR U4486 ( .A(in[1297]), .B(n3873), .Z(n3450) );
  XOR U4487 ( .A(in[1224]), .B(n3647), .Z(n3447) );
  NAND U4488 ( .A(n3450), .B(n3447), .Z(n2821) );
  XNOR U4489 ( .A(n3047), .B(n2821), .Z(out[364]) );
  XNOR U4490 ( .A(in[117]), .B(n4013), .Z(n3049) );
  XOR U4491 ( .A(in[1298]), .B(n3877), .Z(n3454) );
  XOR U4492 ( .A(in[1225]), .B(n3651), .Z(n3451) );
  NAND U4493 ( .A(n3454), .B(n3451), .Z(n2822) );
  XNOR U4494 ( .A(n3049), .B(n2822), .Z(out[365]) );
  XNOR U4495 ( .A(in[118]), .B(n4016), .Z(n3051) );
  XOR U4496 ( .A(in[1299]), .B(n3879), .Z(n3458) );
  XOR U4497 ( .A(in[1226]), .B(n3655), .Z(n3455) );
  NAND U4498 ( .A(n3458), .B(n3455), .Z(n2823) );
  XNOR U4499 ( .A(n3051), .B(n2823), .Z(out[366]) );
  XNOR U4500 ( .A(in[119]), .B(n4019), .Z(n3053) );
  XOR U4501 ( .A(in[1300]), .B(n3881), .Z(n3462) );
  XOR U4502 ( .A(in[1227]), .B(n3659), .Z(n3459) );
  NAND U4503 ( .A(n3462), .B(n3459), .Z(n2824) );
  XNOR U4504 ( .A(n3053), .B(n2824), .Z(out[367]) );
  XNOR U4505 ( .A(in[120]), .B(n4022), .Z(n3055) );
  XOR U4506 ( .A(in[1301]), .B(n3883), .Z(n3466) );
  XOR U4507 ( .A(in[1228]), .B(n3667), .Z(n3463) );
  NAND U4508 ( .A(n3466), .B(n3463), .Z(n2825) );
  XNOR U4509 ( .A(n3055), .B(n2825), .Z(out[368]) );
  XNOR U4510 ( .A(in[121]), .B(n4025), .Z(n3057) );
  XOR U4511 ( .A(in[1302]), .B(n3885), .Z(n3470) );
  XOR U4512 ( .A(in[1229]), .B(n3671), .Z(n3467) );
  NAND U4513 ( .A(n3470), .B(n3467), .Z(n2826) );
  XNOR U4514 ( .A(n3057), .B(n2826), .Z(out[369]) );
  ANDN U4515 ( .B(n2828), .A(n2827), .Z(n2829) );
  XNOR U4516 ( .A(n2830), .B(n2829), .Z(out[36]) );
  XNOR U4517 ( .A(in[122]), .B(n4028), .Z(n3059) );
  XOR U4518 ( .A(in[1303]), .B(n3887), .Z(n3474) );
  XOR U4519 ( .A(in[1230]), .B(n3675), .Z(n3471) );
  NAND U4520 ( .A(n3474), .B(n3471), .Z(n2831) );
  XNOR U4521 ( .A(n3059), .B(n2831), .Z(out[370]) );
  XNOR U4522 ( .A(in[123]), .B(n4031), .Z(n3061) );
  XOR U4523 ( .A(in[1304]), .B(n3889), .Z(n3478) );
  XOR U4524 ( .A(in[1231]), .B(n3679), .Z(n3475) );
  NAND U4525 ( .A(n3478), .B(n3475), .Z(n2832) );
  XNOR U4526 ( .A(n3061), .B(n2832), .Z(out[371]) );
  XNOR U4527 ( .A(in[124]), .B(n4034), .Z(n3069) );
  XOR U4528 ( .A(in[1305]), .B(n3891), .Z(n3482) );
  XOR U4529 ( .A(in[1232]), .B(n3683), .Z(n3479) );
  NAND U4530 ( .A(n3482), .B(n3479), .Z(n2833) );
  XNOR U4531 ( .A(n3069), .B(n2833), .Z(out[372]) );
  XNOR U4532 ( .A(in[125]), .B(n4041), .Z(n3071) );
  XOR U4533 ( .A(in[1306]), .B(n3893), .Z(n3486) );
  XOR U4534 ( .A(in[1233]), .B(n3687), .Z(n3483) );
  NAND U4535 ( .A(n3486), .B(n3483), .Z(n2834) );
  XNOR U4536 ( .A(n3071), .B(n2834), .Z(out[373]) );
  XNOR U4537 ( .A(in[126]), .B(n4044), .Z(n3073) );
  XOR U4538 ( .A(in[1307]), .B(n3895), .Z(n3494) );
  XOR U4539 ( .A(in[1234]), .B(n3691), .Z(n3491) );
  NAND U4540 ( .A(n3494), .B(n3491), .Z(n2835) );
  XNOR U4541 ( .A(n3073), .B(n2835), .Z(out[374]) );
  XNOR U4542 ( .A(in[127]), .B(n4047), .Z(n3075) );
  XOR U4543 ( .A(in[1308]), .B(n3899), .Z(n3498) );
  XOR U4544 ( .A(in[1235]), .B(n3695), .Z(n3495) );
  NAND U4545 ( .A(n3498), .B(n3495), .Z(n2836) );
  XNOR U4546 ( .A(n3075), .B(n2836), .Z(out[375]) );
  XNOR U4547 ( .A(in[64]), .B(n4050), .Z(n3077) );
  XOR U4548 ( .A(in[1309]), .B(n3901), .Z(n3502) );
  XOR U4549 ( .A(in[1236]), .B(n3699), .Z(n3499) );
  NAND U4550 ( .A(n3502), .B(n3499), .Z(n2837) );
  XNOR U4551 ( .A(n3077), .B(n2837), .Z(out[376]) );
  XNOR U4552 ( .A(in[65]), .B(n4053), .Z(n3079) );
  XOR U4553 ( .A(in[1310]), .B(n3903), .Z(n3506) );
  XOR U4554 ( .A(in[1237]), .B(n3703), .Z(n3503) );
  NAND U4555 ( .A(n3506), .B(n3503), .Z(n2838) );
  XNOR U4556 ( .A(n3079), .B(n2838), .Z(out[377]) );
  XNOR U4557 ( .A(in[66]), .B(n4056), .Z(n3081) );
  XOR U4558 ( .A(in[1311]), .B(n3905), .Z(n3510) );
  XOR U4559 ( .A(in[1238]), .B(n3711), .Z(n3507) );
  NAND U4560 ( .A(n3510), .B(n3507), .Z(n2839) );
  XNOR U4561 ( .A(n3081), .B(n2839), .Z(out[378]) );
  XNOR U4562 ( .A(in[67]), .B(n4059), .Z(n3083) );
  XOR U4563 ( .A(in[1312]), .B(n3907), .Z(n3514) );
  XOR U4564 ( .A(in[1239]), .B(n3715), .Z(n3511) );
  NAND U4565 ( .A(n3514), .B(n3511), .Z(n2840) );
  XNOR U4566 ( .A(n3083), .B(n2840), .Z(out[379]) );
  ANDN U4567 ( .B(n2842), .A(n2841), .Z(n2843) );
  XNOR U4568 ( .A(n2844), .B(n2843), .Z(out[37]) );
  XNOR U4569 ( .A(in[68]), .B(n4062), .Z(n3085) );
  XOR U4570 ( .A(in[1313]), .B(n3909), .Z(n3518) );
  XOR U4571 ( .A(in[1240]), .B(n3719), .Z(n3515) );
  NAND U4572 ( .A(n3518), .B(n3515), .Z(n2845) );
  XNOR U4573 ( .A(n3085), .B(n2845), .Z(out[380]) );
  XNOR U4574 ( .A(in[69]), .B(n4065), .Z(n3087) );
  XOR U4575 ( .A(in[1314]), .B(n3911), .Z(n3522) );
  XOR U4576 ( .A(in[1241]), .B(n3723), .Z(n3519) );
  NAND U4577 ( .A(n3522), .B(n3519), .Z(n2846) );
  XNOR U4578 ( .A(n3087), .B(n2846), .Z(out[381]) );
  XNOR U4579 ( .A(in[70]), .B(n4068), .Z(n3093) );
  XOR U4580 ( .A(in[1315]), .B(n3913), .Z(n3526) );
  XOR U4581 ( .A(in[1242]), .B(n3727), .Z(n3523) );
  NAND U4582 ( .A(n3526), .B(n3523), .Z(n2847) );
  XNOR U4583 ( .A(n3093), .B(n2847), .Z(out[382]) );
  XNOR U4584 ( .A(in[71]), .B(n4079), .Z(n3095) );
  XOR U4585 ( .A(in[1316]), .B(n3915), .Z(n3530) );
  XOR U4586 ( .A(in[1243]), .B(n3731), .Z(n3527) );
  NAND U4587 ( .A(n3530), .B(n3527), .Z(n2848) );
  XNOR U4588 ( .A(n3095), .B(n2848), .Z(out[383]) );
  XOR U4589 ( .A(in[497]), .B(n3777), .Z(n3097) );
  NOR U4590 ( .A(n2939), .B(n3252), .Z(n2849) );
  XNOR U4591 ( .A(n3097), .B(n2849), .Z(out[384]) );
  XOR U4592 ( .A(in[498]), .B(n3781), .Z(n3099) );
  NOR U4593 ( .A(n2941), .B(n3256), .Z(n2850) );
  XNOR U4594 ( .A(n3099), .B(n2850), .Z(out[385]) );
  XOR U4595 ( .A(in[499]), .B(n3785), .Z(n3101) );
  NOR U4596 ( .A(n2947), .B(n3260), .Z(n2851) );
  XNOR U4597 ( .A(n3101), .B(n2851), .Z(out[386]) );
  XOR U4598 ( .A(in[500]), .B(n3789), .Z(n3103) );
  NOR U4599 ( .A(n2949), .B(n3264), .Z(n2852) );
  XNOR U4600 ( .A(n3103), .B(n2852), .Z(out[387]) );
  XOR U4601 ( .A(in[501]), .B(n3793), .Z(n3105) );
  NOR U4602 ( .A(n2951), .B(n3272), .Z(n2853) );
  XNOR U4603 ( .A(n3105), .B(n2853), .Z(out[388]) );
  XOR U4604 ( .A(in[502]), .B(n3803), .Z(n3107) );
  NOR U4605 ( .A(n2953), .B(n3276), .Z(n2854) );
  XNOR U4606 ( .A(n3107), .B(n2854), .Z(out[389]) );
  ANDN U4607 ( .B(n2856), .A(n2855), .Z(n2857) );
  XNOR U4608 ( .A(n2858), .B(n2857), .Z(out[38]) );
  XOR U4609 ( .A(in[503]), .B(n3807), .Z(n3109) );
  NOR U4610 ( .A(n2955), .B(n3280), .Z(n2859) );
  XNOR U4611 ( .A(n3109), .B(n2859), .Z(out[390]) );
  XOR U4612 ( .A(in[504]), .B(n3811), .Z(n3111) );
  NOR U4613 ( .A(n2957), .B(n3284), .Z(n2860) );
  XNOR U4614 ( .A(n3111), .B(n2860), .Z(out[391]) );
  XOR U4615 ( .A(in[505]), .B(n3815), .Z(n3117) );
  NOR U4616 ( .A(n2959), .B(n3288), .Z(n2861) );
  XNOR U4617 ( .A(n3117), .B(n2861), .Z(out[392]) );
  XOR U4618 ( .A(in[506]), .B(n3537), .Z(n3119) );
  NOR U4619 ( .A(n2961), .B(n3292), .Z(n2862) );
  XNOR U4620 ( .A(n3119), .B(n2862), .Z(out[393]) );
  XOR U4621 ( .A(in[507]), .B(n3541), .Z(n3121) );
  NOR U4622 ( .A(n2963), .B(n3296), .Z(n2863) );
  XNOR U4623 ( .A(n3121), .B(n2863), .Z(out[394]) );
  XOR U4624 ( .A(in[508]), .B(n3545), .Z(n3123) );
  NOR U4625 ( .A(n2965), .B(n3300), .Z(n2864) );
  XNOR U4626 ( .A(n3123), .B(n2864), .Z(out[395]) );
  XOR U4627 ( .A(in[509]), .B(n3549), .Z(n3125) );
  NOR U4628 ( .A(n2971), .B(n3304), .Z(n2865) );
  XNOR U4629 ( .A(n3125), .B(n2865), .Z(out[396]) );
  XOR U4630 ( .A(in[510]), .B(n3553), .Z(n3127) );
  NOR U4631 ( .A(n2973), .B(n3308), .Z(n2866) );
  XNOR U4632 ( .A(n3127), .B(n2866), .Z(out[397]) );
  XOR U4633 ( .A(in[511]), .B(n3557), .Z(n3129) );
  NOR U4634 ( .A(n2975), .B(n3316), .Z(n2867) );
  XNOR U4635 ( .A(n3129), .B(n2867), .Z(out[398]) );
  XOR U4636 ( .A(in[448]), .B(n3561), .Z(n3131) );
  NOR U4637 ( .A(n2977), .B(n3320), .Z(n2868) );
  XNOR U4638 ( .A(n3131), .B(n2868), .Z(out[399]) );
  ANDN U4639 ( .B(n2870), .A(n2869), .Z(n2871) );
  XNOR U4640 ( .A(n2872), .B(n2871), .Z(out[39]) );
  OR U4641 ( .A(n3708), .B(n2873), .Z(n2874) );
  XNOR U4642 ( .A(n3707), .B(n2874), .Z(out[3]) );
  XOR U4643 ( .A(in[449]), .B(n3565), .Z(n3133) );
  NOR U4644 ( .A(n2979), .B(n3324), .Z(n2875) );
  XNOR U4645 ( .A(n3133), .B(n2875), .Z(out[400]) );
  XNOR U4646 ( .A(n3569), .B(in[450]), .Z(n3135) );
  NOR U4647 ( .A(n2981), .B(n3328), .Z(n2876) );
  XNOR U4648 ( .A(n3135), .B(n2876), .Z(out[401]) );
  XNOR U4649 ( .A(n3573), .B(in[451]), .Z(n3141) );
  NOR U4650 ( .A(n2983), .B(n3332), .Z(n2877) );
  XNOR U4651 ( .A(n3141), .B(n2877), .Z(out[402]) );
  XNOR U4652 ( .A(n3581), .B(in[452]), .Z(n3143) );
  NOR U4653 ( .A(n2985), .B(n3336), .Z(n2878) );
  XNOR U4654 ( .A(n3143), .B(n2878), .Z(out[403]) );
  XNOR U4655 ( .A(n3585), .B(in[453]), .Z(n3145) );
  NOR U4656 ( .A(n2987), .B(n3340), .Z(n2879) );
  XNOR U4657 ( .A(n3145), .B(n2879), .Z(out[404]) );
  XNOR U4658 ( .A(n3589), .B(in[454]), .Z(n3147) );
  NOR U4659 ( .A(n2989), .B(n3344), .Z(n2880) );
  XNOR U4660 ( .A(n3147), .B(n2880), .Z(out[405]) );
  XNOR U4661 ( .A(n3593), .B(in[455]), .Z(n3149) );
  NOR U4662 ( .A(n2995), .B(n3348), .Z(n2881) );
  XNOR U4663 ( .A(n3149), .B(n2881), .Z(out[406]) );
  XNOR U4664 ( .A(n3597), .B(in[456]), .Z(n3151) );
  NOR U4665 ( .A(n2997), .B(n3352), .Z(n2882) );
  XNOR U4666 ( .A(n3151), .B(n2882), .Z(out[407]) );
  XNOR U4667 ( .A(in[457]), .B(n3601), .Z(n3153) );
  NOR U4668 ( .A(n2999), .B(n3362), .Z(n2883) );
  XNOR U4669 ( .A(n3153), .B(n2883), .Z(out[408]) );
  XNOR U4670 ( .A(n3605), .B(in[458]), .Z(n3155) );
  NOR U4671 ( .A(n3001), .B(n3366), .Z(n2884) );
  XNOR U4672 ( .A(n3155), .B(n2884), .Z(out[409]) );
  ANDN U4673 ( .B(n2886), .A(n2885), .Z(n2887) );
  XNOR U4674 ( .A(n2888), .B(n2887), .Z(out[40]) );
  XNOR U4675 ( .A(n3609), .B(in[459]), .Z(n3157) );
  NOR U4676 ( .A(n3003), .B(n3370), .Z(n2889) );
  XNOR U4677 ( .A(n3157), .B(n2889), .Z(out[410]) );
  XNOR U4678 ( .A(in[460]), .B(n3613), .Z(n3159) );
  NOR U4679 ( .A(n3005), .B(n3374), .Z(n2890) );
  XNOR U4680 ( .A(n3159), .B(n2890), .Z(out[411]) );
  XNOR U4681 ( .A(in[461]), .B(n3617), .Z(n3165) );
  NOR U4682 ( .A(n3007), .B(n3378), .Z(n2891) );
  XNOR U4683 ( .A(n3165), .B(n2891), .Z(out[412]) );
  XNOR U4684 ( .A(in[462]), .B(n3625), .Z(n3167) );
  NOR U4685 ( .A(n3009), .B(n3382), .Z(n2892) );
  XNOR U4686 ( .A(n3167), .B(n2892), .Z(out[413]) );
  XNOR U4687 ( .A(in[463]), .B(n3629), .Z(n3169) );
  NOR U4688 ( .A(n3011), .B(n3386), .Z(n2893) );
  XNOR U4689 ( .A(n3169), .B(n2893), .Z(out[414]) );
  XNOR U4690 ( .A(in[464]), .B(n3633), .Z(n3171) );
  NOR U4691 ( .A(n3013), .B(n3390), .Z(n2894) );
  XNOR U4692 ( .A(n3171), .B(n2894), .Z(out[415]) );
  XNOR U4693 ( .A(in[465]), .B(n3637), .Z(n3173) );
  NOR U4694 ( .A(n3019), .B(n3394), .Z(n2895) );
  XNOR U4695 ( .A(n3173), .B(n2895), .Z(out[416]) );
  XNOR U4696 ( .A(in[466]), .B(n3641), .Z(n3175) );
  NOR U4697 ( .A(n3021), .B(n3398), .Z(n2896) );
  XNOR U4698 ( .A(n3175), .B(n2896), .Z(out[417]) );
  XNOR U4699 ( .A(in[467]), .B(n3645), .Z(n3177) );
  NOR U4700 ( .A(n3023), .B(n3406), .Z(n2897) );
  XNOR U4701 ( .A(n3177), .B(n2897), .Z(out[418]) );
  XNOR U4702 ( .A(in[468]), .B(n3649), .Z(n3179) );
  NOR U4703 ( .A(n3025), .B(n3410), .Z(n2898) );
  XNOR U4704 ( .A(n3179), .B(n2898), .Z(out[419]) );
  ANDN U4705 ( .B(n2900), .A(n2899), .Z(n2901) );
  XNOR U4706 ( .A(n2902), .B(n2901), .Z(out[41]) );
  XNOR U4707 ( .A(in[469]), .B(n3653), .Z(n3181) );
  NOR U4708 ( .A(n3027), .B(n3414), .Z(n2903) );
  XNOR U4709 ( .A(n3181), .B(n2903), .Z(out[420]) );
  XNOR U4710 ( .A(in[470]), .B(n3657), .Z(n3183) );
  NOR U4711 ( .A(n3029), .B(n3418), .Z(n2904) );
  XNOR U4712 ( .A(n3183), .B(n2904), .Z(out[421]) );
  XNOR U4713 ( .A(in[471]), .B(n3661), .Z(n3189) );
  NOR U4714 ( .A(n3031), .B(n3422), .Z(n2905) );
  XNOR U4715 ( .A(n3189), .B(n2905), .Z(out[422]) );
  XNOR U4716 ( .A(in[472]), .B(n3669), .Z(n3191) );
  NOR U4717 ( .A(n3033), .B(n3426), .Z(n2906) );
  XNOR U4718 ( .A(n3191), .B(n2906), .Z(out[423]) );
  XNOR U4719 ( .A(in[473]), .B(n3673), .Z(n3193) );
  NOR U4720 ( .A(n3035), .B(n3430), .Z(n2907) );
  XNOR U4721 ( .A(n3193), .B(n2907), .Z(out[424]) );
  XNOR U4722 ( .A(in[474]), .B(n3677), .Z(n3195) );
  NOR U4723 ( .A(n3037), .B(n3434), .Z(n2908) );
  XNOR U4724 ( .A(n3195), .B(n2908), .Z(out[425]) );
  XNOR U4725 ( .A(in[475]), .B(n3681), .Z(n3197) );
  NOR U4726 ( .A(n3043), .B(n3438), .Z(n2909) );
  XNOR U4727 ( .A(n3197), .B(n2909), .Z(out[426]) );
  XNOR U4728 ( .A(in[476]), .B(n3685), .Z(n3199) );
  NOR U4729 ( .A(n3045), .B(n3442), .Z(n2910) );
  XNOR U4730 ( .A(n3199), .B(n2910), .Z(out[427]) );
  XNOR U4731 ( .A(in[477]), .B(n3689), .Z(n3201) );
  NOR U4732 ( .A(n3047), .B(n3450), .Z(n2911) );
  XNOR U4733 ( .A(n3201), .B(n2911), .Z(out[428]) );
  XNOR U4734 ( .A(in[478]), .B(n3693), .Z(n3203) );
  NOR U4735 ( .A(n3049), .B(n3454), .Z(n2912) );
  XNOR U4736 ( .A(n3203), .B(n2912), .Z(out[429]) );
  ANDN U4737 ( .B(n2914), .A(n2913), .Z(n2915) );
  XNOR U4738 ( .A(n2916), .B(n2915), .Z(out[42]) );
  XNOR U4739 ( .A(in[479]), .B(n3697), .Z(n3205) );
  NOR U4740 ( .A(n3051), .B(n3458), .Z(n2917) );
  XNOR U4741 ( .A(n3205), .B(n2917), .Z(out[430]) );
  XNOR U4742 ( .A(in[480]), .B(n3701), .Z(n3207) );
  NOR U4743 ( .A(n3053), .B(n3462), .Z(n2918) );
  XNOR U4744 ( .A(n3207), .B(n2918), .Z(out[431]) );
  XNOR U4745 ( .A(in[481]), .B(n3705), .Z(n3213) );
  NOR U4746 ( .A(n3055), .B(n3466), .Z(n2919) );
  XNOR U4747 ( .A(n3213), .B(n2919), .Z(out[432]) );
  XNOR U4748 ( .A(in[482]), .B(n3713), .Z(n3215) );
  NOR U4749 ( .A(n3057), .B(n3470), .Z(n2920) );
  XNOR U4750 ( .A(n3215), .B(n2920), .Z(out[433]) );
  XNOR U4751 ( .A(in[483]), .B(n3717), .Z(n3217) );
  NOR U4752 ( .A(n3059), .B(n3474), .Z(n2921) );
  XNOR U4753 ( .A(n3217), .B(n2921), .Z(out[434]) );
  XNOR U4754 ( .A(in[484]), .B(n3721), .Z(n3219) );
  NOR U4755 ( .A(n3061), .B(n3478), .Z(n2922) );
  XNOR U4756 ( .A(n3219), .B(n2922), .Z(out[435]) );
  XNOR U4757 ( .A(in[485]), .B(n3725), .Z(n3221) );
  NOR U4758 ( .A(n3069), .B(n3482), .Z(n2923) );
  XNOR U4759 ( .A(n3221), .B(n2923), .Z(out[436]) );
  XOR U4760 ( .A(in[486]), .B(n3729), .Z(n3223) );
  NOR U4761 ( .A(n3071), .B(n3486), .Z(n2924) );
  XNOR U4762 ( .A(n3223), .B(n2924), .Z(out[437]) );
  XOR U4763 ( .A(in[487]), .B(n3733), .Z(n3225) );
  NOR U4764 ( .A(n3073), .B(n3494), .Z(n2925) );
  XNOR U4765 ( .A(n3225), .B(n2925), .Z(out[438]) );
  XOR U4766 ( .A(in[488]), .B(n3737), .Z(n3227) );
  NOR U4767 ( .A(n3075), .B(n3498), .Z(n2926) );
  XNOR U4768 ( .A(n3227), .B(n2926), .Z(out[439]) );
  ANDN U4769 ( .B(n2928), .A(n2927), .Z(n2929) );
  XNOR U4770 ( .A(n2930), .B(n2929), .Z(out[43]) );
  XOR U4771 ( .A(in[489]), .B(n3741), .Z(n3229) );
  NOR U4772 ( .A(n3077), .B(n3502), .Z(n2931) );
  XNOR U4773 ( .A(n3229), .B(n2931), .Z(out[440]) );
  XOR U4774 ( .A(in[490]), .B(n3745), .Z(n3231) );
  NOR U4775 ( .A(n3079), .B(n3506), .Z(n2932) );
  XNOR U4776 ( .A(n3231), .B(n2932), .Z(out[441]) );
  XOR U4777 ( .A(in[491]), .B(n3749), .Z(n3237) );
  NOR U4778 ( .A(n3081), .B(n3510), .Z(n2933) );
  XNOR U4779 ( .A(n3237), .B(n2933), .Z(out[442]) );
  XOR U4780 ( .A(in[492]), .B(n3757), .Z(n3239) );
  NOR U4781 ( .A(n3083), .B(n3514), .Z(n2934) );
  XNOR U4782 ( .A(n3239), .B(n2934), .Z(out[443]) );
  XOR U4783 ( .A(in[493]), .B(n3761), .Z(n3241) );
  NOR U4784 ( .A(n3085), .B(n3518), .Z(n2935) );
  XNOR U4785 ( .A(n3241), .B(n2935), .Z(out[444]) );
  XOR U4786 ( .A(in[494]), .B(n3765), .Z(n3243) );
  NOR U4787 ( .A(n3087), .B(n3522), .Z(n2936) );
  XNOR U4788 ( .A(n3243), .B(n2936), .Z(out[445]) );
  XOR U4789 ( .A(in[495]), .B(n3769), .Z(n3245) );
  NOR U4790 ( .A(n3093), .B(n3526), .Z(n2937) );
  XNOR U4791 ( .A(n3245), .B(n2937), .Z(out[446]) );
  XOR U4792 ( .A(in[496]), .B(n3773), .Z(n3247) );
  NOR U4793 ( .A(n3095), .B(n3530), .Z(n2938) );
  XNOR U4794 ( .A(n3247), .B(n2938), .Z(out[447]) );
  XNOR U4795 ( .A(in[886]), .B(n3776), .Z(n3250) );
  NAND U4796 ( .A(n3097), .B(n2939), .Z(n2940) );
  XNOR U4797 ( .A(n3250), .B(n2940), .Z(out[448]) );
  XNOR U4798 ( .A(in[887]), .B(n3780), .Z(n3254) );
  NAND U4799 ( .A(n3099), .B(n2941), .Z(n2942) );
  XNOR U4800 ( .A(n3254), .B(n2942), .Z(out[449]) );
  ANDN U4801 ( .B(n2944), .A(n2943), .Z(n2945) );
  XNOR U4802 ( .A(n2946), .B(n2945), .Z(out[44]) );
  XNOR U4803 ( .A(in[888]), .B(n3784), .Z(n3258) );
  NAND U4804 ( .A(n3101), .B(n2947), .Z(n2948) );
  XNOR U4805 ( .A(n3258), .B(n2948), .Z(out[450]) );
  XNOR U4806 ( .A(in[889]), .B(n3788), .Z(n3262) );
  NAND U4807 ( .A(n3103), .B(n2949), .Z(n2950) );
  XNOR U4808 ( .A(n3262), .B(n2950), .Z(out[451]) );
  XNOR U4809 ( .A(in[890]), .B(n3792), .Z(n3270) );
  NAND U4810 ( .A(n3105), .B(n2951), .Z(n2952) );
  XNOR U4811 ( .A(n3270), .B(n2952), .Z(out[452]) );
  XOR U4812 ( .A(in[891]), .B(n3802), .Z(n3274) );
  NAND U4813 ( .A(n3107), .B(n2953), .Z(n2954) );
  XNOR U4814 ( .A(n3274), .B(n2954), .Z(out[453]) );
  XOR U4815 ( .A(in[892]), .B(n3806), .Z(n3278) );
  NAND U4816 ( .A(n3109), .B(n2955), .Z(n2956) );
  XNOR U4817 ( .A(n3278), .B(n2956), .Z(out[454]) );
  XOR U4818 ( .A(in[893]), .B(n3810), .Z(n3282) );
  NAND U4819 ( .A(n3111), .B(n2957), .Z(n2958) );
  XNOR U4820 ( .A(n3282), .B(n2958), .Z(out[455]) );
  XNOR U4821 ( .A(in[894]), .B(n3814), .Z(n3286) );
  NAND U4822 ( .A(n3117), .B(n2959), .Z(n2960) );
  XNOR U4823 ( .A(n3286), .B(n2960), .Z(out[456]) );
  XOR U4824 ( .A(in[895]), .B(n3536), .Z(n3290) );
  NAND U4825 ( .A(n3119), .B(n2961), .Z(n2962) );
  XNOR U4826 ( .A(n3290), .B(n2962), .Z(out[457]) );
  XOR U4827 ( .A(in[832]), .B(n3540), .Z(n3294) );
  NAND U4828 ( .A(n3121), .B(n2963), .Z(n2964) );
  XNOR U4829 ( .A(n3294), .B(n2964), .Z(out[458]) );
  XOR U4830 ( .A(in[833]), .B(n3544), .Z(n3298) );
  NAND U4831 ( .A(n3123), .B(n2965), .Z(n2966) );
  XNOR U4832 ( .A(n3298), .B(n2966), .Z(out[459]) );
  ANDN U4833 ( .B(n2968), .A(n2967), .Z(n2969) );
  XNOR U4834 ( .A(n2970), .B(n2969), .Z(out[45]) );
  XOR U4835 ( .A(in[834]), .B(n3548), .Z(n3302) );
  NAND U4836 ( .A(n3125), .B(n2971), .Z(n2972) );
  XNOR U4837 ( .A(n3302), .B(n2972), .Z(out[460]) );
  XOR U4838 ( .A(in[835]), .B(n3552), .Z(n3306) );
  NAND U4839 ( .A(n3127), .B(n2973), .Z(n2974) );
  XNOR U4840 ( .A(n3306), .B(n2974), .Z(out[461]) );
  XOR U4841 ( .A(in[836]), .B(n3556), .Z(n3314) );
  NAND U4842 ( .A(n3129), .B(n2975), .Z(n2976) );
  XNOR U4843 ( .A(n3314), .B(n2976), .Z(out[462]) );
  XOR U4844 ( .A(in[837]), .B(n3560), .Z(n3318) );
  NAND U4845 ( .A(n3131), .B(n2977), .Z(n2978) );
  XNOR U4846 ( .A(n3318), .B(n2978), .Z(out[463]) );
  XOR U4847 ( .A(in[838]), .B(n3564), .Z(n3322) );
  NAND U4848 ( .A(n3133), .B(n2979), .Z(n2980) );
  XNOR U4849 ( .A(n3322), .B(n2980), .Z(out[464]) );
  XOR U4850 ( .A(in[839]), .B(n3568), .Z(n3326) );
  NAND U4851 ( .A(n3135), .B(n2981), .Z(n2982) );
  XNOR U4852 ( .A(n3326), .B(n2982), .Z(out[465]) );
  XOR U4853 ( .A(in[840]), .B(n3572), .Z(n3330) );
  NAND U4854 ( .A(n3141), .B(n2983), .Z(n2984) );
  XNOR U4855 ( .A(n3330), .B(n2984), .Z(out[466]) );
  XOR U4856 ( .A(in[841]), .B(n3580), .Z(n3334) );
  NAND U4857 ( .A(n3143), .B(n2985), .Z(n2986) );
  XNOR U4858 ( .A(n3334), .B(n2986), .Z(out[467]) );
  XOR U4859 ( .A(in[842]), .B(n3584), .Z(n3338) );
  NAND U4860 ( .A(n3145), .B(n2987), .Z(n2988) );
  XNOR U4861 ( .A(n3338), .B(n2988), .Z(out[468]) );
  XOR U4862 ( .A(in[843]), .B(n3588), .Z(n3342) );
  NAND U4863 ( .A(n3147), .B(n2989), .Z(n2990) );
  XNOR U4864 ( .A(n3342), .B(n2990), .Z(out[469]) );
  ANDN U4865 ( .B(n2992), .A(n2991), .Z(n2993) );
  XNOR U4866 ( .A(n2994), .B(n2993), .Z(out[46]) );
  XOR U4867 ( .A(in[844]), .B(n3592), .Z(n3346) );
  NAND U4868 ( .A(n3149), .B(n2995), .Z(n2996) );
  XNOR U4869 ( .A(n3346), .B(n2996), .Z(out[470]) );
  XOR U4870 ( .A(in[845]), .B(n3596), .Z(n3350) );
  NAND U4871 ( .A(n3151), .B(n2997), .Z(n2998) );
  XNOR U4872 ( .A(n3350), .B(n2998), .Z(out[471]) );
  XOR U4873 ( .A(in[846]), .B(n3600), .Z(n3360) );
  NAND U4874 ( .A(n3153), .B(n2999), .Z(n3000) );
  XNOR U4875 ( .A(n3360), .B(n3000), .Z(out[472]) );
  XOR U4876 ( .A(in[847]), .B(n3604), .Z(n3364) );
  NAND U4877 ( .A(n3155), .B(n3001), .Z(n3002) );
  XNOR U4878 ( .A(n3364), .B(n3002), .Z(out[473]) );
  XOR U4879 ( .A(in[848]), .B(n3608), .Z(n3368) );
  NAND U4880 ( .A(n3157), .B(n3003), .Z(n3004) );
  XNOR U4881 ( .A(n3368), .B(n3004), .Z(out[474]) );
  XOR U4882 ( .A(in[849]), .B(n3612), .Z(n3372) );
  NAND U4883 ( .A(n3159), .B(n3005), .Z(n3006) );
  XNOR U4884 ( .A(n3372), .B(n3006), .Z(out[475]) );
  XOR U4885 ( .A(in[850]), .B(n3616), .Z(n3376) );
  NAND U4886 ( .A(n3165), .B(n3007), .Z(n3008) );
  XNOR U4887 ( .A(n3376), .B(n3008), .Z(out[476]) );
  XNOR U4888 ( .A(in[851]), .B(n3624), .Z(n3380) );
  NAND U4889 ( .A(n3167), .B(n3009), .Z(n3010) );
  XNOR U4890 ( .A(n3380), .B(n3010), .Z(out[477]) );
  XNOR U4891 ( .A(in[852]), .B(n3628), .Z(n3384) );
  NAND U4892 ( .A(n3169), .B(n3011), .Z(n3012) );
  XNOR U4893 ( .A(n3384), .B(n3012), .Z(out[478]) );
  XNOR U4894 ( .A(in[853]), .B(n3632), .Z(n3388) );
  NAND U4895 ( .A(n3171), .B(n3013), .Z(n3014) );
  XNOR U4896 ( .A(n3388), .B(n3014), .Z(out[479]) );
  ANDN U4897 ( .B(n3016), .A(n3015), .Z(n3017) );
  XNOR U4898 ( .A(n3018), .B(n3017), .Z(out[47]) );
  XNOR U4899 ( .A(in[854]), .B(n3636), .Z(n3392) );
  NAND U4900 ( .A(n3173), .B(n3019), .Z(n3020) );
  XNOR U4901 ( .A(n3392), .B(n3020), .Z(out[480]) );
  XNOR U4902 ( .A(in[855]), .B(n3640), .Z(n3396) );
  NAND U4903 ( .A(n3175), .B(n3021), .Z(n3022) );
  XNOR U4904 ( .A(n3396), .B(n3022), .Z(out[481]) );
  XNOR U4905 ( .A(in[856]), .B(n3644), .Z(n3404) );
  NAND U4906 ( .A(n3177), .B(n3023), .Z(n3024) );
  XNOR U4907 ( .A(n3404), .B(n3024), .Z(out[482]) );
  XNOR U4908 ( .A(in[857]), .B(n3648), .Z(n3408) );
  NAND U4909 ( .A(n3179), .B(n3025), .Z(n3026) );
  XNOR U4910 ( .A(n3408), .B(n3026), .Z(out[483]) );
  XNOR U4911 ( .A(in[858]), .B(n3652), .Z(n3412) );
  NAND U4912 ( .A(n3181), .B(n3027), .Z(n3028) );
  XNOR U4913 ( .A(n3412), .B(n3028), .Z(out[484]) );
  XNOR U4914 ( .A(in[859]), .B(n3656), .Z(n3416) );
  NAND U4915 ( .A(n3183), .B(n3029), .Z(n3030) );
  XNOR U4916 ( .A(n3416), .B(n3030), .Z(out[485]) );
  XNOR U4917 ( .A(in[860]), .B(n3660), .Z(n3420) );
  NAND U4918 ( .A(n3189), .B(n3031), .Z(n3032) );
  XNOR U4919 ( .A(n3420), .B(n3032), .Z(out[486]) );
  XNOR U4920 ( .A(in[861]), .B(n3668), .Z(n3424) );
  NAND U4921 ( .A(n3191), .B(n3033), .Z(n3034) );
  XNOR U4922 ( .A(n3424), .B(n3034), .Z(out[487]) );
  XNOR U4923 ( .A(in[862]), .B(n3672), .Z(n3428) );
  NAND U4924 ( .A(n3193), .B(n3035), .Z(n3036) );
  XNOR U4925 ( .A(n3428), .B(n3036), .Z(out[488]) );
  XNOR U4926 ( .A(in[863]), .B(n3676), .Z(n3432) );
  NAND U4927 ( .A(n3195), .B(n3037), .Z(n3038) );
  XNOR U4928 ( .A(n3432), .B(n3038), .Z(out[489]) );
  ANDN U4929 ( .B(n3040), .A(n3039), .Z(n3041) );
  XNOR U4930 ( .A(n3042), .B(n3041), .Z(out[48]) );
  XNOR U4931 ( .A(in[864]), .B(n3680), .Z(n3436) );
  NAND U4932 ( .A(n3197), .B(n3043), .Z(n3044) );
  XNOR U4933 ( .A(n3436), .B(n3044), .Z(out[490]) );
  XNOR U4934 ( .A(in[865]), .B(n3684), .Z(n3440) );
  NAND U4935 ( .A(n3199), .B(n3045), .Z(n3046) );
  XNOR U4936 ( .A(n3440), .B(n3046), .Z(out[491]) );
  XOR U4937 ( .A(n3688), .B(in[866]), .Z(n3448) );
  NAND U4938 ( .A(n3201), .B(n3047), .Z(n3048) );
  XNOR U4939 ( .A(n3448), .B(n3048), .Z(out[492]) );
  XOR U4940 ( .A(n3692), .B(in[867]), .Z(n3452) );
  NAND U4941 ( .A(n3203), .B(n3049), .Z(n3050) );
  XNOR U4942 ( .A(n3452), .B(n3050), .Z(out[493]) );
  XOR U4943 ( .A(n3696), .B(in[868]), .Z(n3456) );
  NAND U4944 ( .A(n3205), .B(n3051), .Z(n3052) );
  XNOR U4945 ( .A(n3456), .B(n3052), .Z(out[494]) );
  XOR U4946 ( .A(n3700), .B(in[869]), .Z(n3460) );
  NAND U4947 ( .A(n3207), .B(n3053), .Z(n3054) );
  XNOR U4948 ( .A(n3460), .B(n3054), .Z(out[495]) );
  XNOR U4949 ( .A(in[870]), .B(n3704), .Z(n3464) );
  NAND U4950 ( .A(n3213), .B(n3055), .Z(n3056) );
  XNOR U4951 ( .A(n3464), .B(n3056), .Z(out[496]) );
  XNOR U4952 ( .A(in[871]), .B(n3712), .Z(n3468) );
  NAND U4953 ( .A(n3215), .B(n3057), .Z(n3058) );
  XNOR U4954 ( .A(n3468), .B(n3058), .Z(out[497]) );
  XNOR U4955 ( .A(in[872]), .B(n3716), .Z(n3472) );
  NAND U4956 ( .A(n3217), .B(n3059), .Z(n3060) );
  XNOR U4957 ( .A(n3472), .B(n3060), .Z(out[498]) );
  XNOR U4958 ( .A(in[873]), .B(n3720), .Z(n3476) );
  NAND U4959 ( .A(n3219), .B(n3061), .Z(n3062) );
  XNOR U4960 ( .A(n3476), .B(n3062), .Z(out[499]) );
  ANDN U4961 ( .B(n3064), .A(n3063), .Z(n3065) );
  XNOR U4962 ( .A(n3066), .B(n3065), .Z(out[49]) );
  OR U4963 ( .A(n3752), .B(n3067), .Z(n3068) );
  XNOR U4964 ( .A(n3751), .B(n3068), .Z(out[4]) );
  XNOR U4965 ( .A(in[874]), .B(n3724), .Z(n3480) );
  NAND U4966 ( .A(n3221), .B(n3069), .Z(n3070) );
  XNOR U4967 ( .A(n3480), .B(n3070), .Z(out[500]) );
  XNOR U4968 ( .A(in[875]), .B(n3728), .Z(n3484) );
  NAND U4969 ( .A(n3223), .B(n3071), .Z(n3072) );
  XNOR U4970 ( .A(n3484), .B(n3072), .Z(out[501]) );
  XNOR U4971 ( .A(in[876]), .B(n3732), .Z(n3492) );
  NAND U4972 ( .A(n3225), .B(n3073), .Z(n3074) );
  XNOR U4973 ( .A(n3492), .B(n3074), .Z(out[502]) );
  XNOR U4974 ( .A(in[877]), .B(n3736), .Z(n3496) );
  NAND U4975 ( .A(n3227), .B(n3075), .Z(n3076) );
  XNOR U4976 ( .A(n3496), .B(n3076), .Z(out[503]) );
  XNOR U4977 ( .A(in[878]), .B(n3740), .Z(n3500) );
  NAND U4978 ( .A(n3229), .B(n3077), .Z(n3078) );
  XNOR U4979 ( .A(n3500), .B(n3078), .Z(out[504]) );
  XNOR U4980 ( .A(in[879]), .B(n3744), .Z(n3504) );
  NAND U4981 ( .A(n3231), .B(n3079), .Z(n3080) );
  XNOR U4982 ( .A(n3504), .B(n3080), .Z(out[505]) );
  XNOR U4983 ( .A(in[880]), .B(n3748), .Z(n3508) );
  NAND U4984 ( .A(n3237), .B(n3081), .Z(n3082) );
  XNOR U4985 ( .A(n3508), .B(n3082), .Z(out[506]) );
  XNOR U4986 ( .A(in[881]), .B(n3756), .Z(n3512) );
  NAND U4987 ( .A(n3239), .B(n3083), .Z(n3084) );
  XNOR U4988 ( .A(n3512), .B(n3084), .Z(out[507]) );
  XNOR U4989 ( .A(in[882]), .B(n3760), .Z(n3516) );
  NAND U4990 ( .A(n3241), .B(n3085), .Z(n3086) );
  XNOR U4991 ( .A(n3516), .B(n3086), .Z(out[508]) );
  XNOR U4992 ( .A(in[883]), .B(n3764), .Z(n3520) );
  NAND U4993 ( .A(n3243), .B(n3087), .Z(n3088) );
  XNOR U4994 ( .A(n3520), .B(n3088), .Z(out[509]) );
  ANDN U4995 ( .B(n3090), .A(n3089), .Z(n3091) );
  XNOR U4996 ( .A(n3092), .B(n3091), .Z(out[50]) );
  XNOR U4997 ( .A(in[884]), .B(n3768), .Z(n3524) );
  NAND U4998 ( .A(n3245), .B(n3093), .Z(n3094) );
  XNOR U4999 ( .A(n3524), .B(n3094), .Z(out[510]) );
  XNOR U5000 ( .A(in[885]), .B(n3772), .Z(n3528) );
  NAND U5001 ( .A(n3247), .B(n3095), .Z(n3096) );
  XNOR U5002 ( .A(n3528), .B(n3096), .Z(out[511]) );
  OR U5003 ( .A(n3250), .B(n3097), .Z(n3098) );
  XNOR U5004 ( .A(n3249), .B(n3098), .Z(out[512]) );
  OR U5005 ( .A(n3254), .B(n3099), .Z(n3100) );
  XNOR U5006 ( .A(n3253), .B(n3100), .Z(out[513]) );
  OR U5007 ( .A(n3258), .B(n3101), .Z(n3102) );
  XNOR U5008 ( .A(n3257), .B(n3102), .Z(out[514]) );
  OR U5009 ( .A(n3262), .B(n3103), .Z(n3104) );
  XNOR U5010 ( .A(n3261), .B(n3104), .Z(out[515]) );
  OR U5011 ( .A(n3270), .B(n3105), .Z(n3106) );
  XNOR U5012 ( .A(n3269), .B(n3106), .Z(out[516]) );
  OR U5013 ( .A(n3274), .B(n3107), .Z(n3108) );
  XNOR U5014 ( .A(n3273), .B(n3108), .Z(out[517]) );
  OR U5015 ( .A(n3278), .B(n3109), .Z(n3110) );
  XNOR U5016 ( .A(n3277), .B(n3110), .Z(out[518]) );
  OR U5017 ( .A(n3282), .B(n3111), .Z(n3112) );
  XNOR U5018 ( .A(n3281), .B(n3112), .Z(out[519]) );
  ANDN U5019 ( .B(n3114), .A(n3113), .Z(n3115) );
  XNOR U5020 ( .A(n3116), .B(n3115), .Z(out[51]) );
  OR U5021 ( .A(n3286), .B(n3117), .Z(n3118) );
  XNOR U5022 ( .A(n3285), .B(n3118), .Z(out[520]) );
  OR U5023 ( .A(n3290), .B(n3119), .Z(n3120) );
  XNOR U5024 ( .A(n3289), .B(n3120), .Z(out[521]) );
  OR U5025 ( .A(n3294), .B(n3121), .Z(n3122) );
  XNOR U5026 ( .A(n3293), .B(n3122), .Z(out[522]) );
  OR U5027 ( .A(n3298), .B(n3123), .Z(n3124) );
  XNOR U5028 ( .A(n3297), .B(n3124), .Z(out[523]) );
  OR U5029 ( .A(n3302), .B(n3125), .Z(n3126) );
  XNOR U5030 ( .A(n3301), .B(n3126), .Z(out[524]) );
  OR U5031 ( .A(n3306), .B(n3127), .Z(n3128) );
  XNOR U5032 ( .A(n3305), .B(n3128), .Z(out[525]) );
  OR U5033 ( .A(n3314), .B(n3129), .Z(n3130) );
  XNOR U5034 ( .A(n3313), .B(n3130), .Z(out[526]) );
  OR U5035 ( .A(n3318), .B(n3131), .Z(n3132) );
  XNOR U5036 ( .A(n3317), .B(n3132), .Z(out[527]) );
  OR U5037 ( .A(n3322), .B(n3133), .Z(n3134) );
  XNOR U5038 ( .A(n3321), .B(n3134), .Z(out[528]) );
  OR U5039 ( .A(n3326), .B(n3135), .Z(n3136) );
  XNOR U5040 ( .A(n3325), .B(n3136), .Z(out[529]) );
  ANDN U5041 ( .B(n3138), .A(n3137), .Z(n3139) );
  XNOR U5042 ( .A(n3140), .B(n3139), .Z(out[52]) );
  OR U5043 ( .A(n3330), .B(n3141), .Z(n3142) );
  XNOR U5044 ( .A(n3329), .B(n3142), .Z(out[530]) );
  OR U5045 ( .A(n3334), .B(n3143), .Z(n3144) );
  XNOR U5046 ( .A(n3333), .B(n3144), .Z(out[531]) );
  OR U5047 ( .A(n3338), .B(n3145), .Z(n3146) );
  XNOR U5048 ( .A(n3337), .B(n3146), .Z(out[532]) );
  OR U5049 ( .A(n3342), .B(n3147), .Z(n3148) );
  XNOR U5050 ( .A(n3341), .B(n3148), .Z(out[533]) );
  OR U5051 ( .A(n3346), .B(n3149), .Z(n3150) );
  XNOR U5052 ( .A(n3345), .B(n3150), .Z(out[534]) );
  OR U5053 ( .A(n3350), .B(n3151), .Z(n3152) );
  XNOR U5054 ( .A(n3349), .B(n3152), .Z(out[535]) );
  OR U5055 ( .A(n3360), .B(n3153), .Z(n3154) );
  XNOR U5056 ( .A(n3359), .B(n3154), .Z(out[536]) );
  OR U5057 ( .A(n3364), .B(n3155), .Z(n3156) );
  XNOR U5058 ( .A(n3363), .B(n3156), .Z(out[537]) );
  OR U5059 ( .A(n3368), .B(n3157), .Z(n3158) );
  XNOR U5060 ( .A(n3367), .B(n3158), .Z(out[538]) );
  OR U5061 ( .A(n3372), .B(n3159), .Z(n3160) );
  XNOR U5062 ( .A(n3371), .B(n3160), .Z(out[539]) );
  ANDN U5063 ( .B(n3162), .A(n3161), .Z(n3163) );
  XNOR U5064 ( .A(n3164), .B(n3163), .Z(out[53]) );
  OR U5065 ( .A(n3376), .B(n3165), .Z(n3166) );
  XNOR U5066 ( .A(n3375), .B(n3166), .Z(out[540]) );
  OR U5067 ( .A(n3380), .B(n3167), .Z(n3168) );
  XNOR U5068 ( .A(n3379), .B(n3168), .Z(out[541]) );
  OR U5069 ( .A(n3384), .B(n3169), .Z(n3170) );
  XNOR U5070 ( .A(n3383), .B(n3170), .Z(out[542]) );
  OR U5071 ( .A(n3388), .B(n3171), .Z(n3172) );
  XNOR U5072 ( .A(n3387), .B(n3172), .Z(out[543]) );
  OR U5073 ( .A(n3392), .B(n3173), .Z(n3174) );
  XNOR U5074 ( .A(n3391), .B(n3174), .Z(out[544]) );
  OR U5075 ( .A(n3396), .B(n3175), .Z(n3176) );
  XNOR U5076 ( .A(n3395), .B(n3176), .Z(out[545]) );
  OR U5077 ( .A(n3404), .B(n3177), .Z(n3178) );
  XNOR U5078 ( .A(n3403), .B(n3178), .Z(out[546]) );
  OR U5079 ( .A(n3408), .B(n3179), .Z(n3180) );
  XNOR U5080 ( .A(n3407), .B(n3180), .Z(out[547]) );
  OR U5081 ( .A(n3412), .B(n3181), .Z(n3182) );
  XNOR U5082 ( .A(n3411), .B(n3182), .Z(out[548]) );
  OR U5083 ( .A(n3416), .B(n3183), .Z(n3184) );
  XNOR U5084 ( .A(n3415), .B(n3184), .Z(out[549]) );
  ANDN U5085 ( .B(n3186), .A(n3185), .Z(n3187) );
  XNOR U5086 ( .A(n3188), .B(n3187), .Z(out[54]) );
  OR U5087 ( .A(n3420), .B(n3189), .Z(n3190) );
  XNOR U5088 ( .A(n3419), .B(n3190), .Z(out[550]) );
  OR U5089 ( .A(n3424), .B(n3191), .Z(n3192) );
  XNOR U5090 ( .A(n3423), .B(n3192), .Z(out[551]) );
  OR U5091 ( .A(n3428), .B(n3193), .Z(n3194) );
  XNOR U5092 ( .A(n3427), .B(n3194), .Z(out[552]) );
  OR U5093 ( .A(n3432), .B(n3195), .Z(n3196) );
  XNOR U5094 ( .A(n3431), .B(n3196), .Z(out[553]) );
  OR U5095 ( .A(n3436), .B(n3197), .Z(n3198) );
  XNOR U5096 ( .A(n3435), .B(n3198), .Z(out[554]) );
  OR U5097 ( .A(n3440), .B(n3199), .Z(n3200) );
  XNOR U5098 ( .A(n3439), .B(n3200), .Z(out[555]) );
  OR U5099 ( .A(n3448), .B(n3201), .Z(n3202) );
  XNOR U5100 ( .A(n3447), .B(n3202), .Z(out[556]) );
  OR U5101 ( .A(n3452), .B(n3203), .Z(n3204) );
  XNOR U5102 ( .A(n3451), .B(n3204), .Z(out[557]) );
  OR U5103 ( .A(n3456), .B(n3205), .Z(n3206) );
  XNOR U5104 ( .A(n3455), .B(n3206), .Z(out[558]) );
  OR U5105 ( .A(n3460), .B(n3207), .Z(n3208) );
  XNOR U5106 ( .A(n3459), .B(n3208), .Z(out[559]) );
  ANDN U5107 ( .B(n3210), .A(n3209), .Z(n3211) );
  XNOR U5108 ( .A(n3212), .B(n3211), .Z(out[55]) );
  OR U5109 ( .A(n3464), .B(n3213), .Z(n3214) );
  XNOR U5110 ( .A(n3463), .B(n3214), .Z(out[560]) );
  OR U5111 ( .A(n3468), .B(n3215), .Z(n3216) );
  XNOR U5112 ( .A(n3467), .B(n3216), .Z(out[561]) );
  OR U5113 ( .A(n3472), .B(n3217), .Z(n3218) );
  XNOR U5114 ( .A(n3471), .B(n3218), .Z(out[562]) );
  OR U5115 ( .A(n3476), .B(n3219), .Z(n3220) );
  XNOR U5116 ( .A(n3475), .B(n3220), .Z(out[563]) );
  OR U5117 ( .A(n3480), .B(n3221), .Z(n3222) );
  XNOR U5118 ( .A(n3479), .B(n3222), .Z(out[564]) );
  OR U5119 ( .A(n3484), .B(n3223), .Z(n3224) );
  XNOR U5120 ( .A(n3483), .B(n3224), .Z(out[565]) );
  OR U5121 ( .A(n3492), .B(n3225), .Z(n3226) );
  XNOR U5122 ( .A(n3491), .B(n3226), .Z(out[566]) );
  OR U5123 ( .A(n3496), .B(n3227), .Z(n3228) );
  XNOR U5124 ( .A(n3495), .B(n3228), .Z(out[567]) );
  OR U5125 ( .A(n3500), .B(n3229), .Z(n3230) );
  XNOR U5126 ( .A(n3499), .B(n3230), .Z(out[568]) );
  OR U5127 ( .A(n3504), .B(n3231), .Z(n3232) );
  XNOR U5128 ( .A(n3503), .B(n3232), .Z(out[569]) );
  ANDN U5129 ( .B(n3234), .A(n3233), .Z(n3235) );
  XNOR U5130 ( .A(n3236), .B(n3235), .Z(out[56]) );
  OR U5131 ( .A(n3508), .B(n3237), .Z(n3238) );
  XNOR U5132 ( .A(n3507), .B(n3238), .Z(out[570]) );
  OR U5133 ( .A(n3512), .B(n3239), .Z(n3240) );
  XNOR U5134 ( .A(n3511), .B(n3240), .Z(out[571]) );
  OR U5135 ( .A(n3516), .B(n3241), .Z(n3242) );
  XNOR U5136 ( .A(n3515), .B(n3242), .Z(out[572]) );
  OR U5137 ( .A(n3520), .B(n3243), .Z(n3244) );
  XNOR U5138 ( .A(n3519), .B(n3244), .Z(out[573]) );
  OR U5139 ( .A(n3524), .B(n3245), .Z(n3246) );
  XNOR U5140 ( .A(n3523), .B(n3246), .Z(out[574]) );
  OR U5141 ( .A(n3528), .B(n3247), .Z(n3248) );
  XNOR U5142 ( .A(n3527), .B(n3248), .Z(out[575]) );
  ANDN U5143 ( .B(n3250), .A(n3249), .Z(n3251) );
  XNOR U5144 ( .A(n3252), .B(n3251), .Z(out[576]) );
  ANDN U5145 ( .B(n3254), .A(n3253), .Z(n3255) );
  XNOR U5146 ( .A(n3256), .B(n3255), .Z(out[577]) );
  ANDN U5147 ( .B(n3258), .A(n3257), .Z(n3259) );
  XNOR U5148 ( .A(n3260), .B(n3259), .Z(out[578]) );
  ANDN U5149 ( .B(n3262), .A(n3261), .Z(n3263) );
  XNOR U5150 ( .A(n3264), .B(n3263), .Z(out[579]) );
  ANDN U5151 ( .B(n3266), .A(n3265), .Z(n3267) );
  XNOR U5152 ( .A(n3268), .B(n3267), .Z(out[57]) );
  ANDN U5153 ( .B(n3270), .A(n3269), .Z(n3271) );
  XNOR U5154 ( .A(n3272), .B(n3271), .Z(out[580]) );
  ANDN U5155 ( .B(n3274), .A(n3273), .Z(n3275) );
  XNOR U5156 ( .A(n3276), .B(n3275), .Z(out[581]) );
  ANDN U5157 ( .B(n3278), .A(n3277), .Z(n3279) );
  XNOR U5158 ( .A(n3280), .B(n3279), .Z(out[582]) );
  ANDN U5159 ( .B(n3282), .A(n3281), .Z(n3283) );
  XNOR U5160 ( .A(n3284), .B(n3283), .Z(out[583]) );
  ANDN U5161 ( .B(n3286), .A(n3285), .Z(n3287) );
  XNOR U5162 ( .A(n3288), .B(n3287), .Z(out[584]) );
  ANDN U5163 ( .B(n3290), .A(n3289), .Z(n3291) );
  XNOR U5164 ( .A(n3292), .B(n3291), .Z(out[585]) );
  ANDN U5165 ( .B(n3294), .A(n3293), .Z(n3295) );
  XNOR U5166 ( .A(n3296), .B(n3295), .Z(out[586]) );
  ANDN U5167 ( .B(n3298), .A(n3297), .Z(n3299) );
  XNOR U5168 ( .A(n3300), .B(n3299), .Z(out[587]) );
  ANDN U5169 ( .B(n3302), .A(n3301), .Z(n3303) );
  XNOR U5170 ( .A(n3304), .B(n3303), .Z(out[588]) );
  ANDN U5171 ( .B(n3306), .A(n3305), .Z(n3307) );
  XNOR U5172 ( .A(n3308), .B(n3307), .Z(out[589]) );
  ANDN U5173 ( .B(n3310), .A(n3309), .Z(n3311) );
  XNOR U5174 ( .A(n3312), .B(n3311), .Z(out[58]) );
  ANDN U5175 ( .B(n3314), .A(n3313), .Z(n3315) );
  XNOR U5176 ( .A(n3316), .B(n3315), .Z(out[590]) );
  ANDN U5177 ( .B(n3318), .A(n3317), .Z(n3319) );
  XNOR U5178 ( .A(n3320), .B(n3319), .Z(out[591]) );
  ANDN U5179 ( .B(n3322), .A(n3321), .Z(n3323) );
  XNOR U5180 ( .A(n3324), .B(n3323), .Z(out[592]) );
  ANDN U5181 ( .B(n3326), .A(n3325), .Z(n3327) );
  XNOR U5182 ( .A(n3328), .B(n3327), .Z(out[593]) );
  ANDN U5183 ( .B(n3330), .A(n3329), .Z(n3331) );
  XNOR U5184 ( .A(n3332), .B(n3331), .Z(out[594]) );
  ANDN U5185 ( .B(n3334), .A(n3333), .Z(n3335) );
  XNOR U5186 ( .A(n3336), .B(n3335), .Z(out[595]) );
  ANDN U5187 ( .B(n3338), .A(n3337), .Z(n3339) );
  XNOR U5188 ( .A(n3340), .B(n3339), .Z(out[596]) );
  ANDN U5189 ( .B(n3342), .A(n3341), .Z(n3343) );
  XNOR U5190 ( .A(n3344), .B(n3343), .Z(out[597]) );
  ANDN U5191 ( .B(n3346), .A(n3345), .Z(n3347) );
  XNOR U5192 ( .A(n3348), .B(n3347), .Z(out[598]) );
  ANDN U5193 ( .B(n3350), .A(n3349), .Z(n3351) );
  XNOR U5194 ( .A(n3352), .B(n3351), .Z(out[599]) );
  ANDN U5195 ( .B(n3354), .A(n3353), .Z(n3355) );
  XNOR U5196 ( .A(n3356), .B(n3355), .Z(out[59]) );
  OR U5197 ( .A(n3796), .B(n3357), .Z(n3358) );
  XNOR U5198 ( .A(n3795), .B(n3358), .Z(out[5]) );
  ANDN U5199 ( .B(n3360), .A(n3359), .Z(n3361) );
  XNOR U5200 ( .A(n3362), .B(n3361), .Z(out[600]) );
  ANDN U5201 ( .B(n3364), .A(n3363), .Z(n3365) );
  XNOR U5202 ( .A(n3366), .B(n3365), .Z(out[601]) );
  ANDN U5203 ( .B(n3368), .A(n3367), .Z(n3369) );
  XNOR U5204 ( .A(n3370), .B(n3369), .Z(out[602]) );
  ANDN U5205 ( .B(n3372), .A(n3371), .Z(n3373) );
  XNOR U5206 ( .A(n3374), .B(n3373), .Z(out[603]) );
  ANDN U5207 ( .B(n3376), .A(n3375), .Z(n3377) );
  XNOR U5208 ( .A(n3378), .B(n3377), .Z(out[604]) );
  ANDN U5209 ( .B(n3380), .A(n3379), .Z(n3381) );
  XNOR U5210 ( .A(n3382), .B(n3381), .Z(out[605]) );
  ANDN U5211 ( .B(n3384), .A(n3383), .Z(n3385) );
  XNOR U5212 ( .A(n3386), .B(n3385), .Z(out[606]) );
  ANDN U5213 ( .B(n3388), .A(n3387), .Z(n3389) );
  XNOR U5214 ( .A(n3390), .B(n3389), .Z(out[607]) );
  ANDN U5215 ( .B(n3392), .A(n3391), .Z(n3393) );
  XNOR U5216 ( .A(n3394), .B(n3393), .Z(out[608]) );
  ANDN U5217 ( .B(n3396), .A(n3395), .Z(n3397) );
  XNOR U5218 ( .A(n3398), .B(n3397), .Z(out[609]) );
  ANDN U5219 ( .B(n3400), .A(n3399), .Z(n3401) );
  XNOR U5220 ( .A(n3402), .B(n3401), .Z(out[60]) );
  ANDN U5221 ( .B(n3404), .A(n3403), .Z(n3405) );
  XNOR U5222 ( .A(n3406), .B(n3405), .Z(out[610]) );
  ANDN U5223 ( .B(n3408), .A(n3407), .Z(n3409) );
  XNOR U5224 ( .A(n3410), .B(n3409), .Z(out[611]) );
  ANDN U5225 ( .B(n3412), .A(n3411), .Z(n3413) );
  XNOR U5226 ( .A(n3414), .B(n3413), .Z(out[612]) );
  ANDN U5227 ( .B(n3416), .A(n3415), .Z(n3417) );
  XNOR U5228 ( .A(n3418), .B(n3417), .Z(out[613]) );
  ANDN U5229 ( .B(n3420), .A(n3419), .Z(n3421) );
  XNOR U5230 ( .A(n3422), .B(n3421), .Z(out[614]) );
  ANDN U5231 ( .B(n3424), .A(n3423), .Z(n3425) );
  XNOR U5232 ( .A(n3426), .B(n3425), .Z(out[615]) );
  ANDN U5233 ( .B(n3428), .A(n3427), .Z(n3429) );
  XNOR U5234 ( .A(n3430), .B(n3429), .Z(out[616]) );
  ANDN U5235 ( .B(n3432), .A(n3431), .Z(n3433) );
  XNOR U5236 ( .A(n3434), .B(n3433), .Z(out[617]) );
  ANDN U5237 ( .B(n3436), .A(n3435), .Z(n3437) );
  XNOR U5238 ( .A(n3438), .B(n3437), .Z(out[618]) );
  ANDN U5239 ( .B(n3440), .A(n3439), .Z(n3441) );
  XNOR U5240 ( .A(n3442), .B(n3441), .Z(out[619]) );
  ANDN U5241 ( .B(n3444), .A(n3443), .Z(n3445) );
  XNOR U5242 ( .A(n3446), .B(n3445), .Z(out[61]) );
  ANDN U5243 ( .B(n3448), .A(n3447), .Z(n3449) );
  XNOR U5244 ( .A(n3450), .B(n3449), .Z(out[620]) );
  ANDN U5245 ( .B(n3452), .A(n3451), .Z(n3453) );
  XNOR U5246 ( .A(n3454), .B(n3453), .Z(out[621]) );
  ANDN U5247 ( .B(n3456), .A(n3455), .Z(n3457) );
  XNOR U5248 ( .A(n3458), .B(n3457), .Z(out[622]) );
  ANDN U5249 ( .B(n3460), .A(n3459), .Z(n3461) );
  XNOR U5250 ( .A(n3462), .B(n3461), .Z(out[623]) );
  ANDN U5251 ( .B(n3464), .A(n3463), .Z(n3465) );
  XNOR U5252 ( .A(n3466), .B(n3465), .Z(out[624]) );
  ANDN U5253 ( .B(n3468), .A(n3467), .Z(n3469) );
  XNOR U5254 ( .A(n3470), .B(n3469), .Z(out[625]) );
  ANDN U5255 ( .B(n3472), .A(n3471), .Z(n3473) );
  XNOR U5256 ( .A(n3474), .B(n3473), .Z(out[626]) );
  ANDN U5257 ( .B(n3476), .A(n3475), .Z(n3477) );
  XNOR U5258 ( .A(n3478), .B(n3477), .Z(out[627]) );
  ANDN U5259 ( .B(n3480), .A(n3479), .Z(n3481) );
  XNOR U5260 ( .A(n3482), .B(n3481), .Z(out[628]) );
  ANDN U5261 ( .B(n3484), .A(n3483), .Z(n3485) );
  XNOR U5262 ( .A(n3486), .B(n3485), .Z(out[629]) );
  ANDN U5263 ( .B(n3488), .A(n3487), .Z(n3489) );
  XNOR U5264 ( .A(n3490), .B(n3489), .Z(out[62]) );
  ANDN U5265 ( .B(n3492), .A(n3491), .Z(n3493) );
  XNOR U5266 ( .A(n3494), .B(n3493), .Z(out[630]) );
  ANDN U5267 ( .B(n3496), .A(n3495), .Z(n3497) );
  XNOR U5268 ( .A(n3498), .B(n3497), .Z(out[631]) );
  ANDN U5269 ( .B(n3500), .A(n3499), .Z(n3501) );
  XNOR U5270 ( .A(n3502), .B(n3501), .Z(out[632]) );
  ANDN U5271 ( .B(n3504), .A(n3503), .Z(n3505) );
  XNOR U5272 ( .A(n3506), .B(n3505), .Z(out[633]) );
  ANDN U5273 ( .B(n3508), .A(n3507), .Z(n3509) );
  XNOR U5274 ( .A(n3510), .B(n3509), .Z(out[634]) );
  ANDN U5275 ( .B(n3512), .A(n3511), .Z(n3513) );
  XNOR U5276 ( .A(n3514), .B(n3513), .Z(out[635]) );
  ANDN U5277 ( .B(n3516), .A(n3515), .Z(n3517) );
  XNOR U5278 ( .A(n3518), .B(n3517), .Z(out[636]) );
  ANDN U5279 ( .B(n3520), .A(n3519), .Z(n3521) );
  XNOR U5280 ( .A(n3522), .B(n3521), .Z(out[637]) );
  ANDN U5281 ( .B(n3524), .A(n3523), .Z(n3525) );
  XNOR U5282 ( .A(n3526), .B(n3525), .Z(out[638]) );
  ANDN U5283 ( .B(n3528), .A(n3527), .Z(n3529) );
  XNOR U5284 ( .A(n3530), .B(n3529), .Z(out[639]) );
  ANDN U5285 ( .B(n3532), .A(n3531), .Z(n3533) );
  XNOR U5286 ( .A(n3534), .B(n3533), .Z(out[63]) );
  XNOR U5287 ( .A(in[302]), .B(n3535), .Z(n3964) );
  XNOR U5288 ( .A(in[1535]), .B(n3536), .Z(n4342) );
  XNOR U5289 ( .A(in[1146]), .B(n3537), .Z(n4339) );
  NAND U5290 ( .A(n4342), .B(n4339), .Z(n3538) );
  XNOR U5291 ( .A(n3964), .B(n3538), .Z(out[640]) );
  XNOR U5292 ( .A(in[303]), .B(n3539), .Z(n3967) );
  XNOR U5293 ( .A(in[1472]), .B(n3540), .Z(n4346) );
  XNOR U5294 ( .A(in[1147]), .B(n3541), .Z(n4343) );
  NAND U5295 ( .A(n4346), .B(n4343), .Z(n3542) );
  XNOR U5296 ( .A(n3967), .B(n3542), .Z(out[641]) );
  XNOR U5297 ( .A(in[304]), .B(n3543), .Z(n3974) );
  XNOR U5298 ( .A(in[1473]), .B(n3544), .Z(n4350) );
  XNOR U5299 ( .A(in[1148]), .B(n3545), .Z(n4347) );
  NAND U5300 ( .A(n4350), .B(n4347), .Z(n3546) );
  XNOR U5301 ( .A(n3974), .B(n3546), .Z(out[642]) );
  XNOR U5302 ( .A(in[305]), .B(n3547), .Z(n3977) );
  XNOR U5303 ( .A(in[1474]), .B(n3548), .Z(n4354) );
  XNOR U5304 ( .A(in[1149]), .B(n3549), .Z(n4351) );
  NAND U5305 ( .A(n4354), .B(n4351), .Z(n3550) );
  XNOR U5306 ( .A(n3977), .B(n3550), .Z(out[643]) );
  XNOR U5307 ( .A(in[306]), .B(n3551), .Z(n3980) );
  XNOR U5308 ( .A(in[1475]), .B(n3552), .Z(n4366) );
  XNOR U5309 ( .A(in[1150]), .B(n3553), .Z(n4363) );
  NAND U5310 ( .A(n4366), .B(n4363), .Z(n3554) );
  XNOR U5311 ( .A(n3980), .B(n3554), .Z(out[644]) );
  XNOR U5312 ( .A(in[307]), .B(n3555), .Z(n3983) );
  XNOR U5313 ( .A(in[1476]), .B(n3556), .Z(n4370) );
  XNOR U5314 ( .A(in[1151]), .B(n3557), .Z(n4367) );
  NAND U5315 ( .A(n4370), .B(n4367), .Z(n3558) );
  XNOR U5316 ( .A(n3983), .B(n3558), .Z(out[645]) );
  XNOR U5317 ( .A(in[308]), .B(n3559), .Z(n3986) );
  XNOR U5318 ( .A(in[1477]), .B(n3560), .Z(n4374) );
  XNOR U5319 ( .A(in[1088]), .B(n3561), .Z(n4371) );
  NAND U5320 ( .A(n4374), .B(n4371), .Z(n3562) );
  XNOR U5321 ( .A(n3986), .B(n3562), .Z(out[646]) );
  XNOR U5322 ( .A(in[309]), .B(n3563), .Z(n3989) );
  XNOR U5323 ( .A(in[1478]), .B(n3564), .Z(n4378) );
  XNOR U5324 ( .A(in[1089]), .B(n3565), .Z(n4375) );
  NAND U5325 ( .A(n4378), .B(n4375), .Z(n3566) );
  XNOR U5326 ( .A(n3989), .B(n3566), .Z(out[647]) );
  XNOR U5327 ( .A(in[310]), .B(n3567), .Z(n3992) );
  XNOR U5328 ( .A(in[1479]), .B(n3568), .Z(n4382) );
  XOR U5329 ( .A(n3569), .B(in[1090]), .Z(n4379) );
  NAND U5330 ( .A(n4382), .B(n4379), .Z(n3570) );
  XNOR U5331 ( .A(n3992), .B(n3570), .Z(out[648]) );
  XNOR U5332 ( .A(in[311]), .B(n3571), .Z(n3995) );
  XNOR U5333 ( .A(in[1480]), .B(n3572), .Z(n4386) );
  XOR U5334 ( .A(n3573), .B(in[1091]), .Z(n4383) );
  NAND U5335 ( .A(n4386), .B(n4383), .Z(n3574) );
  XNOR U5336 ( .A(n3995), .B(n3574), .Z(out[649]) );
  NOR U5337 ( .A(n3576), .B(n3575), .Z(n3577) );
  XNOR U5338 ( .A(n3578), .B(n3577), .Z(out[64]) );
  XNOR U5339 ( .A(in[312]), .B(n3579), .Z(n3998) );
  XNOR U5340 ( .A(in[1481]), .B(n3580), .Z(n4390) );
  XOR U5341 ( .A(n3581), .B(in[1092]), .Z(n4387) );
  NAND U5342 ( .A(n4390), .B(n4387), .Z(n3582) );
  XNOR U5343 ( .A(n3998), .B(n3582), .Z(out[650]) );
  XNOR U5344 ( .A(in[313]), .B(n3583), .Z(n4001) );
  XNOR U5345 ( .A(in[1482]), .B(n3584), .Z(n4394) );
  XOR U5346 ( .A(n3585), .B(in[1093]), .Z(n4391) );
  NAND U5347 ( .A(n4394), .B(n4391), .Z(n3586) );
  XNOR U5348 ( .A(n4001), .B(n3586), .Z(out[651]) );
  XNOR U5349 ( .A(in[314]), .B(n3587), .Z(n4008) );
  XNOR U5350 ( .A(in[1483]), .B(n3588), .Z(n4398) );
  XOR U5351 ( .A(n3589), .B(in[1094]), .Z(n4395) );
  NAND U5352 ( .A(n4398), .B(n4395), .Z(n3590) );
  XNOR U5353 ( .A(n4008), .B(n3590), .Z(out[652]) );
  XNOR U5354 ( .A(in[315]), .B(n3591), .Z(n4011) );
  XNOR U5355 ( .A(in[1484]), .B(n3592), .Z(n4402) );
  XOR U5356 ( .A(n3593), .B(in[1095]), .Z(n4399) );
  NAND U5357 ( .A(n4402), .B(n4399), .Z(n3594) );
  XNOR U5358 ( .A(n4011), .B(n3594), .Z(out[653]) );
  XNOR U5359 ( .A(in[316]), .B(n3595), .Z(n4014) );
  XNOR U5360 ( .A(in[1485]), .B(n3596), .Z(n4410) );
  XOR U5361 ( .A(n3597), .B(in[1096]), .Z(n4407) );
  NAND U5362 ( .A(n4410), .B(n4407), .Z(n3598) );
  XNOR U5363 ( .A(n4014), .B(n3598), .Z(out[654]) );
  XNOR U5364 ( .A(in[317]), .B(n3599), .Z(n4017) );
  XNOR U5365 ( .A(in[1486]), .B(n3600), .Z(n4414) );
  XOR U5366 ( .A(in[1097]), .B(n3601), .Z(n4411) );
  NAND U5367 ( .A(n4414), .B(n4411), .Z(n3602) );
  XNOR U5368 ( .A(n4017), .B(n3602), .Z(out[655]) );
  XNOR U5369 ( .A(in[318]), .B(n3603), .Z(n4020) );
  XNOR U5370 ( .A(in[1487]), .B(n3604), .Z(n4418) );
  XOR U5371 ( .A(n3605), .B(in[1098]), .Z(n4415) );
  NAND U5372 ( .A(n4418), .B(n4415), .Z(n3606) );
  XNOR U5373 ( .A(n4020), .B(n3606), .Z(out[656]) );
  XNOR U5374 ( .A(in[319]), .B(n3607), .Z(n4023) );
  XNOR U5375 ( .A(in[1488]), .B(n3608), .Z(n4422) );
  XOR U5376 ( .A(n3609), .B(in[1099]), .Z(n4419) );
  NAND U5377 ( .A(n4422), .B(n4419), .Z(n3610) );
  XNOR U5378 ( .A(n4023), .B(n3610), .Z(out[657]) );
  XNOR U5379 ( .A(in[256]), .B(n3611), .Z(n4026) );
  XNOR U5380 ( .A(in[1489]), .B(n3612), .Z(n4426) );
  XOR U5381 ( .A(in[1100]), .B(n3613), .Z(n4423) );
  NAND U5382 ( .A(n4426), .B(n4423), .Z(n3614) );
  XNOR U5383 ( .A(n4026), .B(n3614), .Z(out[658]) );
  XNOR U5384 ( .A(in[257]), .B(n3615), .Z(n4029) );
  XNOR U5385 ( .A(in[1490]), .B(n3616), .Z(n4430) );
  XOR U5386 ( .A(in[1101]), .B(n3617), .Z(n4427) );
  NAND U5387 ( .A(n4430), .B(n4427), .Z(n3618) );
  XNOR U5388 ( .A(n4029), .B(n3618), .Z(out[659]) );
  NOR U5389 ( .A(n3620), .B(n3619), .Z(n3621) );
  XNOR U5390 ( .A(n3622), .B(n3621), .Z(out[65]) );
  XNOR U5391 ( .A(in[258]), .B(n3623), .Z(n4032) );
  XOR U5392 ( .A(in[1491]), .B(n3624), .Z(n4434) );
  XOR U5393 ( .A(in[1102]), .B(n3625), .Z(n4431) );
  NAND U5394 ( .A(n4434), .B(n4431), .Z(n3626) );
  XNOR U5395 ( .A(n4032), .B(n3626), .Z(out[660]) );
  XNOR U5396 ( .A(in[259]), .B(n3627), .Z(n4035) );
  XOR U5397 ( .A(in[1492]), .B(n3628), .Z(n4438) );
  XOR U5398 ( .A(in[1103]), .B(n3629), .Z(n4435) );
  NAND U5399 ( .A(n4438), .B(n4435), .Z(n3630) );
  XNOR U5400 ( .A(n4035), .B(n3630), .Z(out[661]) );
  XOR U5401 ( .A(in[260]), .B(n3631), .Z(n4042) );
  XOR U5402 ( .A(in[1493]), .B(n3632), .Z(n4442) );
  XOR U5403 ( .A(in[1104]), .B(n3633), .Z(n4439) );
  NAND U5404 ( .A(n4442), .B(n4439), .Z(n3634) );
  XNOR U5405 ( .A(n4042), .B(n3634), .Z(out[662]) );
  XOR U5406 ( .A(in[261]), .B(n3635), .Z(n4045) );
  XOR U5407 ( .A(in[1494]), .B(n3636), .Z(n4446) );
  XOR U5408 ( .A(in[1105]), .B(n3637), .Z(n4443) );
  NAND U5409 ( .A(n4446), .B(n4443), .Z(n3638) );
  XNOR U5410 ( .A(n4045), .B(n3638), .Z(out[663]) );
  XOR U5411 ( .A(in[262]), .B(n3639), .Z(n4048) );
  XOR U5412 ( .A(in[1495]), .B(n3640), .Z(n4454) );
  XOR U5413 ( .A(in[1106]), .B(n3641), .Z(n4451) );
  NAND U5414 ( .A(n4454), .B(n4451), .Z(n3642) );
  XNOR U5415 ( .A(n4048), .B(n3642), .Z(out[664]) );
  XOR U5416 ( .A(in[263]), .B(n3643), .Z(n4051) );
  XOR U5417 ( .A(in[1496]), .B(n3644), .Z(n4458) );
  XOR U5418 ( .A(in[1107]), .B(n3645), .Z(n4455) );
  NAND U5419 ( .A(n4458), .B(n4455), .Z(n3646) );
  XNOR U5420 ( .A(n4051), .B(n3646), .Z(out[665]) );
  XOR U5421 ( .A(in[264]), .B(n3647), .Z(n4054) );
  XOR U5422 ( .A(in[1497]), .B(n3648), .Z(n4462) );
  XOR U5423 ( .A(in[1108]), .B(n3649), .Z(n4459) );
  NAND U5424 ( .A(n4462), .B(n4459), .Z(n3650) );
  XNOR U5425 ( .A(n4054), .B(n3650), .Z(out[666]) );
  XOR U5426 ( .A(in[265]), .B(n3651), .Z(n4057) );
  XOR U5427 ( .A(in[1498]), .B(n3652), .Z(n4466) );
  XOR U5428 ( .A(in[1109]), .B(n3653), .Z(n4463) );
  NAND U5429 ( .A(n4466), .B(n4463), .Z(n3654) );
  XNOR U5430 ( .A(n4057), .B(n3654), .Z(out[667]) );
  XOR U5431 ( .A(in[266]), .B(n3655), .Z(n4060) );
  XOR U5432 ( .A(in[1499]), .B(n3656), .Z(n4470) );
  XOR U5433 ( .A(in[1110]), .B(n3657), .Z(n4467) );
  NAND U5434 ( .A(n4470), .B(n4467), .Z(n3658) );
  XNOR U5435 ( .A(n4060), .B(n3658), .Z(out[668]) );
  XOR U5436 ( .A(in[267]), .B(n3659), .Z(n4063) );
  XOR U5437 ( .A(in[1500]), .B(n3660), .Z(n4474) );
  XOR U5438 ( .A(in[1111]), .B(n3661), .Z(n4471) );
  NAND U5439 ( .A(n4474), .B(n4471), .Z(n3662) );
  XNOR U5440 ( .A(n4063), .B(n3662), .Z(out[669]) );
  ANDN U5441 ( .B(n3664), .A(n3663), .Z(n3665) );
  XNOR U5442 ( .A(n3666), .B(n3665), .Z(out[66]) );
  XOR U5443 ( .A(in[268]), .B(n3667), .Z(n4066) );
  XOR U5444 ( .A(in[1501]), .B(n3668), .Z(n4478) );
  XOR U5445 ( .A(in[1112]), .B(n3669), .Z(n4475) );
  NAND U5446 ( .A(n4478), .B(n4475), .Z(n3670) );
  XNOR U5447 ( .A(n4066), .B(n3670), .Z(out[670]) );
  XOR U5448 ( .A(in[269]), .B(n3671), .Z(n4069) );
  XOR U5449 ( .A(in[1502]), .B(n3672), .Z(n4482) );
  XOR U5450 ( .A(in[1113]), .B(n3673), .Z(n4479) );
  NAND U5451 ( .A(n4482), .B(n4479), .Z(n3674) );
  XNOR U5452 ( .A(n4069), .B(n3674), .Z(out[671]) );
  XOR U5453 ( .A(in[270]), .B(n3675), .Z(n4080) );
  XOR U5454 ( .A(in[1503]), .B(n3676), .Z(n4486) );
  XOR U5455 ( .A(in[1114]), .B(n3677), .Z(n4483) );
  NAND U5456 ( .A(n4486), .B(n4483), .Z(n3678) );
  XNOR U5457 ( .A(n4080), .B(n3678), .Z(out[672]) );
  XOR U5458 ( .A(in[271]), .B(n3679), .Z(n4083) );
  XOR U5459 ( .A(in[1504]), .B(n3680), .Z(n4490) );
  XOR U5460 ( .A(in[1115]), .B(n3681), .Z(n4487) );
  NAND U5461 ( .A(n4490), .B(n4487), .Z(n3682) );
  XNOR U5462 ( .A(n4083), .B(n3682), .Z(out[673]) );
  XOR U5463 ( .A(in[272]), .B(n3683), .Z(n4086) );
  XOR U5464 ( .A(in[1505]), .B(n3684), .Z(n4498) );
  XOR U5465 ( .A(in[1116]), .B(n3685), .Z(n4495) );
  NAND U5466 ( .A(n4498), .B(n4495), .Z(n3686) );
  XNOR U5467 ( .A(n4086), .B(n3686), .Z(out[674]) );
  XOR U5468 ( .A(in[273]), .B(n3687), .Z(n4089) );
  XNOR U5469 ( .A(n3688), .B(in[1506]), .Z(n4502) );
  XOR U5470 ( .A(in[1117]), .B(n3689), .Z(n4499) );
  NAND U5471 ( .A(n4502), .B(n4499), .Z(n3690) );
  XNOR U5472 ( .A(n4089), .B(n3690), .Z(out[675]) );
  XOR U5473 ( .A(in[274]), .B(n3691), .Z(n4092) );
  XNOR U5474 ( .A(n3692), .B(in[1507]), .Z(n4506) );
  XOR U5475 ( .A(in[1118]), .B(n3693), .Z(n4503) );
  NAND U5476 ( .A(n4506), .B(n4503), .Z(n3694) );
  XNOR U5477 ( .A(n4092), .B(n3694), .Z(out[676]) );
  XOR U5478 ( .A(in[275]), .B(n3695), .Z(n4095) );
  XNOR U5479 ( .A(n3696), .B(in[1508]), .Z(n4510) );
  XOR U5480 ( .A(in[1119]), .B(n3697), .Z(n4507) );
  NAND U5481 ( .A(n4510), .B(n4507), .Z(n3698) );
  XNOR U5482 ( .A(n4095), .B(n3698), .Z(out[677]) );
  XOR U5483 ( .A(in[276]), .B(n3699), .Z(n4098) );
  XNOR U5484 ( .A(n3700), .B(in[1509]), .Z(n4514) );
  XOR U5485 ( .A(in[1120]), .B(n3701), .Z(n4511) );
  NAND U5486 ( .A(n4514), .B(n4511), .Z(n3702) );
  XNOR U5487 ( .A(n4098), .B(n3702), .Z(out[678]) );
  XOR U5488 ( .A(in[277]), .B(n3703), .Z(n4101) );
  XOR U5489 ( .A(in[1510]), .B(n3704), .Z(n4518) );
  XOR U5490 ( .A(in[1121]), .B(n3705), .Z(n4515) );
  NAND U5491 ( .A(n4518), .B(n4515), .Z(n3706) );
  XNOR U5492 ( .A(n4101), .B(n3706), .Z(out[679]) );
  ANDN U5493 ( .B(n3708), .A(n3707), .Z(n3709) );
  XNOR U5494 ( .A(n3710), .B(n3709), .Z(out[67]) );
  XOR U5495 ( .A(in[278]), .B(n3711), .Z(n4104) );
  XOR U5496 ( .A(in[1511]), .B(n3712), .Z(n4522) );
  XOR U5497 ( .A(in[1122]), .B(n3713), .Z(n4519) );
  NAND U5498 ( .A(n4522), .B(n4519), .Z(n3714) );
  XNOR U5499 ( .A(n4104), .B(n3714), .Z(out[680]) );
  XOR U5500 ( .A(in[279]), .B(n3715), .Z(n4107) );
  XOR U5501 ( .A(in[1512]), .B(n3716), .Z(n4526) );
  XOR U5502 ( .A(in[1123]), .B(n3717), .Z(n4523) );
  NAND U5503 ( .A(n4526), .B(n4523), .Z(n3718) );
  XNOR U5504 ( .A(n4107), .B(n3718), .Z(out[681]) );
  XOR U5505 ( .A(in[280]), .B(n3719), .Z(n4114) );
  XOR U5506 ( .A(in[1513]), .B(n3720), .Z(n4530) );
  XOR U5507 ( .A(in[1124]), .B(n3721), .Z(n4527) );
  NAND U5508 ( .A(n4530), .B(n4527), .Z(n3722) );
  XNOR U5509 ( .A(n4114), .B(n3722), .Z(out[682]) );
  XOR U5510 ( .A(in[281]), .B(n3723), .Z(n4117) );
  XOR U5511 ( .A(in[1514]), .B(n3724), .Z(n4534) );
  XOR U5512 ( .A(in[1125]), .B(n3725), .Z(n4531) );
  NAND U5513 ( .A(n4534), .B(n4531), .Z(n3726) );
  XNOR U5514 ( .A(n4117), .B(n3726), .Z(out[683]) );
  XOR U5515 ( .A(in[282]), .B(n3727), .Z(n4120) );
  XOR U5516 ( .A(in[1515]), .B(n3728), .Z(n4542) );
  XNOR U5517 ( .A(in[1126]), .B(n3729), .Z(n4539) );
  NAND U5518 ( .A(n4542), .B(n4539), .Z(n3730) );
  XNOR U5519 ( .A(n4120), .B(n3730), .Z(out[684]) );
  XOR U5520 ( .A(in[283]), .B(n3731), .Z(n4123) );
  XOR U5521 ( .A(in[1516]), .B(n3732), .Z(n4546) );
  XNOR U5522 ( .A(in[1127]), .B(n3733), .Z(n4543) );
  NAND U5523 ( .A(n4546), .B(n4543), .Z(n3734) );
  XNOR U5524 ( .A(n4123), .B(n3734), .Z(out[685]) );
  XOR U5525 ( .A(in[284]), .B(n3735), .Z(n4126) );
  XOR U5526 ( .A(in[1517]), .B(n3736), .Z(n4550) );
  XNOR U5527 ( .A(in[1128]), .B(n3737), .Z(n4547) );
  NAND U5528 ( .A(n4550), .B(n4547), .Z(n3738) );
  XNOR U5529 ( .A(n4126), .B(n3738), .Z(out[686]) );
  XOR U5530 ( .A(in[285]), .B(n3739), .Z(n4129) );
  XOR U5531 ( .A(in[1518]), .B(n3740), .Z(n4554) );
  XNOR U5532 ( .A(in[1129]), .B(n3741), .Z(n4551) );
  NAND U5533 ( .A(n4554), .B(n4551), .Z(n3742) );
  XNOR U5534 ( .A(n4129), .B(n3742), .Z(out[687]) );
  XOR U5535 ( .A(in[286]), .B(n3743), .Z(n4132) );
  XOR U5536 ( .A(in[1519]), .B(n3744), .Z(n4558) );
  XNOR U5537 ( .A(in[1130]), .B(n3745), .Z(n4555) );
  NAND U5538 ( .A(n4558), .B(n4555), .Z(n3746) );
  XNOR U5539 ( .A(n4132), .B(n3746), .Z(out[688]) );
  XOR U5540 ( .A(in[287]), .B(n3747), .Z(n4135) );
  XOR U5541 ( .A(in[1520]), .B(n3748), .Z(n4562) );
  XNOR U5542 ( .A(in[1131]), .B(n3749), .Z(n4559) );
  NAND U5543 ( .A(n4562), .B(n4559), .Z(n3750) );
  XNOR U5544 ( .A(n4135), .B(n3750), .Z(out[689]) );
  ANDN U5545 ( .B(n3752), .A(n3751), .Z(n3753) );
  XNOR U5546 ( .A(n3754), .B(n3753), .Z(out[68]) );
  XOR U5547 ( .A(in[288]), .B(n3755), .Z(n4138) );
  XOR U5548 ( .A(in[1521]), .B(n3756), .Z(n4566) );
  XNOR U5549 ( .A(in[1132]), .B(n3757), .Z(n4563) );
  NAND U5550 ( .A(n4566), .B(n4563), .Z(n3758) );
  XNOR U5551 ( .A(n4138), .B(n3758), .Z(out[690]) );
  XOR U5552 ( .A(in[289]), .B(n3759), .Z(n4141) );
  XOR U5553 ( .A(in[1522]), .B(n3760), .Z(n4570) );
  XNOR U5554 ( .A(in[1133]), .B(n3761), .Z(n4567) );
  NAND U5555 ( .A(n4570), .B(n4567), .Z(n3762) );
  XNOR U5556 ( .A(n4141), .B(n3762), .Z(out[691]) );
  XOR U5557 ( .A(in[290]), .B(n3763), .Z(n4148) );
  XOR U5558 ( .A(in[1523]), .B(n3764), .Z(n4574) );
  XNOR U5559 ( .A(in[1134]), .B(n3765), .Z(n4571) );
  NAND U5560 ( .A(n4574), .B(n4571), .Z(n3766) );
  XNOR U5561 ( .A(n4148), .B(n3766), .Z(out[692]) );
  XOR U5562 ( .A(in[291]), .B(n3767), .Z(n4151) );
  XOR U5563 ( .A(in[1524]), .B(n3768), .Z(n4578) );
  XNOR U5564 ( .A(in[1135]), .B(n3769), .Z(n4575) );
  NAND U5565 ( .A(n4578), .B(n4575), .Z(n3770) );
  XNOR U5566 ( .A(n4151), .B(n3770), .Z(out[693]) );
  XOR U5567 ( .A(in[292]), .B(n3771), .Z(n4154) );
  XOR U5568 ( .A(in[1525]), .B(n3772), .Z(n4586) );
  XNOR U5569 ( .A(in[1136]), .B(n3773), .Z(n4583) );
  NAND U5570 ( .A(n4586), .B(n4583), .Z(n3774) );
  XNOR U5571 ( .A(n4154), .B(n3774), .Z(out[694]) );
  XNOR U5572 ( .A(in[293]), .B(n3775), .Z(n4157) );
  XOR U5573 ( .A(in[1526]), .B(n3776), .Z(n4590) );
  XNOR U5574 ( .A(in[1137]), .B(n3777), .Z(n4587) );
  NAND U5575 ( .A(n4590), .B(n4587), .Z(n3778) );
  XNOR U5576 ( .A(n4157), .B(n3778), .Z(out[695]) );
  XNOR U5577 ( .A(in[294]), .B(n3779), .Z(n4160) );
  XOR U5578 ( .A(in[1527]), .B(n3780), .Z(n4594) );
  XNOR U5579 ( .A(in[1138]), .B(n3781), .Z(n4591) );
  NAND U5580 ( .A(n4594), .B(n4591), .Z(n3782) );
  XNOR U5581 ( .A(n4160), .B(n3782), .Z(out[696]) );
  XNOR U5582 ( .A(in[295]), .B(n3783), .Z(n4163) );
  XOR U5583 ( .A(in[1528]), .B(n3784), .Z(n4598) );
  XNOR U5584 ( .A(in[1139]), .B(n3785), .Z(n4595) );
  NAND U5585 ( .A(n4598), .B(n4595), .Z(n3786) );
  XNOR U5586 ( .A(n4163), .B(n3786), .Z(out[697]) );
  XNOR U5587 ( .A(in[296]), .B(n3787), .Z(n4166) );
  XOR U5588 ( .A(in[1529]), .B(n3788), .Z(n4602) );
  XNOR U5589 ( .A(in[1140]), .B(n3789), .Z(n4599) );
  NAND U5590 ( .A(n4602), .B(n4599), .Z(n3790) );
  XNOR U5591 ( .A(n4166), .B(n3790), .Z(out[698]) );
  XNOR U5592 ( .A(in[297]), .B(n3791), .Z(n4169) );
  XOR U5593 ( .A(in[1530]), .B(n3792), .Z(n4606) );
  XNOR U5594 ( .A(in[1141]), .B(n3793), .Z(n4603) );
  NAND U5595 ( .A(n4606), .B(n4603), .Z(n3794) );
  XNOR U5596 ( .A(n4169), .B(n3794), .Z(out[699]) );
  ANDN U5597 ( .B(n3796), .A(n3795), .Z(n3797) );
  XNOR U5598 ( .A(n3798), .B(n3797), .Z(out[69]) );
  OR U5599 ( .A(n3830), .B(n3799), .Z(n3800) );
  XNOR U5600 ( .A(n3829), .B(n3800), .Z(out[6]) );
  XNOR U5601 ( .A(in[298]), .B(n3801), .Z(n4172) );
  XNOR U5602 ( .A(in[1531]), .B(n3802), .Z(n4610) );
  XNOR U5603 ( .A(in[1142]), .B(n3803), .Z(n4607) );
  NAND U5604 ( .A(n4610), .B(n4607), .Z(n3804) );
  XNOR U5605 ( .A(n4172), .B(n3804), .Z(out[700]) );
  XNOR U5606 ( .A(in[299]), .B(n3805), .Z(n4175) );
  XNOR U5607 ( .A(in[1532]), .B(n3806), .Z(n4614) );
  XNOR U5608 ( .A(in[1143]), .B(n3807), .Z(n4611) );
  NAND U5609 ( .A(n4614), .B(n4611), .Z(n3808) );
  XNOR U5610 ( .A(n4175), .B(n3808), .Z(out[701]) );
  XNOR U5611 ( .A(in[300]), .B(n3809), .Z(n4182) );
  XNOR U5612 ( .A(in[1533]), .B(n3810), .Z(n4618) );
  XNOR U5613 ( .A(in[1144]), .B(n3811), .Z(n4615) );
  NAND U5614 ( .A(n4618), .B(n4615), .Z(n3812) );
  XNOR U5615 ( .A(n4182), .B(n3812), .Z(out[702]) );
  XNOR U5616 ( .A(in[301]), .B(n3813), .Z(n4185) );
  XOR U5617 ( .A(in[1534]), .B(n3814), .Z(n4622) );
  XNOR U5618 ( .A(in[1145]), .B(n3815), .Z(n4619) );
  NAND U5619 ( .A(n4622), .B(n4619), .Z(n3816) );
  XNOR U5620 ( .A(n4185), .B(n3816), .Z(out[703]) );
  XOR U5621 ( .A(in[376]), .B(n3817), .Z(n4187) );
  NOR U5622 ( .A(n3964), .B(n4342), .Z(n3818) );
  XNOR U5623 ( .A(n4187), .B(n3818), .Z(out[704]) );
  XOR U5624 ( .A(in[377]), .B(n3819), .Z(n4189) );
  NOR U5625 ( .A(n3967), .B(n4346), .Z(n3820) );
  XNOR U5626 ( .A(n4189), .B(n3820), .Z(out[705]) );
  XOR U5627 ( .A(in[378]), .B(n3821), .Z(n4191) );
  NOR U5628 ( .A(n3974), .B(n4350), .Z(n3822) );
  XNOR U5629 ( .A(n4191), .B(n3822), .Z(out[706]) );
  XOR U5630 ( .A(in[379]), .B(n3823), .Z(n4193) );
  NOR U5631 ( .A(n3977), .B(n4354), .Z(n3824) );
  XNOR U5632 ( .A(n4193), .B(n3824), .Z(out[707]) );
  XOR U5633 ( .A(in[380]), .B(n3825), .Z(n4195) );
  NOR U5634 ( .A(n3980), .B(n4366), .Z(n3826) );
  XNOR U5635 ( .A(n4195), .B(n3826), .Z(out[708]) );
  XOR U5636 ( .A(in[381]), .B(n3827), .Z(n4197) );
  NOR U5637 ( .A(n3983), .B(n4370), .Z(n3828) );
  XNOR U5638 ( .A(n4197), .B(n3828), .Z(out[709]) );
  ANDN U5639 ( .B(n3830), .A(n3829), .Z(n3831) );
  XNOR U5640 ( .A(n3832), .B(n3831), .Z(out[70]) );
  XOR U5641 ( .A(in[382]), .B(n3833), .Z(n4199) );
  NOR U5642 ( .A(n3986), .B(n4374), .Z(n3834) );
  XNOR U5643 ( .A(n4199), .B(n3834), .Z(out[710]) );
  XOR U5644 ( .A(in[383]), .B(n3835), .Z(n4201) );
  NOR U5645 ( .A(n3989), .B(n4378), .Z(n3836) );
  XNOR U5646 ( .A(n4201), .B(n3836), .Z(out[711]) );
  XOR U5647 ( .A(in[320]), .B(n3837), .Z(n4207) );
  NOR U5648 ( .A(n3992), .B(n4382), .Z(n3838) );
  XNOR U5649 ( .A(n4207), .B(n3838), .Z(out[712]) );
  XOR U5650 ( .A(in[321]), .B(n3839), .Z(n4209) );
  NOR U5651 ( .A(n3995), .B(n4386), .Z(n3840) );
  XNOR U5652 ( .A(n4209), .B(n3840), .Z(out[713]) );
  XOR U5653 ( .A(in[322]), .B(n3841), .Z(n4211) );
  NOR U5654 ( .A(n3998), .B(n4390), .Z(n3842) );
  XNOR U5655 ( .A(n4211), .B(n3842), .Z(out[714]) );
  XOR U5656 ( .A(in[323]), .B(n3843), .Z(n4213) );
  NOR U5657 ( .A(n4001), .B(n4394), .Z(n3844) );
  XNOR U5658 ( .A(n4213), .B(n3844), .Z(out[715]) );
  XOR U5659 ( .A(in[324]), .B(n3845), .Z(n4215) );
  NOR U5660 ( .A(n4008), .B(n4398), .Z(n3846) );
  XNOR U5661 ( .A(n4215), .B(n3846), .Z(out[716]) );
  XOR U5662 ( .A(in[325]), .B(n3847), .Z(n4217) );
  NOR U5663 ( .A(n4011), .B(n4402), .Z(n3848) );
  XNOR U5664 ( .A(n4217), .B(n3848), .Z(out[717]) );
  XOR U5665 ( .A(in[326]), .B(n3849), .Z(n4219) );
  NOR U5666 ( .A(n4014), .B(n4410), .Z(n3850) );
  XNOR U5667 ( .A(n4219), .B(n3850), .Z(out[718]) );
  XOR U5668 ( .A(in[327]), .B(n3851), .Z(n4221) );
  NOR U5669 ( .A(n4017), .B(n4414), .Z(n3852) );
  XNOR U5670 ( .A(n4221), .B(n3852), .Z(out[719]) );
  ANDN U5671 ( .B(n4076), .A(n4078), .Z(n3853) );
  XNOR U5672 ( .A(n3854), .B(n3853), .Z(out[71]) );
  XOR U5673 ( .A(in[328]), .B(n3855), .Z(n4223) );
  NOR U5674 ( .A(n4020), .B(n4418), .Z(n3856) );
  XNOR U5675 ( .A(n4223), .B(n3856), .Z(out[720]) );
  XOR U5676 ( .A(in[329]), .B(n3857), .Z(n4225) );
  NOR U5677 ( .A(n4023), .B(n4422), .Z(n3858) );
  XNOR U5678 ( .A(n4225), .B(n3858), .Z(out[721]) );
  XOR U5679 ( .A(in[330]), .B(n3859), .Z(n4231) );
  NOR U5680 ( .A(n4026), .B(n4426), .Z(n3860) );
  XNOR U5681 ( .A(n4231), .B(n3860), .Z(out[722]) );
  XOR U5682 ( .A(in[331]), .B(n3861), .Z(n4233) );
  NOR U5683 ( .A(n4029), .B(n4430), .Z(n3862) );
  XNOR U5684 ( .A(n4233), .B(n3862), .Z(out[723]) );
  XOR U5685 ( .A(in[332]), .B(n3863), .Z(n4235) );
  NOR U5686 ( .A(n4032), .B(n4434), .Z(n3864) );
  XNOR U5687 ( .A(n4235), .B(n3864), .Z(out[724]) );
  XOR U5688 ( .A(in[333]), .B(n3865), .Z(n4237) );
  NOR U5689 ( .A(n4035), .B(n4438), .Z(n3866) );
  XNOR U5690 ( .A(n4237), .B(n3866), .Z(out[725]) );
  XOR U5691 ( .A(in[334]), .B(n3867), .Z(n4239) );
  NOR U5692 ( .A(n4042), .B(n4442), .Z(n3868) );
  XNOR U5693 ( .A(n4239), .B(n3868), .Z(out[726]) );
  XOR U5694 ( .A(in[335]), .B(n3869), .Z(n4241) );
  NOR U5695 ( .A(n4045), .B(n4446), .Z(n3870) );
  XNOR U5696 ( .A(n4241), .B(n3870), .Z(out[727]) );
  XOR U5697 ( .A(in[336]), .B(n3871), .Z(n4243) );
  NOR U5698 ( .A(n4048), .B(n4454), .Z(n3872) );
  XNOR U5699 ( .A(n4243), .B(n3872), .Z(out[728]) );
  XOR U5700 ( .A(in[337]), .B(n3873), .Z(n4245) );
  NOR U5701 ( .A(n4051), .B(n4458), .Z(n3874) );
  XNOR U5702 ( .A(n4245), .B(n3874), .Z(out[729]) );
  ANDN U5703 ( .B(n4360), .A(n4362), .Z(n3875) );
  XNOR U5704 ( .A(n3876), .B(n3875), .Z(out[72]) );
  XOR U5705 ( .A(in[338]), .B(n3877), .Z(n4247) );
  NOR U5706 ( .A(n4054), .B(n4462), .Z(n3878) );
  XNOR U5707 ( .A(n4247), .B(n3878), .Z(out[730]) );
  XOR U5708 ( .A(in[339]), .B(n3879), .Z(n4249) );
  NOR U5709 ( .A(n4057), .B(n4466), .Z(n3880) );
  XNOR U5710 ( .A(n4249), .B(n3880), .Z(out[731]) );
  XOR U5711 ( .A(in[340]), .B(n3881), .Z(n4255) );
  NOR U5712 ( .A(n4060), .B(n4470), .Z(n3882) );
  XNOR U5713 ( .A(n4255), .B(n3882), .Z(out[732]) );
  XOR U5714 ( .A(in[341]), .B(n3883), .Z(n4257) );
  NOR U5715 ( .A(n4063), .B(n4474), .Z(n3884) );
  XNOR U5716 ( .A(n4257), .B(n3884), .Z(out[733]) );
  XOR U5717 ( .A(in[342]), .B(n3885), .Z(n4259) );
  NOR U5718 ( .A(n4066), .B(n4478), .Z(n3886) );
  XNOR U5719 ( .A(n4259), .B(n3886), .Z(out[734]) );
  XOR U5720 ( .A(in[343]), .B(n3887), .Z(n4261) );
  NOR U5721 ( .A(n4069), .B(n4482), .Z(n3888) );
  XNOR U5722 ( .A(n4261), .B(n3888), .Z(out[735]) );
  XOR U5723 ( .A(in[344]), .B(n3889), .Z(n4263) );
  NOR U5724 ( .A(n4080), .B(n4486), .Z(n3890) );
  XNOR U5725 ( .A(n4263), .B(n3890), .Z(out[736]) );
  XOR U5726 ( .A(in[345]), .B(n3891), .Z(n4265) );
  NOR U5727 ( .A(n4083), .B(n4490), .Z(n3892) );
  XNOR U5728 ( .A(n4265), .B(n3892), .Z(out[737]) );
  XOR U5729 ( .A(in[346]), .B(n3893), .Z(n4267) );
  NOR U5730 ( .A(n4086), .B(n4498), .Z(n3894) );
  XNOR U5731 ( .A(n4267), .B(n3894), .Z(out[738]) );
  XOR U5732 ( .A(in[347]), .B(n3895), .Z(n4269) );
  NOR U5733 ( .A(n4089), .B(n4502), .Z(n3896) );
  XNOR U5734 ( .A(n4269), .B(n3896), .Z(out[739]) );
  ANDN U5735 ( .B(n4804), .A(n4806), .Z(n3897) );
  XNOR U5736 ( .A(n3898), .B(n3897), .Z(out[73]) );
  XOR U5737 ( .A(in[348]), .B(n3899), .Z(n4271) );
  NOR U5738 ( .A(n4092), .B(n4506), .Z(n3900) );
  XNOR U5739 ( .A(n4271), .B(n3900), .Z(out[740]) );
  XOR U5740 ( .A(in[349]), .B(n3901), .Z(n4273) );
  NOR U5741 ( .A(n4095), .B(n4510), .Z(n3902) );
  XNOR U5742 ( .A(n4273), .B(n3902), .Z(out[741]) );
  XOR U5743 ( .A(in[350]), .B(n3903), .Z(n4279) );
  NOR U5744 ( .A(n4098), .B(n4514), .Z(n3904) );
  XNOR U5745 ( .A(n4279), .B(n3904), .Z(out[742]) );
  XOR U5746 ( .A(in[351]), .B(n3905), .Z(n4281) );
  NOR U5747 ( .A(n4101), .B(n4518), .Z(n3906) );
  XNOR U5748 ( .A(n4281), .B(n3906), .Z(out[743]) );
  XOR U5749 ( .A(in[352]), .B(n3907), .Z(n4283) );
  NOR U5750 ( .A(n4104), .B(n4522), .Z(n3908) );
  XNOR U5751 ( .A(n4283), .B(n3908), .Z(out[744]) );
  XOR U5752 ( .A(in[353]), .B(n3909), .Z(n4285) );
  NOR U5753 ( .A(n4107), .B(n4526), .Z(n3910) );
  XNOR U5754 ( .A(n4285), .B(n3910), .Z(out[745]) );
  XOR U5755 ( .A(in[354]), .B(n3911), .Z(n4287) );
  NOR U5756 ( .A(n4114), .B(n4530), .Z(n3912) );
  XNOR U5757 ( .A(n4287), .B(n3912), .Z(out[746]) );
  XOR U5758 ( .A(in[355]), .B(n3913), .Z(n4289) );
  NOR U5759 ( .A(n4117), .B(n4534), .Z(n3914) );
  XNOR U5760 ( .A(n4289), .B(n3914), .Z(out[747]) );
  XOR U5761 ( .A(in[356]), .B(n3915), .Z(n4291) );
  NOR U5762 ( .A(n4120), .B(n4542), .Z(n3916) );
  XNOR U5763 ( .A(n4291), .B(n3916), .Z(out[748]) );
  XOR U5764 ( .A(in[357]), .B(n3917), .Z(n4293) );
  NOR U5765 ( .A(n4123), .B(n4546), .Z(n3918) );
  XNOR U5766 ( .A(n4293), .B(n3918), .Z(out[749]) );
  NOR U5767 ( .A(n3920), .B(n3919), .Z(n3921) );
  XNOR U5768 ( .A(n3922), .B(n3921), .Z(out[74]) );
  XOR U5769 ( .A(in[358]), .B(n3923), .Z(n4295) );
  NOR U5770 ( .A(n4126), .B(n4550), .Z(n3924) );
  XNOR U5771 ( .A(n4295), .B(n3924), .Z(out[750]) );
  XOR U5772 ( .A(in[359]), .B(n3925), .Z(n4297) );
  NOR U5773 ( .A(n4129), .B(n4554), .Z(n3926) );
  XNOR U5774 ( .A(n4297), .B(n3926), .Z(out[751]) );
  XOR U5775 ( .A(in[360]), .B(n3927), .Z(n4303) );
  NOR U5776 ( .A(n4132), .B(n4558), .Z(n3928) );
  XNOR U5777 ( .A(n4303), .B(n3928), .Z(out[752]) );
  XOR U5778 ( .A(in[361]), .B(n3929), .Z(n4305) );
  NOR U5779 ( .A(n4135), .B(n4562), .Z(n3930) );
  XNOR U5780 ( .A(n4305), .B(n3930), .Z(out[753]) );
  XOR U5781 ( .A(in[362]), .B(n3931), .Z(n4307) );
  NOR U5782 ( .A(n4138), .B(n4566), .Z(n3932) );
  XNOR U5783 ( .A(n4307), .B(n3932), .Z(out[754]) );
  XOR U5784 ( .A(in[363]), .B(n3933), .Z(n4309) );
  NOR U5785 ( .A(n4141), .B(n4570), .Z(n3934) );
  XNOR U5786 ( .A(n4309), .B(n3934), .Z(out[755]) );
  XOR U5787 ( .A(in[364]), .B(n3935), .Z(n4311) );
  NOR U5788 ( .A(n4148), .B(n4574), .Z(n3936) );
  XNOR U5789 ( .A(n4311), .B(n3936), .Z(out[756]) );
  XOR U5790 ( .A(in[365]), .B(n3937), .Z(n4313) );
  NOR U5791 ( .A(n4151), .B(n4578), .Z(n3938) );
  XNOR U5792 ( .A(n4313), .B(n3938), .Z(out[757]) );
  XOR U5793 ( .A(in[366]), .B(n3939), .Z(n4315) );
  NOR U5794 ( .A(n4154), .B(n4586), .Z(n3940) );
  XNOR U5795 ( .A(n4315), .B(n3940), .Z(out[758]) );
  XOR U5796 ( .A(in[367]), .B(n3941), .Z(n4317) );
  NOR U5797 ( .A(n4157), .B(n4590), .Z(n3942) );
  XNOR U5798 ( .A(n4317), .B(n3942), .Z(out[759]) );
  NOR U5799 ( .A(n3944), .B(n3943), .Z(n3945) );
  XNOR U5800 ( .A(n3946), .B(n3945), .Z(out[75]) );
  XOR U5801 ( .A(in[368]), .B(n3947), .Z(n4319) );
  NOR U5802 ( .A(n4160), .B(n4594), .Z(n3948) );
  XNOR U5803 ( .A(n4319), .B(n3948), .Z(out[760]) );
  XOR U5804 ( .A(in[369]), .B(n3949), .Z(n4321) );
  NOR U5805 ( .A(n4163), .B(n4598), .Z(n3950) );
  XNOR U5806 ( .A(n4321), .B(n3950), .Z(out[761]) );
  XOR U5807 ( .A(in[370]), .B(n3951), .Z(n4327) );
  NOR U5808 ( .A(n4166), .B(n4602), .Z(n3952) );
  XNOR U5809 ( .A(n4327), .B(n3952), .Z(out[762]) );
  XOR U5810 ( .A(in[371]), .B(n3953), .Z(n4329) );
  NOR U5811 ( .A(n4169), .B(n4606), .Z(n3954) );
  XNOR U5812 ( .A(n4329), .B(n3954), .Z(out[763]) );
  XOR U5813 ( .A(in[372]), .B(n3955), .Z(n4331) );
  NOR U5814 ( .A(n4172), .B(n4610), .Z(n3956) );
  XNOR U5815 ( .A(n4331), .B(n3956), .Z(out[764]) );
  XOR U5816 ( .A(in[373]), .B(n3957), .Z(n4333) );
  NOR U5817 ( .A(n4175), .B(n4614), .Z(n3958) );
  XNOR U5818 ( .A(n4333), .B(n3958), .Z(out[765]) );
  XOR U5819 ( .A(in[374]), .B(n3959), .Z(n4335) );
  NOR U5820 ( .A(n4182), .B(n4618), .Z(n3960) );
  XNOR U5821 ( .A(n4335), .B(n3960), .Z(out[766]) );
  XOR U5822 ( .A(in[375]), .B(n3961), .Z(n4337) );
  NOR U5823 ( .A(n4185), .B(n4622), .Z(n3962) );
  XNOR U5824 ( .A(n4337), .B(n3962), .Z(out[767]) );
  XNOR U5825 ( .A(in[743]), .B(n3963), .Z(n4340) );
  NAND U5826 ( .A(n4187), .B(n3964), .Z(n3965) );
  XNOR U5827 ( .A(n4340), .B(n3965), .Z(out[768]) );
  XNOR U5828 ( .A(in[744]), .B(n3966), .Z(n4344) );
  NAND U5829 ( .A(n4189), .B(n3967), .Z(n3968) );
  XNOR U5830 ( .A(n4344), .B(n3968), .Z(out[769]) );
  NOR U5831 ( .A(n3970), .B(n3969), .Z(n3971) );
  XNOR U5832 ( .A(n3972), .B(n3971), .Z(out[76]) );
  XNOR U5833 ( .A(in[745]), .B(n3973), .Z(n4348) );
  NAND U5834 ( .A(n4191), .B(n3974), .Z(n3975) );
  XNOR U5835 ( .A(n4348), .B(n3975), .Z(out[770]) );
  XNOR U5836 ( .A(in[746]), .B(n3976), .Z(n4352) );
  NAND U5837 ( .A(n4193), .B(n3977), .Z(n3978) );
  XNOR U5838 ( .A(n4352), .B(n3978), .Z(out[771]) );
  XNOR U5839 ( .A(in[747]), .B(n3979), .Z(n4364) );
  NAND U5840 ( .A(n4195), .B(n3980), .Z(n3981) );
  XNOR U5841 ( .A(n4364), .B(n3981), .Z(out[772]) );
  XNOR U5842 ( .A(in[748]), .B(n3982), .Z(n4368) );
  NAND U5843 ( .A(n4197), .B(n3983), .Z(n3984) );
  XNOR U5844 ( .A(n4368), .B(n3984), .Z(out[773]) );
  XNOR U5845 ( .A(in[749]), .B(n3985), .Z(n4372) );
  NAND U5846 ( .A(n4199), .B(n3986), .Z(n3987) );
  XNOR U5847 ( .A(n4372), .B(n3987), .Z(out[774]) );
  XNOR U5848 ( .A(in[750]), .B(n3988), .Z(n4376) );
  NAND U5849 ( .A(n4201), .B(n3989), .Z(n3990) );
  XNOR U5850 ( .A(n4376), .B(n3990), .Z(out[775]) );
  XNOR U5851 ( .A(in[751]), .B(n3991), .Z(n4380) );
  NAND U5852 ( .A(n4207), .B(n3992), .Z(n3993) );
  XNOR U5853 ( .A(n4380), .B(n3993), .Z(out[776]) );
  XNOR U5854 ( .A(in[752]), .B(n3994), .Z(n4384) );
  NAND U5855 ( .A(n4209), .B(n3995), .Z(n3996) );
  XNOR U5856 ( .A(n4384), .B(n3996), .Z(out[777]) );
  XNOR U5857 ( .A(in[753]), .B(n3997), .Z(n4388) );
  NAND U5858 ( .A(n4211), .B(n3998), .Z(n3999) );
  XNOR U5859 ( .A(n4388), .B(n3999), .Z(out[778]) );
  XNOR U5860 ( .A(in[754]), .B(n4000), .Z(n4392) );
  NAND U5861 ( .A(n4213), .B(n4001), .Z(n4002) );
  XNOR U5862 ( .A(n4392), .B(n4002), .Z(out[779]) );
  NOR U5863 ( .A(n4004), .B(n4003), .Z(n4005) );
  XNOR U5864 ( .A(n4006), .B(n4005), .Z(out[77]) );
  XNOR U5865 ( .A(in[755]), .B(n4007), .Z(n4396) );
  NAND U5866 ( .A(n4215), .B(n4008), .Z(n4009) );
  XNOR U5867 ( .A(n4396), .B(n4009), .Z(out[780]) );
  XNOR U5868 ( .A(in[756]), .B(n4010), .Z(n4400) );
  NAND U5869 ( .A(n4217), .B(n4011), .Z(n4012) );
  XNOR U5870 ( .A(n4400), .B(n4012), .Z(out[781]) );
  XNOR U5871 ( .A(in[757]), .B(n4013), .Z(n4408) );
  NAND U5872 ( .A(n4219), .B(n4014), .Z(n4015) );
  XNOR U5873 ( .A(n4408), .B(n4015), .Z(out[782]) );
  XNOR U5874 ( .A(in[758]), .B(n4016), .Z(n4412) );
  NAND U5875 ( .A(n4221), .B(n4017), .Z(n4018) );
  XNOR U5876 ( .A(n4412), .B(n4018), .Z(out[783]) );
  XNOR U5877 ( .A(in[759]), .B(n4019), .Z(n4416) );
  NAND U5878 ( .A(n4223), .B(n4020), .Z(n4021) );
  XNOR U5879 ( .A(n4416), .B(n4021), .Z(out[784]) );
  XNOR U5880 ( .A(in[760]), .B(n4022), .Z(n4420) );
  NAND U5881 ( .A(n4225), .B(n4023), .Z(n4024) );
  XNOR U5882 ( .A(n4420), .B(n4024), .Z(out[785]) );
  XNOR U5883 ( .A(in[761]), .B(n4025), .Z(n4424) );
  NAND U5884 ( .A(n4231), .B(n4026), .Z(n4027) );
  XNOR U5885 ( .A(n4424), .B(n4027), .Z(out[786]) );
  XNOR U5886 ( .A(in[762]), .B(n4028), .Z(n4428) );
  NAND U5887 ( .A(n4233), .B(n4029), .Z(n4030) );
  XNOR U5888 ( .A(n4428), .B(n4030), .Z(out[787]) );
  XNOR U5889 ( .A(in[763]), .B(n4031), .Z(n4432) );
  NAND U5890 ( .A(n4235), .B(n4032), .Z(n4033) );
  XNOR U5891 ( .A(n4432), .B(n4033), .Z(out[788]) );
  XNOR U5892 ( .A(in[764]), .B(n4034), .Z(n4436) );
  NAND U5893 ( .A(n4237), .B(n4035), .Z(n4036) );
  XNOR U5894 ( .A(n4436), .B(n4036), .Z(out[789]) );
  NOR U5895 ( .A(n4038), .B(n4037), .Z(n4039) );
  XNOR U5896 ( .A(n4040), .B(n4039), .Z(out[78]) );
  XNOR U5897 ( .A(in[765]), .B(n4041), .Z(n4440) );
  NAND U5898 ( .A(n4239), .B(n4042), .Z(n4043) );
  XNOR U5899 ( .A(n4440), .B(n4043), .Z(out[790]) );
  XNOR U5900 ( .A(in[766]), .B(n4044), .Z(n4444) );
  NAND U5901 ( .A(n4241), .B(n4045), .Z(n4046) );
  XNOR U5902 ( .A(n4444), .B(n4046), .Z(out[791]) );
  XNOR U5903 ( .A(in[767]), .B(n4047), .Z(n4452) );
  NAND U5904 ( .A(n4243), .B(n4048), .Z(n4049) );
  XNOR U5905 ( .A(n4452), .B(n4049), .Z(out[792]) );
  XNOR U5906 ( .A(in[704]), .B(n4050), .Z(n4456) );
  NAND U5907 ( .A(n4245), .B(n4051), .Z(n4052) );
  XNOR U5908 ( .A(n4456), .B(n4052), .Z(out[793]) );
  XNOR U5909 ( .A(in[705]), .B(n4053), .Z(n4460) );
  NAND U5910 ( .A(n4247), .B(n4054), .Z(n4055) );
  XNOR U5911 ( .A(n4460), .B(n4055), .Z(out[794]) );
  XNOR U5912 ( .A(in[706]), .B(n4056), .Z(n4464) );
  NAND U5913 ( .A(n4249), .B(n4057), .Z(n4058) );
  XNOR U5914 ( .A(n4464), .B(n4058), .Z(out[795]) );
  XNOR U5915 ( .A(in[707]), .B(n4059), .Z(n4468) );
  NAND U5916 ( .A(n4255), .B(n4060), .Z(n4061) );
  XNOR U5917 ( .A(n4468), .B(n4061), .Z(out[796]) );
  XNOR U5918 ( .A(in[708]), .B(n4062), .Z(n4472) );
  NAND U5919 ( .A(n4257), .B(n4063), .Z(n4064) );
  XNOR U5920 ( .A(n4472), .B(n4064), .Z(out[797]) );
  XNOR U5921 ( .A(in[709]), .B(n4065), .Z(n4476) );
  NAND U5922 ( .A(n4259), .B(n4066), .Z(n4067) );
  XNOR U5923 ( .A(n4476), .B(n4067), .Z(out[798]) );
  XNOR U5924 ( .A(in[710]), .B(n4068), .Z(n4480) );
  NAND U5925 ( .A(n4261), .B(n4069), .Z(n4070) );
  XNOR U5926 ( .A(n4480), .B(n4070), .Z(out[799]) );
  NOR U5927 ( .A(n4072), .B(n4071), .Z(n4073) );
  XNOR U5928 ( .A(n4074), .B(n4073), .Z(out[79]) );
  OR U5929 ( .A(n4076), .B(n4075), .Z(n4077) );
  XNOR U5930 ( .A(n4078), .B(n4077), .Z(out[7]) );
  XNOR U5931 ( .A(in[711]), .B(n4079), .Z(n4484) );
  NAND U5932 ( .A(n4263), .B(n4080), .Z(n4081) );
  XNOR U5933 ( .A(n4484), .B(n4081), .Z(out[800]) );
  XNOR U5934 ( .A(in[712]), .B(n4082), .Z(n4488) );
  NAND U5935 ( .A(n4265), .B(n4083), .Z(n4084) );
  XNOR U5936 ( .A(n4488), .B(n4084), .Z(out[801]) );
  XNOR U5937 ( .A(in[713]), .B(n4085), .Z(n4496) );
  NAND U5938 ( .A(n4267), .B(n4086), .Z(n4087) );
  XNOR U5939 ( .A(n4496), .B(n4087), .Z(out[802]) );
  XNOR U5940 ( .A(in[714]), .B(n4088), .Z(n4500) );
  NAND U5941 ( .A(n4269), .B(n4089), .Z(n4090) );
  XNOR U5942 ( .A(n4500), .B(n4090), .Z(out[803]) );
  XNOR U5943 ( .A(in[715]), .B(n4091), .Z(n4504) );
  NAND U5944 ( .A(n4271), .B(n4092), .Z(n4093) );
  XNOR U5945 ( .A(n4504), .B(n4093), .Z(out[804]) );
  XOR U5946 ( .A(n4094), .B(in[716]), .Z(n4508) );
  NAND U5947 ( .A(n4273), .B(n4095), .Z(n4096) );
  XNOR U5948 ( .A(n4508), .B(n4096), .Z(out[805]) );
  XOR U5949 ( .A(n4097), .B(in[717]), .Z(n4512) );
  NAND U5950 ( .A(n4279), .B(n4098), .Z(n4099) );
  XNOR U5951 ( .A(n4512), .B(n4099), .Z(out[806]) );
  XOR U5952 ( .A(n4100), .B(in[718]), .Z(n4516) );
  NAND U5953 ( .A(n4281), .B(n4101), .Z(n4102) );
  XNOR U5954 ( .A(n4516), .B(n4102), .Z(out[807]) );
  XOR U5955 ( .A(n4103), .B(in[719]), .Z(n4520) );
  NAND U5956 ( .A(n4283), .B(n4104), .Z(n4105) );
  XNOR U5957 ( .A(n4520), .B(n4105), .Z(out[808]) );
  XOR U5958 ( .A(n4106), .B(in[720]), .Z(n4524) );
  NAND U5959 ( .A(n4285), .B(n4107), .Z(n4108) );
  XNOR U5960 ( .A(n4524), .B(n4108), .Z(out[809]) );
  NOR U5961 ( .A(n4110), .B(n4109), .Z(n4111) );
  XNOR U5962 ( .A(n4112), .B(n4111), .Z(out[80]) );
  XOR U5963 ( .A(n4113), .B(in[721]), .Z(n4528) );
  NAND U5964 ( .A(n4287), .B(n4114), .Z(n4115) );
  XNOR U5965 ( .A(n4528), .B(n4115), .Z(out[810]) );
  XOR U5966 ( .A(n4116), .B(in[722]), .Z(n4532) );
  NAND U5967 ( .A(n4289), .B(n4117), .Z(n4118) );
  XNOR U5968 ( .A(n4532), .B(n4118), .Z(out[811]) );
  XOR U5969 ( .A(n4119), .B(in[723]), .Z(n4540) );
  NAND U5970 ( .A(n4291), .B(n4120), .Z(n4121) );
  XNOR U5971 ( .A(n4540), .B(n4121), .Z(out[812]) );
  XOR U5972 ( .A(in[724]), .B(n4122), .Z(n4544) );
  NAND U5973 ( .A(n4293), .B(n4123), .Z(n4124) );
  XNOR U5974 ( .A(n4544), .B(n4124), .Z(out[813]) );
  XOR U5975 ( .A(in[725]), .B(n4125), .Z(n4548) );
  NAND U5976 ( .A(n4295), .B(n4126), .Z(n4127) );
  XNOR U5977 ( .A(n4548), .B(n4127), .Z(out[814]) );
  XOR U5978 ( .A(in[726]), .B(n4128), .Z(n4552) );
  NAND U5979 ( .A(n4297), .B(n4129), .Z(n4130) );
  XNOR U5980 ( .A(n4552), .B(n4130), .Z(out[815]) );
  XOR U5981 ( .A(in[727]), .B(n4131), .Z(n4556) );
  NAND U5982 ( .A(n4303), .B(n4132), .Z(n4133) );
  XNOR U5983 ( .A(n4556), .B(n4133), .Z(out[816]) );
  XOR U5984 ( .A(in[728]), .B(n4134), .Z(n4560) );
  NAND U5985 ( .A(n4305), .B(n4135), .Z(n4136) );
  XNOR U5986 ( .A(n4560), .B(n4136), .Z(out[817]) );
  XOR U5987 ( .A(in[729]), .B(n4137), .Z(n4564) );
  NAND U5988 ( .A(n4307), .B(n4138), .Z(n4139) );
  XNOR U5989 ( .A(n4564), .B(n4139), .Z(out[818]) );
  XOR U5990 ( .A(in[730]), .B(n4140), .Z(n4568) );
  NAND U5991 ( .A(n4309), .B(n4141), .Z(n4142) );
  XNOR U5992 ( .A(n4568), .B(n4142), .Z(out[819]) );
  NOR U5993 ( .A(n4144), .B(n4143), .Z(n4145) );
  XNOR U5994 ( .A(n4146), .B(n4145), .Z(out[81]) );
  XOR U5995 ( .A(in[731]), .B(n4147), .Z(n4572) );
  NAND U5996 ( .A(n4311), .B(n4148), .Z(n4149) );
  XNOR U5997 ( .A(n4572), .B(n4149), .Z(out[820]) );
  XOR U5998 ( .A(in[732]), .B(n4150), .Z(n4576) );
  NAND U5999 ( .A(n4313), .B(n4151), .Z(n4152) );
  XNOR U6000 ( .A(n4576), .B(n4152), .Z(out[821]) );
  XOR U6001 ( .A(in[733]), .B(n4153), .Z(n4584) );
  NAND U6002 ( .A(n4315), .B(n4154), .Z(n4155) );
  XNOR U6003 ( .A(n4584), .B(n4155), .Z(out[822]) );
  XOR U6004 ( .A(in[734]), .B(n4156), .Z(n4588) );
  NAND U6005 ( .A(n4317), .B(n4157), .Z(n4158) );
  XNOR U6006 ( .A(n4588), .B(n4158), .Z(out[823]) );
  XOR U6007 ( .A(in[735]), .B(n4159), .Z(n4592) );
  NAND U6008 ( .A(n4319), .B(n4160), .Z(n4161) );
  XNOR U6009 ( .A(n4592), .B(n4161), .Z(out[824]) );
  XOR U6010 ( .A(in[736]), .B(n4162), .Z(n4596) );
  NAND U6011 ( .A(n4321), .B(n4163), .Z(n4164) );
  XNOR U6012 ( .A(n4596), .B(n4164), .Z(out[825]) );
  XOR U6013 ( .A(in[737]), .B(n4165), .Z(n4600) );
  NAND U6014 ( .A(n4327), .B(n4166), .Z(n4167) );
  XNOR U6015 ( .A(n4600), .B(n4167), .Z(out[826]) );
  XOR U6016 ( .A(in[738]), .B(n4168), .Z(n4604) );
  NAND U6017 ( .A(n4329), .B(n4169), .Z(n4170) );
  XNOR U6018 ( .A(n4604), .B(n4170), .Z(out[827]) );
  XOR U6019 ( .A(in[739]), .B(n4171), .Z(n4608) );
  NAND U6020 ( .A(n4331), .B(n4172), .Z(n4173) );
  XNOR U6021 ( .A(n4608), .B(n4173), .Z(out[828]) );
  XNOR U6022 ( .A(in[740]), .B(n4174), .Z(n4612) );
  NAND U6023 ( .A(n4333), .B(n4175), .Z(n4176) );
  XNOR U6024 ( .A(n4612), .B(n4176), .Z(out[829]) );
  NOR U6025 ( .A(n4178), .B(n4177), .Z(n4179) );
  XNOR U6026 ( .A(n4180), .B(n4179), .Z(out[82]) );
  XNOR U6027 ( .A(in[741]), .B(n4181), .Z(n4616) );
  NAND U6028 ( .A(n4335), .B(n4182), .Z(n4183) );
  XNOR U6029 ( .A(n4616), .B(n4183), .Z(out[830]) );
  XNOR U6030 ( .A(in[742]), .B(n4184), .Z(n4620) );
  NAND U6031 ( .A(n4337), .B(n4185), .Z(n4186) );
  XNOR U6032 ( .A(n4620), .B(n4186), .Z(out[831]) );
  OR U6033 ( .A(n4340), .B(n4187), .Z(n4188) );
  XNOR U6034 ( .A(n4339), .B(n4188), .Z(out[832]) );
  OR U6035 ( .A(n4344), .B(n4189), .Z(n4190) );
  XNOR U6036 ( .A(n4343), .B(n4190), .Z(out[833]) );
  OR U6037 ( .A(n4348), .B(n4191), .Z(n4192) );
  XNOR U6038 ( .A(n4347), .B(n4192), .Z(out[834]) );
  OR U6039 ( .A(n4352), .B(n4193), .Z(n4194) );
  XNOR U6040 ( .A(n4351), .B(n4194), .Z(out[835]) );
  OR U6041 ( .A(n4364), .B(n4195), .Z(n4196) );
  XNOR U6042 ( .A(n4363), .B(n4196), .Z(out[836]) );
  OR U6043 ( .A(n4368), .B(n4197), .Z(n4198) );
  XNOR U6044 ( .A(n4367), .B(n4198), .Z(out[837]) );
  OR U6045 ( .A(n4372), .B(n4199), .Z(n4200) );
  XNOR U6046 ( .A(n4371), .B(n4200), .Z(out[838]) );
  OR U6047 ( .A(n4376), .B(n4201), .Z(n4202) );
  XNOR U6048 ( .A(n4375), .B(n4202), .Z(out[839]) );
  NOR U6049 ( .A(n4204), .B(n4203), .Z(n4205) );
  XNOR U6050 ( .A(n4206), .B(n4205), .Z(out[83]) );
  OR U6051 ( .A(n4380), .B(n4207), .Z(n4208) );
  XNOR U6052 ( .A(n4379), .B(n4208), .Z(out[840]) );
  OR U6053 ( .A(n4384), .B(n4209), .Z(n4210) );
  XNOR U6054 ( .A(n4383), .B(n4210), .Z(out[841]) );
  OR U6055 ( .A(n4388), .B(n4211), .Z(n4212) );
  XNOR U6056 ( .A(n4387), .B(n4212), .Z(out[842]) );
  OR U6057 ( .A(n4392), .B(n4213), .Z(n4214) );
  XNOR U6058 ( .A(n4391), .B(n4214), .Z(out[843]) );
  OR U6059 ( .A(n4396), .B(n4215), .Z(n4216) );
  XNOR U6060 ( .A(n4395), .B(n4216), .Z(out[844]) );
  OR U6061 ( .A(n4400), .B(n4217), .Z(n4218) );
  XNOR U6062 ( .A(n4399), .B(n4218), .Z(out[845]) );
  OR U6063 ( .A(n4408), .B(n4219), .Z(n4220) );
  XNOR U6064 ( .A(n4407), .B(n4220), .Z(out[846]) );
  OR U6065 ( .A(n4412), .B(n4221), .Z(n4222) );
  XNOR U6066 ( .A(n4411), .B(n4222), .Z(out[847]) );
  OR U6067 ( .A(n4416), .B(n4223), .Z(n4224) );
  XNOR U6068 ( .A(n4415), .B(n4224), .Z(out[848]) );
  OR U6069 ( .A(n4420), .B(n4225), .Z(n4226) );
  XNOR U6070 ( .A(n4419), .B(n4226), .Z(out[849]) );
  NOR U6071 ( .A(n4228), .B(n4227), .Z(n4229) );
  XNOR U6072 ( .A(n4230), .B(n4229), .Z(out[84]) );
  OR U6073 ( .A(n4424), .B(n4231), .Z(n4232) );
  XNOR U6074 ( .A(n4423), .B(n4232), .Z(out[850]) );
  OR U6075 ( .A(n4428), .B(n4233), .Z(n4234) );
  XNOR U6076 ( .A(n4427), .B(n4234), .Z(out[851]) );
  OR U6077 ( .A(n4432), .B(n4235), .Z(n4236) );
  XNOR U6078 ( .A(n4431), .B(n4236), .Z(out[852]) );
  OR U6079 ( .A(n4436), .B(n4237), .Z(n4238) );
  XNOR U6080 ( .A(n4435), .B(n4238), .Z(out[853]) );
  OR U6081 ( .A(n4440), .B(n4239), .Z(n4240) );
  XNOR U6082 ( .A(n4439), .B(n4240), .Z(out[854]) );
  OR U6083 ( .A(n4444), .B(n4241), .Z(n4242) );
  XNOR U6084 ( .A(n4443), .B(n4242), .Z(out[855]) );
  OR U6085 ( .A(n4452), .B(n4243), .Z(n4244) );
  XNOR U6086 ( .A(n4451), .B(n4244), .Z(out[856]) );
  OR U6087 ( .A(n4456), .B(n4245), .Z(n4246) );
  XNOR U6088 ( .A(n4455), .B(n4246), .Z(out[857]) );
  OR U6089 ( .A(n4460), .B(n4247), .Z(n4248) );
  XNOR U6090 ( .A(n4459), .B(n4248), .Z(out[858]) );
  OR U6091 ( .A(n4464), .B(n4249), .Z(n4250) );
  XNOR U6092 ( .A(n4463), .B(n4250), .Z(out[859]) );
  NOR U6093 ( .A(n4252), .B(n4251), .Z(n4253) );
  XNOR U6094 ( .A(n4254), .B(n4253), .Z(out[85]) );
  OR U6095 ( .A(n4468), .B(n4255), .Z(n4256) );
  XNOR U6096 ( .A(n4467), .B(n4256), .Z(out[860]) );
  OR U6097 ( .A(n4472), .B(n4257), .Z(n4258) );
  XNOR U6098 ( .A(n4471), .B(n4258), .Z(out[861]) );
  OR U6099 ( .A(n4476), .B(n4259), .Z(n4260) );
  XNOR U6100 ( .A(n4475), .B(n4260), .Z(out[862]) );
  OR U6101 ( .A(n4480), .B(n4261), .Z(n4262) );
  XNOR U6102 ( .A(n4479), .B(n4262), .Z(out[863]) );
  OR U6103 ( .A(n4484), .B(n4263), .Z(n4264) );
  XNOR U6104 ( .A(n4483), .B(n4264), .Z(out[864]) );
  OR U6105 ( .A(n4488), .B(n4265), .Z(n4266) );
  XNOR U6106 ( .A(n4487), .B(n4266), .Z(out[865]) );
  OR U6107 ( .A(n4496), .B(n4267), .Z(n4268) );
  XNOR U6108 ( .A(n4495), .B(n4268), .Z(out[866]) );
  OR U6109 ( .A(n4500), .B(n4269), .Z(n4270) );
  XNOR U6110 ( .A(n4499), .B(n4270), .Z(out[867]) );
  OR U6111 ( .A(n4504), .B(n4271), .Z(n4272) );
  XNOR U6112 ( .A(n4503), .B(n4272), .Z(out[868]) );
  OR U6113 ( .A(n4508), .B(n4273), .Z(n4274) );
  XNOR U6114 ( .A(n4507), .B(n4274), .Z(out[869]) );
  NOR U6115 ( .A(n4276), .B(n4275), .Z(n4277) );
  XNOR U6116 ( .A(n4278), .B(n4277), .Z(out[86]) );
  OR U6117 ( .A(n4512), .B(n4279), .Z(n4280) );
  XNOR U6118 ( .A(n4511), .B(n4280), .Z(out[870]) );
  OR U6119 ( .A(n4516), .B(n4281), .Z(n4282) );
  XNOR U6120 ( .A(n4515), .B(n4282), .Z(out[871]) );
  OR U6121 ( .A(n4520), .B(n4283), .Z(n4284) );
  XNOR U6122 ( .A(n4519), .B(n4284), .Z(out[872]) );
  OR U6123 ( .A(n4524), .B(n4285), .Z(n4286) );
  XNOR U6124 ( .A(n4523), .B(n4286), .Z(out[873]) );
  OR U6125 ( .A(n4528), .B(n4287), .Z(n4288) );
  XNOR U6126 ( .A(n4527), .B(n4288), .Z(out[874]) );
  OR U6127 ( .A(n4532), .B(n4289), .Z(n4290) );
  XNOR U6128 ( .A(n4531), .B(n4290), .Z(out[875]) );
  OR U6129 ( .A(n4540), .B(n4291), .Z(n4292) );
  XNOR U6130 ( .A(n4539), .B(n4292), .Z(out[876]) );
  OR U6131 ( .A(n4544), .B(n4293), .Z(n4294) );
  XNOR U6132 ( .A(n4543), .B(n4294), .Z(out[877]) );
  OR U6133 ( .A(n4548), .B(n4295), .Z(n4296) );
  XNOR U6134 ( .A(n4547), .B(n4296), .Z(out[878]) );
  OR U6135 ( .A(n4552), .B(n4297), .Z(n4298) );
  XNOR U6136 ( .A(n4551), .B(n4298), .Z(out[879]) );
  NOR U6137 ( .A(n4300), .B(n4299), .Z(n4301) );
  XNOR U6138 ( .A(n4302), .B(n4301), .Z(out[87]) );
  OR U6139 ( .A(n4556), .B(n4303), .Z(n4304) );
  XNOR U6140 ( .A(n4555), .B(n4304), .Z(out[880]) );
  OR U6141 ( .A(n4560), .B(n4305), .Z(n4306) );
  XNOR U6142 ( .A(n4559), .B(n4306), .Z(out[881]) );
  OR U6143 ( .A(n4564), .B(n4307), .Z(n4308) );
  XNOR U6144 ( .A(n4563), .B(n4308), .Z(out[882]) );
  OR U6145 ( .A(n4568), .B(n4309), .Z(n4310) );
  XNOR U6146 ( .A(n4567), .B(n4310), .Z(out[883]) );
  OR U6147 ( .A(n4572), .B(n4311), .Z(n4312) );
  XNOR U6148 ( .A(n4571), .B(n4312), .Z(out[884]) );
  OR U6149 ( .A(n4576), .B(n4313), .Z(n4314) );
  XNOR U6150 ( .A(n4575), .B(n4314), .Z(out[885]) );
  OR U6151 ( .A(n4584), .B(n4315), .Z(n4316) );
  XNOR U6152 ( .A(n4583), .B(n4316), .Z(out[886]) );
  OR U6153 ( .A(n4588), .B(n4317), .Z(n4318) );
  XNOR U6154 ( .A(n4587), .B(n4318), .Z(out[887]) );
  OR U6155 ( .A(n4592), .B(n4319), .Z(n4320) );
  XNOR U6156 ( .A(n4591), .B(n4320), .Z(out[888]) );
  OR U6157 ( .A(n4596), .B(n4321), .Z(n4322) );
  XNOR U6158 ( .A(n4595), .B(n4322), .Z(out[889]) );
  NOR U6159 ( .A(n4324), .B(n4323), .Z(n4325) );
  XNOR U6160 ( .A(n4326), .B(n4325), .Z(out[88]) );
  OR U6161 ( .A(n4600), .B(n4327), .Z(n4328) );
  XNOR U6162 ( .A(n4599), .B(n4328), .Z(out[890]) );
  OR U6163 ( .A(n4604), .B(n4329), .Z(n4330) );
  XNOR U6164 ( .A(n4603), .B(n4330), .Z(out[891]) );
  OR U6165 ( .A(n4608), .B(n4331), .Z(n4332) );
  XNOR U6166 ( .A(n4607), .B(n4332), .Z(out[892]) );
  OR U6167 ( .A(n4612), .B(n4333), .Z(n4334) );
  XNOR U6168 ( .A(n4611), .B(n4334), .Z(out[893]) );
  OR U6169 ( .A(n4616), .B(n4335), .Z(n4336) );
  XNOR U6170 ( .A(n4615), .B(n4336), .Z(out[894]) );
  OR U6171 ( .A(n4620), .B(n4337), .Z(n4338) );
  XNOR U6172 ( .A(n4619), .B(n4338), .Z(out[895]) );
  ANDN U6173 ( .B(n4340), .A(n4339), .Z(n4341) );
  XNOR U6174 ( .A(n4342), .B(n4341), .Z(out[896]) );
  ANDN U6175 ( .B(n4344), .A(n4343), .Z(n4345) );
  XNOR U6176 ( .A(n4346), .B(n4345), .Z(out[897]) );
  ANDN U6177 ( .B(n4348), .A(n4347), .Z(n4349) );
  XNOR U6178 ( .A(n4350), .B(n4349), .Z(out[898]) );
  ANDN U6179 ( .B(n4352), .A(n4351), .Z(n4353) );
  XNOR U6180 ( .A(n4354), .B(n4353), .Z(out[899]) );
  NOR U6181 ( .A(n4356), .B(n4355), .Z(n4357) );
  XNOR U6182 ( .A(n4358), .B(n4357), .Z(out[89]) );
  OR U6183 ( .A(n4360), .B(n4359), .Z(n4361) );
  XNOR U6184 ( .A(n4362), .B(n4361), .Z(out[8]) );
  ANDN U6185 ( .B(n4364), .A(n4363), .Z(n4365) );
  XNOR U6186 ( .A(n4366), .B(n4365), .Z(out[900]) );
  ANDN U6187 ( .B(n4368), .A(n4367), .Z(n4369) );
  XNOR U6188 ( .A(n4370), .B(n4369), .Z(out[901]) );
  ANDN U6189 ( .B(n4372), .A(n4371), .Z(n4373) );
  XNOR U6190 ( .A(n4374), .B(n4373), .Z(out[902]) );
  ANDN U6191 ( .B(n4376), .A(n4375), .Z(n4377) );
  XNOR U6192 ( .A(n4378), .B(n4377), .Z(out[903]) );
  ANDN U6193 ( .B(n4380), .A(n4379), .Z(n4381) );
  XNOR U6194 ( .A(n4382), .B(n4381), .Z(out[904]) );
  ANDN U6195 ( .B(n4384), .A(n4383), .Z(n4385) );
  XNOR U6196 ( .A(n4386), .B(n4385), .Z(out[905]) );
  ANDN U6197 ( .B(n4388), .A(n4387), .Z(n4389) );
  XNOR U6198 ( .A(n4390), .B(n4389), .Z(out[906]) );
  ANDN U6199 ( .B(n4392), .A(n4391), .Z(n4393) );
  XNOR U6200 ( .A(n4394), .B(n4393), .Z(out[907]) );
  ANDN U6201 ( .B(n4396), .A(n4395), .Z(n4397) );
  XNOR U6202 ( .A(n4398), .B(n4397), .Z(out[908]) );
  ANDN U6203 ( .B(n4400), .A(n4399), .Z(n4401) );
  XNOR U6204 ( .A(n4402), .B(n4401), .Z(out[909]) );
  NOR U6205 ( .A(n4404), .B(n4403), .Z(n4405) );
  XNOR U6206 ( .A(n4406), .B(n4405), .Z(out[90]) );
  ANDN U6207 ( .B(n4408), .A(n4407), .Z(n4409) );
  XNOR U6208 ( .A(n4410), .B(n4409), .Z(out[910]) );
  ANDN U6209 ( .B(n4412), .A(n4411), .Z(n4413) );
  XNOR U6210 ( .A(n4414), .B(n4413), .Z(out[911]) );
  ANDN U6211 ( .B(n4416), .A(n4415), .Z(n4417) );
  XNOR U6212 ( .A(n4418), .B(n4417), .Z(out[912]) );
  ANDN U6213 ( .B(n4420), .A(n4419), .Z(n4421) );
  XNOR U6214 ( .A(n4422), .B(n4421), .Z(out[913]) );
  ANDN U6215 ( .B(n4424), .A(n4423), .Z(n4425) );
  XNOR U6216 ( .A(n4426), .B(n4425), .Z(out[914]) );
  ANDN U6217 ( .B(n4428), .A(n4427), .Z(n4429) );
  XNOR U6218 ( .A(n4430), .B(n4429), .Z(out[915]) );
  ANDN U6219 ( .B(n4432), .A(n4431), .Z(n4433) );
  XNOR U6220 ( .A(n4434), .B(n4433), .Z(out[916]) );
  ANDN U6221 ( .B(n4436), .A(n4435), .Z(n4437) );
  XNOR U6222 ( .A(n4438), .B(n4437), .Z(out[917]) );
  ANDN U6223 ( .B(n4440), .A(n4439), .Z(n4441) );
  XNOR U6224 ( .A(n4442), .B(n4441), .Z(out[918]) );
  ANDN U6225 ( .B(n4444), .A(n4443), .Z(n4445) );
  XNOR U6226 ( .A(n4446), .B(n4445), .Z(out[919]) );
  NOR U6227 ( .A(n4448), .B(n4447), .Z(n4449) );
  XNOR U6228 ( .A(n4450), .B(n4449), .Z(out[91]) );
  ANDN U6229 ( .B(n4452), .A(n4451), .Z(n4453) );
  XNOR U6230 ( .A(n4454), .B(n4453), .Z(out[920]) );
  ANDN U6231 ( .B(n4456), .A(n4455), .Z(n4457) );
  XNOR U6232 ( .A(n4458), .B(n4457), .Z(out[921]) );
  ANDN U6233 ( .B(n4460), .A(n4459), .Z(n4461) );
  XNOR U6234 ( .A(n4462), .B(n4461), .Z(out[922]) );
  ANDN U6235 ( .B(n4464), .A(n4463), .Z(n4465) );
  XNOR U6236 ( .A(n4466), .B(n4465), .Z(out[923]) );
  ANDN U6237 ( .B(n4468), .A(n4467), .Z(n4469) );
  XNOR U6238 ( .A(n4470), .B(n4469), .Z(out[924]) );
  ANDN U6239 ( .B(n4472), .A(n4471), .Z(n4473) );
  XNOR U6240 ( .A(n4474), .B(n4473), .Z(out[925]) );
  ANDN U6241 ( .B(n4476), .A(n4475), .Z(n4477) );
  XNOR U6242 ( .A(n4478), .B(n4477), .Z(out[926]) );
  ANDN U6243 ( .B(n4480), .A(n4479), .Z(n4481) );
  XNOR U6244 ( .A(n4482), .B(n4481), .Z(out[927]) );
  ANDN U6245 ( .B(n4484), .A(n4483), .Z(n4485) );
  XNOR U6246 ( .A(n4486), .B(n4485), .Z(out[928]) );
  ANDN U6247 ( .B(n4488), .A(n4487), .Z(n4489) );
  XNOR U6248 ( .A(n4490), .B(n4489), .Z(out[929]) );
  ANDN U6249 ( .B(n4492), .A(n4491), .Z(n4493) );
  XNOR U6250 ( .A(n4494), .B(n4493), .Z(out[92]) );
  ANDN U6251 ( .B(n4496), .A(n4495), .Z(n4497) );
  XNOR U6252 ( .A(n4498), .B(n4497), .Z(out[930]) );
  ANDN U6253 ( .B(n4500), .A(n4499), .Z(n4501) );
  XNOR U6254 ( .A(n4502), .B(n4501), .Z(out[931]) );
  ANDN U6255 ( .B(n4504), .A(n4503), .Z(n4505) );
  XNOR U6256 ( .A(n4506), .B(n4505), .Z(out[932]) );
  ANDN U6257 ( .B(n4508), .A(n4507), .Z(n4509) );
  XNOR U6258 ( .A(n4510), .B(n4509), .Z(out[933]) );
  ANDN U6259 ( .B(n4512), .A(n4511), .Z(n4513) );
  XNOR U6260 ( .A(n4514), .B(n4513), .Z(out[934]) );
  ANDN U6261 ( .B(n4516), .A(n4515), .Z(n4517) );
  XNOR U6262 ( .A(n4518), .B(n4517), .Z(out[935]) );
  ANDN U6263 ( .B(n4520), .A(n4519), .Z(n4521) );
  XNOR U6264 ( .A(n4522), .B(n4521), .Z(out[936]) );
  ANDN U6265 ( .B(n4524), .A(n4523), .Z(n4525) );
  XNOR U6266 ( .A(n4526), .B(n4525), .Z(out[937]) );
  ANDN U6267 ( .B(n4528), .A(n4527), .Z(n4529) );
  XNOR U6268 ( .A(n4530), .B(n4529), .Z(out[938]) );
  ANDN U6269 ( .B(n4532), .A(n4531), .Z(n4533) );
  XNOR U6270 ( .A(n4534), .B(n4533), .Z(out[939]) );
  ANDN U6271 ( .B(n4536), .A(n4535), .Z(n4537) );
  XNOR U6272 ( .A(n4538), .B(n4537), .Z(out[93]) );
  ANDN U6273 ( .B(n4540), .A(n4539), .Z(n4541) );
  XNOR U6274 ( .A(n4542), .B(n4541), .Z(out[940]) );
  ANDN U6275 ( .B(n4544), .A(n4543), .Z(n4545) );
  XNOR U6276 ( .A(n4546), .B(n4545), .Z(out[941]) );
  ANDN U6277 ( .B(n4548), .A(n4547), .Z(n4549) );
  XNOR U6278 ( .A(n4550), .B(n4549), .Z(out[942]) );
  ANDN U6279 ( .B(n4552), .A(n4551), .Z(n4553) );
  XNOR U6280 ( .A(n4554), .B(n4553), .Z(out[943]) );
  ANDN U6281 ( .B(n4556), .A(n4555), .Z(n4557) );
  XNOR U6282 ( .A(n4558), .B(n4557), .Z(out[944]) );
  ANDN U6283 ( .B(n4560), .A(n4559), .Z(n4561) );
  XNOR U6284 ( .A(n4562), .B(n4561), .Z(out[945]) );
  ANDN U6285 ( .B(n4564), .A(n4563), .Z(n4565) );
  XNOR U6286 ( .A(n4566), .B(n4565), .Z(out[946]) );
  ANDN U6287 ( .B(n4568), .A(n4567), .Z(n4569) );
  XNOR U6288 ( .A(n4570), .B(n4569), .Z(out[947]) );
  ANDN U6289 ( .B(n4572), .A(n4571), .Z(n4573) );
  XNOR U6290 ( .A(n4574), .B(n4573), .Z(out[948]) );
  ANDN U6291 ( .B(n4576), .A(n4575), .Z(n4577) );
  XNOR U6292 ( .A(n4578), .B(n4577), .Z(out[949]) );
  ANDN U6293 ( .B(n4580), .A(n4579), .Z(n4581) );
  XNOR U6294 ( .A(n4582), .B(n4581), .Z(out[94]) );
  ANDN U6295 ( .B(n4584), .A(n4583), .Z(n4585) );
  XNOR U6296 ( .A(n4586), .B(n4585), .Z(out[950]) );
  ANDN U6297 ( .B(n4588), .A(n4587), .Z(n4589) );
  XNOR U6298 ( .A(n4590), .B(n4589), .Z(out[951]) );
  ANDN U6299 ( .B(n4592), .A(n4591), .Z(n4593) );
  XNOR U6300 ( .A(n4594), .B(n4593), .Z(out[952]) );
  ANDN U6301 ( .B(n4596), .A(n4595), .Z(n4597) );
  XNOR U6302 ( .A(n4598), .B(n4597), .Z(out[953]) );
  ANDN U6303 ( .B(n4600), .A(n4599), .Z(n4601) );
  XNOR U6304 ( .A(n4602), .B(n4601), .Z(out[954]) );
  ANDN U6305 ( .B(n4604), .A(n4603), .Z(n4605) );
  XNOR U6306 ( .A(n4606), .B(n4605), .Z(out[955]) );
  ANDN U6307 ( .B(n4608), .A(n4607), .Z(n4609) );
  XNOR U6308 ( .A(n4610), .B(n4609), .Z(out[956]) );
  ANDN U6309 ( .B(n4612), .A(n4611), .Z(n4613) );
  XNOR U6310 ( .A(n4614), .B(n4613), .Z(out[957]) );
  ANDN U6311 ( .B(n4616), .A(n4615), .Z(n4617) );
  XNOR U6312 ( .A(n4618), .B(n4617), .Z(out[958]) );
  ANDN U6313 ( .B(n4620), .A(n4619), .Z(n4621) );
  XNOR U6314 ( .A(n4622), .B(n4621), .Z(out[959]) );
  ANDN U6315 ( .B(n4624), .A(n4623), .Z(n4625) );
  XNOR U6316 ( .A(n4626), .B(n4625), .Z(out[95]) );
  ANDN U6317 ( .B(n4628), .A(n4627), .Z(n4629) );
  XNOR U6318 ( .A(n4630), .B(n4629), .Z(out[960]) );
  ANDN U6319 ( .B(n4632), .A(n4631), .Z(n4633) );
  XNOR U6320 ( .A(n4634), .B(n4633), .Z(out[961]) );
  ANDN U6321 ( .B(n4636), .A(n4635), .Z(n4637) );
  XNOR U6322 ( .A(n4638), .B(n4637), .Z(out[962]) );
  ANDN U6323 ( .B(n4640), .A(n4639), .Z(n4641) );
  XNOR U6324 ( .A(n4642), .B(n4641), .Z(out[963]) );
  ANDN U6325 ( .B(n4644), .A(n4643), .Z(n4645) );
  XNOR U6326 ( .A(n4646), .B(n4645), .Z(out[964]) );
  ANDN U6327 ( .B(n4648), .A(n4647), .Z(n4649) );
  XNOR U6328 ( .A(n4650), .B(n4649), .Z(out[965]) );
  ANDN U6329 ( .B(n4652), .A(n4651), .Z(n4653) );
  XNOR U6330 ( .A(n4654), .B(n4653), .Z(out[966]) );
  ANDN U6331 ( .B(n4656), .A(n4655), .Z(n4657) );
  XNOR U6332 ( .A(n4658), .B(n4657), .Z(out[967]) );
  ANDN U6333 ( .B(n4660), .A(n4659), .Z(n4661) );
  XNOR U6334 ( .A(n4662), .B(n4661), .Z(out[968]) );
  ANDN U6335 ( .B(n4664), .A(n4663), .Z(n4665) );
  XNOR U6336 ( .A(n4666), .B(n4665), .Z(out[969]) );
  ANDN U6337 ( .B(n4668), .A(n4667), .Z(n4669) );
  XNOR U6338 ( .A(n4670), .B(n4669), .Z(out[96]) );
  ANDN U6339 ( .B(n4672), .A(n4671), .Z(n4673) );
  XNOR U6340 ( .A(n4674), .B(n4673), .Z(out[970]) );
  ANDN U6341 ( .B(n4676), .A(n4675), .Z(n4677) );
  XNOR U6342 ( .A(n4678), .B(n4677), .Z(out[971]) );
  ANDN U6343 ( .B(n4680), .A(n4679), .Z(n4681) );
  XNOR U6344 ( .A(n4682), .B(n4681), .Z(out[972]) );
  ANDN U6345 ( .B(n4684), .A(n4683), .Z(n4685) );
  XNOR U6346 ( .A(n4686), .B(n4685), .Z(out[973]) );
  ANDN U6347 ( .B(n4688), .A(n4687), .Z(n4689) );
  XNOR U6348 ( .A(n4690), .B(n4689), .Z(out[974]) );
  ANDN U6349 ( .B(n4692), .A(n4691), .Z(n4693) );
  XNOR U6350 ( .A(n4694), .B(n4693), .Z(out[975]) );
  ANDN U6351 ( .B(n4696), .A(n4695), .Z(n4697) );
  XNOR U6352 ( .A(n4698), .B(n4697), .Z(out[976]) );
  ANDN U6353 ( .B(n4700), .A(n4699), .Z(n4701) );
  XNOR U6354 ( .A(n4702), .B(n4701), .Z(out[977]) );
  ANDN U6355 ( .B(n4704), .A(n4703), .Z(n4705) );
  XNOR U6356 ( .A(n4706), .B(n4705), .Z(out[978]) );
  ANDN U6357 ( .B(n4708), .A(n4707), .Z(n4709) );
  XNOR U6358 ( .A(n4710), .B(n4709), .Z(out[979]) );
  ANDN U6359 ( .B(n4712), .A(n4711), .Z(n4713) );
  XNOR U6360 ( .A(n4714), .B(n4713), .Z(out[97]) );
  ANDN U6361 ( .B(n4716), .A(n4715), .Z(n4717) );
  XNOR U6362 ( .A(n4718), .B(n4717), .Z(out[980]) );
  ANDN U6363 ( .B(n4720), .A(n4719), .Z(n4721) );
  XNOR U6364 ( .A(n4722), .B(n4721), .Z(out[981]) );
  ANDN U6365 ( .B(n4724), .A(n4723), .Z(n4725) );
  XNOR U6366 ( .A(n4726), .B(n4725), .Z(out[982]) );
  ANDN U6367 ( .B(n4728), .A(n4727), .Z(n4729) );
  XNOR U6368 ( .A(n4730), .B(n4729), .Z(out[983]) );
  ANDN U6369 ( .B(n4732), .A(n4731), .Z(n4733) );
  XNOR U6370 ( .A(n4734), .B(n4733), .Z(out[984]) );
  ANDN U6371 ( .B(n4736), .A(n4735), .Z(n4737) );
  XNOR U6372 ( .A(n4738), .B(n4737), .Z(out[985]) );
  ANDN U6373 ( .B(n4740), .A(n4739), .Z(n4741) );
  XNOR U6374 ( .A(n4742), .B(n4741), .Z(out[986]) );
  ANDN U6375 ( .B(n4744), .A(n4743), .Z(n4745) );
  XNOR U6376 ( .A(n4746), .B(n4745), .Z(out[987]) );
  ANDN U6377 ( .B(n4748), .A(n4747), .Z(n4749) );
  XNOR U6378 ( .A(n4750), .B(n4749), .Z(out[988]) );
  ANDN U6379 ( .B(n4752), .A(n4751), .Z(n4753) );
  XNOR U6380 ( .A(n4754), .B(n4753), .Z(out[989]) );
  ANDN U6381 ( .B(n4756), .A(n4755), .Z(n4757) );
  XNOR U6382 ( .A(n4758), .B(n4757), .Z(out[98]) );
  ANDN U6383 ( .B(n4760), .A(n4759), .Z(n4761) );
  XNOR U6384 ( .A(n4762), .B(n4761), .Z(out[990]) );
  ANDN U6385 ( .B(n4764), .A(n4763), .Z(n4765) );
  XNOR U6386 ( .A(n4766), .B(n4765), .Z(out[991]) );
  ANDN U6387 ( .B(n4768), .A(n4767), .Z(n4769) );
  XNOR U6388 ( .A(n4770), .B(n4769), .Z(out[992]) );
  ANDN U6389 ( .B(n4772), .A(n4771), .Z(n4773) );
  XNOR U6390 ( .A(n4774), .B(n4773), .Z(out[993]) );
  ANDN U6391 ( .B(n4776), .A(n4775), .Z(n4777) );
  XNOR U6392 ( .A(n4778), .B(n4777), .Z(out[994]) );
  ANDN U6393 ( .B(n4780), .A(n4779), .Z(n4781) );
  XNOR U6394 ( .A(n4782), .B(n4781), .Z(out[995]) );
  ANDN U6395 ( .B(n4784), .A(n4783), .Z(n4785) );
  XNOR U6396 ( .A(n4786), .B(n4785), .Z(out[996]) );
  ANDN U6397 ( .B(n4788), .A(n4787), .Z(n4789) );
  XNOR U6398 ( .A(n4790), .B(n4789), .Z(out[997]) );
  ANDN U6399 ( .B(n4792), .A(n4791), .Z(n4793) );
  XNOR U6400 ( .A(n4794), .B(n4793), .Z(out[998]) );
  ANDN U6401 ( .B(n4796), .A(n4795), .Z(n4797) );
  XNOR U6402 ( .A(n4798), .B(n4797), .Z(out[999]) );
  ANDN U6403 ( .B(n4800), .A(n4799), .Z(n4801) );
  XNOR U6404 ( .A(n4802), .B(n4801), .Z(out[99]) );
  OR U6405 ( .A(n4804), .B(n4803), .Z(n4805) );
  XNOR U6406 ( .A(n4806), .B(n4805), .Z(out[9]) );
endmodule


module round_4 ( in, round_const, out );
  input [1599:0] in;
  input [63:0] round_const;
  output [1599:0] out;
  wire   round_const_31, round_const_15, round_const_7, round_const_3, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807;
  assign round_const_31 = round_const[31];
  assign round_const_15 = round_const[15];
  assign round_const_7 = round_const[7];
  assign round_const_3 = round_const[3];

  XOR U1 ( .A(in[1469]), .B(in[509]), .Z(n2) );
  XNOR U2 ( .A(in[829]), .B(in[189]), .Z(n1) );
  XNOR U3 ( .A(n2), .B(n1), .Z(n3) );
  XOR U4 ( .A(in[1149]), .B(n3), .Z(n872) );
  XOR U5 ( .A(in[1598]), .B(in[638]), .Z(n5) );
  XNOR U6 ( .A(in[958]), .B(in[318]), .Z(n4) );
  XNOR U7 ( .A(n5), .B(n4), .Z(n6) );
  XOR U8 ( .A(in[1278]), .B(n6), .Z(n1473) );
  XNOR U9 ( .A(n872), .B(n1473), .Z(n3815) );
  XNOR U10 ( .A(in[254]), .B(n3815), .Z(n3577) );
  XOR U11 ( .A(in[1345]), .B(in[65]), .Z(n8) );
  XNOR U12 ( .A(in[1025]), .B(in[385]), .Z(n7) );
  XNOR U13 ( .A(n8), .B(n7), .Z(n9) );
  XOR U14 ( .A(in[705]), .B(n9), .Z(n1481) );
  XOR U15 ( .A(in[1474]), .B(in[514]), .Z(n11) );
  XNOR U16 ( .A(in[834]), .B(in[194]), .Z(n10) );
  XNOR U17 ( .A(n11), .B(n10), .Z(n12) );
  XNOR U18 ( .A(in[1154]), .B(n12), .Z(n1188) );
  XNOR U19 ( .A(n1481), .B(n1188), .Z(n3570) );
  XNOR U20 ( .A(in[1410]), .B(n3570), .Z(n3576) );
  XOR U21 ( .A(in[137]), .B(in[457]), .Z(n14) );
  XNOR U22 ( .A(in[777]), .B(in[1417]), .Z(n13) );
  XNOR U23 ( .A(n14), .B(n13), .Z(n15) );
  XOR U24 ( .A(in[1097]), .B(n15), .Z(n1141) );
  XOR U25 ( .A(in[328]), .B(in[8]), .Z(n17) );
  XNOR U26 ( .A(in[968]), .B(in[648]), .Z(n16) );
  XNOR U27 ( .A(n17), .B(n16), .Z(n18) );
  XOR U28 ( .A(in[1288]), .B(n18), .Z(n1209) );
  XNOR U29 ( .A(n1141), .B(n1209), .Z(n4086) );
  XNOR U30 ( .A(in[1033]), .B(n4086), .Z(n2609) );
  NAND U31 ( .A(n3576), .B(n2609), .Z(n19) );
  XNOR U32 ( .A(n3577), .B(n19), .Z(out[0]) );
  XOR U33 ( .A(in[1386]), .B(in[106]), .Z(n21) );
  XNOR U34 ( .A(in[1066]), .B(in[746]), .Z(n20) );
  XNOR U35 ( .A(n21), .B(n20), .Z(n22) );
  XOR U36 ( .A(in[426]), .B(n22), .Z(n475) );
  XOR U37 ( .A(in[1515]), .B(in[555]), .Z(n24) );
  XNOR U38 ( .A(in[875]), .B(in[235]), .Z(n23) );
  XNOR U39 ( .A(n24), .B(n23), .Z(n25) );
  XOR U40 ( .A(in[1195]), .B(n25), .Z(n1329) );
  XNOR U41 ( .A(n475), .B(n1329), .Z(n3750) );
  XNOR U42 ( .A(in[171]), .B(n3750), .Z(n1301) );
  XOR U43 ( .A(in[971]), .B(in[1291]), .Z(n27) );
  XNOR U44 ( .A(in[11]), .B(in[331]), .Z(n26) );
  XNOR U45 ( .A(n27), .B(n26), .Z(n28) );
  XOR U46 ( .A(in[651]), .B(n28), .Z(n1220) );
  XOR U47 ( .A(in[140]), .B(in[460]), .Z(n30) );
  XNOR U48 ( .A(in[1100]), .B(in[1420]), .Z(n29) );
  XNOR U49 ( .A(n30), .B(n29), .Z(n31) );
  XNOR U50 ( .A(in[780]), .B(n31), .Z(n1159) );
  XNOR U51 ( .A(n1220), .B(n1159), .Z(n4095) );
  XNOR U52 ( .A(in[1356]), .B(n4095), .Z(n1696) );
  XOR U53 ( .A(in[1364]), .B(in[724]), .Z(n33) );
  XNOR U54 ( .A(in[84]), .B(in[404]), .Z(n32) );
  XNOR U55 ( .A(n33), .B(n32), .Z(n34) );
  XOR U56 ( .A(in[1044]), .B(n34), .Z(n777) );
  XOR U57 ( .A(in[1555]), .B(in[595]), .Z(n36) );
  XNOR U58 ( .A(in[915]), .B(in[275]), .Z(n35) );
  XNOR U59 ( .A(n36), .B(n35), .Z(n37) );
  XOR U60 ( .A(in[1235]), .B(n37), .Z(n489) );
  XNOR U61 ( .A(n777), .B(n489), .Z(n3882) );
  XNOR U62 ( .A(in[980]), .B(n3882), .Z(n1693) );
  NAND U63 ( .A(n1696), .B(n1693), .Z(n38) );
  XNOR U64 ( .A(n1301), .B(n38), .Z(out[1000]) );
  XOR U65 ( .A(in[1387]), .B(in[107]), .Z(n40) );
  XNOR U66 ( .A(in[1067]), .B(in[747]), .Z(n39) );
  XNOR U67 ( .A(n40), .B(n39), .Z(n41) );
  XOR U68 ( .A(in[427]), .B(n41), .Z(n486) );
  XOR U69 ( .A(in[1516]), .B(in[556]), .Z(n43) );
  XNOR U70 ( .A(in[876]), .B(in[236]), .Z(n42) );
  XNOR U71 ( .A(n43), .B(n42), .Z(n44) );
  XOR U72 ( .A(in[1196]), .B(n44), .Z(n1333) );
  XNOR U73 ( .A(n486), .B(n1333), .Z(n3758) );
  XNOR U74 ( .A(in[172]), .B(n3758), .Z(n1305) );
  XOR U75 ( .A(in[972]), .B(in[12]), .Z(n46) );
  XNOR U76 ( .A(in[1292]), .B(in[332]), .Z(n45) );
  XNOR U77 ( .A(n46), .B(n45), .Z(n47) );
  XOR U78 ( .A(in[652]), .B(n47), .Z(n1223) );
  XOR U79 ( .A(in[141]), .B(in[461]), .Z(n49) );
  XNOR U80 ( .A(in[1101]), .B(in[1421]), .Z(n48) );
  XNOR U81 ( .A(n49), .B(n48), .Z(n50) );
  XNOR U82 ( .A(in[781]), .B(n50), .Z(n1164) );
  XNOR U83 ( .A(n1223), .B(n1164), .Z(n4098) );
  XNOR U84 ( .A(in[1357]), .B(n4098), .Z(n1700) );
  XOR U85 ( .A(in[1365]), .B(in[725]), .Z(n52) );
  XNOR U86 ( .A(in[85]), .B(in[405]), .Z(n51) );
  XNOR U87 ( .A(n52), .B(n51), .Z(n53) );
  XOR U88 ( .A(in[1045]), .B(n53), .Z(n790) );
  XOR U89 ( .A(in[1556]), .B(in[596]), .Z(n55) );
  XNOR U90 ( .A(in[916]), .B(in[276]), .Z(n54) );
  XNOR U91 ( .A(n55), .B(n54), .Z(n56) );
  XOR U92 ( .A(in[1236]), .B(n56), .Z(n504) );
  XNOR U93 ( .A(n790), .B(n504), .Z(n3884) );
  XNOR U94 ( .A(in[981]), .B(n3884), .Z(n1697) );
  NAND U95 ( .A(n1700), .B(n1697), .Z(n57) );
  XNOR U96 ( .A(n1305), .B(n57), .Z(out[1001]) );
  XOR U97 ( .A(in[1388]), .B(in[108]), .Z(n59) );
  XNOR U98 ( .A(in[1068]), .B(in[748]), .Z(n58) );
  XNOR U99 ( .A(n59), .B(n58), .Z(n60) );
  XOR U100 ( .A(in[428]), .B(n60), .Z(n1395) );
  XOR U101 ( .A(in[1517]), .B(in[557]), .Z(n62) );
  XNOR U102 ( .A(in[877]), .B(in[237]), .Z(n61) );
  XNOR U103 ( .A(n62), .B(n61), .Z(n63) );
  XOR U104 ( .A(in[1197]), .B(n63), .Z(n1337) );
  XNOR U105 ( .A(n1395), .B(n1337), .Z(n3762) );
  XNOR U106 ( .A(in[173]), .B(n3762), .Z(n1310) );
  XOR U107 ( .A(in[973]), .B(in[13]), .Z(n65) );
  XNOR U108 ( .A(in[1293]), .B(in[333]), .Z(n64) );
  XNOR U109 ( .A(n65), .B(n64), .Z(n66) );
  XOR U110 ( .A(in[653]), .B(n66), .Z(n1226) );
  XOR U111 ( .A(in[142]), .B(in[1422]), .Z(n68) );
  XNOR U112 ( .A(in[1102]), .B(in[782]), .Z(n67) );
  XNOR U113 ( .A(n68), .B(n67), .Z(n69) );
  XNOR U114 ( .A(in[462]), .B(n69), .Z(n1169) );
  XNOR U115 ( .A(n1226), .B(n1169), .Z(n4101) );
  XNOR U116 ( .A(in[1358]), .B(n4101), .Z(n1704) );
  XOR U117 ( .A(in[1366]), .B(in[726]), .Z(n71) );
  XNOR U118 ( .A(in[86]), .B(in[406]), .Z(n70) );
  XNOR U119 ( .A(n71), .B(n70), .Z(n72) );
  XOR U120 ( .A(in[1046]), .B(n72), .Z(n803) );
  XOR U121 ( .A(in[1557]), .B(in[597]), .Z(n74) );
  XNOR U122 ( .A(in[917]), .B(in[277]), .Z(n73) );
  XNOR U123 ( .A(n74), .B(n73), .Z(n75) );
  XOR U124 ( .A(in[1237]), .B(n75), .Z(n519) );
  XNOR U125 ( .A(n803), .B(n519), .Z(n3886) );
  XNOR U126 ( .A(in[982]), .B(n3886), .Z(n1701) );
  NAND U127 ( .A(n1704), .B(n1701), .Z(n76) );
  XNOR U128 ( .A(n1310), .B(n76), .Z(out[1002]) );
  XOR U129 ( .A(in[1389]), .B(in[109]), .Z(n78) );
  XNOR U130 ( .A(in[1069]), .B(in[749]), .Z(n77) );
  XNOR U131 ( .A(n78), .B(n77), .Z(n79) );
  XOR U132 ( .A(in[429]), .B(n79), .Z(n1399) );
  XOR U133 ( .A(in[1518]), .B(in[558]), .Z(n81) );
  XNOR U134 ( .A(in[878]), .B(in[238]), .Z(n80) );
  XNOR U135 ( .A(n81), .B(n80), .Z(n82) );
  XOR U136 ( .A(in[1198]), .B(n82), .Z(n1341) );
  XNOR U137 ( .A(n1399), .B(n1341), .Z(n3766) );
  XNOR U138 ( .A(in[174]), .B(n3766), .Z(n1314) );
  XOR U139 ( .A(in[974]), .B(in[14]), .Z(n84) );
  XNOR U140 ( .A(in[1294]), .B(in[334]), .Z(n83) );
  XNOR U141 ( .A(n84), .B(n83), .Z(n85) );
  XOR U142 ( .A(in[654]), .B(n85), .Z(n1229) );
  XOR U143 ( .A(in[143]), .B(in[1423]), .Z(n87) );
  XNOR U144 ( .A(in[1103]), .B(in[783]), .Z(n86) );
  XNOR U145 ( .A(n87), .B(n86), .Z(n88) );
  XNOR U146 ( .A(in[463]), .B(n88), .Z(n1174) );
  XNOR U147 ( .A(n1229), .B(n1174), .Z(n4104) );
  XNOR U148 ( .A(in[1359]), .B(n4104), .Z(n1708) );
  XOR U149 ( .A(in[1367]), .B(in[727]), .Z(n90) );
  XNOR U150 ( .A(in[87]), .B(in[407]), .Z(n89) );
  XNOR U151 ( .A(n90), .B(n89), .Z(n91) );
  XOR U152 ( .A(in[1047]), .B(n91), .Z(n816) );
  XOR U153 ( .A(in[1558]), .B(in[598]), .Z(n93) );
  XNOR U154 ( .A(in[918]), .B(in[278]), .Z(n92) );
  XNOR U155 ( .A(n93), .B(n92), .Z(n94) );
  XOR U156 ( .A(in[1238]), .B(n94), .Z(n534) );
  XNOR U157 ( .A(n816), .B(n534), .Z(n3888) );
  XNOR U158 ( .A(in[983]), .B(n3888), .Z(n1705) );
  NAND U159 ( .A(n1708), .B(n1705), .Z(n95) );
  XNOR U160 ( .A(n1314), .B(n95), .Z(out[1003]) );
  XOR U161 ( .A(in[1390]), .B(in[110]), .Z(n97) );
  XNOR U162 ( .A(in[1070]), .B(in[750]), .Z(n96) );
  XNOR U163 ( .A(n97), .B(n96), .Z(n98) );
  XOR U164 ( .A(in[430]), .B(n98), .Z(n1403) );
  XOR U165 ( .A(in[1519]), .B(in[559]), .Z(n100) );
  XNOR U166 ( .A(in[879]), .B(in[239]), .Z(n99) );
  XNOR U167 ( .A(n100), .B(n99), .Z(n101) );
  XOR U168 ( .A(in[1199]), .B(n101), .Z(n1345) );
  XNOR U169 ( .A(n1403), .B(n1345), .Z(n3770) );
  XNOR U170 ( .A(in[175]), .B(n3770), .Z(n1318) );
  XOR U171 ( .A(in[975]), .B(in[15]), .Z(n103) );
  XNOR U172 ( .A(in[1295]), .B(in[335]), .Z(n102) );
  XNOR U173 ( .A(n103), .B(n102), .Z(n104) );
  XOR U174 ( .A(in[655]), .B(n104), .Z(n1232) );
  XOR U175 ( .A(in[144]), .B(in[1424]), .Z(n106) );
  XNOR U176 ( .A(in[1104]), .B(in[784]), .Z(n105) );
  XNOR U177 ( .A(n106), .B(n105), .Z(n107) );
  XNOR U178 ( .A(in[464]), .B(n107), .Z(n1179) );
  XNOR U179 ( .A(n1232), .B(n1179), .Z(n4107) );
  XNOR U180 ( .A(in[1360]), .B(n4107), .Z(n1713) );
  XOR U181 ( .A(in[1368]), .B(in[728]), .Z(n109) );
  XNOR U182 ( .A(in[88]), .B(in[408]), .Z(n108) );
  XNOR U183 ( .A(n109), .B(n108), .Z(n110) );
  XOR U184 ( .A(in[1048]), .B(n110), .Z(n829) );
  XOR U185 ( .A(in[1559]), .B(in[599]), .Z(n112) );
  XNOR U186 ( .A(in[919]), .B(in[279]), .Z(n111) );
  XNOR U187 ( .A(n112), .B(n111), .Z(n113) );
  XOR U188 ( .A(in[1239]), .B(n113), .Z(n549) );
  XNOR U189 ( .A(n829), .B(n549), .Z(n3890) );
  XNOR U190 ( .A(in[984]), .B(n3890), .Z(n1710) );
  NAND U191 ( .A(n1713), .B(n1710), .Z(n114) );
  XNOR U192 ( .A(n1318), .B(n114), .Z(out[1004]) );
  XOR U193 ( .A(in[1391]), .B(in[111]), .Z(n116) );
  XNOR U194 ( .A(in[1071]), .B(in[751]), .Z(n115) );
  XNOR U195 ( .A(n116), .B(n115), .Z(n117) );
  XOR U196 ( .A(in[431]), .B(n117), .Z(n1407) );
  XOR U197 ( .A(in[1520]), .B(in[560]), .Z(n119) );
  XNOR U198 ( .A(in[880]), .B(in[240]), .Z(n118) );
  XNOR U199 ( .A(n119), .B(n118), .Z(n120) );
  XOR U200 ( .A(in[1200]), .B(n120), .Z(n1350) );
  XNOR U201 ( .A(n1407), .B(n1350), .Z(n3774) );
  XNOR U202 ( .A(in[176]), .B(n3774), .Z(n1322) );
  XOR U203 ( .A(in[976]), .B(in[16]), .Z(n122) );
  XNOR U204 ( .A(in[1296]), .B(in[336]), .Z(n121) );
  XNOR U205 ( .A(n122), .B(n121), .Z(n123) );
  XOR U206 ( .A(in[656]), .B(n123), .Z(n1235) );
  XOR U207 ( .A(in[145]), .B(in[1425]), .Z(n125) );
  XNOR U208 ( .A(in[1105]), .B(in[785]), .Z(n124) );
  XNOR U209 ( .A(n125), .B(n124), .Z(n126) );
  XNOR U210 ( .A(in[465]), .B(n126), .Z(n1184) );
  XNOR U211 ( .A(n1235), .B(n1184), .Z(n4114) );
  XNOR U212 ( .A(in[1361]), .B(n4114), .Z(n1717) );
  XOR U213 ( .A(in[1369]), .B(in[729]), .Z(n128) );
  XNOR U214 ( .A(in[89]), .B(in[409]), .Z(n127) );
  XNOR U215 ( .A(n128), .B(n127), .Z(n129) );
  XOR U216 ( .A(in[1049]), .B(n129), .Z(n842) );
  XOR U217 ( .A(in[1560]), .B(in[600]), .Z(n131) );
  XNOR U218 ( .A(in[920]), .B(in[280]), .Z(n130) );
  XNOR U219 ( .A(n131), .B(n130), .Z(n132) );
  XOR U220 ( .A(in[1240]), .B(n132), .Z(n564) );
  XNOR U221 ( .A(n842), .B(n564), .Z(n3892) );
  XNOR U222 ( .A(in[985]), .B(n3892), .Z(n1714) );
  NAND U223 ( .A(n1717), .B(n1714), .Z(n133) );
  XNOR U224 ( .A(n1322), .B(n133), .Z(out[1005]) );
  XOR U225 ( .A(in[1392]), .B(in[112]), .Z(n135) );
  XNOR U226 ( .A(in[1072]), .B(in[752]), .Z(n134) );
  XNOR U227 ( .A(n135), .B(n134), .Z(n136) );
  XOR U228 ( .A(in[432]), .B(n136), .Z(n1411) );
  XOR U229 ( .A(in[1521]), .B(in[561]), .Z(n138) );
  XNOR U230 ( .A(in[881]), .B(in[241]), .Z(n137) );
  XNOR U231 ( .A(n138), .B(n137), .Z(n139) );
  XOR U232 ( .A(in[1201]), .B(n139), .Z(n1354) );
  XNOR U233 ( .A(n1411), .B(n1354), .Z(n3778) );
  XNOR U234 ( .A(in[177]), .B(n3778), .Z(n1326) );
  XOR U235 ( .A(in[1426]), .B(in[466]), .Z(n141) );
  XNOR U236 ( .A(in[786]), .B(in[146]), .Z(n140) );
  XNOR U237 ( .A(n141), .B(n140), .Z(n142) );
  XOR U238 ( .A(in[1106]), .B(n142), .Z(n488) );
  XOR U239 ( .A(in[17]), .B(in[657]), .Z(n144) );
  XNOR U240 ( .A(in[977]), .B(in[337]), .Z(n143) );
  XNOR U241 ( .A(n144), .B(n143), .Z(n145) );
  XNOR U242 ( .A(in[1297]), .B(n145), .Z(n1238) );
  XNOR U243 ( .A(n488), .B(n1238), .Z(n4117) );
  XNOR U244 ( .A(n4117), .B(in[1362]), .Z(n1721) );
  XOR U245 ( .A(in[1370]), .B(in[730]), .Z(n147) );
  XNOR U246 ( .A(in[90]), .B(in[410]), .Z(n146) );
  XNOR U247 ( .A(n147), .B(n146), .Z(n148) );
  XOR U248 ( .A(in[1050]), .B(n148), .Z(n857) );
  XOR U249 ( .A(in[1561]), .B(in[601]), .Z(n150) );
  XNOR U250 ( .A(in[921]), .B(in[281]), .Z(n149) );
  XNOR U251 ( .A(n150), .B(n149), .Z(n151) );
  XOR U252 ( .A(in[1241]), .B(n151), .Z(n590) );
  XNOR U253 ( .A(n857), .B(n590), .Z(n3894) );
  XNOR U254 ( .A(in[986]), .B(n3894), .Z(n1718) );
  NAND U255 ( .A(n1721), .B(n1718), .Z(n152) );
  XNOR U256 ( .A(n1326), .B(n152), .Z(out[1006]) );
  XOR U257 ( .A(in[1393]), .B(in[113]), .Z(n154) );
  XNOR U258 ( .A(in[1073]), .B(in[753]), .Z(n153) );
  XNOR U259 ( .A(n154), .B(n153), .Z(n155) );
  XOR U260 ( .A(in[433]), .B(n155), .Z(n1415) );
  XOR U261 ( .A(in[1522]), .B(in[562]), .Z(n157) );
  XNOR U262 ( .A(in[882]), .B(in[242]), .Z(n156) );
  XNOR U263 ( .A(n157), .B(n156), .Z(n158) );
  XOR U264 ( .A(in[1202]), .B(n158), .Z(n1358) );
  XNOR U265 ( .A(n1415), .B(n1358), .Z(n3782) );
  XNOR U266 ( .A(in[178]), .B(n3782), .Z(n1330) );
  XOR U267 ( .A(in[147]), .B(in[1427]), .Z(n160) );
  XNOR U268 ( .A(in[1107]), .B(in[787]), .Z(n159) );
  XNOR U269 ( .A(n160), .B(n159), .Z(n161) );
  XOR U270 ( .A(in[467]), .B(n161), .Z(n503) );
  XOR U271 ( .A(in[978]), .B(in[18]), .Z(n163) );
  XNOR U272 ( .A(in[1298]), .B(in[338]), .Z(n162) );
  XNOR U273 ( .A(n163), .B(n162), .Z(n164) );
  XNOR U274 ( .A(in[658]), .B(n164), .Z(n1241) );
  XNOR U275 ( .A(n503), .B(n1241), .Z(n4120) );
  XNOR U276 ( .A(in[1363]), .B(n4120), .Z(n1725) );
  XOR U277 ( .A(in[1371]), .B(in[731]), .Z(n166) );
  XNOR U278 ( .A(in[91]), .B(in[411]), .Z(n165) );
  XNOR U279 ( .A(n166), .B(n165), .Z(n167) );
  XOR U280 ( .A(in[1051]), .B(n167), .Z(n870) );
  XOR U281 ( .A(in[1562]), .B(in[602]), .Z(n169) );
  XNOR U282 ( .A(in[922]), .B(in[282]), .Z(n168) );
  XNOR U283 ( .A(n169), .B(n168), .Z(n170) );
  XOR U284 ( .A(in[1242]), .B(n170), .Z(n605) );
  XNOR U285 ( .A(n870), .B(n605), .Z(n3896) );
  XNOR U286 ( .A(in[987]), .B(n3896), .Z(n1722) );
  NAND U287 ( .A(n1725), .B(n1722), .Z(n171) );
  XNOR U288 ( .A(n1330), .B(n171), .Z(out[1007]) );
  XOR U289 ( .A(in[1394]), .B(in[114]), .Z(n173) );
  XNOR U290 ( .A(in[1074]), .B(in[754]), .Z(n172) );
  XNOR U291 ( .A(n173), .B(n172), .Z(n174) );
  XOR U292 ( .A(in[434]), .B(n174), .Z(n1419) );
  XOR U293 ( .A(in[1523]), .B(in[563]), .Z(n176) );
  XNOR U294 ( .A(in[883]), .B(in[243]), .Z(n175) );
  XNOR U295 ( .A(n176), .B(n175), .Z(n177) );
  XOR U296 ( .A(in[1203]), .B(n177), .Z(n1362) );
  XNOR U297 ( .A(n1419), .B(n1362), .Z(n3786) );
  XNOR U298 ( .A(in[179]), .B(n3786), .Z(n1334) );
  XOR U299 ( .A(in[979]), .B(in[19]), .Z(n179) );
  XNOR U300 ( .A(in[1299]), .B(in[339]), .Z(n178) );
  XNOR U301 ( .A(n179), .B(n178), .Z(n180) );
  XOR U302 ( .A(in[659]), .B(n180), .Z(n1245) );
  XOR U303 ( .A(in[148]), .B(in[1428]), .Z(n182) );
  XNOR U304 ( .A(in[1108]), .B(in[788]), .Z(n181) );
  XNOR U305 ( .A(n182), .B(n181), .Z(n183) );
  XNOR U306 ( .A(in[468]), .B(n183), .Z(n518) );
  XNOR U307 ( .A(n1245), .B(n518), .Z(n4123) );
  XNOR U308 ( .A(in[1364]), .B(n4123), .Z(n1729) );
  XOR U309 ( .A(in[1372]), .B(in[732]), .Z(n185) );
  XNOR U310 ( .A(in[92]), .B(in[412]), .Z(n184) );
  XNOR U311 ( .A(n185), .B(n184), .Z(n186) );
  XOR U312 ( .A(in[1052]), .B(n186), .Z(n890) );
  XOR U313 ( .A(in[1563]), .B(in[603]), .Z(n188) );
  XNOR U314 ( .A(in[923]), .B(in[283]), .Z(n187) );
  XNOR U315 ( .A(n188), .B(n187), .Z(n189) );
  XOR U316 ( .A(in[1243]), .B(n189), .Z(n620) );
  XNOR U317 ( .A(n890), .B(n620), .Z(n3900) );
  XNOR U318 ( .A(in[988]), .B(n3900), .Z(n1726) );
  NAND U319 ( .A(n1729), .B(n1726), .Z(n190) );
  XNOR U320 ( .A(n1334), .B(n190), .Z(out[1008]) );
  XOR U321 ( .A(in[1395]), .B(in[115]), .Z(n192) );
  XNOR U322 ( .A(in[1075]), .B(in[755]), .Z(n191) );
  XNOR U323 ( .A(n192), .B(n191), .Z(n193) );
  XOR U324 ( .A(in[435]), .B(n193), .Z(n1423) );
  XOR U325 ( .A(in[1524]), .B(in[564]), .Z(n195) );
  XNOR U326 ( .A(in[884]), .B(in[244]), .Z(n194) );
  XNOR U327 ( .A(n195), .B(n194), .Z(n196) );
  XOR U328 ( .A(in[1204]), .B(n196), .Z(n1366) );
  XNOR U329 ( .A(n1423), .B(n1366), .Z(n3790) );
  XNOR U330 ( .A(in[180]), .B(n3790), .Z(n1338) );
  XOR U331 ( .A(in[149]), .B(in[1429]), .Z(n198) );
  XNOR U332 ( .A(in[1109]), .B(in[789]), .Z(n197) );
  XNOR U333 ( .A(n198), .B(n197), .Z(n199) );
  XOR U334 ( .A(in[469]), .B(n199), .Z(n533) );
  XOR U335 ( .A(in[340]), .B(in[660]), .Z(n201) );
  XNOR U336 ( .A(in[20]), .B(in[1300]), .Z(n200) );
  XNOR U337 ( .A(n201), .B(n200), .Z(n202) );
  XNOR U338 ( .A(in[980]), .B(n202), .Z(n1248) );
  XNOR U339 ( .A(n533), .B(n1248), .Z(n4126) );
  XNOR U340 ( .A(in[1365]), .B(n4126), .Z(n1733) );
  XOR U341 ( .A(in[1373]), .B(in[733]), .Z(n204) );
  XNOR U342 ( .A(in[93]), .B(in[413]), .Z(n203) );
  XNOR U343 ( .A(n204), .B(n203), .Z(n205) );
  XOR U344 ( .A(in[1053]), .B(n205), .Z(n903) );
  XOR U345 ( .A(in[1564]), .B(in[604]), .Z(n207) );
  XNOR U346 ( .A(in[924]), .B(in[284]), .Z(n206) );
  XNOR U347 ( .A(n207), .B(n206), .Z(n208) );
  XOR U348 ( .A(in[1244]), .B(n208), .Z(n635) );
  XNOR U349 ( .A(n903), .B(n635), .Z(n3902) );
  XNOR U350 ( .A(in[989]), .B(n3902), .Z(n1730) );
  NAND U351 ( .A(n1733), .B(n1730), .Z(n209) );
  XNOR U352 ( .A(n1338), .B(n209), .Z(out[1009]) );
  XOR U353 ( .A(in[1339]), .B(in[59]), .Z(n211) );
  XNOR U354 ( .A(in[699]), .B(in[379]), .Z(n210) );
  XNOR U355 ( .A(n211), .B(n210), .Z(n212) );
  XOR U356 ( .A(in[1019]), .B(n212), .Z(n861) );
  XOR U357 ( .A(in[1530]), .B(in[570]), .Z(n214) );
  XNOR U358 ( .A(in[1210]), .B(in[250]), .Z(n213) );
  XNOR U359 ( .A(n214), .B(n213), .Z(n215) );
  XOR U360 ( .A(in[890]), .B(n215), .Z(n327) );
  XNOR U361 ( .A(n861), .B(n327), .Z(n3592) );
  XNOR U362 ( .A(in[635]), .B(n3592), .Z(n2550) );
  XOR U363 ( .A(in[161]), .B(in[1441]), .Z(n217) );
  XNOR U364 ( .A(in[801]), .B(in[1121]), .Z(n216) );
  XNOR U365 ( .A(n217), .B(n216), .Z(n218) );
  XOR U366 ( .A(in[481]), .B(n218), .Z(n454) );
  XOR U367 ( .A(in[1570]), .B(in[610]), .Z(n220) );
  XNOR U368 ( .A(in[930]), .B(in[290]), .Z(n219) );
  XNOR U369 ( .A(n220), .B(n219), .Z(n221) );
  XNOR U370 ( .A(in[1250]), .B(n221), .Z(n337) );
  XNOR U371 ( .A(n454), .B(n337), .Z(n3689) );
  XNOR U372 ( .A(in[226]), .B(n3689), .Z(n2831) );
  XOR U373 ( .A(in[1061]), .B(in[421]), .Z(n223) );
  XNOR U374 ( .A(in[741]), .B(in[1381]), .Z(n222) );
  XNOR U375 ( .A(n223), .B(n222), .Z(n224) );
  XOR U376 ( .A(in[101]), .B(n224), .Z(n373) );
  XOR U377 ( .A(in[1510]), .B(in[550]), .Z(n226) );
  XNOR U378 ( .A(in[870]), .B(in[230]), .Z(n225) );
  XNOR U379 ( .A(n226), .B(n225), .Z(n227) );
  XOR U380 ( .A(in[1190]), .B(n227), .Z(n1309) );
  XNOR U381 ( .A(n373), .B(n1309), .Z(n3730) );
  XNOR U382 ( .A(in[1446]), .B(n3730), .Z(n2828) );
  NAND U383 ( .A(n2831), .B(n2828), .Z(n228) );
  XNOR U384 ( .A(n2550), .B(n228), .Z(out[100]) );
  XOR U385 ( .A(in[1396]), .B(in[116]), .Z(n230) );
  XNOR U386 ( .A(in[1076]), .B(in[756]), .Z(n229) );
  XNOR U387 ( .A(n230), .B(n229), .Z(n231) );
  XOR U388 ( .A(in[436]), .B(n231), .Z(n1428) );
  XOR U389 ( .A(in[1525]), .B(in[565]), .Z(n233) );
  XNOR U390 ( .A(in[885]), .B(in[245]), .Z(n232) );
  XNOR U391 ( .A(n233), .B(n232), .Z(n234) );
  XOR U392 ( .A(in[1205]), .B(n234), .Z(n1370) );
  XNOR U393 ( .A(n1428), .B(n1370), .Z(n3794) );
  XNOR U394 ( .A(in[181]), .B(n3794), .Z(n1342) );
  XOR U395 ( .A(in[341]), .B(in[661]), .Z(n236) );
  XNOR U396 ( .A(in[21]), .B(in[1301]), .Z(n235) );
  XNOR U397 ( .A(n236), .B(n235), .Z(n237) );
  XOR U398 ( .A(in[981]), .B(n237), .Z(n1251) );
  XOR U399 ( .A(in[150]), .B(in[1430]), .Z(n239) );
  XNOR U400 ( .A(in[1110]), .B(in[790]), .Z(n238) );
  XNOR U401 ( .A(n239), .B(n238), .Z(n240) );
  XNOR U402 ( .A(in[470]), .B(n240), .Z(n548) );
  XNOR U403 ( .A(n1251), .B(n548), .Z(n4129) );
  XNOR U404 ( .A(in[1366]), .B(n4129), .Z(n1737) );
  XOR U405 ( .A(in[1374]), .B(in[734]), .Z(n242) );
  XNOR U406 ( .A(in[94]), .B(in[414]), .Z(n241) );
  XNOR U407 ( .A(n242), .B(n241), .Z(n243) );
  XOR U408 ( .A(in[1054]), .B(n243), .Z(n916) );
  XOR U409 ( .A(in[1565]), .B(in[605]), .Z(n245) );
  XNOR U410 ( .A(in[925]), .B(in[285]), .Z(n244) );
  XNOR U411 ( .A(n245), .B(n244), .Z(n246) );
  XOR U412 ( .A(in[1245]), .B(n246), .Z(n650) );
  XNOR U413 ( .A(n916), .B(n650), .Z(n3904) );
  XNOR U414 ( .A(in[990]), .B(n3904), .Z(n1734) );
  NAND U415 ( .A(n1737), .B(n1734), .Z(n247) );
  XNOR U416 ( .A(n1342), .B(n247), .Z(out[1010]) );
  XOR U417 ( .A(in[1526]), .B(in[566]), .Z(n249) );
  XNOR U418 ( .A(in[886]), .B(in[246]), .Z(n248) );
  XNOR U419 ( .A(n249), .B(n248), .Z(n250) );
  XOR U420 ( .A(in[1206]), .B(n250), .Z(n1374) );
  XOR U421 ( .A(in[1397]), .B(in[117]), .Z(n252) );
  XNOR U422 ( .A(in[1077]), .B(in[757]), .Z(n251) );
  XNOR U423 ( .A(n252), .B(n251), .Z(n253) );
  XOR U424 ( .A(in[437]), .B(n253), .Z(n1432) );
  XNOR U425 ( .A(n1374), .B(n1432), .Z(n3804) );
  XNOR U426 ( .A(in[182]), .B(n3804), .Z(n1346) );
  XOR U427 ( .A(in[151]), .B(in[1431]), .Z(n255) );
  XNOR U428 ( .A(in[1111]), .B(in[791]), .Z(n254) );
  XNOR U429 ( .A(n255), .B(n254), .Z(n256) );
  XOR U430 ( .A(in[471]), .B(n256), .Z(n563) );
  XOR U431 ( .A(in[342]), .B(in[662]), .Z(n258) );
  XNOR U432 ( .A(in[22]), .B(in[1302]), .Z(n257) );
  XNOR U433 ( .A(n258), .B(n257), .Z(n259) );
  XNOR U434 ( .A(in[982]), .B(n259), .Z(n1254) );
  XNOR U435 ( .A(n563), .B(n1254), .Z(n4132) );
  XNOR U436 ( .A(in[1367]), .B(n4132), .Z(n1741) );
  XOR U437 ( .A(in[1375]), .B(in[735]), .Z(n261) );
  XNOR U438 ( .A(in[95]), .B(in[415]), .Z(n260) );
  XNOR U439 ( .A(n261), .B(n260), .Z(n262) );
  XOR U440 ( .A(in[1055]), .B(n262), .Z(n929) );
  XOR U441 ( .A(in[1566]), .B(in[606]), .Z(n264) );
  XNOR U442 ( .A(in[926]), .B(in[286]), .Z(n263) );
  XNOR U443 ( .A(n264), .B(n263), .Z(n265) );
  XOR U444 ( .A(in[1246]), .B(n265), .Z(n665) );
  XNOR U445 ( .A(n929), .B(n665), .Z(n3906) );
  XNOR U446 ( .A(in[991]), .B(n3906), .Z(n1738) );
  NAND U447 ( .A(n1741), .B(n1738), .Z(n266) );
  XNOR U448 ( .A(n1346), .B(n266), .Z(out[1011]) );
  XOR U449 ( .A(in[1527]), .B(in[567]), .Z(n268) );
  XNOR U450 ( .A(in[887]), .B(in[247]), .Z(n267) );
  XNOR U451 ( .A(n268), .B(n267), .Z(n269) );
  XOR U452 ( .A(in[1207]), .B(n269), .Z(n1378) );
  XOR U453 ( .A(in[1398]), .B(in[118]), .Z(n271) );
  XNOR U454 ( .A(in[1078]), .B(in[758]), .Z(n270) );
  XNOR U455 ( .A(n271), .B(n270), .Z(n272) );
  XOR U456 ( .A(in[438]), .B(n272), .Z(n1436) );
  XNOR U457 ( .A(n1378), .B(n1436), .Z(n3808) );
  XNOR U458 ( .A(in[183]), .B(n3808), .Z(n1351) );
  XOR U459 ( .A(in[343]), .B(in[663]), .Z(n274) );
  XNOR U460 ( .A(in[23]), .B(in[1303]), .Z(n273) );
  XNOR U461 ( .A(n274), .B(n273), .Z(n275) );
  XOR U462 ( .A(in[983]), .B(n275), .Z(n1257) );
  XOR U463 ( .A(in[152]), .B(in[1432]), .Z(n277) );
  XNOR U464 ( .A(in[1112]), .B(in[792]), .Z(n276) );
  XNOR U465 ( .A(n277), .B(n276), .Z(n278) );
  XNOR U466 ( .A(in[472]), .B(n278), .Z(n589) );
  XNOR U467 ( .A(n1257), .B(n589), .Z(n4135) );
  XNOR U468 ( .A(in[1368]), .B(n4135), .Z(n1745) );
  XOR U469 ( .A(in[1376]), .B(in[736]), .Z(n280) );
  XNOR U470 ( .A(in[96]), .B(in[416]), .Z(n279) );
  XNOR U471 ( .A(n280), .B(n279), .Z(n281) );
  XOR U472 ( .A(in[1056]), .B(n281), .Z(n944) );
  XOR U473 ( .A(in[1567]), .B(in[607]), .Z(n283) );
  XNOR U474 ( .A(in[927]), .B(in[287]), .Z(n282) );
  XNOR U475 ( .A(n283), .B(n282), .Z(n284) );
  XOR U476 ( .A(in[1247]), .B(n284), .Z(n680) );
  XNOR U477 ( .A(n944), .B(n680), .Z(n3908) );
  XNOR U478 ( .A(in[992]), .B(n3908), .Z(n1742) );
  NAND U479 ( .A(n1745), .B(n1742), .Z(n285) );
  XNOR U480 ( .A(n1351), .B(n285), .Z(out[1012]) );
  XOR U481 ( .A(in[1528]), .B(in[568]), .Z(n287) );
  XNOR U482 ( .A(in[888]), .B(in[248]), .Z(n286) );
  XNOR U483 ( .A(n287), .B(n286), .Z(n288) );
  XOR U484 ( .A(in[1208]), .B(n288), .Z(n1382) );
  XOR U485 ( .A(in[1399]), .B(in[119]), .Z(n290) );
  XNOR U486 ( .A(in[1079]), .B(in[759]), .Z(n289) );
  XNOR U487 ( .A(n290), .B(n289), .Z(n291) );
  XOR U488 ( .A(in[439]), .B(n291), .Z(n1440) );
  XNOR U489 ( .A(n1382), .B(n1440), .Z(n3812) );
  XNOR U490 ( .A(in[184]), .B(n3812), .Z(n1355) );
  XOR U491 ( .A(in[344]), .B(in[664]), .Z(n293) );
  XNOR U492 ( .A(in[24]), .B(in[1304]), .Z(n292) );
  XNOR U493 ( .A(n293), .B(n292), .Z(n294) );
  XOR U494 ( .A(in[984]), .B(n294), .Z(n1260) );
  XOR U495 ( .A(in[153]), .B(in[1433]), .Z(n296) );
  XNOR U496 ( .A(in[1113]), .B(in[793]), .Z(n295) );
  XNOR U497 ( .A(n296), .B(n295), .Z(n297) );
  XNOR U498 ( .A(in[473]), .B(n297), .Z(n604) );
  XNOR U499 ( .A(n1260), .B(n604), .Z(n4138) );
  XNOR U500 ( .A(in[1369]), .B(n4138), .Z(n1749) );
  XOR U501 ( .A(in[1377]), .B(in[737]), .Z(n299) );
  XNOR U502 ( .A(in[97]), .B(in[417]), .Z(n298) );
  XNOR U503 ( .A(n299), .B(n298), .Z(n300) );
  XOR U504 ( .A(in[1057]), .B(n300), .Z(n959) );
  XOR U505 ( .A(in[1568]), .B(in[608]), .Z(n302) );
  XNOR U506 ( .A(in[928]), .B(in[288]), .Z(n301) );
  XNOR U507 ( .A(n302), .B(n301), .Z(n303) );
  XOR U508 ( .A(in[1248]), .B(n303), .Z(n695) );
  XNOR U509 ( .A(n959), .B(n695), .Z(n3910) );
  XNOR U510 ( .A(in[993]), .B(n3910), .Z(n1746) );
  NAND U511 ( .A(n1749), .B(n1746), .Z(n304) );
  XNOR U512 ( .A(n1355), .B(n304), .Z(out[1013]) );
  XOR U513 ( .A(in[1529]), .B(in[569]), .Z(n306) );
  XNOR U514 ( .A(in[889]), .B(in[249]), .Z(n305) );
  XNOR U515 ( .A(n306), .B(n305), .Z(n307) );
  XOR U516 ( .A(in[1209]), .B(n307), .Z(n1386) );
  XOR U517 ( .A(in[1400]), .B(in[120]), .Z(n309) );
  XNOR U518 ( .A(in[1080]), .B(in[760]), .Z(n308) );
  XNOR U519 ( .A(n309), .B(n308), .Z(n310) );
  XOR U520 ( .A(in[440]), .B(n310), .Z(n1444) );
  XNOR U521 ( .A(n1386), .B(n1444), .Z(n3816) );
  XNOR U522 ( .A(in[185]), .B(n3816), .Z(n1359) );
  XOR U523 ( .A(in[345]), .B(in[665]), .Z(n312) );
  XNOR U524 ( .A(in[25]), .B(in[1305]), .Z(n311) );
  XNOR U525 ( .A(n312), .B(n311), .Z(n313) );
  XOR U526 ( .A(in[985]), .B(n313), .Z(n1263) );
  XOR U527 ( .A(in[154]), .B(in[1434]), .Z(n315) );
  XNOR U528 ( .A(in[1114]), .B(in[794]), .Z(n314) );
  XNOR U529 ( .A(n315), .B(n314), .Z(n316) );
  XNOR U530 ( .A(in[474]), .B(n316), .Z(n619) );
  XNOR U531 ( .A(n1263), .B(n619), .Z(n4141) );
  XNOR U532 ( .A(in[1370]), .B(n4141), .Z(n1754) );
  XOR U533 ( .A(in[1569]), .B(in[609]), .Z(n318) );
  XNOR U534 ( .A(in[929]), .B(in[289]), .Z(n317) );
  XNOR U535 ( .A(n318), .B(n317), .Z(n319) );
  XOR U536 ( .A(in[1249]), .B(n319), .Z(n710) );
  XOR U537 ( .A(in[1378]), .B(in[738]), .Z(n321) );
  XNOR U538 ( .A(in[98]), .B(in[418]), .Z(n320) );
  XNOR U539 ( .A(n321), .B(n320), .Z(n322) );
  XOR U540 ( .A(in[1058]), .B(n322), .Z(n974) );
  XNOR U541 ( .A(n710), .B(n974), .Z(n3912) );
  XNOR U542 ( .A(in[994]), .B(n3912), .Z(n1751) );
  NAND U543 ( .A(n1754), .B(n1751), .Z(n323) );
  XNOR U544 ( .A(n1359), .B(n323), .Z(out[1014]) );
  XOR U545 ( .A(in[1401]), .B(in[121]), .Z(n325) );
  XNOR U546 ( .A(in[1081]), .B(in[761]), .Z(n324) );
  XNOR U547 ( .A(n325), .B(n324), .Z(n326) );
  XOR U548 ( .A(in[441]), .B(n326), .Z(n1448) );
  XNOR U549 ( .A(n327), .B(n1448), .Z(n3538) );
  XNOR U550 ( .A(in[186]), .B(n3538), .Z(n1363) );
  XOR U551 ( .A(in[155]), .B(in[1435]), .Z(n329) );
  XNOR U552 ( .A(in[1115]), .B(in[795]), .Z(n328) );
  XNOR U553 ( .A(n329), .B(n328), .Z(n330) );
  XOR U554 ( .A(in[475]), .B(n330), .Z(n634) );
  XOR U555 ( .A(in[346]), .B(in[666]), .Z(n332) );
  XNOR U556 ( .A(in[26]), .B(in[1306]), .Z(n331) );
  XNOR U557 ( .A(n332), .B(n331), .Z(n333) );
  XNOR U558 ( .A(in[986]), .B(n333), .Z(n1266) );
  XNOR U559 ( .A(n634), .B(n1266), .Z(n4148) );
  XNOR U560 ( .A(in[1371]), .B(n4148), .Z(n1758) );
  XOR U561 ( .A(in[1379]), .B(in[739]), .Z(n335) );
  XNOR U562 ( .A(in[99]), .B(in[419]), .Z(n334) );
  XNOR U563 ( .A(n335), .B(n334), .Z(n336) );
  XNOR U564 ( .A(in[1059]), .B(n336), .Z(n989) );
  XNOR U565 ( .A(n337), .B(n989), .Z(n3914) );
  XNOR U566 ( .A(in[995]), .B(n3914), .Z(n1755) );
  NAND U567 ( .A(n1758), .B(n1755), .Z(n338) );
  XNOR U568 ( .A(n1363), .B(n338), .Z(out[1015]) );
  XOR U569 ( .A(in[1402]), .B(in[122]), .Z(n340) );
  XNOR U570 ( .A(in[1082]), .B(in[762]), .Z(n339) );
  XNOR U571 ( .A(n340), .B(n339), .Z(n341) );
  XOR U572 ( .A(in[442]), .B(n341), .Z(n1452) );
  XOR U573 ( .A(in[1531]), .B(in[571]), .Z(n343) );
  XNOR U574 ( .A(in[1211]), .B(in[251]), .Z(n342) );
  XNOR U575 ( .A(n343), .B(n342), .Z(n344) );
  XOR U576 ( .A(in[891]), .B(n344), .Z(n416) );
  XNOR U577 ( .A(n1452), .B(n416), .Z(n3542) );
  XNOR U578 ( .A(in[187]), .B(n3542), .Z(n1367) );
  XOR U579 ( .A(in[156]), .B(in[1436]), .Z(n346) );
  XNOR U580 ( .A(in[1116]), .B(in[796]), .Z(n345) );
  XNOR U581 ( .A(n346), .B(n345), .Z(n347) );
  XOR U582 ( .A(in[476]), .B(n347), .Z(n649) );
  XOR U583 ( .A(in[347]), .B(in[667]), .Z(n349) );
  XNOR U584 ( .A(in[27]), .B(in[1307]), .Z(n348) );
  XNOR U585 ( .A(n349), .B(n348), .Z(n350) );
  XNOR U586 ( .A(in[987]), .B(n350), .Z(n1269) );
  XNOR U587 ( .A(n649), .B(n1269), .Z(n4151) );
  XNOR U588 ( .A(in[1372]), .B(n4151), .Z(n1762) );
  XOR U589 ( .A(in[1060]), .B(in[420]), .Z(n352) );
  XNOR U590 ( .A(in[740]), .B(in[1380]), .Z(n351) );
  XNOR U591 ( .A(n352), .B(n351), .Z(n353) );
  XOR U592 ( .A(in[100]), .B(n353), .Z(n1004) );
  XOR U593 ( .A(in[1571]), .B(in[611]), .Z(n355) );
  XNOR U594 ( .A(in[931]), .B(in[291]), .Z(n354) );
  XNOR U595 ( .A(n355), .B(n354), .Z(n356) );
  XOR U596 ( .A(in[1251]), .B(n356), .Z(n420) );
  XNOR U597 ( .A(n1004), .B(n420), .Z(n3916) );
  XNOR U598 ( .A(in[996]), .B(n3916), .Z(n1759) );
  NAND U599 ( .A(n1762), .B(n1759), .Z(n357) );
  XNOR U600 ( .A(n1367), .B(n357), .Z(out[1016]) );
  XOR U601 ( .A(in[1403]), .B(in[123]), .Z(n359) );
  XNOR U602 ( .A(in[1083]), .B(in[763]), .Z(n358) );
  XNOR U603 ( .A(n359), .B(n358), .Z(n360) );
  XOR U604 ( .A(in[443]), .B(n360), .Z(n1456) );
  XOR U605 ( .A(in[1532]), .B(in[572]), .Z(n362) );
  XNOR U606 ( .A(in[1212]), .B(in[252]), .Z(n361) );
  XNOR U607 ( .A(n362), .B(n361), .Z(n363) );
  XOR U608 ( .A(in[892]), .B(n363), .Z(n581) );
  XNOR U609 ( .A(n1456), .B(n581), .Z(n3546) );
  XNOR U610 ( .A(in[188]), .B(n3546), .Z(n1371) );
  XOR U611 ( .A(in[157]), .B(in[1437]), .Z(n365) );
  XNOR U612 ( .A(in[1117]), .B(in[797]), .Z(n364) );
  XNOR U613 ( .A(n365), .B(n364), .Z(n366) );
  XOR U614 ( .A(in[477]), .B(n366), .Z(n664) );
  XOR U615 ( .A(in[348]), .B(in[668]), .Z(n368) );
  XNOR U616 ( .A(in[28]), .B(in[1308]), .Z(n367) );
  XNOR U617 ( .A(n368), .B(n367), .Z(n369) );
  XNOR U618 ( .A(in[988]), .B(n369), .Z(n1272) );
  XNOR U619 ( .A(n664), .B(n1272), .Z(n4154) );
  XNOR U620 ( .A(in[1373]), .B(n4154), .Z(n1766) );
  XOR U621 ( .A(in[1572]), .B(in[612]), .Z(n371) );
  XNOR U622 ( .A(in[932]), .B(in[292]), .Z(n370) );
  XNOR U623 ( .A(n371), .B(n370), .Z(n372) );
  XOR U624 ( .A(in[1252]), .B(n372), .Z(n583) );
  XNOR U625 ( .A(n373), .B(n583), .Z(n3918) );
  XNOR U626 ( .A(in[997]), .B(n3918), .Z(n1763) );
  NAND U627 ( .A(n1766), .B(n1763), .Z(n374) );
  XNOR U628 ( .A(n1371), .B(n374), .Z(out[1017]) );
  XOR U629 ( .A(in[1404]), .B(in[124]), .Z(n376) );
  XNOR U630 ( .A(in[1084]), .B(in[764]), .Z(n375) );
  XNOR U631 ( .A(n376), .B(n375), .Z(n377) );
  XOR U632 ( .A(in[444]), .B(n377), .Z(n1460) );
  XOR U633 ( .A(in[1533]), .B(in[573]), .Z(n379) );
  XNOR U634 ( .A(in[1213]), .B(in[253]), .Z(n378) );
  XNOR U635 ( .A(n379), .B(n378), .Z(n380) );
  XOR U636 ( .A(in[893]), .B(n380), .Z(n740) );
  XNOR U637 ( .A(n1460), .B(n740), .Z(n3550) );
  XNOR U638 ( .A(in[189]), .B(n3550), .Z(n1375) );
  XOR U639 ( .A(in[158]), .B(in[1438]), .Z(n382) );
  XNOR U640 ( .A(in[1118]), .B(in[798]), .Z(n381) );
  XNOR U641 ( .A(n382), .B(n381), .Z(n383) );
  XOR U642 ( .A(in[478]), .B(n383), .Z(n679) );
  XOR U643 ( .A(in[349]), .B(in[669]), .Z(n385) );
  XNOR U644 ( .A(in[29]), .B(in[1309]), .Z(n384) );
  XNOR U645 ( .A(n385), .B(n384), .Z(n386) );
  XNOR U646 ( .A(in[989]), .B(n386), .Z(n1276) );
  XNOR U647 ( .A(n679), .B(n1276), .Z(n4157) );
  XNOR U648 ( .A(in[1374]), .B(n4157), .Z(n1770) );
  XOR U649 ( .A(in[1062]), .B(in[422]), .Z(n388) );
  XNOR U650 ( .A(in[742]), .B(in[1382]), .Z(n387) );
  XNOR U651 ( .A(n388), .B(n387), .Z(n389) );
  XOR U652 ( .A(in[102]), .B(n389), .Z(n424) );
  XOR U653 ( .A(in[1573]), .B(in[613]), .Z(n391) );
  XNOR U654 ( .A(in[933]), .B(in[293]), .Z(n390) );
  XNOR U655 ( .A(n391), .B(n390), .Z(n392) );
  XOR U656 ( .A(in[1253]), .B(n392), .Z(n742) );
  XNOR U657 ( .A(n424), .B(n742), .Z(n3924) );
  XNOR U658 ( .A(in[998]), .B(n3924), .Z(n1767) );
  NAND U659 ( .A(n1770), .B(n1767), .Z(n393) );
  XNOR U660 ( .A(n1375), .B(n393), .Z(out[1018]) );
  XOR U661 ( .A(in[1405]), .B(in[125]), .Z(n395) );
  XNOR U662 ( .A(in[1085]), .B(in[765]), .Z(n394) );
  XNOR U663 ( .A(n395), .B(n394), .Z(n396) );
  XOR U664 ( .A(in[445]), .B(n396), .Z(n1464) );
  XOR U665 ( .A(in[1534]), .B(in[894]), .Z(n398) );
  XNOR U666 ( .A(in[574]), .B(in[1214]), .Z(n397) );
  XNOR U667 ( .A(n398), .B(n397), .Z(n399) );
  XOR U668 ( .A(in[254]), .B(n399), .Z(n877) );
  XNOR U669 ( .A(n1464), .B(n877), .Z(n3554) );
  XNOR U670 ( .A(in[190]), .B(n3554), .Z(n1379) );
  XOR U671 ( .A(in[1439]), .B(in[479]), .Z(n401) );
  XNOR U672 ( .A(in[799]), .B(in[159]), .Z(n400) );
  XNOR U673 ( .A(n401), .B(n400), .Z(n402) );
  XOR U674 ( .A(in[1119]), .B(n402), .Z(n694) );
  XOR U675 ( .A(in[350]), .B(in[670]), .Z(n404) );
  XNOR U676 ( .A(in[30]), .B(in[1310]), .Z(n403) );
  XNOR U677 ( .A(n404), .B(n403), .Z(n405) );
  XNOR U678 ( .A(in[990]), .B(n405), .Z(n1279) );
  XNOR U679 ( .A(n694), .B(n1279), .Z(n4160) );
  XNOR U680 ( .A(in[1375]), .B(n4160), .Z(n1774) );
  XOR U681 ( .A(in[1063]), .B(in[423]), .Z(n407) );
  XNOR U682 ( .A(in[743]), .B(in[1383]), .Z(n406) );
  XNOR U683 ( .A(n407), .B(n406), .Z(n408) );
  XOR U684 ( .A(in[103]), .B(n408), .Z(n587) );
  XOR U685 ( .A(in[1574]), .B(in[614]), .Z(n410) );
  XNOR U686 ( .A(in[934]), .B(in[294]), .Z(n409) );
  XNOR U687 ( .A(n410), .B(n409), .Z(n411) );
  XOR U688 ( .A(in[1254]), .B(n411), .Z(n786) );
  XNOR U689 ( .A(n587), .B(n786), .Z(n3926) );
  XNOR U690 ( .A(in[999]), .B(n3926), .Z(n1771) );
  NAND U691 ( .A(n1774), .B(n1771), .Z(n412) );
  XNOR U692 ( .A(n1379), .B(n412), .Z(out[1019]) );
  XOR U693 ( .A(in[1340]), .B(in[60]), .Z(n414) );
  XNOR U694 ( .A(in[700]), .B(in[380]), .Z(n413) );
  XNOR U695 ( .A(n414), .B(n413), .Z(n415) );
  XOR U696 ( .A(in[1020]), .B(n415), .Z(n871) );
  XNOR U697 ( .A(n416), .B(n871), .Z(n3596) );
  XNOR U698 ( .A(in[636]), .B(n3596), .Z(n2552) );
  XOR U699 ( .A(in[162]), .B(in[1442]), .Z(n418) );
  XNOR U700 ( .A(in[802]), .B(in[1122]), .Z(n417) );
  XNOR U701 ( .A(n418), .B(n417), .Z(n419) );
  XNOR U702 ( .A(in[482]), .B(n419), .Z(n471) );
  XNOR U703 ( .A(n420), .B(n471), .Z(n3693) );
  XNOR U704 ( .A(in[227]), .B(n3693), .Z(n2845) );
  XOR U705 ( .A(in[1511]), .B(in[551]), .Z(n422) );
  XNOR U706 ( .A(in[871]), .B(in[231]), .Z(n421) );
  XNOR U707 ( .A(n422), .B(n421), .Z(n423) );
  XOR U708 ( .A(in[1191]), .B(n423), .Z(n1313) );
  XNOR U709 ( .A(n424), .B(n1313), .Z(n3734) );
  XNOR U710 ( .A(in[1447]), .B(n3734), .Z(n2842) );
  NAND U711 ( .A(n2845), .B(n2842), .Z(n425) );
  XNOR U712 ( .A(n2552), .B(n425), .Z(out[101]) );
  XOR U713 ( .A(in[1406]), .B(in[126]), .Z(n427) );
  XNOR U714 ( .A(in[1086]), .B(in[766]), .Z(n426) );
  XNOR U715 ( .A(n427), .B(n426), .Z(n428) );
  XOR U716 ( .A(in[446]), .B(n428), .Z(n1469) );
  XOR U717 ( .A(in[1535]), .B(in[575]), .Z(n430) );
  XNOR U718 ( .A(in[895]), .B(in[255]), .Z(n429) );
  XNOR U719 ( .A(n430), .B(n429), .Z(n431) );
  XOR U720 ( .A(in[1215]), .B(n431), .Z(n1024) );
  XNOR U721 ( .A(n1469), .B(n1024), .Z(n3558) );
  XNOR U722 ( .A(in[191]), .B(n3558), .Z(n1383) );
  XOR U723 ( .A(in[1440]), .B(in[480]), .Z(n433) );
  XNOR U724 ( .A(in[800]), .B(in[160]), .Z(n432) );
  XNOR U725 ( .A(n433), .B(n432), .Z(n434) );
  XOR U726 ( .A(in[1120]), .B(n434), .Z(n709) );
  XOR U727 ( .A(in[351]), .B(in[671]), .Z(n436) );
  XNOR U728 ( .A(in[31]), .B(in[1311]), .Z(n435) );
  XNOR U729 ( .A(n436), .B(n435), .Z(n437) );
  XNOR U730 ( .A(in[991]), .B(n437), .Z(n1282) );
  XNOR U731 ( .A(n709), .B(n1282), .Z(n4163) );
  XNOR U732 ( .A(in[1376]), .B(n4163), .Z(n1778) );
  XOR U733 ( .A(in[1064]), .B(in[424]), .Z(n439) );
  XNOR U734 ( .A(in[744]), .B(in[1384]), .Z(n438) );
  XNOR U735 ( .A(n439), .B(n438), .Z(n440) );
  XOR U736 ( .A(in[104]), .B(n440), .Z(n746) );
  XOR U737 ( .A(in[1575]), .B(in[615]), .Z(n442) );
  XNOR U738 ( .A(in[935]), .B(in[295]), .Z(n441) );
  XNOR U739 ( .A(n442), .B(n441), .Z(n443) );
  XOR U740 ( .A(in[1255]), .B(n443), .Z(n799) );
  XNOR U741 ( .A(n746), .B(n799), .Z(n3928) );
  XNOR U742 ( .A(in[1000]), .B(n3928), .Z(n1775) );
  NAND U743 ( .A(n1778), .B(n1775), .Z(n444) );
  XNOR U744 ( .A(n1383), .B(n444), .Z(out[1020]) );
  XOR U745 ( .A(in[1407]), .B(in[127]), .Z(n446) );
  XNOR U746 ( .A(in[1087]), .B(in[767]), .Z(n445) );
  XNOR U747 ( .A(n446), .B(n445), .Z(n447) );
  XOR U748 ( .A(in[447]), .B(n447), .Z(n1472) );
  XOR U749 ( .A(in[1472]), .B(in[512]), .Z(n449) );
  XNOR U750 ( .A(in[832]), .B(in[192]), .Z(n448) );
  XNOR U751 ( .A(n449), .B(n448), .Z(n450) );
  XOR U752 ( .A(in[1152]), .B(n450), .Z(n1091) );
  XNOR U753 ( .A(n1472), .B(n1091), .Z(n3562) );
  XNOR U754 ( .A(in[128]), .B(n3562), .Z(n1387) );
  XOR U755 ( .A(in[352]), .B(in[672]), .Z(n452) );
  XNOR U756 ( .A(in[32]), .B(in[1312]), .Z(n451) );
  XNOR U757 ( .A(n452), .B(n451), .Z(n453) );
  XNOR U758 ( .A(in[992]), .B(n453), .Z(n1285) );
  XNOR U759 ( .A(n454), .B(n1285), .Z(n4166) );
  XNOR U760 ( .A(in[1377]), .B(n4166), .Z(n1782) );
  XOR U761 ( .A(in[1065]), .B(in[425]), .Z(n456) );
  XNOR U762 ( .A(in[745]), .B(in[1385]), .Z(n455) );
  XNOR U763 ( .A(n456), .B(n455), .Z(n457) );
  XOR U764 ( .A(in[105]), .B(n457), .Z(n881) );
  XOR U765 ( .A(in[1576]), .B(in[616]), .Z(n459) );
  XNOR U766 ( .A(in[936]), .B(in[296]), .Z(n458) );
  XNOR U767 ( .A(n459), .B(n458), .Z(n460) );
  XOR U768 ( .A(in[1256]), .B(n460), .Z(n812) );
  XNOR U769 ( .A(n881), .B(n812), .Z(n3930) );
  XNOR U770 ( .A(in[1001]), .B(n3930), .Z(n1779) );
  NAND U771 ( .A(n1782), .B(n1779), .Z(n461) );
  XNOR U772 ( .A(n1387), .B(n461), .Z(out[1021]) );
  XOR U773 ( .A(in[1344]), .B(in[64]), .Z(n463) );
  XNOR U774 ( .A(in[1024]), .B(in[384]), .Z(n462) );
  XNOR U775 ( .A(n463), .B(n462), .Z(n464) );
  XOR U776 ( .A(in[704]), .B(n464), .Z(n1477) );
  XOR U777 ( .A(in[1473]), .B(in[513]), .Z(n466) );
  XNOR U778 ( .A(in[833]), .B(in[193]), .Z(n465) );
  XNOR U779 ( .A(n466), .B(n465), .Z(n467) );
  XOR U780 ( .A(in[1153]), .B(n467), .Z(n1144) );
  XNOR U781 ( .A(n1477), .B(n1144), .Z(n3566) );
  XNOR U782 ( .A(in[129]), .B(n3566), .Z(n1390) );
  XOR U783 ( .A(in[353]), .B(in[673]), .Z(n469) );
  XNOR U784 ( .A(in[33]), .B(in[1313]), .Z(n468) );
  XNOR U785 ( .A(n469), .B(n468), .Z(n470) );
  XOR U786 ( .A(in[993]), .B(n470), .Z(n1288) );
  XNOR U787 ( .A(n1288), .B(n471), .Z(n4169) );
  XNOR U788 ( .A(in[1378]), .B(n4169), .Z(n1786) );
  XOR U789 ( .A(in[1577]), .B(in[617]), .Z(n473) );
  XNOR U790 ( .A(in[937]), .B(in[297]), .Z(n472) );
  XNOR U791 ( .A(n473), .B(n472), .Z(n474) );
  XOR U792 ( .A(in[1257]), .B(n474), .Z(n825) );
  XNOR U793 ( .A(n475), .B(n825), .Z(n3932) );
  XNOR U794 ( .A(in[1002]), .B(n3932), .Z(n1783) );
  NAND U795 ( .A(n1786), .B(n1783), .Z(n476) );
  XNOR U796 ( .A(n1390), .B(n476), .Z(out[1022]) );
  XOR U797 ( .A(n3570), .B(in[130]), .Z(n1392) );
  XOR U798 ( .A(in[163]), .B(in[1443]), .Z(n478) );
  XNOR U799 ( .A(in[803]), .B(in[1123]), .Z(n477) );
  XNOR U800 ( .A(n478), .B(n477), .Z(n479) );
  XOR U801 ( .A(in[483]), .B(n479), .Z(n582) );
  XOR U802 ( .A(in[354]), .B(in[674]), .Z(n481) );
  XNOR U803 ( .A(in[34]), .B(in[1314]), .Z(n480) );
  XNOR U804 ( .A(n481), .B(n480), .Z(n482) );
  XNOR U805 ( .A(in[994]), .B(n482), .Z(n1291) );
  XNOR U806 ( .A(n582), .B(n1291), .Z(n4172) );
  XNOR U807 ( .A(in[1379]), .B(n4172), .Z(n1790) );
  XOR U808 ( .A(in[1578]), .B(in[618]), .Z(n484) );
  XNOR U809 ( .A(in[938]), .B(in[298]), .Z(n483) );
  XNOR U810 ( .A(n484), .B(n483), .Z(n485) );
  XOR U811 ( .A(in[1258]), .B(n485), .Z(n838) );
  XNOR U812 ( .A(n486), .B(n838), .Z(n3934) );
  XNOR U813 ( .A(in[1003]), .B(n3934), .Z(n1787) );
  NAND U814 ( .A(n1790), .B(n1787), .Z(n487) );
  XNOR U815 ( .A(n1392), .B(n487), .Z(out[1023]) );
  XNOR U816 ( .A(n489), .B(n488), .Z(n3625) );
  XNOR U817 ( .A(in[531]), .B(n3625), .Z(n1396) );
  XOR U818 ( .A(in[1346]), .B(in[66]), .Z(n491) );
  XNOR U819 ( .A(in[1026]), .B(in[386]), .Z(n490) );
  XNOR U820 ( .A(n491), .B(n490), .Z(n492) );
  XOR U821 ( .A(in[706]), .B(n492), .Z(n1485) );
  XOR U822 ( .A(in[1475]), .B(in[515]), .Z(n494) );
  XNOR U823 ( .A(in[835]), .B(in[195]), .Z(n493) );
  XNOR U824 ( .A(n494), .B(n493), .Z(n495) );
  XNOR U825 ( .A(in[1155]), .B(n495), .Z(n1196) );
  XNOR U826 ( .A(n1485), .B(n1196), .Z(n3574) );
  XNOR U827 ( .A(in[131]), .B(n3574), .Z(n4631) );
  XOR U828 ( .A(in[35]), .B(in[675]), .Z(n497) );
  XNOR U829 ( .A(in[355]), .B(in[1315]), .Z(n496) );
  XNOR U830 ( .A(n497), .B(n496), .Z(n498) );
  XOR U831 ( .A(in[995]), .B(n498), .Z(n1294) );
  XOR U832 ( .A(in[164]), .B(in[1444]), .Z(n500) );
  XNOR U833 ( .A(in[804]), .B(in[1124]), .Z(n499) );
  XNOR U834 ( .A(n500), .B(n499), .Z(n501) );
  XOR U835 ( .A(in[484]), .B(n501), .Z(n741) );
  XNOR U836 ( .A(n1294), .B(n741), .Z(n4175) );
  XNOR U837 ( .A(in[1380]), .B(n4175), .Z(n4628) );
  NAND U838 ( .A(n4631), .B(n4628), .Z(n502) );
  XNOR U839 ( .A(n1396), .B(n502), .Z(out[1024]) );
  XNOR U840 ( .A(n504), .B(n503), .Z(n3629) );
  XNOR U841 ( .A(in[532]), .B(n3629), .Z(n1400) );
  XOR U842 ( .A(in[1347]), .B(in[67]), .Z(n506) );
  XNOR U843 ( .A(in[1027]), .B(in[387]), .Z(n505) );
  XNOR U844 ( .A(n506), .B(n505), .Z(n507) );
  XOR U845 ( .A(in[707]), .B(n507), .Z(n1489) );
  XOR U846 ( .A(in[1476]), .B(in[516]), .Z(n509) );
  XNOR U847 ( .A(in[836]), .B(in[196]), .Z(n508) );
  XNOR U848 ( .A(n509), .B(n508), .Z(n510) );
  XNOR U849 ( .A(in[1156]), .B(n510), .Z(n1199) );
  XNOR U850 ( .A(n1489), .B(n1199), .Z(n3582) );
  XNOR U851 ( .A(in[132]), .B(n3582), .Z(n4635) );
  XOR U852 ( .A(in[36]), .B(in[676]), .Z(n512) );
  XNOR U853 ( .A(in[356]), .B(in[1316]), .Z(n511) );
  XNOR U854 ( .A(n512), .B(n511), .Z(n513) );
  XOR U855 ( .A(in[996]), .B(n513), .Z(n1297) );
  XOR U856 ( .A(in[1445]), .B(in[165]), .Z(n515) );
  XNOR U857 ( .A(in[805]), .B(in[1125]), .Z(n514) );
  XNOR U858 ( .A(n515), .B(n514), .Z(n516) );
  XOR U859 ( .A(in[485]), .B(n516), .Z(n785) );
  XNOR U860 ( .A(n1297), .B(n785), .Z(n4182) );
  XNOR U861 ( .A(in[1381]), .B(n4182), .Z(n4632) );
  NAND U862 ( .A(n4635), .B(n4632), .Z(n517) );
  XNOR U863 ( .A(n1400), .B(n517), .Z(out[1025]) );
  XOR U864 ( .A(n519), .B(n518), .Z(n3633) );
  XNOR U865 ( .A(in[533]), .B(n3633), .Z(n1404) );
  XOR U866 ( .A(in[1348]), .B(in[68]), .Z(n521) );
  XNOR U867 ( .A(in[1028]), .B(in[388]), .Z(n520) );
  XNOR U868 ( .A(n521), .B(n520), .Z(n522) );
  XOR U869 ( .A(in[708]), .B(n522), .Z(n1493) );
  XOR U870 ( .A(in[1477]), .B(in[517]), .Z(n524) );
  XNOR U871 ( .A(in[837]), .B(in[197]), .Z(n523) );
  XNOR U872 ( .A(n524), .B(n523), .Z(n525) );
  XNOR U873 ( .A(in[1157]), .B(n525), .Z(n1202) );
  XNOR U874 ( .A(n1493), .B(n1202), .Z(n3586) );
  XNOR U875 ( .A(in[133]), .B(n3586), .Z(n4639) );
  XOR U876 ( .A(in[166]), .B(in[806]), .Z(n527) );
  XNOR U877 ( .A(in[1126]), .B(in[486]), .Z(n526) );
  XNOR U878 ( .A(n527), .B(n526), .Z(n528) );
  XOR U879 ( .A(in[1446]), .B(n528), .Z(n798) );
  XOR U880 ( .A(in[37]), .B(in[677]), .Z(n530) );
  XNOR U881 ( .A(in[357]), .B(in[1317]), .Z(n529) );
  XNOR U882 ( .A(n530), .B(n529), .Z(n531) );
  XOR U883 ( .A(in[997]), .B(n531), .Z(n1300) );
  XNOR U884 ( .A(n798), .B(n1300), .Z(n4185) );
  XNOR U885 ( .A(in[1382]), .B(n4185), .Z(n4636) );
  NAND U886 ( .A(n4639), .B(n4636), .Z(n532) );
  XNOR U887 ( .A(n1404), .B(n532), .Z(out[1026]) );
  XNOR U888 ( .A(n534), .B(n533), .Z(n3637) );
  XNOR U889 ( .A(in[534]), .B(n3637), .Z(n1408) );
  XOR U890 ( .A(in[1349]), .B(in[69]), .Z(n536) );
  XNOR U891 ( .A(in[1029]), .B(in[389]), .Z(n535) );
  XNOR U892 ( .A(n536), .B(n535), .Z(n537) );
  XOR U893 ( .A(in[709]), .B(n537), .Z(n1497) );
  XOR U894 ( .A(in[1478]), .B(in[518]), .Z(n539) );
  XNOR U895 ( .A(in[838]), .B(in[198]), .Z(n538) );
  XNOR U896 ( .A(n539), .B(n538), .Z(n540) );
  XNOR U897 ( .A(in[1158]), .B(n540), .Z(n1205) );
  XNOR U898 ( .A(n1497), .B(n1205), .Z(n3590) );
  XNOR U899 ( .A(in[134]), .B(n3590), .Z(n4643) );
  XOR U900 ( .A(in[38]), .B(in[678]), .Z(n542) );
  XNOR U901 ( .A(in[358]), .B(in[1318]), .Z(n541) );
  XNOR U902 ( .A(n542), .B(n541), .Z(n543) );
  XOR U903 ( .A(in[998]), .B(n543), .Z(n1304) );
  XOR U904 ( .A(in[167]), .B(in[807]), .Z(n545) );
  XNOR U905 ( .A(in[1127]), .B(in[487]), .Z(n544) );
  XNOR U906 ( .A(n545), .B(n544), .Z(n546) );
  XOR U907 ( .A(in[1447]), .B(n546), .Z(n811) );
  XNOR U908 ( .A(n1304), .B(n811), .Z(n3964) );
  XNOR U909 ( .A(in[1383]), .B(n3964), .Z(n4640) );
  NAND U910 ( .A(n4643), .B(n4640), .Z(n547) );
  XNOR U911 ( .A(n1408), .B(n547), .Z(out[1027]) );
  XOR U912 ( .A(n549), .B(n548), .Z(n3641) );
  XNOR U913 ( .A(in[535]), .B(n3641), .Z(n1412) );
  XOR U914 ( .A(in[1350]), .B(in[70]), .Z(n551) );
  XNOR U915 ( .A(in[1030]), .B(in[390]), .Z(n550) );
  XNOR U916 ( .A(n551), .B(n550), .Z(n552) );
  XOR U917 ( .A(in[710]), .B(n552), .Z(n1501) );
  XOR U918 ( .A(in[199]), .B(in[1479]), .Z(n554) );
  XNOR U919 ( .A(in[1159]), .B(in[839]), .Z(n553) );
  XNOR U920 ( .A(n554), .B(n553), .Z(n555) );
  XNOR U921 ( .A(in[519]), .B(n555), .Z(n1208) );
  XNOR U922 ( .A(n1501), .B(n1208), .Z(n3594) );
  XNOR U923 ( .A(in[135]), .B(n3594), .Z(n4647) );
  XOR U924 ( .A(in[168]), .B(in[1448]), .Z(n557) );
  XNOR U925 ( .A(in[1128]), .B(in[808]), .Z(n556) );
  XNOR U926 ( .A(n557), .B(n556), .Z(n558) );
  XOR U927 ( .A(in[488]), .B(n558), .Z(n824) );
  XOR U928 ( .A(in[39]), .B(in[679]), .Z(n560) );
  XNOR U929 ( .A(in[359]), .B(in[1319]), .Z(n559) );
  XNOR U930 ( .A(n560), .B(n559), .Z(n561) );
  XOR U931 ( .A(in[999]), .B(n561), .Z(n1308) );
  XNOR U932 ( .A(n824), .B(n1308), .Z(n3967) );
  XNOR U933 ( .A(in[1384]), .B(n3967), .Z(n4644) );
  NAND U934 ( .A(n4647), .B(n4644), .Z(n562) );
  XNOR U935 ( .A(n1412), .B(n562), .Z(out[1028]) );
  XNOR U936 ( .A(n564), .B(n563), .Z(n3645) );
  XNOR U937 ( .A(in[536]), .B(n3645), .Z(n1416) );
  XOR U938 ( .A(in[1351]), .B(in[711]), .Z(n566) );
  XNOR U939 ( .A(in[1031]), .B(in[391]), .Z(n565) );
  XNOR U940 ( .A(n566), .B(n565), .Z(n567) );
  XOR U941 ( .A(in[71]), .B(n567), .Z(n1505) );
  XOR U942 ( .A(in[1480]), .B(in[520]), .Z(n569) );
  XNOR U943 ( .A(in[840]), .B(in[200]), .Z(n568) );
  XNOR U944 ( .A(n569), .B(n568), .Z(n570) );
  XNOR U945 ( .A(in[1160]), .B(n570), .Z(n1213) );
  XNOR U946 ( .A(n1505), .B(n1213), .Z(n3598) );
  XNOR U947 ( .A(in[136]), .B(n3598), .Z(n4651) );
  XOR U948 ( .A(in[169]), .B(in[1449]), .Z(n572) );
  XNOR U949 ( .A(in[1129]), .B(in[809]), .Z(n571) );
  XNOR U950 ( .A(n572), .B(n571), .Z(n573) );
  XOR U951 ( .A(in[489]), .B(n573), .Z(n837) );
  XOR U952 ( .A(in[680]), .B(in[1320]), .Z(n575) );
  XNOR U953 ( .A(in[40]), .B(in[360]), .Z(n574) );
  XNOR U954 ( .A(n575), .B(n574), .Z(n576) );
  XOR U955 ( .A(in[1000]), .B(n576), .Z(n1312) );
  XNOR U956 ( .A(n837), .B(n1312), .Z(n3974) );
  XNOR U957 ( .A(in[1385]), .B(n3974), .Z(n4648) );
  NAND U958 ( .A(n4651), .B(n4648), .Z(n577) );
  XNOR U959 ( .A(n1416), .B(n577), .Z(out[1029]) );
  XOR U960 ( .A(in[1341]), .B(in[61]), .Z(n579) );
  XNOR U961 ( .A(in[701]), .B(in[381]), .Z(n578) );
  XNOR U962 ( .A(n579), .B(n578), .Z(n580) );
  XOR U963 ( .A(in[1021]), .B(n580), .Z(n894) );
  XNOR U964 ( .A(n581), .B(n894), .Z(n3600) );
  XNOR U965 ( .A(in[637]), .B(n3600), .Z(n2555) );
  XOR U966 ( .A(n583), .B(n582), .Z(n3697) );
  XNOR U967 ( .A(in[228]), .B(n3697), .Z(n2859) );
  XOR U968 ( .A(in[1512]), .B(in[552]), .Z(n585) );
  XNOR U969 ( .A(in[872]), .B(in[232]), .Z(n584) );
  XNOR U970 ( .A(n585), .B(n584), .Z(n586) );
  XOR U971 ( .A(in[1192]), .B(n586), .Z(n1317) );
  XNOR U972 ( .A(n587), .B(n1317), .Z(n3738) );
  XNOR U973 ( .A(in[1448]), .B(n3738), .Z(n2856) );
  NAND U974 ( .A(n2859), .B(n2856), .Z(n588) );
  XNOR U975 ( .A(n2555), .B(n588), .Z(out[102]) );
  XOR U976 ( .A(n590), .B(n589), .Z(n3649) );
  XNOR U977 ( .A(in[537]), .B(n3649), .Z(n1420) );
  XOR U978 ( .A(in[1352]), .B(in[712]), .Z(n592) );
  XNOR U979 ( .A(in[1032]), .B(in[392]), .Z(n591) );
  XNOR U980 ( .A(n592), .B(n591), .Z(n593) );
  XOR U981 ( .A(in[72]), .B(n593), .Z(n1510) );
  XOR U982 ( .A(in[1481]), .B(in[521]), .Z(n595) );
  XNOR U983 ( .A(in[841]), .B(in[201]), .Z(n594) );
  XNOR U984 ( .A(n595), .B(n594), .Z(n596) );
  XNOR U985 ( .A(in[1161]), .B(n596), .Z(n1216) );
  XNOR U986 ( .A(n1510), .B(n1216), .Z(n3602) );
  XNOR U987 ( .A(in[137]), .B(n3602), .Z(n4655) );
  XOR U988 ( .A(in[170]), .B(in[1450]), .Z(n598) );
  XNOR U989 ( .A(in[1130]), .B(in[810]), .Z(n597) );
  XNOR U990 ( .A(n598), .B(n597), .Z(n599) );
  XOR U991 ( .A(in[490]), .B(n599), .Z(n853) );
  XOR U992 ( .A(in[681]), .B(in[1321]), .Z(n601) );
  XNOR U993 ( .A(in[41]), .B(in[361]), .Z(n600) );
  XNOR U994 ( .A(n601), .B(n600), .Z(n602) );
  XOR U995 ( .A(in[1001]), .B(n602), .Z(n1316) );
  XNOR U996 ( .A(n853), .B(n1316), .Z(n3977) );
  XNOR U997 ( .A(in[1386]), .B(n3977), .Z(n4652) );
  NAND U998 ( .A(n4655), .B(n4652), .Z(n603) );
  XNOR U999 ( .A(n1420), .B(n603), .Z(out[1030]) );
  XOR U1000 ( .A(n605), .B(n604), .Z(n3653) );
  XNOR U1001 ( .A(in[538]), .B(n3653), .Z(n1424) );
  XOR U1002 ( .A(in[1353]), .B(in[393]), .Z(n607) );
  XNOR U1003 ( .A(in[713]), .B(in[73]), .Z(n606) );
  XNOR U1004 ( .A(n607), .B(n606), .Z(n608) );
  XOR U1005 ( .A(in[1033]), .B(n608), .Z(n1514) );
  XOR U1006 ( .A(in[1482]), .B(in[522]), .Z(n610) );
  XNOR U1007 ( .A(in[842]), .B(in[202]), .Z(n609) );
  XNOR U1008 ( .A(n610), .B(n609), .Z(n611) );
  XNOR U1009 ( .A(in[1162]), .B(n611), .Z(n1219) );
  XNOR U1010 ( .A(n1514), .B(n1219), .Z(n3606) );
  XNOR U1011 ( .A(in[138]), .B(n3606), .Z(n4659) );
  XOR U1012 ( .A(in[811]), .B(in[491]), .Z(n613) );
  XNOR U1013 ( .A(in[1451]), .B(in[1131]), .Z(n612) );
  XNOR U1014 ( .A(n613), .B(n612), .Z(n614) );
  XOR U1015 ( .A(in[171]), .B(n614), .Z(n866) );
  XOR U1016 ( .A(in[682]), .B(in[1322]), .Z(n616) );
  XNOR U1017 ( .A(in[42]), .B(in[362]), .Z(n615) );
  XNOR U1018 ( .A(n616), .B(n615), .Z(n617) );
  XOR U1019 ( .A(in[1002]), .B(n617), .Z(n1321) );
  XNOR U1020 ( .A(n866), .B(n1321), .Z(n3980) );
  XNOR U1021 ( .A(in[1387]), .B(n3980), .Z(n4656) );
  NAND U1022 ( .A(n4659), .B(n4656), .Z(n618) );
  XNOR U1023 ( .A(n1424), .B(n618), .Z(out[1031]) );
  XOR U1024 ( .A(n620), .B(n619), .Z(n3657) );
  XNOR U1025 ( .A(in[539]), .B(n3657), .Z(n1429) );
  XOR U1026 ( .A(in[1354]), .B(in[714]), .Z(n622) );
  XNOR U1027 ( .A(in[74]), .B(in[394]), .Z(n621) );
  XNOR U1028 ( .A(n622), .B(n621), .Z(n623) );
  XOR U1029 ( .A(in[1034]), .B(n623), .Z(n1518) );
  XOR U1030 ( .A(in[1483]), .B(in[523]), .Z(n625) );
  XNOR U1031 ( .A(in[843]), .B(in[203]), .Z(n624) );
  XNOR U1032 ( .A(n625), .B(n624), .Z(n626) );
  XNOR U1033 ( .A(in[1163]), .B(n626), .Z(n1222) );
  XNOR U1034 ( .A(n1518), .B(n1222), .Z(n3610) );
  XNOR U1035 ( .A(n3610), .B(in[139]), .Z(n4663) );
  XOR U1036 ( .A(in[812]), .B(in[492]), .Z(n628) );
  XNOR U1037 ( .A(in[1452]), .B(in[1132]), .Z(n627) );
  XNOR U1038 ( .A(n628), .B(n627), .Z(n629) );
  XOR U1039 ( .A(in[172]), .B(n629), .Z(n886) );
  XOR U1040 ( .A(in[683]), .B(in[1323]), .Z(n631) );
  XNOR U1041 ( .A(in[43]), .B(in[363]), .Z(n630) );
  XNOR U1042 ( .A(n631), .B(n630), .Z(n632) );
  XOR U1043 ( .A(in[1003]), .B(n632), .Z(n1325) );
  XNOR U1044 ( .A(n886), .B(n1325), .Z(n3983) );
  XNOR U1045 ( .A(in[1388]), .B(n3983), .Z(n4660) );
  NAND U1046 ( .A(n4663), .B(n4660), .Z(n633) );
  XNOR U1047 ( .A(n1429), .B(n633), .Z(out[1032]) );
  XNOR U1048 ( .A(n635), .B(n634), .Z(n3661) );
  XNOR U1049 ( .A(in[540]), .B(n3661), .Z(n1433) );
  XOR U1050 ( .A(in[1355]), .B(in[715]), .Z(n637) );
  XNOR U1051 ( .A(in[1035]), .B(in[395]), .Z(n636) );
  XNOR U1052 ( .A(n637), .B(n636), .Z(n638) );
  XOR U1053 ( .A(in[75]), .B(n638), .Z(n1522) );
  XOR U1054 ( .A(in[1484]), .B(in[524]), .Z(n640) );
  XNOR U1055 ( .A(in[844]), .B(in[204]), .Z(n639) );
  XNOR U1056 ( .A(n640), .B(n639), .Z(n641) );
  XNOR U1057 ( .A(in[1164]), .B(n641), .Z(n1225) );
  XNOR U1058 ( .A(n1522), .B(n1225), .Z(n3614) );
  XNOR U1059 ( .A(in[140]), .B(n3614), .Z(n4667) );
  XOR U1060 ( .A(in[1324]), .B(in[44]), .Z(n643) );
  XNOR U1061 ( .A(in[684]), .B(in[364]), .Z(n642) );
  XNOR U1062 ( .A(n643), .B(n642), .Z(n644) );
  XOR U1063 ( .A(in[1004]), .B(n644), .Z(n1328) );
  XOR U1064 ( .A(in[813]), .B(in[493]), .Z(n646) );
  XNOR U1065 ( .A(in[1453]), .B(in[1133]), .Z(n645) );
  XNOR U1066 ( .A(n646), .B(n645), .Z(n647) );
  XOR U1067 ( .A(in[173]), .B(n647), .Z(n899) );
  XNOR U1068 ( .A(n1328), .B(n899), .Z(n3986) );
  XNOR U1069 ( .A(in[1389]), .B(n3986), .Z(n4664) );
  NAND U1070 ( .A(n4667), .B(n4664), .Z(n648) );
  XNOR U1071 ( .A(n1433), .B(n648), .Z(out[1033]) );
  XNOR U1072 ( .A(n650), .B(n649), .Z(n3669) );
  XNOR U1073 ( .A(in[541]), .B(n3669), .Z(n1437) );
  XOR U1074 ( .A(in[76]), .B(in[1036]), .Z(n652) );
  XNOR U1075 ( .A(in[716]), .B(in[396]), .Z(n651) );
  XNOR U1076 ( .A(n652), .B(n651), .Z(n653) );
  XOR U1077 ( .A(in[1356]), .B(n653), .Z(n1526) );
  XOR U1078 ( .A(in[1485]), .B(in[525]), .Z(n655) );
  XNOR U1079 ( .A(in[845]), .B(in[205]), .Z(n654) );
  XNOR U1080 ( .A(n655), .B(n654), .Z(n656) );
  XNOR U1081 ( .A(in[1165]), .B(n656), .Z(n1228) );
  XNOR U1082 ( .A(n1526), .B(n1228), .Z(n3618) );
  XNOR U1083 ( .A(in[141]), .B(n3618), .Z(n4675) );
  XOR U1084 ( .A(in[1325]), .B(in[45]), .Z(n658) );
  XNOR U1085 ( .A(in[685]), .B(in[365]), .Z(n657) );
  XNOR U1086 ( .A(n658), .B(n657), .Z(n659) );
  XOR U1087 ( .A(in[1005]), .B(n659), .Z(n1332) );
  XOR U1088 ( .A(in[814]), .B(in[494]), .Z(n661) );
  XNOR U1089 ( .A(in[1454]), .B(in[1134]), .Z(n660) );
  XNOR U1090 ( .A(n661), .B(n660), .Z(n662) );
  XOR U1091 ( .A(in[174]), .B(n662), .Z(n912) );
  XNOR U1092 ( .A(n1332), .B(n912), .Z(n3989) );
  XNOR U1093 ( .A(in[1390]), .B(n3989), .Z(n4672) );
  NAND U1094 ( .A(n4675), .B(n4672), .Z(n663) );
  XNOR U1095 ( .A(n1437), .B(n663), .Z(out[1034]) );
  XNOR U1096 ( .A(n665), .B(n664), .Z(n3673) );
  XNOR U1097 ( .A(in[542]), .B(n3673), .Z(n1441) );
  XOR U1098 ( .A(in[77]), .B(in[1037]), .Z(n667) );
  XNOR U1099 ( .A(in[717]), .B(in[397]), .Z(n666) );
  XNOR U1100 ( .A(n667), .B(n666), .Z(n668) );
  XOR U1101 ( .A(in[1357]), .B(n668), .Z(n1530) );
  XOR U1102 ( .A(in[1486]), .B(in[526]), .Z(n670) );
  XNOR U1103 ( .A(in[846]), .B(in[206]), .Z(n669) );
  XNOR U1104 ( .A(n670), .B(n669), .Z(n671) );
  XNOR U1105 ( .A(in[1166]), .B(n671), .Z(n1231) );
  XNOR U1106 ( .A(n1530), .B(n1231), .Z(n3626) );
  XNOR U1107 ( .A(in[142]), .B(n3626), .Z(n4679) );
  XOR U1108 ( .A(in[815]), .B(in[495]), .Z(n673) );
  XNOR U1109 ( .A(in[1455]), .B(in[1135]), .Z(n672) );
  XNOR U1110 ( .A(n673), .B(n672), .Z(n674) );
  XOR U1111 ( .A(in[175]), .B(n674), .Z(n925) );
  XOR U1112 ( .A(in[1326]), .B(in[46]), .Z(n676) );
  XNOR U1113 ( .A(in[686]), .B(in[366]), .Z(n675) );
  XNOR U1114 ( .A(n676), .B(n675), .Z(n677) );
  XOR U1115 ( .A(in[1006]), .B(n677), .Z(n1336) );
  XNOR U1116 ( .A(n925), .B(n1336), .Z(n3992) );
  XNOR U1117 ( .A(in[1391]), .B(n3992), .Z(n4676) );
  NAND U1118 ( .A(n4679), .B(n4676), .Z(n678) );
  XNOR U1119 ( .A(n1441), .B(n678), .Z(out[1035]) );
  XNOR U1120 ( .A(n680), .B(n679), .Z(n3677) );
  XNOR U1121 ( .A(in[543]), .B(n3677), .Z(n1445) );
  XOR U1122 ( .A(in[78]), .B(in[1038]), .Z(n682) );
  XNOR U1123 ( .A(in[718]), .B(in[398]), .Z(n681) );
  XNOR U1124 ( .A(n682), .B(n681), .Z(n683) );
  XOR U1125 ( .A(in[1358]), .B(n683), .Z(n1534) );
  XOR U1126 ( .A(in[1487]), .B(in[527]), .Z(n685) );
  XNOR U1127 ( .A(in[847]), .B(in[207]), .Z(n684) );
  XNOR U1128 ( .A(n685), .B(n684), .Z(n686) );
  XNOR U1129 ( .A(in[1167]), .B(n686), .Z(n1234) );
  XNOR U1130 ( .A(n1534), .B(n1234), .Z(n3630) );
  XNOR U1131 ( .A(in[143]), .B(n3630), .Z(n4683) );
  XOR U1132 ( .A(in[816]), .B(in[496]), .Z(n688) );
  XNOR U1133 ( .A(in[1456]), .B(in[1136]), .Z(n687) );
  XNOR U1134 ( .A(n688), .B(n687), .Z(n689) );
  XOR U1135 ( .A(in[176]), .B(n689), .Z(n940) );
  XOR U1136 ( .A(in[1327]), .B(in[47]), .Z(n691) );
  XNOR U1137 ( .A(in[687]), .B(in[367]), .Z(n690) );
  XNOR U1138 ( .A(n691), .B(n690), .Z(n692) );
  XOR U1139 ( .A(in[1007]), .B(n692), .Z(n1340) );
  XNOR U1140 ( .A(n940), .B(n1340), .Z(n3995) );
  XNOR U1141 ( .A(in[1392]), .B(n3995), .Z(n4680) );
  NAND U1142 ( .A(n4683), .B(n4680), .Z(n693) );
  XNOR U1143 ( .A(n1445), .B(n693), .Z(out[1036]) );
  XNOR U1144 ( .A(n695), .B(n694), .Z(n3681) );
  XNOR U1145 ( .A(in[544]), .B(n3681), .Z(n1449) );
  XOR U1146 ( .A(in[79]), .B(in[1039]), .Z(n697) );
  XNOR U1147 ( .A(in[719]), .B(in[399]), .Z(n696) );
  XNOR U1148 ( .A(n697), .B(n696), .Z(n698) );
  XOR U1149 ( .A(in[1359]), .B(n698), .Z(n1538) );
  XOR U1150 ( .A(in[1488]), .B(in[528]), .Z(n700) );
  XNOR U1151 ( .A(in[848]), .B(in[208]), .Z(n699) );
  XNOR U1152 ( .A(n700), .B(n699), .Z(n701) );
  XNOR U1153 ( .A(in[1168]), .B(n701), .Z(n1237) );
  XNOR U1154 ( .A(n1538), .B(n1237), .Z(n3634) );
  XNOR U1155 ( .A(in[144]), .B(n3634), .Z(n4687) );
  XOR U1156 ( .A(in[1328]), .B(in[48]), .Z(n703) );
  XNOR U1157 ( .A(in[688]), .B(in[368]), .Z(n702) );
  XNOR U1158 ( .A(n703), .B(n702), .Z(n704) );
  XOR U1159 ( .A(in[1008]), .B(n704), .Z(n1344) );
  XOR U1160 ( .A(in[817]), .B(in[497]), .Z(n706) );
  XNOR U1161 ( .A(in[1457]), .B(in[1137]), .Z(n705) );
  XNOR U1162 ( .A(n706), .B(n705), .Z(n707) );
  XOR U1163 ( .A(in[177]), .B(n707), .Z(n955) );
  XNOR U1164 ( .A(n1344), .B(n955), .Z(n3998) );
  XNOR U1165 ( .A(in[1393]), .B(n3998), .Z(n4684) );
  NAND U1166 ( .A(n4687), .B(n4684), .Z(n708) );
  XNOR U1167 ( .A(n1449), .B(n708), .Z(out[1037]) );
  XNOR U1168 ( .A(n710), .B(n709), .Z(n3685) );
  XNOR U1169 ( .A(in[545]), .B(n3685), .Z(n1453) );
  XOR U1170 ( .A(in[80]), .B(in[1040]), .Z(n712) );
  XNOR U1171 ( .A(in[720]), .B(in[400]), .Z(n711) );
  XNOR U1172 ( .A(n712), .B(n711), .Z(n713) );
  XOR U1173 ( .A(in[1360]), .B(n713), .Z(n1542) );
  XOR U1174 ( .A(in[1489]), .B(in[529]), .Z(n715) );
  XNOR U1175 ( .A(in[849]), .B(in[209]), .Z(n714) );
  XNOR U1176 ( .A(n715), .B(n714), .Z(n716) );
  XNOR U1177 ( .A(in[1169]), .B(n716), .Z(n1240) );
  XNOR U1178 ( .A(n1542), .B(n1240), .Z(n3638) );
  XNOR U1179 ( .A(in[145]), .B(n3638), .Z(n4691) );
  XOR U1180 ( .A(in[818]), .B(in[498]), .Z(n718) );
  XNOR U1181 ( .A(in[1458]), .B(in[1138]), .Z(n717) );
  XNOR U1182 ( .A(n718), .B(n717), .Z(n719) );
  XOR U1183 ( .A(in[178]), .B(n719), .Z(n970) );
  XOR U1184 ( .A(in[1329]), .B(in[49]), .Z(n721) );
  XNOR U1185 ( .A(in[689]), .B(in[369]), .Z(n720) );
  XNOR U1186 ( .A(n721), .B(n720), .Z(n722) );
  XOR U1187 ( .A(in[1009]), .B(n722), .Z(n1349) );
  XNOR U1188 ( .A(n970), .B(n1349), .Z(n4001) );
  XNOR U1189 ( .A(in[1394]), .B(n4001), .Z(n4688) );
  NAND U1190 ( .A(n4691), .B(n4688), .Z(n723) );
  XNOR U1191 ( .A(n1453), .B(n723), .Z(out[1038]) );
  XOR U1192 ( .A(n3689), .B(in[546]), .Z(n1457) );
  XOR U1193 ( .A(in[81]), .B(in[1041]), .Z(n725) );
  XNOR U1194 ( .A(in[721]), .B(in[401]), .Z(n724) );
  XNOR U1195 ( .A(n725), .B(n724), .Z(n726) );
  XOR U1196 ( .A(in[1361]), .B(n726), .Z(n1546) );
  XOR U1197 ( .A(in[1490]), .B(in[530]), .Z(n728) );
  XNOR U1198 ( .A(in[850]), .B(in[210]), .Z(n727) );
  XNOR U1199 ( .A(n728), .B(n727), .Z(n729) );
  XNOR U1200 ( .A(in[1170]), .B(n729), .Z(n1244) );
  XNOR U1201 ( .A(n1546), .B(n1244), .Z(n3642) );
  XNOR U1202 ( .A(in[146]), .B(n3642), .Z(n4695) );
  XOR U1203 ( .A(in[819]), .B(in[499]), .Z(n731) );
  XNOR U1204 ( .A(in[1459]), .B(in[1139]), .Z(n730) );
  XNOR U1205 ( .A(n731), .B(n730), .Z(n732) );
  XOR U1206 ( .A(in[179]), .B(n732), .Z(n985) );
  XOR U1207 ( .A(in[1330]), .B(in[50]), .Z(n734) );
  XNOR U1208 ( .A(in[690]), .B(in[370]), .Z(n733) );
  XNOR U1209 ( .A(n734), .B(n733), .Z(n735) );
  XOR U1210 ( .A(in[1010]), .B(n735), .Z(n1353) );
  XNOR U1211 ( .A(n985), .B(n1353), .Z(n4008) );
  XNOR U1212 ( .A(in[1395]), .B(n4008), .Z(n4692) );
  NAND U1213 ( .A(n4695), .B(n4692), .Z(n736) );
  XNOR U1214 ( .A(n1457), .B(n736), .Z(out[1039]) );
  XOR U1215 ( .A(in[1342]), .B(in[62]), .Z(n738) );
  XNOR U1216 ( .A(in[702]), .B(in[382]), .Z(n737) );
  XNOR U1217 ( .A(n738), .B(n737), .Z(n739) );
  XOR U1218 ( .A(in[1022]), .B(n739), .Z(n907) );
  XNOR U1219 ( .A(n740), .B(n907), .Z(n3604) );
  XNOR U1220 ( .A(in[638]), .B(n3604), .Z(n2557) );
  XOR U1221 ( .A(n742), .B(n741), .Z(n3701) );
  XNOR U1222 ( .A(in[229]), .B(n3701), .Z(n2873) );
  XOR U1223 ( .A(in[1513]), .B(in[553]), .Z(n744) );
  XNOR U1224 ( .A(in[873]), .B(in[233]), .Z(n743) );
  XNOR U1225 ( .A(n744), .B(n743), .Z(n745) );
  XOR U1226 ( .A(in[1193]), .B(n745), .Z(n1320) );
  XNOR U1227 ( .A(n746), .B(n1320), .Z(n3742) );
  XNOR U1228 ( .A(in[1449]), .B(n3742), .Z(n2870) );
  NAND U1229 ( .A(n2873), .B(n2870), .Z(n747) );
  XNOR U1230 ( .A(n2557), .B(n747), .Z(out[103]) );
  XOR U1231 ( .A(n3693), .B(in[547]), .Z(n1461) );
  XOR U1232 ( .A(in[1042]), .B(in[402]), .Z(n749) );
  XNOR U1233 ( .A(in[722]), .B(in[82]), .Z(n748) );
  XNOR U1234 ( .A(n749), .B(n748), .Z(n750) );
  XOR U1235 ( .A(in[1362]), .B(n750), .Z(n1551) );
  XOR U1236 ( .A(in[851]), .B(in[1171]), .Z(n752) );
  XNOR U1237 ( .A(in[1491]), .B(in[211]), .Z(n751) );
  XNOR U1238 ( .A(n752), .B(n751), .Z(n753) );
  XNOR U1239 ( .A(in[531]), .B(n753), .Z(n1247) );
  XNOR U1240 ( .A(n1551), .B(n1247), .Z(n3646) );
  XNOR U1241 ( .A(in[147]), .B(n3646), .Z(n4699) );
  XOR U1242 ( .A(in[820]), .B(in[500]), .Z(n755) );
  XNOR U1243 ( .A(in[1460]), .B(in[1140]), .Z(n754) );
  XNOR U1244 ( .A(n755), .B(n754), .Z(n756) );
  XOR U1245 ( .A(in[180]), .B(n756), .Z(n1000) );
  XOR U1246 ( .A(in[1331]), .B(in[51]), .Z(n758) );
  XNOR U1247 ( .A(in[691]), .B(in[371]), .Z(n757) );
  XNOR U1248 ( .A(n758), .B(n757), .Z(n759) );
  XOR U1249 ( .A(in[1011]), .B(n759), .Z(n1357) );
  XNOR U1250 ( .A(n1000), .B(n1357), .Z(n4011) );
  XNOR U1251 ( .A(in[1396]), .B(n4011), .Z(n4696) );
  NAND U1252 ( .A(n4699), .B(n4696), .Z(n760) );
  XNOR U1253 ( .A(n1461), .B(n760), .Z(out[1040]) );
  XOR U1254 ( .A(n3697), .B(in[548]), .Z(n1465) );
  XOR U1255 ( .A(in[83]), .B(in[1043]), .Z(n762) );
  XNOR U1256 ( .A(in[723]), .B(in[403]), .Z(n761) );
  XNOR U1257 ( .A(n762), .B(n761), .Z(n763) );
  XOR U1258 ( .A(in[1363]), .B(n763), .Z(n1555) );
  XOR U1259 ( .A(in[852]), .B(in[1172]), .Z(n765) );
  XNOR U1260 ( .A(in[1492]), .B(in[212]), .Z(n764) );
  XNOR U1261 ( .A(n765), .B(n764), .Z(n766) );
  XNOR U1262 ( .A(in[532]), .B(n766), .Z(n1250) );
  XNOR U1263 ( .A(n1555), .B(n1250), .Z(n3650) );
  XNOR U1264 ( .A(in[148]), .B(n3650), .Z(n4703) );
  XOR U1265 ( .A(in[821]), .B(in[501]), .Z(n768) );
  XNOR U1266 ( .A(in[1461]), .B(in[1141]), .Z(n767) );
  XNOR U1267 ( .A(n768), .B(n767), .Z(n769) );
  XOR U1268 ( .A(in[181]), .B(n769), .Z(n1015) );
  XOR U1269 ( .A(in[1332]), .B(in[52]), .Z(n771) );
  XNOR U1270 ( .A(in[692]), .B(in[372]), .Z(n770) );
  XNOR U1271 ( .A(n771), .B(n770), .Z(n772) );
  XOR U1272 ( .A(in[1012]), .B(n772), .Z(n1361) );
  XNOR U1273 ( .A(n1015), .B(n1361), .Z(n4014) );
  XNOR U1274 ( .A(in[1397]), .B(n4014), .Z(n4700) );
  NAND U1275 ( .A(n4703), .B(n4700), .Z(n773) );
  XNOR U1276 ( .A(n1465), .B(n773), .Z(out[1041]) );
  XOR U1277 ( .A(n3701), .B(in[549]), .Z(n1470) );
  XOR U1278 ( .A(in[853]), .B(in[1173]), .Z(n775) );
  XNOR U1279 ( .A(in[1493]), .B(in[213]), .Z(n774) );
  XNOR U1280 ( .A(n775), .B(n774), .Z(n776) );
  XNOR U1281 ( .A(in[533]), .B(n776), .Z(n1253) );
  XNOR U1282 ( .A(n777), .B(n1253), .Z(n3654) );
  XNOR U1283 ( .A(in[149]), .B(n3654), .Z(n4707) );
  XOR U1284 ( .A(in[1333]), .B(in[53]), .Z(n779) );
  XNOR U1285 ( .A(in[693]), .B(in[373]), .Z(n778) );
  XNOR U1286 ( .A(n779), .B(n778), .Z(n780) );
  XOR U1287 ( .A(in[1013]), .B(n780), .Z(n1365) );
  XOR U1288 ( .A(in[822]), .B(in[502]), .Z(n782) );
  XNOR U1289 ( .A(in[1462]), .B(in[1142]), .Z(n781) );
  XNOR U1290 ( .A(n782), .B(n781), .Z(n783) );
  XOR U1291 ( .A(in[182]), .B(n783), .Z(n1029) );
  XNOR U1292 ( .A(n1365), .B(n1029), .Z(n4017) );
  XNOR U1293 ( .A(in[1398]), .B(n4017), .Z(n4704) );
  NAND U1294 ( .A(n4707), .B(n4704), .Z(n784) );
  XNOR U1295 ( .A(n1470), .B(n784), .Z(out[1042]) );
  XNOR U1296 ( .A(n786), .B(n785), .Z(n3705) );
  XNOR U1297 ( .A(in[550]), .B(n3705), .Z(n1474) );
  XOR U1298 ( .A(in[854]), .B(in[1174]), .Z(n788) );
  XNOR U1299 ( .A(in[1494]), .B(in[214]), .Z(n787) );
  XNOR U1300 ( .A(n788), .B(n787), .Z(n789) );
  XNOR U1301 ( .A(in[534]), .B(n789), .Z(n1256) );
  XNOR U1302 ( .A(n790), .B(n1256), .Z(n3658) );
  XNOR U1303 ( .A(in[150]), .B(n3658), .Z(n4711) );
  XOR U1304 ( .A(in[1334]), .B(in[54]), .Z(n792) );
  XNOR U1305 ( .A(in[694]), .B(in[374]), .Z(n791) );
  XNOR U1306 ( .A(n792), .B(n791), .Z(n793) );
  XOR U1307 ( .A(in[1014]), .B(n793), .Z(n1369) );
  XOR U1308 ( .A(in[823]), .B(in[503]), .Z(n795) );
  XNOR U1309 ( .A(in[1463]), .B(in[1143]), .Z(n794) );
  XNOR U1310 ( .A(n795), .B(n794), .Z(n796) );
  XOR U1311 ( .A(in[183]), .B(n796), .Z(n1040) );
  XNOR U1312 ( .A(n1369), .B(n1040), .Z(n4020) );
  XNOR U1313 ( .A(in[1399]), .B(n4020), .Z(n4708) );
  NAND U1314 ( .A(n4711), .B(n4708), .Z(n797) );
  XNOR U1315 ( .A(n1474), .B(n797), .Z(out[1043]) );
  XNOR U1316 ( .A(n799), .B(n798), .Z(n3713) );
  XNOR U1317 ( .A(in[551]), .B(n3713), .Z(n1478) );
  XOR U1318 ( .A(in[855]), .B(in[1175]), .Z(n801) );
  XNOR U1319 ( .A(in[1495]), .B(in[215]), .Z(n800) );
  XNOR U1320 ( .A(n801), .B(n800), .Z(n802) );
  XNOR U1321 ( .A(in[535]), .B(n802), .Z(n1259) );
  XNOR U1322 ( .A(n803), .B(n1259), .Z(n3662) );
  XNOR U1323 ( .A(in[151]), .B(n3662), .Z(n4719) );
  XOR U1324 ( .A(in[824]), .B(in[504]), .Z(n805) );
  XNOR U1325 ( .A(in[1464]), .B(in[1144]), .Z(n804) );
  XNOR U1326 ( .A(n805), .B(n804), .Z(n806) );
  XOR U1327 ( .A(in[184]), .B(n806), .Z(n1045) );
  XOR U1328 ( .A(in[1335]), .B(in[55]), .Z(n808) );
  XNOR U1329 ( .A(in[695]), .B(in[375]), .Z(n807) );
  XNOR U1330 ( .A(n808), .B(n807), .Z(n809) );
  XOR U1331 ( .A(in[1015]), .B(n809), .Z(n1373) );
  XNOR U1332 ( .A(n1045), .B(n1373), .Z(n4023) );
  XNOR U1333 ( .A(in[1400]), .B(n4023), .Z(n4716) );
  NAND U1334 ( .A(n4719), .B(n4716), .Z(n810) );
  XNOR U1335 ( .A(n1478), .B(n810), .Z(out[1044]) );
  XNOR U1336 ( .A(n812), .B(n811), .Z(n3717) );
  XNOR U1337 ( .A(in[552]), .B(n3717), .Z(n1482) );
  XOR U1338 ( .A(in[856]), .B(in[1176]), .Z(n814) );
  XNOR U1339 ( .A(in[1496]), .B(in[216]), .Z(n813) );
  XNOR U1340 ( .A(n814), .B(n813), .Z(n815) );
  XNOR U1341 ( .A(in[536]), .B(n815), .Z(n1262) );
  XNOR U1342 ( .A(n816), .B(n1262), .Z(n3670) );
  XNOR U1343 ( .A(in[152]), .B(n3670), .Z(n4723) );
  XOR U1344 ( .A(in[825]), .B(in[505]), .Z(n818) );
  XNOR U1345 ( .A(in[1465]), .B(in[1145]), .Z(n817) );
  XNOR U1346 ( .A(n818), .B(n817), .Z(n819) );
  XOR U1347 ( .A(in[185]), .B(n819), .Z(n1056) );
  XOR U1348 ( .A(in[1336]), .B(in[56]), .Z(n821) );
  XNOR U1349 ( .A(in[696]), .B(in[376]), .Z(n820) );
  XNOR U1350 ( .A(n821), .B(n820), .Z(n822) );
  XOR U1351 ( .A(in[1016]), .B(n822), .Z(n1377) );
  XNOR U1352 ( .A(n1056), .B(n1377), .Z(n4026) );
  XNOR U1353 ( .A(in[1401]), .B(n4026), .Z(n4720) );
  NAND U1354 ( .A(n4723), .B(n4720), .Z(n823) );
  XNOR U1355 ( .A(n1482), .B(n823), .Z(out[1045]) );
  XNOR U1356 ( .A(n825), .B(n824), .Z(n3721) );
  XNOR U1357 ( .A(in[553]), .B(n3721), .Z(n1486) );
  XOR U1358 ( .A(in[857]), .B(in[1177]), .Z(n827) );
  XNOR U1359 ( .A(in[1497]), .B(in[217]), .Z(n826) );
  XNOR U1360 ( .A(n827), .B(n826), .Z(n828) );
  XNOR U1361 ( .A(in[537]), .B(n828), .Z(n1265) );
  XNOR U1362 ( .A(n829), .B(n1265), .Z(n3674) );
  XNOR U1363 ( .A(in[153]), .B(n3674), .Z(n4727) );
  XOR U1364 ( .A(in[1337]), .B(in[57]), .Z(n831) );
  XNOR U1365 ( .A(in[697]), .B(in[377]), .Z(n830) );
  XNOR U1366 ( .A(n831), .B(n830), .Z(n832) );
  XOR U1367 ( .A(in[1017]), .B(n832), .Z(n1381) );
  XOR U1368 ( .A(in[826]), .B(in[506]), .Z(n834) );
  XNOR U1369 ( .A(in[1466]), .B(in[1146]), .Z(n833) );
  XNOR U1370 ( .A(n834), .B(n833), .Z(n835) );
  XOR U1371 ( .A(in[186]), .B(n835), .Z(n1067) );
  XNOR U1372 ( .A(n1381), .B(n1067), .Z(n4029) );
  XNOR U1373 ( .A(in[1402]), .B(n4029), .Z(n4724) );
  NAND U1374 ( .A(n4727), .B(n4724), .Z(n836) );
  XNOR U1375 ( .A(n1486), .B(n836), .Z(out[1046]) );
  XNOR U1376 ( .A(n838), .B(n837), .Z(n3725) );
  XNOR U1377 ( .A(in[554]), .B(n3725), .Z(n1490) );
  XOR U1378 ( .A(in[858]), .B(in[1178]), .Z(n840) );
  XNOR U1379 ( .A(in[1498]), .B(in[218]), .Z(n839) );
  XNOR U1380 ( .A(n840), .B(n839), .Z(n841) );
  XNOR U1381 ( .A(in[538]), .B(n841), .Z(n1268) );
  XNOR U1382 ( .A(n842), .B(n1268), .Z(n3678) );
  XNOR U1383 ( .A(in[154]), .B(n3678), .Z(n4731) );
  XOR U1384 ( .A(in[1338]), .B(in[58]), .Z(n844) );
  XNOR U1385 ( .A(in[698]), .B(in[378]), .Z(n843) );
  XNOR U1386 ( .A(n844), .B(n843), .Z(n845) );
  XOR U1387 ( .A(in[1018]), .B(n845), .Z(n1385) );
  XOR U1388 ( .A(in[827]), .B(in[507]), .Z(n847) );
  XNOR U1389 ( .A(in[1467]), .B(in[1147]), .Z(n846) );
  XNOR U1390 ( .A(n847), .B(n846), .Z(n848) );
  XOR U1391 ( .A(in[187]), .B(n848), .Z(n1072) );
  XNOR U1392 ( .A(n1385), .B(n1072), .Z(n4032) );
  XNOR U1393 ( .A(in[1403]), .B(n4032), .Z(n4728) );
  NAND U1394 ( .A(n4731), .B(n4728), .Z(n849) );
  XNOR U1395 ( .A(n1490), .B(n849), .Z(out[1047]) );
  XOR U1396 ( .A(in[1579]), .B(in[619]), .Z(n851) );
  XNOR U1397 ( .A(in[939]), .B(in[299]), .Z(n850) );
  XNOR U1398 ( .A(n851), .B(n850), .Z(n852) );
  XOR U1399 ( .A(in[1259]), .B(n852), .Z(n1394) );
  XNOR U1400 ( .A(n853), .B(n1394), .Z(n3729) );
  XNOR U1401 ( .A(in[555]), .B(n3729), .Z(n1494) );
  XOR U1402 ( .A(in[859]), .B(in[1179]), .Z(n855) );
  XNOR U1403 ( .A(in[1499]), .B(in[219]), .Z(n854) );
  XNOR U1404 ( .A(n855), .B(n854), .Z(n856) );
  XNOR U1405 ( .A(in[539]), .B(n856), .Z(n1271) );
  XNOR U1406 ( .A(n857), .B(n1271), .Z(n3682) );
  XNOR U1407 ( .A(in[155]), .B(n3682), .Z(n4735) );
  XOR U1408 ( .A(in[828]), .B(in[508]), .Z(n859) );
  XNOR U1409 ( .A(in[1468]), .B(in[1148]), .Z(n858) );
  XNOR U1410 ( .A(n859), .B(n858), .Z(n860) );
  XOR U1411 ( .A(in[188]), .B(n860), .Z(n1077) );
  XNOR U1412 ( .A(n861), .B(n1077), .Z(n4035) );
  XNOR U1413 ( .A(in[1404]), .B(n4035), .Z(n4732) );
  NAND U1414 ( .A(n4735), .B(n4732), .Z(n862) );
  XNOR U1415 ( .A(n1494), .B(n862), .Z(out[1048]) );
  XOR U1416 ( .A(in[1580]), .B(in[620]), .Z(n864) );
  XNOR U1417 ( .A(in[940]), .B(in[300]), .Z(n863) );
  XNOR U1418 ( .A(n864), .B(n863), .Z(n865) );
  XOR U1419 ( .A(in[1260]), .B(n865), .Z(n1398) );
  XNOR U1420 ( .A(n866), .B(n1398), .Z(n3733) );
  XNOR U1421 ( .A(in[556]), .B(n3733), .Z(n1498) );
  XOR U1422 ( .A(in[860]), .B(in[1180]), .Z(n868) );
  XNOR U1423 ( .A(in[1500]), .B(in[220]), .Z(n867) );
  XNOR U1424 ( .A(n868), .B(n867), .Z(n869) );
  XNOR U1425 ( .A(in[540]), .B(n869), .Z(n1275) );
  XNOR U1426 ( .A(n870), .B(n1275), .Z(n3686) );
  XNOR U1427 ( .A(in[156]), .B(n3686), .Z(n4739) );
  XNOR U1428 ( .A(n872), .B(n871), .Z(n4042) );
  XNOR U1429 ( .A(in[1405]), .B(n4042), .Z(n4736) );
  NAND U1430 ( .A(n4739), .B(n4736), .Z(n873) );
  XNOR U1431 ( .A(n1498), .B(n873), .Z(out[1049]) );
  XOR U1432 ( .A(in[1343]), .B(in[63]), .Z(n875) );
  XNOR U1433 ( .A(in[703]), .B(in[383]), .Z(n874) );
  XNOR U1434 ( .A(n875), .B(n874), .Z(n876) );
  XOR U1435 ( .A(in[1023]), .B(n876), .Z(n920) );
  XNOR U1436 ( .A(n877), .B(n920), .Z(n3608) );
  XNOR U1437 ( .A(in[639]), .B(n3608), .Z(n2559) );
  XOR U1438 ( .A(in[230]), .B(n3705), .Z(n2889) );
  XOR U1439 ( .A(in[874]), .B(in[1194]), .Z(n879) );
  XNOR U1440 ( .A(in[1514]), .B(in[234]), .Z(n878) );
  XNOR U1441 ( .A(n879), .B(n878), .Z(n880) );
  XOR U1442 ( .A(in[554]), .B(n880), .Z(n1324) );
  XNOR U1443 ( .A(n881), .B(n1324), .Z(n3746) );
  XNOR U1444 ( .A(in[1450]), .B(n3746), .Z(n2886) );
  NAND U1445 ( .A(n2889), .B(n2886), .Z(n882) );
  XNOR U1446 ( .A(n2559), .B(n882), .Z(out[104]) );
  XOR U1447 ( .A(in[1581]), .B(in[621]), .Z(n884) );
  XNOR U1448 ( .A(in[941]), .B(in[301]), .Z(n883) );
  XNOR U1449 ( .A(n884), .B(n883), .Z(n885) );
  XOR U1450 ( .A(in[1261]), .B(n885), .Z(n1402) );
  XNOR U1451 ( .A(n886), .B(n1402), .Z(n3737) );
  XNOR U1452 ( .A(in[557]), .B(n3737), .Z(n1502) );
  XOR U1453 ( .A(in[861]), .B(in[1181]), .Z(n888) );
  XNOR U1454 ( .A(in[1501]), .B(in[221]), .Z(n887) );
  XNOR U1455 ( .A(n888), .B(n887), .Z(n889) );
  XNOR U1456 ( .A(in[541]), .B(n889), .Z(n1278) );
  XNOR U1457 ( .A(n890), .B(n1278), .Z(n3690) );
  XNOR U1458 ( .A(in[157]), .B(n3690), .Z(n4743) );
  XOR U1459 ( .A(in[830]), .B(in[510]), .Z(n892) );
  XNOR U1460 ( .A(in[1470]), .B(in[1150]), .Z(n891) );
  XNOR U1461 ( .A(n892), .B(n891), .Z(n893) );
  XOR U1462 ( .A(in[190]), .B(n893), .Z(n1083) );
  XNOR U1463 ( .A(n894), .B(n1083), .Z(n4045) );
  XNOR U1464 ( .A(in[1406]), .B(n4045), .Z(n4740) );
  NAND U1465 ( .A(n4743), .B(n4740), .Z(n895) );
  XNOR U1466 ( .A(n1502), .B(n895), .Z(out[1050]) );
  XOR U1467 ( .A(in[1582]), .B(in[622]), .Z(n897) );
  XNOR U1468 ( .A(in[942]), .B(in[302]), .Z(n896) );
  XNOR U1469 ( .A(n897), .B(n896), .Z(n898) );
  XOR U1470 ( .A(in[1262]), .B(n898), .Z(n1406) );
  XNOR U1471 ( .A(n899), .B(n1406), .Z(n3741) );
  XNOR U1472 ( .A(in[558]), .B(n3741), .Z(n1506) );
  XOR U1473 ( .A(in[862]), .B(in[1182]), .Z(n901) );
  XNOR U1474 ( .A(in[1502]), .B(in[222]), .Z(n900) );
  XNOR U1475 ( .A(n901), .B(n900), .Z(n902) );
  XNOR U1476 ( .A(in[542]), .B(n902), .Z(n1281) );
  XNOR U1477 ( .A(n903), .B(n1281), .Z(n3694) );
  XNOR U1478 ( .A(in[158]), .B(n3694), .Z(n4747) );
  XOR U1479 ( .A(in[831]), .B(in[511]), .Z(n905) );
  XNOR U1480 ( .A(in[1471]), .B(in[1151]), .Z(n904) );
  XNOR U1481 ( .A(n905), .B(n904), .Z(n906) );
  XOR U1482 ( .A(in[191]), .B(n906), .Z(n1088) );
  XNOR U1483 ( .A(n907), .B(n1088), .Z(n4048) );
  XNOR U1484 ( .A(in[1407]), .B(n4048), .Z(n4744) );
  NAND U1485 ( .A(n4747), .B(n4744), .Z(n908) );
  XNOR U1486 ( .A(n1506), .B(n908), .Z(out[1051]) );
  XOR U1487 ( .A(in[1583]), .B(in[623]), .Z(n910) );
  XNOR U1488 ( .A(in[943]), .B(in[303]), .Z(n909) );
  XNOR U1489 ( .A(n910), .B(n909), .Z(n911) );
  XOR U1490 ( .A(in[1263]), .B(n911), .Z(n1410) );
  XNOR U1491 ( .A(n912), .B(n1410), .Z(n3745) );
  XNOR U1492 ( .A(in[559]), .B(n3745), .Z(n1511) );
  XOR U1493 ( .A(in[863]), .B(in[1183]), .Z(n914) );
  XNOR U1494 ( .A(in[1503]), .B(in[223]), .Z(n913) );
  XNOR U1495 ( .A(n914), .B(n913), .Z(n915) );
  XNOR U1496 ( .A(in[543]), .B(n915), .Z(n1284) );
  XNOR U1497 ( .A(n916), .B(n1284), .Z(n3698) );
  XNOR U1498 ( .A(in[159]), .B(n3698), .Z(n4751) );
  XOR U1499 ( .A(in[768]), .B(in[1088]), .Z(n918) );
  XNOR U1500 ( .A(in[448]), .B(in[1408]), .Z(n917) );
  XNOR U1501 ( .A(n918), .B(n917), .Z(n919) );
  XOR U1502 ( .A(in[128]), .B(n919), .Z(n1096) );
  XNOR U1503 ( .A(n920), .B(n1096), .Z(n4051) );
  XNOR U1504 ( .A(in[1344]), .B(n4051), .Z(n4748) );
  NAND U1505 ( .A(n4751), .B(n4748), .Z(n921) );
  XNOR U1506 ( .A(n1511), .B(n921), .Z(out[1052]) );
  XOR U1507 ( .A(in[1584]), .B(in[624]), .Z(n923) );
  XNOR U1508 ( .A(in[944]), .B(in[304]), .Z(n922) );
  XNOR U1509 ( .A(n923), .B(n922), .Z(n924) );
  XOR U1510 ( .A(in[1264]), .B(n924), .Z(n1414) );
  XNOR U1511 ( .A(n925), .B(n1414), .Z(n3749) );
  XNOR U1512 ( .A(in[560]), .B(n3749), .Z(n1515) );
  XOR U1513 ( .A(in[224]), .B(in[864]), .Z(n927) );
  XNOR U1514 ( .A(in[1184]), .B(in[1504]), .Z(n926) );
  XNOR U1515 ( .A(n927), .B(n926), .Z(n928) );
  XNOR U1516 ( .A(in[544]), .B(n928), .Z(n1287) );
  XNOR U1517 ( .A(n929), .B(n1287), .Z(n3702) );
  XNOR U1518 ( .A(in[160]), .B(n3702), .Z(n4755) );
  XOR U1519 ( .A(in[1280]), .B(in[640]), .Z(n931) );
  XNOR U1520 ( .A(in[960]), .B(in[320]), .Z(n930) );
  XNOR U1521 ( .A(n931), .B(n930), .Z(n932) );
  XOR U1522 ( .A(in[0]), .B(n932), .Z(n1023) );
  XOR U1523 ( .A(in[769]), .B(in[1089]), .Z(n934) );
  XNOR U1524 ( .A(in[449]), .B(in[1409]), .Z(n933) );
  XNOR U1525 ( .A(n934), .B(n933), .Z(n935) );
  XOR U1526 ( .A(in[129]), .B(n935), .Z(n1101) );
  XNOR U1527 ( .A(n1023), .B(n1101), .Z(n4054) );
  XNOR U1528 ( .A(in[1345]), .B(n4054), .Z(n4752) );
  NAND U1529 ( .A(n4755), .B(n4752), .Z(n936) );
  XNOR U1530 ( .A(n1515), .B(n936), .Z(out[1053]) );
  XOR U1531 ( .A(in[1585]), .B(in[625]), .Z(n938) );
  XNOR U1532 ( .A(in[945]), .B(in[305]), .Z(n937) );
  XNOR U1533 ( .A(n938), .B(n937), .Z(n939) );
  XOR U1534 ( .A(in[1265]), .B(n939), .Z(n1418) );
  XNOR U1535 ( .A(n940), .B(n1418), .Z(n3757) );
  XNOR U1536 ( .A(in[561]), .B(n3757), .Z(n1519) );
  XOR U1537 ( .A(in[225]), .B(in[865]), .Z(n942) );
  XNOR U1538 ( .A(in[1185]), .B(in[1505]), .Z(n941) );
  XNOR U1539 ( .A(n942), .B(n941), .Z(n943) );
  XNOR U1540 ( .A(in[545]), .B(n943), .Z(n1290) );
  XNOR U1541 ( .A(n944), .B(n1290), .Z(n3706) );
  XNOR U1542 ( .A(in[161]), .B(n3706), .Z(n4763) );
  XOR U1543 ( .A(in[1090]), .B(in[450]), .Z(n946) );
  XNOR U1544 ( .A(in[130]), .B(in[770]), .Z(n945) );
  XNOR U1545 ( .A(n946), .B(n945), .Z(n947) );
  XOR U1546 ( .A(in[1410]), .B(n947), .Z(n1106) );
  XOR U1547 ( .A(in[1]), .B(in[641]), .Z(n949) );
  XNOR U1548 ( .A(in[961]), .B(in[321]), .Z(n948) );
  XNOR U1549 ( .A(n949), .B(n948), .Z(n950) );
  XOR U1550 ( .A(in[1281]), .B(n950), .Z(n1090) );
  XNOR U1551 ( .A(n1106), .B(n1090), .Z(n4057) );
  XNOR U1552 ( .A(in[1346]), .B(n4057), .Z(n4760) );
  NAND U1553 ( .A(n4763), .B(n4760), .Z(n951) );
  XNOR U1554 ( .A(n1519), .B(n951), .Z(out[1054]) );
  XOR U1555 ( .A(in[1586]), .B(in[626]), .Z(n953) );
  XNOR U1556 ( .A(in[946]), .B(in[306]), .Z(n952) );
  XNOR U1557 ( .A(n953), .B(n952), .Z(n954) );
  XOR U1558 ( .A(in[1266]), .B(n954), .Z(n1422) );
  XNOR U1559 ( .A(n955), .B(n1422), .Z(n3761) );
  XNOR U1560 ( .A(in[562]), .B(n3761), .Z(n1523) );
  XOR U1561 ( .A(in[1186]), .B(in[1506]), .Z(n957) );
  XNOR U1562 ( .A(in[546]), .B(in[866]), .Z(n956) );
  XNOR U1563 ( .A(n957), .B(n956), .Z(n958) );
  XNOR U1564 ( .A(in[226]), .B(n958), .Z(n1293) );
  XNOR U1565 ( .A(n959), .B(n1293), .Z(n3714) );
  XNOR U1566 ( .A(in[162]), .B(n3714), .Z(n4767) );
  XOR U1567 ( .A(in[2]), .B(in[642]), .Z(n961) );
  XNOR U1568 ( .A(in[962]), .B(in[322]), .Z(n960) );
  XNOR U1569 ( .A(n961), .B(n960), .Z(n962) );
  XOR U1570 ( .A(in[1282]), .B(n962), .Z(n1143) );
  XOR U1571 ( .A(in[771]), .B(in[1091]), .Z(n964) );
  XNOR U1572 ( .A(in[451]), .B(in[1411]), .Z(n963) );
  XNOR U1573 ( .A(n964), .B(n963), .Z(n965) );
  XOR U1574 ( .A(in[131]), .B(n965), .Z(n1111) );
  XNOR U1575 ( .A(n1143), .B(n1111), .Z(n4060) );
  XNOR U1576 ( .A(in[1347]), .B(n4060), .Z(n4764) );
  NAND U1577 ( .A(n4767), .B(n4764), .Z(n966) );
  XNOR U1578 ( .A(n1523), .B(n966), .Z(out[1055]) );
  XOR U1579 ( .A(in[1587]), .B(in[627]), .Z(n968) );
  XNOR U1580 ( .A(in[947]), .B(in[307]), .Z(n967) );
  XNOR U1581 ( .A(n968), .B(n967), .Z(n969) );
  XOR U1582 ( .A(in[1267]), .B(n969), .Z(n1427) );
  XNOR U1583 ( .A(n970), .B(n1427), .Z(n3765) );
  XNOR U1584 ( .A(in[563]), .B(n3765), .Z(n1527) );
  XOR U1585 ( .A(in[1187]), .B(in[1507]), .Z(n972) );
  XNOR U1586 ( .A(in[547]), .B(in[867]), .Z(n971) );
  XNOR U1587 ( .A(n972), .B(n971), .Z(n973) );
  XNOR U1588 ( .A(in[227]), .B(n973), .Z(n1296) );
  XNOR U1589 ( .A(n974), .B(n1296), .Z(n3718) );
  XNOR U1590 ( .A(in[163]), .B(n3718), .Z(n4771) );
  XOR U1591 ( .A(in[772]), .B(in[1092]), .Z(n976) );
  XNOR U1592 ( .A(in[452]), .B(in[1412]), .Z(n975) );
  XNOR U1593 ( .A(n976), .B(n975), .Z(n977) );
  XOR U1594 ( .A(in[132]), .B(n977), .Z(n1116) );
  XOR U1595 ( .A(in[323]), .B(in[643]), .Z(n979) );
  XNOR U1596 ( .A(in[963]), .B(in[3]), .Z(n978) );
  XNOR U1597 ( .A(n979), .B(n978), .Z(n980) );
  XOR U1598 ( .A(in[1283]), .B(n980), .Z(n1189) );
  XNOR U1599 ( .A(n1116), .B(n1189), .Z(n4063) );
  XNOR U1600 ( .A(in[1348]), .B(n4063), .Z(n4768) );
  NAND U1601 ( .A(n4771), .B(n4768), .Z(n981) );
  XNOR U1602 ( .A(n1527), .B(n981), .Z(out[1056]) );
  XOR U1603 ( .A(in[1588]), .B(in[628]), .Z(n983) );
  XNOR U1604 ( .A(in[948]), .B(in[308]), .Z(n982) );
  XNOR U1605 ( .A(n983), .B(n982), .Z(n984) );
  XOR U1606 ( .A(in[1268]), .B(n984), .Z(n1431) );
  XNOR U1607 ( .A(n985), .B(n1431), .Z(n3769) );
  XNOR U1608 ( .A(in[564]), .B(n3769), .Z(n1531) );
  XOR U1609 ( .A(in[1188]), .B(in[1508]), .Z(n987) );
  XNOR U1610 ( .A(in[548]), .B(in[868]), .Z(n986) );
  XNOR U1611 ( .A(n987), .B(n986), .Z(n988) );
  XOR U1612 ( .A(in[228]), .B(n988), .Z(n1299) );
  XNOR U1613 ( .A(n1299), .B(n989), .Z(n3722) );
  XNOR U1614 ( .A(in[164]), .B(n3722), .Z(n4775) );
  XOR U1615 ( .A(in[773]), .B(in[1093]), .Z(n991) );
  XNOR U1616 ( .A(in[453]), .B(in[1413]), .Z(n990) );
  XNOR U1617 ( .A(n991), .B(n990), .Z(n992) );
  XOR U1618 ( .A(in[133]), .B(n992), .Z(n1121) );
  XOR U1619 ( .A(in[324]), .B(in[644]), .Z(n994) );
  XNOR U1620 ( .A(in[964]), .B(in[4]), .Z(n993) );
  XNOR U1621 ( .A(n994), .B(n993), .Z(n995) );
  XOR U1622 ( .A(in[1284]), .B(n995), .Z(n1197) );
  XNOR U1623 ( .A(n1121), .B(n1197), .Z(n4066) );
  XNOR U1624 ( .A(in[1349]), .B(n4066), .Z(n4772) );
  NAND U1625 ( .A(n4775), .B(n4772), .Z(n996) );
  XNOR U1626 ( .A(n1531), .B(n996), .Z(out[1057]) );
  XOR U1627 ( .A(in[1589]), .B(in[629]), .Z(n998) );
  XNOR U1628 ( .A(in[949]), .B(in[309]), .Z(n997) );
  XNOR U1629 ( .A(n998), .B(n997), .Z(n999) );
  XOR U1630 ( .A(in[1269]), .B(n999), .Z(n1435) );
  XNOR U1631 ( .A(n1000), .B(n1435), .Z(n3773) );
  XNOR U1632 ( .A(in[565]), .B(n3773), .Z(n1535) );
  XOR U1633 ( .A(in[1189]), .B(in[1509]), .Z(n1002) );
  XNOR U1634 ( .A(in[549]), .B(in[869]), .Z(n1001) );
  XNOR U1635 ( .A(n1002), .B(n1001), .Z(n1003) );
  XNOR U1636 ( .A(in[229]), .B(n1003), .Z(n1303) );
  XNOR U1637 ( .A(n1004), .B(n1303), .Z(n3726) );
  XNOR U1638 ( .A(in[165]), .B(n3726), .Z(n4779) );
  XOR U1639 ( .A(in[774]), .B(in[1094]), .Z(n1006) );
  XNOR U1640 ( .A(in[454]), .B(in[1414]), .Z(n1005) );
  XNOR U1641 ( .A(n1006), .B(n1005), .Z(n1007) );
  XOR U1642 ( .A(in[134]), .B(n1007), .Z(n1126) );
  XOR U1643 ( .A(in[325]), .B(in[645]), .Z(n1009) );
  XNOR U1644 ( .A(in[965]), .B(in[5]), .Z(n1008) );
  XNOR U1645 ( .A(n1009), .B(n1008), .Z(n1010) );
  XOR U1646 ( .A(in[1285]), .B(n1010), .Z(n1200) );
  XNOR U1647 ( .A(n1126), .B(n1200), .Z(n4069) );
  XNOR U1648 ( .A(in[1350]), .B(n4069), .Z(n4776) );
  NAND U1649 ( .A(n4779), .B(n4776), .Z(n1011) );
  XNOR U1650 ( .A(n1535), .B(n1011), .Z(out[1058]) );
  XOR U1651 ( .A(in[1590]), .B(in[630]), .Z(n1013) );
  XNOR U1652 ( .A(in[950]), .B(in[310]), .Z(n1012) );
  XNOR U1653 ( .A(n1013), .B(n1012), .Z(n1014) );
  XOR U1654 ( .A(in[1270]), .B(n1014), .Z(n1439) );
  XNOR U1655 ( .A(n1015), .B(n1439), .Z(n3777) );
  XNOR U1656 ( .A(in[566]), .B(n3777), .Z(n1539) );
  XOR U1657 ( .A(in[166]), .B(n3730), .Z(n4783) );
  XOR U1658 ( .A(in[775]), .B(in[1095]), .Z(n1017) );
  XNOR U1659 ( .A(in[455]), .B(in[1415]), .Z(n1016) );
  XNOR U1660 ( .A(n1017), .B(n1016), .Z(n1018) );
  XOR U1661 ( .A(in[135]), .B(n1018), .Z(n1131) );
  XOR U1662 ( .A(in[326]), .B(in[6]), .Z(n1020) );
  XNOR U1663 ( .A(in[966]), .B(in[646]), .Z(n1019) );
  XNOR U1664 ( .A(n1020), .B(n1019), .Z(n1021) );
  XOR U1665 ( .A(in[1286]), .B(n1021), .Z(n1203) );
  XNOR U1666 ( .A(n1131), .B(n1203), .Z(n4080) );
  XNOR U1667 ( .A(in[1351]), .B(n4080), .Z(n4780) );
  NAND U1668 ( .A(n4783), .B(n4780), .Z(n1022) );
  XNOR U1669 ( .A(n1539), .B(n1022), .Z(out[1059]) );
  XNOR U1670 ( .A(n1024), .B(n1023), .Z(n3612) );
  XNOR U1671 ( .A(in[576]), .B(n3612), .Z(n2561) );
  XOR U1672 ( .A(in[231]), .B(n3713), .Z(n2903) );
  XNOR U1673 ( .A(in[1451]), .B(n3750), .Z(n2900) );
  NAND U1674 ( .A(n2903), .B(n2900), .Z(n1025) );
  XNOR U1675 ( .A(n2561), .B(n1025), .Z(out[105]) );
  XOR U1676 ( .A(in[1591]), .B(in[631]), .Z(n1027) );
  XNOR U1677 ( .A(in[951]), .B(in[311]), .Z(n1026) );
  XNOR U1678 ( .A(n1027), .B(n1026), .Z(n1028) );
  XOR U1679 ( .A(in[1271]), .B(n1028), .Z(n1443) );
  XNOR U1680 ( .A(n1029), .B(n1443), .Z(n3781) );
  XNOR U1681 ( .A(in[567]), .B(n3781), .Z(n1543) );
  XOR U1682 ( .A(in[167]), .B(n3734), .Z(n4787) );
  XOR U1683 ( .A(in[776]), .B(in[1096]), .Z(n1031) );
  XNOR U1684 ( .A(in[456]), .B(in[1416]), .Z(n1030) );
  XNOR U1685 ( .A(n1031), .B(n1030), .Z(n1032) );
  XOR U1686 ( .A(in[136]), .B(n1032), .Z(n1136) );
  XOR U1687 ( .A(in[327]), .B(in[7]), .Z(n1034) );
  XNOR U1688 ( .A(in[967]), .B(in[647]), .Z(n1033) );
  XNOR U1689 ( .A(n1034), .B(n1033), .Z(n1035) );
  XOR U1690 ( .A(in[1287]), .B(n1035), .Z(n1206) );
  XNOR U1691 ( .A(n1136), .B(n1206), .Z(n4083) );
  XNOR U1692 ( .A(in[1352]), .B(n4083), .Z(n4784) );
  NAND U1693 ( .A(n4787), .B(n4784), .Z(n1036) );
  XNOR U1694 ( .A(n1543), .B(n1036), .Z(out[1060]) );
  XOR U1695 ( .A(in[632]), .B(in[1592]), .Z(n1038) );
  XNOR U1696 ( .A(in[1272]), .B(in[312]), .Z(n1037) );
  XNOR U1697 ( .A(n1038), .B(n1037), .Z(n1039) );
  XOR U1698 ( .A(in[952]), .B(n1039), .Z(n1447) );
  XNOR U1699 ( .A(n1040), .B(n1447), .Z(n3785) );
  XNOR U1700 ( .A(in[568]), .B(n3785), .Z(n1547) );
  XOR U1701 ( .A(in[168]), .B(n3738), .Z(n4791) );
  XNOR U1702 ( .A(in[1353]), .B(n4086), .Z(n4788) );
  NAND U1703 ( .A(n4791), .B(n4788), .Z(n1041) );
  XNOR U1704 ( .A(n1547), .B(n1041), .Z(out[1061]) );
  XOR U1705 ( .A(in[633]), .B(in[1593]), .Z(n1043) );
  XNOR U1706 ( .A(in[1273]), .B(in[313]), .Z(n1042) );
  XNOR U1707 ( .A(n1043), .B(n1042), .Z(n1044) );
  XOR U1708 ( .A(in[953]), .B(n1044), .Z(n1451) );
  XNOR U1709 ( .A(n1045), .B(n1451), .Z(n3789) );
  XNOR U1710 ( .A(in[569]), .B(n3789), .Z(n1552) );
  XOR U1711 ( .A(in[169]), .B(n3742), .Z(n4795) );
  XOR U1712 ( .A(in[329]), .B(in[969]), .Z(n1047) );
  XNOR U1713 ( .A(in[9]), .B(in[649]), .Z(n1046) );
  XNOR U1714 ( .A(n1047), .B(n1046), .Z(n1048) );
  XOR U1715 ( .A(in[1289]), .B(n1048), .Z(n1214) );
  XOR U1716 ( .A(in[778]), .B(in[1098]), .Z(n1050) );
  XNOR U1717 ( .A(in[458]), .B(in[1418]), .Z(n1049) );
  XNOR U1718 ( .A(n1050), .B(n1049), .Z(n1051) );
  XOR U1719 ( .A(in[138]), .B(n1051), .Z(n1149) );
  XNOR U1720 ( .A(n1214), .B(n1149), .Z(n4089) );
  XNOR U1721 ( .A(in[1354]), .B(n4089), .Z(n4792) );
  NAND U1722 ( .A(n4795), .B(n4792), .Z(n1052) );
  XNOR U1723 ( .A(n1552), .B(n1052), .Z(out[1062]) );
  XOR U1724 ( .A(in[634]), .B(in[1594]), .Z(n1054) );
  XNOR U1725 ( .A(in[1274]), .B(in[314]), .Z(n1053) );
  XNOR U1726 ( .A(n1054), .B(n1053), .Z(n1055) );
  XOR U1727 ( .A(in[954]), .B(n1055), .Z(n1455) );
  XNOR U1728 ( .A(n1056), .B(n1455), .Z(n3793) );
  XNOR U1729 ( .A(in[570]), .B(n3793), .Z(n1556) );
  XOR U1730 ( .A(in[170]), .B(n3746), .Z(n4799) );
  XOR U1731 ( .A(in[1419]), .B(in[779]), .Z(n1058) );
  XNOR U1732 ( .A(in[1099]), .B(in[459]), .Z(n1057) );
  XNOR U1733 ( .A(n1058), .B(n1057), .Z(n1059) );
  XOR U1734 ( .A(in[139]), .B(n1059), .Z(n1154) );
  XOR U1735 ( .A(in[1290]), .B(in[650]), .Z(n1061) );
  XNOR U1736 ( .A(in[970]), .B(in[330]), .Z(n1060) );
  XNOR U1737 ( .A(n1061), .B(n1060), .Z(n1062) );
  XOR U1738 ( .A(in[10]), .B(n1062), .Z(n1217) );
  XNOR U1739 ( .A(n1154), .B(n1217), .Z(n4092) );
  XNOR U1740 ( .A(in[1355]), .B(n4092), .Z(n4796) );
  NAND U1741 ( .A(n4799), .B(n4796), .Z(n1063) );
  XNOR U1742 ( .A(n1556), .B(n1063), .Z(out[1063]) );
  XOR U1743 ( .A(in[955]), .B(in[1275]), .Z(n1065) );
  XNOR U1744 ( .A(in[1595]), .B(in[315]), .Z(n1064) );
  XNOR U1745 ( .A(n1065), .B(n1064), .Z(n1066) );
  XNOR U1746 ( .A(in[635]), .B(n1066), .Z(n1459) );
  XNOR U1747 ( .A(n1067), .B(n1459), .Z(n3803) );
  XNOR U1748 ( .A(in[571]), .B(n3803), .Z(n1558) );
  NOR U1749 ( .A(n1301), .B(n1696), .Z(n1068) );
  XNOR U1750 ( .A(n1558), .B(n1068), .Z(out[1064]) );
  XOR U1751 ( .A(in[956]), .B(in[1276]), .Z(n1070) );
  XNOR U1752 ( .A(in[1596]), .B(in[316]), .Z(n1069) );
  XNOR U1753 ( .A(n1070), .B(n1069), .Z(n1071) );
  XNOR U1754 ( .A(in[636]), .B(n1071), .Z(n1463) );
  XNOR U1755 ( .A(n1072), .B(n1463), .Z(n3807) );
  XNOR U1756 ( .A(in[572]), .B(n3807), .Z(n1560) );
  NOR U1757 ( .A(n1305), .B(n1700), .Z(n1073) );
  XNOR U1758 ( .A(n1560), .B(n1073), .Z(out[1065]) );
  XOR U1759 ( .A(in[957]), .B(in[1277]), .Z(n1075) );
  XNOR U1760 ( .A(in[1597]), .B(in[317]), .Z(n1074) );
  XNOR U1761 ( .A(n1075), .B(n1074), .Z(n1076) );
  XNOR U1762 ( .A(in[637]), .B(n1076), .Z(n1468) );
  XNOR U1763 ( .A(n1077), .B(n1468), .Z(n3811) );
  XNOR U1764 ( .A(in[573]), .B(n3811), .Z(n1562) );
  NOR U1765 ( .A(n1310), .B(n1704), .Z(n1078) );
  XNOR U1766 ( .A(n1562), .B(n1078), .Z(out[1066]) );
  XOR U1767 ( .A(in[574]), .B(n3815), .Z(n1564) );
  NOR U1768 ( .A(n1314), .B(n1708), .Z(n1079) );
  XNOR U1769 ( .A(n1564), .B(n1079), .Z(out[1067]) );
  XOR U1770 ( .A(in[959]), .B(in[1279]), .Z(n1081) );
  XNOR U1771 ( .A(in[1599]), .B(in[319]), .Z(n1080) );
  XNOR U1772 ( .A(n1081), .B(n1080), .Z(n1082) );
  XNOR U1773 ( .A(in[639]), .B(n1082), .Z(n1476) );
  XNOR U1774 ( .A(n1083), .B(n1476), .Z(n3537) );
  XNOR U1775 ( .A(in[575]), .B(n3537), .Z(n1566) );
  NOR U1776 ( .A(n1318), .B(n1713), .Z(n1084) );
  XNOR U1777 ( .A(n1566), .B(n1084), .Z(out[1068]) );
  XOR U1778 ( .A(in[896]), .B(in[1216]), .Z(n1086) );
  XNOR U1779 ( .A(in[1536]), .B(in[256]), .Z(n1085) );
  XNOR U1780 ( .A(n1086), .B(n1085), .Z(n1087) );
  XNOR U1781 ( .A(in[576]), .B(n1087), .Z(n1480) );
  XNOR U1782 ( .A(n1088), .B(n1480), .Z(n3541) );
  XNOR U1783 ( .A(in[512]), .B(n3541), .Z(n1568) );
  NOR U1784 ( .A(n1322), .B(n1717), .Z(n1089) );
  XNOR U1785 ( .A(n1568), .B(n1089), .Z(out[1069]) );
  XNOR U1786 ( .A(n1091), .B(n1090), .Z(n3616) );
  XNOR U1787 ( .A(in[577]), .B(n3616), .Z(n2563) );
  XOR U1788 ( .A(in[232]), .B(n3717), .Z(n2917) );
  XNOR U1789 ( .A(in[1452]), .B(n3758), .Z(n2914) );
  NAND U1790 ( .A(n2917), .B(n2914), .Z(n1092) );
  XNOR U1791 ( .A(n2563), .B(n1092), .Z(out[106]) );
  XOR U1792 ( .A(in[897]), .B(in[1217]), .Z(n1094) );
  XNOR U1793 ( .A(in[1537]), .B(in[257]), .Z(n1093) );
  XNOR U1794 ( .A(n1094), .B(n1093), .Z(n1095) );
  XNOR U1795 ( .A(in[577]), .B(n1095), .Z(n1484) );
  XNOR U1796 ( .A(n1096), .B(n1484), .Z(n3545) );
  XNOR U1797 ( .A(in[513]), .B(n3545), .Z(n1570) );
  NOR U1798 ( .A(n1326), .B(n1721), .Z(n1097) );
  XNOR U1799 ( .A(n1570), .B(n1097), .Z(out[1070]) );
  XOR U1800 ( .A(in[1538]), .B(in[578]), .Z(n1099) );
  XNOR U1801 ( .A(in[898]), .B(in[258]), .Z(n1098) );
  XNOR U1802 ( .A(n1099), .B(n1098), .Z(n1100) );
  XNOR U1803 ( .A(in[1218]), .B(n1100), .Z(n1488) );
  XNOR U1804 ( .A(n1101), .B(n1488), .Z(n3549) );
  XNOR U1805 ( .A(in[514]), .B(n3549), .Z(n1572) );
  NOR U1806 ( .A(n1330), .B(n1725), .Z(n1102) );
  XNOR U1807 ( .A(n1572), .B(n1102), .Z(out[1071]) );
  XOR U1808 ( .A(in[1539]), .B(in[579]), .Z(n1104) );
  XNOR U1809 ( .A(in[899]), .B(in[259]), .Z(n1103) );
  XNOR U1810 ( .A(n1104), .B(n1103), .Z(n1105) );
  XNOR U1811 ( .A(in[1219]), .B(n1105), .Z(n1492) );
  XNOR U1812 ( .A(n1106), .B(n1492), .Z(n3553) );
  XNOR U1813 ( .A(in[515]), .B(n3553), .Z(n1576) );
  NOR U1814 ( .A(n1334), .B(n1729), .Z(n1107) );
  XNOR U1815 ( .A(n1576), .B(n1107), .Z(out[1072]) );
  XOR U1816 ( .A(in[1540]), .B(in[580]), .Z(n1109) );
  XNOR U1817 ( .A(in[900]), .B(in[260]), .Z(n1108) );
  XNOR U1818 ( .A(n1109), .B(n1108), .Z(n1110) );
  XNOR U1819 ( .A(in[1220]), .B(n1110), .Z(n1496) );
  XNOR U1820 ( .A(n1111), .B(n1496), .Z(n3557) );
  XNOR U1821 ( .A(in[516]), .B(n3557), .Z(n1578) );
  NOR U1822 ( .A(n1338), .B(n1733), .Z(n1112) );
  XNOR U1823 ( .A(n1578), .B(n1112), .Z(out[1073]) );
  XOR U1824 ( .A(in[1541]), .B(in[581]), .Z(n1114) );
  XNOR U1825 ( .A(in[901]), .B(in[261]), .Z(n1113) );
  XNOR U1826 ( .A(n1114), .B(n1113), .Z(n1115) );
  XNOR U1827 ( .A(in[1221]), .B(n1115), .Z(n1500) );
  XNOR U1828 ( .A(n1116), .B(n1500), .Z(n3561) );
  XNOR U1829 ( .A(in[517]), .B(n3561), .Z(n1580) );
  NOR U1830 ( .A(n1342), .B(n1737), .Z(n1117) );
  XNOR U1831 ( .A(n1580), .B(n1117), .Z(out[1074]) );
  XOR U1832 ( .A(in[1542]), .B(in[582]), .Z(n1119) );
  XNOR U1833 ( .A(in[902]), .B(in[262]), .Z(n1118) );
  XNOR U1834 ( .A(n1119), .B(n1118), .Z(n1120) );
  XNOR U1835 ( .A(in[1222]), .B(n1120), .Z(n1504) );
  XNOR U1836 ( .A(n1121), .B(n1504), .Z(n3565) );
  XNOR U1837 ( .A(in[518]), .B(n3565), .Z(n1582) );
  NOR U1838 ( .A(n1346), .B(n1741), .Z(n1122) );
  XNOR U1839 ( .A(n1582), .B(n1122), .Z(out[1075]) );
  XOR U1840 ( .A(in[1543]), .B(in[583]), .Z(n1124) );
  XNOR U1841 ( .A(in[903]), .B(in[263]), .Z(n1123) );
  XNOR U1842 ( .A(n1124), .B(n1123), .Z(n1125) );
  XNOR U1843 ( .A(in[1223]), .B(n1125), .Z(n1509) );
  XNOR U1844 ( .A(n1126), .B(n1509), .Z(n3569) );
  XNOR U1845 ( .A(in[519]), .B(n3569), .Z(n1584) );
  NOR U1846 ( .A(n1351), .B(n1745), .Z(n1127) );
  XNOR U1847 ( .A(n1584), .B(n1127), .Z(out[1076]) );
  XOR U1848 ( .A(in[1544]), .B(in[584]), .Z(n1129) );
  XNOR U1849 ( .A(in[904]), .B(in[264]), .Z(n1128) );
  XNOR U1850 ( .A(n1129), .B(n1128), .Z(n1130) );
  XNOR U1851 ( .A(in[1224]), .B(n1130), .Z(n1513) );
  XNOR U1852 ( .A(n1131), .B(n1513), .Z(n3573) );
  XNOR U1853 ( .A(in[520]), .B(n3573), .Z(n1586) );
  NOR U1854 ( .A(n1355), .B(n1749), .Z(n1132) );
  XNOR U1855 ( .A(n1586), .B(n1132), .Z(out[1077]) );
  XOR U1856 ( .A(in[1545]), .B(in[585]), .Z(n1134) );
  XNOR U1857 ( .A(in[905]), .B(in[265]), .Z(n1133) );
  XNOR U1858 ( .A(n1134), .B(n1133), .Z(n1135) );
  XNOR U1859 ( .A(in[1225]), .B(n1135), .Z(n1517) );
  XNOR U1860 ( .A(n1136), .B(n1517), .Z(n3581) );
  XNOR U1861 ( .A(in[521]), .B(n3581), .Z(n1588) );
  NOR U1862 ( .A(n1359), .B(n1754), .Z(n1137) );
  XNOR U1863 ( .A(n1588), .B(n1137), .Z(out[1078]) );
  XOR U1864 ( .A(in[1546]), .B(in[586]), .Z(n1139) );
  XNOR U1865 ( .A(in[906]), .B(in[266]), .Z(n1138) );
  XNOR U1866 ( .A(n1139), .B(n1138), .Z(n1140) );
  XNOR U1867 ( .A(in[1226]), .B(n1140), .Z(n1521) );
  XNOR U1868 ( .A(n1141), .B(n1521), .Z(n3585) );
  XNOR U1869 ( .A(in[522]), .B(n3585), .Z(n1590) );
  NOR U1870 ( .A(n1363), .B(n1758), .Z(n1142) );
  XNOR U1871 ( .A(n1590), .B(n1142), .Z(out[1079]) );
  XNOR U1872 ( .A(n1144), .B(n1143), .Z(n3624) );
  XNOR U1873 ( .A(in[578]), .B(n3624), .Z(n2565) );
  XOR U1874 ( .A(in[233]), .B(n3721), .Z(n2931) );
  XNOR U1875 ( .A(in[1453]), .B(n3762), .Z(n2928) );
  NAND U1876 ( .A(n2931), .B(n2928), .Z(n1145) );
  XNOR U1877 ( .A(n2565), .B(n1145), .Z(out[107]) );
  XOR U1878 ( .A(in[1547]), .B(in[587]), .Z(n1147) );
  XNOR U1879 ( .A(in[907]), .B(in[267]), .Z(n1146) );
  XNOR U1880 ( .A(n1147), .B(n1146), .Z(n1148) );
  XNOR U1881 ( .A(in[1227]), .B(n1148), .Z(n1525) );
  XNOR U1882 ( .A(n1149), .B(n1525), .Z(n3589) );
  XNOR U1883 ( .A(in[523]), .B(n3589), .Z(n1592) );
  NOR U1884 ( .A(n1367), .B(n1762), .Z(n1150) );
  XNOR U1885 ( .A(n1592), .B(n1150), .Z(out[1080]) );
  XOR U1886 ( .A(in[1548]), .B(in[588]), .Z(n1152) );
  XNOR U1887 ( .A(in[908]), .B(in[268]), .Z(n1151) );
  XNOR U1888 ( .A(n1152), .B(n1151), .Z(n1153) );
  XNOR U1889 ( .A(in[1228]), .B(n1153), .Z(n1529) );
  XNOR U1890 ( .A(n1154), .B(n1529), .Z(n3593) );
  XNOR U1891 ( .A(in[524]), .B(n3593), .Z(n1594) );
  NOR U1892 ( .A(n1371), .B(n1766), .Z(n1155) );
  XNOR U1893 ( .A(n1594), .B(n1155), .Z(out[1081]) );
  XOR U1894 ( .A(in[1549]), .B(in[589]), .Z(n1157) );
  XNOR U1895 ( .A(in[909]), .B(in[269]), .Z(n1156) );
  XNOR U1896 ( .A(n1157), .B(n1156), .Z(n1158) );
  XOR U1897 ( .A(in[1229]), .B(n1158), .Z(n1533) );
  XNOR U1898 ( .A(n1533), .B(n1159), .Z(n3597) );
  XNOR U1899 ( .A(in[525]), .B(n3597), .Z(n1597) );
  NOR U1900 ( .A(n1375), .B(n1770), .Z(n1160) );
  XNOR U1901 ( .A(n1597), .B(n1160), .Z(out[1082]) );
  XOR U1902 ( .A(in[1550]), .B(in[590]), .Z(n1162) );
  XNOR U1903 ( .A(in[910]), .B(in[270]), .Z(n1161) );
  XNOR U1904 ( .A(n1162), .B(n1161), .Z(n1163) );
  XOR U1905 ( .A(in[1230]), .B(n1163), .Z(n1537) );
  XNOR U1906 ( .A(n1537), .B(n1164), .Z(n3601) );
  XNOR U1907 ( .A(in[526]), .B(n3601), .Z(n1599) );
  NOR U1908 ( .A(n1379), .B(n1774), .Z(n1165) );
  XNOR U1909 ( .A(n1599), .B(n1165), .Z(out[1083]) );
  XOR U1910 ( .A(in[1551]), .B(in[591]), .Z(n1167) );
  XNOR U1911 ( .A(in[911]), .B(in[271]), .Z(n1166) );
  XNOR U1912 ( .A(n1167), .B(n1166), .Z(n1168) );
  XOR U1913 ( .A(in[1231]), .B(n1168), .Z(n1541) );
  XNOR U1914 ( .A(n1541), .B(n1169), .Z(n3605) );
  XNOR U1915 ( .A(in[527]), .B(n3605), .Z(n1601) );
  NOR U1916 ( .A(n1383), .B(n1778), .Z(n1170) );
  XNOR U1917 ( .A(n1601), .B(n1170), .Z(out[1084]) );
  XOR U1918 ( .A(in[1552]), .B(in[592]), .Z(n1172) );
  XNOR U1919 ( .A(in[912]), .B(in[272]), .Z(n1171) );
  XNOR U1920 ( .A(n1172), .B(n1171), .Z(n1173) );
  XOR U1921 ( .A(in[1232]), .B(n1173), .Z(n1545) );
  XNOR U1922 ( .A(n1545), .B(n1174), .Z(n3609) );
  XNOR U1923 ( .A(in[528]), .B(n3609), .Z(n1603) );
  NOR U1924 ( .A(n1387), .B(n1782), .Z(n1175) );
  XNOR U1925 ( .A(n1603), .B(n1175), .Z(out[1085]) );
  XOR U1926 ( .A(in[1553]), .B(in[593]), .Z(n1177) );
  XNOR U1927 ( .A(in[913]), .B(in[273]), .Z(n1176) );
  XNOR U1928 ( .A(n1177), .B(n1176), .Z(n1178) );
  XOR U1929 ( .A(in[1233]), .B(n1178), .Z(n1550) );
  XNOR U1930 ( .A(n1550), .B(n1179), .Z(n3613) );
  XNOR U1931 ( .A(in[529]), .B(n3613), .Z(n1605) );
  NOR U1932 ( .A(n1390), .B(n1786), .Z(n1180) );
  XNOR U1933 ( .A(n1605), .B(n1180), .Z(out[1086]) );
  XOR U1934 ( .A(in[1554]), .B(in[594]), .Z(n1182) );
  XNOR U1935 ( .A(in[914]), .B(in[274]), .Z(n1181) );
  XNOR U1936 ( .A(n1182), .B(n1181), .Z(n1183) );
  XOR U1937 ( .A(in[1234]), .B(n1183), .Z(n1554) );
  XNOR U1938 ( .A(n1554), .B(n1184), .Z(n3617) );
  XNOR U1939 ( .A(in[530]), .B(n3617), .Z(n1607) );
  NOR U1940 ( .A(n1392), .B(n1790), .Z(n1185) );
  XNOR U1941 ( .A(n1607), .B(n1185), .Z(out[1087]) );
  XOR U1942 ( .A(in[957]), .B(n3600), .Z(n1609) );
  NOR U1943 ( .A(n1396), .B(n4631), .Z(n1186) );
  XNOR U1944 ( .A(n1609), .B(n1186), .Z(out[1088]) );
  XOR U1945 ( .A(in[958]), .B(n3604), .Z(n1611) );
  NOR U1946 ( .A(n1400), .B(n4635), .Z(n1187) );
  XNOR U1947 ( .A(n1611), .B(n1187), .Z(out[1089]) );
  XOR U1948 ( .A(n1189), .B(n1188), .Z(n3628) );
  XNOR U1949 ( .A(in[579]), .B(n3628), .Z(n2567) );
  XOR U1950 ( .A(in[234]), .B(n3725), .Z(n2947) );
  XNOR U1951 ( .A(in[1454]), .B(n3766), .Z(n2944) );
  NAND U1952 ( .A(n2947), .B(n2944), .Z(n1190) );
  XNOR U1953 ( .A(n2567), .B(n1190), .Z(out[108]) );
  XOR U1954 ( .A(in[959]), .B(n3608), .Z(n1613) );
  NOR U1955 ( .A(n1404), .B(n4639), .Z(n1191) );
  XNOR U1956 ( .A(n1613), .B(n1191), .Z(out[1090]) );
  XOR U1957 ( .A(in[896]), .B(n3612), .Z(n1615) );
  NOR U1958 ( .A(n1408), .B(n4643), .Z(n1192) );
  XNOR U1959 ( .A(n1615), .B(n1192), .Z(out[1091]) );
  XOR U1960 ( .A(in[897]), .B(n3616), .Z(n1618) );
  NOR U1961 ( .A(n1412), .B(n4647), .Z(n1193) );
  XNOR U1962 ( .A(n1618), .B(n1193), .Z(out[1092]) );
  XOR U1963 ( .A(in[898]), .B(n3624), .Z(n1620) );
  NOR U1964 ( .A(n1416), .B(n4651), .Z(n1194) );
  XNOR U1965 ( .A(n1620), .B(n1194), .Z(out[1093]) );
  XOR U1966 ( .A(in[899]), .B(n3628), .Z(n1622) );
  NOR U1967 ( .A(n1420), .B(n4655), .Z(n1195) );
  XNOR U1968 ( .A(n1622), .B(n1195), .Z(out[1094]) );
  XNOR U1969 ( .A(n1197), .B(n1196), .Z(n3632) );
  XNOR U1970 ( .A(in[900]), .B(n3632), .Z(n1624) );
  NOR U1971 ( .A(n1424), .B(n4659), .Z(n1198) );
  XNOR U1972 ( .A(n1624), .B(n1198), .Z(out[1095]) );
  XNOR U1973 ( .A(n1200), .B(n1199), .Z(n3636) );
  XNOR U1974 ( .A(in[901]), .B(n3636), .Z(n1626) );
  NOR U1975 ( .A(n1429), .B(n4663), .Z(n1201) );
  XNOR U1976 ( .A(n1626), .B(n1201), .Z(out[1096]) );
  XNOR U1977 ( .A(n1203), .B(n1202), .Z(n3640) );
  XNOR U1978 ( .A(in[902]), .B(n3640), .Z(n1628) );
  NOR U1979 ( .A(n1433), .B(n4667), .Z(n1204) );
  XNOR U1980 ( .A(n1628), .B(n1204), .Z(out[1097]) );
  XNOR U1981 ( .A(n1206), .B(n1205), .Z(n3644) );
  XNOR U1982 ( .A(in[903]), .B(n3644), .Z(n1630) );
  NOR U1983 ( .A(n1437), .B(n4675), .Z(n1207) );
  XNOR U1984 ( .A(n1630), .B(n1207), .Z(out[1098]) );
  XNOR U1985 ( .A(n1209), .B(n1208), .Z(n3648) );
  XNOR U1986 ( .A(in[904]), .B(n3648), .Z(n1632) );
  NOR U1987 ( .A(n1441), .B(n4679), .Z(n1210) );
  XNOR U1988 ( .A(n1632), .B(n1210), .Z(out[1099]) );
  XOR U1989 ( .A(in[580]), .B(n3632), .Z(n2569) );
  XOR U1990 ( .A(in[235]), .B(n3729), .Z(n2971) );
  XNOR U1991 ( .A(in[1455]), .B(n3770), .Z(n2968) );
  NAND U1992 ( .A(n2971), .B(n2968), .Z(n1211) );
  XNOR U1993 ( .A(n2569), .B(n1211), .Z(out[109]) );
  XOR U1994 ( .A(in[200]), .B(n3573), .Z(n3921) );
  XNOR U1995 ( .A(in[1420]), .B(n3614), .Z(n3920) );
  XOR U1996 ( .A(n4120), .B(in[1043]), .Z(n2632) );
  NAND U1997 ( .A(n3920), .B(n2632), .Z(n1212) );
  XNOR U1998 ( .A(n3921), .B(n1212), .Z(out[10]) );
  XNOR U1999 ( .A(n1214), .B(n1213), .Z(n3652) );
  XNOR U2000 ( .A(in[905]), .B(n3652), .Z(n1634) );
  NOR U2001 ( .A(n1445), .B(n4683), .Z(n1215) );
  XNOR U2002 ( .A(n1634), .B(n1215), .Z(out[1100]) );
  XNOR U2003 ( .A(n1217), .B(n1216), .Z(n3656) );
  XNOR U2004 ( .A(in[906]), .B(n3656), .Z(n1636) );
  NOR U2005 ( .A(n1449), .B(n4687), .Z(n1218) );
  XNOR U2006 ( .A(n1636), .B(n1218), .Z(out[1101]) );
  XNOR U2007 ( .A(n1220), .B(n1219), .Z(n3660) );
  XNOR U2008 ( .A(in[907]), .B(n3660), .Z(n1639) );
  NOR U2009 ( .A(n1453), .B(n4691), .Z(n1221) );
  XNOR U2010 ( .A(n1639), .B(n1221), .Z(out[1102]) );
  XNOR U2011 ( .A(n1223), .B(n1222), .Z(n3668) );
  XNOR U2012 ( .A(in[908]), .B(n3668), .Z(n1641) );
  NOR U2013 ( .A(n1457), .B(n4695), .Z(n1224) );
  XNOR U2014 ( .A(n1641), .B(n1224), .Z(out[1103]) );
  XNOR U2015 ( .A(n1226), .B(n1225), .Z(n3672) );
  XNOR U2016 ( .A(in[909]), .B(n3672), .Z(n1643) );
  NOR U2017 ( .A(n1461), .B(n4699), .Z(n1227) );
  XNOR U2018 ( .A(n1643), .B(n1227), .Z(out[1104]) );
  XNOR U2019 ( .A(n1229), .B(n1228), .Z(n3676) );
  XNOR U2020 ( .A(in[910]), .B(n3676), .Z(n1645) );
  NOR U2021 ( .A(n1465), .B(n4703), .Z(n1230) );
  XNOR U2022 ( .A(n1645), .B(n1230), .Z(out[1105]) );
  XNOR U2023 ( .A(n1232), .B(n1231), .Z(n3680) );
  XNOR U2024 ( .A(in[911]), .B(n3680), .Z(n1647) );
  NOR U2025 ( .A(n1470), .B(n4707), .Z(n1233) );
  XNOR U2026 ( .A(n1647), .B(n1233), .Z(out[1106]) );
  XNOR U2027 ( .A(n1235), .B(n1234), .Z(n3684) );
  XNOR U2028 ( .A(in[912]), .B(n3684), .Z(n1649) );
  NOR U2029 ( .A(n1474), .B(n4711), .Z(n1236) );
  XNOR U2030 ( .A(n1649), .B(n1236), .Z(out[1107]) );
  XOR U2031 ( .A(n1238), .B(n1237), .Z(n3688) );
  XNOR U2032 ( .A(in[913]), .B(n3688), .Z(n1651) );
  NOR U2033 ( .A(n1478), .B(n4719), .Z(n1239) );
  XNOR U2034 ( .A(n1651), .B(n1239), .Z(out[1108]) );
  XOR U2035 ( .A(n1241), .B(n1240), .Z(n3692) );
  XNOR U2036 ( .A(in[914]), .B(n3692), .Z(n1653) );
  NOR U2037 ( .A(n1482), .B(n4723), .Z(n1242) );
  XNOR U2038 ( .A(n1653), .B(n1242), .Z(out[1109]) );
  XOR U2039 ( .A(in[581]), .B(n3636), .Z(n2571) );
  XOR U2040 ( .A(in[236]), .B(n3733), .Z(n2995) );
  XNOR U2041 ( .A(in[1456]), .B(n3774), .Z(n2992) );
  NAND U2042 ( .A(n2995), .B(n2992), .Z(n1243) );
  XNOR U2043 ( .A(n2571), .B(n1243), .Z(out[110]) );
  XNOR U2044 ( .A(n1245), .B(n1244), .Z(n3696) );
  XNOR U2045 ( .A(in[915]), .B(n3696), .Z(n1655) );
  NOR U2046 ( .A(n1486), .B(n4727), .Z(n1246) );
  XNOR U2047 ( .A(n1655), .B(n1246), .Z(out[1110]) );
  XOR U2048 ( .A(n1248), .B(n1247), .Z(n3700) );
  XNOR U2049 ( .A(in[916]), .B(n3700), .Z(n1657) );
  NOR U2050 ( .A(n1490), .B(n4731), .Z(n1249) );
  XNOR U2051 ( .A(n1657), .B(n1249), .Z(out[1111]) );
  XNOR U2052 ( .A(n1251), .B(n1250), .Z(n3704) );
  XNOR U2053 ( .A(in[917]), .B(n3704), .Z(n1660) );
  NOR U2054 ( .A(n1494), .B(n4735), .Z(n1252) );
  XNOR U2055 ( .A(n1660), .B(n1252), .Z(out[1112]) );
  XOR U2056 ( .A(n1254), .B(n1253), .Z(n3712) );
  XNOR U2057 ( .A(in[918]), .B(n3712), .Z(n1662) );
  NOR U2058 ( .A(n1498), .B(n4739), .Z(n1255) );
  XNOR U2059 ( .A(n1662), .B(n1255), .Z(out[1113]) );
  XNOR U2060 ( .A(n1257), .B(n1256), .Z(n3716) );
  XNOR U2061 ( .A(in[919]), .B(n3716), .Z(n1664) );
  NOR U2062 ( .A(n1502), .B(n4743), .Z(n1258) );
  XNOR U2063 ( .A(n1664), .B(n1258), .Z(out[1114]) );
  XNOR U2064 ( .A(n1260), .B(n1259), .Z(n3720) );
  XNOR U2065 ( .A(in[920]), .B(n3720), .Z(n1666) );
  NOR U2066 ( .A(n1506), .B(n4747), .Z(n1261) );
  XNOR U2067 ( .A(n1666), .B(n1261), .Z(out[1115]) );
  XNOR U2068 ( .A(n1263), .B(n1262), .Z(n3724) );
  XNOR U2069 ( .A(in[921]), .B(n3724), .Z(n1668) );
  NOR U2070 ( .A(n1511), .B(n4751), .Z(n1264) );
  XNOR U2071 ( .A(n1668), .B(n1264), .Z(out[1116]) );
  XOR U2072 ( .A(n1266), .B(n1265), .Z(n3728) );
  XNOR U2073 ( .A(in[922]), .B(n3728), .Z(n1670) );
  NOR U2074 ( .A(n1515), .B(n4755), .Z(n1267) );
  XNOR U2075 ( .A(n1670), .B(n1267), .Z(out[1117]) );
  XOR U2076 ( .A(n1269), .B(n1268), .Z(n3732) );
  XNOR U2077 ( .A(in[923]), .B(n3732), .Z(n1672) );
  NOR U2078 ( .A(n1519), .B(n4763), .Z(n1270) );
  XNOR U2079 ( .A(n1672), .B(n1270), .Z(out[1118]) );
  XOR U2080 ( .A(n1272), .B(n1271), .Z(n3736) );
  XNOR U2081 ( .A(in[924]), .B(n3736), .Z(n1674) );
  NOR U2082 ( .A(n1523), .B(n4767), .Z(n1273) );
  XNOR U2083 ( .A(n1674), .B(n1273), .Z(out[1119]) );
  XOR U2084 ( .A(in[582]), .B(n3640), .Z(n2573) );
  XOR U2085 ( .A(in[237]), .B(n3737), .Z(n3019) );
  XNOR U2086 ( .A(in[1457]), .B(n3778), .Z(n3016) );
  NAND U2087 ( .A(n3019), .B(n3016), .Z(n1274) );
  XNOR U2088 ( .A(n2573), .B(n1274), .Z(out[111]) );
  XOR U2089 ( .A(n1276), .B(n1275), .Z(n3740) );
  XNOR U2090 ( .A(in[925]), .B(n3740), .Z(n1676) );
  NOR U2091 ( .A(n1527), .B(n4771), .Z(n1277) );
  XNOR U2092 ( .A(n1676), .B(n1277), .Z(out[1120]) );
  XOR U2093 ( .A(n1279), .B(n1278), .Z(n3744) );
  XNOR U2094 ( .A(in[926]), .B(n3744), .Z(n1678) );
  NOR U2095 ( .A(n1531), .B(n4775), .Z(n1280) );
  XNOR U2096 ( .A(n1678), .B(n1280), .Z(out[1121]) );
  XOR U2097 ( .A(n1282), .B(n1281), .Z(n3748) );
  XNOR U2098 ( .A(in[927]), .B(n3748), .Z(n1681) );
  NOR U2099 ( .A(n1535), .B(n4779), .Z(n1283) );
  XNOR U2100 ( .A(n1681), .B(n1283), .Z(out[1122]) );
  XOR U2101 ( .A(n1285), .B(n1284), .Z(n3756) );
  XNOR U2102 ( .A(in[928]), .B(n3756), .Z(n1683) );
  NOR U2103 ( .A(n1539), .B(n4783), .Z(n1286) );
  XNOR U2104 ( .A(n1683), .B(n1286), .Z(out[1123]) );
  XNOR U2105 ( .A(n1288), .B(n1287), .Z(n3760) );
  XNOR U2106 ( .A(in[929]), .B(n3760), .Z(n1685) );
  NOR U2107 ( .A(n1543), .B(n4787), .Z(n1289) );
  XNOR U2108 ( .A(n1685), .B(n1289), .Z(out[1124]) );
  XOR U2109 ( .A(n1291), .B(n1290), .Z(n3764) );
  XNOR U2110 ( .A(in[930]), .B(n3764), .Z(n1687) );
  NOR U2111 ( .A(n1547), .B(n4791), .Z(n1292) );
  XNOR U2112 ( .A(n1687), .B(n1292), .Z(out[1125]) );
  XNOR U2113 ( .A(n1294), .B(n1293), .Z(n3768) );
  XNOR U2114 ( .A(in[931]), .B(n3768), .Z(n1689) );
  NOR U2115 ( .A(n1552), .B(n4795), .Z(n1295) );
  XNOR U2116 ( .A(n1689), .B(n1295), .Z(out[1126]) );
  XNOR U2117 ( .A(n1297), .B(n1296), .Z(n3772) );
  XNOR U2118 ( .A(in[932]), .B(n3772), .Z(n1691) );
  NOR U2119 ( .A(n1556), .B(n4799), .Z(n1298) );
  XNOR U2120 ( .A(n1691), .B(n1298), .Z(out[1127]) );
  XNOR U2121 ( .A(n1300), .B(n1299), .Z(n3776) );
  XNOR U2122 ( .A(in[933]), .B(n3776), .Z(n1694) );
  NAND U2123 ( .A(n1558), .B(n1301), .Z(n1302) );
  XNOR U2124 ( .A(n1694), .B(n1302), .Z(out[1128]) );
  XOR U2125 ( .A(n1304), .B(n1303), .Z(n3780) );
  XNOR U2126 ( .A(in[934]), .B(n3780), .Z(n1698) );
  NAND U2127 ( .A(n1560), .B(n1305), .Z(n1306) );
  XNOR U2128 ( .A(n1698), .B(n1306), .Z(out[1129]) );
  XOR U2129 ( .A(in[583]), .B(n3644), .Z(n2576) );
  XOR U2130 ( .A(in[238]), .B(n3741), .Z(n3043) );
  XNOR U2131 ( .A(in[1458]), .B(n3782), .Z(n3040) );
  NAND U2132 ( .A(n3043), .B(n3040), .Z(n1307) );
  XNOR U2133 ( .A(n2576), .B(n1307), .Z(out[112]) );
  XNOR U2134 ( .A(n1309), .B(n1308), .Z(n3784) );
  XNOR U2135 ( .A(in[935]), .B(n3784), .Z(n1702) );
  NAND U2136 ( .A(n1562), .B(n1310), .Z(n1311) );
  XNOR U2137 ( .A(n1702), .B(n1311), .Z(out[1130]) );
  XNOR U2138 ( .A(n1313), .B(n1312), .Z(n3788) );
  XNOR U2139 ( .A(in[936]), .B(n3788), .Z(n1706) );
  NAND U2140 ( .A(n1564), .B(n1314), .Z(n1315) );
  XNOR U2141 ( .A(n1706), .B(n1315), .Z(out[1131]) );
  XNOR U2142 ( .A(n1317), .B(n1316), .Z(n3792) );
  XNOR U2143 ( .A(in[937]), .B(n3792), .Z(n1711) );
  NAND U2144 ( .A(n1566), .B(n1318), .Z(n1319) );
  XNOR U2145 ( .A(n1711), .B(n1319), .Z(out[1132]) );
  XNOR U2146 ( .A(n1321), .B(n1320), .Z(n3802) );
  XNOR U2147 ( .A(in[938]), .B(n3802), .Z(n1715) );
  NAND U2148 ( .A(n1568), .B(n1322), .Z(n1323) );
  XNOR U2149 ( .A(n1715), .B(n1323), .Z(out[1133]) );
  XNOR U2150 ( .A(n1325), .B(n1324), .Z(n3806) );
  XNOR U2151 ( .A(in[939]), .B(n3806), .Z(n1719) );
  NAND U2152 ( .A(n1570), .B(n1326), .Z(n1327) );
  XNOR U2153 ( .A(n1719), .B(n1327), .Z(out[1134]) );
  XNOR U2154 ( .A(n1329), .B(n1328), .Z(n3810) );
  XNOR U2155 ( .A(in[940]), .B(n3810), .Z(n1723) );
  NAND U2156 ( .A(n1572), .B(n1330), .Z(n1331) );
  XNOR U2157 ( .A(n1723), .B(n1331), .Z(out[1135]) );
  XNOR U2158 ( .A(n1333), .B(n1332), .Z(n3814) );
  XNOR U2159 ( .A(in[941]), .B(n3814), .Z(n1727) );
  NAND U2160 ( .A(n1576), .B(n1334), .Z(n1335) );
  XNOR U2161 ( .A(n1727), .B(n1335), .Z(out[1136]) );
  XNOR U2162 ( .A(n1337), .B(n1336), .Z(n3536) );
  XNOR U2163 ( .A(in[942]), .B(n3536), .Z(n1731) );
  NAND U2164 ( .A(n1578), .B(n1338), .Z(n1339) );
  XNOR U2165 ( .A(n1731), .B(n1339), .Z(out[1137]) );
  XNOR U2166 ( .A(n1341), .B(n1340), .Z(n3540) );
  XNOR U2167 ( .A(in[943]), .B(n3540), .Z(n1735) );
  NAND U2168 ( .A(n1580), .B(n1342), .Z(n1343) );
  XNOR U2169 ( .A(n1735), .B(n1343), .Z(out[1138]) );
  XNOR U2170 ( .A(n1345), .B(n1344), .Z(n3544) );
  XNOR U2171 ( .A(in[944]), .B(n3544), .Z(n1739) );
  NAND U2172 ( .A(n1582), .B(n1346), .Z(n1347) );
  XNOR U2173 ( .A(n1739), .B(n1347), .Z(out[1139]) );
  XOR U2174 ( .A(in[584]), .B(n3648), .Z(n2578) );
  XOR U2175 ( .A(in[239]), .B(n3745), .Z(n3067) );
  XNOR U2176 ( .A(in[1459]), .B(n3786), .Z(n3064) );
  NAND U2177 ( .A(n3067), .B(n3064), .Z(n1348) );
  XNOR U2178 ( .A(n2578), .B(n1348), .Z(out[113]) );
  XNOR U2179 ( .A(n1350), .B(n1349), .Z(n3548) );
  XNOR U2180 ( .A(in[945]), .B(n3548), .Z(n1743) );
  NAND U2181 ( .A(n1584), .B(n1351), .Z(n1352) );
  XNOR U2182 ( .A(n1743), .B(n1352), .Z(out[1140]) );
  XNOR U2183 ( .A(n1354), .B(n1353), .Z(n3552) );
  XNOR U2184 ( .A(in[946]), .B(n3552), .Z(n1747) );
  NAND U2185 ( .A(n1586), .B(n1355), .Z(n1356) );
  XNOR U2186 ( .A(n1747), .B(n1356), .Z(out[1141]) );
  XNOR U2187 ( .A(n1358), .B(n1357), .Z(n3556) );
  XNOR U2188 ( .A(in[947]), .B(n3556), .Z(n1752) );
  NAND U2189 ( .A(n1588), .B(n1359), .Z(n1360) );
  XNOR U2190 ( .A(n1752), .B(n1360), .Z(out[1142]) );
  XNOR U2191 ( .A(n1362), .B(n1361), .Z(n3560) );
  XNOR U2192 ( .A(in[948]), .B(n3560), .Z(n1756) );
  NAND U2193 ( .A(n1590), .B(n1363), .Z(n1364) );
  XNOR U2194 ( .A(n1756), .B(n1364), .Z(out[1143]) );
  XNOR U2195 ( .A(n1366), .B(n1365), .Z(n3564) );
  XNOR U2196 ( .A(in[949]), .B(n3564), .Z(n1760) );
  NAND U2197 ( .A(n1592), .B(n1367), .Z(n1368) );
  XNOR U2198 ( .A(n1760), .B(n1368), .Z(out[1144]) );
  XNOR U2199 ( .A(n1370), .B(n1369), .Z(n3568) );
  XNOR U2200 ( .A(in[950]), .B(n3568), .Z(n1764) );
  NAND U2201 ( .A(n1594), .B(n1371), .Z(n1372) );
  XNOR U2202 ( .A(n1764), .B(n1372), .Z(out[1145]) );
  XNOR U2203 ( .A(n1374), .B(n1373), .Z(n3572) );
  XNOR U2204 ( .A(in[951]), .B(n3572), .Z(n1768) );
  NAND U2205 ( .A(n1597), .B(n1375), .Z(n1376) );
  XNOR U2206 ( .A(n1768), .B(n1376), .Z(out[1146]) );
  XNOR U2207 ( .A(n1378), .B(n1377), .Z(n3580) );
  XNOR U2208 ( .A(in[952]), .B(n3580), .Z(n1772) );
  NAND U2209 ( .A(n1599), .B(n1379), .Z(n1380) );
  XNOR U2210 ( .A(n1772), .B(n1380), .Z(out[1147]) );
  XNOR U2211 ( .A(n1382), .B(n1381), .Z(n3584) );
  XNOR U2212 ( .A(in[953]), .B(n3584), .Z(n1776) );
  NAND U2213 ( .A(n1601), .B(n1383), .Z(n1384) );
  XNOR U2214 ( .A(n1776), .B(n1384), .Z(out[1148]) );
  XNOR U2215 ( .A(n1386), .B(n1385), .Z(n3588) );
  XNOR U2216 ( .A(in[954]), .B(n3588), .Z(n1780) );
  NAND U2217 ( .A(n1603), .B(n1387), .Z(n1388) );
  XNOR U2218 ( .A(n1780), .B(n1388), .Z(out[1149]) );
  XOR U2219 ( .A(in[585]), .B(n3652), .Z(n2580) );
  XOR U2220 ( .A(in[240]), .B(n3749), .Z(n3093) );
  XNOR U2221 ( .A(in[1460]), .B(n3790), .Z(n3090) );
  NAND U2222 ( .A(n3093), .B(n3090), .Z(n1389) );
  XNOR U2223 ( .A(n2580), .B(n1389), .Z(out[114]) );
  XNOR U2224 ( .A(in[955]), .B(n3592), .Z(n1784) );
  NAND U2225 ( .A(n1605), .B(n1390), .Z(n1391) );
  XNOR U2226 ( .A(n1784), .B(n1391), .Z(out[1150]) );
  XNOR U2227 ( .A(in[956]), .B(n3596), .Z(n1788) );
  NAND U2228 ( .A(n1607), .B(n1392), .Z(n1393) );
  XNOR U2229 ( .A(n1788), .B(n1393), .Z(out[1151]) );
  XNOR U2230 ( .A(n1395), .B(n1394), .Z(n3936) );
  XNOR U2231 ( .A(in[1004]), .B(n3936), .Z(n4629) );
  NAND U2232 ( .A(n1609), .B(n1396), .Z(n1397) );
  XNOR U2233 ( .A(n4629), .B(n1397), .Z(out[1152]) );
  XNOR U2234 ( .A(n1399), .B(n1398), .Z(n3938) );
  XNOR U2235 ( .A(in[1005]), .B(n3938), .Z(n4633) );
  NAND U2236 ( .A(n1611), .B(n1400), .Z(n1401) );
  XNOR U2237 ( .A(n4633), .B(n1401), .Z(out[1153]) );
  XNOR U2238 ( .A(n1403), .B(n1402), .Z(n3940) );
  XNOR U2239 ( .A(in[1006]), .B(n3940), .Z(n4637) );
  NAND U2240 ( .A(n1613), .B(n1404), .Z(n1405) );
  XNOR U2241 ( .A(n4637), .B(n1405), .Z(out[1154]) );
  XNOR U2242 ( .A(n1407), .B(n1406), .Z(n3942) );
  XNOR U2243 ( .A(in[1007]), .B(n3942), .Z(n4641) );
  NAND U2244 ( .A(n1615), .B(n1408), .Z(n1409) );
  XNOR U2245 ( .A(n4641), .B(n1409), .Z(out[1155]) );
  XNOR U2246 ( .A(n1411), .B(n1410), .Z(n3948) );
  XNOR U2247 ( .A(in[1008]), .B(n3948), .Z(n4645) );
  NAND U2248 ( .A(n1618), .B(n1412), .Z(n1413) );
  XNOR U2249 ( .A(n4645), .B(n1413), .Z(out[1156]) );
  XNOR U2250 ( .A(n1415), .B(n1414), .Z(n3950) );
  XNOR U2251 ( .A(in[1009]), .B(n3950), .Z(n4649) );
  NAND U2252 ( .A(n1620), .B(n1416), .Z(n1417) );
  XNOR U2253 ( .A(n4649), .B(n1417), .Z(out[1157]) );
  XNOR U2254 ( .A(n1419), .B(n1418), .Z(n3952) );
  XNOR U2255 ( .A(in[1010]), .B(n3952), .Z(n4653) );
  NAND U2256 ( .A(n1622), .B(n1420), .Z(n1421) );
  XNOR U2257 ( .A(n4653), .B(n1421), .Z(out[1158]) );
  XNOR U2258 ( .A(n1423), .B(n1422), .Z(n3954) );
  XNOR U2259 ( .A(in[1011]), .B(n3954), .Z(n4657) );
  NAND U2260 ( .A(n1624), .B(n1424), .Z(n1425) );
  XNOR U2261 ( .A(n4657), .B(n1425), .Z(out[1159]) );
  XOR U2262 ( .A(in[586]), .B(n3656), .Z(n2582) );
  XOR U2263 ( .A(in[241]), .B(n3757), .Z(n3117) );
  XNOR U2264 ( .A(in[1461]), .B(n3794), .Z(n3114) );
  NAND U2265 ( .A(n3117), .B(n3114), .Z(n1426) );
  XNOR U2266 ( .A(n2582), .B(n1426), .Z(out[115]) );
  XNOR U2267 ( .A(n1428), .B(n1427), .Z(n3956) );
  XNOR U2268 ( .A(in[1012]), .B(n3956), .Z(n4661) );
  NAND U2269 ( .A(n1626), .B(n1429), .Z(n1430) );
  XNOR U2270 ( .A(n4661), .B(n1430), .Z(out[1160]) );
  XNOR U2271 ( .A(n1432), .B(n1431), .Z(n3958) );
  XNOR U2272 ( .A(in[1013]), .B(n3958), .Z(n4665) );
  NAND U2273 ( .A(n1628), .B(n1433), .Z(n1434) );
  XNOR U2274 ( .A(n4665), .B(n1434), .Z(out[1161]) );
  XNOR U2275 ( .A(n1436), .B(n1435), .Z(n3960) );
  XNOR U2276 ( .A(in[1014]), .B(n3960), .Z(n4673) );
  NAND U2277 ( .A(n1630), .B(n1437), .Z(n1438) );
  XNOR U2278 ( .A(n4673), .B(n1438), .Z(out[1162]) );
  XNOR U2279 ( .A(n1440), .B(n1439), .Z(n3962) );
  XNOR U2280 ( .A(in[1015]), .B(n3962), .Z(n4677) );
  NAND U2281 ( .A(n1632), .B(n1441), .Z(n1442) );
  XNOR U2282 ( .A(n4677), .B(n1442), .Z(out[1163]) );
  XNOR U2283 ( .A(n1444), .B(n1443), .Z(n3818) );
  XNOR U2284 ( .A(in[1016]), .B(n3818), .Z(n4681) );
  NAND U2285 ( .A(n1634), .B(n1445), .Z(n1446) );
  XNOR U2286 ( .A(n4681), .B(n1446), .Z(out[1164]) );
  XNOR U2287 ( .A(n1448), .B(n1447), .Z(n3820) );
  XNOR U2288 ( .A(in[1017]), .B(n3820), .Z(n4685) );
  NAND U2289 ( .A(n1636), .B(n1449), .Z(n1450) );
  XNOR U2290 ( .A(n4685), .B(n1450), .Z(out[1165]) );
  XNOR U2291 ( .A(n1452), .B(n1451), .Z(n3822) );
  XNOR U2292 ( .A(in[1018]), .B(n3822), .Z(n4689) );
  NAND U2293 ( .A(n1639), .B(n1453), .Z(n1454) );
  XNOR U2294 ( .A(n4689), .B(n1454), .Z(out[1166]) );
  XNOR U2295 ( .A(n1456), .B(n1455), .Z(n3824) );
  XNOR U2296 ( .A(in[1019]), .B(n3824), .Z(n4693) );
  NAND U2297 ( .A(n1641), .B(n1457), .Z(n1458) );
  XNOR U2298 ( .A(n4693), .B(n1458), .Z(out[1167]) );
  XOR U2299 ( .A(n1460), .B(n1459), .Z(n3826) );
  XNOR U2300 ( .A(in[1020]), .B(n3826), .Z(n4697) );
  NAND U2301 ( .A(n1643), .B(n1461), .Z(n1462) );
  XNOR U2302 ( .A(n4697), .B(n1462), .Z(out[1168]) );
  XOR U2303 ( .A(n1464), .B(n1463), .Z(n3828) );
  XNOR U2304 ( .A(in[1021]), .B(n3828), .Z(n4701) );
  NAND U2305 ( .A(n1645), .B(n1465), .Z(n1466) );
  XNOR U2306 ( .A(n4701), .B(n1466), .Z(out[1169]) );
  XOR U2307 ( .A(in[587]), .B(n3660), .Z(n2584) );
  XOR U2308 ( .A(in[242]), .B(n3761), .Z(n3141) );
  XNOR U2309 ( .A(in[1462]), .B(n3804), .Z(n3138) );
  NAND U2310 ( .A(n3141), .B(n3138), .Z(n1467) );
  XNOR U2311 ( .A(n2584), .B(n1467), .Z(out[116]) );
  XOR U2312 ( .A(n1469), .B(n1468), .Z(n3834) );
  XNOR U2313 ( .A(in[1022]), .B(n3834), .Z(n4705) );
  NAND U2314 ( .A(n1647), .B(n1470), .Z(n1471) );
  XNOR U2315 ( .A(n4705), .B(n1471), .Z(out[1170]) );
  XNOR U2316 ( .A(n1473), .B(n1472), .Z(n3836) );
  XNOR U2317 ( .A(in[1023]), .B(n3836), .Z(n4709) );
  NAND U2318 ( .A(n1649), .B(n1474), .Z(n1475) );
  XNOR U2319 ( .A(n4709), .B(n1475), .Z(out[1171]) );
  XOR U2320 ( .A(n1477), .B(n1476), .Z(n3838) );
  XNOR U2321 ( .A(in[960]), .B(n3838), .Z(n4717) );
  NAND U2322 ( .A(n1651), .B(n1478), .Z(n1479) );
  XNOR U2323 ( .A(n4717), .B(n1479), .Z(out[1172]) );
  XOR U2324 ( .A(n1481), .B(n1480), .Z(n3840) );
  XNOR U2325 ( .A(in[961]), .B(n3840), .Z(n4721) );
  NAND U2326 ( .A(n1653), .B(n1482), .Z(n1483) );
  XNOR U2327 ( .A(n4721), .B(n1483), .Z(out[1173]) );
  XOR U2328 ( .A(n1485), .B(n1484), .Z(n3842) );
  XNOR U2329 ( .A(in[962]), .B(n3842), .Z(n4725) );
  NAND U2330 ( .A(n1655), .B(n1486), .Z(n1487) );
  XNOR U2331 ( .A(n4725), .B(n1487), .Z(out[1174]) );
  XOR U2332 ( .A(n1489), .B(n1488), .Z(n3844) );
  XNOR U2333 ( .A(in[963]), .B(n3844), .Z(n4729) );
  NAND U2334 ( .A(n1657), .B(n1490), .Z(n1491) );
  XNOR U2335 ( .A(n4729), .B(n1491), .Z(out[1175]) );
  XOR U2336 ( .A(n1493), .B(n1492), .Z(n3846) );
  XNOR U2337 ( .A(in[964]), .B(n3846), .Z(n4733) );
  NAND U2338 ( .A(n1660), .B(n1494), .Z(n1495) );
  XNOR U2339 ( .A(n4733), .B(n1495), .Z(out[1176]) );
  XOR U2340 ( .A(n1497), .B(n1496), .Z(n3848) );
  XNOR U2341 ( .A(in[965]), .B(n3848), .Z(n4737) );
  NAND U2342 ( .A(n1662), .B(n1498), .Z(n1499) );
  XNOR U2343 ( .A(n4737), .B(n1499), .Z(out[1177]) );
  XOR U2344 ( .A(n1501), .B(n1500), .Z(n3850) );
  XNOR U2345 ( .A(in[966]), .B(n3850), .Z(n4741) );
  NAND U2346 ( .A(n1664), .B(n1502), .Z(n1503) );
  XNOR U2347 ( .A(n4741), .B(n1503), .Z(out[1178]) );
  XOR U2348 ( .A(n1505), .B(n1504), .Z(n3852) );
  XNOR U2349 ( .A(in[967]), .B(n3852), .Z(n4745) );
  NAND U2350 ( .A(n1666), .B(n1506), .Z(n1507) );
  XNOR U2351 ( .A(n4745), .B(n1507), .Z(out[1179]) );
  XOR U2352 ( .A(in[588]), .B(n3668), .Z(n2586) );
  XOR U2353 ( .A(in[243]), .B(n3765), .Z(n3165) );
  XNOR U2354 ( .A(in[1463]), .B(n3808), .Z(n3162) );
  NAND U2355 ( .A(n3165), .B(n3162), .Z(n1508) );
  XNOR U2356 ( .A(n2586), .B(n1508), .Z(out[117]) );
  XOR U2357 ( .A(n1510), .B(n1509), .Z(n3856) );
  XNOR U2358 ( .A(in[968]), .B(n3856), .Z(n4749) );
  NAND U2359 ( .A(n1668), .B(n1511), .Z(n1512) );
  XNOR U2360 ( .A(n4749), .B(n1512), .Z(out[1180]) );
  XOR U2361 ( .A(n1514), .B(n1513), .Z(n3858) );
  XNOR U2362 ( .A(in[969]), .B(n3858), .Z(n4753) );
  NAND U2363 ( .A(n1670), .B(n1515), .Z(n1516) );
  XNOR U2364 ( .A(n4753), .B(n1516), .Z(out[1181]) );
  XOR U2365 ( .A(n1518), .B(n1517), .Z(n3860) );
  XNOR U2366 ( .A(in[970]), .B(n3860), .Z(n4761) );
  NAND U2367 ( .A(n1672), .B(n1519), .Z(n1520) );
  XNOR U2368 ( .A(n4761), .B(n1520), .Z(out[1182]) );
  XOR U2369 ( .A(n1522), .B(n1521), .Z(n3862) );
  XNOR U2370 ( .A(in[971]), .B(n3862), .Z(n4765) );
  NAND U2371 ( .A(n1674), .B(n1523), .Z(n1524) );
  XNOR U2372 ( .A(n4765), .B(n1524), .Z(out[1183]) );
  XOR U2373 ( .A(n1526), .B(n1525), .Z(n3864) );
  XNOR U2374 ( .A(in[972]), .B(n3864), .Z(n4769) );
  NAND U2375 ( .A(n1676), .B(n1527), .Z(n1528) );
  XNOR U2376 ( .A(n4769), .B(n1528), .Z(out[1184]) );
  XOR U2377 ( .A(n1530), .B(n1529), .Z(n3866) );
  XNOR U2378 ( .A(in[973]), .B(n3866), .Z(n4773) );
  NAND U2379 ( .A(n1678), .B(n1531), .Z(n1532) );
  XNOR U2380 ( .A(n4773), .B(n1532), .Z(out[1185]) );
  XNOR U2381 ( .A(n1534), .B(n1533), .Z(n3868) );
  XNOR U2382 ( .A(in[974]), .B(n3868), .Z(n4777) );
  NAND U2383 ( .A(n1681), .B(n1535), .Z(n1536) );
  XNOR U2384 ( .A(n4777), .B(n1536), .Z(out[1186]) );
  XNOR U2385 ( .A(n1538), .B(n1537), .Z(n3870) );
  XNOR U2386 ( .A(in[975]), .B(n3870), .Z(n4781) );
  NAND U2387 ( .A(n1683), .B(n1539), .Z(n1540) );
  XNOR U2388 ( .A(n4781), .B(n1540), .Z(out[1187]) );
  XNOR U2389 ( .A(n1542), .B(n1541), .Z(n3872) );
  XNOR U2390 ( .A(in[976]), .B(n3872), .Z(n4785) );
  NAND U2391 ( .A(n1685), .B(n1543), .Z(n1544) );
  XNOR U2392 ( .A(n4785), .B(n1544), .Z(out[1188]) );
  XNOR U2393 ( .A(n1546), .B(n1545), .Z(n3874) );
  XNOR U2394 ( .A(in[977]), .B(n3874), .Z(n4789) );
  NAND U2395 ( .A(n1687), .B(n1547), .Z(n1548) );
  XNOR U2396 ( .A(n4789), .B(n1548), .Z(out[1189]) );
  XOR U2397 ( .A(in[589]), .B(n3672), .Z(n2588) );
  XOR U2398 ( .A(in[244]), .B(n3769), .Z(n3189) );
  XNOR U2399 ( .A(in[1464]), .B(n3812), .Z(n3186) );
  NAND U2400 ( .A(n3189), .B(n3186), .Z(n1549) );
  XNOR U2401 ( .A(n2588), .B(n1549), .Z(out[118]) );
  XNOR U2402 ( .A(n1551), .B(n1550), .Z(n3878) );
  XNOR U2403 ( .A(in[978]), .B(n3878), .Z(n4793) );
  NAND U2404 ( .A(n1689), .B(n1552), .Z(n1553) );
  XNOR U2405 ( .A(n4793), .B(n1553), .Z(out[1190]) );
  XNOR U2406 ( .A(n1555), .B(n1554), .Z(n3880) );
  XNOR U2407 ( .A(in[979]), .B(n3880), .Z(n4797) );
  NAND U2408 ( .A(n1691), .B(n1556), .Z(n1557) );
  XNOR U2409 ( .A(n4797), .B(n1557), .Z(out[1191]) );
  OR U2410 ( .A(n1694), .B(n1558), .Z(n1559) );
  XNOR U2411 ( .A(n1693), .B(n1559), .Z(out[1192]) );
  OR U2412 ( .A(n1698), .B(n1560), .Z(n1561) );
  XNOR U2413 ( .A(n1697), .B(n1561), .Z(out[1193]) );
  OR U2414 ( .A(n1702), .B(n1562), .Z(n1563) );
  XNOR U2415 ( .A(n1701), .B(n1563), .Z(out[1194]) );
  OR U2416 ( .A(n1706), .B(n1564), .Z(n1565) );
  XNOR U2417 ( .A(n1705), .B(n1565), .Z(out[1195]) );
  OR U2418 ( .A(n1711), .B(n1566), .Z(n1567) );
  XNOR U2419 ( .A(n1710), .B(n1567), .Z(out[1196]) );
  OR U2420 ( .A(n1715), .B(n1568), .Z(n1569) );
  XNOR U2421 ( .A(n1714), .B(n1569), .Z(out[1197]) );
  OR U2422 ( .A(n1719), .B(n1570), .Z(n1571) );
  XNOR U2423 ( .A(n1718), .B(n1571), .Z(out[1198]) );
  OR U2424 ( .A(n1723), .B(n1572), .Z(n1573) );
  XNOR U2425 ( .A(n1722), .B(n1573), .Z(out[1199]) );
  XOR U2426 ( .A(in[590]), .B(n3676), .Z(n2590) );
  XOR U2427 ( .A(in[245]), .B(n3773), .Z(n3213) );
  XNOR U2428 ( .A(in[1465]), .B(n3816), .Z(n3210) );
  NAND U2429 ( .A(n3213), .B(n3210), .Z(n1574) );
  XNOR U2430 ( .A(n2590), .B(n1574), .Z(out[119]) );
  XOR U2431 ( .A(in[201]), .B(n3581), .Z(n3945) );
  XNOR U2432 ( .A(in[1421]), .B(n3618), .Z(n3944) );
  XOR U2433 ( .A(in[1044]), .B(n4123), .Z(n2635) );
  NAND U2434 ( .A(n3944), .B(n2635), .Z(n1575) );
  XNOR U2435 ( .A(n3945), .B(n1575), .Z(out[11]) );
  OR U2436 ( .A(n1727), .B(n1576), .Z(n1577) );
  XNOR U2437 ( .A(n1726), .B(n1577), .Z(out[1200]) );
  OR U2438 ( .A(n1731), .B(n1578), .Z(n1579) );
  XNOR U2439 ( .A(n1730), .B(n1579), .Z(out[1201]) );
  OR U2440 ( .A(n1735), .B(n1580), .Z(n1581) );
  XNOR U2441 ( .A(n1734), .B(n1581), .Z(out[1202]) );
  OR U2442 ( .A(n1739), .B(n1582), .Z(n1583) );
  XNOR U2443 ( .A(n1738), .B(n1583), .Z(out[1203]) );
  OR U2444 ( .A(n1743), .B(n1584), .Z(n1585) );
  XNOR U2445 ( .A(n1742), .B(n1585), .Z(out[1204]) );
  OR U2446 ( .A(n1747), .B(n1586), .Z(n1587) );
  XNOR U2447 ( .A(n1746), .B(n1587), .Z(out[1205]) );
  OR U2448 ( .A(n1752), .B(n1588), .Z(n1589) );
  XNOR U2449 ( .A(n1751), .B(n1589), .Z(out[1206]) );
  OR U2450 ( .A(n1756), .B(n1590), .Z(n1591) );
  XNOR U2451 ( .A(n1755), .B(n1591), .Z(out[1207]) );
  OR U2452 ( .A(n1760), .B(n1592), .Z(n1593) );
  XNOR U2453 ( .A(n1759), .B(n1593), .Z(out[1208]) );
  OR U2454 ( .A(n1764), .B(n1594), .Z(n1595) );
  XNOR U2455 ( .A(n1763), .B(n1595), .Z(out[1209]) );
  XOR U2456 ( .A(in[591]), .B(n3680), .Z(n2592) );
  XOR U2457 ( .A(in[246]), .B(n3777), .Z(n3237) );
  XNOR U2458 ( .A(in[1466]), .B(n3538), .Z(n3234) );
  NAND U2459 ( .A(n3237), .B(n3234), .Z(n1596) );
  XNOR U2460 ( .A(n2592), .B(n1596), .Z(out[120]) );
  OR U2461 ( .A(n1768), .B(n1597), .Z(n1598) );
  XNOR U2462 ( .A(n1767), .B(n1598), .Z(out[1210]) );
  OR U2463 ( .A(n1772), .B(n1599), .Z(n1600) );
  XNOR U2464 ( .A(n1771), .B(n1600), .Z(out[1211]) );
  OR U2465 ( .A(n1776), .B(n1601), .Z(n1602) );
  XNOR U2466 ( .A(n1775), .B(n1602), .Z(out[1212]) );
  OR U2467 ( .A(n1780), .B(n1603), .Z(n1604) );
  XNOR U2468 ( .A(n1779), .B(n1604), .Z(out[1213]) );
  OR U2469 ( .A(n1784), .B(n1605), .Z(n1606) );
  XNOR U2470 ( .A(n1783), .B(n1606), .Z(out[1214]) );
  OR U2471 ( .A(n1788), .B(n1607), .Z(n1608) );
  XNOR U2472 ( .A(n1787), .B(n1608), .Z(out[1215]) );
  OR U2473 ( .A(n4629), .B(n1609), .Z(n1610) );
  XNOR U2474 ( .A(n4628), .B(n1610), .Z(out[1216]) );
  OR U2475 ( .A(n4633), .B(n1611), .Z(n1612) );
  XNOR U2476 ( .A(n4632), .B(n1612), .Z(out[1217]) );
  OR U2477 ( .A(n4637), .B(n1613), .Z(n1614) );
  XNOR U2478 ( .A(n4636), .B(n1614), .Z(out[1218]) );
  OR U2479 ( .A(n4641), .B(n1615), .Z(n1616) );
  XNOR U2480 ( .A(n4640), .B(n1616), .Z(out[1219]) );
  XOR U2481 ( .A(in[592]), .B(n3684), .Z(n2594) );
  XOR U2482 ( .A(in[247]), .B(n3781), .Z(n3269) );
  XNOR U2483 ( .A(in[1467]), .B(n3542), .Z(n3266) );
  NAND U2484 ( .A(n3269), .B(n3266), .Z(n1617) );
  XNOR U2485 ( .A(n2594), .B(n1617), .Z(out[121]) );
  OR U2486 ( .A(n4645), .B(n1618), .Z(n1619) );
  XNOR U2487 ( .A(n4644), .B(n1619), .Z(out[1220]) );
  OR U2488 ( .A(n4649), .B(n1620), .Z(n1621) );
  XNOR U2489 ( .A(n4648), .B(n1621), .Z(out[1221]) );
  OR U2490 ( .A(n4653), .B(n1622), .Z(n1623) );
  XNOR U2491 ( .A(n4652), .B(n1623), .Z(out[1222]) );
  OR U2492 ( .A(n4657), .B(n1624), .Z(n1625) );
  XNOR U2493 ( .A(n4656), .B(n1625), .Z(out[1223]) );
  OR U2494 ( .A(n4661), .B(n1626), .Z(n1627) );
  XNOR U2495 ( .A(n4660), .B(n1627), .Z(out[1224]) );
  OR U2496 ( .A(n4665), .B(n1628), .Z(n1629) );
  XNOR U2497 ( .A(n4664), .B(n1629), .Z(out[1225]) );
  OR U2498 ( .A(n4673), .B(n1630), .Z(n1631) );
  XNOR U2499 ( .A(n4672), .B(n1631), .Z(out[1226]) );
  OR U2500 ( .A(n4677), .B(n1632), .Z(n1633) );
  XNOR U2501 ( .A(n4676), .B(n1633), .Z(out[1227]) );
  OR U2502 ( .A(n4681), .B(n1634), .Z(n1635) );
  XNOR U2503 ( .A(n4680), .B(n1635), .Z(out[1228]) );
  OR U2504 ( .A(n4685), .B(n1636), .Z(n1637) );
  XNOR U2505 ( .A(n4684), .B(n1637), .Z(out[1229]) );
  XOR U2506 ( .A(in[593]), .B(n3688), .Z(n2597) );
  XOR U2507 ( .A(in[248]), .B(n3785), .Z(n3313) );
  XNOR U2508 ( .A(in[1468]), .B(n3546), .Z(n3310) );
  NAND U2509 ( .A(n3313), .B(n3310), .Z(n1638) );
  XNOR U2510 ( .A(n2597), .B(n1638), .Z(out[122]) );
  OR U2511 ( .A(n4689), .B(n1639), .Z(n1640) );
  XNOR U2512 ( .A(n4688), .B(n1640), .Z(out[1230]) );
  OR U2513 ( .A(n4693), .B(n1641), .Z(n1642) );
  XNOR U2514 ( .A(n4692), .B(n1642), .Z(out[1231]) );
  OR U2515 ( .A(n4697), .B(n1643), .Z(n1644) );
  XNOR U2516 ( .A(n4696), .B(n1644), .Z(out[1232]) );
  OR U2517 ( .A(n4701), .B(n1645), .Z(n1646) );
  XNOR U2518 ( .A(n4700), .B(n1646), .Z(out[1233]) );
  OR U2519 ( .A(n4705), .B(n1647), .Z(n1648) );
  XNOR U2520 ( .A(n4704), .B(n1648), .Z(out[1234]) );
  OR U2521 ( .A(n4709), .B(n1649), .Z(n1650) );
  XNOR U2522 ( .A(n4708), .B(n1650), .Z(out[1235]) );
  OR U2523 ( .A(n4717), .B(n1651), .Z(n1652) );
  XNOR U2524 ( .A(n4716), .B(n1652), .Z(out[1236]) );
  OR U2525 ( .A(n4721), .B(n1653), .Z(n1654) );
  XNOR U2526 ( .A(n4720), .B(n1654), .Z(out[1237]) );
  OR U2527 ( .A(n4725), .B(n1655), .Z(n1656) );
  XNOR U2528 ( .A(n4724), .B(n1656), .Z(out[1238]) );
  OR U2529 ( .A(n4729), .B(n1657), .Z(n1658) );
  XNOR U2530 ( .A(n4728), .B(n1658), .Z(out[1239]) );
  XOR U2531 ( .A(in[594]), .B(n3692), .Z(n2599) );
  XOR U2532 ( .A(in[249]), .B(n3789), .Z(n3357) );
  XNOR U2533 ( .A(in[1469]), .B(n3550), .Z(n3354) );
  NAND U2534 ( .A(n3357), .B(n3354), .Z(n1659) );
  XNOR U2535 ( .A(n2599), .B(n1659), .Z(out[123]) );
  OR U2536 ( .A(n4733), .B(n1660), .Z(n1661) );
  XNOR U2537 ( .A(n4732), .B(n1661), .Z(out[1240]) );
  OR U2538 ( .A(n4737), .B(n1662), .Z(n1663) );
  XNOR U2539 ( .A(n4736), .B(n1663), .Z(out[1241]) );
  OR U2540 ( .A(n4741), .B(n1664), .Z(n1665) );
  XNOR U2541 ( .A(n4740), .B(n1665), .Z(out[1242]) );
  OR U2542 ( .A(n4745), .B(n1666), .Z(n1667) );
  XNOR U2543 ( .A(n4744), .B(n1667), .Z(out[1243]) );
  OR U2544 ( .A(n4749), .B(n1668), .Z(n1669) );
  XNOR U2545 ( .A(n4748), .B(n1669), .Z(out[1244]) );
  OR U2546 ( .A(n4753), .B(n1670), .Z(n1671) );
  XNOR U2547 ( .A(n4752), .B(n1671), .Z(out[1245]) );
  OR U2548 ( .A(n4761), .B(n1672), .Z(n1673) );
  XNOR U2549 ( .A(n4760), .B(n1673), .Z(out[1246]) );
  OR U2550 ( .A(n4765), .B(n1674), .Z(n1675) );
  XNOR U2551 ( .A(n4764), .B(n1675), .Z(out[1247]) );
  OR U2552 ( .A(n4769), .B(n1676), .Z(n1677) );
  XNOR U2553 ( .A(n4768), .B(n1677), .Z(out[1248]) );
  OR U2554 ( .A(n4773), .B(n1678), .Z(n1679) );
  XNOR U2555 ( .A(n4772), .B(n1679), .Z(out[1249]) );
  XOR U2556 ( .A(in[595]), .B(n3696), .Z(n2601) );
  XOR U2557 ( .A(in[250]), .B(n3793), .Z(n3403) );
  XNOR U2558 ( .A(in[1470]), .B(n3554), .Z(n3400) );
  NAND U2559 ( .A(n3403), .B(n3400), .Z(n1680) );
  XNOR U2560 ( .A(n2601), .B(n1680), .Z(out[124]) );
  OR U2561 ( .A(n4777), .B(n1681), .Z(n1682) );
  XNOR U2562 ( .A(n4776), .B(n1682), .Z(out[1250]) );
  OR U2563 ( .A(n4781), .B(n1683), .Z(n1684) );
  XNOR U2564 ( .A(n4780), .B(n1684), .Z(out[1251]) );
  OR U2565 ( .A(n4785), .B(n1685), .Z(n1686) );
  XNOR U2566 ( .A(n4784), .B(n1686), .Z(out[1252]) );
  OR U2567 ( .A(n4789), .B(n1687), .Z(n1688) );
  XNOR U2568 ( .A(n4788), .B(n1688), .Z(out[1253]) );
  OR U2569 ( .A(n4793), .B(n1689), .Z(n1690) );
  XNOR U2570 ( .A(n4792), .B(n1690), .Z(out[1254]) );
  OR U2571 ( .A(n4797), .B(n1691), .Z(n1692) );
  XNOR U2572 ( .A(n4796), .B(n1692), .Z(out[1255]) );
  ANDN U2573 ( .B(n1694), .A(n1693), .Z(n1695) );
  XNOR U2574 ( .A(n1696), .B(n1695), .Z(out[1256]) );
  ANDN U2575 ( .B(n1698), .A(n1697), .Z(n1699) );
  XNOR U2576 ( .A(n1700), .B(n1699), .Z(out[1257]) );
  ANDN U2577 ( .B(n1702), .A(n1701), .Z(n1703) );
  XNOR U2578 ( .A(n1704), .B(n1703), .Z(out[1258]) );
  ANDN U2579 ( .B(n1706), .A(n1705), .Z(n1707) );
  XNOR U2580 ( .A(n1708), .B(n1707), .Z(out[1259]) );
  XOR U2581 ( .A(in[596]), .B(n3700), .Z(n2603) );
  XNOR U2582 ( .A(in[251]), .B(n3803), .Z(n3447) );
  XNOR U2583 ( .A(in[1471]), .B(n3558), .Z(n3444) );
  NAND U2584 ( .A(n3447), .B(n3444), .Z(n1709) );
  XNOR U2585 ( .A(n2603), .B(n1709), .Z(out[125]) );
  ANDN U2586 ( .B(n1711), .A(n1710), .Z(n1712) );
  XNOR U2587 ( .A(n1713), .B(n1712), .Z(out[1260]) );
  ANDN U2588 ( .B(n1715), .A(n1714), .Z(n1716) );
  XNOR U2589 ( .A(n1717), .B(n1716), .Z(out[1261]) );
  ANDN U2590 ( .B(n1719), .A(n1718), .Z(n1720) );
  XNOR U2591 ( .A(n1721), .B(n1720), .Z(out[1262]) );
  ANDN U2592 ( .B(n1723), .A(n1722), .Z(n1724) );
  XNOR U2593 ( .A(n1725), .B(n1724), .Z(out[1263]) );
  ANDN U2594 ( .B(n1727), .A(n1726), .Z(n1728) );
  XNOR U2595 ( .A(n1729), .B(n1728), .Z(out[1264]) );
  ANDN U2596 ( .B(n1731), .A(n1730), .Z(n1732) );
  XNOR U2597 ( .A(n1733), .B(n1732), .Z(out[1265]) );
  ANDN U2598 ( .B(n1735), .A(n1734), .Z(n1736) );
  XNOR U2599 ( .A(n1737), .B(n1736), .Z(out[1266]) );
  ANDN U2600 ( .B(n1739), .A(n1738), .Z(n1740) );
  XNOR U2601 ( .A(n1741), .B(n1740), .Z(out[1267]) );
  ANDN U2602 ( .B(n1743), .A(n1742), .Z(n1744) );
  XNOR U2603 ( .A(n1745), .B(n1744), .Z(out[1268]) );
  ANDN U2604 ( .B(n1747), .A(n1746), .Z(n1748) );
  XNOR U2605 ( .A(n1749), .B(n1748), .Z(out[1269]) );
  XOR U2606 ( .A(in[597]), .B(n3704), .Z(n2605) );
  XNOR U2607 ( .A(in[252]), .B(n3807), .Z(n3491) );
  XNOR U2608 ( .A(in[1408]), .B(n3562), .Z(n3488) );
  NAND U2609 ( .A(n3491), .B(n3488), .Z(n1750) );
  XNOR U2610 ( .A(n2605), .B(n1750), .Z(out[126]) );
  ANDN U2611 ( .B(n1752), .A(n1751), .Z(n1753) );
  XNOR U2612 ( .A(n1754), .B(n1753), .Z(out[1270]) );
  ANDN U2613 ( .B(n1756), .A(n1755), .Z(n1757) );
  XNOR U2614 ( .A(n1758), .B(n1757), .Z(out[1271]) );
  ANDN U2615 ( .B(n1760), .A(n1759), .Z(n1761) );
  XNOR U2616 ( .A(n1762), .B(n1761), .Z(out[1272]) );
  ANDN U2617 ( .B(n1764), .A(n1763), .Z(n1765) );
  XNOR U2618 ( .A(n1766), .B(n1765), .Z(out[1273]) );
  ANDN U2619 ( .B(n1768), .A(n1767), .Z(n1769) );
  XNOR U2620 ( .A(n1770), .B(n1769), .Z(out[1274]) );
  ANDN U2621 ( .B(n1772), .A(n1771), .Z(n1773) );
  XNOR U2622 ( .A(n1774), .B(n1773), .Z(out[1275]) );
  ANDN U2623 ( .B(n1776), .A(n1775), .Z(n1777) );
  XNOR U2624 ( .A(n1778), .B(n1777), .Z(out[1276]) );
  ANDN U2625 ( .B(n1780), .A(n1779), .Z(n1781) );
  XNOR U2626 ( .A(n1782), .B(n1781), .Z(out[1277]) );
  ANDN U2627 ( .B(n1784), .A(n1783), .Z(n1785) );
  XNOR U2628 ( .A(n1786), .B(n1785), .Z(out[1278]) );
  ANDN U2629 ( .B(n1788), .A(n1787), .Z(n1789) );
  XNOR U2630 ( .A(n1790), .B(n1789), .Z(out[1279]) );
  XOR U2631 ( .A(in[598]), .B(n3712), .Z(n2607) );
  XNOR U2632 ( .A(in[253]), .B(n3811), .Z(n3535) );
  XNOR U2633 ( .A(in[1409]), .B(n3566), .Z(n3532) );
  NAND U2634 ( .A(n3535), .B(n3532), .Z(n1791) );
  XNOR U2635 ( .A(n2607), .B(n1791), .Z(out[127]) );
  XNOR U2636 ( .A(in[50]), .B(n3952), .Z(n1934) );
  XOR U2637 ( .A(in[1536]), .B(n3612), .Z(n2206) );
  XNOR U2638 ( .A(in[1172]), .B(n3629), .Z(n2204) );
  NAND U2639 ( .A(n2206), .B(n2204), .Z(n1792) );
  XNOR U2640 ( .A(n1934), .B(n1792), .Z(out[1280]) );
  XNOR U2641 ( .A(in[51]), .B(n3954), .Z(n1936) );
  XOR U2642 ( .A(in[1537]), .B(n3616), .Z(n2211) );
  XNOR U2643 ( .A(in[1173]), .B(n3633), .Z(n2209) );
  NAND U2644 ( .A(n2211), .B(n2209), .Z(n1793) );
  XNOR U2645 ( .A(n1936), .B(n1793), .Z(out[1281]) );
  XNOR U2646 ( .A(in[52]), .B(n3956), .Z(n1939) );
  XOR U2647 ( .A(in[1538]), .B(n3624), .Z(n2217) );
  XNOR U2648 ( .A(in[1174]), .B(n3637), .Z(n2214) );
  NAND U2649 ( .A(n2217), .B(n2214), .Z(n1794) );
  XNOR U2650 ( .A(n1939), .B(n1794), .Z(out[1282]) );
  XNOR U2651 ( .A(in[53]), .B(n3958), .Z(n1941) );
  XOR U2652 ( .A(in[1539]), .B(n3628), .Z(n2220) );
  XNOR U2653 ( .A(in[1175]), .B(n3641), .Z(n2218) );
  NAND U2654 ( .A(n2220), .B(n2218), .Z(n1795) );
  XNOR U2655 ( .A(n1941), .B(n1795), .Z(out[1283]) );
  XNOR U2656 ( .A(in[54]), .B(n3960), .Z(n1943) );
  XNOR U2657 ( .A(in[1540]), .B(n3632), .Z(n2227) );
  XNOR U2658 ( .A(in[1176]), .B(n3645), .Z(n2224) );
  NAND U2659 ( .A(n2227), .B(n2224), .Z(n1796) );
  XNOR U2660 ( .A(n1943), .B(n1796), .Z(out[1284]) );
  XNOR U2661 ( .A(in[55]), .B(n3962), .Z(n1945) );
  XNOR U2662 ( .A(in[1541]), .B(n3636), .Z(n2231) );
  XNOR U2663 ( .A(in[1177]), .B(n3649), .Z(n2228) );
  NAND U2664 ( .A(n2231), .B(n2228), .Z(n1797) );
  XNOR U2665 ( .A(n1945), .B(n1797), .Z(out[1285]) );
  XNOR U2666 ( .A(in[56]), .B(n3818), .Z(n1947) );
  XNOR U2667 ( .A(in[1542]), .B(n3640), .Z(n2235) );
  XNOR U2668 ( .A(in[1178]), .B(n3653), .Z(n2232) );
  NAND U2669 ( .A(n2235), .B(n2232), .Z(n1798) );
  XNOR U2670 ( .A(n1947), .B(n1798), .Z(out[1286]) );
  XNOR U2671 ( .A(in[57]), .B(n3820), .Z(n1949) );
  XNOR U2672 ( .A(in[1543]), .B(n3644), .Z(n2238) );
  XNOR U2673 ( .A(in[1179]), .B(n3657), .Z(n2236) );
  NAND U2674 ( .A(n2238), .B(n2236), .Z(n1799) );
  XNOR U2675 ( .A(n1949), .B(n1799), .Z(out[1287]) );
  XNOR U2676 ( .A(in[58]), .B(n3822), .Z(n1951) );
  XNOR U2677 ( .A(in[1544]), .B(n3648), .Z(n2244) );
  XNOR U2678 ( .A(in[1180]), .B(n3661), .Z(n2241) );
  NAND U2679 ( .A(n2244), .B(n2241), .Z(n1800) );
  XNOR U2680 ( .A(n1951), .B(n1800), .Z(out[1288]) );
  XNOR U2681 ( .A(in[59]), .B(n3824), .Z(n1953) );
  XNOR U2682 ( .A(in[1545]), .B(n3652), .Z(n2248) );
  XNOR U2683 ( .A(in[1181]), .B(n3669), .Z(n2245) );
  NAND U2684 ( .A(n2248), .B(n2245), .Z(n1801) );
  XNOR U2685 ( .A(n1953), .B(n1801), .Z(out[1289]) );
  XNOR U2686 ( .A(in[665]), .B(n3892), .Z(n2610) );
  XNOR U2687 ( .A(in[599]), .B(n3716), .Z(n3579) );
  NAND U2688 ( .A(n3579), .B(n3577), .Z(n1802) );
  XNOR U2689 ( .A(n2610), .B(n1802), .Z(out[128]) );
  XNOR U2690 ( .A(in[60]), .B(n3826), .Z(n1955) );
  XNOR U2691 ( .A(in[1546]), .B(n3656), .Z(n2252) );
  XNOR U2692 ( .A(in[1182]), .B(n3673), .Z(n2249) );
  NAND U2693 ( .A(n2252), .B(n2249), .Z(n1803) );
  XNOR U2694 ( .A(n1955), .B(n1803), .Z(out[1290]) );
  XNOR U2695 ( .A(in[61]), .B(n3828), .Z(n1957) );
  XNOR U2696 ( .A(in[1547]), .B(n3660), .Z(n2256) );
  XNOR U2697 ( .A(in[1183]), .B(n3677), .Z(n2253) );
  NAND U2698 ( .A(n2256), .B(n2253), .Z(n1804) );
  XNOR U2699 ( .A(n1957), .B(n1804), .Z(out[1291]) );
  XNOR U2700 ( .A(in[62]), .B(n3834), .Z(n1960) );
  XNOR U2701 ( .A(in[1548]), .B(n3668), .Z(n2260) );
  XNOR U2702 ( .A(in[1184]), .B(n3681), .Z(n2257) );
  NAND U2703 ( .A(n2260), .B(n2257), .Z(n1805) );
  XNOR U2704 ( .A(n1960), .B(n1805), .Z(out[1292]) );
  XNOR U2705 ( .A(in[63]), .B(n3836), .Z(n1962) );
  XNOR U2706 ( .A(in[1549]), .B(n3672), .Z(n2264) );
  XNOR U2707 ( .A(in[1185]), .B(n3685), .Z(n2261) );
  NAND U2708 ( .A(n2264), .B(n2261), .Z(n1806) );
  XNOR U2709 ( .A(n1962), .B(n1806), .Z(out[1293]) );
  XNOR U2710 ( .A(in[0]), .B(n3838), .Z(n1964) );
  XNOR U2711 ( .A(in[1550]), .B(n3676), .Z(n2269) );
  XOR U2712 ( .A(n3689), .B(in[1186]), .Z(n2266) );
  NAND U2713 ( .A(n2269), .B(n2266), .Z(n1807) );
  XNOR U2714 ( .A(n1964), .B(n1807), .Z(out[1294]) );
  XNOR U2715 ( .A(in[1]), .B(n3840), .Z(n1966) );
  XNOR U2716 ( .A(in[1551]), .B(n3680), .Z(n2272) );
  XOR U2717 ( .A(n3693), .B(in[1187]), .Z(n2270) );
  NAND U2718 ( .A(n2272), .B(n2270), .Z(n1808) );
  XNOR U2719 ( .A(n1966), .B(n1808), .Z(out[1295]) );
  XNOR U2720 ( .A(in[2]), .B(n3842), .Z(n1968) );
  XNOR U2721 ( .A(in[1552]), .B(n3684), .Z(n2278) );
  XOR U2722 ( .A(n3697), .B(in[1188]), .Z(n2275) );
  NAND U2723 ( .A(n2278), .B(n2275), .Z(n1809) );
  XNOR U2724 ( .A(n1968), .B(n1809), .Z(out[1296]) );
  XNOR U2725 ( .A(in[3]), .B(n3844), .Z(n1970) );
  XNOR U2726 ( .A(in[1553]), .B(n3688), .Z(n2282) );
  XOR U2727 ( .A(n3701), .B(in[1189]), .Z(n2279) );
  NAND U2728 ( .A(n2282), .B(n2279), .Z(n1810) );
  XNOR U2729 ( .A(n1970), .B(n1810), .Z(out[1297]) );
  XNOR U2730 ( .A(in[4]), .B(n3846), .Z(n1972) );
  XNOR U2731 ( .A(in[1554]), .B(n3692), .Z(n2286) );
  XNOR U2732 ( .A(in[1190]), .B(n3705), .Z(n2283) );
  NAND U2733 ( .A(n2286), .B(n2283), .Z(n1811) );
  XNOR U2734 ( .A(n1972), .B(n1811), .Z(out[1298]) );
  XNOR U2735 ( .A(in[5]), .B(n3848), .Z(n1974) );
  XNOR U2736 ( .A(in[1555]), .B(n3696), .Z(n2290) );
  XNOR U2737 ( .A(in[1191]), .B(n3713), .Z(n2287) );
  NAND U2738 ( .A(n2290), .B(n2287), .Z(n1812) );
  XNOR U2739 ( .A(n1974), .B(n1812), .Z(out[1299]) );
  XNOR U2740 ( .A(in[666]), .B(n3894), .Z(n2612) );
  XNOR U2741 ( .A(in[600]), .B(n3720), .Z(n3623) );
  XOR U2742 ( .A(in[255]), .B(n3537), .Z(n3621) );
  NAND U2743 ( .A(n3623), .B(n3621), .Z(n1813) );
  XNOR U2744 ( .A(n2612), .B(n1813), .Z(out[129]) );
  XOR U2745 ( .A(in[202]), .B(n3585), .Z(n3971) );
  XNOR U2746 ( .A(in[1422]), .B(n3626), .Z(n3970) );
  XOR U2747 ( .A(in[1045]), .B(n4126), .Z(n2638) );
  NAND U2748 ( .A(n3970), .B(n2638), .Z(n1814) );
  XNOR U2749 ( .A(n3971), .B(n1814), .Z(out[12]) );
  XNOR U2750 ( .A(in[6]), .B(n3850), .Z(n1976) );
  XNOR U2751 ( .A(in[1556]), .B(n3700), .Z(n2294) );
  XNOR U2752 ( .A(in[1192]), .B(n3717), .Z(n2291) );
  NAND U2753 ( .A(n2294), .B(n2291), .Z(n1815) );
  XNOR U2754 ( .A(n1976), .B(n1815), .Z(out[1300]) );
  XNOR U2755 ( .A(in[7]), .B(n3852), .Z(n1978) );
  XNOR U2756 ( .A(in[1557]), .B(n3704), .Z(n2298) );
  XNOR U2757 ( .A(in[1193]), .B(n3721), .Z(n2295) );
  NAND U2758 ( .A(n2298), .B(n2295), .Z(n1816) );
  XNOR U2759 ( .A(n1978), .B(n1816), .Z(out[1301]) );
  XNOR U2760 ( .A(in[8]), .B(n3856), .Z(n1981) );
  XNOR U2761 ( .A(in[1558]), .B(n3712), .Z(n2302) );
  XNOR U2762 ( .A(in[1194]), .B(n3725), .Z(n2299) );
  NAND U2763 ( .A(n2302), .B(n2299), .Z(n1817) );
  XNOR U2764 ( .A(n1981), .B(n1817), .Z(out[1302]) );
  XNOR U2765 ( .A(in[9]), .B(n3858), .Z(n1983) );
  XNOR U2766 ( .A(in[1559]), .B(n3716), .Z(n2306) );
  XNOR U2767 ( .A(in[1195]), .B(n3729), .Z(n2303) );
  NAND U2768 ( .A(n2306), .B(n2303), .Z(n1818) );
  XNOR U2769 ( .A(n1983), .B(n1818), .Z(out[1303]) );
  XNOR U2770 ( .A(in[10]), .B(n3860), .Z(n1985) );
  XNOR U2771 ( .A(in[1560]), .B(n3720), .Z(n2311) );
  XNOR U2772 ( .A(in[1196]), .B(n3733), .Z(n2308) );
  NAND U2773 ( .A(n2311), .B(n2308), .Z(n1819) );
  XNOR U2774 ( .A(n1985), .B(n1819), .Z(out[1304]) );
  XNOR U2775 ( .A(in[11]), .B(n3862), .Z(n1987) );
  XNOR U2776 ( .A(in[1561]), .B(n3724), .Z(n2315) );
  XNOR U2777 ( .A(in[1197]), .B(n3737), .Z(n2312) );
  NAND U2778 ( .A(n2315), .B(n2312), .Z(n1820) );
  XNOR U2779 ( .A(n1987), .B(n1820), .Z(out[1305]) );
  XNOR U2780 ( .A(in[12]), .B(n3864), .Z(n1989) );
  XNOR U2781 ( .A(in[1562]), .B(n3728), .Z(n2319) );
  XNOR U2782 ( .A(in[1198]), .B(n3741), .Z(n2316) );
  NAND U2783 ( .A(n2319), .B(n2316), .Z(n1821) );
  XNOR U2784 ( .A(n1989), .B(n1821), .Z(out[1306]) );
  XNOR U2785 ( .A(in[13]), .B(n3866), .Z(n1991) );
  XNOR U2786 ( .A(in[1563]), .B(n3732), .Z(n2323) );
  XNOR U2787 ( .A(in[1199]), .B(n3745), .Z(n2320) );
  NAND U2788 ( .A(n2323), .B(n2320), .Z(n1822) );
  XNOR U2789 ( .A(n1991), .B(n1822), .Z(out[1307]) );
  XNOR U2790 ( .A(in[14]), .B(n3868), .Z(n1993) );
  XNOR U2791 ( .A(in[1564]), .B(n3736), .Z(n2327) );
  XNOR U2792 ( .A(in[1200]), .B(n3749), .Z(n2324) );
  NAND U2793 ( .A(n2327), .B(n2324), .Z(n1823) );
  XNOR U2794 ( .A(n1993), .B(n1823), .Z(out[1308]) );
  XNOR U2795 ( .A(in[15]), .B(n3870), .Z(n1995) );
  XNOR U2796 ( .A(in[1565]), .B(n3740), .Z(n2331) );
  XNOR U2797 ( .A(in[1201]), .B(n3757), .Z(n2328) );
  NAND U2798 ( .A(n2331), .B(n2328), .Z(n1824) );
  XNOR U2799 ( .A(n1995), .B(n1824), .Z(out[1309]) );
  XNOR U2800 ( .A(in[667]), .B(n3896), .Z(n2615) );
  XNOR U2801 ( .A(in[601]), .B(n3724), .Z(n3667) );
  XOR U2802 ( .A(in[192]), .B(n3541), .Z(n3664) );
  NAND U2803 ( .A(n3667), .B(n3664), .Z(n1825) );
  XNOR U2804 ( .A(n2615), .B(n1825), .Z(out[130]) );
  XNOR U2805 ( .A(in[16]), .B(n3872), .Z(n1997) );
  XNOR U2806 ( .A(in[1566]), .B(n3744), .Z(n2335) );
  XNOR U2807 ( .A(in[1202]), .B(n3761), .Z(n2332) );
  NAND U2808 ( .A(n2335), .B(n2332), .Z(n1826) );
  XNOR U2809 ( .A(n1997), .B(n1826), .Z(out[1310]) );
  XNOR U2810 ( .A(in[17]), .B(n3874), .Z(n1999) );
  XNOR U2811 ( .A(in[1567]), .B(n3748), .Z(n2338) );
  XNOR U2812 ( .A(in[1203]), .B(n3765), .Z(n2336) );
  NAND U2813 ( .A(n2338), .B(n2336), .Z(n1827) );
  XNOR U2814 ( .A(n1999), .B(n1827), .Z(out[1311]) );
  XNOR U2815 ( .A(in[18]), .B(n3878), .Z(n2002) );
  XNOR U2816 ( .A(in[1568]), .B(n3756), .Z(n2344) );
  XNOR U2817 ( .A(in[1204]), .B(n3769), .Z(n2341) );
  NAND U2818 ( .A(n2344), .B(n2341), .Z(n1828) );
  XNOR U2819 ( .A(n2002), .B(n1828), .Z(out[1312]) );
  XNOR U2820 ( .A(in[19]), .B(n3880), .Z(n2004) );
  XNOR U2821 ( .A(in[1569]), .B(n3760), .Z(n2348) );
  XNOR U2822 ( .A(in[1205]), .B(n3773), .Z(n2345) );
  NAND U2823 ( .A(n2348), .B(n2345), .Z(n1829) );
  XNOR U2824 ( .A(n2004), .B(n1829), .Z(out[1313]) );
  XNOR U2825 ( .A(in[20]), .B(n3882), .Z(n2006) );
  XNOR U2826 ( .A(in[1570]), .B(n3764), .Z(n2353) );
  XNOR U2827 ( .A(in[1206]), .B(n3777), .Z(n2350) );
  NAND U2828 ( .A(n2353), .B(n2350), .Z(n1830) );
  XNOR U2829 ( .A(n2006), .B(n1830), .Z(out[1314]) );
  XNOR U2830 ( .A(in[21]), .B(n3884), .Z(n2008) );
  XNOR U2831 ( .A(in[1571]), .B(n3768), .Z(n2357) );
  XNOR U2832 ( .A(in[1207]), .B(n3781), .Z(n2354) );
  NAND U2833 ( .A(n2357), .B(n2354), .Z(n1831) );
  XNOR U2834 ( .A(n2008), .B(n1831), .Z(out[1315]) );
  XNOR U2835 ( .A(in[22]), .B(n3886), .Z(n2010) );
  XNOR U2836 ( .A(in[1572]), .B(n3772), .Z(n2361) );
  XNOR U2837 ( .A(in[1208]), .B(n3785), .Z(n2358) );
  NAND U2838 ( .A(n2361), .B(n2358), .Z(n1832) );
  XNOR U2839 ( .A(n2010), .B(n1832), .Z(out[1316]) );
  XNOR U2840 ( .A(in[23]), .B(n3888), .Z(n2012) );
  XOR U2841 ( .A(in[1573]), .B(n3776), .Z(n2365) );
  XNOR U2842 ( .A(in[1209]), .B(n3789), .Z(n2362) );
  NAND U2843 ( .A(n2365), .B(n2362), .Z(n1833) );
  XNOR U2844 ( .A(n2012), .B(n1833), .Z(out[1317]) );
  XNOR U2845 ( .A(in[24]), .B(n3890), .Z(n2014) );
  XOR U2846 ( .A(in[1574]), .B(n3780), .Z(n2369) );
  XNOR U2847 ( .A(in[1210]), .B(n3793), .Z(n2366) );
  NAND U2848 ( .A(n2369), .B(n2366), .Z(n1834) );
  XNOR U2849 ( .A(n2014), .B(n1834), .Z(out[1318]) );
  XNOR U2850 ( .A(in[25]), .B(n3892), .Z(n2016) );
  XOR U2851 ( .A(in[1575]), .B(n3784), .Z(n2373) );
  XOR U2852 ( .A(in[1211]), .B(n3803), .Z(n2370) );
  NAND U2853 ( .A(n2373), .B(n2370), .Z(n1835) );
  XNOR U2854 ( .A(n2016), .B(n1835), .Z(out[1319]) );
  XNOR U2855 ( .A(in[668]), .B(n3900), .Z(n2617) );
  XNOR U2856 ( .A(in[602]), .B(n3728), .Z(n3711) );
  XOR U2857 ( .A(in[193]), .B(n3545), .Z(n3708) );
  NAND U2858 ( .A(n3711), .B(n3708), .Z(n1836) );
  XNOR U2859 ( .A(n2617), .B(n1836), .Z(out[131]) );
  XNOR U2860 ( .A(in[26]), .B(n3894), .Z(n2018) );
  XOR U2861 ( .A(in[1576]), .B(n3788), .Z(n2377) );
  XOR U2862 ( .A(in[1212]), .B(n3807), .Z(n2374) );
  NAND U2863 ( .A(n2377), .B(n2374), .Z(n1837) );
  XNOR U2864 ( .A(n2018), .B(n1837), .Z(out[1320]) );
  XNOR U2865 ( .A(in[27]), .B(n3896), .Z(n2020) );
  XOR U2866 ( .A(in[1577]), .B(n3792), .Z(n2381) );
  XOR U2867 ( .A(in[1213]), .B(n3811), .Z(n2378) );
  NAND U2868 ( .A(n2381), .B(n2378), .Z(n1838) );
  XNOR U2869 ( .A(n2020), .B(n1838), .Z(out[1321]) );
  XNOR U2870 ( .A(in[28]), .B(n3900), .Z(n2023) );
  XOR U2871 ( .A(in[1578]), .B(n3802), .Z(n2385) );
  XNOR U2872 ( .A(in[1214]), .B(n3815), .Z(n2382) );
  NAND U2873 ( .A(n2385), .B(n2382), .Z(n1839) );
  XNOR U2874 ( .A(n2023), .B(n1839), .Z(out[1322]) );
  XNOR U2875 ( .A(in[29]), .B(n3902), .Z(n2025) );
  XOR U2876 ( .A(in[1579]), .B(n3806), .Z(n2389) );
  XOR U2877 ( .A(in[1215]), .B(n3537), .Z(n2386) );
  NAND U2878 ( .A(n2389), .B(n2386), .Z(n1840) );
  XNOR U2879 ( .A(n2025), .B(n1840), .Z(out[1323]) );
  XNOR U2880 ( .A(in[30]), .B(n3904), .Z(n2027) );
  XOR U2881 ( .A(in[1580]), .B(n3810), .Z(n2394) );
  XOR U2882 ( .A(in[1152]), .B(n3541), .Z(n2391) );
  NAND U2883 ( .A(n2394), .B(n2391), .Z(n1841) );
  XNOR U2884 ( .A(n2027), .B(n1841), .Z(out[1324]) );
  XNOR U2885 ( .A(in[31]), .B(n3906), .Z(n2029) );
  XOR U2886 ( .A(in[1581]), .B(n3814), .Z(n2398) );
  XOR U2887 ( .A(in[1153]), .B(n3545), .Z(n2395) );
  NAND U2888 ( .A(n2398), .B(n2395), .Z(n1842) );
  XNOR U2889 ( .A(n2029), .B(n1842), .Z(out[1325]) );
  XNOR U2890 ( .A(in[32]), .B(n3908), .Z(n2031) );
  XOR U2891 ( .A(in[1582]), .B(n3536), .Z(n2402) );
  XOR U2892 ( .A(in[1154]), .B(n3549), .Z(n2399) );
  NAND U2893 ( .A(n2402), .B(n2399), .Z(n1843) );
  XNOR U2894 ( .A(n2031), .B(n1843), .Z(out[1326]) );
  XNOR U2895 ( .A(in[33]), .B(n3910), .Z(n2033) );
  XOR U2896 ( .A(in[1583]), .B(n3540), .Z(n2406) );
  XOR U2897 ( .A(in[1155]), .B(n3553), .Z(n2403) );
  NAND U2898 ( .A(n2406), .B(n2403), .Z(n1844) );
  XNOR U2899 ( .A(n2033), .B(n1844), .Z(out[1327]) );
  XNOR U2900 ( .A(in[34]), .B(n3912), .Z(n2035) );
  XOR U2901 ( .A(in[1584]), .B(n3544), .Z(n2410) );
  XOR U2902 ( .A(in[1156]), .B(n3557), .Z(n2407) );
  NAND U2903 ( .A(n2410), .B(n2407), .Z(n1845) );
  XNOR U2904 ( .A(n2035), .B(n1845), .Z(out[1328]) );
  XNOR U2905 ( .A(in[35]), .B(n3914), .Z(n2037) );
  XOR U2906 ( .A(in[1585]), .B(n3548), .Z(n2414) );
  XOR U2907 ( .A(in[1157]), .B(n3561), .Z(n2411) );
  NAND U2908 ( .A(n2414), .B(n2411), .Z(n1846) );
  XNOR U2909 ( .A(n2037), .B(n1846), .Z(out[1329]) );
  XNOR U2910 ( .A(in[669]), .B(n3902), .Z(n2620) );
  XNOR U2911 ( .A(in[603]), .B(n3732), .Z(n3755) );
  XOR U2912 ( .A(in[194]), .B(n3549), .Z(n3752) );
  NAND U2913 ( .A(n3755), .B(n3752), .Z(n1847) );
  XNOR U2914 ( .A(n2620), .B(n1847), .Z(out[132]) );
  XNOR U2915 ( .A(in[36]), .B(n3916), .Z(n2039) );
  XOR U2916 ( .A(in[1586]), .B(n3552), .Z(n2418) );
  XOR U2917 ( .A(in[1158]), .B(n3565), .Z(n2415) );
  NAND U2918 ( .A(n2418), .B(n2415), .Z(n1848) );
  XNOR U2919 ( .A(n2039), .B(n1848), .Z(out[1330]) );
  XNOR U2920 ( .A(in[37]), .B(n3918), .Z(n2041) );
  XOR U2921 ( .A(in[1587]), .B(n3556), .Z(n2422) );
  XOR U2922 ( .A(in[1159]), .B(n3569), .Z(n2419) );
  NAND U2923 ( .A(n2422), .B(n2419), .Z(n1849) );
  XNOR U2924 ( .A(n2041), .B(n1849), .Z(out[1331]) );
  XNOR U2925 ( .A(in[38]), .B(n3924), .Z(n2044) );
  XOR U2926 ( .A(in[1588]), .B(n3560), .Z(n2426) );
  XOR U2927 ( .A(in[1160]), .B(n3573), .Z(n2423) );
  NAND U2928 ( .A(n2426), .B(n2423), .Z(n1850) );
  XNOR U2929 ( .A(n2044), .B(n1850), .Z(out[1332]) );
  XNOR U2930 ( .A(in[39]), .B(n3926), .Z(n2046) );
  XOR U2931 ( .A(in[1589]), .B(n3564), .Z(n2430) );
  XOR U2932 ( .A(in[1161]), .B(n3581), .Z(n2427) );
  NAND U2933 ( .A(n2430), .B(n2427), .Z(n1851) );
  XNOR U2934 ( .A(n2046), .B(n1851), .Z(out[1333]) );
  XNOR U2935 ( .A(in[40]), .B(n3928), .Z(n2048) );
  XOR U2936 ( .A(in[1590]), .B(n3568), .Z(n2435) );
  XOR U2937 ( .A(in[1162]), .B(n3585), .Z(n2432) );
  NAND U2938 ( .A(n2435), .B(n2432), .Z(n1852) );
  XNOR U2939 ( .A(n2048), .B(n1852), .Z(out[1334]) );
  XNOR U2940 ( .A(in[41]), .B(n3930), .Z(n2050) );
  XOR U2941 ( .A(in[1591]), .B(n3572), .Z(n2439) );
  XOR U2942 ( .A(in[1163]), .B(n3589), .Z(n2436) );
  NAND U2943 ( .A(n2439), .B(n2436), .Z(n1853) );
  XNOR U2944 ( .A(n2050), .B(n1853), .Z(out[1335]) );
  XNOR U2945 ( .A(in[42]), .B(n3932), .Z(n2052) );
  XOR U2946 ( .A(in[1592]), .B(n3580), .Z(n2443) );
  XOR U2947 ( .A(in[1164]), .B(n3593), .Z(n2440) );
  NAND U2948 ( .A(n2443), .B(n2440), .Z(n1854) );
  XNOR U2949 ( .A(n2052), .B(n1854), .Z(out[1336]) );
  XNOR U2950 ( .A(in[43]), .B(n3934), .Z(n2054) );
  XOR U2951 ( .A(in[1593]), .B(n3584), .Z(n2447) );
  XOR U2952 ( .A(in[1165]), .B(n3597), .Z(n2444) );
  NAND U2953 ( .A(n2447), .B(n2444), .Z(n1855) );
  XNOR U2954 ( .A(n2054), .B(n1855), .Z(out[1337]) );
  XNOR U2955 ( .A(in[44]), .B(n3936), .Z(n2056) );
  XOR U2956 ( .A(in[1594]), .B(n3588), .Z(n2451) );
  XOR U2957 ( .A(in[1166]), .B(n3601), .Z(n2448) );
  NAND U2958 ( .A(n2451), .B(n2448), .Z(n1856) );
  XNOR U2959 ( .A(n2056), .B(n1856), .Z(out[1338]) );
  XNOR U2960 ( .A(in[45]), .B(n3938), .Z(n2058) );
  XOR U2961 ( .A(in[1595]), .B(n3592), .Z(n2455) );
  XOR U2962 ( .A(in[1167]), .B(n3605), .Z(n2452) );
  NAND U2963 ( .A(n2455), .B(n2452), .Z(n1857) );
  XNOR U2964 ( .A(n2058), .B(n1857), .Z(out[1339]) );
  XNOR U2965 ( .A(in[670]), .B(n3904), .Z(n2622) );
  XNOR U2966 ( .A(in[604]), .B(n3736), .Z(n3799) );
  XOR U2967 ( .A(in[195]), .B(n3553), .Z(n3796) );
  NAND U2968 ( .A(n3799), .B(n3796), .Z(n1858) );
  XNOR U2969 ( .A(n2622), .B(n1858), .Z(out[133]) );
  XNOR U2970 ( .A(in[46]), .B(n3940), .Z(n2060) );
  XOR U2971 ( .A(in[1596]), .B(n3596), .Z(n2459) );
  XOR U2972 ( .A(in[1168]), .B(n3609), .Z(n2456) );
  NAND U2973 ( .A(n2459), .B(n2456), .Z(n1859) );
  XNOR U2974 ( .A(n2060), .B(n1859), .Z(out[1340]) );
  XNOR U2975 ( .A(in[47]), .B(n3942), .Z(n2062) );
  XOR U2976 ( .A(in[1597]), .B(n3600), .Z(n2463) );
  XOR U2977 ( .A(in[1169]), .B(n3613), .Z(n2460) );
  NAND U2978 ( .A(n2463), .B(n2460), .Z(n1860) );
  XNOR U2979 ( .A(n2062), .B(n1860), .Z(out[1341]) );
  XNOR U2980 ( .A(in[48]), .B(n3948), .Z(n2065) );
  XOR U2981 ( .A(in[1598]), .B(n3604), .Z(n2467) );
  XOR U2982 ( .A(in[1170]), .B(n3617), .Z(n2464) );
  NAND U2983 ( .A(n2467), .B(n2464), .Z(n1861) );
  XNOR U2984 ( .A(n2065), .B(n1861), .Z(out[1342]) );
  XNOR U2985 ( .A(in[49]), .B(n3950), .Z(n2067) );
  XOR U2986 ( .A(in[1599]), .B(n3608), .Z(n2470) );
  XNOR U2987 ( .A(in[1171]), .B(n3625), .Z(n2468) );
  NAND U2988 ( .A(n2470), .B(n2468), .Z(n1862) );
  XNOR U2989 ( .A(n2067), .B(n1862), .Z(out[1343]) );
  XOR U2990 ( .A(in[427]), .B(n3980), .Z(n2069) );
  NOR U2991 ( .A(n1934), .B(n2206), .Z(n1863) );
  XNOR U2992 ( .A(n2069), .B(n1863), .Z(out[1344]) );
  XOR U2993 ( .A(in[428]), .B(n3983), .Z(n2071) );
  NOR U2994 ( .A(n1936), .B(n2211), .Z(n1864) );
  XNOR U2995 ( .A(n2071), .B(n1864), .Z(out[1345]) );
  XOR U2996 ( .A(in[429]), .B(n3986), .Z(n2073) );
  NOR U2997 ( .A(n1939), .B(n2217), .Z(n1865) );
  XNOR U2998 ( .A(n2073), .B(n1865), .Z(out[1346]) );
  XOR U2999 ( .A(in[430]), .B(n3989), .Z(n2075) );
  NOR U3000 ( .A(n1941), .B(n2220), .Z(n1866) );
  XNOR U3001 ( .A(n2075), .B(n1866), .Z(out[1347]) );
  XOR U3002 ( .A(in[431]), .B(n3992), .Z(n2077) );
  NOR U3003 ( .A(n1943), .B(n2227), .Z(n1867) );
  XNOR U3004 ( .A(n2077), .B(n1867), .Z(out[1348]) );
  XOR U3005 ( .A(in[432]), .B(n3995), .Z(n2079) );
  NOR U3006 ( .A(n1945), .B(n2231), .Z(n1868) );
  XNOR U3007 ( .A(n2079), .B(n1868), .Z(out[1349]) );
  XNOR U3008 ( .A(in[671]), .B(n3906), .Z(n2624) );
  XNOR U3009 ( .A(in[605]), .B(n3740), .Z(n3833) );
  XOR U3010 ( .A(in[196]), .B(n3557), .Z(n3830) );
  NAND U3011 ( .A(n3833), .B(n3830), .Z(n1869) );
  XNOR U3012 ( .A(n2624), .B(n1869), .Z(out[134]) );
  XOR U3013 ( .A(in[433]), .B(n3998), .Z(n2081) );
  NOR U3014 ( .A(n1947), .B(n2235), .Z(n1870) );
  XNOR U3015 ( .A(n2081), .B(n1870), .Z(out[1350]) );
  XOR U3016 ( .A(in[434]), .B(n4001), .Z(n2083) );
  NOR U3017 ( .A(n1949), .B(n2238), .Z(n1871) );
  XNOR U3018 ( .A(n2083), .B(n1871), .Z(out[1351]) );
  XOR U3019 ( .A(in[435]), .B(n4008), .Z(n2086) );
  NOR U3020 ( .A(n1951), .B(n2244), .Z(n1872) );
  XNOR U3021 ( .A(n2086), .B(n1872), .Z(out[1352]) );
  XOR U3022 ( .A(in[436]), .B(n4011), .Z(n2088) );
  NOR U3023 ( .A(n1953), .B(n2248), .Z(n1873) );
  XNOR U3024 ( .A(n2088), .B(n1873), .Z(out[1353]) );
  XOR U3025 ( .A(in[437]), .B(n4014), .Z(n2090) );
  NOR U3026 ( .A(n1955), .B(n2252), .Z(n1874) );
  XNOR U3027 ( .A(n2090), .B(n1874), .Z(out[1354]) );
  XOR U3028 ( .A(in[438]), .B(n4017), .Z(n2092) );
  NOR U3029 ( .A(n1957), .B(n2256), .Z(n1875) );
  XNOR U3030 ( .A(n2092), .B(n1875), .Z(out[1355]) );
  XOR U3031 ( .A(in[439]), .B(n4020), .Z(n2094) );
  NOR U3032 ( .A(n1960), .B(n2260), .Z(n1876) );
  XNOR U3033 ( .A(n2094), .B(n1876), .Z(out[1356]) );
  XOR U3034 ( .A(in[440]), .B(n4023), .Z(n2096) );
  NOR U3035 ( .A(n1962), .B(n2264), .Z(n1877) );
  XNOR U3036 ( .A(n2096), .B(n1877), .Z(out[1357]) );
  XOR U3037 ( .A(in[441]), .B(n4026), .Z(n2098) );
  NOR U3038 ( .A(n1964), .B(n2269), .Z(n1878) );
  XNOR U3039 ( .A(n2098), .B(n1878), .Z(out[1358]) );
  XOR U3040 ( .A(in[442]), .B(n4029), .Z(n2100) );
  NOR U3041 ( .A(n1966), .B(n2272), .Z(n1879) );
  XNOR U3042 ( .A(n2100), .B(n1879), .Z(out[1359]) );
  XNOR U3043 ( .A(in[672]), .B(n3908), .Z(n2626) );
  XNOR U3044 ( .A(in[606]), .B(n3744), .Z(n3855) );
  XOR U3045 ( .A(in[197]), .B(n3561), .Z(n4079) );
  NAND U3046 ( .A(n3855), .B(n4079), .Z(n1880) );
  XNOR U3047 ( .A(n2626), .B(n1880), .Z(out[135]) );
  XOR U3048 ( .A(in[443]), .B(n4032), .Z(n2102) );
  NOR U3049 ( .A(n1968), .B(n2278), .Z(n1881) );
  XNOR U3050 ( .A(n2102), .B(n1881), .Z(out[1360]) );
  XOR U3051 ( .A(in[444]), .B(n4035), .Z(n2104) );
  NOR U3052 ( .A(n1970), .B(n2282), .Z(n1882) );
  XNOR U3053 ( .A(n2104), .B(n1882), .Z(out[1361]) );
  XOR U3054 ( .A(in[445]), .B(n4042), .Z(n2107) );
  NOR U3055 ( .A(n1972), .B(n2286), .Z(n1883) );
  XNOR U3056 ( .A(n2107), .B(n1883), .Z(out[1362]) );
  XOR U3057 ( .A(in[446]), .B(n4045), .Z(n2109) );
  NOR U3058 ( .A(n1974), .B(n2290), .Z(n1884) );
  XNOR U3059 ( .A(n2109), .B(n1884), .Z(out[1363]) );
  XOR U3060 ( .A(in[447]), .B(n4048), .Z(n2111) );
  NOR U3061 ( .A(n1976), .B(n2294), .Z(n1885) );
  XNOR U3062 ( .A(n2111), .B(n1885), .Z(out[1364]) );
  XOR U3063 ( .A(in[384]), .B(n4051), .Z(n2113) );
  NOR U3064 ( .A(n1978), .B(n2298), .Z(n1886) );
  XNOR U3065 ( .A(n2113), .B(n1886), .Z(out[1365]) );
  XOR U3066 ( .A(in[385]), .B(n4054), .Z(n2115) );
  NOR U3067 ( .A(n1981), .B(n2302), .Z(n1887) );
  XNOR U3068 ( .A(n2115), .B(n1887), .Z(out[1366]) );
  XOR U3069 ( .A(in[386]), .B(n4057), .Z(n2117) );
  NOR U3070 ( .A(n1983), .B(n2306), .Z(n1888) );
  XNOR U3071 ( .A(n2117), .B(n1888), .Z(out[1367]) );
  XOR U3072 ( .A(in[387]), .B(n4060), .Z(n2119) );
  NOR U3073 ( .A(n1985), .B(n2311), .Z(n1889) );
  XNOR U3074 ( .A(n2119), .B(n1889), .Z(out[1368]) );
  XOR U3075 ( .A(in[388]), .B(n4063), .Z(n2121) );
  NOR U3076 ( .A(n1987), .B(n2315), .Z(n1890) );
  XNOR U3077 ( .A(n2121), .B(n1890), .Z(out[1369]) );
  XNOR U3078 ( .A(in[673]), .B(n3910), .Z(n2628) );
  XNOR U3079 ( .A(in[607]), .B(n3748), .Z(n3877) );
  XOR U3080 ( .A(in[198]), .B(n3565), .Z(n4363) );
  NAND U3081 ( .A(n3877), .B(n4363), .Z(n1891) );
  XNOR U3082 ( .A(n2628), .B(n1891), .Z(out[136]) );
  XOR U3083 ( .A(in[389]), .B(n4066), .Z(n2123) );
  NOR U3084 ( .A(n1989), .B(n2319), .Z(n1892) );
  XNOR U3085 ( .A(n2123), .B(n1892), .Z(out[1370]) );
  XOR U3086 ( .A(in[390]), .B(n4069), .Z(n2125) );
  NOR U3087 ( .A(n1991), .B(n2323), .Z(n1893) );
  XNOR U3088 ( .A(n2125), .B(n1893), .Z(out[1371]) );
  XOR U3089 ( .A(in[391]), .B(n4080), .Z(n2129) );
  NOR U3090 ( .A(n1993), .B(n2327), .Z(n1894) );
  XNOR U3091 ( .A(n2129), .B(n1894), .Z(out[1372]) );
  XOR U3092 ( .A(in[392]), .B(n4083), .Z(n2131) );
  NOR U3093 ( .A(n1995), .B(n2331), .Z(n1895) );
  XNOR U3094 ( .A(n2131), .B(n1895), .Z(out[1373]) );
  XOR U3095 ( .A(in[393]), .B(n4086), .Z(n2133) );
  NOR U3096 ( .A(n1997), .B(n2335), .Z(n1896) );
  XNOR U3097 ( .A(n2133), .B(n1896), .Z(out[1374]) );
  XOR U3098 ( .A(in[394]), .B(n4089), .Z(n2135) );
  NOR U3099 ( .A(n1999), .B(n2338), .Z(n1897) );
  XNOR U3100 ( .A(n2135), .B(n1897), .Z(out[1375]) );
  XOR U3101 ( .A(in[395]), .B(n4092), .Z(n2137) );
  NOR U3102 ( .A(n2002), .B(n2344), .Z(n1898) );
  XNOR U3103 ( .A(n2137), .B(n1898), .Z(out[1376]) );
  XNOR U3104 ( .A(n4095), .B(in[396]), .Z(n2139) );
  NOR U3105 ( .A(n2004), .B(n2348), .Z(n1899) );
  XNOR U3106 ( .A(n2139), .B(n1899), .Z(out[1377]) );
  XNOR U3107 ( .A(n4098), .B(in[397]), .Z(n2141) );
  NOR U3108 ( .A(n2006), .B(n2353), .Z(n1900) );
  XNOR U3109 ( .A(n2141), .B(n1900), .Z(out[1378]) );
  XNOR U3110 ( .A(n4101), .B(in[398]), .Z(n2143) );
  NOR U3111 ( .A(n2008), .B(n2357), .Z(n1901) );
  XNOR U3112 ( .A(n2143), .B(n1901), .Z(out[1379]) );
  XNOR U3113 ( .A(in[674]), .B(n3912), .Z(n2630) );
  XNOR U3114 ( .A(in[608]), .B(n3756), .Z(n3899) );
  XOR U3115 ( .A(in[199]), .B(n3569), .Z(n4807) );
  NAND U3116 ( .A(n3899), .B(n4807), .Z(n1902) );
  XNOR U3117 ( .A(n2630), .B(n1902), .Z(out[137]) );
  XNOR U3118 ( .A(n4104), .B(in[399]), .Z(n2145) );
  NOR U3119 ( .A(n2010), .B(n2361), .Z(n1903) );
  XNOR U3120 ( .A(n2145), .B(n1903), .Z(out[1380]) );
  XNOR U3121 ( .A(n4107), .B(in[400]), .Z(n2147) );
  NOR U3122 ( .A(n2012), .B(n2365), .Z(n1904) );
  XNOR U3123 ( .A(n2147), .B(n1904), .Z(out[1381]) );
  XNOR U3124 ( .A(n4114), .B(in[401]), .Z(n2150) );
  NOR U3125 ( .A(n2014), .B(n2369), .Z(n1905) );
  XNOR U3126 ( .A(n2150), .B(n1905), .Z(out[1382]) );
  XNOR U3127 ( .A(n4117), .B(in[402]), .Z(n2152) );
  NOR U3128 ( .A(n2016), .B(n2373), .Z(n1906) );
  XNOR U3129 ( .A(n2152), .B(n1906), .Z(out[1383]) );
  XNOR U3130 ( .A(n4120), .B(in[403]), .Z(n2154) );
  NOR U3131 ( .A(n2018), .B(n2377), .Z(n1907) );
  XNOR U3132 ( .A(n2154), .B(n1907), .Z(out[1384]) );
  XNOR U3133 ( .A(in[404]), .B(n4123), .Z(n2156) );
  NOR U3134 ( .A(n2020), .B(n2381), .Z(n1908) );
  XNOR U3135 ( .A(n2156), .B(n1908), .Z(out[1385]) );
  XNOR U3136 ( .A(in[405]), .B(n4126), .Z(n2158) );
  NOR U3137 ( .A(n2023), .B(n2385), .Z(n1909) );
  XNOR U3138 ( .A(n2158), .B(n1909), .Z(out[1386]) );
  XNOR U3139 ( .A(in[406]), .B(n4129), .Z(n2160) );
  NOR U3140 ( .A(n2025), .B(n2389), .Z(n1910) );
  XNOR U3141 ( .A(n2160), .B(n1910), .Z(out[1387]) );
  XNOR U3142 ( .A(in[407]), .B(n4132), .Z(n2162) );
  NOR U3143 ( .A(n2027), .B(n2394), .Z(n1911) );
  XNOR U3144 ( .A(n2162), .B(n1911), .Z(out[1388]) );
  XNOR U3145 ( .A(in[408]), .B(n4135), .Z(n2164) );
  NOR U3146 ( .A(n2029), .B(n2398), .Z(n1912) );
  XNOR U3147 ( .A(n2164), .B(n1912), .Z(out[1389]) );
  XNOR U3148 ( .A(in[675]), .B(n3914), .Z(n2633) );
  XNOR U3149 ( .A(in[609]), .B(n3760), .Z(n3923) );
  NAND U3150 ( .A(n3923), .B(n3921), .Z(n1913) );
  XNOR U3151 ( .A(n2633), .B(n1913), .Z(out[138]) );
  XNOR U3152 ( .A(in[409]), .B(n4138), .Z(n2166) );
  NOR U3153 ( .A(n2031), .B(n2402), .Z(n1914) );
  XNOR U3154 ( .A(n2166), .B(n1914), .Z(out[1390]) );
  XNOR U3155 ( .A(in[410]), .B(n4141), .Z(n2168) );
  NOR U3156 ( .A(n2033), .B(n2406), .Z(n1915) );
  XNOR U3157 ( .A(n2168), .B(n1915), .Z(out[1391]) );
  XNOR U3158 ( .A(in[411]), .B(n4148), .Z(n2171) );
  NOR U3159 ( .A(n2035), .B(n2410), .Z(n1916) );
  XNOR U3160 ( .A(n2171), .B(n1916), .Z(out[1392]) );
  XNOR U3161 ( .A(in[412]), .B(n4151), .Z(n2173) );
  NOR U3162 ( .A(n2037), .B(n2414), .Z(n1917) );
  XNOR U3163 ( .A(n2173), .B(n1917), .Z(out[1393]) );
  XNOR U3164 ( .A(in[413]), .B(n4154), .Z(n2175) );
  NOR U3165 ( .A(n2039), .B(n2418), .Z(n1918) );
  XNOR U3166 ( .A(n2175), .B(n1918), .Z(out[1394]) );
  XNOR U3167 ( .A(in[414]), .B(n4157), .Z(n2177) );
  NOR U3168 ( .A(n2041), .B(n2422), .Z(n1919) );
  XNOR U3169 ( .A(n2177), .B(n1919), .Z(out[1395]) );
  XNOR U3170 ( .A(in[415]), .B(n4160), .Z(n2179) );
  NOR U3171 ( .A(n2044), .B(n2426), .Z(n1920) );
  XNOR U3172 ( .A(n2179), .B(n1920), .Z(out[1396]) );
  XNOR U3173 ( .A(in[416]), .B(n4163), .Z(n2181) );
  NOR U3174 ( .A(n2046), .B(n2430), .Z(n1921) );
  XNOR U3175 ( .A(n2181), .B(n1921), .Z(out[1397]) );
  XNOR U3176 ( .A(in[417]), .B(n4166), .Z(n2183) );
  NOR U3177 ( .A(n2048), .B(n2435), .Z(n1922) );
  XNOR U3178 ( .A(n2183), .B(n1922), .Z(out[1398]) );
  XNOR U3179 ( .A(in[418]), .B(n4169), .Z(n2185) );
  NOR U3180 ( .A(n2050), .B(n2439), .Z(n1923) );
  XNOR U3181 ( .A(n2185), .B(n1923), .Z(out[1399]) );
  XNOR U3182 ( .A(in[676]), .B(n3916), .Z(n2636) );
  XNOR U3183 ( .A(in[610]), .B(n3764), .Z(n3947) );
  NAND U3184 ( .A(n3947), .B(n3945), .Z(n1924) );
  XNOR U3185 ( .A(n2636), .B(n1924), .Z(out[139]) );
  XOR U3186 ( .A(in[203]), .B(n3589), .Z(n4005) );
  XNOR U3187 ( .A(in[1423]), .B(n3630), .Z(n4004) );
  XOR U3188 ( .A(in[1046]), .B(n4129), .Z(n2641) );
  NAND U3189 ( .A(n4004), .B(n2641), .Z(n1925) );
  XNOR U3190 ( .A(n4005), .B(n1925), .Z(out[13]) );
  XNOR U3191 ( .A(in[419]), .B(n4172), .Z(n2187) );
  NOR U3192 ( .A(n2052), .B(n2443), .Z(n1926) );
  XNOR U3193 ( .A(n2187), .B(n1926), .Z(out[1400]) );
  XOR U3194 ( .A(in[420]), .B(n4175), .Z(n2189) );
  NOR U3195 ( .A(n2054), .B(n2447), .Z(n1927) );
  XNOR U3196 ( .A(n2189), .B(n1927), .Z(out[1401]) );
  XOR U3197 ( .A(in[421]), .B(n4182), .Z(n2192) );
  NOR U3198 ( .A(n2056), .B(n2451), .Z(n1928) );
  XNOR U3199 ( .A(n2192), .B(n1928), .Z(out[1402]) );
  XOR U3200 ( .A(in[422]), .B(n4185), .Z(n2194) );
  NOR U3201 ( .A(n2058), .B(n2455), .Z(n1929) );
  XNOR U3202 ( .A(n2194), .B(n1929), .Z(out[1403]) );
  XOR U3203 ( .A(in[423]), .B(n3964), .Z(n2196) );
  NOR U3204 ( .A(n2060), .B(n2459), .Z(n1930) );
  XNOR U3205 ( .A(n2196), .B(n1930), .Z(out[1404]) );
  XOR U3206 ( .A(in[424]), .B(n3967), .Z(n2198) );
  NOR U3207 ( .A(n2062), .B(n2463), .Z(n1931) );
  XNOR U3208 ( .A(n2198), .B(n1931), .Z(out[1405]) );
  XOR U3209 ( .A(in[425]), .B(n3974), .Z(n2200) );
  NOR U3210 ( .A(n2065), .B(n2467), .Z(n1932) );
  XNOR U3211 ( .A(n2200), .B(n1932), .Z(out[1406]) );
  XOR U3212 ( .A(in[426]), .B(n3977), .Z(n2202) );
  NOR U3213 ( .A(n2067), .B(n2470), .Z(n1933) );
  XNOR U3214 ( .A(n2202), .B(n1933), .Z(out[1407]) );
  XOR U3215 ( .A(in[789]), .B(n3654), .Z(n2205) );
  NAND U3216 ( .A(n2069), .B(n1934), .Z(n1935) );
  XNOR U3217 ( .A(n2205), .B(n1935), .Z(out[1408]) );
  XOR U3218 ( .A(in[790]), .B(n3658), .Z(n2210) );
  NAND U3219 ( .A(n2071), .B(n1936), .Z(n1937) );
  XNOR U3220 ( .A(n2210), .B(n1937), .Z(out[1409]) );
  XNOR U3221 ( .A(in[677]), .B(n3918), .Z(n2639) );
  XNOR U3222 ( .A(in[611]), .B(n3768), .Z(n3973) );
  NAND U3223 ( .A(n3973), .B(n3971), .Z(n1938) );
  XNOR U3224 ( .A(n2639), .B(n1938), .Z(out[140]) );
  XOR U3225 ( .A(in[791]), .B(n3662), .Z(n2215) );
  NAND U3226 ( .A(n2073), .B(n1939), .Z(n1940) );
  XNOR U3227 ( .A(n2215), .B(n1940), .Z(out[1410]) );
  XOR U3228 ( .A(in[792]), .B(n3670), .Z(n2219) );
  NAND U3229 ( .A(n2075), .B(n1941), .Z(n1942) );
  XNOR U3230 ( .A(n2219), .B(n1942), .Z(out[1411]) );
  XOR U3231 ( .A(in[793]), .B(n3674), .Z(n2225) );
  NAND U3232 ( .A(n2077), .B(n1943), .Z(n1944) );
  XNOR U3233 ( .A(n2225), .B(n1944), .Z(out[1412]) );
  XOR U3234 ( .A(in[794]), .B(n3678), .Z(n2229) );
  NAND U3235 ( .A(n2079), .B(n1945), .Z(n1946) );
  XNOR U3236 ( .A(n2229), .B(n1946), .Z(out[1413]) );
  XOR U3237 ( .A(in[795]), .B(n3682), .Z(n2233) );
  NAND U3238 ( .A(n2081), .B(n1947), .Z(n1948) );
  XNOR U3239 ( .A(n2233), .B(n1948), .Z(out[1414]) );
  XOR U3240 ( .A(in[796]), .B(n3686), .Z(n2237) );
  NAND U3241 ( .A(n2083), .B(n1949), .Z(n1950) );
  XNOR U3242 ( .A(n2237), .B(n1950), .Z(out[1415]) );
  XOR U3243 ( .A(in[797]), .B(n3690), .Z(n2242) );
  NAND U3244 ( .A(n2086), .B(n1951), .Z(n1952) );
  XNOR U3245 ( .A(n2242), .B(n1952), .Z(out[1416]) );
  XOR U3246 ( .A(in[798]), .B(n3694), .Z(n2246) );
  NAND U3247 ( .A(n2088), .B(n1953), .Z(n1954) );
  XNOR U3248 ( .A(n2246), .B(n1954), .Z(out[1417]) );
  XOR U3249 ( .A(in[799]), .B(n3698), .Z(n2250) );
  NAND U3250 ( .A(n2090), .B(n1955), .Z(n1956) );
  XNOR U3251 ( .A(n2250), .B(n1956), .Z(out[1418]) );
  XOR U3252 ( .A(in[800]), .B(n3702), .Z(n2254) );
  NAND U3253 ( .A(n2092), .B(n1957), .Z(n1958) );
  XNOR U3254 ( .A(n2254), .B(n1958), .Z(out[1419]) );
  XNOR U3255 ( .A(in[678]), .B(n3924), .Z(n2642) );
  XNOR U3256 ( .A(in[612]), .B(n3772), .Z(n4007) );
  NAND U3257 ( .A(n4007), .B(n4005), .Z(n1959) );
  XNOR U3258 ( .A(n2642), .B(n1959), .Z(out[141]) );
  XOR U3259 ( .A(in[801]), .B(n3706), .Z(n2258) );
  NAND U3260 ( .A(n2094), .B(n1960), .Z(n1961) );
  XNOR U3261 ( .A(n2258), .B(n1961), .Z(out[1420]) );
  XOR U3262 ( .A(in[802]), .B(n3714), .Z(n2262) );
  NAND U3263 ( .A(n2096), .B(n1962), .Z(n1963) );
  XNOR U3264 ( .A(n2262), .B(n1963), .Z(out[1421]) );
  XOR U3265 ( .A(in[803]), .B(n3718), .Z(n2267) );
  NAND U3266 ( .A(n2098), .B(n1964), .Z(n1965) );
  XNOR U3267 ( .A(n2267), .B(n1965), .Z(out[1422]) );
  XOR U3268 ( .A(in[804]), .B(n3722), .Z(n2271) );
  NAND U3269 ( .A(n2100), .B(n1966), .Z(n1967) );
  XNOR U3270 ( .A(n2271), .B(n1967), .Z(out[1423]) );
  XOR U3271 ( .A(in[805]), .B(n3726), .Z(n2276) );
  NAND U3272 ( .A(n2102), .B(n1968), .Z(n1969) );
  XNOR U3273 ( .A(n2276), .B(n1969), .Z(out[1424]) );
  XNOR U3274 ( .A(in[806]), .B(n3730), .Z(n2280) );
  NAND U3275 ( .A(n2104), .B(n1970), .Z(n1971) );
  XNOR U3276 ( .A(n2280), .B(n1971), .Z(out[1425]) );
  XNOR U3277 ( .A(in[807]), .B(n3734), .Z(n2284) );
  NAND U3278 ( .A(n2107), .B(n1972), .Z(n1973) );
  XNOR U3279 ( .A(n2284), .B(n1973), .Z(out[1426]) );
  XNOR U3280 ( .A(in[808]), .B(n3738), .Z(n2288) );
  NAND U3281 ( .A(n2109), .B(n1974), .Z(n1975) );
  XNOR U3282 ( .A(n2288), .B(n1975), .Z(out[1427]) );
  XNOR U3283 ( .A(in[809]), .B(n3742), .Z(n2292) );
  NAND U3284 ( .A(n2111), .B(n1976), .Z(n1977) );
  XNOR U3285 ( .A(n2292), .B(n1977), .Z(out[1428]) );
  XNOR U3286 ( .A(in[810]), .B(n3746), .Z(n2296) );
  NAND U3287 ( .A(n2113), .B(n1978), .Z(n1979) );
  XNOR U3288 ( .A(n2296), .B(n1979), .Z(out[1429]) );
  XNOR U3289 ( .A(in[679]), .B(n3926), .Z(n2646) );
  XOR U3290 ( .A(in[613]), .B(n3776), .Z(n4041) );
  XOR U3291 ( .A(in[204]), .B(n3593), .Z(n4039) );
  NAND U3292 ( .A(n4041), .B(n4039), .Z(n1980) );
  XNOR U3293 ( .A(n2646), .B(n1980), .Z(out[142]) );
  XNOR U3294 ( .A(in[811]), .B(n3750), .Z(n2300) );
  NAND U3295 ( .A(n2115), .B(n1981), .Z(n1982) );
  XNOR U3296 ( .A(n2300), .B(n1982), .Z(out[1430]) );
  XNOR U3297 ( .A(in[812]), .B(n3758), .Z(n2304) );
  NAND U3298 ( .A(n2117), .B(n1983), .Z(n1984) );
  XNOR U3299 ( .A(n2304), .B(n1984), .Z(out[1431]) );
  XNOR U3300 ( .A(in[813]), .B(n3762), .Z(n2309) );
  NAND U3301 ( .A(n2119), .B(n1985), .Z(n1986) );
  XNOR U3302 ( .A(n2309), .B(n1986), .Z(out[1432]) );
  XNOR U3303 ( .A(in[814]), .B(n3766), .Z(n2313) );
  NAND U3304 ( .A(n2121), .B(n1987), .Z(n1988) );
  XNOR U3305 ( .A(n2313), .B(n1988), .Z(out[1433]) );
  XNOR U3306 ( .A(in[815]), .B(n3770), .Z(n2317) );
  NAND U3307 ( .A(n2123), .B(n1989), .Z(n1990) );
  XNOR U3308 ( .A(n2317), .B(n1990), .Z(out[1434]) );
  XNOR U3309 ( .A(in[816]), .B(n3774), .Z(n2321) );
  NAND U3310 ( .A(n2125), .B(n1991), .Z(n1992) );
  XNOR U3311 ( .A(n2321), .B(n1992), .Z(out[1435]) );
  XNOR U3312 ( .A(in[817]), .B(n3778), .Z(n2325) );
  NAND U3313 ( .A(n2129), .B(n1993), .Z(n1994) );
  XNOR U3314 ( .A(n2325), .B(n1994), .Z(out[1436]) );
  XNOR U3315 ( .A(in[818]), .B(n3782), .Z(n2329) );
  NAND U3316 ( .A(n2131), .B(n1995), .Z(n1996) );
  XNOR U3317 ( .A(n2329), .B(n1996), .Z(out[1437]) );
  XNOR U3318 ( .A(in[819]), .B(n3786), .Z(n2333) );
  NAND U3319 ( .A(n2133), .B(n1997), .Z(n1998) );
  XNOR U3320 ( .A(n2333), .B(n1998), .Z(out[1438]) );
  XNOR U3321 ( .A(in[820]), .B(n3790), .Z(n2337) );
  NAND U3322 ( .A(n2135), .B(n1999), .Z(n2000) );
  XNOR U3323 ( .A(n2337), .B(n2000), .Z(out[1439]) );
  XNOR U3324 ( .A(in[680]), .B(n3928), .Z(n2649) );
  XOR U3325 ( .A(in[614]), .B(n3780), .Z(n4075) );
  XOR U3326 ( .A(in[205]), .B(n3597), .Z(n4073) );
  NAND U3327 ( .A(n4075), .B(n4073), .Z(n2001) );
  XNOR U3328 ( .A(n2649), .B(n2001), .Z(out[143]) );
  XNOR U3329 ( .A(in[821]), .B(n3794), .Z(n2342) );
  NAND U3330 ( .A(n2137), .B(n2002), .Z(n2003) );
  XNOR U3331 ( .A(n2342), .B(n2003), .Z(out[1440]) );
  XNOR U3332 ( .A(in[822]), .B(n3804), .Z(n2346) );
  NAND U3333 ( .A(n2139), .B(n2004), .Z(n2005) );
  XNOR U3334 ( .A(n2346), .B(n2005), .Z(out[1441]) );
  XNOR U3335 ( .A(in[823]), .B(n3808), .Z(n2351) );
  NAND U3336 ( .A(n2141), .B(n2006), .Z(n2007) );
  XNOR U3337 ( .A(n2351), .B(n2007), .Z(out[1442]) );
  XNOR U3338 ( .A(in[824]), .B(n3812), .Z(n2355) );
  NAND U3339 ( .A(n2143), .B(n2008), .Z(n2009) );
  XNOR U3340 ( .A(n2355), .B(n2009), .Z(out[1443]) );
  XNOR U3341 ( .A(in[825]), .B(n3816), .Z(n2359) );
  NAND U3342 ( .A(n2145), .B(n2010), .Z(n2011) );
  XNOR U3343 ( .A(n2359), .B(n2011), .Z(out[1444]) );
  XNOR U3344 ( .A(in[826]), .B(n3538), .Z(n2363) );
  NAND U3345 ( .A(n2147), .B(n2012), .Z(n2013) );
  XNOR U3346 ( .A(n2363), .B(n2013), .Z(out[1445]) );
  XNOR U3347 ( .A(in[827]), .B(n3542), .Z(n2367) );
  NAND U3348 ( .A(n2150), .B(n2014), .Z(n2015) );
  XNOR U3349 ( .A(n2367), .B(n2015), .Z(out[1446]) );
  XNOR U3350 ( .A(in[828]), .B(n3546), .Z(n2371) );
  NAND U3351 ( .A(n2152), .B(n2016), .Z(n2017) );
  XNOR U3352 ( .A(n2371), .B(n2017), .Z(out[1447]) );
  XNOR U3353 ( .A(in[829]), .B(n3550), .Z(n2375) );
  NAND U3354 ( .A(n2154), .B(n2018), .Z(n2019) );
  XNOR U3355 ( .A(n2375), .B(n2019), .Z(out[1448]) );
  XNOR U3356 ( .A(in[830]), .B(n3554), .Z(n2379) );
  NAND U3357 ( .A(n2156), .B(n2020), .Z(n2021) );
  XNOR U3358 ( .A(n2379), .B(n2021), .Z(out[1449]) );
  XNOR U3359 ( .A(in[681]), .B(n3930), .Z(n2652) );
  XOR U3360 ( .A(in[615]), .B(n3784), .Z(n4113) );
  XOR U3361 ( .A(in[206]), .B(n3601), .Z(n4111) );
  NAND U3362 ( .A(n4113), .B(n4111), .Z(n2022) );
  XNOR U3363 ( .A(n2652), .B(n2022), .Z(out[144]) );
  XNOR U3364 ( .A(in[831]), .B(n3558), .Z(n2383) );
  NAND U3365 ( .A(n2158), .B(n2023), .Z(n2024) );
  XNOR U3366 ( .A(n2383), .B(n2024), .Z(out[1450]) );
  XNOR U3367 ( .A(in[768]), .B(n3562), .Z(n2387) );
  NAND U3368 ( .A(n2160), .B(n2025), .Z(n2026) );
  XNOR U3369 ( .A(n2387), .B(n2026), .Z(out[1451]) );
  XNOR U3370 ( .A(in[769]), .B(n3566), .Z(n2392) );
  NAND U3371 ( .A(n2162), .B(n2027), .Z(n2028) );
  XNOR U3372 ( .A(n2392), .B(n2028), .Z(out[1452]) );
  XOR U3373 ( .A(n3570), .B(in[770]), .Z(n2396) );
  NAND U3374 ( .A(n2164), .B(n2029), .Z(n2030) );
  XNOR U3375 ( .A(n2396), .B(n2030), .Z(out[1453]) );
  XOR U3376 ( .A(n3574), .B(in[771]), .Z(n2400) );
  NAND U3377 ( .A(n2166), .B(n2031), .Z(n2032) );
  XNOR U3378 ( .A(n2400), .B(n2032), .Z(out[1454]) );
  XOR U3379 ( .A(n3582), .B(in[772]), .Z(n2404) );
  NAND U3380 ( .A(n2168), .B(n2033), .Z(n2034) );
  XNOR U3381 ( .A(n2404), .B(n2034), .Z(out[1455]) );
  XOR U3382 ( .A(n3586), .B(in[773]), .Z(n2408) );
  NAND U3383 ( .A(n2171), .B(n2035), .Z(n2036) );
  XNOR U3384 ( .A(n2408), .B(n2036), .Z(out[1456]) );
  XOR U3385 ( .A(n3590), .B(in[774]), .Z(n2412) );
  NAND U3386 ( .A(n2173), .B(n2037), .Z(n2038) );
  XNOR U3387 ( .A(n2412), .B(n2038), .Z(out[1457]) );
  XOR U3388 ( .A(n3594), .B(in[775]), .Z(n2416) );
  NAND U3389 ( .A(n2175), .B(n2039), .Z(n2040) );
  XNOR U3390 ( .A(n2416), .B(n2040), .Z(out[1458]) );
  XOR U3391 ( .A(n3598), .B(in[776]), .Z(n2420) );
  NAND U3392 ( .A(n2177), .B(n2041), .Z(n2042) );
  XNOR U3393 ( .A(n2420), .B(n2042), .Z(out[1459]) );
  XNOR U3394 ( .A(in[682]), .B(n3932), .Z(n2655) );
  XOR U3395 ( .A(in[616]), .B(n3788), .Z(n4147) );
  XOR U3396 ( .A(in[207]), .B(n3605), .Z(n4145) );
  NAND U3397 ( .A(n4147), .B(n4145), .Z(n2043) );
  XNOR U3398 ( .A(n2655), .B(n2043), .Z(out[145]) );
  XOR U3399 ( .A(in[777]), .B(n3602), .Z(n2424) );
  NAND U3400 ( .A(n2179), .B(n2044), .Z(n2045) );
  XNOR U3401 ( .A(n2424), .B(n2045), .Z(out[1460]) );
  XOR U3402 ( .A(n3606), .B(in[778]), .Z(n2428) );
  NAND U3403 ( .A(n2181), .B(n2046), .Z(n2047) );
  XNOR U3404 ( .A(n2428), .B(n2047), .Z(out[1461]) );
  XOR U3405 ( .A(n3610), .B(in[779]), .Z(n2433) );
  NAND U3406 ( .A(n2183), .B(n2048), .Z(n2049) );
  XNOR U3407 ( .A(n2433), .B(n2049), .Z(out[1462]) );
  XOR U3408 ( .A(in[780]), .B(n3614), .Z(n2437) );
  NAND U3409 ( .A(n2185), .B(n2050), .Z(n2051) );
  XNOR U3410 ( .A(n2437), .B(n2051), .Z(out[1463]) );
  XOR U3411 ( .A(in[781]), .B(n3618), .Z(n2441) );
  NAND U3412 ( .A(n2187), .B(n2052), .Z(n2053) );
  XNOR U3413 ( .A(n2441), .B(n2053), .Z(out[1464]) );
  XOR U3414 ( .A(in[782]), .B(n3626), .Z(n2445) );
  NAND U3415 ( .A(n2189), .B(n2054), .Z(n2055) );
  XNOR U3416 ( .A(n2445), .B(n2055), .Z(out[1465]) );
  XOR U3417 ( .A(in[783]), .B(n3630), .Z(n2449) );
  NAND U3418 ( .A(n2192), .B(n2056), .Z(n2057) );
  XNOR U3419 ( .A(n2449), .B(n2057), .Z(out[1466]) );
  XOR U3420 ( .A(in[784]), .B(n3634), .Z(n2453) );
  NAND U3421 ( .A(n2194), .B(n2058), .Z(n2059) );
  XNOR U3422 ( .A(n2453), .B(n2059), .Z(out[1467]) );
  XOR U3423 ( .A(in[785]), .B(n3638), .Z(n2457) );
  NAND U3424 ( .A(n2196), .B(n2060), .Z(n2061) );
  XNOR U3425 ( .A(n2457), .B(n2061), .Z(out[1468]) );
  XOR U3426 ( .A(in[786]), .B(n3642), .Z(n2461) );
  NAND U3427 ( .A(n2198), .B(n2062), .Z(n2063) );
  XNOR U3428 ( .A(n2461), .B(n2063), .Z(out[1469]) );
  XNOR U3429 ( .A(in[683]), .B(n3934), .Z(n2658) );
  XOR U3430 ( .A(in[617]), .B(n3792), .Z(n4181) );
  XOR U3431 ( .A(in[208]), .B(n3609), .Z(n4179) );
  NAND U3432 ( .A(n4181), .B(n4179), .Z(n2064) );
  XNOR U3433 ( .A(n2658), .B(n2064), .Z(out[146]) );
  XOR U3434 ( .A(in[787]), .B(n3646), .Z(n2465) );
  NAND U3435 ( .A(n2200), .B(n2065), .Z(n2066) );
  XNOR U3436 ( .A(n2465), .B(n2066), .Z(out[1470]) );
  XOR U3437 ( .A(in[788]), .B(n3650), .Z(n2469) );
  NAND U3438 ( .A(n2202), .B(n2067), .Z(n2068) );
  XNOR U3439 ( .A(n2469), .B(n2068), .Z(out[1471]) );
  OR U3440 ( .A(n2205), .B(n2069), .Z(n2070) );
  XNOR U3441 ( .A(n2204), .B(n2070), .Z(out[1472]) );
  OR U3442 ( .A(n2210), .B(n2071), .Z(n2072) );
  XNOR U3443 ( .A(n2209), .B(n2072), .Z(out[1473]) );
  OR U3444 ( .A(n2215), .B(n2073), .Z(n2074) );
  XNOR U3445 ( .A(n2214), .B(n2074), .Z(out[1474]) );
  OR U3446 ( .A(n2219), .B(n2075), .Z(n2076) );
  XNOR U3447 ( .A(n2218), .B(n2076), .Z(out[1475]) );
  OR U3448 ( .A(n2225), .B(n2077), .Z(n2078) );
  XNOR U3449 ( .A(n2224), .B(n2078), .Z(out[1476]) );
  OR U3450 ( .A(n2229), .B(n2079), .Z(n2080) );
  XNOR U3451 ( .A(n2228), .B(n2080), .Z(out[1477]) );
  OR U3452 ( .A(n2233), .B(n2081), .Z(n2082) );
  XNOR U3453 ( .A(n2232), .B(n2082), .Z(out[1478]) );
  OR U3454 ( .A(n2237), .B(n2083), .Z(n2084) );
  XNOR U3455 ( .A(n2236), .B(n2084), .Z(out[1479]) );
  XNOR U3456 ( .A(in[684]), .B(n3936), .Z(n2661) );
  XOR U3457 ( .A(in[618]), .B(n3802), .Z(n4207) );
  XOR U3458 ( .A(in[209]), .B(n3613), .Z(n4205) );
  NAND U3459 ( .A(n4207), .B(n4205), .Z(n2085) );
  XNOR U3460 ( .A(n2661), .B(n2085), .Z(out[147]) );
  OR U3461 ( .A(n2242), .B(n2086), .Z(n2087) );
  XNOR U3462 ( .A(n2241), .B(n2087), .Z(out[1480]) );
  OR U3463 ( .A(n2246), .B(n2088), .Z(n2089) );
  XNOR U3464 ( .A(n2245), .B(n2089), .Z(out[1481]) );
  OR U3465 ( .A(n2250), .B(n2090), .Z(n2091) );
  XNOR U3466 ( .A(n2249), .B(n2091), .Z(out[1482]) );
  OR U3467 ( .A(n2254), .B(n2092), .Z(n2093) );
  XNOR U3468 ( .A(n2253), .B(n2093), .Z(out[1483]) );
  OR U3469 ( .A(n2258), .B(n2094), .Z(n2095) );
  XNOR U3470 ( .A(n2257), .B(n2095), .Z(out[1484]) );
  OR U3471 ( .A(n2262), .B(n2096), .Z(n2097) );
  XNOR U3472 ( .A(n2261), .B(n2097), .Z(out[1485]) );
  OR U3473 ( .A(n2267), .B(n2098), .Z(n2099) );
  XNOR U3474 ( .A(n2266), .B(n2099), .Z(out[1486]) );
  OR U3475 ( .A(n2271), .B(n2100), .Z(n2101) );
  XNOR U3476 ( .A(n2270), .B(n2101), .Z(out[1487]) );
  OR U3477 ( .A(n2276), .B(n2102), .Z(n2103) );
  XNOR U3478 ( .A(n2275), .B(n2103), .Z(out[1488]) );
  OR U3479 ( .A(n2280), .B(n2104), .Z(n2105) );
  XNOR U3480 ( .A(n2279), .B(n2105), .Z(out[1489]) );
  XNOR U3481 ( .A(in[685]), .B(n3938), .Z(n2664) );
  XOR U3482 ( .A(in[619]), .B(n3806), .Z(n4231) );
  XOR U3483 ( .A(in[210]), .B(n3617), .Z(n4229) );
  NAND U3484 ( .A(n4231), .B(n4229), .Z(n2106) );
  XNOR U3485 ( .A(n2664), .B(n2106), .Z(out[148]) );
  OR U3486 ( .A(n2284), .B(n2107), .Z(n2108) );
  XNOR U3487 ( .A(n2283), .B(n2108), .Z(out[1490]) );
  OR U3488 ( .A(n2288), .B(n2109), .Z(n2110) );
  XNOR U3489 ( .A(n2287), .B(n2110), .Z(out[1491]) );
  OR U3490 ( .A(n2292), .B(n2111), .Z(n2112) );
  XNOR U3491 ( .A(n2291), .B(n2112), .Z(out[1492]) );
  OR U3492 ( .A(n2296), .B(n2113), .Z(n2114) );
  XNOR U3493 ( .A(n2295), .B(n2114), .Z(out[1493]) );
  OR U3494 ( .A(n2300), .B(n2115), .Z(n2116) );
  XNOR U3495 ( .A(n2299), .B(n2116), .Z(out[1494]) );
  OR U3496 ( .A(n2304), .B(n2117), .Z(n2118) );
  XNOR U3497 ( .A(n2303), .B(n2118), .Z(out[1495]) );
  OR U3498 ( .A(n2309), .B(n2119), .Z(n2120) );
  XNOR U3499 ( .A(n2308), .B(n2120), .Z(out[1496]) );
  OR U3500 ( .A(n2313), .B(n2121), .Z(n2122) );
  XNOR U3501 ( .A(n2312), .B(n2122), .Z(out[1497]) );
  OR U3502 ( .A(n2317), .B(n2123), .Z(n2124) );
  XNOR U3503 ( .A(n2316), .B(n2124), .Z(out[1498]) );
  OR U3504 ( .A(n2321), .B(n2125), .Z(n2126) );
  XNOR U3505 ( .A(n2320), .B(n2126), .Z(out[1499]) );
  XNOR U3506 ( .A(in[686]), .B(n3940), .Z(n2666) );
  XOR U3507 ( .A(in[620]), .B(n3810), .Z(n4255) );
  XNOR U3508 ( .A(in[211]), .B(n3625), .Z(n4253) );
  NAND U3509 ( .A(n4255), .B(n4253), .Z(n2127) );
  XNOR U3510 ( .A(n2666), .B(n2127), .Z(out[149]) );
  XNOR U3511 ( .A(in[1424]), .B(n3634), .Z(n4038) );
  XOR U3512 ( .A(in[1047]), .B(n4132), .Z(n2645) );
  NAND U3513 ( .A(n4038), .B(n2645), .Z(n2128) );
  XNOR U3514 ( .A(n4039), .B(n2128), .Z(out[14]) );
  OR U3515 ( .A(n2325), .B(n2129), .Z(n2130) );
  XNOR U3516 ( .A(n2324), .B(n2130), .Z(out[1500]) );
  OR U3517 ( .A(n2329), .B(n2131), .Z(n2132) );
  XNOR U3518 ( .A(n2328), .B(n2132), .Z(out[1501]) );
  OR U3519 ( .A(n2333), .B(n2133), .Z(n2134) );
  XNOR U3520 ( .A(n2332), .B(n2134), .Z(out[1502]) );
  OR U3521 ( .A(n2337), .B(n2135), .Z(n2136) );
  XNOR U3522 ( .A(n2336), .B(n2136), .Z(out[1503]) );
  OR U3523 ( .A(n2342), .B(n2137), .Z(n2138) );
  XNOR U3524 ( .A(n2341), .B(n2138), .Z(out[1504]) );
  OR U3525 ( .A(n2346), .B(n2139), .Z(n2140) );
  XNOR U3526 ( .A(n2345), .B(n2140), .Z(out[1505]) );
  OR U3527 ( .A(n2351), .B(n2141), .Z(n2142) );
  XNOR U3528 ( .A(n2350), .B(n2142), .Z(out[1506]) );
  OR U3529 ( .A(n2355), .B(n2143), .Z(n2144) );
  XNOR U3530 ( .A(n2354), .B(n2144), .Z(out[1507]) );
  OR U3531 ( .A(n2359), .B(n2145), .Z(n2146) );
  XNOR U3532 ( .A(n2358), .B(n2146), .Z(out[1508]) );
  OR U3533 ( .A(n2363), .B(n2147), .Z(n2148) );
  XNOR U3534 ( .A(n2362), .B(n2148), .Z(out[1509]) );
  XNOR U3535 ( .A(in[687]), .B(n3942), .Z(n2669) );
  XOR U3536 ( .A(in[621]), .B(n3814), .Z(n4279) );
  XNOR U3537 ( .A(in[212]), .B(n3629), .Z(n4277) );
  NAND U3538 ( .A(n4279), .B(n4277), .Z(n2149) );
  XNOR U3539 ( .A(n2669), .B(n2149), .Z(out[150]) );
  OR U3540 ( .A(n2367), .B(n2150), .Z(n2151) );
  XNOR U3541 ( .A(n2366), .B(n2151), .Z(out[1510]) );
  OR U3542 ( .A(n2371), .B(n2152), .Z(n2153) );
  XNOR U3543 ( .A(n2370), .B(n2153), .Z(out[1511]) );
  OR U3544 ( .A(n2375), .B(n2154), .Z(n2155) );
  XNOR U3545 ( .A(n2374), .B(n2155), .Z(out[1512]) );
  OR U3546 ( .A(n2379), .B(n2156), .Z(n2157) );
  XNOR U3547 ( .A(n2378), .B(n2157), .Z(out[1513]) );
  OR U3548 ( .A(n2383), .B(n2158), .Z(n2159) );
  XNOR U3549 ( .A(n2382), .B(n2159), .Z(out[1514]) );
  OR U3550 ( .A(n2387), .B(n2160), .Z(n2161) );
  XNOR U3551 ( .A(n2386), .B(n2161), .Z(out[1515]) );
  OR U3552 ( .A(n2392), .B(n2162), .Z(n2163) );
  XNOR U3553 ( .A(n2391), .B(n2163), .Z(out[1516]) );
  OR U3554 ( .A(n2396), .B(n2164), .Z(n2165) );
  XNOR U3555 ( .A(n2395), .B(n2165), .Z(out[1517]) );
  OR U3556 ( .A(n2400), .B(n2166), .Z(n2167) );
  XNOR U3557 ( .A(n2399), .B(n2167), .Z(out[1518]) );
  OR U3558 ( .A(n2404), .B(n2168), .Z(n2169) );
  XNOR U3559 ( .A(n2403), .B(n2169), .Z(out[1519]) );
  XNOR U3560 ( .A(in[688]), .B(n3948), .Z(n2672) );
  XOR U3561 ( .A(in[622]), .B(n3536), .Z(n4303) );
  XNOR U3562 ( .A(in[213]), .B(n3633), .Z(n4301) );
  NAND U3563 ( .A(n4303), .B(n4301), .Z(n2170) );
  XNOR U3564 ( .A(n2672), .B(n2170), .Z(out[151]) );
  OR U3565 ( .A(n2408), .B(n2171), .Z(n2172) );
  XNOR U3566 ( .A(n2407), .B(n2172), .Z(out[1520]) );
  OR U3567 ( .A(n2412), .B(n2173), .Z(n2174) );
  XNOR U3568 ( .A(n2411), .B(n2174), .Z(out[1521]) );
  OR U3569 ( .A(n2416), .B(n2175), .Z(n2176) );
  XNOR U3570 ( .A(n2415), .B(n2176), .Z(out[1522]) );
  OR U3571 ( .A(n2420), .B(n2177), .Z(n2178) );
  XNOR U3572 ( .A(n2419), .B(n2178), .Z(out[1523]) );
  OR U3573 ( .A(n2424), .B(n2179), .Z(n2180) );
  XNOR U3574 ( .A(n2423), .B(n2180), .Z(out[1524]) );
  OR U3575 ( .A(n2428), .B(n2181), .Z(n2182) );
  XNOR U3576 ( .A(n2427), .B(n2182), .Z(out[1525]) );
  OR U3577 ( .A(n2433), .B(n2183), .Z(n2184) );
  XNOR U3578 ( .A(n2432), .B(n2184), .Z(out[1526]) );
  OR U3579 ( .A(n2437), .B(n2185), .Z(n2186) );
  XNOR U3580 ( .A(n2436), .B(n2186), .Z(out[1527]) );
  OR U3581 ( .A(n2441), .B(n2187), .Z(n2188) );
  XNOR U3582 ( .A(n2440), .B(n2188), .Z(out[1528]) );
  OR U3583 ( .A(n2445), .B(n2189), .Z(n2190) );
  XNOR U3584 ( .A(n2444), .B(n2190), .Z(out[1529]) );
  XNOR U3585 ( .A(in[689]), .B(n3950), .Z(n2676) );
  XOR U3586 ( .A(in[623]), .B(n3540), .Z(n4327) );
  XNOR U3587 ( .A(in[214]), .B(n3637), .Z(n4325) );
  NAND U3588 ( .A(n4327), .B(n4325), .Z(n2191) );
  XNOR U3589 ( .A(n2676), .B(n2191), .Z(out[152]) );
  OR U3590 ( .A(n2449), .B(n2192), .Z(n2193) );
  XNOR U3591 ( .A(n2448), .B(n2193), .Z(out[1530]) );
  OR U3592 ( .A(n2453), .B(n2194), .Z(n2195) );
  XNOR U3593 ( .A(n2452), .B(n2195), .Z(out[1531]) );
  OR U3594 ( .A(n2457), .B(n2196), .Z(n2197) );
  XNOR U3595 ( .A(n2456), .B(n2197), .Z(out[1532]) );
  OR U3596 ( .A(n2461), .B(n2198), .Z(n2199) );
  XNOR U3597 ( .A(n2460), .B(n2199), .Z(out[1533]) );
  OR U3598 ( .A(n2465), .B(n2200), .Z(n2201) );
  XNOR U3599 ( .A(n2464), .B(n2201), .Z(out[1534]) );
  OR U3600 ( .A(n2469), .B(n2202), .Z(n2203) );
  XNOR U3601 ( .A(n2468), .B(n2203), .Z(out[1535]) );
  ANDN U3602 ( .B(n2205), .A(n2204), .Z(n2208) );
  XOR U3603 ( .A(n2206), .B(round_const[0]), .Z(n2207) );
  XNOR U3604 ( .A(n2208), .B(n2207), .Z(out[1536]) );
  ANDN U3605 ( .B(n2210), .A(n2209), .Z(n2213) );
  XOR U3606 ( .A(n2211), .B(round_const[1]), .Z(n2212) );
  XNOR U3607 ( .A(n2213), .B(n2212), .Z(out[1537]) );
  ANDN U3608 ( .B(n2215), .A(n2214), .Z(n2216) );
  XNOR U3609 ( .A(n2217), .B(n2216), .Z(out[1538]) );
  ANDN U3610 ( .B(n2219), .A(n2218), .Z(n2222) );
  XOR U3611 ( .A(n2220), .B(round_const_3), .Z(n2221) );
  XNOR U3612 ( .A(n2222), .B(n2221), .Z(out[1539]) );
  XNOR U3613 ( .A(in[690]), .B(n3952), .Z(n2679) );
  XOR U3614 ( .A(in[624]), .B(n3544), .Z(n4359) );
  XNOR U3615 ( .A(in[215]), .B(n3641), .Z(n4357) );
  NAND U3616 ( .A(n4359), .B(n4357), .Z(n2223) );
  XNOR U3617 ( .A(n2679), .B(n2223), .Z(out[153]) );
  ANDN U3618 ( .B(n2225), .A(n2224), .Z(n2226) );
  XNOR U3619 ( .A(n2227), .B(n2226), .Z(out[1540]) );
  ANDN U3620 ( .B(n2229), .A(n2228), .Z(n2230) );
  XNOR U3621 ( .A(n2231), .B(n2230), .Z(out[1541]) );
  ANDN U3622 ( .B(n2233), .A(n2232), .Z(n2234) );
  XNOR U3623 ( .A(n2235), .B(n2234), .Z(out[1542]) );
  ANDN U3624 ( .B(n2237), .A(n2236), .Z(n2240) );
  XOR U3625 ( .A(n2238), .B(round_const_7), .Z(n2239) );
  XNOR U3626 ( .A(n2240), .B(n2239), .Z(out[1543]) );
  ANDN U3627 ( .B(n2242), .A(n2241), .Z(n2243) );
  XNOR U3628 ( .A(n2244), .B(n2243), .Z(out[1544]) );
  ANDN U3629 ( .B(n2246), .A(n2245), .Z(n2247) );
  XNOR U3630 ( .A(n2248), .B(n2247), .Z(out[1545]) );
  ANDN U3631 ( .B(n2250), .A(n2249), .Z(n2251) );
  XNOR U3632 ( .A(n2252), .B(n2251), .Z(out[1546]) );
  ANDN U3633 ( .B(n2254), .A(n2253), .Z(n2255) );
  XNOR U3634 ( .A(n2256), .B(n2255), .Z(out[1547]) );
  ANDN U3635 ( .B(n2258), .A(n2257), .Z(n2259) );
  XNOR U3636 ( .A(n2260), .B(n2259), .Z(out[1548]) );
  ANDN U3637 ( .B(n2262), .A(n2261), .Z(n2263) );
  XNOR U3638 ( .A(n2264), .B(n2263), .Z(out[1549]) );
  XNOR U3639 ( .A(in[691]), .B(n3954), .Z(n2682) );
  XOR U3640 ( .A(in[625]), .B(n3548), .Z(n4407) );
  XNOR U3641 ( .A(in[216]), .B(n3645), .Z(n4405) );
  NAND U3642 ( .A(n4407), .B(n4405), .Z(n2265) );
  XNOR U3643 ( .A(n2682), .B(n2265), .Z(out[154]) );
  ANDN U3644 ( .B(n2267), .A(n2266), .Z(n2268) );
  XNOR U3645 ( .A(n2269), .B(n2268), .Z(out[1550]) );
  ANDN U3646 ( .B(n2271), .A(n2270), .Z(n2274) );
  XOR U3647 ( .A(n2272), .B(round_const_15), .Z(n2273) );
  XNOR U3648 ( .A(n2274), .B(n2273), .Z(out[1551]) );
  ANDN U3649 ( .B(n2276), .A(n2275), .Z(n2277) );
  XNOR U3650 ( .A(n2278), .B(n2277), .Z(out[1552]) );
  ANDN U3651 ( .B(n2280), .A(n2279), .Z(n2281) );
  XNOR U3652 ( .A(n2282), .B(n2281), .Z(out[1553]) );
  ANDN U3653 ( .B(n2284), .A(n2283), .Z(n2285) );
  XNOR U3654 ( .A(n2286), .B(n2285), .Z(out[1554]) );
  ANDN U3655 ( .B(n2288), .A(n2287), .Z(n2289) );
  XNOR U3656 ( .A(n2290), .B(n2289), .Z(out[1555]) );
  ANDN U3657 ( .B(n2292), .A(n2291), .Z(n2293) );
  XNOR U3658 ( .A(n2294), .B(n2293), .Z(out[1556]) );
  ANDN U3659 ( .B(n2296), .A(n2295), .Z(n2297) );
  XNOR U3660 ( .A(n2298), .B(n2297), .Z(out[1557]) );
  ANDN U3661 ( .B(n2300), .A(n2299), .Z(n2301) );
  XNOR U3662 ( .A(n2302), .B(n2301), .Z(out[1558]) );
  ANDN U3663 ( .B(n2304), .A(n2303), .Z(n2305) );
  XNOR U3664 ( .A(n2306), .B(n2305), .Z(out[1559]) );
  XNOR U3665 ( .A(in[692]), .B(n3956), .Z(n2685) );
  XOR U3666 ( .A(in[626]), .B(n3552), .Z(n4451) );
  XNOR U3667 ( .A(in[217]), .B(n3649), .Z(n4449) );
  NAND U3668 ( .A(n4451), .B(n4449), .Z(n2307) );
  XNOR U3669 ( .A(n2685), .B(n2307), .Z(out[155]) );
  ANDN U3670 ( .B(n2309), .A(n2308), .Z(n2310) );
  XNOR U3671 ( .A(n2311), .B(n2310), .Z(out[1560]) );
  ANDN U3672 ( .B(n2313), .A(n2312), .Z(n2314) );
  XNOR U3673 ( .A(n2315), .B(n2314), .Z(out[1561]) );
  ANDN U3674 ( .B(n2317), .A(n2316), .Z(n2318) );
  XNOR U3675 ( .A(n2319), .B(n2318), .Z(out[1562]) );
  ANDN U3676 ( .B(n2321), .A(n2320), .Z(n2322) );
  XNOR U3677 ( .A(n2323), .B(n2322), .Z(out[1563]) );
  ANDN U3678 ( .B(n2325), .A(n2324), .Z(n2326) );
  XNOR U3679 ( .A(n2327), .B(n2326), .Z(out[1564]) );
  ANDN U3680 ( .B(n2329), .A(n2328), .Z(n2330) );
  XNOR U3681 ( .A(n2331), .B(n2330), .Z(out[1565]) );
  ANDN U3682 ( .B(n2333), .A(n2332), .Z(n2334) );
  XNOR U3683 ( .A(n2335), .B(n2334), .Z(out[1566]) );
  ANDN U3684 ( .B(n2337), .A(n2336), .Z(n2340) );
  XOR U3685 ( .A(n2338), .B(round_const_31), .Z(n2339) );
  XNOR U3686 ( .A(n2340), .B(n2339), .Z(out[1567]) );
  ANDN U3687 ( .B(n2342), .A(n2341), .Z(n2343) );
  XNOR U3688 ( .A(n2344), .B(n2343), .Z(out[1568]) );
  ANDN U3689 ( .B(n2346), .A(n2345), .Z(n2347) );
  XNOR U3690 ( .A(n2348), .B(n2347), .Z(out[1569]) );
  XNOR U3691 ( .A(in[693]), .B(n3958), .Z(n2688) );
  XOR U3692 ( .A(in[627]), .B(n3556), .Z(n4495) );
  XNOR U3693 ( .A(in[218]), .B(n3653), .Z(n4492) );
  NAND U3694 ( .A(n4495), .B(n4492), .Z(n2349) );
  XNOR U3695 ( .A(n2688), .B(n2349), .Z(out[156]) );
  ANDN U3696 ( .B(n2351), .A(n2350), .Z(n2352) );
  XNOR U3697 ( .A(n2353), .B(n2352), .Z(out[1570]) );
  ANDN U3698 ( .B(n2355), .A(n2354), .Z(n2356) );
  XNOR U3699 ( .A(n2357), .B(n2356), .Z(out[1571]) );
  ANDN U3700 ( .B(n2359), .A(n2358), .Z(n2360) );
  XNOR U3701 ( .A(n2361), .B(n2360), .Z(out[1572]) );
  ANDN U3702 ( .B(n2363), .A(n2362), .Z(n2364) );
  XNOR U3703 ( .A(n2365), .B(n2364), .Z(out[1573]) );
  ANDN U3704 ( .B(n2367), .A(n2366), .Z(n2368) );
  XNOR U3705 ( .A(n2369), .B(n2368), .Z(out[1574]) );
  ANDN U3706 ( .B(n2371), .A(n2370), .Z(n2372) );
  XNOR U3707 ( .A(n2373), .B(n2372), .Z(out[1575]) );
  ANDN U3708 ( .B(n2375), .A(n2374), .Z(n2376) );
  XNOR U3709 ( .A(n2377), .B(n2376), .Z(out[1576]) );
  ANDN U3710 ( .B(n2379), .A(n2378), .Z(n2380) );
  XNOR U3711 ( .A(n2381), .B(n2380), .Z(out[1577]) );
  ANDN U3712 ( .B(n2383), .A(n2382), .Z(n2384) );
  XNOR U3713 ( .A(n2385), .B(n2384), .Z(out[1578]) );
  ANDN U3714 ( .B(n2387), .A(n2386), .Z(n2388) );
  XNOR U3715 ( .A(n2389), .B(n2388), .Z(out[1579]) );
  XNOR U3716 ( .A(in[694]), .B(n3960), .Z(n2690) );
  XOR U3717 ( .A(in[628]), .B(n3560), .Z(n4539) );
  XNOR U3718 ( .A(in[219]), .B(n3657), .Z(n4536) );
  NAND U3719 ( .A(n4539), .B(n4536), .Z(n2390) );
  XNOR U3720 ( .A(n2690), .B(n2390), .Z(out[157]) );
  ANDN U3721 ( .B(n2392), .A(n2391), .Z(n2393) );
  XNOR U3722 ( .A(n2394), .B(n2393), .Z(out[1580]) );
  ANDN U3723 ( .B(n2396), .A(n2395), .Z(n2397) );
  XNOR U3724 ( .A(n2398), .B(n2397), .Z(out[1581]) );
  ANDN U3725 ( .B(n2400), .A(n2399), .Z(n2401) );
  XNOR U3726 ( .A(n2402), .B(n2401), .Z(out[1582]) );
  ANDN U3727 ( .B(n2404), .A(n2403), .Z(n2405) );
  XNOR U3728 ( .A(n2406), .B(n2405), .Z(out[1583]) );
  ANDN U3729 ( .B(n2408), .A(n2407), .Z(n2409) );
  XNOR U3730 ( .A(n2410), .B(n2409), .Z(out[1584]) );
  ANDN U3731 ( .B(n2412), .A(n2411), .Z(n2413) );
  XNOR U3732 ( .A(n2414), .B(n2413), .Z(out[1585]) );
  ANDN U3733 ( .B(n2416), .A(n2415), .Z(n2417) );
  XNOR U3734 ( .A(n2418), .B(n2417), .Z(out[1586]) );
  ANDN U3735 ( .B(n2420), .A(n2419), .Z(n2421) );
  XNOR U3736 ( .A(n2422), .B(n2421), .Z(out[1587]) );
  ANDN U3737 ( .B(n2424), .A(n2423), .Z(n2425) );
  XNOR U3738 ( .A(n2426), .B(n2425), .Z(out[1588]) );
  ANDN U3739 ( .B(n2428), .A(n2427), .Z(n2429) );
  XNOR U3740 ( .A(n2430), .B(n2429), .Z(out[1589]) );
  XNOR U3741 ( .A(in[695]), .B(n3962), .Z(n2692) );
  XOR U3742 ( .A(in[629]), .B(n3564), .Z(n4583) );
  XNOR U3743 ( .A(in[220]), .B(n3661), .Z(n4580) );
  NAND U3744 ( .A(n4583), .B(n4580), .Z(n2431) );
  XNOR U3745 ( .A(n2692), .B(n2431), .Z(out[158]) );
  ANDN U3746 ( .B(n2433), .A(n2432), .Z(n2434) );
  XNOR U3747 ( .A(n2435), .B(n2434), .Z(out[1590]) );
  ANDN U3748 ( .B(n2437), .A(n2436), .Z(n2438) );
  XNOR U3749 ( .A(n2439), .B(n2438), .Z(out[1591]) );
  ANDN U3750 ( .B(n2441), .A(n2440), .Z(n2442) );
  XNOR U3751 ( .A(n2443), .B(n2442), .Z(out[1592]) );
  ANDN U3752 ( .B(n2445), .A(n2444), .Z(n2446) );
  XNOR U3753 ( .A(n2447), .B(n2446), .Z(out[1593]) );
  ANDN U3754 ( .B(n2449), .A(n2448), .Z(n2450) );
  XNOR U3755 ( .A(n2451), .B(n2450), .Z(out[1594]) );
  ANDN U3756 ( .B(n2453), .A(n2452), .Z(n2454) );
  XNOR U3757 ( .A(n2455), .B(n2454), .Z(out[1595]) );
  ANDN U3758 ( .B(n2457), .A(n2456), .Z(n2458) );
  XNOR U3759 ( .A(n2459), .B(n2458), .Z(out[1596]) );
  ANDN U3760 ( .B(n2461), .A(n2460), .Z(n2462) );
  XNOR U3761 ( .A(n2463), .B(n2462), .Z(out[1597]) );
  ANDN U3762 ( .B(n2465), .A(n2464), .Z(n2466) );
  XNOR U3763 ( .A(n2467), .B(n2466), .Z(out[1598]) );
  ANDN U3764 ( .B(n2469), .A(n2468), .Z(n2472) );
  XOR U3765 ( .A(n2470), .B(round_const_7), .Z(n2471) );
  XNOR U3766 ( .A(n2472), .B(n2471), .Z(out[1599]) );
  XNOR U3767 ( .A(in[696]), .B(n3818), .Z(n2694) );
  XOR U3768 ( .A(in[630]), .B(n3568), .Z(n4627) );
  XNOR U3769 ( .A(in[221]), .B(n3669), .Z(n4624) );
  NAND U3770 ( .A(n4627), .B(n4624), .Z(n2473) );
  XNOR U3771 ( .A(n2694), .B(n2473), .Z(out[159]) );
  XNOR U3772 ( .A(in[1425]), .B(n3638), .Z(n4072) );
  XOR U3773 ( .A(in[1048]), .B(n4135), .Z(n2648) );
  NAND U3774 ( .A(n4072), .B(n2648), .Z(n2474) );
  XNOR U3775 ( .A(n4073), .B(n2474), .Z(out[15]) );
  XNOR U3776 ( .A(in[697]), .B(n3820), .Z(n2696) );
  XOR U3777 ( .A(in[631]), .B(n3572), .Z(n4671) );
  XNOR U3778 ( .A(in[222]), .B(n3673), .Z(n4668) );
  NAND U3779 ( .A(n4671), .B(n4668), .Z(n2475) );
  XNOR U3780 ( .A(n2696), .B(n2475), .Z(out[160]) );
  XNOR U3781 ( .A(in[698]), .B(n3822), .Z(n2698) );
  XOR U3782 ( .A(in[632]), .B(n3580), .Z(n4715) );
  XNOR U3783 ( .A(in[223]), .B(n3677), .Z(n4712) );
  NAND U3784 ( .A(n4715), .B(n4712), .Z(n2476) );
  XNOR U3785 ( .A(n2698), .B(n2476), .Z(out[161]) );
  XNOR U3786 ( .A(in[699]), .B(n3824), .Z(n2702) );
  XOR U3787 ( .A(in[633]), .B(n3584), .Z(n4759) );
  XNOR U3788 ( .A(in[224]), .B(n3681), .Z(n4756) );
  NAND U3789 ( .A(n4759), .B(n4756), .Z(n2477) );
  XNOR U3790 ( .A(n2702), .B(n2477), .Z(out[162]) );
  XNOR U3791 ( .A(in[700]), .B(n3826), .Z(n2704) );
  XOR U3792 ( .A(in[634]), .B(n3588), .Z(n4803) );
  XNOR U3793 ( .A(in[225]), .B(n3685), .Z(n4800) );
  NAND U3794 ( .A(n4803), .B(n4800), .Z(n2478) );
  XNOR U3795 ( .A(n2704), .B(n2478), .Z(out[163]) );
  XOR U3796 ( .A(in[701]), .B(n3828), .Z(n2706) );
  NOR U3797 ( .A(n2550), .B(n2831), .Z(n2479) );
  XNOR U3798 ( .A(n2706), .B(n2479), .Z(out[164]) );
  XOR U3799 ( .A(in[702]), .B(n3834), .Z(n2708) );
  NOR U3800 ( .A(n2552), .B(n2845), .Z(n2480) );
  XNOR U3801 ( .A(n2708), .B(n2480), .Z(out[165]) );
  XOR U3802 ( .A(in[703]), .B(n3836), .Z(n2710) );
  NOR U3803 ( .A(n2555), .B(n2859), .Z(n2481) );
  XNOR U3804 ( .A(n2710), .B(n2481), .Z(out[166]) );
  XOR U3805 ( .A(in[640]), .B(n3838), .Z(n2712) );
  NOR U3806 ( .A(n2557), .B(n2873), .Z(n2482) );
  XNOR U3807 ( .A(n2712), .B(n2482), .Z(out[167]) );
  XOR U3808 ( .A(in[641]), .B(n3840), .Z(n2714) );
  NOR U3809 ( .A(n2559), .B(n2889), .Z(n2483) );
  XNOR U3810 ( .A(n2714), .B(n2483), .Z(out[168]) );
  XOR U3811 ( .A(in[642]), .B(n3842), .Z(n2716) );
  NOR U3812 ( .A(n2561), .B(n2903), .Z(n2484) );
  XNOR U3813 ( .A(n2716), .B(n2484), .Z(out[169]) );
  XNOR U3814 ( .A(in[1426]), .B(n3642), .Z(n4110) );
  XOR U3815 ( .A(in[1049]), .B(n4138), .Z(n2651) );
  NAND U3816 ( .A(n4110), .B(n2651), .Z(n2485) );
  XNOR U3817 ( .A(n4111), .B(n2485), .Z(out[16]) );
  XOR U3818 ( .A(in[643]), .B(n3844), .Z(n2718) );
  NOR U3819 ( .A(n2563), .B(n2917), .Z(n2486) );
  XNOR U3820 ( .A(n2718), .B(n2486), .Z(out[170]) );
  XOR U3821 ( .A(in[644]), .B(n3846), .Z(n2720) );
  NOR U3822 ( .A(n2565), .B(n2931), .Z(n2487) );
  XNOR U3823 ( .A(n2720), .B(n2487), .Z(out[171]) );
  XOR U3824 ( .A(in[645]), .B(n3848), .Z(n2726) );
  NOR U3825 ( .A(n2567), .B(n2947), .Z(n2488) );
  XNOR U3826 ( .A(n2726), .B(n2488), .Z(out[172]) );
  XOR U3827 ( .A(in[646]), .B(n3850), .Z(n2728) );
  NOR U3828 ( .A(n2569), .B(n2971), .Z(n2489) );
  XNOR U3829 ( .A(n2728), .B(n2489), .Z(out[173]) );
  XOR U3830 ( .A(in[647]), .B(n3852), .Z(n2730) );
  NOR U3831 ( .A(n2571), .B(n2995), .Z(n2490) );
  XNOR U3832 ( .A(n2730), .B(n2490), .Z(out[174]) );
  XOR U3833 ( .A(in[648]), .B(n3856), .Z(n2732) );
  NOR U3834 ( .A(n2573), .B(n3019), .Z(n2491) );
  XNOR U3835 ( .A(n2732), .B(n2491), .Z(out[175]) );
  XOR U3836 ( .A(in[649]), .B(n3858), .Z(n2734) );
  NOR U3837 ( .A(n2576), .B(n3043), .Z(n2492) );
  XNOR U3838 ( .A(n2734), .B(n2492), .Z(out[176]) );
  XOR U3839 ( .A(in[650]), .B(n3860), .Z(n2736) );
  NOR U3840 ( .A(n2578), .B(n3067), .Z(n2493) );
  XNOR U3841 ( .A(n2736), .B(n2493), .Z(out[177]) );
  XOR U3842 ( .A(in[651]), .B(n3862), .Z(n2738) );
  NOR U3843 ( .A(n2580), .B(n3093), .Z(n2494) );
  XNOR U3844 ( .A(n2738), .B(n2494), .Z(out[178]) );
  XOR U3845 ( .A(in[652]), .B(n3864), .Z(n2740) );
  NOR U3846 ( .A(n2582), .B(n3117), .Z(n2495) );
  XNOR U3847 ( .A(n2740), .B(n2495), .Z(out[179]) );
  XNOR U3848 ( .A(in[1427]), .B(n3646), .Z(n4144) );
  XOR U3849 ( .A(in[1050]), .B(n4141), .Z(n2654) );
  NAND U3850 ( .A(n4144), .B(n2654), .Z(n2496) );
  XNOR U3851 ( .A(n4145), .B(n2496), .Z(out[17]) );
  XOR U3852 ( .A(in[653]), .B(n3866), .Z(n2742) );
  NOR U3853 ( .A(n2584), .B(n3141), .Z(n2497) );
  XNOR U3854 ( .A(n2742), .B(n2497), .Z(out[180]) );
  XOR U3855 ( .A(in[654]), .B(n3868), .Z(n2744) );
  NOR U3856 ( .A(n2586), .B(n3165), .Z(n2498) );
  XNOR U3857 ( .A(n2744), .B(n2498), .Z(out[181]) );
  XOR U3858 ( .A(in[655]), .B(n3870), .Z(n2748) );
  NOR U3859 ( .A(n2588), .B(n3189), .Z(n2499) );
  XNOR U3860 ( .A(n2748), .B(n2499), .Z(out[182]) );
  XOR U3861 ( .A(in[656]), .B(n3872), .Z(n2750) );
  NOR U3862 ( .A(n2590), .B(n3213), .Z(n2500) );
  XNOR U3863 ( .A(n2750), .B(n2500), .Z(out[183]) );
  XOR U3864 ( .A(in[657]), .B(n3874), .Z(n2752) );
  NOR U3865 ( .A(n2592), .B(n3237), .Z(n2501) );
  XNOR U3866 ( .A(n2752), .B(n2501), .Z(out[184]) );
  XOR U3867 ( .A(in[658]), .B(n3878), .Z(n2754) );
  NOR U3868 ( .A(n2594), .B(n3269), .Z(n2502) );
  XNOR U3869 ( .A(n2754), .B(n2502), .Z(out[185]) );
  XOR U3870 ( .A(in[659]), .B(n3880), .Z(n2756) );
  NOR U3871 ( .A(n2597), .B(n3313), .Z(n2503) );
  XNOR U3872 ( .A(n2756), .B(n2503), .Z(out[186]) );
  XOR U3873 ( .A(in[660]), .B(n3882), .Z(n2758) );
  NOR U3874 ( .A(n2599), .B(n3357), .Z(n2504) );
  XNOR U3875 ( .A(n2758), .B(n2504), .Z(out[187]) );
  XOR U3876 ( .A(in[661]), .B(n3884), .Z(n2760) );
  NOR U3877 ( .A(n2601), .B(n3403), .Z(n2505) );
  XNOR U3878 ( .A(n2760), .B(n2505), .Z(out[188]) );
  XOR U3879 ( .A(in[662]), .B(n3886), .Z(n2762) );
  NOR U3880 ( .A(n2603), .B(n3447), .Z(n2506) );
  XNOR U3881 ( .A(n2762), .B(n2506), .Z(out[189]) );
  XNOR U3882 ( .A(in[1428]), .B(n3650), .Z(n4178) );
  XOR U3883 ( .A(in[1051]), .B(n4148), .Z(n2657) );
  NAND U3884 ( .A(n4178), .B(n2657), .Z(n2507) );
  XNOR U3885 ( .A(n4179), .B(n2507), .Z(out[18]) );
  XOR U3886 ( .A(in[663]), .B(n3888), .Z(n2764) );
  NOR U3887 ( .A(n2605), .B(n3491), .Z(n2508) );
  XNOR U3888 ( .A(n2764), .B(n2508), .Z(out[190]) );
  XOR U3889 ( .A(in[664]), .B(n3890), .Z(n2766) );
  NOR U3890 ( .A(n2607), .B(n3535), .Z(n2509) );
  XNOR U3891 ( .A(n2766), .B(n2509), .Z(out[191]) );
  OR U3892 ( .A(n2610), .B(n3579), .Z(n2510) );
  XNOR U3893 ( .A(n2609), .B(n2510), .Z(out[192]) );
  XOR U3894 ( .A(in[1034]), .B(n4089), .Z(n2613) );
  NOR U3895 ( .A(n2612), .B(n3623), .Z(n2511) );
  XNOR U3896 ( .A(n2613), .B(n2511), .Z(out[193]) );
  XOR U3897 ( .A(in[1035]), .B(n4092), .Z(n2724) );
  NOR U3898 ( .A(n2615), .B(n3667), .Z(n2512) );
  XNOR U3899 ( .A(n2724), .B(n2512), .Z(out[194]) );
  XNOR U3900 ( .A(n4095), .B(in[1036]), .Z(n2874) );
  NOR U3901 ( .A(n2617), .B(n3711), .Z(n2513) );
  XNOR U3902 ( .A(n2874), .B(n2513), .Z(out[195]) );
  XNOR U3903 ( .A(n4098), .B(in[1037]), .Z(n3068) );
  NOR U3904 ( .A(n2620), .B(n3755), .Z(n2514) );
  XNOR U3905 ( .A(n3068), .B(n2514), .Z(out[196]) );
  XNOR U3906 ( .A(n4101), .B(in[1038]), .Z(n3358) );
  NOR U3907 ( .A(n2622), .B(n3799), .Z(n2515) );
  XNOR U3908 ( .A(n3358), .B(n2515), .Z(out[197]) );
  XNOR U3909 ( .A(n4104), .B(in[1039]), .Z(n3800) );
  NOR U3910 ( .A(n2624), .B(n3833), .Z(n2516) );
  XNOR U3911 ( .A(n3800), .B(n2516), .Z(out[198]) );
  XNOR U3912 ( .A(n4107), .B(in[1040]), .Z(n4076) );
  NOR U3913 ( .A(n2626), .B(n3855), .Z(n2517) );
  XNOR U3914 ( .A(n4076), .B(n2517), .Z(out[199]) );
  XNOR U3915 ( .A(in[1429]), .B(n3654), .Z(n4204) );
  XOR U3916 ( .A(in[1052]), .B(n4151), .Z(n2660) );
  NAND U3917 ( .A(n4204), .B(n2660), .Z(n2518) );
  XNOR U3918 ( .A(n4205), .B(n2518), .Z(out[19]) );
  XNOR U3919 ( .A(n3574), .B(in[1411]), .Z(n3620) );
  NANDN U3920 ( .A(n2613), .B(n3620), .Z(n2519) );
  XNOR U3921 ( .A(n3621), .B(n2519), .Z(out[1]) );
  XNOR U3922 ( .A(n4114), .B(in[1041]), .Z(n4360) );
  NOR U3923 ( .A(n2628), .B(n3877), .Z(n2520) );
  XNOR U3924 ( .A(n4360), .B(n2520), .Z(out[200]) );
  XNOR U3925 ( .A(n4117), .B(in[1042]), .Z(n4804) );
  NOR U3926 ( .A(n2630), .B(n3899), .Z(n2521) );
  XNOR U3927 ( .A(n4804), .B(n2521), .Z(out[201]) );
  OR U3928 ( .A(n2633), .B(n3923), .Z(n2522) );
  XNOR U3929 ( .A(n2632), .B(n2522), .Z(out[202]) );
  OR U3930 ( .A(n2636), .B(n3947), .Z(n2523) );
  XNOR U3931 ( .A(n2635), .B(n2523), .Z(out[203]) );
  OR U3932 ( .A(n2639), .B(n3973), .Z(n2524) );
  XNOR U3933 ( .A(n2638), .B(n2524), .Z(out[204]) );
  OR U3934 ( .A(n2642), .B(n4007), .Z(n2525) );
  XNOR U3935 ( .A(n2641), .B(n2525), .Z(out[205]) );
  OR U3936 ( .A(n2646), .B(n4041), .Z(n2526) );
  XNOR U3937 ( .A(n2645), .B(n2526), .Z(out[206]) );
  OR U3938 ( .A(n2649), .B(n4075), .Z(n2527) );
  XNOR U3939 ( .A(n2648), .B(n2527), .Z(out[207]) );
  OR U3940 ( .A(n2652), .B(n4113), .Z(n2528) );
  XNOR U3941 ( .A(n2651), .B(n2528), .Z(out[208]) );
  OR U3942 ( .A(n2655), .B(n4147), .Z(n2529) );
  XNOR U3943 ( .A(n2654), .B(n2529), .Z(out[209]) );
  XNOR U3944 ( .A(in[1430]), .B(n3658), .Z(n4228) );
  XOR U3945 ( .A(in[1053]), .B(n4154), .Z(n2663) );
  NAND U3946 ( .A(n4228), .B(n2663), .Z(n2530) );
  XNOR U3947 ( .A(n4229), .B(n2530), .Z(out[20]) );
  OR U3948 ( .A(n2658), .B(n4181), .Z(n2531) );
  XNOR U3949 ( .A(n2657), .B(n2531), .Z(out[210]) );
  OR U3950 ( .A(n2661), .B(n4207), .Z(n2532) );
  XNOR U3951 ( .A(n2660), .B(n2532), .Z(out[211]) );
  OR U3952 ( .A(n2664), .B(n4231), .Z(n2533) );
  XNOR U3953 ( .A(n2663), .B(n2533), .Z(out[212]) );
  XNOR U3954 ( .A(in[1054]), .B(n4157), .Z(n2667) );
  NOR U3955 ( .A(n2666), .B(n4255), .Z(n2534) );
  XNOR U3956 ( .A(n2667), .B(n2534), .Z(out[213]) );
  XNOR U3957 ( .A(in[1055]), .B(n4160), .Z(n2670) );
  NOR U3958 ( .A(n2669), .B(n4279), .Z(n2535) );
  XNOR U3959 ( .A(n2670), .B(n2535), .Z(out[214]) );
  XNOR U3960 ( .A(in[1056]), .B(n4163), .Z(n2673) );
  NOR U3961 ( .A(n2672), .B(n4303), .Z(n2536) );
  XNOR U3962 ( .A(n2673), .B(n2536), .Z(out[215]) );
  XNOR U3963 ( .A(in[1057]), .B(n4166), .Z(n2677) );
  NOR U3964 ( .A(n2676), .B(n4327), .Z(n2537) );
  XNOR U3965 ( .A(n2677), .B(n2537), .Z(out[216]) );
  XNOR U3966 ( .A(in[1058]), .B(n4169), .Z(n2680) );
  NOR U3967 ( .A(n2679), .B(n4359), .Z(n2538) );
  XNOR U3968 ( .A(n2680), .B(n2538), .Z(out[217]) );
  XNOR U3969 ( .A(in[1059]), .B(n4172), .Z(n2683) );
  NOR U3970 ( .A(n2682), .B(n4407), .Z(n2539) );
  XNOR U3971 ( .A(n2683), .B(n2539), .Z(out[218]) );
  XOR U3972 ( .A(in[1060]), .B(n4175), .Z(n2686) );
  NOR U3973 ( .A(n2685), .B(n4451), .Z(n2540) );
  XNOR U3974 ( .A(n2686), .B(n2540), .Z(out[219]) );
  XNOR U3975 ( .A(in[1431]), .B(n3662), .Z(n4252) );
  NANDN U3976 ( .A(n2667), .B(n4252), .Z(n2541) );
  XNOR U3977 ( .A(n4253), .B(n2541), .Z(out[21]) );
  XOR U3978 ( .A(in[1061]), .B(n4182), .Z(n2700) );
  NOR U3979 ( .A(n2688), .B(n4495), .Z(n2542) );
  XNOR U3980 ( .A(n2700), .B(n2542), .Z(out[220]) );
  XOR U3981 ( .A(in[1062]), .B(n4185), .Z(n2722) );
  NOR U3982 ( .A(n2690), .B(n4539), .Z(n2543) );
  XNOR U3983 ( .A(n2722), .B(n2543), .Z(out[221]) );
  XOR U3984 ( .A(in[1063]), .B(n3964), .Z(n2746) );
  NOR U3985 ( .A(n2692), .B(n4583), .Z(n2544) );
  XNOR U3986 ( .A(n2746), .B(n2544), .Z(out[222]) );
  XOR U3987 ( .A(in[1064]), .B(n3967), .Z(n2768) );
  NOR U3988 ( .A(n2694), .B(n4627), .Z(n2545) );
  XNOR U3989 ( .A(n2768), .B(n2545), .Z(out[223]) );
  XOR U3990 ( .A(in[1065]), .B(n3974), .Z(n2780) );
  NOR U3991 ( .A(n2696), .B(n4671), .Z(n2546) );
  XNOR U3992 ( .A(n2780), .B(n2546), .Z(out[224]) );
  XOR U3993 ( .A(in[1066]), .B(n3977), .Z(n2792) );
  NOR U3994 ( .A(n2698), .B(n4715), .Z(n2547) );
  XNOR U3995 ( .A(n2792), .B(n2547), .Z(out[225]) );
  XOR U3996 ( .A(in[1067]), .B(n3980), .Z(n2804) );
  NOR U3997 ( .A(n2702), .B(n4759), .Z(n2548) );
  XNOR U3998 ( .A(n2804), .B(n2548), .Z(out[226]) );
  XOR U3999 ( .A(in[1068]), .B(n3983), .Z(n2816) );
  NOR U4000 ( .A(n2704), .B(n4803), .Z(n2549) );
  XNOR U4001 ( .A(n2816), .B(n2549), .Z(out[227]) );
  XNOR U4002 ( .A(in[1069]), .B(n3986), .Z(n2829) );
  NAND U4003 ( .A(n2706), .B(n2550), .Z(n2551) );
  XNOR U4004 ( .A(n2829), .B(n2551), .Z(out[228]) );
  XNOR U4005 ( .A(in[1070]), .B(n3989), .Z(n2843) );
  NAND U4006 ( .A(n2708), .B(n2552), .Z(n2553) );
  XNOR U4007 ( .A(n2843), .B(n2553), .Z(out[229]) );
  XNOR U4008 ( .A(in[1432]), .B(n3670), .Z(n4276) );
  NANDN U4009 ( .A(n2670), .B(n4276), .Z(n2554) );
  XNOR U4010 ( .A(n4277), .B(n2554), .Z(out[22]) );
  XNOR U4011 ( .A(in[1071]), .B(n3992), .Z(n2857) );
  NAND U4012 ( .A(n2710), .B(n2555), .Z(n2556) );
  XNOR U4013 ( .A(n2857), .B(n2556), .Z(out[230]) );
  XNOR U4014 ( .A(in[1072]), .B(n3995), .Z(n2871) );
  NAND U4015 ( .A(n2712), .B(n2557), .Z(n2558) );
  XNOR U4016 ( .A(n2871), .B(n2558), .Z(out[231]) );
  XNOR U4017 ( .A(in[1073]), .B(n3998), .Z(n2887) );
  NAND U4018 ( .A(n2714), .B(n2559), .Z(n2560) );
  XNOR U4019 ( .A(n2887), .B(n2560), .Z(out[232]) );
  XNOR U4020 ( .A(in[1074]), .B(n4001), .Z(n2901) );
  NAND U4021 ( .A(n2716), .B(n2561), .Z(n2562) );
  XNOR U4022 ( .A(n2901), .B(n2562), .Z(out[233]) );
  XNOR U4023 ( .A(in[1075]), .B(n4008), .Z(n2915) );
  NAND U4024 ( .A(n2718), .B(n2563), .Z(n2564) );
  XNOR U4025 ( .A(n2915), .B(n2564), .Z(out[234]) );
  XNOR U4026 ( .A(in[1076]), .B(n4011), .Z(n2929) );
  NAND U4027 ( .A(n2720), .B(n2565), .Z(n2566) );
  XNOR U4028 ( .A(n2929), .B(n2566), .Z(out[235]) );
  XNOR U4029 ( .A(in[1077]), .B(n4014), .Z(n2945) );
  NAND U4030 ( .A(n2726), .B(n2567), .Z(n2568) );
  XNOR U4031 ( .A(n2945), .B(n2568), .Z(out[236]) );
  XNOR U4032 ( .A(in[1078]), .B(n4017), .Z(n2969) );
  NAND U4033 ( .A(n2728), .B(n2569), .Z(n2570) );
  XNOR U4034 ( .A(n2969), .B(n2570), .Z(out[237]) );
  XNOR U4035 ( .A(in[1079]), .B(n4020), .Z(n2993) );
  NAND U4036 ( .A(n2730), .B(n2571), .Z(n2572) );
  XNOR U4037 ( .A(n2993), .B(n2572), .Z(out[238]) );
  XNOR U4038 ( .A(in[1080]), .B(n4023), .Z(n3017) );
  NAND U4039 ( .A(n2732), .B(n2573), .Z(n2574) );
  XNOR U4040 ( .A(n3017), .B(n2574), .Z(out[239]) );
  XNOR U4041 ( .A(in[1433]), .B(n3674), .Z(n4300) );
  NANDN U4042 ( .A(n2673), .B(n4300), .Z(n2575) );
  XNOR U4043 ( .A(n4301), .B(n2575), .Z(out[23]) );
  XNOR U4044 ( .A(in[1081]), .B(n4026), .Z(n3041) );
  NAND U4045 ( .A(n2734), .B(n2576), .Z(n2577) );
  XNOR U4046 ( .A(n3041), .B(n2577), .Z(out[240]) );
  XNOR U4047 ( .A(in[1082]), .B(n4029), .Z(n3065) );
  NAND U4048 ( .A(n2736), .B(n2578), .Z(n2579) );
  XNOR U4049 ( .A(n3065), .B(n2579), .Z(out[241]) );
  XNOR U4050 ( .A(in[1083]), .B(n4032), .Z(n3091) );
  NAND U4051 ( .A(n2738), .B(n2580), .Z(n2581) );
  XNOR U4052 ( .A(n3091), .B(n2581), .Z(out[242]) );
  XNOR U4053 ( .A(in[1084]), .B(n4035), .Z(n3115) );
  NAND U4054 ( .A(n2740), .B(n2582), .Z(n2583) );
  XNOR U4055 ( .A(n3115), .B(n2583), .Z(out[243]) );
  XNOR U4056 ( .A(in[1085]), .B(n4042), .Z(n3139) );
  NAND U4057 ( .A(n2742), .B(n2584), .Z(n2585) );
  XNOR U4058 ( .A(n3139), .B(n2585), .Z(out[244]) );
  XNOR U4059 ( .A(in[1086]), .B(n4045), .Z(n3163) );
  NAND U4060 ( .A(n2744), .B(n2586), .Z(n2587) );
  XNOR U4061 ( .A(n3163), .B(n2587), .Z(out[245]) );
  XNOR U4062 ( .A(in[1087]), .B(n4048), .Z(n3187) );
  NAND U4063 ( .A(n2748), .B(n2588), .Z(n2589) );
  XNOR U4064 ( .A(n3187), .B(n2589), .Z(out[246]) );
  XNOR U4065 ( .A(in[1024]), .B(n4051), .Z(n3211) );
  NAND U4066 ( .A(n2750), .B(n2590), .Z(n2591) );
  XNOR U4067 ( .A(n3211), .B(n2591), .Z(out[247]) );
  XNOR U4068 ( .A(in[1025]), .B(n4054), .Z(n3235) );
  NAND U4069 ( .A(n2752), .B(n2592), .Z(n2593) );
  XNOR U4070 ( .A(n3235), .B(n2593), .Z(out[248]) );
  XNOR U4071 ( .A(in[1026]), .B(n4057), .Z(n3267) );
  NAND U4072 ( .A(n2754), .B(n2594), .Z(n2595) );
  XNOR U4073 ( .A(n3267), .B(n2595), .Z(out[249]) );
  XNOR U4074 ( .A(in[1434]), .B(n3678), .Z(n4324) );
  NANDN U4075 ( .A(n2677), .B(n4324), .Z(n2596) );
  XNOR U4076 ( .A(n4325), .B(n2596), .Z(out[24]) );
  XNOR U4077 ( .A(in[1027]), .B(n4060), .Z(n3311) );
  NAND U4078 ( .A(n2756), .B(n2597), .Z(n2598) );
  XNOR U4079 ( .A(n3311), .B(n2598), .Z(out[250]) );
  XNOR U4080 ( .A(in[1028]), .B(n4063), .Z(n3355) );
  NAND U4081 ( .A(n2758), .B(n2599), .Z(n2600) );
  XNOR U4082 ( .A(n3355), .B(n2600), .Z(out[251]) );
  XNOR U4083 ( .A(in[1029]), .B(n4066), .Z(n3401) );
  NAND U4084 ( .A(n2760), .B(n2601), .Z(n2602) );
  XNOR U4085 ( .A(n3401), .B(n2602), .Z(out[252]) );
  XNOR U4086 ( .A(in[1030]), .B(n4069), .Z(n3445) );
  NAND U4087 ( .A(n2762), .B(n2603), .Z(n2604) );
  XNOR U4088 ( .A(n3445), .B(n2604), .Z(out[253]) );
  XNOR U4089 ( .A(in[1031]), .B(n4080), .Z(n3489) );
  NAND U4090 ( .A(n2764), .B(n2605), .Z(n2606) );
  XNOR U4091 ( .A(n3489), .B(n2606), .Z(out[254]) );
  XNOR U4092 ( .A(in[1032]), .B(n4083), .Z(n3533) );
  NAND U4093 ( .A(n2766), .B(n2607), .Z(n2608) );
  XNOR U4094 ( .A(n3533), .B(n2608), .Z(out[255]) );
  ANDN U4095 ( .B(n2610), .A(n2609), .Z(n2611) );
  XNOR U4096 ( .A(n3576), .B(n2611), .Z(out[256]) );
  AND U4097 ( .A(n2613), .B(n2612), .Z(n2614) );
  XNOR U4098 ( .A(n3620), .B(n2614), .Z(out[257]) );
  XOR U4099 ( .A(n3582), .B(in[1412]), .Z(n3665) );
  NAND U4100 ( .A(n2724), .B(n2615), .Z(n2616) );
  XNOR U4101 ( .A(n3665), .B(n2616), .Z(out[258]) );
  XOR U4102 ( .A(n3586), .B(in[1413]), .Z(n3709) );
  NAND U4103 ( .A(n2874), .B(n2617), .Z(n2618) );
  XNOR U4104 ( .A(n3709), .B(n2618), .Z(out[259]) );
  XNOR U4105 ( .A(in[1435]), .B(n3682), .Z(n4356) );
  NANDN U4106 ( .A(n2680), .B(n4356), .Z(n2619) );
  XNOR U4107 ( .A(n4357), .B(n2619), .Z(out[25]) );
  XOR U4108 ( .A(n3590), .B(in[1414]), .Z(n3753) );
  NAND U4109 ( .A(n3068), .B(n2620), .Z(n2621) );
  XNOR U4110 ( .A(n3753), .B(n2621), .Z(out[260]) );
  XOR U4111 ( .A(n3594), .B(in[1415]), .Z(n3797) );
  NAND U4112 ( .A(n3358), .B(n2622), .Z(n2623) );
  XNOR U4113 ( .A(n3797), .B(n2623), .Z(out[261]) );
  XOR U4114 ( .A(n3598), .B(in[1416]), .Z(n3831) );
  NAND U4115 ( .A(n3800), .B(n2624), .Z(n2625) );
  XNOR U4116 ( .A(n3831), .B(n2625), .Z(out[262]) );
  XOR U4117 ( .A(in[1417]), .B(n3602), .Z(n4077) );
  NAND U4118 ( .A(n4076), .B(n2626), .Z(n2627) );
  XNOR U4119 ( .A(n4077), .B(n2627), .Z(out[263]) );
  XOR U4120 ( .A(n3606), .B(in[1418]), .Z(n4361) );
  NAND U4121 ( .A(n4360), .B(n2628), .Z(n2629) );
  XNOR U4122 ( .A(n4361), .B(n2629), .Z(out[264]) );
  XOR U4123 ( .A(n3610), .B(in[1419]), .Z(n4805) );
  NAND U4124 ( .A(n4804), .B(n2630), .Z(n2631) );
  XNOR U4125 ( .A(n4805), .B(n2631), .Z(out[265]) );
  ANDN U4126 ( .B(n2633), .A(n2632), .Z(n2634) );
  XNOR U4127 ( .A(n3920), .B(n2634), .Z(out[266]) );
  ANDN U4128 ( .B(n2636), .A(n2635), .Z(n2637) );
  XNOR U4129 ( .A(n3944), .B(n2637), .Z(out[267]) );
  ANDN U4130 ( .B(n2639), .A(n2638), .Z(n2640) );
  XNOR U4131 ( .A(n3970), .B(n2640), .Z(out[268]) );
  ANDN U4132 ( .B(n2642), .A(n2641), .Z(n2643) );
  XNOR U4133 ( .A(n4004), .B(n2643), .Z(out[269]) );
  XNOR U4134 ( .A(in[1436]), .B(n3686), .Z(n4404) );
  NANDN U4135 ( .A(n2683), .B(n4404), .Z(n2644) );
  XNOR U4136 ( .A(n4405), .B(n2644), .Z(out[26]) );
  ANDN U4137 ( .B(n2646), .A(n2645), .Z(n2647) );
  XNOR U4138 ( .A(n4038), .B(n2647), .Z(out[270]) );
  ANDN U4139 ( .B(n2649), .A(n2648), .Z(n2650) );
  XNOR U4140 ( .A(n4072), .B(n2650), .Z(out[271]) );
  ANDN U4141 ( .B(n2652), .A(n2651), .Z(n2653) );
  XNOR U4142 ( .A(n4110), .B(n2653), .Z(out[272]) );
  ANDN U4143 ( .B(n2655), .A(n2654), .Z(n2656) );
  XNOR U4144 ( .A(n4144), .B(n2656), .Z(out[273]) );
  ANDN U4145 ( .B(n2658), .A(n2657), .Z(n2659) );
  XNOR U4146 ( .A(n4178), .B(n2659), .Z(out[274]) );
  ANDN U4147 ( .B(n2661), .A(n2660), .Z(n2662) );
  XNOR U4148 ( .A(n4204), .B(n2662), .Z(out[275]) );
  ANDN U4149 ( .B(n2664), .A(n2663), .Z(n2665) );
  XNOR U4150 ( .A(n4228), .B(n2665), .Z(out[276]) );
  AND U4151 ( .A(n2667), .B(n2666), .Z(n2668) );
  XNOR U4152 ( .A(n4252), .B(n2668), .Z(out[277]) );
  AND U4153 ( .A(n2670), .B(n2669), .Z(n2671) );
  XNOR U4154 ( .A(n4276), .B(n2671), .Z(out[278]) );
  AND U4155 ( .A(n2673), .B(n2672), .Z(n2674) );
  XNOR U4156 ( .A(n4300), .B(n2674), .Z(out[279]) );
  XNOR U4157 ( .A(in[1437]), .B(n3690), .Z(n4448) );
  NANDN U4158 ( .A(n2686), .B(n4448), .Z(n2675) );
  XNOR U4159 ( .A(n4449), .B(n2675), .Z(out[27]) );
  AND U4160 ( .A(n2677), .B(n2676), .Z(n2678) );
  XNOR U4161 ( .A(n4324), .B(n2678), .Z(out[280]) );
  AND U4162 ( .A(n2680), .B(n2679), .Z(n2681) );
  XNOR U4163 ( .A(n4356), .B(n2681), .Z(out[281]) );
  AND U4164 ( .A(n2683), .B(n2682), .Z(n2684) );
  XNOR U4165 ( .A(n4404), .B(n2684), .Z(out[282]) );
  AND U4166 ( .A(n2686), .B(n2685), .Z(n2687) );
  XNOR U4167 ( .A(n4448), .B(n2687), .Z(out[283]) );
  XOR U4168 ( .A(in[1438]), .B(n3694), .Z(n4493) );
  NAND U4169 ( .A(n2700), .B(n2688), .Z(n2689) );
  XNOR U4170 ( .A(n4493), .B(n2689), .Z(out[284]) );
  XOR U4171 ( .A(in[1439]), .B(n3698), .Z(n4537) );
  NAND U4172 ( .A(n2722), .B(n2690), .Z(n2691) );
  XNOR U4173 ( .A(n4537), .B(n2691), .Z(out[285]) );
  XOR U4174 ( .A(in[1440]), .B(n3702), .Z(n4581) );
  NAND U4175 ( .A(n2746), .B(n2692), .Z(n2693) );
  XNOR U4176 ( .A(n4581), .B(n2693), .Z(out[286]) );
  XOR U4177 ( .A(in[1441]), .B(n3706), .Z(n4625) );
  NAND U4178 ( .A(n2768), .B(n2694), .Z(n2695) );
  XNOR U4179 ( .A(n4625), .B(n2695), .Z(out[287]) );
  XOR U4180 ( .A(in[1442]), .B(n3714), .Z(n4669) );
  NAND U4181 ( .A(n2780), .B(n2696), .Z(n2697) );
  XNOR U4182 ( .A(n4669), .B(n2697), .Z(out[288]) );
  XOR U4183 ( .A(in[1443]), .B(n3718), .Z(n4713) );
  NAND U4184 ( .A(n2792), .B(n2698), .Z(n2699) );
  XNOR U4185 ( .A(n4713), .B(n2699), .Z(out[289]) );
  OR U4186 ( .A(n4493), .B(n2700), .Z(n2701) );
  XNOR U4187 ( .A(n4492), .B(n2701), .Z(out[28]) );
  XOR U4188 ( .A(in[1444]), .B(n3722), .Z(n4757) );
  NAND U4189 ( .A(n2804), .B(n2702), .Z(n2703) );
  XNOR U4190 ( .A(n4757), .B(n2703), .Z(out[290]) );
  XOR U4191 ( .A(in[1445]), .B(n3726), .Z(n4801) );
  NAND U4192 ( .A(n2816), .B(n2704), .Z(n2705) );
  XNOR U4193 ( .A(n4801), .B(n2705), .Z(out[291]) );
  OR U4194 ( .A(n2829), .B(n2706), .Z(n2707) );
  XNOR U4195 ( .A(n2828), .B(n2707), .Z(out[292]) );
  OR U4196 ( .A(n2843), .B(n2708), .Z(n2709) );
  XNOR U4197 ( .A(n2842), .B(n2709), .Z(out[293]) );
  OR U4198 ( .A(n2857), .B(n2710), .Z(n2711) );
  XNOR U4199 ( .A(n2856), .B(n2711), .Z(out[294]) );
  OR U4200 ( .A(n2871), .B(n2712), .Z(n2713) );
  XNOR U4201 ( .A(n2870), .B(n2713), .Z(out[295]) );
  OR U4202 ( .A(n2887), .B(n2714), .Z(n2715) );
  XNOR U4203 ( .A(n2886), .B(n2715), .Z(out[296]) );
  OR U4204 ( .A(n2901), .B(n2716), .Z(n2717) );
  XNOR U4205 ( .A(n2900), .B(n2717), .Z(out[297]) );
  OR U4206 ( .A(n2915), .B(n2718), .Z(n2719) );
  XNOR U4207 ( .A(n2914), .B(n2719), .Z(out[298]) );
  OR U4208 ( .A(n2929), .B(n2720), .Z(n2721) );
  XNOR U4209 ( .A(n2928), .B(n2721), .Z(out[299]) );
  OR U4210 ( .A(n4537), .B(n2722), .Z(n2723) );
  XNOR U4211 ( .A(n4536), .B(n2723), .Z(out[29]) );
  OR U4212 ( .A(n3665), .B(n2724), .Z(n2725) );
  XNOR U4213 ( .A(n3664), .B(n2725), .Z(out[2]) );
  OR U4214 ( .A(n2945), .B(n2726), .Z(n2727) );
  XNOR U4215 ( .A(n2944), .B(n2727), .Z(out[300]) );
  OR U4216 ( .A(n2969), .B(n2728), .Z(n2729) );
  XNOR U4217 ( .A(n2968), .B(n2729), .Z(out[301]) );
  OR U4218 ( .A(n2993), .B(n2730), .Z(n2731) );
  XNOR U4219 ( .A(n2992), .B(n2731), .Z(out[302]) );
  OR U4220 ( .A(n3017), .B(n2732), .Z(n2733) );
  XNOR U4221 ( .A(n3016), .B(n2733), .Z(out[303]) );
  OR U4222 ( .A(n3041), .B(n2734), .Z(n2735) );
  XNOR U4223 ( .A(n3040), .B(n2735), .Z(out[304]) );
  OR U4224 ( .A(n3065), .B(n2736), .Z(n2737) );
  XNOR U4225 ( .A(n3064), .B(n2737), .Z(out[305]) );
  OR U4226 ( .A(n3091), .B(n2738), .Z(n2739) );
  XNOR U4227 ( .A(n3090), .B(n2739), .Z(out[306]) );
  OR U4228 ( .A(n3115), .B(n2740), .Z(n2741) );
  XNOR U4229 ( .A(n3114), .B(n2741), .Z(out[307]) );
  OR U4230 ( .A(n3139), .B(n2742), .Z(n2743) );
  XNOR U4231 ( .A(n3138), .B(n2743), .Z(out[308]) );
  OR U4232 ( .A(n3163), .B(n2744), .Z(n2745) );
  XNOR U4233 ( .A(n3162), .B(n2745), .Z(out[309]) );
  OR U4234 ( .A(n4581), .B(n2746), .Z(n2747) );
  XNOR U4235 ( .A(n4580), .B(n2747), .Z(out[30]) );
  OR U4236 ( .A(n3187), .B(n2748), .Z(n2749) );
  XNOR U4237 ( .A(n3186), .B(n2749), .Z(out[310]) );
  OR U4238 ( .A(n3211), .B(n2750), .Z(n2751) );
  XNOR U4239 ( .A(n3210), .B(n2751), .Z(out[311]) );
  OR U4240 ( .A(n3235), .B(n2752), .Z(n2753) );
  XNOR U4241 ( .A(n3234), .B(n2753), .Z(out[312]) );
  OR U4242 ( .A(n3267), .B(n2754), .Z(n2755) );
  XNOR U4243 ( .A(n3266), .B(n2755), .Z(out[313]) );
  OR U4244 ( .A(n3311), .B(n2756), .Z(n2757) );
  XNOR U4245 ( .A(n3310), .B(n2757), .Z(out[314]) );
  OR U4246 ( .A(n3355), .B(n2758), .Z(n2759) );
  XNOR U4247 ( .A(n3354), .B(n2759), .Z(out[315]) );
  OR U4248 ( .A(n3401), .B(n2760), .Z(n2761) );
  XNOR U4249 ( .A(n3400), .B(n2761), .Z(out[316]) );
  OR U4250 ( .A(n3445), .B(n2762), .Z(n2763) );
  XNOR U4251 ( .A(n3444), .B(n2763), .Z(out[317]) );
  OR U4252 ( .A(n3489), .B(n2764), .Z(n2765) );
  XNOR U4253 ( .A(n3488), .B(n2765), .Z(out[318]) );
  OR U4254 ( .A(n3533), .B(n2766), .Z(n2767) );
  XNOR U4255 ( .A(n3532), .B(n2767), .Z(out[319]) );
  OR U4256 ( .A(n4625), .B(n2768), .Z(n2769) );
  XNOR U4257 ( .A(n4624), .B(n2769), .Z(out[31]) );
  XNOR U4258 ( .A(in[72]), .B(n4083), .Z(n2940) );
  XOR U4259 ( .A(in[1317]), .B(n3918), .Z(n3253) );
  XOR U4260 ( .A(in[1244]), .B(n3736), .Z(n3250) );
  NAND U4261 ( .A(n3253), .B(n3250), .Z(n2770) );
  XNOR U4262 ( .A(n2940), .B(n2770), .Z(out[320]) );
  XNOR U4263 ( .A(in[73]), .B(n4086), .Z(n2942) );
  XOR U4264 ( .A(in[1318]), .B(n3924), .Z(n3257) );
  XOR U4265 ( .A(in[1245]), .B(n3740), .Z(n3254) );
  NAND U4266 ( .A(n3257), .B(n3254), .Z(n2771) );
  XNOR U4267 ( .A(n2942), .B(n2771), .Z(out[321]) );
  XNOR U4268 ( .A(in[74]), .B(n4089), .Z(n2948) );
  XOR U4269 ( .A(in[1319]), .B(n3926), .Z(n3261) );
  XOR U4270 ( .A(in[1246]), .B(n3744), .Z(n3258) );
  NAND U4271 ( .A(n3261), .B(n3258), .Z(n2772) );
  XNOR U4272 ( .A(n2948), .B(n2772), .Z(out[322]) );
  XNOR U4273 ( .A(in[75]), .B(n4092), .Z(n2950) );
  XOR U4274 ( .A(in[1320]), .B(n3928), .Z(n3265) );
  XOR U4275 ( .A(in[1247]), .B(n3748), .Z(n3262) );
  NAND U4276 ( .A(n3265), .B(n3262), .Z(n2773) );
  XNOR U4277 ( .A(n2950), .B(n2773), .Z(out[323]) );
  XOR U4278 ( .A(n4095), .B(in[76]), .Z(n2952) );
  XOR U4279 ( .A(in[1321]), .B(n3930), .Z(n3273) );
  XOR U4280 ( .A(in[1248]), .B(n3756), .Z(n3270) );
  NAND U4281 ( .A(n3273), .B(n3270), .Z(n2774) );
  XNOR U4282 ( .A(n2952), .B(n2774), .Z(out[324]) );
  XOR U4283 ( .A(n4098), .B(in[77]), .Z(n2954) );
  XOR U4284 ( .A(in[1322]), .B(n3932), .Z(n3277) );
  XOR U4285 ( .A(in[1249]), .B(n3760), .Z(n3274) );
  NAND U4286 ( .A(n3277), .B(n3274), .Z(n2775) );
  XNOR U4287 ( .A(n2954), .B(n2775), .Z(out[325]) );
  XOR U4288 ( .A(n4101), .B(in[78]), .Z(n2956) );
  XOR U4289 ( .A(in[1323]), .B(n3934), .Z(n3281) );
  XOR U4290 ( .A(in[1250]), .B(n3764), .Z(n3278) );
  NAND U4291 ( .A(n3281), .B(n3278), .Z(n2776) );
  XNOR U4292 ( .A(n2956), .B(n2776), .Z(out[326]) );
  XOR U4293 ( .A(n4104), .B(in[79]), .Z(n2958) );
  XOR U4294 ( .A(in[1324]), .B(n3936), .Z(n3285) );
  XOR U4295 ( .A(in[1251]), .B(n3768), .Z(n3282) );
  NAND U4296 ( .A(n3285), .B(n3282), .Z(n2777) );
  XNOR U4297 ( .A(n2958), .B(n2777), .Z(out[327]) );
  XOR U4298 ( .A(n4107), .B(in[80]), .Z(n2960) );
  XOR U4299 ( .A(in[1325]), .B(n3938), .Z(n3289) );
  XOR U4300 ( .A(in[1252]), .B(n3772), .Z(n3286) );
  NAND U4301 ( .A(n3289), .B(n3286), .Z(n2778) );
  XNOR U4302 ( .A(n2960), .B(n2778), .Z(out[328]) );
  XOR U4303 ( .A(n4114), .B(in[81]), .Z(n2962) );
  XOR U4304 ( .A(in[1326]), .B(n3940), .Z(n3293) );
  XNOR U4305 ( .A(in[1253]), .B(n3776), .Z(n3290) );
  NAND U4306 ( .A(n3293), .B(n3290), .Z(n2779) );
  XNOR U4307 ( .A(n2962), .B(n2779), .Z(out[329]) );
  OR U4308 ( .A(n4669), .B(n2780), .Z(n2781) );
  XNOR U4309 ( .A(n4668), .B(n2781), .Z(out[32]) );
  XOR U4310 ( .A(n4117), .B(in[82]), .Z(n2964) );
  XOR U4311 ( .A(in[1327]), .B(n3942), .Z(n3297) );
  XNOR U4312 ( .A(in[1254]), .B(n3780), .Z(n3294) );
  NAND U4313 ( .A(n3297), .B(n3294), .Z(n2782) );
  XNOR U4314 ( .A(n2964), .B(n2782), .Z(out[330]) );
  XOR U4315 ( .A(n4120), .B(in[83]), .Z(n2966) );
  XOR U4316 ( .A(in[1328]), .B(n3948), .Z(n3301) );
  XNOR U4317 ( .A(in[1255]), .B(n3784), .Z(n3298) );
  NAND U4318 ( .A(n3301), .B(n3298), .Z(n2783) );
  XNOR U4319 ( .A(n2966), .B(n2783), .Z(out[331]) );
  XOR U4320 ( .A(in[84]), .B(n4123), .Z(n2972) );
  XOR U4321 ( .A(in[1329]), .B(n3950), .Z(n3305) );
  XNOR U4322 ( .A(in[1256]), .B(n3788), .Z(n3302) );
  NAND U4323 ( .A(n3305), .B(n3302), .Z(n2784) );
  XNOR U4324 ( .A(n2972), .B(n2784), .Z(out[332]) );
  XOR U4325 ( .A(in[85]), .B(n4126), .Z(n2974) );
  XOR U4326 ( .A(in[1330]), .B(n3952), .Z(n3309) );
  XNOR U4327 ( .A(in[1257]), .B(n3792), .Z(n3306) );
  NAND U4328 ( .A(n3309), .B(n3306), .Z(n2785) );
  XNOR U4329 ( .A(n2974), .B(n2785), .Z(out[333]) );
  XOR U4330 ( .A(in[86]), .B(n4129), .Z(n2976) );
  XOR U4331 ( .A(in[1331]), .B(n3954), .Z(n3317) );
  XNOR U4332 ( .A(in[1258]), .B(n3802), .Z(n3314) );
  NAND U4333 ( .A(n3317), .B(n3314), .Z(n2786) );
  XNOR U4334 ( .A(n2976), .B(n2786), .Z(out[334]) );
  XOR U4335 ( .A(in[87]), .B(n4132), .Z(n2978) );
  XOR U4336 ( .A(in[1332]), .B(n3956), .Z(n3321) );
  XNOR U4337 ( .A(in[1259]), .B(n3806), .Z(n3318) );
  NAND U4338 ( .A(n3321), .B(n3318), .Z(n2787) );
  XNOR U4339 ( .A(n2978), .B(n2787), .Z(out[335]) );
  XOR U4340 ( .A(in[88]), .B(n4135), .Z(n2980) );
  XOR U4341 ( .A(in[1333]), .B(n3958), .Z(n3325) );
  XNOR U4342 ( .A(in[1260]), .B(n3810), .Z(n3322) );
  NAND U4343 ( .A(n3325), .B(n3322), .Z(n2788) );
  XNOR U4344 ( .A(n2980), .B(n2788), .Z(out[336]) );
  XOR U4345 ( .A(in[89]), .B(n4138), .Z(n2982) );
  XOR U4346 ( .A(in[1334]), .B(n3960), .Z(n3329) );
  XNOR U4347 ( .A(in[1261]), .B(n3814), .Z(n3326) );
  NAND U4348 ( .A(n3329), .B(n3326), .Z(n2789) );
  XNOR U4349 ( .A(n2982), .B(n2789), .Z(out[337]) );
  XOR U4350 ( .A(in[90]), .B(n4141), .Z(n2984) );
  XOR U4351 ( .A(in[1335]), .B(n3962), .Z(n3333) );
  XNOR U4352 ( .A(in[1262]), .B(n3536), .Z(n3330) );
  NAND U4353 ( .A(n3333), .B(n3330), .Z(n2790) );
  XNOR U4354 ( .A(n2984), .B(n2790), .Z(out[338]) );
  XOR U4355 ( .A(in[91]), .B(n4148), .Z(n2986) );
  XOR U4356 ( .A(in[1336]), .B(n3818), .Z(n3337) );
  XNOR U4357 ( .A(in[1263]), .B(n3540), .Z(n3334) );
  NAND U4358 ( .A(n3337), .B(n3334), .Z(n2791) );
  XNOR U4359 ( .A(n2986), .B(n2791), .Z(out[339]) );
  OR U4360 ( .A(n4713), .B(n2792), .Z(n2793) );
  XNOR U4361 ( .A(n4712), .B(n2793), .Z(out[33]) );
  XOR U4362 ( .A(in[92]), .B(n4151), .Z(n2988) );
  XOR U4363 ( .A(in[1337]), .B(n3820), .Z(n3341) );
  XNOR U4364 ( .A(in[1264]), .B(n3544), .Z(n3338) );
  NAND U4365 ( .A(n3341), .B(n3338), .Z(n2794) );
  XNOR U4366 ( .A(n2988), .B(n2794), .Z(out[340]) );
  XOR U4367 ( .A(in[93]), .B(n4154), .Z(n2990) );
  XOR U4368 ( .A(in[1338]), .B(n3822), .Z(n3345) );
  XNOR U4369 ( .A(in[1265]), .B(n3548), .Z(n3342) );
  NAND U4370 ( .A(n3345), .B(n3342), .Z(n2795) );
  XNOR U4371 ( .A(n2990), .B(n2795), .Z(out[341]) );
  XOR U4372 ( .A(in[94]), .B(n4157), .Z(n2996) );
  XOR U4373 ( .A(in[1339]), .B(n3824), .Z(n3349) );
  XNOR U4374 ( .A(in[1266]), .B(n3552), .Z(n3346) );
  NAND U4375 ( .A(n3349), .B(n3346), .Z(n2796) );
  XNOR U4376 ( .A(n2996), .B(n2796), .Z(out[342]) );
  XOR U4377 ( .A(in[95]), .B(n4160), .Z(n2998) );
  XOR U4378 ( .A(in[1340]), .B(n3826), .Z(n3353) );
  XNOR U4379 ( .A(in[1267]), .B(n3556), .Z(n3350) );
  NAND U4380 ( .A(n3353), .B(n3350), .Z(n2797) );
  XNOR U4381 ( .A(n2998), .B(n2797), .Z(out[343]) );
  XOR U4382 ( .A(in[96]), .B(n4163), .Z(n3000) );
  XOR U4383 ( .A(in[1341]), .B(n3828), .Z(n3363) );
  XNOR U4384 ( .A(in[1268]), .B(n3560), .Z(n3360) );
  NAND U4385 ( .A(n3363), .B(n3360), .Z(n2798) );
  XNOR U4386 ( .A(n3000), .B(n2798), .Z(out[344]) );
  XOR U4387 ( .A(in[97]), .B(n4166), .Z(n3002) );
  XOR U4388 ( .A(in[1342]), .B(n3834), .Z(n3367) );
  XNOR U4389 ( .A(in[1269]), .B(n3564), .Z(n3364) );
  NAND U4390 ( .A(n3367), .B(n3364), .Z(n2799) );
  XNOR U4391 ( .A(n3002), .B(n2799), .Z(out[345]) );
  XOR U4392 ( .A(in[98]), .B(n4169), .Z(n3004) );
  XOR U4393 ( .A(in[1343]), .B(n3836), .Z(n3371) );
  XNOR U4394 ( .A(in[1270]), .B(n3568), .Z(n3368) );
  NAND U4395 ( .A(n3371), .B(n3368), .Z(n2800) );
  XNOR U4396 ( .A(n3004), .B(n2800), .Z(out[346]) );
  XOR U4397 ( .A(in[99]), .B(n4172), .Z(n3006) );
  XOR U4398 ( .A(in[1280]), .B(n3838), .Z(n3375) );
  XNOR U4399 ( .A(in[1271]), .B(n3572), .Z(n3372) );
  NAND U4400 ( .A(n3375), .B(n3372), .Z(n2801) );
  XNOR U4401 ( .A(n3006), .B(n2801), .Z(out[347]) );
  XNOR U4402 ( .A(in[100]), .B(n4175), .Z(n3008) );
  XOR U4403 ( .A(in[1281]), .B(n3840), .Z(n3379) );
  XNOR U4404 ( .A(in[1272]), .B(n3580), .Z(n3376) );
  NAND U4405 ( .A(n3379), .B(n3376), .Z(n2802) );
  XNOR U4406 ( .A(n3008), .B(n2802), .Z(out[348]) );
  XNOR U4407 ( .A(in[101]), .B(n4182), .Z(n3010) );
  XOR U4408 ( .A(in[1282]), .B(n3842), .Z(n3383) );
  XNOR U4409 ( .A(in[1273]), .B(n3584), .Z(n3380) );
  NAND U4410 ( .A(n3383), .B(n3380), .Z(n2803) );
  XNOR U4411 ( .A(n3010), .B(n2803), .Z(out[349]) );
  OR U4412 ( .A(n4757), .B(n2804), .Z(n2805) );
  XNOR U4413 ( .A(n4756), .B(n2805), .Z(out[34]) );
  XNOR U4414 ( .A(in[102]), .B(n4185), .Z(n3012) );
  XOR U4415 ( .A(in[1283]), .B(n3844), .Z(n3387) );
  XNOR U4416 ( .A(in[1274]), .B(n3588), .Z(n3384) );
  NAND U4417 ( .A(n3387), .B(n3384), .Z(n2806) );
  XNOR U4418 ( .A(n3012), .B(n2806), .Z(out[350]) );
  XNOR U4419 ( .A(in[103]), .B(n3964), .Z(n3014) );
  XOR U4420 ( .A(in[1284]), .B(n3846), .Z(n3391) );
  XNOR U4421 ( .A(in[1275]), .B(n3592), .Z(n3388) );
  NAND U4422 ( .A(n3391), .B(n3388), .Z(n2807) );
  XNOR U4423 ( .A(n3014), .B(n2807), .Z(out[351]) );
  XNOR U4424 ( .A(in[104]), .B(n3967), .Z(n3020) );
  XOR U4425 ( .A(in[1285]), .B(n3848), .Z(n3395) );
  XNOR U4426 ( .A(in[1276]), .B(n3596), .Z(n3392) );
  NAND U4427 ( .A(n3395), .B(n3392), .Z(n2808) );
  XNOR U4428 ( .A(n3020), .B(n2808), .Z(out[352]) );
  XNOR U4429 ( .A(in[105]), .B(n3974), .Z(n3022) );
  XOR U4430 ( .A(in[1286]), .B(n3850), .Z(n3399) );
  XNOR U4431 ( .A(in[1277]), .B(n3600), .Z(n3396) );
  NAND U4432 ( .A(n3399), .B(n3396), .Z(n2809) );
  XNOR U4433 ( .A(n3022), .B(n2809), .Z(out[353]) );
  XNOR U4434 ( .A(in[106]), .B(n3977), .Z(n3024) );
  XOR U4435 ( .A(in[1287]), .B(n3852), .Z(n3407) );
  XNOR U4436 ( .A(in[1278]), .B(n3604), .Z(n3404) );
  NAND U4437 ( .A(n3407), .B(n3404), .Z(n2810) );
  XNOR U4438 ( .A(n3024), .B(n2810), .Z(out[354]) );
  XNOR U4439 ( .A(in[107]), .B(n3980), .Z(n3026) );
  XOR U4440 ( .A(in[1288]), .B(n3856), .Z(n3411) );
  XNOR U4441 ( .A(in[1279]), .B(n3608), .Z(n3408) );
  NAND U4442 ( .A(n3411), .B(n3408), .Z(n2811) );
  XNOR U4443 ( .A(n3026), .B(n2811), .Z(out[355]) );
  XNOR U4444 ( .A(in[108]), .B(n3983), .Z(n3028) );
  XOR U4445 ( .A(in[1289]), .B(n3858), .Z(n3415) );
  XNOR U4446 ( .A(in[1216]), .B(n3612), .Z(n3412) );
  NAND U4447 ( .A(n3415), .B(n3412), .Z(n2812) );
  XNOR U4448 ( .A(n3028), .B(n2812), .Z(out[356]) );
  XNOR U4449 ( .A(in[109]), .B(n3986), .Z(n3030) );
  XOR U4450 ( .A(in[1290]), .B(n3860), .Z(n3419) );
  XNOR U4451 ( .A(in[1217]), .B(n3616), .Z(n3416) );
  NAND U4452 ( .A(n3419), .B(n3416), .Z(n2813) );
  XNOR U4453 ( .A(n3030), .B(n2813), .Z(out[357]) );
  XNOR U4454 ( .A(in[110]), .B(n3989), .Z(n3032) );
  XOR U4455 ( .A(in[1291]), .B(n3862), .Z(n3423) );
  XNOR U4456 ( .A(in[1218]), .B(n3624), .Z(n3420) );
  NAND U4457 ( .A(n3423), .B(n3420), .Z(n2814) );
  XNOR U4458 ( .A(n3032), .B(n2814), .Z(out[358]) );
  XNOR U4459 ( .A(in[111]), .B(n3992), .Z(n3034) );
  XOR U4460 ( .A(in[1292]), .B(n3864), .Z(n3427) );
  XNOR U4461 ( .A(in[1219]), .B(n3628), .Z(n3424) );
  NAND U4462 ( .A(n3427), .B(n3424), .Z(n2815) );
  XNOR U4463 ( .A(n3034), .B(n2815), .Z(out[359]) );
  OR U4464 ( .A(n4801), .B(n2816), .Z(n2817) );
  XNOR U4465 ( .A(n4800), .B(n2817), .Z(out[35]) );
  XNOR U4466 ( .A(in[112]), .B(n3995), .Z(n3036) );
  XOR U4467 ( .A(in[1293]), .B(n3866), .Z(n3431) );
  XOR U4468 ( .A(in[1220]), .B(n3632), .Z(n3428) );
  NAND U4469 ( .A(n3431), .B(n3428), .Z(n2818) );
  XNOR U4470 ( .A(n3036), .B(n2818), .Z(out[360]) );
  XNOR U4471 ( .A(in[113]), .B(n3998), .Z(n3038) );
  XOR U4472 ( .A(in[1294]), .B(n3868), .Z(n3435) );
  XOR U4473 ( .A(in[1221]), .B(n3636), .Z(n3432) );
  NAND U4474 ( .A(n3435), .B(n3432), .Z(n2819) );
  XNOR U4475 ( .A(n3038), .B(n2819), .Z(out[361]) );
  XNOR U4476 ( .A(in[114]), .B(n4001), .Z(n3044) );
  XOR U4477 ( .A(in[1295]), .B(n3870), .Z(n3439) );
  XOR U4478 ( .A(in[1222]), .B(n3640), .Z(n3436) );
  NAND U4479 ( .A(n3439), .B(n3436), .Z(n2820) );
  XNOR U4480 ( .A(n3044), .B(n2820), .Z(out[362]) );
  XNOR U4481 ( .A(in[115]), .B(n4008), .Z(n3046) );
  XOR U4482 ( .A(in[1296]), .B(n3872), .Z(n3443) );
  XOR U4483 ( .A(in[1223]), .B(n3644), .Z(n3440) );
  NAND U4484 ( .A(n3443), .B(n3440), .Z(n2821) );
  XNOR U4485 ( .A(n3046), .B(n2821), .Z(out[363]) );
  XNOR U4486 ( .A(in[116]), .B(n4011), .Z(n3048) );
  XOR U4487 ( .A(in[1297]), .B(n3874), .Z(n3451) );
  XOR U4488 ( .A(in[1224]), .B(n3648), .Z(n3448) );
  NAND U4489 ( .A(n3451), .B(n3448), .Z(n2822) );
  XNOR U4490 ( .A(n3048), .B(n2822), .Z(out[364]) );
  XNOR U4491 ( .A(in[117]), .B(n4014), .Z(n3050) );
  XOR U4492 ( .A(in[1298]), .B(n3878), .Z(n3455) );
  XOR U4493 ( .A(in[1225]), .B(n3652), .Z(n3452) );
  NAND U4494 ( .A(n3455), .B(n3452), .Z(n2823) );
  XNOR U4495 ( .A(n3050), .B(n2823), .Z(out[365]) );
  XNOR U4496 ( .A(in[118]), .B(n4017), .Z(n3052) );
  XOR U4497 ( .A(in[1299]), .B(n3880), .Z(n3459) );
  XOR U4498 ( .A(in[1226]), .B(n3656), .Z(n3456) );
  NAND U4499 ( .A(n3459), .B(n3456), .Z(n2824) );
  XNOR U4500 ( .A(n3052), .B(n2824), .Z(out[366]) );
  XNOR U4501 ( .A(in[119]), .B(n4020), .Z(n3054) );
  XOR U4502 ( .A(in[1300]), .B(n3882), .Z(n3463) );
  XOR U4503 ( .A(in[1227]), .B(n3660), .Z(n3460) );
  NAND U4504 ( .A(n3463), .B(n3460), .Z(n2825) );
  XNOR U4505 ( .A(n3054), .B(n2825), .Z(out[367]) );
  XNOR U4506 ( .A(in[120]), .B(n4023), .Z(n3056) );
  XOR U4507 ( .A(in[1301]), .B(n3884), .Z(n3467) );
  XOR U4508 ( .A(in[1228]), .B(n3668), .Z(n3464) );
  NAND U4509 ( .A(n3467), .B(n3464), .Z(n2826) );
  XNOR U4510 ( .A(n3056), .B(n2826), .Z(out[368]) );
  XNOR U4511 ( .A(in[121]), .B(n4026), .Z(n3058) );
  XOR U4512 ( .A(in[1302]), .B(n3886), .Z(n3471) );
  XOR U4513 ( .A(in[1229]), .B(n3672), .Z(n3468) );
  NAND U4514 ( .A(n3471), .B(n3468), .Z(n2827) );
  XNOR U4515 ( .A(n3058), .B(n2827), .Z(out[369]) );
  ANDN U4516 ( .B(n2829), .A(n2828), .Z(n2830) );
  XNOR U4517 ( .A(n2831), .B(n2830), .Z(out[36]) );
  XNOR U4518 ( .A(in[122]), .B(n4029), .Z(n3060) );
  XOR U4519 ( .A(in[1303]), .B(n3888), .Z(n3475) );
  XOR U4520 ( .A(in[1230]), .B(n3676), .Z(n3472) );
  NAND U4521 ( .A(n3475), .B(n3472), .Z(n2832) );
  XNOR U4522 ( .A(n3060), .B(n2832), .Z(out[370]) );
  XNOR U4523 ( .A(in[123]), .B(n4032), .Z(n3062) );
  XOR U4524 ( .A(in[1304]), .B(n3890), .Z(n3479) );
  XOR U4525 ( .A(in[1231]), .B(n3680), .Z(n3476) );
  NAND U4526 ( .A(n3479), .B(n3476), .Z(n2833) );
  XNOR U4527 ( .A(n3062), .B(n2833), .Z(out[371]) );
  XNOR U4528 ( .A(in[124]), .B(n4035), .Z(n3070) );
  XOR U4529 ( .A(in[1305]), .B(n3892), .Z(n3483) );
  XOR U4530 ( .A(in[1232]), .B(n3684), .Z(n3480) );
  NAND U4531 ( .A(n3483), .B(n3480), .Z(n2834) );
  XNOR U4532 ( .A(n3070), .B(n2834), .Z(out[372]) );
  XNOR U4533 ( .A(in[125]), .B(n4042), .Z(n3072) );
  XOR U4534 ( .A(in[1306]), .B(n3894), .Z(n3487) );
  XOR U4535 ( .A(in[1233]), .B(n3688), .Z(n3484) );
  NAND U4536 ( .A(n3487), .B(n3484), .Z(n2835) );
  XNOR U4537 ( .A(n3072), .B(n2835), .Z(out[373]) );
  XNOR U4538 ( .A(in[126]), .B(n4045), .Z(n3074) );
  XOR U4539 ( .A(in[1307]), .B(n3896), .Z(n3495) );
  XOR U4540 ( .A(in[1234]), .B(n3692), .Z(n3492) );
  NAND U4541 ( .A(n3495), .B(n3492), .Z(n2836) );
  XNOR U4542 ( .A(n3074), .B(n2836), .Z(out[374]) );
  XNOR U4543 ( .A(in[127]), .B(n4048), .Z(n3076) );
  XOR U4544 ( .A(in[1308]), .B(n3900), .Z(n3499) );
  XOR U4545 ( .A(in[1235]), .B(n3696), .Z(n3496) );
  NAND U4546 ( .A(n3499), .B(n3496), .Z(n2837) );
  XNOR U4547 ( .A(n3076), .B(n2837), .Z(out[375]) );
  XNOR U4548 ( .A(in[64]), .B(n4051), .Z(n3078) );
  XOR U4549 ( .A(in[1309]), .B(n3902), .Z(n3503) );
  XOR U4550 ( .A(in[1236]), .B(n3700), .Z(n3500) );
  NAND U4551 ( .A(n3503), .B(n3500), .Z(n2838) );
  XNOR U4552 ( .A(n3078), .B(n2838), .Z(out[376]) );
  XNOR U4553 ( .A(in[65]), .B(n4054), .Z(n3080) );
  XOR U4554 ( .A(in[1310]), .B(n3904), .Z(n3507) );
  XOR U4555 ( .A(in[1237]), .B(n3704), .Z(n3504) );
  NAND U4556 ( .A(n3507), .B(n3504), .Z(n2839) );
  XNOR U4557 ( .A(n3080), .B(n2839), .Z(out[377]) );
  XNOR U4558 ( .A(in[66]), .B(n4057), .Z(n3082) );
  XOR U4559 ( .A(in[1311]), .B(n3906), .Z(n3511) );
  XOR U4560 ( .A(in[1238]), .B(n3712), .Z(n3508) );
  NAND U4561 ( .A(n3511), .B(n3508), .Z(n2840) );
  XNOR U4562 ( .A(n3082), .B(n2840), .Z(out[378]) );
  XNOR U4563 ( .A(in[67]), .B(n4060), .Z(n3084) );
  XOR U4564 ( .A(in[1312]), .B(n3908), .Z(n3515) );
  XOR U4565 ( .A(in[1239]), .B(n3716), .Z(n3512) );
  NAND U4566 ( .A(n3515), .B(n3512), .Z(n2841) );
  XNOR U4567 ( .A(n3084), .B(n2841), .Z(out[379]) );
  ANDN U4568 ( .B(n2843), .A(n2842), .Z(n2844) );
  XNOR U4569 ( .A(n2845), .B(n2844), .Z(out[37]) );
  XNOR U4570 ( .A(in[68]), .B(n4063), .Z(n3086) );
  XOR U4571 ( .A(in[1313]), .B(n3910), .Z(n3519) );
  XOR U4572 ( .A(in[1240]), .B(n3720), .Z(n3516) );
  NAND U4573 ( .A(n3519), .B(n3516), .Z(n2846) );
  XNOR U4574 ( .A(n3086), .B(n2846), .Z(out[380]) );
  XNOR U4575 ( .A(in[69]), .B(n4066), .Z(n3088) );
  XOR U4576 ( .A(in[1314]), .B(n3912), .Z(n3523) );
  XOR U4577 ( .A(in[1241]), .B(n3724), .Z(n3520) );
  NAND U4578 ( .A(n3523), .B(n3520), .Z(n2847) );
  XNOR U4579 ( .A(n3088), .B(n2847), .Z(out[381]) );
  XNOR U4580 ( .A(in[70]), .B(n4069), .Z(n3094) );
  XOR U4581 ( .A(in[1315]), .B(n3914), .Z(n3527) );
  XOR U4582 ( .A(in[1242]), .B(n3728), .Z(n3524) );
  NAND U4583 ( .A(n3527), .B(n3524), .Z(n2848) );
  XNOR U4584 ( .A(n3094), .B(n2848), .Z(out[382]) );
  XNOR U4585 ( .A(in[71]), .B(n4080), .Z(n3096) );
  XOR U4586 ( .A(in[1316]), .B(n3916), .Z(n3531) );
  XOR U4587 ( .A(in[1243]), .B(n3732), .Z(n3528) );
  NAND U4588 ( .A(n3531), .B(n3528), .Z(n2849) );
  XNOR U4589 ( .A(n3096), .B(n2849), .Z(out[383]) );
  XOR U4590 ( .A(in[497]), .B(n3778), .Z(n3098) );
  NOR U4591 ( .A(n2940), .B(n3253), .Z(n2850) );
  XNOR U4592 ( .A(n3098), .B(n2850), .Z(out[384]) );
  XOR U4593 ( .A(in[498]), .B(n3782), .Z(n3100) );
  NOR U4594 ( .A(n2942), .B(n3257), .Z(n2851) );
  XNOR U4595 ( .A(n3100), .B(n2851), .Z(out[385]) );
  XOR U4596 ( .A(in[499]), .B(n3786), .Z(n3102) );
  NOR U4597 ( .A(n2948), .B(n3261), .Z(n2852) );
  XNOR U4598 ( .A(n3102), .B(n2852), .Z(out[386]) );
  XOR U4599 ( .A(in[500]), .B(n3790), .Z(n3104) );
  NOR U4600 ( .A(n2950), .B(n3265), .Z(n2853) );
  XNOR U4601 ( .A(n3104), .B(n2853), .Z(out[387]) );
  XOR U4602 ( .A(in[501]), .B(n3794), .Z(n3106) );
  NOR U4603 ( .A(n2952), .B(n3273), .Z(n2854) );
  XNOR U4604 ( .A(n3106), .B(n2854), .Z(out[388]) );
  XOR U4605 ( .A(in[502]), .B(n3804), .Z(n3108) );
  NOR U4606 ( .A(n2954), .B(n3277), .Z(n2855) );
  XNOR U4607 ( .A(n3108), .B(n2855), .Z(out[389]) );
  ANDN U4608 ( .B(n2857), .A(n2856), .Z(n2858) );
  XNOR U4609 ( .A(n2859), .B(n2858), .Z(out[38]) );
  XOR U4610 ( .A(in[503]), .B(n3808), .Z(n3110) );
  NOR U4611 ( .A(n2956), .B(n3281), .Z(n2860) );
  XNOR U4612 ( .A(n3110), .B(n2860), .Z(out[390]) );
  XOR U4613 ( .A(in[504]), .B(n3812), .Z(n3112) );
  NOR U4614 ( .A(n2958), .B(n3285), .Z(n2861) );
  XNOR U4615 ( .A(n3112), .B(n2861), .Z(out[391]) );
  XOR U4616 ( .A(in[505]), .B(n3816), .Z(n3118) );
  NOR U4617 ( .A(n2960), .B(n3289), .Z(n2862) );
  XNOR U4618 ( .A(n3118), .B(n2862), .Z(out[392]) );
  XOR U4619 ( .A(in[506]), .B(n3538), .Z(n3120) );
  NOR U4620 ( .A(n2962), .B(n3293), .Z(n2863) );
  XNOR U4621 ( .A(n3120), .B(n2863), .Z(out[393]) );
  XOR U4622 ( .A(in[507]), .B(n3542), .Z(n3122) );
  NOR U4623 ( .A(n2964), .B(n3297), .Z(n2864) );
  XNOR U4624 ( .A(n3122), .B(n2864), .Z(out[394]) );
  XOR U4625 ( .A(in[508]), .B(n3546), .Z(n3124) );
  NOR U4626 ( .A(n2966), .B(n3301), .Z(n2865) );
  XNOR U4627 ( .A(n3124), .B(n2865), .Z(out[395]) );
  XOR U4628 ( .A(in[509]), .B(n3550), .Z(n3126) );
  NOR U4629 ( .A(n2972), .B(n3305), .Z(n2866) );
  XNOR U4630 ( .A(n3126), .B(n2866), .Z(out[396]) );
  XOR U4631 ( .A(in[510]), .B(n3554), .Z(n3128) );
  NOR U4632 ( .A(n2974), .B(n3309), .Z(n2867) );
  XNOR U4633 ( .A(n3128), .B(n2867), .Z(out[397]) );
  XOR U4634 ( .A(in[511]), .B(n3558), .Z(n3130) );
  NOR U4635 ( .A(n2976), .B(n3317), .Z(n2868) );
  XNOR U4636 ( .A(n3130), .B(n2868), .Z(out[398]) );
  XOR U4637 ( .A(in[448]), .B(n3562), .Z(n3132) );
  NOR U4638 ( .A(n2978), .B(n3321), .Z(n2869) );
  XNOR U4639 ( .A(n3132), .B(n2869), .Z(out[399]) );
  ANDN U4640 ( .B(n2871), .A(n2870), .Z(n2872) );
  XNOR U4641 ( .A(n2873), .B(n2872), .Z(out[39]) );
  OR U4642 ( .A(n3709), .B(n2874), .Z(n2875) );
  XNOR U4643 ( .A(n3708), .B(n2875), .Z(out[3]) );
  XOR U4644 ( .A(in[449]), .B(n3566), .Z(n3134) );
  NOR U4645 ( .A(n2980), .B(n3325), .Z(n2876) );
  XNOR U4646 ( .A(n3134), .B(n2876), .Z(out[400]) );
  XNOR U4647 ( .A(n3570), .B(in[450]), .Z(n3136) );
  NOR U4648 ( .A(n2982), .B(n3329), .Z(n2877) );
  XNOR U4649 ( .A(n3136), .B(n2877), .Z(out[401]) );
  XNOR U4650 ( .A(n3574), .B(in[451]), .Z(n3142) );
  NOR U4651 ( .A(n2984), .B(n3333), .Z(n2878) );
  XNOR U4652 ( .A(n3142), .B(n2878), .Z(out[402]) );
  XNOR U4653 ( .A(n3582), .B(in[452]), .Z(n3144) );
  NOR U4654 ( .A(n2986), .B(n3337), .Z(n2879) );
  XNOR U4655 ( .A(n3144), .B(n2879), .Z(out[403]) );
  XNOR U4656 ( .A(n3586), .B(in[453]), .Z(n3146) );
  NOR U4657 ( .A(n2988), .B(n3341), .Z(n2880) );
  XNOR U4658 ( .A(n3146), .B(n2880), .Z(out[404]) );
  XNOR U4659 ( .A(n3590), .B(in[454]), .Z(n3148) );
  NOR U4660 ( .A(n2990), .B(n3345), .Z(n2881) );
  XNOR U4661 ( .A(n3148), .B(n2881), .Z(out[405]) );
  XNOR U4662 ( .A(n3594), .B(in[455]), .Z(n3150) );
  NOR U4663 ( .A(n2996), .B(n3349), .Z(n2882) );
  XNOR U4664 ( .A(n3150), .B(n2882), .Z(out[406]) );
  XNOR U4665 ( .A(n3598), .B(in[456]), .Z(n3152) );
  NOR U4666 ( .A(n2998), .B(n3353), .Z(n2883) );
  XNOR U4667 ( .A(n3152), .B(n2883), .Z(out[407]) );
  XNOR U4668 ( .A(in[457]), .B(n3602), .Z(n3154) );
  NOR U4669 ( .A(n3000), .B(n3363), .Z(n2884) );
  XNOR U4670 ( .A(n3154), .B(n2884), .Z(out[408]) );
  XNOR U4671 ( .A(n3606), .B(in[458]), .Z(n3156) );
  NOR U4672 ( .A(n3002), .B(n3367), .Z(n2885) );
  XNOR U4673 ( .A(n3156), .B(n2885), .Z(out[409]) );
  ANDN U4674 ( .B(n2887), .A(n2886), .Z(n2888) );
  XNOR U4675 ( .A(n2889), .B(n2888), .Z(out[40]) );
  XNOR U4676 ( .A(n3610), .B(in[459]), .Z(n3158) );
  NOR U4677 ( .A(n3004), .B(n3371), .Z(n2890) );
  XNOR U4678 ( .A(n3158), .B(n2890), .Z(out[410]) );
  XNOR U4679 ( .A(in[460]), .B(n3614), .Z(n3160) );
  NOR U4680 ( .A(n3006), .B(n3375), .Z(n2891) );
  XNOR U4681 ( .A(n3160), .B(n2891), .Z(out[411]) );
  XNOR U4682 ( .A(in[461]), .B(n3618), .Z(n3166) );
  NOR U4683 ( .A(n3008), .B(n3379), .Z(n2892) );
  XNOR U4684 ( .A(n3166), .B(n2892), .Z(out[412]) );
  XNOR U4685 ( .A(in[462]), .B(n3626), .Z(n3168) );
  NOR U4686 ( .A(n3010), .B(n3383), .Z(n2893) );
  XNOR U4687 ( .A(n3168), .B(n2893), .Z(out[413]) );
  XNOR U4688 ( .A(in[463]), .B(n3630), .Z(n3170) );
  NOR U4689 ( .A(n3012), .B(n3387), .Z(n2894) );
  XNOR U4690 ( .A(n3170), .B(n2894), .Z(out[414]) );
  XNOR U4691 ( .A(in[464]), .B(n3634), .Z(n3172) );
  NOR U4692 ( .A(n3014), .B(n3391), .Z(n2895) );
  XNOR U4693 ( .A(n3172), .B(n2895), .Z(out[415]) );
  XNOR U4694 ( .A(in[465]), .B(n3638), .Z(n3174) );
  NOR U4695 ( .A(n3020), .B(n3395), .Z(n2896) );
  XNOR U4696 ( .A(n3174), .B(n2896), .Z(out[416]) );
  XNOR U4697 ( .A(in[466]), .B(n3642), .Z(n3176) );
  NOR U4698 ( .A(n3022), .B(n3399), .Z(n2897) );
  XNOR U4699 ( .A(n3176), .B(n2897), .Z(out[417]) );
  XNOR U4700 ( .A(in[467]), .B(n3646), .Z(n3178) );
  NOR U4701 ( .A(n3024), .B(n3407), .Z(n2898) );
  XNOR U4702 ( .A(n3178), .B(n2898), .Z(out[418]) );
  XNOR U4703 ( .A(in[468]), .B(n3650), .Z(n3180) );
  NOR U4704 ( .A(n3026), .B(n3411), .Z(n2899) );
  XNOR U4705 ( .A(n3180), .B(n2899), .Z(out[419]) );
  ANDN U4706 ( .B(n2901), .A(n2900), .Z(n2902) );
  XNOR U4707 ( .A(n2903), .B(n2902), .Z(out[41]) );
  XNOR U4708 ( .A(in[469]), .B(n3654), .Z(n3182) );
  NOR U4709 ( .A(n3028), .B(n3415), .Z(n2904) );
  XNOR U4710 ( .A(n3182), .B(n2904), .Z(out[420]) );
  XNOR U4711 ( .A(in[470]), .B(n3658), .Z(n3184) );
  NOR U4712 ( .A(n3030), .B(n3419), .Z(n2905) );
  XNOR U4713 ( .A(n3184), .B(n2905), .Z(out[421]) );
  XNOR U4714 ( .A(in[471]), .B(n3662), .Z(n3190) );
  NOR U4715 ( .A(n3032), .B(n3423), .Z(n2906) );
  XNOR U4716 ( .A(n3190), .B(n2906), .Z(out[422]) );
  XNOR U4717 ( .A(in[472]), .B(n3670), .Z(n3192) );
  NOR U4718 ( .A(n3034), .B(n3427), .Z(n2907) );
  XNOR U4719 ( .A(n3192), .B(n2907), .Z(out[423]) );
  XNOR U4720 ( .A(in[473]), .B(n3674), .Z(n3194) );
  NOR U4721 ( .A(n3036), .B(n3431), .Z(n2908) );
  XNOR U4722 ( .A(n3194), .B(n2908), .Z(out[424]) );
  XNOR U4723 ( .A(in[474]), .B(n3678), .Z(n3196) );
  NOR U4724 ( .A(n3038), .B(n3435), .Z(n2909) );
  XNOR U4725 ( .A(n3196), .B(n2909), .Z(out[425]) );
  XNOR U4726 ( .A(in[475]), .B(n3682), .Z(n3198) );
  NOR U4727 ( .A(n3044), .B(n3439), .Z(n2910) );
  XNOR U4728 ( .A(n3198), .B(n2910), .Z(out[426]) );
  XNOR U4729 ( .A(in[476]), .B(n3686), .Z(n3200) );
  NOR U4730 ( .A(n3046), .B(n3443), .Z(n2911) );
  XNOR U4731 ( .A(n3200), .B(n2911), .Z(out[427]) );
  XNOR U4732 ( .A(in[477]), .B(n3690), .Z(n3202) );
  NOR U4733 ( .A(n3048), .B(n3451), .Z(n2912) );
  XNOR U4734 ( .A(n3202), .B(n2912), .Z(out[428]) );
  XNOR U4735 ( .A(in[478]), .B(n3694), .Z(n3204) );
  NOR U4736 ( .A(n3050), .B(n3455), .Z(n2913) );
  XNOR U4737 ( .A(n3204), .B(n2913), .Z(out[429]) );
  ANDN U4738 ( .B(n2915), .A(n2914), .Z(n2916) );
  XNOR U4739 ( .A(n2917), .B(n2916), .Z(out[42]) );
  XNOR U4740 ( .A(in[479]), .B(n3698), .Z(n3206) );
  NOR U4741 ( .A(n3052), .B(n3459), .Z(n2918) );
  XNOR U4742 ( .A(n3206), .B(n2918), .Z(out[430]) );
  XNOR U4743 ( .A(in[480]), .B(n3702), .Z(n3208) );
  NOR U4744 ( .A(n3054), .B(n3463), .Z(n2919) );
  XNOR U4745 ( .A(n3208), .B(n2919), .Z(out[431]) );
  XNOR U4746 ( .A(in[481]), .B(n3706), .Z(n3214) );
  NOR U4747 ( .A(n3056), .B(n3467), .Z(n2920) );
  XNOR U4748 ( .A(n3214), .B(n2920), .Z(out[432]) );
  XNOR U4749 ( .A(in[482]), .B(n3714), .Z(n3216) );
  NOR U4750 ( .A(n3058), .B(n3471), .Z(n2921) );
  XNOR U4751 ( .A(n3216), .B(n2921), .Z(out[433]) );
  XNOR U4752 ( .A(in[483]), .B(n3718), .Z(n3218) );
  NOR U4753 ( .A(n3060), .B(n3475), .Z(n2922) );
  XNOR U4754 ( .A(n3218), .B(n2922), .Z(out[434]) );
  XNOR U4755 ( .A(in[484]), .B(n3722), .Z(n3220) );
  NOR U4756 ( .A(n3062), .B(n3479), .Z(n2923) );
  XNOR U4757 ( .A(n3220), .B(n2923), .Z(out[435]) );
  XNOR U4758 ( .A(in[485]), .B(n3726), .Z(n3222) );
  NOR U4759 ( .A(n3070), .B(n3483), .Z(n2924) );
  XNOR U4760 ( .A(n3222), .B(n2924), .Z(out[436]) );
  XOR U4761 ( .A(in[486]), .B(n3730), .Z(n3224) );
  NOR U4762 ( .A(n3072), .B(n3487), .Z(n2925) );
  XNOR U4763 ( .A(n3224), .B(n2925), .Z(out[437]) );
  XOR U4764 ( .A(in[487]), .B(n3734), .Z(n3226) );
  NOR U4765 ( .A(n3074), .B(n3495), .Z(n2926) );
  XNOR U4766 ( .A(n3226), .B(n2926), .Z(out[438]) );
  XOR U4767 ( .A(in[488]), .B(n3738), .Z(n3228) );
  NOR U4768 ( .A(n3076), .B(n3499), .Z(n2927) );
  XNOR U4769 ( .A(n3228), .B(n2927), .Z(out[439]) );
  ANDN U4770 ( .B(n2929), .A(n2928), .Z(n2930) );
  XNOR U4771 ( .A(n2931), .B(n2930), .Z(out[43]) );
  XOR U4772 ( .A(in[489]), .B(n3742), .Z(n3230) );
  NOR U4773 ( .A(n3078), .B(n3503), .Z(n2932) );
  XNOR U4774 ( .A(n3230), .B(n2932), .Z(out[440]) );
  XOR U4775 ( .A(in[490]), .B(n3746), .Z(n3232) );
  NOR U4776 ( .A(n3080), .B(n3507), .Z(n2933) );
  XNOR U4777 ( .A(n3232), .B(n2933), .Z(out[441]) );
  XOR U4778 ( .A(in[491]), .B(n3750), .Z(n3238) );
  NOR U4779 ( .A(n3082), .B(n3511), .Z(n2934) );
  XNOR U4780 ( .A(n3238), .B(n2934), .Z(out[442]) );
  XOR U4781 ( .A(in[492]), .B(n3758), .Z(n3240) );
  NOR U4782 ( .A(n3084), .B(n3515), .Z(n2935) );
  XNOR U4783 ( .A(n3240), .B(n2935), .Z(out[443]) );
  XOR U4784 ( .A(in[493]), .B(n3762), .Z(n3242) );
  NOR U4785 ( .A(n3086), .B(n3519), .Z(n2936) );
  XNOR U4786 ( .A(n3242), .B(n2936), .Z(out[444]) );
  XOR U4787 ( .A(in[494]), .B(n3766), .Z(n3244) );
  NOR U4788 ( .A(n3088), .B(n3523), .Z(n2937) );
  XNOR U4789 ( .A(n3244), .B(n2937), .Z(out[445]) );
  XOR U4790 ( .A(in[495]), .B(n3770), .Z(n3246) );
  NOR U4791 ( .A(n3094), .B(n3527), .Z(n2938) );
  XNOR U4792 ( .A(n3246), .B(n2938), .Z(out[446]) );
  XOR U4793 ( .A(in[496]), .B(n3774), .Z(n3248) );
  NOR U4794 ( .A(n3096), .B(n3531), .Z(n2939) );
  XNOR U4795 ( .A(n3248), .B(n2939), .Z(out[447]) );
  XNOR U4796 ( .A(in[886]), .B(n3777), .Z(n3251) );
  NAND U4797 ( .A(n3098), .B(n2940), .Z(n2941) );
  XNOR U4798 ( .A(n3251), .B(n2941), .Z(out[448]) );
  XNOR U4799 ( .A(in[887]), .B(n3781), .Z(n3255) );
  NAND U4800 ( .A(n3100), .B(n2942), .Z(n2943) );
  XNOR U4801 ( .A(n3255), .B(n2943), .Z(out[449]) );
  ANDN U4802 ( .B(n2945), .A(n2944), .Z(n2946) );
  XNOR U4803 ( .A(n2947), .B(n2946), .Z(out[44]) );
  XNOR U4804 ( .A(in[888]), .B(n3785), .Z(n3259) );
  NAND U4805 ( .A(n3102), .B(n2948), .Z(n2949) );
  XNOR U4806 ( .A(n3259), .B(n2949), .Z(out[450]) );
  XNOR U4807 ( .A(in[889]), .B(n3789), .Z(n3263) );
  NAND U4808 ( .A(n3104), .B(n2950), .Z(n2951) );
  XNOR U4809 ( .A(n3263), .B(n2951), .Z(out[451]) );
  XNOR U4810 ( .A(in[890]), .B(n3793), .Z(n3271) );
  NAND U4811 ( .A(n3106), .B(n2952), .Z(n2953) );
  XNOR U4812 ( .A(n3271), .B(n2953), .Z(out[452]) );
  XOR U4813 ( .A(in[891]), .B(n3803), .Z(n3275) );
  NAND U4814 ( .A(n3108), .B(n2954), .Z(n2955) );
  XNOR U4815 ( .A(n3275), .B(n2955), .Z(out[453]) );
  XOR U4816 ( .A(in[892]), .B(n3807), .Z(n3279) );
  NAND U4817 ( .A(n3110), .B(n2956), .Z(n2957) );
  XNOR U4818 ( .A(n3279), .B(n2957), .Z(out[454]) );
  XOR U4819 ( .A(in[893]), .B(n3811), .Z(n3283) );
  NAND U4820 ( .A(n3112), .B(n2958), .Z(n2959) );
  XNOR U4821 ( .A(n3283), .B(n2959), .Z(out[455]) );
  XNOR U4822 ( .A(in[894]), .B(n3815), .Z(n3287) );
  NAND U4823 ( .A(n3118), .B(n2960), .Z(n2961) );
  XNOR U4824 ( .A(n3287), .B(n2961), .Z(out[456]) );
  XOR U4825 ( .A(in[895]), .B(n3537), .Z(n3291) );
  NAND U4826 ( .A(n3120), .B(n2962), .Z(n2963) );
  XNOR U4827 ( .A(n3291), .B(n2963), .Z(out[457]) );
  XOR U4828 ( .A(in[832]), .B(n3541), .Z(n3295) );
  NAND U4829 ( .A(n3122), .B(n2964), .Z(n2965) );
  XNOR U4830 ( .A(n3295), .B(n2965), .Z(out[458]) );
  XOR U4831 ( .A(in[833]), .B(n3545), .Z(n3299) );
  NAND U4832 ( .A(n3124), .B(n2966), .Z(n2967) );
  XNOR U4833 ( .A(n3299), .B(n2967), .Z(out[459]) );
  ANDN U4834 ( .B(n2969), .A(n2968), .Z(n2970) );
  XNOR U4835 ( .A(n2971), .B(n2970), .Z(out[45]) );
  XOR U4836 ( .A(in[834]), .B(n3549), .Z(n3303) );
  NAND U4837 ( .A(n3126), .B(n2972), .Z(n2973) );
  XNOR U4838 ( .A(n3303), .B(n2973), .Z(out[460]) );
  XOR U4839 ( .A(in[835]), .B(n3553), .Z(n3307) );
  NAND U4840 ( .A(n3128), .B(n2974), .Z(n2975) );
  XNOR U4841 ( .A(n3307), .B(n2975), .Z(out[461]) );
  XOR U4842 ( .A(in[836]), .B(n3557), .Z(n3315) );
  NAND U4843 ( .A(n3130), .B(n2976), .Z(n2977) );
  XNOR U4844 ( .A(n3315), .B(n2977), .Z(out[462]) );
  XOR U4845 ( .A(in[837]), .B(n3561), .Z(n3319) );
  NAND U4846 ( .A(n3132), .B(n2978), .Z(n2979) );
  XNOR U4847 ( .A(n3319), .B(n2979), .Z(out[463]) );
  XOR U4848 ( .A(in[838]), .B(n3565), .Z(n3323) );
  NAND U4849 ( .A(n3134), .B(n2980), .Z(n2981) );
  XNOR U4850 ( .A(n3323), .B(n2981), .Z(out[464]) );
  XOR U4851 ( .A(in[839]), .B(n3569), .Z(n3327) );
  NAND U4852 ( .A(n3136), .B(n2982), .Z(n2983) );
  XNOR U4853 ( .A(n3327), .B(n2983), .Z(out[465]) );
  XOR U4854 ( .A(in[840]), .B(n3573), .Z(n3331) );
  NAND U4855 ( .A(n3142), .B(n2984), .Z(n2985) );
  XNOR U4856 ( .A(n3331), .B(n2985), .Z(out[466]) );
  XOR U4857 ( .A(in[841]), .B(n3581), .Z(n3335) );
  NAND U4858 ( .A(n3144), .B(n2986), .Z(n2987) );
  XNOR U4859 ( .A(n3335), .B(n2987), .Z(out[467]) );
  XOR U4860 ( .A(in[842]), .B(n3585), .Z(n3339) );
  NAND U4861 ( .A(n3146), .B(n2988), .Z(n2989) );
  XNOR U4862 ( .A(n3339), .B(n2989), .Z(out[468]) );
  XOR U4863 ( .A(in[843]), .B(n3589), .Z(n3343) );
  NAND U4864 ( .A(n3148), .B(n2990), .Z(n2991) );
  XNOR U4865 ( .A(n3343), .B(n2991), .Z(out[469]) );
  ANDN U4866 ( .B(n2993), .A(n2992), .Z(n2994) );
  XNOR U4867 ( .A(n2995), .B(n2994), .Z(out[46]) );
  XOR U4868 ( .A(in[844]), .B(n3593), .Z(n3347) );
  NAND U4869 ( .A(n3150), .B(n2996), .Z(n2997) );
  XNOR U4870 ( .A(n3347), .B(n2997), .Z(out[470]) );
  XOR U4871 ( .A(in[845]), .B(n3597), .Z(n3351) );
  NAND U4872 ( .A(n3152), .B(n2998), .Z(n2999) );
  XNOR U4873 ( .A(n3351), .B(n2999), .Z(out[471]) );
  XOR U4874 ( .A(in[846]), .B(n3601), .Z(n3361) );
  NAND U4875 ( .A(n3154), .B(n3000), .Z(n3001) );
  XNOR U4876 ( .A(n3361), .B(n3001), .Z(out[472]) );
  XOR U4877 ( .A(in[847]), .B(n3605), .Z(n3365) );
  NAND U4878 ( .A(n3156), .B(n3002), .Z(n3003) );
  XNOR U4879 ( .A(n3365), .B(n3003), .Z(out[473]) );
  XOR U4880 ( .A(in[848]), .B(n3609), .Z(n3369) );
  NAND U4881 ( .A(n3158), .B(n3004), .Z(n3005) );
  XNOR U4882 ( .A(n3369), .B(n3005), .Z(out[474]) );
  XOR U4883 ( .A(in[849]), .B(n3613), .Z(n3373) );
  NAND U4884 ( .A(n3160), .B(n3006), .Z(n3007) );
  XNOR U4885 ( .A(n3373), .B(n3007), .Z(out[475]) );
  XOR U4886 ( .A(in[850]), .B(n3617), .Z(n3377) );
  NAND U4887 ( .A(n3166), .B(n3008), .Z(n3009) );
  XNOR U4888 ( .A(n3377), .B(n3009), .Z(out[476]) );
  XNOR U4889 ( .A(in[851]), .B(n3625), .Z(n3381) );
  NAND U4890 ( .A(n3168), .B(n3010), .Z(n3011) );
  XNOR U4891 ( .A(n3381), .B(n3011), .Z(out[477]) );
  XNOR U4892 ( .A(in[852]), .B(n3629), .Z(n3385) );
  NAND U4893 ( .A(n3170), .B(n3012), .Z(n3013) );
  XNOR U4894 ( .A(n3385), .B(n3013), .Z(out[478]) );
  XNOR U4895 ( .A(in[853]), .B(n3633), .Z(n3389) );
  NAND U4896 ( .A(n3172), .B(n3014), .Z(n3015) );
  XNOR U4897 ( .A(n3389), .B(n3015), .Z(out[479]) );
  ANDN U4898 ( .B(n3017), .A(n3016), .Z(n3018) );
  XNOR U4899 ( .A(n3019), .B(n3018), .Z(out[47]) );
  XNOR U4900 ( .A(in[854]), .B(n3637), .Z(n3393) );
  NAND U4901 ( .A(n3174), .B(n3020), .Z(n3021) );
  XNOR U4902 ( .A(n3393), .B(n3021), .Z(out[480]) );
  XNOR U4903 ( .A(in[855]), .B(n3641), .Z(n3397) );
  NAND U4904 ( .A(n3176), .B(n3022), .Z(n3023) );
  XNOR U4905 ( .A(n3397), .B(n3023), .Z(out[481]) );
  XNOR U4906 ( .A(in[856]), .B(n3645), .Z(n3405) );
  NAND U4907 ( .A(n3178), .B(n3024), .Z(n3025) );
  XNOR U4908 ( .A(n3405), .B(n3025), .Z(out[482]) );
  XNOR U4909 ( .A(in[857]), .B(n3649), .Z(n3409) );
  NAND U4910 ( .A(n3180), .B(n3026), .Z(n3027) );
  XNOR U4911 ( .A(n3409), .B(n3027), .Z(out[483]) );
  XNOR U4912 ( .A(in[858]), .B(n3653), .Z(n3413) );
  NAND U4913 ( .A(n3182), .B(n3028), .Z(n3029) );
  XNOR U4914 ( .A(n3413), .B(n3029), .Z(out[484]) );
  XNOR U4915 ( .A(in[859]), .B(n3657), .Z(n3417) );
  NAND U4916 ( .A(n3184), .B(n3030), .Z(n3031) );
  XNOR U4917 ( .A(n3417), .B(n3031), .Z(out[485]) );
  XNOR U4918 ( .A(in[860]), .B(n3661), .Z(n3421) );
  NAND U4919 ( .A(n3190), .B(n3032), .Z(n3033) );
  XNOR U4920 ( .A(n3421), .B(n3033), .Z(out[486]) );
  XNOR U4921 ( .A(in[861]), .B(n3669), .Z(n3425) );
  NAND U4922 ( .A(n3192), .B(n3034), .Z(n3035) );
  XNOR U4923 ( .A(n3425), .B(n3035), .Z(out[487]) );
  XNOR U4924 ( .A(in[862]), .B(n3673), .Z(n3429) );
  NAND U4925 ( .A(n3194), .B(n3036), .Z(n3037) );
  XNOR U4926 ( .A(n3429), .B(n3037), .Z(out[488]) );
  XNOR U4927 ( .A(in[863]), .B(n3677), .Z(n3433) );
  NAND U4928 ( .A(n3196), .B(n3038), .Z(n3039) );
  XNOR U4929 ( .A(n3433), .B(n3039), .Z(out[489]) );
  ANDN U4930 ( .B(n3041), .A(n3040), .Z(n3042) );
  XNOR U4931 ( .A(n3043), .B(n3042), .Z(out[48]) );
  XNOR U4932 ( .A(in[864]), .B(n3681), .Z(n3437) );
  NAND U4933 ( .A(n3198), .B(n3044), .Z(n3045) );
  XNOR U4934 ( .A(n3437), .B(n3045), .Z(out[490]) );
  XNOR U4935 ( .A(in[865]), .B(n3685), .Z(n3441) );
  NAND U4936 ( .A(n3200), .B(n3046), .Z(n3047) );
  XNOR U4937 ( .A(n3441), .B(n3047), .Z(out[491]) );
  XOR U4938 ( .A(n3689), .B(in[866]), .Z(n3449) );
  NAND U4939 ( .A(n3202), .B(n3048), .Z(n3049) );
  XNOR U4940 ( .A(n3449), .B(n3049), .Z(out[492]) );
  XOR U4941 ( .A(n3693), .B(in[867]), .Z(n3453) );
  NAND U4942 ( .A(n3204), .B(n3050), .Z(n3051) );
  XNOR U4943 ( .A(n3453), .B(n3051), .Z(out[493]) );
  XOR U4944 ( .A(n3697), .B(in[868]), .Z(n3457) );
  NAND U4945 ( .A(n3206), .B(n3052), .Z(n3053) );
  XNOR U4946 ( .A(n3457), .B(n3053), .Z(out[494]) );
  XOR U4947 ( .A(n3701), .B(in[869]), .Z(n3461) );
  NAND U4948 ( .A(n3208), .B(n3054), .Z(n3055) );
  XNOR U4949 ( .A(n3461), .B(n3055), .Z(out[495]) );
  XNOR U4950 ( .A(in[870]), .B(n3705), .Z(n3465) );
  NAND U4951 ( .A(n3214), .B(n3056), .Z(n3057) );
  XNOR U4952 ( .A(n3465), .B(n3057), .Z(out[496]) );
  XNOR U4953 ( .A(in[871]), .B(n3713), .Z(n3469) );
  NAND U4954 ( .A(n3216), .B(n3058), .Z(n3059) );
  XNOR U4955 ( .A(n3469), .B(n3059), .Z(out[497]) );
  XNOR U4956 ( .A(in[872]), .B(n3717), .Z(n3473) );
  NAND U4957 ( .A(n3218), .B(n3060), .Z(n3061) );
  XNOR U4958 ( .A(n3473), .B(n3061), .Z(out[498]) );
  XNOR U4959 ( .A(in[873]), .B(n3721), .Z(n3477) );
  NAND U4960 ( .A(n3220), .B(n3062), .Z(n3063) );
  XNOR U4961 ( .A(n3477), .B(n3063), .Z(out[499]) );
  ANDN U4962 ( .B(n3065), .A(n3064), .Z(n3066) );
  XNOR U4963 ( .A(n3067), .B(n3066), .Z(out[49]) );
  OR U4964 ( .A(n3753), .B(n3068), .Z(n3069) );
  XNOR U4965 ( .A(n3752), .B(n3069), .Z(out[4]) );
  XNOR U4966 ( .A(in[874]), .B(n3725), .Z(n3481) );
  NAND U4967 ( .A(n3222), .B(n3070), .Z(n3071) );
  XNOR U4968 ( .A(n3481), .B(n3071), .Z(out[500]) );
  XNOR U4969 ( .A(in[875]), .B(n3729), .Z(n3485) );
  NAND U4970 ( .A(n3224), .B(n3072), .Z(n3073) );
  XNOR U4971 ( .A(n3485), .B(n3073), .Z(out[501]) );
  XNOR U4972 ( .A(in[876]), .B(n3733), .Z(n3493) );
  NAND U4973 ( .A(n3226), .B(n3074), .Z(n3075) );
  XNOR U4974 ( .A(n3493), .B(n3075), .Z(out[502]) );
  XNOR U4975 ( .A(in[877]), .B(n3737), .Z(n3497) );
  NAND U4976 ( .A(n3228), .B(n3076), .Z(n3077) );
  XNOR U4977 ( .A(n3497), .B(n3077), .Z(out[503]) );
  XNOR U4978 ( .A(in[878]), .B(n3741), .Z(n3501) );
  NAND U4979 ( .A(n3230), .B(n3078), .Z(n3079) );
  XNOR U4980 ( .A(n3501), .B(n3079), .Z(out[504]) );
  XNOR U4981 ( .A(in[879]), .B(n3745), .Z(n3505) );
  NAND U4982 ( .A(n3232), .B(n3080), .Z(n3081) );
  XNOR U4983 ( .A(n3505), .B(n3081), .Z(out[505]) );
  XNOR U4984 ( .A(in[880]), .B(n3749), .Z(n3509) );
  NAND U4985 ( .A(n3238), .B(n3082), .Z(n3083) );
  XNOR U4986 ( .A(n3509), .B(n3083), .Z(out[506]) );
  XNOR U4987 ( .A(in[881]), .B(n3757), .Z(n3513) );
  NAND U4988 ( .A(n3240), .B(n3084), .Z(n3085) );
  XNOR U4989 ( .A(n3513), .B(n3085), .Z(out[507]) );
  XNOR U4990 ( .A(in[882]), .B(n3761), .Z(n3517) );
  NAND U4991 ( .A(n3242), .B(n3086), .Z(n3087) );
  XNOR U4992 ( .A(n3517), .B(n3087), .Z(out[508]) );
  XNOR U4993 ( .A(in[883]), .B(n3765), .Z(n3521) );
  NAND U4994 ( .A(n3244), .B(n3088), .Z(n3089) );
  XNOR U4995 ( .A(n3521), .B(n3089), .Z(out[509]) );
  ANDN U4996 ( .B(n3091), .A(n3090), .Z(n3092) );
  XNOR U4997 ( .A(n3093), .B(n3092), .Z(out[50]) );
  XNOR U4998 ( .A(in[884]), .B(n3769), .Z(n3525) );
  NAND U4999 ( .A(n3246), .B(n3094), .Z(n3095) );
  XNOR U5000 ( .A(n3525), .B(n3095), .Z(out[510]) );
  XNOR U5001 ( .A(in[885]), .B(n3773), .Z(n3529) );
  NAND U5002 ( .A(n3248), .B(n3096), .Z(n3097) );
  XNOR U5003 ( .A(n3529), .B(n3097), .Z(out[511]) );
  OR U5004 ( .A(n3251), .B(n3098), .Z(n3099) );
  XNOR U5005 ( .A(n3250), .B(n3099), .Z(out[512]) );
  OR U5006 ( .A(n3255), .B(n3100), .Z(n3101) );
  XNOR U5007 ( .A(n3254), .B(n3101), .Z(out[513]) );
  OR U5008 ( .A(n3259), .B(n3102), .Z(n3103) );
  XNOR U5009 ( .A(n3258), .B(n3103), .Z(out[514]) );
  OR U5010 ( .A(n3263), .B(n3104), .Z(n3105) );
  XNOR U5011 ( .A(n3262), .B(n3105), .Z(out[515]) );
  OR U5012 ( .A(n3271), .B(n3106), .Z(n3107) );
  XNOR U5013 ( .A(n3270), .B(n3107), .Z(out[516]) );
  OR U5014 ( .A(n3275), .B(n3108), .Z(n3109) );
  XNOR U5015 ( .A(n3274), .B(n3109), .Z(out[517]) );
  OR U5016 ( .A(n3279), .B(n3110), .Z(n3111) );
  XNOR U5017 ( .A(n3278), .B(n3111), .Z(out[518]) );
  OR U5018 ( .A(n3283), .B(n3112), .Z(n3113) );
  XNOR U5019 ( .A(n3282), .B(n3113), .Z(out[519]) );
  ANDN U5020 ( .B(n3115), .A(n3114), .Z(n3116) );
  XNOR U5021 ( .A(n3117), .B(n3116), .Z(out[51]) );
  OR U5022 ( .A(n3287), .B(n3118), .Z(n3119) );
  XNOR U5023 ( .A(n3286), .B(n3119), .Z(out[520]) );
  OR U5024 ( .A(n3291), .B(n3120), .Z(n3121) );
  XNOR U5025 ( .A(n3290), .B(n3121), .Z(out[521]) );
  OR U5026 ( .A(n3295), .B(n3122), .Z(n3123) );
  XNOR U5027 ( .A(n3294), .B(n3123), .Z(out[522]) );
  OR U5028 ( .A(n3299), .B(n3124), .Z(n3125) );
  XNOR U5029 ( .A(n3298), .B(n3125), .Z(out[523]) );
  OR U5030 ( .A(n3303), .B(n3126), .Z(n3127) );
  XNOR U5031 ( .A(n3302), .B(n3127), .Z(out[524]) );
  OR U5032 ( .A(n3307), .B(n3128), .Z(n3129) );
  XNOR U5033 ( .A(n3306), .B(n3129), .Z(out[525]) );
  OR U5034 ( .A(n3315), .B(n3130), .Z(n3131) );
  XNOR U5035 ( .A(n3314), .B(n3131), .Z(out[526]) );
  OR U5036 ( .A(n3319), .B(n3132), .Z(n3133) );
  XNOR U5037 ( .A(n3318), .B(n3133), .Z(out[527]) );
  OR U5038 ( .A(n3323), .B(n3134), .Z(n3135) );
  XNOR U5039 ( .A(n3322), .B(n3135), .Z(out[528]) );
  OR U5040 ( .A(n3327), .B(n3136), .Z(n3137) );
  XNOR U5041 ( .A(n3326), .B(n3137), .Z(out[529]) );
  ANDN U5042 ( .B(n3139), .A(n3138), .Z(n3140) );
  XNOR U5043 ( .A(n3141), .B(n3140), .Z(out[52]) );
  OR U5044 ( .A(n3331), .B(n3142), .Z(n3143) );
  XNOR U5045 ( .A(n3330), .B(n3143), .Z(out[530]) );
  OR U5046 ( .A(n3335), .B(n3144), .Z(n3145) );
  XNOR U5047 ( .A(n3334), .B(n3145), .Z(out[531]) );
  OR U5048 ( .A(n3339), .B(n3146), .Z(n3147) );
  XNOR U5049 ( .A(n3338), .B(n3147), .Z(out[532]) );
  OR U5050 ( .A(n3343), .B(n3148), .Z(n3149) );
  XNOR U5051 ( .A(n3342), .B(n3149), .Z(out[533]) );
  OR U5052 ( .A(n3347), .B(n3150), .Z(n3151) );
  XNOR U5053 ( .A(n3346), .B(n3151), .Z(out[534]) );
  OR U5054 ( .A(n3351), .B(n3152), .Z(n3153) );
  XNOR U5055 ( .A(n3350), .B(n3153), .Z(out[535]) );
  OR U5056 ( .A(n3361), .B(n3154), .Z(n3155) );
  XNOR U5057 ( .A(n3360), .B(n3155), .Z(out[536]) );
  OR U5058 ( .A(n3365), .B(n3156), .Z(n3157) );
  XNOR U5059 ( .A(n3364), .B(n3157), .Z(out[537]) );
  OR U5060 ( .A(n3369), .B(n3158), .Z(n3159) );
  XNOR U5061 ( .A(n3368), .B(n3159), .Z(out[538]) );
  OR U5062 ( .A(n3373), .B(n3160), .Z(n3161) );
  XNOR U5063 ( .A(n3372), .B(n3161), .Z(out[539]) );
  ANDN U5064 ( .B(n3163), .A(n3162), .Z(n3164) );
  XNOR U5065 ( .A(n3165), .B(n3164), .Z(out[53]) );
  OR U5066 ( .A(n3377), .B(n3166), .Z(n3167) );
  XNOR U5067 ( .A(n3376), .B(n3167), .Z(out[540]) );
  OR U5068 ( .A(n3381), .B(n3168), .Z(n3169) );
  XNOR U5069 ( .A(n3380), .B(n3169), .Z(out[541]) );
  OR U5070 ( .A(n3385), .B(n3170), .Z(n3171) );
  XNOR U5071 ( .A(n3384), .B(n3171), .Z(out[542]) );
  OR U5072 ( .A(n3389), .B(n3172), .Z(n3173) );
  XNOR U5073 ( .A(n3388), .B(n3173), .Z(out[543]) );
  OR U5074 ( .A(n3393), .B(n3174), .Z(n3175) );
  XNOR U5075 ( .A(n3392), .B(n3175), .Z(out[544]) );
  OR U5076 ( .A(n3397), .B(n3176), .Z(n3177) );
  XNOR U5077 ( .A(n3396), .B(n3177), .Z(out[545]) );
  OR U5078 ( .A(n3405), .B(n3178), .Z(n3179) );
  XNOR U5079 ( .A(n3404), .B(n3179), .Z(out[546]) );
  OR U5080 ( .A(n3409), .B(n3180), .Z(n3181) );
  XNOR U5081 ( .A(n3408), .B(n3181), .Z(out[547]) );
  OR U5082 ( .A(n3413), .B(n3182), .Z(n3183) );
  XNOR U5083 ( .A(n3412), .B(n3183), .Z(out[548]) );
  OR U5084 ( .A(n3417), .B(n3184), .Z(n3185) );
  XNOR U5085 ( .A(n3416), .B(n3185), .Z(out[549]) );
  ANDN U5086 ( .B(n3187), .A(n3186), .Z(n3188) );
  XNOR U5087 ( .A(n3189), .B(n3188), .Z(out[54]) );
  OR U5088 ( .A(n3421), .B(n3190), .Z(n3191) );
  XNOR U5089 ( .A(n3420), .B(n3191), .Z(out[550]) );
  OR U5090 ( .A(n3425), .B(n3192), .Z(n3193) );
  XNOR U5091 ( .A(n3424), .B(n3193), .Z(out[551]) );
  OR U5092 ( .A(n3429), .B(n3194), .Z(n3195) );
  XNOR U5093 ( .A(n3428), .B(n3195), .Z(out[552]) );
  OR U5094 ( .A(n3433), .B(n3196), .Z(n3197) );
  XNOR U5095 ( .A(n3432), .B(n3197), .Z(out[553]) );
  OR U5096 ( .A(n3437), .B(n3198), .Z(n3199) );
  XNOR U5097 ( .A(n3436), .B(n3199), .Z(out[554]) );
  OR U5098 ( .A(n3441), .B(n3200), .Z(n3201) );
  XNOR U5099 ( .A(n3440), .B(n3201), .Z(out[555]) );
  OR U5100 ( .A(n3449), .B(n3202), .Z(n3203) );
  XNOR U5101 ( .A(n3448), .B(n3203), .Z(out[556]) );
  OR U5102 ( .A(n3453), .B(n3204), .Z(n3205) );
  XNOR U5103 ( .A(n3452), .B(n3205), .Z(out[557]) );
  OR U5104 ( .A(n3457), .B(n3206), .Z(n3207) );
  XNOR U5105 ( .A(n3456), .B(n3207), .Z(out[558]) );
  OR U5106 ( .A(n3461), .B(n3208), .Z(n3209) );
  XNOR U5107 ( .A(n3460), .B(n3209), .Z(out[559]) );
  ANDN U5108 ( .B(n3211), .A(n3210), .Z(n3212) );
  XNOR U5109 ( .A(n3213), .B(n3212), .Z(out[55]) );
  OR U5110 ( .A(n3465), .B(n3214), .Z(n3215) );
  XNOR U5111 ( .A(n3464), .B(n3215), .Z(out[560]) );
  OR U5112 ( .A(n3469), .B(n3216), .Z(n3217) );
  XNOR U5113 ( .A(n3468), .B(n3217), .Z(out[561]) );
  OR U5114 ( .A(n3473), .B(n3218), .Z(n3219) );
  XNOR U5115 ( .A(n3472), .B(n3219), .Z(out[562]) );
  OR U5116 ( .A(n3477), .B(n3220), .Z(n3221) );
  XNOR U5117 ( .A(n3476), .B(n3221), .Z(out[563]) );
  OR U5118 ( .A(n3481), .B(n3222), .Z(n3223) );
  XNOR U5119 ( .A(n3480), .B(n3223), .Z(out[564]) );
  OR U5120 ( .A(n3485), .B(n3224), .Z(n3225) );
  XNOR U5121 ( .A(n3484), .B(n3225), .Z(out[565]) );
  OR U5122 ( .A(n3493), .B(n3226), .Z(n3227) );
  XNOR U5123 ( .A(n3492), .B(n3227), .Z(out[566]) );
  OR U5124 ( .A(n3497), .B(n3228), .Z(n3229) );
  XNOR U5125 ( .A(n3496), .B(n3229), .Z(out[567]) );
  OR U5126 ( .A(n3501), .B(n3230), .Z(n3231) );
  XNOR U5127 ( .A(n3500), .B(n3231), .Z(out[568]) );
  OR U5128 ( .A(n3505), .B(n3232), .Z(n3233) );
  XNOR U5129 ( .A(n3504), .B(n3233), .Z(out[569]) );
  ANDN U5130 ( .B(n3235), .A(n3234), .Z(n3236) );
  XNOR U5131 ( .A(n3237), .B(n3236), .Z(out[56]) );
  OR U5132 ( .A(n3509), .B(n3238), .Z(n3239) );
  XNOR U5133 ( .A(n3508), .B(n3239), .Z(out[570]) );
  OR U5134 ( .A(n3513), .B(n3240), .Z(n3241) );
  XNOR U5135 ( .A(n3512), .B(n3241), .Z(out[571]) );
  OR U5136 ( .A(n3517), .B(n3242), .Z(n3243) );
  XNOR U5137 ( .A(n3516), .B(n3243), .Z(out[572]) );
  OR U5138 ( .A(n3521), .B(n3244), .Z(n3245) );
  XNOR U5139 ( .A(n3520), .B(n3245), .Z(out[573]) );
  OR U5140 ( .A(n3525), .B(n3246), .Z(n3247) );
  XNOR U5141 ( .A(n3524), .B(n3247), .Z(out[574]) );
  OR U5142 ( .A(n3529), .B(n3248), .Z(n3249) );
  XNOR U5143 ( .A(n3528), .B(n3249), .Z(out[575]) );
  ANDN U5144 ( .B(n3251), .A(n3250), .Z(n3252) );
  XNOR U5145 ( .A(n3253), .B(n3252), .Z(out[576]) );
  ANDN U5146 ( .B(n3255), .A(n3254), .Z(n3256) );
  XNOR U5147 ( .A(n3257), .B(n3256), .Z(out[577]) );
  ANDN U5148 ( .B(n3259), .A(n3258), .Z(n3260) );
  XNOR U5149 ( .A(n3261), .B(n3260), .Z(out[578]) );
  ANDN U5150 ( .B(n3263), .A(n3262), .Z(n3264) );
  XNOR U5151 ( .A(n3265), .B(n3264), .Z(out[579]) );
  ANDN U5152 ( .B(n3267), .A(n3266), .Z(n3268) );
  XNOR U5153 ( .A(n3269), .B(n3268), .Z(out[57]) );
  ANDN U5154 ( .B(n3271), .A(n3270), .Z(n3272) );
  XNOR U5155 ( .A(n3273), .B(n3272), .Z(out[580]) );
  ANDN U5156 ( .B(n3275), .A(n3274), .Z(n3276) );
  XNOR U5157 ( .A(n3277), .B(n3276), .Z(out[581]) );
  ANDN U5158 ( .B(n3279), .A(n3278), .Z(n3280) );
  XNOR U5159 ( .A(n3281), .B(n3280), .Z(out[582]) );
  ANDN U5160 ( .B(n3283), .A(n3282), .Z(n3284) );
  XNOR U5161 ( .A(n3285), .B(n3284), .Z(out[583]) );
  ANDN U5162 ( .B(n3287), .A(n3286), .Z(n3288) );
  XNOR U5163 ( .A(n3289), .B(n3288), .Z(out[584]) );
  ANDN U5164 ( .B(n3291), .A(n3290), .Z(n3292) );
  XNOR U5165 ( .A(n3293), .B(n3292), .Z(out[585]) );
  ANDN U5166 ( .B(n3295), .A(n3294), .Z(n3296) );
  XNOR U5167 ( .A(n3297), .B(n3296), .Z(out[586]) );
  ANDN U5168 ( .B(n3299), .A(n3298), .Z(n3300) );
  XNOR U5169 ( .A(n3301), .B(n3300), .Z(out[587]) );
  ANDN U5170 ( .B(n3303), .A(n3302), .Z(n3304) );
  XNOR U5171 ( .A(n3305), .B(n3304), .Z(out[588]) );
  ANDN U5172 ( .B(n3307), .A(n3306), .Z(n3308) );
  XNOR U5173 ( .A(n3309), .B(n3308), .Z(out[589]) );
  ANDN U5174 ( .B(n3311), .A(n3310), .Z(n3312) );
  XNOR U5175 ( .A(n3313), .B(n3312), .Z(out[58]) );
  ANDN U5176 ( .B(n3315), .A(n3314), .Z(n3316) );
  XNOR U5177 ( .A(n3317), .B(n3316), .Z(out[590]) );
  ANDN U5178 ( .B(n3319), .A(n3318), .Z(n3320) );
  XNOR U5179 ( .A(n3321), .B(n3320), .Z(out[591]) );
  ANDN U5180 ( .B(n3323), .A(n3322), .Z(n3324) );
  XNOR U5181 ( .A(n3325), .B(n3324), .Z(out[592]) );
  ANDN U5182 ( .B(n3327), .A(n3326), .Z(n3328) );
  XNOR U5183 ( .A(n3329), .B(n3328), .Z(out[593]) );
  ANDN U5184 ( .B(n3331), .A(n3330), .Z(n3332) );
  XNOR U5185 ( .A(n3333), .B(n3332), .Z(out[594]) );
  ANDN U5186 ( .B(n3335), .A(n3334), .Z(n3336) );
  XNOR U5187 ( .A(n3337), .B(n3336), .Z(out[595]) );
  ANDN U5188 ( .B(n3339), .A(n3338), .Z(n3340) );
  XNOR U5189 ( .A(n3341), .B(n3340), .Z(out[596]) );
  ANDN U5190 ( .B(n3343), .A(n3342), .Z(n3344) );
  XNOR U5191 ( .A(n3345), .B(n3344), .Z(out[597]) );
  ANDN U5192 ( .B(n3347), .A(n3346), .Z(n3348) );
  XNOR U5193 ( .A(n3349), .B(n3348), .Z(out[598]) );
  ANDN U5194 ( .B(n3351), .A(n3350), .Z(n3352) );
  XNOR U5195 ( .A(n3353), .B(n3352), .Z(out[599]) );
  ANDN U5196 ( .B(n3355), .A(n3354), .Z(n3356) );
  XNOR U5197 ( .A(n3357), .B(n3356), .Z(out[59]) );
  OR U5198 ( .A(n3797), .B(n3358), .Z(n3359) );
  XNOR U5199 ( .A(n3796), .B(n3359), .Z(out[5]) );
  ANDN U5200 ( .B(n3361), .A(n3360), .Z(n3362) );
  XNOR U5201 ( .A(n3363), .B(n3362), .Z(out[600]) );
  ANDN U5202 ( .B(n3365), .A(n3364), .Z(n3366) );
  XNOR U5203 ( .A(n3367), .B(n3366), .Z(out[601]) );
  ANDN U5204 ( .B(n3369), .A(n3368), .Z(n3370) );
  XNOR U5205 ( .A(n3371), .B(n3370), .Z(out[602]) );
  ANDN U5206 ( .B(n3373), .A(n3372), .Z(n3374) );
  XNOR U5207 ( .A(n3375), .B(n3374), .Z(out[603]) );
  ANDN U5208 ( .B(n3377), .A(n3376), .Z(n3378) );
  XNOR U5209 ( .A(n3379), .B(n3378), .Z(out[604]) );
  ANDN U5210 ( .B(n3381), .A(n3380), .Z(n3382) );
  XNOR U5211 ( .A(n3383), .B(n3382), .Z(out[605]) );
  ANDN U5212 ( .B(n3385), .A(n3384), .Z(n3386) );
  XNOR U5213 ( .A(n3387), .B(n3386), .Z(out[606]) );
  ANDN U5214 ( .B(n3389), .A(n3388), .Z(n3390) );
  XNOR U5215 ( .A(n3391), .B(n3390), .Z(out[607]) );
  ANDN U5216 ( .B(n3393), .A(n3392), .Z(n3394) );
  XNOR U5217 ( .A(n3395), .B(n3394), .Z(out[608]) );
  ANDN U5218 ( .B(n3397), .A(n3396), .Z(n3398) );
  XNOR U5219 ( .A(n3399), .B(n3398), .Z(out[609]) );
  ANDN U5220 ( .B(n3401), .A(n3400), .Z(n3402) );
  XNOR U5221 ( .A(n3403), .B(n3402), .Z(out[60]) );
  ANDN U5222 ( .B(n3405), .A(n3404), .Z(n3406) );
  XNOR U5223 ( .A(n3407), .B(n3406), .Z(out[610]) );
  ANDN U5224 ( .B(n3409), .A(n3408), .Z(n3410) );
  XNOR U5225 ( .A(n3411), .B(n3410), .Z(out[611]) );
  ANDN U5226 ( .B(n3413), .A(n3412), .Z(n3414) );
  XNOR U5227 ( .A(n3415), .B(n3414), .Z(out[612]) );
  ANDN U5228 ( .B(n3417), .A(n3416), .Z(n3418) );
  XNOR U5229 ( .A(n3419), .B(n3418), .Z(out[613]) );
  ANDN U5230 ( .B(n3421), .A(n3420), .Z(n3422) );
  XNOR U5231 ( .A(n3423), .B(n3422), .Z(out[614]) );
  ANDN U5232 ( .B(n3425), .A(n3424), .Z(n3426) );
  XNOR U5233 ( .A(n3427), .B(n3426), .Z(out[615]) );
  ANDN U5234 ( .B(n3429), .A(n3428), .Z(n3430) );
  XNOR U5235 ( .A(n3431), .B(n3430), .Z(out[616]) );
  ANDN U5236 ( .B(n3433), .A(n3432), .Z(n3434) );
  XNOR U5237 ( .A(n3435), .B(n3434), .Z(out[617]) );
  ANDN U5238 ( .B(n3437), .A(n3436), .Z(n3438) );
  XNOR U5239 ( .A(n3439), .B(n3438), .Z(out[618]) );
  ANDN U5240 ( .B(n3441), .A(n3440), .Z(n3442) );
  XNOR U5241 ( .A(n3443), .B(n3442), .Z(out[619]) );
  ANDN U5242 ( .B(n3445), .A(n3444), .Z(n3446) );
  XNOR U5243 ( .A(n3447), .B(n3446), .Z(out[61]) );
  ANDN U5244 ( .B(n3449), .A(n3448), .Z(n3450) );
  XNOR U5245 ( .A(n3451), .B(n3450), .Z(out[620]) );
  ANDN U5246 ( .B(n3453), .A(n3452), .Z(n3454) );
  XNOR U5247 ( .A(n3455), .B(n3454), .Z(out[621]) );
  ANDN U5248 ( .B(n3457), .A(n3456), .Z(n3458) );
  XNOR U5249 ( .A(n3459), .B(n3458), .Z(out[622]) );
  ANDN U5250 ( .B(n3461), .A(n3460), .Z(n3462) );
  XNOR U5251 ( .A(n3463), .B(n3462), .Z(out[623]) );
  ANDN U5252 ( .B(n3465), .A(n3464), .Z(n3466) );
  XNOR U5253 ( .A(n3467), .B(n3466), .Z(out[624]) );
  ANDN U5254 ( .B(n3469), .A(n3468), .Z(n3470) );
  XNOR U5255 ( .A(n3471), .B(n3470), .Z(out[625]) );
  ANDN U5256 ( .B(n3473), .A(n3472), .Z(n3474) );
  XNOR U5257 ( .A(n3475), .B(n3474), .Z(out[626]) );
  ANDN U5258 ( .B(n3477), .A(n3476), .Z(n3478) );
  XNOR U5259 ( .A(n3479), .B(n3478), .Z(out[627]) );
  ANDN U5260 ( .B(n3481), .A(n3480), .Z(n3482) );
  XNOR U5261 ( .A(n3483), .B(n3482), .Z(out[628]) );
  ANDN U5262 ( .B(n3485), .A(n3484), .Z(n3486) );
  XNOR U5263 ( .A(n3487), .B(n3486), .Z(out[629]) );
  ANDN U5264 ( .B(n3489), .A(n3488), .Z(n3490) );
  XNOR U5265 ( .A(n3491), .B(n3490), .Z(out[62]) );
  ANDN U5266 ( .B(n3493), .A(n3492), .Z(n3494) );
  XNOR U5267 ( .A(n3495), .B(n3494), .Z(out[630]) );
  ANDN U5268 ( .B(n3497), .A(n3496), .Z(n3498) );
  XNOR U5269 ( .A(n3499), .B(n3498), .Z(out[631]) );
  ANDN U5270 ( .B(n3501), .A(n3500), .Z(n3502) );
  XNOR U5271 ( .A(n3503), .B(n3502), .Z(out[632]) );
  ANDN U5272 ( .B(n3505), .A(n3504), .Z(n3506) );
  XNOR U5273 ( .A(n3507), .B(n3506), .Z(out[633]) );
  ANDN U5274 ( .B(n3509), .A(n3508), .Z(n3510) );
  XNOR U5275 ( .A(n3511), .B(n3510), .Z(out[634]) );
  ANDN U5276 ( .B(n3513), .A(n3512), .Z(n3514) );
  XNOR U5277 ( .A(n3515), .B(n3514), .Z(out[635]) );
  ANDN U5278 ( .B(n3517), .A(n3516), .Z(n3518) );
  XNOR U5279 ( .A(n3519), .B(n3518), .Z(out[636]) );
  ANDN U5280 ( .B(n3521), .A(n3520), .Z(n3522) );
  XNOR U5281 ( .A(n3523), .B(n3522), .Z(out[637]) );
  ANDN U5282 ( .B(n3525), .A(n3524), .Z(n3526) );
  XNOR U5283 ( .A(n3527), .B(n3526), .Z(out[638]) );
  ANDN U5284 ( .B(n3529), .A(n3528), .Z(n3530) );
  XNOR U5285 ( .A(n3531), .B(n3530), .Z(out[639]) );
  ANDN U5286 ( .B(n3533), .A(n3532), .Z(n3534) );
  XNOR U5287 ( .A(n3535), .B(n3534), .Z(out[63]) );
  XNOR U5288 ( .A(in[302]), .B(n3536), .Z(n3965) );
  XNOR U5289 ( .A(in[1535]), .B(n3537), .Z(n4343) );
  XNOR U5290 ( .A(in[1146]), .B(n3538), .Z(n4340) );
  NAND U5291 ( .A(n4343), .B(n4340), .Z(n3539) );
  XNOR U5292 ( .A(n3965), .B(n3539), .Z(out[640]) );
  XNOR U5293 ( .A(in[303]), .B(n3540), .Z(n3968) );
  XNOR U5294 ( .A(in[1472]), .B(n3541), .Z(n4347) );
  XNOR U5295 ( .A(in[1147]), .B(n3542), .Z(n4344) );
  NAND U5296 ( .A(n4347), .B(n4344), .Z(n3543) );
  XNOR U5297 ( .A(n3968), .B(n3543), .Z(out[641]) );
  XNOR U5298 ( .A(in[304]), .B(n3544), .Z(n3975) );
  XNOR U5299 ( .A(in[1473]), .B(n3545), .Z(n4351) );
  XNOR U5300 ( .A(in[1148]), .B(n3546), .Z(n4348) );
  NAND U5301 ( .A(n4351), .B(n4348), .Z(n3547) );
  XNOR U5302 ( .A(n3975), .B(n3547), .Z(out[642]) );
  XNOR U5303 ( .A(in[305]), .B(n3548), .Z(n3978) );
  XNOR U5304 ( .A(in[1474]), .B(n3549), .Z(n4355) );
  XNOR U5305 ( .A(in[1149]), .B(n3550), .Z(n4352) );
  NAND U5306 ( .A(n4355), .B(n4352), .Z(n3551) );
  XNOR U5307 ( .A(n3978), .B(n3551), .Z(out[643]) );
  XNOR U5308 ( .A(in[306]), .B(n3552), .Z(n3981) );
  XNOR U5309 ( .A(in[1475]), .B(n3553), .Z(n4367) );
  XNOR U5310 ( .A(in[1150]), .B(n3554), .Z(n4364) );
  NAND U5311 ( .A(n4367), .B(n4364), .Z(n3555) );
  XNOR U5312 ( .A(n3981), .B(n3555), .Z(out[644]) );
  XNOR U5313 ( .A(in[307]), .B(n3556), .Z(n3984) );
  XNOR U5314 ( .A(in[1476]), .B(n3557), .Z(n4371) );
  XNOR U5315 ( .A(in[1151]), .B(n3558), .Z(n4368) );
  NAND U5316 ( .A(n4371), .B(n4368), .Z(n3559) );
  XNOR U5317 ( .A(n3984), .B(n3559), .Z(out[645]) );
  XNOR U5318 ( .A(in[308]), .B(n3560), .Z(n3987) );
  XNOR U5319 ( .A(in[1477]), .B(n3561), .Z(n4375) );
  XNOR U5320 ( .A(in[1088]), .B(n3562), .Z(n4372) );
  NAND U5321 ( .A(n4375), .B(n4372), .Z(n3563) );
  XNOR U5322 ( .A(n3987), .B(n3563), .Z(out[646]) );
  XNOR U5323 ( .A(in[309]), .B(n3564), .Z(n3990) );
  XNOR U5324 ( .A(in[1478]), .B(n3565), .Z(n4379) );
  XNOR U5325 ( .A(in[1089]), .B(n3566), .Z(n4376) );
  NAND U5326 ( .A(n4379), .B(n4376), .Z(n3567) );
  XNOR U5327 ( .A(n3990), .B(n3567), .Z(out[647]) );
  XNOR U5328 ( .A(in[310]), .B(n3568), .Z(n3993) );
  XNOR U5329 ( .A(in[1479]), .B(n3569), .Z(n4383) );
  XOR U5330 ( .A(n3570), .B(in[1090]), .Z(n4380) );
  NAND U5331 ( .A(n4383), .B(n4380), .Z(n3571) );
  XNOR U5332 ( .A(n3993), .B(n3571), .Z(out[648]) );
  XNOR U5333 ( .A(in[311]), .B(n3572), .Z(n3996) );
  XNOR U5334 ( .A(in[1480]), .B(n3573), .Z(n4387) );
  XOR U5335 ( .A(n3574), .B(in[1091]), .Z(n4384) );
  NAND U5336 ( .A(n4387), .B(n4384), .Z(n3575) );
  XNOR U5337 ( .A(n3996), .B(n3575), .Z(out[649]) );
  NOR U5338 ( .A(n3577), .B(n3576), .Z(n3578) );
  XNOR U5339 ( .A(n3579), .B(n3578), .Z(out[64]) );
  XNOR U5340 ( .A(in[312]), .B(n3580), .Z(n3999) );
  XNOR U5341 ( .A(in[1481]), .B(n3581), .Z(n4391) );
  XOR U5342 ( .A(n3582), .B(in[1092]), .Z(n4388) );
  NAND U5343 ( .A(n4391), .B(n4388), .Z(n3583) );
  XNOR U5344 ( .A(n3999), .B(n3583), .Z(out[650]) );
  XNOR U5345 ( .A(in[313]), .B(n3584), .Z(n4002) );
  XNOR U5346 ( .A(in[1482]), .B(n3585), .Z(n4395) );
  XOR U5347 ( .A(n3586), .B(in[1093]), .Z(n4392) );
  NAND U5348 ( .A(n4395), .B(n4392), .Z(n3587) );
  XNOR U5349 ( .A(n4002), .B(n3587), .Z(out[651]) );
  XNOR U5350 ( .A(in[314]), .B(n3588), .Z(n4009) );
  XNOR U5351 ( .A(in[1483]), .B(n3589), .Z(n4399) );
  XOR U5352 ( .A(n3590), .B(in[1094]), .Z(n4396) );
  NAND U5353 ( .A(n4399), .B(n4396), .Z(n3591) );
  XNOR U5354 ( .A(n4009), .B(n3591), .Z(out[652]) );
  XNOR U5355 ( .A(in[315]), .B(n3592), .Z(n4012) );
  XNOR U5356 ( .A(in[1484]), .B(n3593), .Z(n4403) );
  XOR U5357 ( .A(n3594), .B(in[1095]), .Z(n4400) );
  NAND U5358 ( .A(n4403), .B(n4400), .Z(n3595) );
  XNOR U5359 ( .A(n4012), .B(n3595), .Z(out[653]) );
  XNOR U5360 ( .A(in[316]), .B(n3596), .Z(n4015) );
  XNOR U5361 ( .A(in[1485]), .B(n3597), .Z(n4411) );
  XOR U5362 ( .A(n3598), .B(in[1096]), .Z(n4408) );
  NAND U5363 ( .A(n4411), .B(n4408), .Z(n3599) );
  XNOR U5364 ( .A(n4015), .B(n3599), .Z(out[654]) );
  XNOR U5365 ( .A(in[317]), .B(n3600), .Z(n4018) );
  XNOR U5366 ( .A(in[1486]), .B(n3601), .Z(n4415) );
  XOR U5367 ( .A(in[1097]), .B(n3602), .Z(n4412) );
  NAND U5368 ( .A(n4415), .B(n4412), .Z(n3603) );
  XNOR U5369 ( .A(n4018), .B(n3603), .Z(out[655]) );
  XNOR U5370 ( .A(in[318]), .B(n3604), .Z(n4021) );
  XNOR U5371 ( .A(in[1487]), .B(n3605), .Z(n4419) );
  XOR U5372 ( .A(n3606), .B(in[1098]), .Z(n4416) );
  NAND U5373 ( .A(n4419), .B(n4416), .Z(n3607) );
  XNOR U5374 ( .A(n4021), .B(n3607), .Z(out[656]) );
  XNOR U5375 ( .A(in[319]), .B(n3608), .Z(n4024) );
  XNOR U5376 ( .A(in[1488]), .B(n3609), .Z(n4423) );
  XOR U5377 ( .A(n3610), .B(in[1099]), .Z(n4420) );
  NAND U5378 ( .A(n4423), .B(n4420), .Z(n3611) );
  XNOR U5379 ( .A(n4024), .B(n3611), .Z(out[657]) );
  XNOR U5380 ( .A(in[256]), .B(n3612), .Z(n4027) );
  XNOR U5381 ( .A(in[1489]), .B(n3613), .Z(n4427) );
  XOR U5382 ( .A(in[1100]), .B(n3614), .Z(n4424) );
  NAND U5383 ( .A(n4427), .B(n4424), .Z(n3615) );
  XNOR U5384 ( .A(n4027), .B(n3615), .Z(out[658]) );
  XNOR U5385 ( .A(in[257]), .B(n3616), .Z(n4030) );
  XNOR U5386 ( .A(in[1490]), .B(n3617), .Z(n4431) );
  XOR U5387 ( .A(in[1101]), .B(n3618), .Z(n4428) );
  NAND U5388 ( .A(n4431), .B(n4428), .Z(n3619) );
  XNOR U5389 ( .A(n4030), .B(n3619), .Z(out[659]) );
  NOR U5390 ( .A(n3621), .B(n3620), .Z(n3622) );
  XNOR U5391 ( .A(n3623), .B(n3622), .Z(out[65]) );
  XNOR U5392 ( .A(in[258]), .B(n3624), .Z(n4033) );
  XOR U5393 ( .A(in[1491]), .B(n3625), .Z(n4435) );
  XOR U5394 ( .A(in[1102]), .B(n3626), .Z(n4432) );
  NAND U5395 ( .A(n4435), .B(n4432), .Z(n3627) );
  XNOR U5396 ( .A(n4033), .B(n3627), .Z(out[660]) );
  XNOR U5397 ( .A(in[259]), .B(n3628), .Z(n4036) );
  XOR U5398 ( .A(in[1492]), .B(n3629), .Z(n4439) );
  XOR U5399 ( .A(in[1103]), .B(n3630), .Z(n4436) );
  NAND U5400 ( .A(n4439), .B(n4436), .Z(n3631) );
  XNOR U5401 ( .A(n4036), .B(n3631), .Z(out[661]) );
  XOR U5402 ( .A(in[260]), .B(n3632), .Z(n4043) );
  XOR U5403 ( .A(in[1493]), .B(n3633), .Z(n4443) );
  XOR U5404 ( .A(in[1104]), .B(n3634), .Z(n4440) );
  NAND U5405 ( .A(n4443), .B(n4440), .Z(n3635) );
  XNOR U5406 ( .A(n4043), .B(n3635), .Z(out[662]) );
  XOR U5407 ( .A(in[261]), .B(n3636), .Z(n4046) );
  XOR U5408 ( .A(in[1494]), .B(n3637), .Z(n4447) );
  XOR U5409 ( .A(in[1105]), .B(n3638), .Z(n4444) );
  NAND U5410 ( .A(n4447), .B(n4444), .Z(n3639) );
  XNOR U5411 ( .A(n4046), .B(n3639), .Z(out[663]) );
  XOR U5412 ( .A(in[262]), .B(n3640), .Z(n4049) );
  XOR U5413 ( .A(in[1495]), .B(n3641), .Z(n4455) );
  XOR U5414 ( .A(in[1106]), .B(n3642), .Z(n4452) );
  NAND U5415 ( .A(n4455), .B(n4452), .Z(n3643) );
  XNOR U5416 ( .A(n4049), .B(n3643), .Z(out[664]) );
  XOR U5417 ( .A(in[263]), .B(n3644), .Z(n4052) );
  XOR U5418 ( .A(in[1496]), .B(n3645), .Z(n4459) );
  XOR U5419 ( .A(in[1107]), .B(n3646), .Z(n4456) );
  NAND U5420 ( .A(n4459), .B(n4456), .Z(n3647) );
  XNOR U5421 ( .A(n4052), .B(n3647), .Z(out[665]) );
  XOR U5422 ( .A(in[264]), .B(n3648), .Z(n4055) );
  XOR U5423 ( .A(in[1497]), .B(n3649), .Z(n4463) );
  XOR U5424 ( .A(in[1108]), .B(n3650), .Z(n4460) );
  NAND U5425 ( .A(n4463), .B(n4460), .Z(n3651) );
  XNOR U5426 ( .A(n4055), .B(n3651), .Z(out[666]) );
  XOR U5427 ( .A(in[265]), .B(n3652), .Z(n4058) );
  XOR U5428 ( .A(in[1498]), .B(n3653), .Z(n4467) );
  XOR U5429 ( .A(in[1109]), .B(n3654), .Z(n4464) );
  NAND U5430 ( .A(n4467), .B(n4464), .Z(n3655) );
  XNOR U5431 ( .A(n4058), .B(n3655), .Z(out[667]) );
  XOR U5432 ( .A(in[266]), .B(n3656), .Z(n4061) );
  XOR U5433 ( .A(in[1499]), .B(n3657), .Z(n4471) );
  XOR U5434 ( .A(in[1110]), .B(n3658), .Z(n4468) );
  NAND U5435 ( .A(n4471), .B(n4468), .Z(n3659) );
  XNOR U5436 ( .A(n4061), .B(n3659), .Z(out[668]) );
  XOR U5437 ( .A(in[267]), .B(n3660), .Z(n4064) );
  XOR U5438 ( .A(in[1500]), .B(n3661), .Z(n4475) );
  XOR U5439 ( .A(in[1111]), .B(n3662), .Z(n4472) );
  NAND U5440 ( .A(n4475), .B(n4472), .Z(n3663) );
  XNOR U5441 ( .A(n4064), .B(n3663), .Z(out[669]) );
  ANDN U5442 ( .B(n3665), .A(n3664), .Z(n3666) );
  XNOR U5443 ( .A(n3667), .B(n3666), .Z(out[66]) );
  XOR U5444 ( .A(in[268]), .B(n3668), .Z(n4067) );
  XOR U5445 ( .A(in[1501]), .B(n3669), .Z(n4479) );
  XOR U5446 ( .A(in[1112]), .B(n3670), .Z(n4476) );
  NAND U5447 ( .A(n4479), .B(n4476), .Z(n3671) );
  XNOR U5448 ( .A(n4067), .B(n3671), .Z(out[670]) );
  XOR U5449 ( .A(in[269]), .B(n3672), .Z(n4070) );
  XOR U5450 ( .A(in[1502]), .B(n3673), .Z(n4483) );
  XOR U5451 ( .A(in[1113]), .B(n3674), .Z(n4480) );
  NAND U5452 ( .A(n4483), .B(n4480), .Z(n3675) );
  XNOR U5453 ( .A(n4070), .B(n3675), .Z(out[671]) );
  XOR U5454 ( .A(in[270]), .B(n3676), .Z(n4081) );
  XOR U5455 ( .A(in[1503]), .B(n3677), .Z(n4487) );
  XOR U5456 ( .A(in[1114]), .B(n3678), .Z(n4484) );
  NAND U5457 ( .A(n4487), .B(n4484), .Z(n3679) );
  XNOR U5458 ( .A(n4081), .B(n3679), .Z(out[672]) );
  XOR U5459 ( .A(in[271]), .B(n3680), .Z(n4084) );
  XOR U5460 ( .A(in[1504]), .B(n3681), .Z(n4491) );
  XOR U5461 ( .A(in[1115]), .B(n3682), .Z(n4488) );
  NAND U5462 ( .A(n4491), .B(n4488), .Z(n3683) );
  XNOR U5463 ( .A(n4084), .B(n3683), .Z(out[673]) );
  XOR U5464 ( .A(in[272]), .B(n3684), .Z(n4087) );
  XOR U5465 ( .A(in[1505]), .B(n3685), .Z(n4499) );
  XOR U5466 ( .A(in[1116]), .B(n3686), .Z(n4496) );
  NAND U5467 ( .A(n4499), .B(n4496), .Z(n3687) );
  XNOR U5468 ( .A(n4087), .B(n3687), .Z(out[674]) );
  XOR U5469 ( .A(in[273]), .B(n3688), .Z(n4090) );
  XNOR U5470 ( .A(n3689), .B(in[1506]), .Z(n4503) );
  XOR U5471 ( .A(in[1117]), .B(n3690), .Z(n4500) );
  NAND U5472 ( .A(n4503), .B(n4500), .Z(n3691) );
  XNOR U5473 ( .A(n4090), .B(n3691), .Z(out[675]) );
  XOR U5474 ( .A(in[274]), .B(n3692), .Z(n4093) );
  XNOR U5475 ( .A(n3693), .B(in[1507]), .Z(n4507) );
  XOR U5476 ( .A(in[1118]), .B(n3694), .Z(n4504) );
  NAND U5477 ( .A(n4507), .B(n4504), .Z(n3695) );
  XNOR U5478 ( .A(n4093), .B(n3695), .Z(out[676]) );
  XOR U5479 ( .A(in[275]), .B(n3696), .Z(n4096) );
  XNOR U5480 ( .A(n3697), .B(in[1508]), .Z(n4511) );
  XOR U5481 ( .A(in[1119]), .B(n3698), .Z(n4508) );
  NAND U5482 ( .A(n4511), .B(n4508), .Z(n3699) );
  XNOR U5483 ( .A(n4096), .B(n3699), .Z(out[677]) );
  XOR U5484 ( .A(in[276]), .B(n3700), .Z(n4099) );
  XNOR U5485 ( .A(n3701), .B(in[1509]), .Z(n4515) );
  XOR U5486 ( .A(in[1120]), .B(n3702), .Z(n4512) );
  NAND U5487 ( .A(n4515), .B(n4512), .Z(n3703) );
  XNOR U5488 ( .A(n4099), .B(n3703), .Z(out[678]) );
  XOR U5489 ( .A(in[277]), .B(n3704), .Z(n4102) );
  XOR U5490 ( .A(in[1510]), .B(n3705), .Z(n4519) );
  XOR U5491 ( .A(in[1121]), .B(n3706), .Z(n4516) );
  NAND U5492 ( .A(n4519), .B(n4516), .Z(n3707) );
  XNOR U5493 ( .A(n4102), .B(n3707), .Z(out[679]) );
  ANDN U5494 ( .B(n3709), .A(n3708), .Z(n3710) );
  XNOR U5495 ( .A(n3711), .B(n3710), .Z(out[67]) );
  XOR U5496 ( .A(in[278]), .B(n3712), .Z(n4105) );
  XOR U5497 ( .A(in[1511]), .B(n3713), .Z(n4523) );
  XOR U5498 ( .A(in[1122]), .B(n3714), .Z(n4520) );
  NAND U5499 ( .A(n4523), .B(n4520), .Z(n3715) );
  XNOR U5500 ( .A(n4105), .B(n3715), .Z(out[680]) );
  XOR U5501 ( .A(in[279]), .B(n3716), .Z(n4108) );
  XOR U5502 ( .A(in[1512]), .B(n3717), .Z(n4527) );
  XOR U5503 ( .A(in[1123]), .B(n3718), .Z(n4524) );
  NAND U5504 ( .A(n4527), .B(n4524), .Z(n3719) );
  XNOR U5505 ( .A(n4108), .B(n3719), .Z(out[681]) );
  XOR U5506 ( .A(in[280]), .B(n3720), .Z(n4115) );
  XOR U5507 ( .A(in[1513]), .B(n3721), .Z(n4531) );
  XOR U5508 ( .A(in[1124]), .B(n3722), .Z(n4528) );
  NAND U5509 ( .A(n4531), .B(n4528), .Z(n3723) );
  XNOR U5510 ( .A(n4115), .B(n3723), .Z(out[682]) );
  XOR U5511 ( .A(in[281]), .B(n3724), .Z(n4118) );
  XOR U5512 ( .A(in[1514]), .B(n3725), .Z(n4535) );
  XOR U5513 ( .A(in[1125]), .B(n3726), .Z(n4532) );
  NAND U5514 ( .A(n4535), .B(n4532), .Z(n3727) );
  XNOR U5515 ( .A(n4118), .B(n3727), .Z(out[683]) );
  XOR U5516 ( .A(in[282]), .B(n3728), .Z(n4121) );
  XOR U5517 ( .A(in[1515]), .B(n3729), .Z(n4543) );
  XNOR U5518 ( .A(in[1126]), .B(n3730), .Z(n4540) );
  NAND U5519 ( .A(n4543), .B(n4540), .Z(n3731) );
  XNOR U5520 ( .A(n4121), .B(n3731), .Z(out[684]) );
  XOR U5521 ( .A(in[283]), .B(n3732), .Z(n4124) );
  XOR U5522 ( .A(in[1516]), .B(n3733), .Z(n4547) );
  XNOR U5523 ( .A(in[1127]), .B(n3734), .Z(n4544) );
  NAND U5524 ( .A(n4547), .B(n4544), .Z(n3735) );
  XNOR U5525 ( .A(n4124), .B(n3735), .Z(out[685]) );
  XOR U5526 ( .A(in[284]), .B(n3736), .Z(n4127) );
  XOR U5527 ( .A(in[1517]), .B(n3737), .Z(n4551) );
  XNOR U5528 ( .A(in[1128]), .B(n3738), .Z(n4548) );
  NAND U5529 ( .A(n4551), .B(n4548), .Z(n3739) );
  XNOR U5530 ( .A(n4127), .B(n3739), .Z(out[686]) );
  XOR U5531 ( .A(in[285]), .B(n3740), .Z(n4130) );
  XOR U5532 ( .A(in[1518]), .B(n3741), .Z(n4555) );
  XNOR U5533 ( .A(in[1129]), .B(n3742), .Z(n4552) );
  NAND U5534 ( .A(n4555), .B(n4552), .Z(n3743) );
  XNOR U5535 ( .A(n4130), .B(n3743), .Z(out[687]) );
  XOR U5536 ( .A(in[286]), .B(n3744), .Z(n4133) );
  XOR U5537 ( .A(in[1519]), .B(n3745), .Z(n4559) );
  XNOR U5538 ( .A(in[1130]), .B(n3746), .Z(n4556) );
  NAND U5539 ( .A(n4559), .B(n4556), .Z(n3747) );
  XNOR U5540 ( .A(n4133), .B(n3747), .Z(out[688]) );
  XOR U5541 ( .A(in[287]), .B(n3748), .Z(n4136) );
  XOR U5542 ( .A(in[1520]), .B(n3749), .Z(n4563) );
  XNOR U5543 ( .A(in[1131]), .B(n3750), .Z(n4560) );
  NAND U5544 ( .A(n4563), .B(n4560), .Z(n3751) );
  XNOR U5545 ( .A(n4136), .B(n3751), .Z(out[689]) );
  ANDN U5546 ( .B(n3753), .A(n3752), .Z(n3754) );
  XNOR U5547 ( .A(n3755), .B(n3754), .Z(out[68]) );
  XOR U5548 ( .A(in[288]), .B(n3756), .Z(n4139) );
  XOR U5549 ( .A(in[1521]), .B(n3757), .Z(n4567) );
  XNOR U5550 ( .A(in[1132]), .B(n3758), .Z(n4564) );
  NAND U5551 ( .A(n4567), .B(n4564), .Z(n3759) );
  XNOR U5552 ( .A(n4139), .B(n3759), .Z(out[690]) );
  XOR U5553 ( .A(in[289]), .B(n3760), .Z(n4142) );
  XOR U5554 ( .A(in[1522]), .B(n3761), .Z(n4571) );
  XNOR U5555 ( .A(in[1133]), .B(n3762), .Z(n4568) );
  NAND U5556 ( .A(n4571), .B(n4568), .Z(n3763) );
  XNOR U5557 ( .A(n4142), .B(n3763), .Z(out[691]) );
  XOR U5558 ( .A(in[290]), .B(n3764), .Z(n4149) );
  XOR U5559 ( .A(in[1523]), .B(n3765), .Z(n4575) );
  XNOR U5560 ( .A(in[1134]), .B(n3766), .Z(n4572) );
  NAND U5561 ( .A(n4575), .B(n4572), .Z(n3767) );
  XNOR U5562 ( .A(n4149), .B(n3767), .Z(out[692]) );
  XOR U5563 ( .A(in[291]), .B(n3768), .Z(n4152) );
  XOR U5564 ( .A(in[1524]), .B(n3769), .Z(n4579) );
  XNOR U5565 ( .A(in[1135]), .B(n3770), .Z(n4576) );
  NAND U5566 ( .A(n4579), .B(n4576), .Z(n3771) );
  XNOR U5567 ( .A(n4152), .B(n3771), .Z(out[693]) );
  XOR U5568 ( .A(in[292]), .B(n3772), .Z(n4155) );
  XOR U5569 ( .A(in[1525]), .B(n3773), .Z(n4587) );
  XNOR U5570 ( .A(in[1136]), .B(n3774), .Z(n4584) );
  NAND U5571 ( .A(n4587), .B(n4584), .Z(n3775) );
  XNOR U5572 ( .A(n4155), .B(n3775), .Z(out[694]) );
  XNOR U5573 ( .A(in[293]), .B(n3776), .Z(n4158) );
  XOR U5574 ( .A(in[1526]), .B(n3777), .Z(n4591) );
  XNOR U5575 ( .A(in[1137]), .B(n3778), .Z(n4588) );
  NAND U5576 ( .A(n4591), .B(n4588), .Z(n3779) );
  XNOR U5577 ( .A(n4158), .B(n3779), .Z(out[695]) );
  XNOR U5578 ( .A(in[294]), .B(n3780), .Z(n4161) );
  XOR U5579 ( .A(in[1527]), .B(n3781), .Z(n4595) );
  XNOR U5580 ( .A(in[1138]), .B(n3782), .Z(n4592) );
  NAND U5581 ( .A(n4595), .B(n4592), .Z(n3783) );
  XNOR U5582 ( .A(n4161), .B(n3783), .Z(out[696]) );
  XNOR U5583 ( .A(in[295]), .B(n3784), .Z(n4164) );
  XOR U5584 ( .A(in[1528]), .B(n3785), .Z(n4599) );
  XNOR U5585 ( .A(in[1139]), .B(n3786), .Z(n4596) );
  NAND U5586 ( .A(n4599), .B(n4596), .Z(n3787) );
  XNOR U5587 ( .A(n4164), .B(n3787), .Z(out[697]) );
  XNOR U5588 ( .A(in[296]), .B(n3788), .Z(n4167) );
  XOR U5589 ( .A(in[1529]), .B(n3789), .Z(n4603) );
  XNOR U5590 ( .A(in[1140]), .B(n3790), .Z(n4600) );
  NAND U5591 ( .A(n4603), .B(n4600), .Z(n3791) );
  XNOR U5592 ( .A(n4167), .B(n3791), .Z(out[698]) );
  XNOR U5593 ( .A(in[297]), .B(n3792), .Z(n4170) );
  XOR U5594 ( .A(in[1530]), .B(n3793), .Z(n4607) );
  XNOR U5595 ( .A(in[1141]), .B(n3794), .Z(n4604) );
  NAND U5596 ( .A(n4607), .B(n4604), .Z(n3795) );
  XNOR U5597 ( .A(n4170), .B(n3795), .Z(out[699]) );
  ANDN U5598 ( .B(n3797), .A(n3796), .Z(n3798) );
  XNOR U5599 ( .A(n3799), .B(n3798), .Z(out[69]) );
  OR U5600 ( .A(n3831), .B(n3800), .Z(n3801) );
  XNOR U5601 ( .A(n3830), .B(n3801), .Z(out[6]) );
  XNOR U5602 ( .A(in[298]), .B(n3802), .Z(n4173) );
  XNOR U5603 ( .A(in[1531]), .B(n3803), .Z(n4611) );
  XNOR U5604 ( .A(in[1142]), .B(n3804), .Z(n4608) );
  NAND U5605 ( .A(n4611), .B(n4608), .Z(n3805) );
  XNOR U5606 ( .A(n4173), .B(n3805), .Z(out[700]) );
  XNOR U5607 ( .A(in[299]), .B(n3806), .Z(n4176) );
  XNOR U5608 ( .A(in[1532]), .B(n3807), .Z(n4615) );
  XNOR U5609 ( .A(in[1143]), .B(n3808), .Z(n4612) );
  NAND U5610 ( .A(n4615), .B(n4612), .Z(n3809) );
  XNOR U5611 ( .A(n4176), .B(n3809), .Z(out[701]) );
  XNOR U5612 ( .A(in[300]), .B(n3810), .Z(n4183) );
  XNOR U5613 ( .A(in[1533]), .B(n3811), .Z(n4619) );
  XNOR U5614 ( .A(in[1144]), .B(n3812), .Z(n4616) );
  NAND U5615 ( .A(n4619), .B(n4616), .Z(n3813) );
  XNOR U5616 ( .A(n4183), .B(n3813), .Z(out[702]) );
  XNOR U5617 ( .A(in[301]), .B(n3814), .Z(n4186) );
  XOR U5618 ( .A(in[1534]), .B(n3815), .Z(n4623) );
  XNOR U5619 ( .A(in[1145]), .B(n3816), .Z(n4620) );
  NAND U5620 ( .A(n4623), .B(n4620), .Z(n3817) );
  XNOR U5621 ( .A(n4186), .B(n3817), .Z(out[703]) );
  XOR U5622 ( .A(in[376]), .B(n3818), .Z(n4188) );
  NOR U5623 ( .A(n3965), .B(n4343), .Z(n3819) );
  XNOR U5624 ( .A(n4188), .B(n3819), .Z(out[704]) );
  XOR U5625 ( .A(in[377]), .B(n3820), .Z(n4190) );
  NOR U5626 ( .A(n3968), .B(n4347), .Z(n3821) );
  XNOR U5627 ( .A(n4190), .B(n3821), .Z(out[705]) );
  XOR U5628 ( .A(in[378]), .B(n3822), .Z(n4192) );
  NOR U5629 ( .A(n3975), .B(n4351), .Z(n3823) );
  XNOR U5630 ( .A(n4192), .B(n3823), .Z(out[706]) );
  XOR U5631 ( .A(in[379]), .B(n3824), .Z(n4194) );
  NOR U5632 ( .A(n3978), .B(n4355), .Z(n3825) );
  XNOR U5633 ( .A(n4194), .B(n3825), .Z(out[707]) );
  XOR U5634 ( .A(in[380]), .B(n3826), .Z(n4196) );
  NOR U5635 ( .A(n3981), .B(n4367), .Z(n3827) );
  XNOR U5636 ( .A(n4196), .B(n3827), .Z(out[708]) );
  XOR U5637 ( .A(in[381]), .B(n3828), .Z(n4198) );
  NOR U5638 ( .A(n3984), .B(n4371), .Z(n3829) );
  XNOR U5639 ( .A(n4198), .B(n3829), .Z(out[709]) );
  ANDN U5640 ( .B(n3831), .A(n3830), .Z(n3832) );
  XNOR U5641 ( .A(n3833), .B(n3832), .Z(out[70]) );
  XOR U5642 ( .A(in[382]), .B(n3834), .Z(n4200) );
  NOR U5643 ( .A(n3987), .B(n4375), .Z(n3835) );
  XNOR U5644 ( .A(n4200), .B(n3835), .Z(out[710]) );
  XOR U5645 ( .A(in[383]), .B(n3836), .Z(n4202) );
  NOR U5646 ( .A(n3990), .B(n4379), .Z(n3837) );
  XNOR U5647 ( .A(n4202), .B(n3837), .Z(out[711]) );
  XOR U5648 ( .A(in[320]), .B(n3838), .Z(n4208) );
  NOR U5649 ( .A(n3993), .B(n4383), .Z(n3839) );
  XNOR U5650 ( .A(n4208), .B(n3839), .Z(out[712]) );
  XOR U5651 ( .A(in[321]), .B(n3840), .Z(n4210) );
  NOR U5652 ( .A(n3996), .B(n4387), .Z(n3841) );
  XNOR U5653 ( .A(n4210), .B(n3841), .Z(out[713]) );
  XOR U5654 ( .A(in[322]), .B(n3842), .Z(n4212) );
  NOR U5655 ( .A(n3999), .B(n4391), .Z(n3843) );
  XNOR U5656 ( .A(n4212), .B(n3843), .Z(out[714]) );
  XOR U5657 ( .A(in[323]), .B(n3844), .Z(n4214) );
  NOR U5658 ( .A(n4002), .B(n4395), .Z(n3845) );
  XNOR U5659 ( .A(n4214), .B(n3845), .Z(out[715]) );
  XOR U5660 ( .A(in[324]), .B(n3846), .Z(n4216) );
  NOR U5661 ( .A(n4009), .B(n4399), .Z(n3847) );
  XNOR U5662 ( .A(n4216), .B(n3847), .Z(out[716]) );
  XOR U5663 ( .A(in[325]), .B(n3848), .Z(n4218) );
  NOR U5664 ( .A(n4012), .B(n4403), .Z(n3849) );
  XNOR U5665 ( .A(n4218), .B(n3849), .Z(out[717]) );
  XOR U5666 ( .A(in[326]), .B(n3850), .Z(n4220) );
  NOR U5667 ( .A(n4015), .B(n4411), .Z(n3851) );
  XNOR U5668 ( .A(n4220), .B(n3851), .Z(out[718]) );
  XOR U5669 ( .A(in[327]), .B(n3852), .Z(n4222) );
  NOR U5670 ( .A(n4018), .B(n4415), .Z(n3853) );
  XNOR U5671 ( .A(n4222), .B(n3853), .Z(out[719]) );
  ANDN U5672 ( .B(n4077), .A(n4079), .Z(n3854) );
  XNOR U5673 ( .A(n3855), .B(n3854), .Z(out[71]) );
  XOR U5674 ( .A(in[328]), .B(n3856), .Z(n4224) );
  NOR U5675 ( .A(n4021), .B(n4419), .Z(n3857) );
  XNOR U5676 ( .A(n4224), .B(n3857), .Z(out[720]) );
  XOR U5677 ( .A(in[329]), .B(n3858), .Z(n4226) );
  NOR U5678 ( .A(n4024), .B(n4423), .Z(n3859) );
  XNOR U5679 ( .A(n4226), .B(n3859), .Z(out[721]) );
  XOR U5680 ( .A(in[330]), .B(n3860), .Z(n4232) );
  NOR U5681 ( .A(n4027), .B(n4427), .Z(n3861) );
  XNOR U5682 ( .A(n4232), .B(n3861), .Z(out[722]) );
  XOR U5683 ( .A(in[331]), .B(n3862), .Z(n4234) );
  NOR U5684 ( .A(n4030), .B(n4431), .Z(n3863) );
  XNOR U5685 ( .A(n4234), .B(n3863), .Z(out[723]) );
  XOR U5686 ( .A(in[332]), .B(n3864), .Z(n4236) );
  NOR U5687 ( .A(n4033), .B(n4435), .Z(n3865) );
  XNOR U5688 ( .A(n4236), .B(n3865), .Z(out[724]) );
  XOR U5689 ( .A(in[333]), .B(n3866), .Z(n4238) );
  NOR U5690 ( .A(n4036), .B(n4439), .Z(n3867) );
  XNOR U5691 ( .A(n4238), .B(n3867), .Z(out[725]) );
  XOR U5692 ( .A(in[334]), .B(n3868), .Z(n4240) );
  NOR U5693 ( .A(n4043), .B(n4443), .Z(n3869) );
  XNOR U5694 ( .A(n4240), .B(n3869), .Z(out[726]) );
  XOR U5695 ( .A(in[335]), .B(n3870), .Z(n4242) );
  NOR U5696 ( .A(n4046), .B(n4447), .Z(n3871) );
  XNOR U5697 ( .A(n4242), .B(n3871), .Z(out[727]) );
  XOR U5698 ( .A(in[336]), .B(n3872), .Z(n4244) );
  NOR U5699 ( .A(n4049), .B(n4455), .Z(n3873) );
  XNOR U5700 ( .A(n4244), .B(n3873), .Z(out[728]) );
  XOR U5701 ( .A(in[337]), .B(n3874), .Z(n4246) );
  NOR U5702 ( .A(n4052), .B(n4459), .Z(n3875) );
  XNOR U5703 ( .A(n4246), .B(n3875), .Z(out[729]) );
  ANDN U5704 ( .B(n4361), .A(n4363), .Z(n3876) );
  XNOR U5705 ( .A(n3877), .B(n3876), .Z(out[72]) );
  XOR U5706 ( .A(in[338]), .B(n3878), .Z(n4248) );
  NOR U5707 ( .A(n4055), .B(n4463), .Z(n3879) );
  XNOR U5708 ( .A(n4248), .B(n3879), .Z(out[730]) );
  XOR U5709 ( .A(in[339]), .B(n3880), .Z(n4250) );
  NOR U5710 ( .A(n4058), .B(n4467), .Z(n3881) );
  XNOR U5711 ( .A(n4250), .B(n3881), .Z(out[731]) );
  XOR U5712 ( .A(in[340]), .B(n3882), .Z(n4256) );
  NOR U5713 ( .A(n4061), .B(n4471), .Z(n3883) );
  XNOR U5714 ( .A(n4256), .B(n3883), .Z(out[732]) );
  XOR U5715 ( .A(in[341]), .B(n3884), .Z(n4258) );
  NOR U5716 ( .A(n4064), .B(n4475), .Z(n3885) );
  XNOR U5717 ( .A(n4258), .B(n3885), .Z(out[733]) );
  XOR U5718 ( .A(in[342]), .B(n3886), .Z(n4260) );
  NOR U5719 ( .A(n4067), .B(n4479), .Z(n3887) );
  XNOR U5720 ( .A(n4260), .B(n3887), .Z(out[734]) );
  XOR U5721 ( .A(in[343]), .B(n3888), .Z(n4262) );
  NOR U5722 ( .A(n4070), .B(n4483), .Z(n3889) );
  XNOR U5723 ( .A(n4262), .B(n3889), .Z(out[735]) );
  XOR U5724 ( .A(in[344]), .B(n3890), .Z(n4264) );
  NOR U5725 ( .A(n4081), .B(n4487), .Z(n3891) );
  XNOR U5726 ( .A(n4264), .B(n3891), .Z(out[736]) );
  XOR U5727 ( .A(in[345]), .B(n3892), .Z(n4266) );
  NOR U5728 ( .A(n4084), .B(n4491), .Z(n3893) );
  XNOR U5729 ( .A(n4266), .B(n3893), .Z(out[737]) );
  XOR U5730 ( .A(in[346]), .B(n3894), .Z(n4268) );
  NOR U5731 ( .A(n4087), .B(n4499), .Z(n3895) );
  XNOR U5732 ( .A(n4268), .B(n3895), .Z(out[738]) );
  XOR U5733 ( .A(in[347]), .B(n3896), .Z(n4270) );
  NOR U5734 ( .A(n4090), .B(n4503), .Z(n3897) );
  XNOR U5735 ( .A(n4270), .B(n3897), .Z(out[739]) );
  ANDN U5736 ( .B(n4805), .A(n4807), .Z(n3898) );
  XNOR U5737 ( .A(n3899), .B(n3898), .Z(out[73]) );
  XOR U5738 ( .A(in[348]), .B(n3900), .Z(n4272) );
  NOR U5739 ( .A(n4093), .B(n4507), .Z(n3901) );
  XNOR U5740 ( .A(n4272), .B(n3901), .Z(out[740]) );
  XOR U5741 ( .A(in[349]), .B(n3902), .Z(n4274) );
  NOR U5742 ( .A(n4096), .B(n4511), .Z(n3903) );
  XNOR U5743 ( .A(n4274), .B(n3903), .Z(out[741]) );
  XOR U5744 ( .A(in[350]), .B(n3904), .Z(n4280) );
  NOR U5745 ( .A(n4099), .B(n4515), .Z(n3905) );
  XNOR U5746 ( .A(n4280), .B(n3905), .Z(out[742]) );
  XOR U5747 ( .A(in[351]), .B(n3906), .Z(n4282) );
  NOR U5748 ( .A(n4102), .B(n4519), .Z(n3907) );
  XNOR U5749 ( .A(n4282), .B(n3907), .Z(out[743]) );
  XOR U5750 ( .A(in[352]), .B(n3908), .Z(n4284) );
  NOR U5751 ( .A(n4105), .B(n4523), .Z(n3909) );
  XNOR U5752 ( .A(n4284), .B(n3909), .Z(out[744]) );
  XOR U5753 ( .A(in[353]), .B(n3910), .Z(n4286) );
  NOR U5754 ( .A(n4108), .B(n4527), .Z(n3911) );
  XNOR U5755 ( .A(n4286), .B(n3911), .Z(out[745]) );
  XOR U5756 ( .A(in[354]), .B(n3912), .Z(n4288) );
  NOR U5757 ( .A(n4115), .B(n4531), .Z(n3913) );
  XNOR U5758 ( .A(n4288), .B(n3913), .Z(out[746]) );
  XOR U5759 ( .A(in[355]), .B(n3914), .Z(n4290) );
  NOR U5760 ( .A(n4118), .B(n4535), .Z(n3915) );
  XNOR U5761 ( .A(n4290), .B(n3915), .Z(out[747]) );
  XOR U5762 ( .A(in[356]), .B(n3916), .Z(n4292) );
  NOR U5763 ( .A(n4121), .B(n4543), .Z(n3917) );
  XNOR U5764 ( .A(n4292), .B(n3917), .Z(out[748]) );
  XOR U5765 ( .A(in[357]), .B(n3918), .Z(n4294) );
  NOR U5766 ( .A(n4124), .B(n4547), .Z(n3919) );
  XNOR U5767 ( .A(n4294), .B(n3919), .Z(out[749]) );
  NOR U5768 ( .A(n3921), .B(n3920), .Z(n3922) );
  XNOR U5769 ( .A(n3923), .B(n3922), .Z(out[74]) );
  XOR U5770 ( .A(in[358]), .B(n3924), .Z(n4296) );
  NOR U5771 ( .A(n4127), .B(n4551), .Z(n3925) );
  XNOR U5772 ( .A(n4296), .B(n3925), .Z(out[750]) );
  XOR U5773 ( .A(in[359]), .B(n3926), .Z(n4298) );
  NOR U5774 ( .A(n4130), .B(n4555), .Z(n3927) );
  XNOR U5775 ( .A(n4298), .B(n3927), .Z(out[751]) );
  XOR U5776 ( .A(in[360]), .B(n3928), .Z(n4304) );
  NOR U5777 ( .A(n4133), .B(n4559), .Z(n3929) );
  XNOR U5778 ( .A(n4304), .B(n3929), .Z(out[752]) );
  XOR U5779 ( .A(in[361]), .B(n3930), .Z(n4306) );
  NOR U5780 ( .A(n4136), .B(n4563), .Z(n3931) );
  XNOR U5781 ( .A(n4306), .B(n3931), .Z(out[753]) );
  XOR U5782 ( .A(in[362]), .B(n3932), .Z(n4308) );
  NOR U5783 ( .A(n4139), .B(n4567), .Z(n3933) );
  XNOR U5784 ( .A(n4308), .B(n3933), .Z(out[754]) );
  XOR U5785 ( .A(in[363]), .B(n3934), .Z(n4310) );
  NOR U5786 ( .A(n4142), .B(n4571), .Z(n3935) );
  XNOR U5787 ( .A(n4310), .B(n3935), .Z(out[755]) );
  XOR U5788 ( .A(in[364]), .B(n3936), .Z(n4312) );
  NOR U5789 ( .A(n4149), .B(n4575), .Z(n3937) );
  XNOR U5790 ( .A(n4312), .B(n3937), .Z(out[756]) );
  XOR U5791 ( .A(in[365]), .B(n3938), .Z(n4314) );
  NOR U5792 ( .A(n4152), .B(n4579), .Z(n3939) );
  XNOR U5793 ( .A(n4314), .B(n3939), .Z(out[757]) );
  XOR U5794 ( .A(in[366]), .B(n3940), .Z(n4316) );
  NOR U5795 ( .A(n4155), .B(n4587), .Z(n3941) );
  XNOR U5796 ( .A(n4316), .B(n3941), .Z(out[758]) );
  XOR U5797 ( .A(in[367]), .B(n3942), .Z(n4318) );
  NOR U5798 ( .A(n4158), .B(n4591), .Z(n3943) );
  XNOR U5799 ( .A(n4318), .B(n3943), .Z(out[759]) );
  NOR U5800 ( .A(n3945), .B(n3944), .Z(n3946) );
  XNOR U5801 ( .A(n3947), .B(n3946), .Z(out[75]) );
  XOR U5802 ( .A(in[368]), .B(n3948), .Z(n4320) );
  NOR U5803 ( .A(n4161), .B(n4595), .Z(n3949) );
  XNOR U5804 ( .A(n4320), .B(n3949), .Z(out[760]) );
  XOR U5805 ( .A(in[369]), .B(n3950), .Z(n4322) );
  NOR U5806 ( .A(n4164), .B(n4599), .Z(n3951) );
  XNOR U5807 ( .A(n4322), .B(n3951), .Z(out[761]) );
  XOR U5808 ( .A(in[370]), .B(n3952), .Z(n4328) );
  NOR U5809 ( .A(n4167), .B(n4603), .Z(n3953) );
  XNOR U5810 ( .A(n4328), .B(n3953), .Z(out[762]) );
  XOR U5811 ( .A(in[371]), .B(n3954), .Z(n4330) );
  NOR U5812 ( .A(n4170), .B(n4607), .Z(n3955) );
  XNOR U5813 ( .A(n4330), .B(n3955), .Z(out[763]) );
  XOR U5814 ( .A(in[372]), .B(n3956), .Z(n4332) );
  NOR U5815 ( .A(n4173), .B(n4611), .Z(n3957) );
  XNOR U5816 ( .A(n4332), .B(n3957), .Z(out[764]) );
  XOR U5817 ( .A(in[373]), .B(n3958), .Z(n4334) );
  NOR U5818 ( .A(n4176), .B(n4615), .Z(n3959) );
  XNOR U5819 ( .A(n4334), .B(n3959), .Z(out[765]) );
  XOR U5820 ( .A(in[374]), .B(n3960), .Z(n4336) );
  NOR U5821 ( .A(n4183), .B(n4619), .Z(n3961) );
  XNOR U5822 ( .A(n4336), .B(n3961), .Z(out[766]) );
  XOR U5823 ( .A(in[375]), .B(n3962), .Z(n4338) );
  NOR U5824 ( .A(n4186), .B(n4623), .Z(n3963) );
  XNOR U5825 ( .A(n4338), .B(n3963), .Z(out[767]) );
  XNOR U5826 ( .A(in[743]), .B(n3964), .Z(n4341) );
  NAND U5827 ( .A(n4188), .B(n3965), .Z(n3966) );
  XNOR U5828 ( .A(n4341), .B(n3966), .Z(out[768]) );
  XNOR U5829 ( .A(in[744]), .B(n3967), .Z(n4345) );
  NAND U5830 ( .A(n4190), .B(n3968), .Z(n3969) );
  XNOR U5831 ( .A(n4345), .B(n3969), .Z(out[769]) );
  NOR U5832 ( .A(n3971), .B(n3970), .Z(n3972) );
  XNOR U5833 ( .A(n3973), .B(n3972), .Z(out[76]) );
  XNOR U5834 ( .A(in[745]), .B(n3974), .Z(n4349) );
  NAND U5835 ( .A(n4192), .B(n3975), .Z(n3976) );
  XNOR U5836 ( .A(n4349), .B(n3976), .Z(out[770]) );
  XNOR U5837 ( .A(in[746]), .B(n3977), .Z(n4353) );
  NAND U5838 ( .A(n4194), .B(n3978), .Z(n3979) );
  XNOR U5839 ( .A(n4353), .B(n3979), .Z(out[771]) );
  XNOR U5840 ( .A(in[747]), .B(n3980), .Z(n4365) );
  NAND U5841 ( .A(n4196), .B(n3981), .Z(n3982) );
  XNOR U5842 ( .A(n4365), .B(n3982), .Z(out[772]) );
  XNOR U5843 ( .A(in[748]), .B(n3983), .Z(n4369) );
  NAND U5844 ( .A(n4198), .B(n3984), .Z(n3985) );
  XNOR U5845 ( .A(n4369), .B(n3985), .Z(out[773]) );
  XNOR U5846 ( .A(in[749]), .B(n3986), .Z(n4373) );
  NAND U5847 ( .A(n4200), .B(n3987), .Z(n3988) );
  XNOR U5848 ( .A(n4373), .B(n3988), .Z(out[774]) );
  XNOR U5849 ( .A(in[750]), .B(n3989), .Z(n4377) );
  NAND U5850 ( .A(n4202), .B(n3990), .Z(n3991) );
  XNOR U5851 ( .A(n4377), .B(n3991), .Z(out[775]) );
  XNOR U5852 ( .A(in[751]), .B(n3992), .Z(n4381) );
  NAND U5853 ( .A(n4208), .B(n3993), .Z(n3994) );
  XNOR U5854 ( .A(n4381), .B(n3994), .Z(out[776]) );
  XNOR U5855 ( .A(in[752]), .B(n3995), .Z(n4385) );
  NAND U5856 ( .A(n4210), .B(n3996), .Z(n3997) );
  XNOR U5857 ( .A(n4385), .B(n3997), .Z(out[777]) );
  XNOR U5858 ( .A(in[753]), .B(n3998), .Z(n4389) );
  NAND U5859 ( .A(n4212), .B(n3999), .Z(n4000) );
  XNOR U5860 ( .A(n4389), .B(n4000), .Z(out[778]) );
  XNOR U5861 ( .A(in[754]), .B(n4001), .Z(n4393) );
  NAND U5862 ( .A(n4214), .B(n4002), .Z(n4003) );
  XNOR U5863 ( .A(n4393), .B(n4003), .Z(out[779]) );
  NOR U5864 ( .A(n4005), .B(n4004), .Z(n4006) );
  XNOR U5865 ( .A(n4007), .B(n4006), .Z(out[77]) );
  XNOR U5866 ( .A(in[755]), .B(n4008), .Z(n4397) );
  NAND U5867 ( .A(n4216), .B(n4009), .Z(n4010) );
  XNOR U5868 ( .A(n4397), .B(n4010), .Z(out[780]) );
  XNOR U5869 ( .A(in[756]), .B(n4011), .Z(n4401) );
  NAND U5870 ( .A(n4218), .B(n4012), .Z(n4013) );
  XNOR U5871 ( .A(n4401), .B(n4013), .Z(out[781]) );
  XNOR U5872 ( .A(in[757]), .B(n4014), .Z(n4409) );
  NAND U5873 ( .A(n4220), .B(n4015), .Z(n4016) );
  XNOR U5874 ( .A(n4409), .B(n4016), .Z(out[782]) );
  XNOR U5875 ( .A(in[758]), .B(n4017), .Z(n4413) );
  NAND U5876 ( .A(n4222), .B(n4018), .Z(n4019) );
  XNOR U5877 ( .A(n4413), .B(n4019), .Z(out[783]) );
  XNOR U5878 ( .A(in[759]), .B(n4020), .Z(n4417) );
  NAND U5879 ( .A(n4224), .B(n4021), .Z(n4022) );
  XNOR U5880 ( .A(n4417), .B(n4022), .Z(out[784]) );
  XNOR U5881 ( .A(in[760]), .B(n4023), .Z(n4421) );
  NAND U5882 ( .A(n4226), .B(n4024), .Z(n4025) );
  XNOR U5883 ( .A(n4421), .B(n4025), .Z(out[785]) );
  XNOR U5884 ( .A(in[761]), .B(n4026), .Z(n4425) );
  NAND U5885 ( .A(n4232), .B(n4027), .Z(n4028) );
  XNOR U5886 ( .A(n4425), .B(n4028), .Z(out[786]) );
  XNOR U5887 ( .A(in[762]), .B(n4029), .Z(n4429) );
  NAND U5888 ( .A(n4234), .B(n4030), .Z(n4031) );
  XNOR U5889 ( .A(n4429), .B(n4031), .Z(out[787]) );
  XNOR U5890 ( .A(in[763]), .B(n4032), .Z(n4433) );
  NAND U5891 ( .A(n4236), .B(n4033), .Z(n4034) );
  XNOR U5892 ( .A(n4433), .B(n4034), .Z(out[788]) );
  XNOR U5893 ( .A(in[764]), .B(n4035), .Z(n4437) );
  NAND U5894 ( .A(n4238), .B(n4036), .Z(n4037) );
  XNOR U5895 ( .A(n4437), .B(n4037), .Z(out[789]) );
  NOR U5896 ( .A(n4039), .B(n4038), .Z(n4040) );
  XNOR U5897 ( .A(n4041), .B(n4040), .Z(out[78]) );
  XNOR U5898 ( .A(in[765]), .B(n4042), .Z(n4441) );
  NAND U5899 ( .A(n4240), .B(n4043), .Z(n4044) );
  XNOR U5900 ( .A(n4441), .B(n4044), .Z(out[790]) );
  XNOR U5901 ( .A(in[766]), .B(n4045), .Z(n4445) );
  NAND U5902 ( .A(n4242), .B(n4046), .Z(n4047) );
  XNOR U5903 ( .A(n4445), .B(n4047), .Z(out[791]) );
  XNOR U5904 ( .A(in[767]), .B(n4048), .Z(n4453) );
  NAND U5905 ( .A(n4244), .B(n4049), .Z(n4050) );
  XNOR U5906 ( .A(n4453), .B(n4050), .Z(out[792]) );
  XNOR U5907 ( .A(in[704]), .B(n4051), .Z(n4457) );
  NAND U5908 ( .A(n4246), .B(n4052), .Z(n4053) );
  XNOR U5909 ( .A(n4457), .B(n4053), .Z(out[793]) );
  XNOR U5910 ( .A(in[705]), .B(n4054), .Z(n4461) );
  NAND U5911 ( .A(n4248), .B(n4055), .Z(n4056) );
  XNOR U5912 ( .A(n4461), .B(n4056), .Z(out[794]) );
  XNOR U5913 ( .A(in[706]), .B(n4057), .Z(n4465) );
  NAND U5914 ( .A(n4250), .B(n4058), .Z(n4059) );
  XNOR U5915 ( .A(n4465), .B(n4059), .Z(out[795]) );
  XNOR U5916 ( .A(in[707]), .B(n4060), .Z(n4469) );
  NAND U5917 ( .A(n4256), .B(n4061), .Z(n4062) );
  XNOR U5918 ( .A(n4469), .B(n4062), .Z(out[796]) );
  XNOR U5919 ( .A(in[708]), .B(n4063), .Z(n4473) );
  NAND U5920 ( .A(n4258), .B(n4064), .Z(n4065) );
  XNOR U5921 ( .A(n4473), .B(n4065), .Z(out[797]) );
  XNOR U5922 ( .A(in[709]), .B(n4066), .Z(n4477) );
  NAND U5923 ( .A(n4260), .B(n4067), .Z(n4068) );
  XNOR U5924 ( .A(n4477), .B(n4068), .Z(out[798]) );
  XNOR U5925 ( .A(in[710]), .B(n4069), .Z(n4481) );
  NAND U5926 ( .A(n4262), .B(n4070), .Z(n4071) );
  XNOR U5927 ( .A(n4481), .B(n4071), .Z(out[799]) );
  NOR U5928 ( .A(n4073), .B(n4072), .Z(n4074) );
  XNOR U5929 ( .A(n4075), .B(n4074), .Z(out[79]) );
  OR U5930 ( .A(n4077), .B(n4076), .Z(n4078) );
  XNOR U5931 ( .A(n4079), .B(n4078), .Z(out[7]) );
  XNOR U5932 ( .A(in[711]), .B(n4080), .Z(n4485) );
  NAND U5933 ( .A(n4264), .B(n4081), .Z(n4082) );
  XNOR U5934 ( .A(n4485), .B(n4082), .Z(out[800]) );
  XNOR U5935 ( .A(in[712]), .B(n4083), .Z(n4489) );
  NAND U5936 ( .A(n4266), .B(n4084), .Z(n4085) );
  XNOR U5937 ( .A(n4489), .B(n4085), .Z(out[801]) );
  XNOR U5938 ( .A(in[713]), .B(n4086), .Z(n4497) );
  NAND U5939 ( .A(n4268), .B(n4087), .Z(n4088) );
  XNOR U5940 ( .A(n4497), .B(n4088), .Z(out[802]) );
  XNOR U5941 ( .A(in[714]), .B(n4089), .Z(n4501) );
  NAND U5942 ( .A(n4270), .B(n4090), .Z(n4091) );
  XNOR U5943 ( .A(n4501), .B(n4091), .Z(out[803]) );
  XNOR U5944 ( .A(in[715]), .B(n4092), .Z(n4505) );
  NAND U5945 ( .A(n4272), .B(n4093), .Z(n4094) );
  XNOR U5946 ( .A(n4505), .B(n4094), .Z(out[804]) );
  XOR U5947 ( .A(n4095), .B(in[716]), .Z(n4509) );
  NAND U5948 ( .A(n4274), .B(n4096), .Z(n4097) );
  XNOR U5949 ( .A(n4509), .B(n4097), .Z(out[805]) );
  XOR U5950 ( .A(n4098), .B(in[717]), .Z(n4513) );
  NAND U5951 ( .A(n4280), .B(n4099), .Z(n4100) );
  XNOR U5952 ( .A(n4513), .B(n4100), .Z(out[806]) );
  XOR U5953 ( .A(n4101), .B(in[718]), .Z(n4517) );
  NAND U5954 ( .A(n4282), .B(n4102), .Z(n4103) );
  XNOR U5955 ( .A(n4517), .B(n4103), .Z(out[807]) );
  XOR U5956 ( .A(n4104), .B(in[719]), .Z(n4521) );
  NAND U5957 ( .A(n4284), .B(n4105), .Z(n4106) );
  XNOR U5958 ( .A(n4521), .B(n4106), .Z(out[808]) );
  XOR U5959 ( .A(n4107), .B(in[720]), .Z(n4525) );
  NAND U5960 ( .A(n4286), .B(n4108), .Z(n4109) );
  XNOR U5961 ( .A(n4525), .B(n4109), .Z(out[809]) );
  NOR U5962 ( .A(n4111), .B(n4110), .Z(n4112) );
  XNOR U5963 ( .A(n4113), .B(n4112), .Z(out[80]) );
  XOR U5964 ( .A(n4114), .B(in[721]), .Z(n4529) );
  NAND U5965 ( .A(n4288), .B(n4115), .Z(n4116) );
  XNOR U5966 ( .A(n4529), .B(n4116), .Z(out[810]) );
  XOR U5967 ( .A(n4117), .B(in[722]), .Z(n4533) );
  NAND U5968 ( .A(n4290), .B(n4118), .Z(n4119) );
  XNOR U5969 ( .A(n4533), .B(n4119), .Z(out[811]) );
  XOR U5970 ( .A(n4120), .B(in[723]), .Z(n4541) );
  NAND U5971 ( .A(n4292), .B(n4121), .Z(n4122) );
  XNOR U5972 ( .A(n4541), .B(n4122), .Z(out[812]) );
  XOR U5973 ( .A(in[724]), .B(n4123), .Z(n4545) );
  NAND U5974 ( .A(n4294), .B(n4124), .Z(n4125) );
  XNOR U5975 ( .A(n4545), .B(n4125), .Z(out[813]) );
  XOR U5976 ( .A(in[725]), .B(n4126), .Z(n4549) );
  NAND U5977 ( .A(n4296), .B(n4127), .Z(n4128) );
  XNOR U5978 ( .A(n4549), .B(n4128), .Z(out[814]) );
  XOR U5979 ( .A(in[726]), .B(n4129), .Z(n4553) );
  NAND U5980 ( .A(n4298), .B(n4130), .Z(n4131) );
  XNOR U5981 ( .A(n4553), .B(n4131), .Z(out[815]) );
  XOR U5982 ( .A(in[727]), .B(n4132), .Z(n4557) );
  NAND U5983 ( .A(n4304), .B(n4133), .Z(n4134) );
  XNOR U5984 ( .A(n4557), .B(n4134), .Z(out[816]) );
  XOR U5985 ( .A(in[728]), .B(n4135), .Z(n4561) );
  NAND U5986 ( .A(n4306), .B(n4136), .Z(n4137) );
  XNOR U5987 ( .A(n4561), .B(n4137), .Z(out[817]) );
  XOR U5988 ( .A(in[729]), .B(n4138), .Z(n4565) );
  NAND U5989 ( .A(n4308), .B(n4139), .Z(n4140) );
  XNOR U5990 ( .A(n4565), .B(n4140), .Z(out[818]) );
  XOR U5991 ( .A(in[730]), .B(n4141), .Z(n4569) );
  NAND U5992 ( .A(n4310), .B(n4142), .Z(n4143) );
  XNOR U5993 ( .A(n4569), .B(n4143), .Z(out[819]) );
  NOR U5994 ( .A(n4145), .B(n4144), .Z(n4146) );
  XNOR U5995 ( .A(n4147), .B(n4146), .Z(out[81]) );
  XOR U5996 ( .A(in[731]), .B(n4148), .Z(n4573) );
  NAND U5997 ( .A(n4312), .B(n4149), .Z(n4150) );
  XNOR U5998 ( .A(n4573), .B(n4150), .Z(out[820]) );
  XOR U5999 ( .A(in[732]), .B(n4151), .Z(n4577) );
  NAND U6000 ( .A(n4314), .B(n4152), .Z(n4153) );
  XNOR U6001 ( .A(n4577), .B(n4153), .Z(out[821]) );
  XOR U6002 ( .A(in[733]), .B(n4154), .Z(n4585) );
  NAND U6003 ( .A(n4316), .B(n4155), .Z(n4156) );
  XNOR U6004 ( .A(n4585), .B(n4156), .Z(out[822]) );
  XOR U6005 ( .A(in[734]), .B(n4157), .Z(n4589) );
  NAND U6006 ( .A(n4318), .B(n4158), .Z(n4159) );
  XNOR U6007 ( .A(n4589), .B(n4159), .Z(out[823]) );
  XOR U6008 ( .A(in[735]), .B(n4160), .Z(n4593) );
  NAND U6009 ( .A(n4320), .B(n4161), .Z(n4162) );
  XNOR U6010 ( .A(n4593), .B(n4162), .Z(out[824]) );
  XOR U6011 ( .A(in[736]), .B(n4163), .Z(n4597) );
  NAND U6012 ( .A(n4322), .B(n4164), .Z(n4165) );
  XNOR U6013 ( .A(n4597), .B(n4165), .Z(out[825]) );
  XOR U6014 ( .A(in[737]), .B(n4166), .Z(n4601) );
  NAND U6015 ( .A(n4328), .B(n4167), .Z(n4168) );
  XNOR U6016 ( .A(n4601), .B(n4168), .Z(out[826]) );
  XOR U6017 ( .A(in[738]), .B(n4169), .Z(n4605) );
  NAND U6018 ( .A(n4330), .B(n4170), .Z(n4171) );
  XNOR U6019 ( .A(n4605), .B(n4171), .Z(out[827]) );
  XOR U6020 ( .A(in[739]), .B(n4172), .Z(n4609) );
  NAND U6021 ( .A(n4332), .B(n4173), .Z(n4174) );
  XNOR U6022 ( .A(n4609), .B(n4174), .Z(out[828]) );
  XNOR U6023 ( .A(in[740]), .B(n4175), .Z(n4613) );
  NAND U6024 ( .A(n4334), .B(n4176), .Z(n4177) );
  XNOR U6025 ( .A(n4613), .B(n4177), .Z(out[829]) );
  NOR U6026 ( .A(n4179), .B(n4178), .Z(n4180) );
  XNOR U6027 ( .A(n4181), .B(n4180), .Z(out[82]) );
  XNOR U6028 ( .A(in[741]), .B(n4182), .Z(n4617) );
  NAND U6029 ( .A(n4336), .B(n4183), .Z(n4184) );
  XNOR U6030 ( .A(n4617), .B(n4184), .Z(out[830]) );
  XNOR U6031 ( .A(in[742]), .B(n4185), .Z(n4621) );
  NAND U6032 ( .A(n4338), .B(n4186), .Z(n4187) );
  XNOR U6033 ( .A(n4621), .B(n4187), .Z(out[831]) );
  OR U6034 ( .A(n4341), .B(n4188), .Z(n4189) );
  XNOR U6035 ( .A(n4340), .B(n4189), .Z(out[832]) );
  OR U6036 ( .A(n4345), .B(n4190), .Z(n4191) );
  XNOR U6037 ( .A(n4344), .B(n4191), .Z(out[833]) );
  OR U6038 ( .A(n4349), .B(n4192), .Z(n4193) );
  XNOR U6039 ( .A(n4348), .B(n4193), .Z(out[834]) );
  OR U6040 ( .A(n4353), .B(n4194), .Z(n4195) );
  XNOR U6041 ( .A(n4352), .B(n4195), .Z(out[835]) );
  OR U6042 ( .A(n4365), .B(n4196), .Z(n4197) );
  XNOR U6043 ( .A(n4364), .B(n4197), .Z(out[836]) );
  OR U6044 ( .A(n4369), .B(n4198), .Z(n4199) );
  XNOR U6045 ( .A(n4368), .B(n4199), .Z(out[837]) );
  OR U6046 ( .A(n4373), .B(n4200), .Z(n4201) );
  XNOR U6047 ( .A(n4372), .B(n4201), .Z(out[838]) );
  OR U6048 ( .A(n4377), .B(n4202), .Z(n4203) );
  XNOR U6049 ( .A(n4376), .B(n4203), .Z(out[839]) );
  NOR U6050 ( .A(n4205), .B(n4204), .Z(n4206) );
  XNOR U6051 ( .A(n4207), .B(n4206), .Z(out[83]) );
  OR U6052 ( .A(n4381), .B(n4208), .Z(n4209) );
  XNOR U6053 ( .A(n4380), .B(n4209), .Z(out[840]) );
  OR U6054 ( .A(n4385), .B(n4210), .Z(n4211) );
  XNOR U6055 ( .A(n4384), .B(n4211), .Z(out[841]) );
  OR U6056 ( .A(n4389), .B(n4212), .Z(n4213) );
  XNOR U6057 ( .A(n4388), .B(n4213), .Z(out[842]) );
  OR U6058 ( .A(n4393), .B(n4214), .Z(n4215) );
  XNOR U6059 ( .A(n4392), .B(n4215), .Z(out[843]) );
  OR U6060 ( .A(n4397), .B(n4216), .Z(n4217) );
  XNOR U6061 ( .A(n4396), .B(n4217), .Z(out[844]) );
  OR U6062 ( .A(n4401), .B(n4218), .Z(n4219) );
  XNOR U6063 ( .A(n4400), .B(n4219), .Z(out[845]) );
  OR U6064 ( .A(n4409), .B(n4220), .Z(n4221) );
  XNOR U6065 ( .A(n4408), .B(n4221), .Z(out[846]) );
  OR U6066 ( .A(n4413), .B(n4222), .Z(n4223) );
  XNOR U6067 ( .A(n4412), .B(n4223), .Z(out[847]) );
  OR U6068 ( .A(n4417), .B(n4224), .Z(n4225) );
  XNOR U6069 ( .A(n4416), .B(n4225), .Z(out[848]) );
  OR U6070 ( .A(n4421), .B(n4226), .Z(n4227) );
  XNOR U6071 ( .A(n4420), .B(n4227), .Z(out[849]) );
  NOR U6072 ( .A(n4229), .B(n4228), .Z(n4230) );
  XNOR U6073 ( .A(n4231), .B(n4230), .Z(out[84]) );
  OR U6074 ( .A(n4425), .B(n4232), .Z(n4233) );
  XNOR U6075 ( .A(n4424), .B(n4233), .Z(out[850]) );
  OR U6076 ( .A(n4429), .B(n4234), .Z(n4235) );
  XNOR U6077 ( .A(n4428), .B(n4235), .Z(out[851]) );
  OR U6078 ( .A(n4433), .B(n4236), .Z(n4237) );
  XNOR U6079 ( .A(n4432), .B(n4237), .Z(out[852]) );
  OR U6080 ( .A(n4437), .B(n4238), .Z(n4239) );
  XNOR U6081 ( .A(n4436), .B(n4239), .Z(out[853]) );
  OR U6082 ( .A(n4441), .B(n4240), .Z(n4241) );
  XNOR U6083 ( .A(n4440), .B(n4241), .Z(out[854]) );
  OR U6084 ( .A(n4445), .B(n4242), .Z(n4243) );
  XNOR U6085 ( .A(n4444), .B(n4243), .Z(out[855]) );
  OR U6086 ( .A(n4453), .B(n4244), .Z(n4245) );
  XNOR U6087 ( .A(n4452), .B(n4245), .Z(out[856]) );
  OR U6088 ( .A(n4457), .B(n4246), .Z(n4247) );
  XNOR U6089 ( .A(n4456), .B(n4247), .Z(out[857]) );
  OR U6090 ( .A(n4461), .B(n4248), .Z(n4249) );
  XNOR U6091 ( .A(n4460), .B(n4249), .Z(out[858]) );
  OR U6092 ( .A(n4465), .B(n4250), .Z(n4251) );
  XNOR U6093 ( .A(n4464), .B(n4251), .Z(out[859]) );
  NOR U6094 ( .A(n4253), .B(n4252), .Z(n4254) );
  XNOR U6095 ( .A(n4255), .B(n4254), .Z(out[85]) );
  OR U6096 ( .A(n4469), .B(n4256), .Z(n4257) );
  XNOR U6097 ( .A(n4468), .B(n4257), .Z(out[860]) );
  OR U6098 ( .A(n4473), .B(n4258), .Z(n4259) );
  XNOR U6099 ( .A(n4472), .B(n4259), .Z(out[861]) );
  OR U6100 ( .A(n4477), .B(n4260), .Z(n4261) );
  XNOR U6101 ( .A(n4476), .B(n4261), .Z(out[862]) );
  OR U6102 ( .A(n4481), .B(n4262), .Z(n4263) );
  XNOR U6103 ( .A(n4480), .B(n4263), .Z(out[863]) );
  OR U6104 ( .A(n4485), .B(n4264), .Z(n4265) );
  XNOR U6105 ( .A(n4484), .B(n4265), .Z(out[864]) );
  OR U6106 ( .A(n4489), .B(n4266), .Z(n4267) );
  XNOR U6107 ( .A(n4488), .B(n4267), .Z(out[865]) );
  OR U6108 ( .A(n4497), .B(n4268), .Z(n4269) );
  XNOR U6109 ( .A(n4496), .B(n4269), .Z(out[866]) );
  OR U6110 ( .A(n4501), .B(n4270), .Z(n4271) );
  XNOR U6111 ( .A(n4500), .B(n4271), .Z(out[867]) );
  OR U6112 ( .A(n4505), .B(n4272), .Z(n4273) );
  XNOR U6113 ( .A(n4504), .B(n4273), .Z(out[868]) );
  OR U6114 ( .A(n4509), .B(n4274), .Z(n4275) );
  XNOR U6115 ( .A(n4508), .B(n4275), .Z(out[869]) );
  NOR U6116 ( .A(n4277), .B(n4276), .Z(n4278) );
  XNOR U6117 ( .A(n4279), .B(n4278), .Z(out[86]) );
  OR U6118 ( .A(n4513), .B(n4280), .Z(n4281) );
  XNOR U6119 ( .A(n4512), .B(n4281), .Z(out[870]) );
  OR U6120 ( .A(n4517), .B(n4282), .Z(n4283) );
  XNOR U6121 ( .A(n4516), .B(n4283), .Z(out[871]) );
  OR U6122 ( .A(n4521), .B(n4284), .Z(n4285) );
  XNOR U6123 ( .A(n4520), .B(n4285), .Z(out[872]) );
  OR U6124 ( .A(n4525), .B(n4286), .Z(n4287) );
  XNOR U6125 ( .A(n4524), .B(n4287), .Z(out[873]) );
  OR U6126 ( .A(n4529), .B(n4288), .Z(n4289) );
  XNOR U6127 ( .A(n4528), .B(n4289), .Z(out[874]) );
  OR U6128 ( .A(n4533), .B(n4290), .Z(n4291) );
  XNOR U6129 ( .A(n4532), .B(n4291), .Z(out[875]) );
  OR U6130 ( .A(n4541), .B(n4292), .Z(n4293) );
  XNOR U6131 ( .A(n4540), .B(n4293), .Z(out[876]) );
  OR U6132 ( .A(n4545), .B(n4294), .Z(n4295) );
  XNOR U6133 ( .A(n4544), .B(n4295), .Z(out[877]) );
  OR U6134 ( .A(n4549), .B(n4296), .Z(n4297) );
  XNOR U6135 ( .A(n4548), .B(n4297), .Z(out[878]) );
  OR U6136 ( .A(n4553), .B(n4298), .Z(n4299) );
  XNOR U6137 ( .A(n4552), .B(n4299), .Z(out[879]) );
  NOR U6138 ( .A(n4301), .B(n4300), .Z(n4302) );
  XNOR U6139 ( .A(n4303), .B(n4302), .Z(out[87]) );
  OR U6140 ( .A(n4557), .B(n4304), .Z(n4305) );
  XNOR U6141 ( .A(n4556), .B(n4305), .Z(out[880]) );
  OR U6142 ( .A(n4561), .B(n4306), .Z(n4307) );
  XNOR U6143 ( .A(n4560), .B(n4307), .Z(out[881]) );
  OR U6144 ( .A(n4565), .B(n4308), .Z(n4309) );
  XNOR U6145 ( .A(n4564), .B(n4309), .Z(out[882]) );
  OR U6146 ( .A(n4569), .B(n4310), .Z(n4311) );
  XNOR U6147 ( .A(n4568), .B(n4311), .Z(out[883]) );
  OR U6148 ( .A(n4573), .B(n4312), .Z(n4313) );
  XNOR U6149 ( .A(n4572), .B(n4313), .Z(out[884]) );
  OR U6150 ( .A(n4577), .B(n4314), .Z(n4315) );
  XNOR U6151 ( .A(n4576), .B(n4315), .Z(out[885]) );
  OR U6152 ( .A(n4585), .B(n4316), .Z(n4317) );
  XNOR U6153 ( .A(n4584), .B(n4317), .Z(out[886]) );
  OR U6154 ( .A(n4589), .B(n4318), .Z(n4319) );
  XNOR U6155 ( .A(n4588), .B(n4319), .Z(out[887]) );
  OR U6156 ( .A(n4593), .B(n4320), .Z(n4321) );
  XNOR U6157 ( .A(n4592), .B(n4321), .Z(out[888]) );
  OR U6158 ( .A(n4597), .B(n4322), .Z(n4323) );
  XNOR U6159 ( .A(n4596), .B(n4323), .Z(out[889]) );
  NOR U6160 ( .A(n4325), .B(n4324), .Z(n4326) );
  XNOR U6161 ( .A(n4327), .B(n4326), .Z(out[88]) );
  OR U6162 ( .A(n4601), .B(n4328), .Z(n4329) );
  XNOR U6163 ( .A(n4600), .B(n4329), .Z(out[890]) );
  OR U6164 ( .A(n4605), .B(n4330), .Z(n4331) );
  XNOR U6165 ( .A(n4604), .B(n4331), .Z(out[891]) );
  OR U6166 ( .A(n4609), .B(n4332), .Z(n4333) );
  XNOR U6167 ( .A(n4608), .B(n4333), .Z(out[892]) );
  OR U6168 ( .A(n4613), .B(n4334), .Z(n4335) );
  XNOR U6169 ( .A(n4612), .B(n4335), .Z(out[893]) );
  OR U6170 ( .A(n4617), .B(n4336), .Z(n4337) );
  XNOR U6171 ( .A(n4616), .B(n4337), .Z(out[894]) );
  OR U6172 ( .A(n4621), .B(n4338), .Z(n4339) );
  XNOR U6173 ( .A(n4620), .B(n4339), .Z(out[895]) );
  ANDN U6174 ( .B(n4341), .A(n4340), .Z(n4342) );
  XNOR U6175 ( .A(n4343), .B(n4342), .Z(out[896]) );
  ANDN U6176 ( .B(n4345), .A(n4344), .Z(n4346) );
  XNOR U6177 ( .A(n4347), .B(n4346), .Z(out[897]) );
  ANDN U6178 ( .B(n4349), .A(n4348), .Z(n4350) );
  XNOR U6179 ( .A(n4351), .B(n4350), .Z(out[898]) );
  ANDN U6180 ( .B(n4353), .A(n4352), .Z(n4354) );
  XNOR U6181 ( .A(n4355), .B(n4354), .Z(out[899]) );
  NOR U6182 ( .A(n4357), .B(n4356), .Z(n4358) );
  XNOR U6183 ( .A(n4359), .B(n4358), .Z(out[89]) );
  OR U6184 ( .A(n4361), .B(n4360), .Z(n4362) );
  XNOR U6185 ( .A(n4363), .B(n4362), .Z(out[8]) );
  ANDN U6186 ( .B(n4365), .A(n4364), .Z(n4366) );
  XNOR U6187 ( .A(n4367), .B(n4366), .Z(out[900]) );
  ANDN U6188 ( .B(n4369), .A(n4368), .Z(n4370) );
  XNOR U6189 ( .A(n4371), .B(n4370), .Z(out[901]) );
  ANDN U6190 ( .B(n4373), .A(n4372), .Z(n4374) );
  XNOR U6191 ( .A(n4375), .B(n4374), .Z(out[902]) );
  ANDN U6192 ( .B(n4377), .A(n4376), .Z(n4378) );
  XNOR U6193 ( .A(n4379), .B(n4378), .Z(out[903]) );
  ANDN U6194 ( .B(n4381), .A(n4380), .Z(n4382) );
  XNOR U6195 ( .A(n4383), .B(n4382), .Z(out[904]) );
  ANDN U6196 ( .B(n4385), .A(n4384), .Z(n4386) );
  XNOR U6197 ( .A(n4387), .B(n4386), .Z(out[905]) );
  ANDN U6198 ( .B(n4389), .A(n4388), .Z(n4390) );
  XNOR U6199 ( .A(n4391), .B(n4390), .Z(out[906]) );
  ANDN U6200 ( .B(n4393), .A(n4392), .Z(n4394) );
  XNOR U6201 ( .A(n4395), .B(n4394), .Z(out[907]) );
  ANDN U6202 ( .B(n4397), .A(n4396), .Z(n4398) );
  XNOR U6203 ( .A(n4399), .B(n4398), .Z(out[908]) );
  ANDN U6204 ( .B(n4401), .A(n4400), .Z(n4402) );
  XNOR U6205 ( .A(n4403), .B(n4402), .Z(out[909]) );
  NOR U6206 ( .A(n4405), .B(n4404), .Z(n4406) );
  XNOR U6207 ( .A(n4407), .B(n4406), .Z(out[90]) );
  ANDN U6208 ( .B(n4409), .A(n4408), .Z(n4410) );
  XNOR U6209 ( .A(n4411), .B(n4410), .Z(out[910]) );
  ANDN U6210 ( .B(n4413), .A(n4412), .Z(n4414) );
  XNOR U6211 ( .A(n4415), .B(n4414), .Z(out[911]) );
  ANDN U6212 ( .B(n4417), .A(n4416), .Z(n4418) );
  XNOR U6213 ( .A(n4419), .B(n4418), .Z(out[912]) );
  ANDN U6214 ( .B(n4421), .A(n4420), .Z(n4422) );
  XNOR U6215 ( .A(n4423), .B(n4422), .Z(out[913]) );
  ANDN U6216 ( .B(n4425), .A(n4424), .Z(n4426) );
  XNOR U6217 ( .A(n4427), .B(n4426), .Z(out[914]) );
  ANDN U6218 ( .B(n4429), .A(n4428), .Z(n4430) );
  XNOR U6219 ( .A(n4431), .B(n4430), .Z(out[915]) );
  ANDN U6220 ( .B(n4433), .A(n4432), .Z(n4434) );
  XNOR U6221 ( .A(n4435), .B(n4434), .Z(out[916]) );
  ANDN U6222 ( .B(n4437), .A(n4436), .Z(n4438) );
  XNOR U6223 ( .A(n4439), .B(n4438), .Z(out[917]) );
  ANDN U6224 ( .B(n4441), .A(n4440), .Z(n4442) );
  XNOR U6225 ( .A(n4443), .B(n4442), .Z(out[918]) );
  ANDN U6226 ( .B(n4445), .A(n4444), .Z(n4446) );
  XNOR U6227 ( .A(n4447), .B(n4446), .Z(out[919]) );
  NOR U6228 ( .A(n4449), .B(n4448), .Z(n4450) );
  XNOR U6229 ( .A(n4451), .B(n4450), .Z(out[91]) );
  ANDN U6230 ( .B(n4453), .A(n4452), .Z(n4454) );
  XNOR U6231 ( .A(n4455), .B(n4454), .Z(out[920]) );
  ANDN U6232 ( .B(n4457), .A(n4456), .Z(n4458) );
  XNOR U6233 ( .A(n4459), .B(n4458), .Z(out[921]) );
  ANDN U6234 ( .B(n4461), .A(n4460), .Z(n4462) );
  XNOR U6235 ( .A(n4463), .B(n4462), .Z(out[922]) );
  ANDN U6236 ( .B(n4465), .A(n4464), .Z(n4466) );
  XNOR U6237 ( .A(n4467), .B(n4466), .Z(out[923]) );
  ANDN U6238 ( .B(n4469), .A(n4468), .Z(n4470) );
  XNOR U6239 ( .A(n4471), .B(n4470), .Z(out[924]) );
  ANDN U6240 ( .B(n4473), .A(n4472), .Z(n4474) );
  XNOR U6241 ( .A(n4475), .B(n4474), .Z(out[925]) );
  ANDN U6242 ( .B(n4477), .A(n4476), .Z(n4478) );
  XNOR U6243 ( .A(n4479), .B(n4478), .Z(out[926]) );
  ANDN U6244 ( .B(n4481), .A(n4480), .Z(n4482) );
  XNOR U6245 ( .A(n4483), .B(n4482), .Z(out[927]) );
  ANDN U6246 ( .B(n4485), .A(n4484), .Z(n4486) );
  XNOR U6247 ( .A(n4487), .B(n4486), .Z(out[928]) );
  ANDN U6248 ( .B(n4489), .A(n4488), .Z(n4490) );
  XNOR U6249 ( .A(n4491), .B(n4490), .Z(out[929]) );
  ANDN U6250 ( .B(n4493), .A(n4492), .Z(n4494) );
  XNOR U6251 ( .A(n4495), .B(n4494), .Z(out[92]) );
  ANDN U6252 ( .B(n4497), .A(n4496), .Z(n4498) );
  XNOR U6253 ( .A(n4499), .B(n4498), .Z(out[930]) );
  ANDN U6254 ( .B(n4501), .A(n4500), .Z(n4502) );
  XNOR U6255 ( .A(n4503), .B(n4502), .Z(out[931]) );
  ANDN U6256 ( .B(n4505), .A(n4504), .Z(n4506) );
  XNOR U6257 ( .A(n4507), .B(n4506), .Z(out[932]) );
  ANDN U6258 ( .B(n4509), .A(n4508), .Z(n4510) );
  XNOR U6259 ( .A(n4511), .B(n4510), .Z(out[933]) );
  ANDN U6260 ( .B(n4513), .A(n4512), .Z(n4514) );
  XNOR U6261 ( .A(n4515), .B(n4514), .Z(out[934]) );
  ANDN U6262 ( .B(n4517), .A(n4516), .Z(n4518) );
  XNOR U6263 ( .A(n4519), .B(n4518), .Z(out[935]) );
  ANDN U6264 ( .B(n4521), .A(n4520), .Z(n4522) );
  XNOR U6265 ( .A(n4523), .B(n4522), .Z(out[936]) );
  ANDN U6266 ( .B(n4525), .A(n4524), .Z(n4526) );
  XNOR U6267 ( .A(n4527), .B(n4526), .Z(out[937]) );
  ANDN U6268 ( .B(n4529), .A(n4528), .Z(n4530) );
  XNOR U6269 ( .A(n4531), .B(n4530), .Z(out[938]) );
  ANDN U6270 ( .B(n4533), .A(n4532), .Z(n4534) );
  XNOR U6271 ( .A(n4535), .B(n4534), .Z(out[939]) );
  ANDN U6272 ( .B(n4537), .A(n4536), .Z(n4538) );
  XNOR U6273 ( .A(n4539), .B(n4538), .Z(out[93]) );
  ANDN U6274 ( .B(n4541), .A(n4540), .Z(n4542) );
  XNOR U6275 ( .A(n4543), .B(n4542), .Z(out[940]) );
  ANDN U6276 ( .B(n4545), .A(n4544), .Z(n4546) );
  XNOR U6277 ( .A(n4547), .B(n4546), .Z(out[941]) );
  ANDN U6278 ( .B(n4549), .A(n4548), .Z(n4550) );
  XNOR U6279 ( .A(n4551), .B(n4550), .Z(out[942]) );
  ANDN U6280 ( .B(n4553), .A(n4552), .Z(n4554) );
  XNOR U6281 ( .A(n4555), .B(n4554), .Z(out[943]) );
  ANDN U6282 ( .B(n4557), .A(n4556), .Z(n4558) );
  XNOR U6283 ( .A(n4559), .B(n4558), .Z(out[944]) );
  ANDN U6284 ( .B(n4561), .A(n4560), .Z(n4562) );
  XNOR U6285 ( .A(n4563), .B(n4562), .Z(out[945]) );
  ANDN U6286 ( .B(n4565), .A(n4564), .Z(n4566) );
  XNOR U6287 ( .A(n4567), .B(n4566), .Z(out[946]) );
  ANDN U6288 ( .B(n4569), .A(n4568), .Z(n4570) );
  XNOR U6289 ( .A(n4571), .B(n4570), .Z(out[947]) );
  ANDN U6290 ( .B(n4573), .A(n4572), .Z(n4574) );
  XNOR U6291 ( .A(n4575), .B(n4574), .Z(out[948]) );
  ANDN U6292 ( .B(n4577), .A(n4576), .Z(n4578) );
  XNOR U6293 ( .A(n4579), .B(n4578), .Z(out[949]) );
  ANDN U6294 ( .B(n4581), .A(n4580), .Z(n4582) );
  XNOR U6295 ( .A(n4583), .B(n4582), .Z(out[94]) );
  ANDN U6296 ( .B(n4585), .A(n4584), .Z(n4586) );
  XNOR U6297 ( .A(n4587), .B(n4586), .Z(out[950]) );
  ANDN U6298 ( .B(n4589), .A(n4588), .Z(n4590) );
  XNOR U6299 ( .A(n4591), .B(n4590), .Z(out[951]) );
  ANDN U6300 ( .B(n4593), .A(n4592), .Z(n4594) );
  XNOR U6301 ( .A(n4595), .B(n4594), .Z(out[952]) );
  ANDN U6302 ( .B(n4597), .A(n4596), .Z(n4598) );
  XNOR U6303 ( .A(n4599), .B(n4598), .Z(out[953]) );
  ANDN U6304 ( .B(n4601), .A(n4600), .Z(n4602) );
  XNOR U6305 ( .A(n4603), .B(n4602), .Z(out[954]) );
  ANDN U6306 ( .B(n4605), .A(n4604), .Z(n4606) );
  XNOR U6307 ( .A(n4607), .B(n4606), .Z(out[955]) );
  ANDN U6308 ( .B(n4609), .A(n4608), .Z(n4610) );
  XNOR U6309 ( .A(n4611), .B(n4610), .Z(out[956]) );
  ANDN U6310 ( .B(n4613), .A(n4612), .Z(n4614) );
  XNOR U6311 ( .A(n4615), .B(n4614), .Z(out[957]) );
  ANDN U6312 ( .B(n4617), .A(n4616), .Z(n4618) );
  XNOR U6313 ( .A(n4619), .B(n4618), .Z(out[958]) );
  ANDN U6314 ( .B(n4621), .A(n4620), .Z(n4622) );
  XNOR U6315 ( .A(n4623), .B(n4622), .Z(out[959]) );
  ANDN U6316 ( .B(n4625), .A(n4624), .Z(n4626) );
  XNOR U6317 ( .A(n4627), .B(n4626), .Z(out[95]) );
  ANDN U6318 ( .B(n4629), .A(n4628), .Z(n4630) );
  XNOR U6319 ( .A(n4631), .B(n4630), .Z(out[960]) );
  ANDN U6320 ( .B(n4633), .A(n4632), .Z(n4634) );
  XNOR U6321 ( .A(n4635), .B(n4634), .Z(out[961]) );
  ANDN U6322 ( .B(n4637), .A(n4636), .Z(n4638) );
  XNOR U6323 ( .A(n4639), .B(n4638), .Z(out[962]) );
  ANDN U6324 ( .B(n4641), .A(n4640), .Z(n4642) );
  XNOR U6325 ( .A(n4643), .B(n4642), .Z(out[963]) );
  ANDN U6326 ( .B(n4645), .A(n4644), .Z(n4646) );
  XNOR U6327 ( .A(n4647), .B(n4646), .Z(out[964]) );
  ANDN U6328 ( .B(n4649), .A(n4648), .Z(n4650) );
  XNOR U6329 ( .A(n4651), .B(n4650), .Z(out[965]) );
  ANDN U6330 ( .B(n4653), .A(n4652), .Z(n4654) );
  XNOR U6331 ( .A(n4655), .B(n4654), .Z(out[966]) );
  ANDN U6332 ( .B(n4657), .A(n4656), .Z(n4658) );
  XNOR U6333 ( .A(n4659), .B(n4658), .Z(out[967]) );
  ANDN U6334 ( .B(n4661), .A(n4660), .Z(n4662) );
  XNOR U6335 ( .A(n4663), .B(n4662), .Z(out[968]) );
  ANDN U6336 ( .B(n4665), .A(n4664), .Z(n4666) );
  XNOR U6337 ( .A(n4667), .B(n4666), .Z(out[969]) );
  ANDN U6338 ( .B(n4669), .A(n4668), .Z(n4670) );
  XNOR U6339 ( .A(n4671), .B(n4670), .Z(out[96]) );
  ANDN U6340 ( .B(n4673), .A(n4672), .Z(n4674) );
  XNOR U6341 ( .A(n4675), .B(n4674), .Z(out[970]) );
  ANDN U6342 ( .B(n4677), .A(n4676), .Z(n4678) );
  XNOR U6343 ( .A(n4679), .B(n4678), .Z(out[971]) );
  ANDN U6344 ( .B(n4681), .A(n4680), .Z(n4682) );
  XNOR U6345 ( .A(n4683), .B(n4682), .Z(out[972]) );
  ANDN U6346 ( .B(n4685), .A(n4684), .Z(n4686) );
  XNOR U6347 ( .A(n4687), .B(n4686), .Z(out[973]) );
  ANDN U6348 ( .B(n4689), .A(n4688), .Z(n4690) );
  XNOR U6349 ( .A(n4691), .B(n4690), .Z(out[974]) );
  ANDN U6350 ( .B(n4693), .A(n4692), .Z(n4694) );
  XNOR U6351 ( .A(n4695), .B(n4694), .Z(out[975]) );
  ANDN U6352 ( .B(n4697), .A(n4696), .Z(n4698) );
  XNOR U6353 ( .A(n4699), .B(n4698), .Z(out[976]) );
  ANDN U6354 ( .B(n4701), .A(n4700), .Z(n4702) );
  XNOR U6355 ( .A(n4703), .B(n4702), .Z(out[977]) );
  ANDN U6356 ( .B(n4705), .A(n4704), .Z(n4706) );
  XNOR U6357 ( .A(n4707), .B(n4706), .Z(out[978]) );
  ANDN U6358 ( .B(n4709), .A(n4708), .Z(n4710) );
  XNOR U6359 ( .A(n4711), .B(n4710), .Z(out[979]) );
  ANDN U6360 ( .B(n4713), .A(n4712), .Z(n4714) );
  XNOR U6361 ( .A(n4715), .B(n4714), .Z(out[97]) );
  ANDN U6362 ( .B(n4717), .A(n4716), .Z(n4718) );
  XNOR U6363 ( .A(n4719), .B(n4718), .Z(out[980]) );
  ANDN U6364 ( .B(n4721), .A(n4720), .Z(n4722) );
  XNOR U6365 ( .A(n4723), .B(n4722), .Z(out[981]) );
  ANDN U6366 ( .B(n4725), .A(n4724), .Z(n4726) );
  XNOR U6367 ( .A(n4727), .B(n4726), .Z(out[982]) );
  ANDN U6368 ( .B(n4729), .A(n4728), .Z(n4730) );
  XNOR U6369 ( .A(n4731), .B(n4730), .Z(out[983]) );
  ANDN U6370 ( .B(n4733), .A(n4732), .Z(n4734) );
  XNOR U6371 ( .A(n4735), .B(n4734), .Z(out[984]) );
  ANDN U6372 ( .B(n4737), .A(n4736), .Z(n4738) );
  XNOR U6373 ( .A(n4739), .B(n4738), .Z(out[985]) );
  ANDN U6374 ( .B(n4741), .A(n4740), .Z(n4742) );
  XNOR U6375 ( .A(n4743), .B(n4742), .Z(out[986]) );
  ANDN U6376 ( .B(n4745), .A(n4744), .Z(n4746) );
  XNOR U6377 ( .A(n4747), .B(n4746), .Z(out[987]) );
  ANDN U6378 ( .B(n4749), .A(n4748), .Z(n4750) );
  XNOR U6379 ( .A(n4751), .B(n4750), .Z(out[988]) );
  ANDN U6380 ( .B(n4753), .A(n4752), .Z(n4754) );
  XNOR U6381 ( .A(n4755), .B(n4754), .Z(out[989]) );
  ANDN U6382 ( .B(n4757), .A(n4756), .Z(n4758) );
  XNOR U6383 ( .A(n4759), .B(n4758), .Z(out[98]) );
  ANDN U6384 ( .B(n4761), .A(n4760), .Z(n4762) );
  XNOR U6385 ( .A(n4763), .B(n4762), .Z(out[990]) );
  ANDN U6386 ( .B(n4765), .A(n4764), .Z(n4766) );
  XNOR U6387 ( .A(n4767), .B(n4766), .Z(out[991]) );
  ANDN U6388 ( .B(n4769), .A(n4768), .Z(n4770) );
  XNOR U6389 ( .A(n4771), .B(n4770), .Z(out[992]) );
  ANDN U6390 ( .B(n4773), .A(n4772), .Z(n4774) );
  XNOR U6391 ( .A(n4775), .B(n4774), .Z(out[993]) );
  ANDN U6392 ( .B(n4777), .A(n4776), .Z(n4778) );
  XNOR U6393 ( .A(n4779), .B(n4778), .Z(out[994]) );
  ANDN U6394 ( .B(n4781), .A(n4780), .Z(n4782) );
  XNOR U6395 ( .A(n4783), .B(n4782), .Z(out[995]) );
  ANDN U6396 ( .B(n4785), .A(n4784), .Z(n4786) );
  XNOR U6397 ( .A(n4787), .B(n4786), .Z(out[996]) );
  ANDN U6398 ( .B(n4789), .A(n4788), .Z(n4790) );
  XNOR U6399 ( .A(n4791), .B(n4790), .Z(out[997]) );
  ANDN U6400 ( .B(n4793), .A(n4792), .Z(n4794) );
  XNOR U6401 ( .A(n4795), .B(n4794), .Z(out[998]) );
  ANDN U6402 ( .B(n4797), .A(n4796), .Z(n4798) );
  XNOR U6403 ( .A(n4799), .B(n4798), .Z(out[999]) );
  ANDN U6404 ( .B(n4801), .A(n4800), .Z(n4802) );
  XNOR U6405 ( .A(n4803), .B(n4802), .Z(out[99]) );
  OR U6406 ( .A(n4805), .B(n4804), .Z(n4806) );
  XNOR U6407 ( .A(n4807), .B(n4806), .Z(out[9]) );
endmodule


module round_5 ( in, round_const, out );
  input [1599:0] in;
  input [63:0] round_const;
  output [1599:0] out;
  wire   round_const_63, round_const_31, round_const_15, round_const_7,
         round_const_3, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
         n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
         n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
         n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
         n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
         n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
         n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
         n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
         n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
         n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
         n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
         n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
         n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807;
  assign round_const_63 = round_const[63];
  assign round_const_31 = round_const[31];
  assign round_const_15 = round_const[15];
  assign round_const_7 = round_const[7];
  assign round_const_3 = round_const[3];

  XOR U1 ( .A(in[1469]), .B(in[509]), .Z(n2) );
  XNOR U2 ( .A(in[829]), .B(in[189]), .Z(n1) );
  XNOR U3 ( .A(n2), .B(n1), .Z(n3) );
  XOR U4 ( .A(in[1149]), .B(n3), .Z(n872) );
  XOR U5 ( .A(in[1598]), .B(in[638]), .Z(n5) );
  XNOR U6 ( .A(in[958]), .B(in[318]), .Z(n4) );
  XNOR U7 ( .A(n5), .B(n4), .Z(n6) );
  XOR U8 ( .A(in[1278]), .B(n6), .Z(n1473) );
  XNOR U9 ( .A(n872), .B(n1473), .Z(n3815) );
  XNOR U10 ( .A(in[254]), .B(n3815), .Z(n3577) );
  XOR U11 ( .A(in[1345]), .B(in[65]), .Z(n8) );
  XNOR U12 ( .A(in[1025]), .B(in[385]), .Z(n7) );
  XNOR U13 ( .A(n8), .B(n7), .Z(n9) );
  XOR U14 ( .A(in[705]), .B(n9), .Z(n1481) );
  XOR U15 ( .A(in[1474]), .B(in[514]), .Z(n11) );
  XNOR U16 ( .A(in[834]), .B(in[194]), .Z(n10) );
  XNOR U17 ( .A(n11), .B(n10), .Z(n12) );
  XNOR U18 ( .A(in[1154]), .B(n12), .Z(n1188) );
  XNOR U19 ( .A(n1481), .B(n1188), .Z(n3570) );
  XNOR U20 ( .A(in[1410]), .B(n3570), .Z(n3576) );
  XOR U21 ( .A(in[328]), .B(in[8]), .Z(n14) );
  XNOR U22 ( .A(in[968]), .B(in[648]), .Z(n13) );
  XNOR U23 ( .A(n14), .B(n13), .Z(n15) );
  XOR U24 ( .A(in[1288]), .B(n15), .Z(n1209) );
  XOR U25 ( .A(in[137]), .B(in[457]), .Z(n17) );
  XNOR U26 ( .A(in[777]), .B(in[1417]), .Z(n16) );
  XNOR U27 ( .A(n17), .B(n16), .Z(n18) );
  XOR U28 ( .A(in[1097]), .B(n18), .Z(n1141) );
  XNOR U29 ( .A(n1209), .B(n1141), .Z(n4086) );
  XNOR U30 ( .A(in[1033]), .B(n4086), .Z(n2609) );
  NAND U31 ( .A(n3576), .B(n2609), .Z(n19) );
  XNOR U32 ( .A(n3577), .B(n19), .Z(out[0]) );
  XOR U33 ( .A(in[1515]), .B(in[555]), .Z(n21) );
  XNOR U34 ( .A(in[875]), .B(in[235]), .Z(n20) );
  XNOR U35 ( .A(n21), .B(n20), .Z(n22) );
  XOR U36 ( .A(in[1195]), .B(n22), .Z(n1329) );
  XOR U37 ( .A(in[1386]), .B(in[106]), .Z(n24) );
  XNOR U38 ( .A(in[1066]), .B(in[746]), .Z(n23) );
  XNOR U39 ( .A(n24), .B(n23), .Z(n25) );
  XOR U40 ( .A(in[426]), .B(n25), .Z(n475) );
  XNOR U41 ( .A(n1329), .B(n475), .Z(n3750) );
  XNOR U42 ( .A(in[171]), .B(n3750), .Z(n1301) );
  XOR U43 ( .A(in[140]), .B(in[460]), .Z(n27) );
  XNOR U44 ( .A(in[1100]), .B(in[1420]), .Z(n26) );
  XNOR U45 ( .A(n27), .B(n26), .Z(n28) );
  XOR U46 ( .A(in[780]), .B(n28), .Z(n1159) );
  XOR U47 ( .A(in[971]), .B(in[1291]), .Z(n30) );
  XNOR U48 ( .A(in[11]), .B(in[331]), .Z(n29) );
  XNOR U49 ( .A(n30), .B(n29), .Z(n31) );
  XNOR U50 ( .A(in[651]), .B(n31), .Z(n1220) );
  XNOR U51 ( .A(n1159), .B(n1220), .Z(n4095) );
  XNOR U52 ( .A(in[1356]), .B(n4095), .Z(n1696) );
  XOR U53 ( .A(in[1364]), .B(in[724]), .Z(n33) );
  XNOR U54 ( .A(in[84]), .B(in[404]), .Z(n32) );
  XNOR U55 ( .A(n33), .B(n32), .Z(n34) );
  XOR U56 ( .A(in[1044]), .B(n34), .Z(n777) );
  XOR U57 ( .A(in[1555]), .B(in[595]), .Z(n36) );
  XNOR U58 ( .A(in[915]), .B(in[275]), .Z(n35) );
  XNOR U59 ( .A(n36), .B(n35), .Z(n37) );
  XOR U60 ( .A(in[1235]), .B(n37), .Z(n489) );
  XNOR U61 ( .A(n777), .B(n489), .Z(n3882) );
  XNOR U62 ( .A(in[980]), .B(n3882), .Z(n1693) );
  NAND U63 ( .A(n1696), .B(n1693), .Z(n38) );
  XNOR U64 ( .A(n1301), .B(n38), .Z(out[1000]) );
  XOR U65 ( .A(in[1516]), .B(in[556]), .Z(n40) );
  XNOR U66 ( .A(in[876]), .B(in[236]), .Z(n39) );
  XNOR U67 ( .A(n40), .B(n39), .Z(n41) );
  XOR U68 ( .A(in[1196]), .B(n41), .Z(n1333) );
  XOR U69 ( .A(in[1387]), .B(in[107]), .Z(n43) );
  XNOR U70 ( .A(in[1067]), .B(in[747]), .Z(n42) );
  XNOR U71 ( .A(n43), .B(n42), .Z(n44) );
  XOR U72 ( .A(in[427]), .B(n44), .Z(n486) );
  XNOR U73 ( .A(n1333), .B(n486), .Z(n3758) );
  XNOR U74 ( .A(in[172]), .B(n3758), .Z(n1305) );
  XOR U75 ( .A(in[972]), .B(in[12]), .Z(n46) );
  XNOR U76 ( .A(in[1292]), .B(in[332]), .Z(n45) );
  XNOR U77 ( .A(n46), .B(n45), .Z(n47) );
  XOR U78 ( .A(in[652]), .B(n47), .Z(n1223) );
  XOR U79 ( .A(in[141]), .B(in[461]), .Z(n49) );
  XNOR U80 ( .A(in[1101]), .B(in[1421]), .Z(n48) );
  XNOR U81 ( .A(n49), .B(n48), .Z(n50) );
  XNOR U82 ( .A(in[781]), .B(n50), .Z(n1164) );
  XNOR U83 ( .A(n1223), .B(n1164), .Z(n4098) );
  XNOR U84 ( .A(in[1357]), .B(n4098), .Z(n1700) );
  XOR U85 ( .A(in[1365]), .B(in[725]), .Z(n52) );
  XNOR U86 ( .A(in[85]), .B(in[405]), .Z(n51) );
  XNOR U87 ( .A(n52), .B(n51), .Z(n53) );
  XOR U88 ( .A(in[1045]), .B(n53), .Z(n790) );
  XOR U89 ( .A(in[1556]), .B(in[596]), .Z(n55) );
  XNOR U90 ( .A(in[916]), .B(in[276]), .Z(n54) );
  XNOR U91 ( .A(n55), .B(n54), .Z(n56) );
  XOR U92 ( .A(in[1236]), .B(n56), .Z(n504) );
  XNOR U93 ( .A(n790), .B(n504), .Z(n3884) );
  XNOR U94 ( .A(in[981]), .B(n3884), .Z(n1697) );
  NAND U95 ( .A(n1700), .B(n1697), .Z(n57) );
  XNOR U96 ( .A(n1305), .B(n57), .Z(out[1001]) );
  XOR U97 ( .A(in[1388]), .B(in[108]), .Z(n59) );
  XNOR U98 ( .A(in[1068]), .B(in[748]), .Z(n58) );
  XNOR U99 ( .A(n59), .B(n58), .Z(n60) );
  XOR U100 ( .A(in[428]), .B(n60), .Z(n1395) );
  XOR U101 ( .A(in[1517]), .B(in[557]), .Z(n62) );
  XNOR U102 ( .A(in[877]), .B(in[237]), .Z(n61) );
  XNOR U103 ( .A(n62), .B(n61), .Z(n63) );
  XOR U104 ( .A(in[1197]), .B(n63), .Z(n1337) );
  XNOR U105 ( .A(n1395), .B(n1337), .Z(n3762) );
  XNOR U106 ( .A(in[173]), .B(n3762), .Z(n1310) );
  XOR U107 ( .A(in[973]), .B(in[13]), .Z(n65) );
  XNOR U108 ( .A(in[1293]), .B(in[333]), .Z(n64) );
  XNOR U109 ( .A(n65), .B(n64), .Z(n66) );
  XOR U110 ( .A(in[653]), .B(n66), .Z(n1226) );
  XOR U111 ( .A(in[142]), .B(in[1422]), .Z(n68) );
  XNOR U112 ( .A(in[1102]), .B(in[782]), .Z(n67) );
  XNOR U113 ( .A(n68), .B(n67), .Z(n69) );
  XNOR U114 ( .A(in[462]), .B(n69), .Z(n1169) );
  XNOR U115 ( .A(n1226), .B(n1169), .Z(n4101) );
  XNOR U116 ( .A(in[1358]), .B(n4101), .Z(n1704) );
  XOR U117 ( .A(in[1366]), .B(in[726]), .Z(n71) );
  XNOR U118 ( .A(in[86]), .B(in[406]), .Z(n70) );
  XNOR U119 ( .A(n71), .B(n70), .Z(n72) );
  XOR U120 ( .A(in[1046]), .B(n72), .Z(n803) );
  XOR U121 ( .A(in[1557]), .B(in[597]), .Z(n74) );
  XNOR U122 ( .A(in[917]), .B(in[277]), .Z(n73) );
  XNOR U123 ( .A(n74), .B(n73), .Z(n75) );
  XOR U124 ( .A(in[1237]), .B(n75), .Z(n519) );
  XNOR U125 ( .A(n803), .B(n519), .Z(n3886) );
  XNOR U126 ( .A(in[982]), .B(n3886), .Z(n1701) );
  NAND U127 ( .A(n1704), .B(n1701), .Z(n76) );
  XNOR U128 ( .A(n1310), .B(n76), .Z(out[1002]) );
  XOR U129 ( .A(in[1389]), .B(in[109]), .Z(n78) );
  XNOR U130 ( .A(in[1069]), .B(in[749]), .Z(n77) );
  XNOR U131 ( .A(n78), .B(n77), .Z(n79) );
  XOR U132 ( .A(in[429]), .B(n79), .Z(n1399) );
  XOR U133 ( .A(in[1518]), .B(in[558]), .Z(n81) );
  XNOR U134 ( .A(in[878]), .B(in[238]), .Z(n80) );
  XNOR U135 ( .A(n81), .B(n80), .Z(n82) );
  XOR U136 ( .A(in[1198]), .B(n82), .Z(n1341) );
  XNOR U137 ( .A(n1399), .B(n1341), .Z(n3766) );
  XNOR U138 ( .A(in[174]), .B(n3766), .Z(n1314) );
  XOR U139 ( .A(in[143]), .B(in[1423]), .Z(n84) );
  XNOR U140 ( .A(in[1103]), .B(in[783]), .Z(n83) );
  XNOR U141 ( .A(n84), .B(n83), .Z(n85) );
  XOR U142 ( .A(in[463]), .B(n85), .Z(n1174) );
  XOR U143 ( .A(in[974]), .B(in[14]), .Z(n87) );
  XNOR U144 ( .A(in[1294]), .B(in[334]), .Z(n86) );
  XNOR U145 ( .A(n87), .B(n86), .Z(n88) );
  XNOR U146 ( .A(in[654]), .B(n88), .Z(n1229) );
  XNOR U147 ( .A(n1174), .B(n1229), .Z(n4104) );
  XNOR U148 ( .A(in[1359]), .B(n4104), .Z(n1708) );
  XOR U149 ( .A(in[1367]), .B(in[727]), .Z(n90) );
  XNOR U150 ( .A(in[87]), .B(in[407]), .Z(n89) );
  XNOR U151 ( .A(n90), .B(n89), .Z(n91) );
  XOR U152 ( .A(in[1047]), .B(n91), .Z(n816) );
  XOR U153 ( .A(in[1558]), .B(in[598]), .Z(n93) );
  XNOR U154 ( .A(in[918]), .B(in[278]), .Z(n92) );
  XNOR U155 ( .A(n93), .B(n92), .Z(n94) );
  XOR U156 ( .A(in[1238]), .B(n94), .Z(n534) );
  XNOR U157 ( .A(n816), .B(n534), .Z(n3888) );
  XNOR U158 ( .A(in[983]), .B(n3888), .Z(n1705) );
  NAND U159 ( .A(n1708), .B(n1705), .Z(n95) );
  XNOR U160 ( .A(n1314), .B(n95), .Z(out[1003]) );
  XOR U161 ( .A(in[1390]), .B(in[110]), .Z(n97) );
  XNOR U162 ( .A(in[1070]), .B(in[750]), .Z(n96) );
  XNOR U163 ( .A(n97), .B(n96), .Z(n98) );
  XOR U164 ( .A(in[430]), .B(n98), .Z(n1403) );
  XOR U165 ( .A(in[1519]), .B(in[559]), .Z(n100) );
  XNOR U166 ( .A(in[879]), .B(in[239]), .Z(n99) );
  XNOR U167 ( .A(n100), .B(n99), .Z(n101) );
  XOR U168 ( .A(in[1199]), .B(n101), .Z(n1345) );
  XNOR U169 ( .A(n1403), .B(n1345), .Z(n3770) );
  XNOR U170 ( .A(in[175]), .B(n3770), .Z(n1318) );
  XOR U171 ( .A(in[144]), .B(in[1424]), .Z(n103) );
  XNOR U172 ( .A(in[1104]), .B(in[784]), .Z(n102) );
  XNOR U173 ( .A(n103), .B(n102), .Z(n104) );
  XOR U174 ( .A(in[464]), .B(n104), .Z(n1179) );
  XOR U175 ( .A(in[975]), .B(in[15]), .Z(n106) );
  XNOR U176 ( .A(in[1295]), .B(in[335]), .Z(n105) );
  XNOR U177 ( .A(n106), .B(n105), .Z(n107) );
  XNOR U178 ( .A(in[655]), .B(n107), .Z(n1232) );
  XNOR U179 ( .A(n1179), .B(n1232), .Z(n4107) );
  XNOR U180 ( .A(in[1360]), .B(n4107), .Z(n1713) );
  XOR U181 ( .A(in[1368]), .B(in[728]), .Z(n109) );
  XNOR U182 ( .A(in[88]), .B(in[408]), .Z(n108) );
  XNOR U183 ( .A(n109), .B(n108), .Z(n110) );
  XOR U184 ( .A(in[1048]), .B(n110), .Z(n829) );
  XOR U185 ( .A(in[1559]), .B(in[599]), .Z(n112) );
  XNOR U186 ( .A(in[919]), .B(in[279]), .Z(n111) );
  XNOR U187 ( .A(n112), .B(n111), .Z(n113) );
  XOR U188 ( .A(in[1239]), .B(n113), .Z(n549) );
  XNOR U189 ( .A(n829), .B(n549), .Z(n3890) );
  XNOR U190 ( .A(in[984]), .B(n3890), .Z(n1710) );
  NAND U191 ( .A(n1713), .B(n1710), .Z(n114) );
  XNOR U192 ( .A(n1318), .B(n114), .Z(out[1004]) );
  XOR U193 ( .A(in[1391]), .B(in[111]), .Z(n116) );
  XNOR U194 ( .A(in[1071]), .B(in[751]), .Z(n115) );
  XNOR U195 ( .A(n116), .B(n115), .Z(n117) );
  XOR U196 ( .A(in[431]), .B(n117), .Z(n1407) );
  XOR U197 ( .A(in[1520]), .B(in[560]), .Z(n119) );
  XNOR U198 ( .A(in[880]), .B(in[240]), .Z(n118) );
  XNOR U199 ( .A(n119), .B(n118), .Z(n120) );
  XOR U200 ( .A(in[1200]), .B(n120), .Z(n1350) );
  XNOR U201 ( .A(n1407), .B(n1350), .Z(n3774) );
  XNOR U202 ( .A(in[176]), .B(n3774), .Z(n1322) );
  XOR U203 ( .A(in[976]), .B(in[16]), .Z(n122) );
  XNOR U204 ( .A(in[1296]), .B(in[336]), .Z(n121) );
  XNOR U205 ( .A(n122), .B(n121), .Z(n123) );
  XOR U206 ( .A(in[656]), .B(n123), .Z(n1235) );
  XOR U207 ( .A(in[145]), .B(in[1425]), .Z(n125) );
  XNOR U208 ( .A(in[1105]), .B(in[785]), .Z(n124) );
  XNOR U209 ( .A(n125), .B(n124), .Z(n126) );
  XNOR U210 ( .A(in[465]), .B(n126), .Z(n1184) );
  XNOR U211 ( .A(n1235), .B(n1184), .Z(n4114) );
  XNOR U212 ( .A(in[1361]), .B(n4114), .Z(n1717) );
  XOR U213 ( .A(in[1369]), .B(in[729]), .Z(n128) );
  XNOR U214 ( .A(in[89]), .B(in[409]), .Z(n127) );
  XNOR U215 ( .A(n128), .B(n127), .Z(n129) );
  XOR U216 ( .A(in[1049]), .B(n129), .Z(n842) );
  XOR U217 ( .A(in[1560]), .B(in[600]), .Z(n131) );
  XNOR U218 ( .A(in[920]), .B(in[280]), .Z(n130) );
  XNOR U219 ( .A(n131), .B(n130), .Z(n132) );
  XOR U220 ( .A(in[1240]), .B(n132), .Z(n564) );
  XNOR U221 ( .A(n842), .B(n564), .Z(n3892) );
  XNOR U222 ( .A(in[985]), .B(n3892), .Z(n1714) );
  NAND U223 ( .A(n1717), .B(n1714), .Z(n133) );
  XNOR U224 ( .A(n1322), .B(n133), .Z(out[1005]) );
  XOR U225 ( .A(in[1392]), .B(in[112]), .Z(n135) );
  XNOR U226 ( .A(in[1072]), .B(in[752]), .Z(n134) );
  XNOR U227 ( .A(n135), .B(n134), .Z(n136) );
  XOR U228 ( .A(in[432]), .B(n136), .Z(n1411) );
  XOR U229 ( .A(in[1521]), .B(in[561]), .Z(n138) );
  XNOR U230 ( .A(in[881]), .B(in[241]), .Z(n137) );
  XNOR U231 ( .A(n138), .B(n137), .Z(n139) );
  XOR U232 ( .A(in[1201]), .B(n139), .Z(n1354) );
  XNOR U233 ( .A(n1411), .B(n1354), .Z(n3778) );
  XNOR U234 ( .A(in[177]), .B(n3778), .Z(n1326) );
  XOR U235 ( .A(in[1426]), .B(in[466]), .Z(n141) );
  XNOR U236 ( .A(in[786]), .B(in[146]), .Z(n140) );
  XNOR U237 ( .A(n141), .B(n140), .Z(n142) );
  XOR U238 ( .A(in[1106]), .B(n142), .Z(n488) );
  XOR U239 ( .A(in[17]), .B(in[657]), .Z(n144) );
  XNOR U240 ( .A(in[977]), .B(in[337]), .Z(n143) );
  XNOR U241 ( .A(n144), .B(n143), .Z(n145) );
  XNOR U242 ( .A(in[1297]), .B(n145), .Z(n1238) );
  XNOR U243 ( .A(n488), .B(n1238), .Z(n4117) );
  XNOR U244 ( .A(n4117), .B(in[1362]), .Z(n1721) );
  XOR U245 ( .A(in[1370]), .B(in[730]), .Z(n147) );
  XNOR U246 ( .A(in[90]), .B(in[410]), .Z(n146) );
  XNOR U247 ( .A(n147), .B(n146), .Z(n148) );
  XOR U248 ( .A(in[1050]), .B(n148), .Z(n857) );
  XOR U249 ( .A(in[1561]), .B(in[601]), .Z(n150) );
  XNOR U250 ( .A(in[921]), .B(in[281]), .Z(n149) );
  XNOR U251 ( .A(n150), .B(n149), .Z(n151) );
  XOR U252 ( .A(in[1241]), .B(n151), .Z(n590) );
  XNOR U253 ( .A(n857), .B(n590), .Z(n3894) );
  XNOR U254 ( .A(in[986]), .B(n3894), .Z(n1718) );
  NAND U255 ( .A(n1721), .B(n1718), .Z(n152) );
  XNOR U256 ( .A(n1326), .B(n152), .Z(out[1006]) );
  XOR U257 ( .A(in[1393]), .B(in[113]), .Z(n154) );
  XNOR U258 ( .A(in[1073]), .B(in[753]), .Z(n153) );
  XNOR U259 ( .A(n154), .B(n153), .Z(n155) );
  XOR U260 ( .A(in[433]), .B(n155), .Z(n1415) );
  XOR U261 ( .A(in[1522]), .B(in[562]), .Z(n157) );
  XNOR U262 ( .A(in[882]), .B(in[242]), .Z(n156) );
  XNOR U263 ( .A(n157), .B(n156), .Z(n158) );
  XOR U264 ( .A(in[1202]), .B(n158), .Z(n1358) );
  XNOR U265 ( .A(n1415), .B(n1358), .Z(n3782) );
  XNOR U266 ( .A(in[178]), .B(n3782), .Z(n1330) );
  XOR U267 ( .A(in[978]), .B(in[18]), .Z(n160) );
  XNOR U268 ( .A(in[1298]), .B(in[338]), .Z(n159) );
  XNOR U269 ( .A(n160), .B(n159), .Z(n161) );
  XOR U270 ( .A(in[658]), .B(n161), .Z(n1241) );
  XOR U271 ( .A(in[147]), .B(in[1427]), .Z(n163) );
  XNOR U272 ( .A(in[1107]), .B(in[787]), .Z(n162) );
  XNOR U273 ( .A(n163), .B(n162), .Z(n164) );
  XNOR U274 ( .A(in[467]), .B(n164), .Z(n503) );
  XNOR U275 ( .A(n1241), .B(n503), .Z(n4120) );
  XNOR U276 ( .A(in[1363]), .B(n4120), .Z(n1725) );
  XOR U277 ( .A(in[1371]), .B(in[731]), .Z(n166) );
  XNOR U278 ( .A(in[91]), .B(in[411]), .Z(n165) );
  XNOR U279 ( .A(n166), .B(n165), .Z(n167) );
  XOR U280 ( .A(in[1051]), .B(n167), .Z(n870) );
  XOR U281 ( .A(in[1562]), .B(in[602]), .Z(n169) );
  XNOR U282 ( .A(in[922]), .B(in[282]), .Z(n168) );
  XNOR U283 ( .A(n169), .B(n168), .Z(n170) );
  XOR U284 ( .A(in[1242]), .B(n170), .Z(n605) );
  XNOR U285 ( .A(n870), .B(n605), .Z(n3896) );
  XNOR U286 ( .A(in[987]), .B(n3896), .Z(n1722) );
  NAND U287 ( .A(n1725), .B(n1722), .Z(n171) );
  XNOR U288 ( .A(n1330), .B(n171), .Z(out[1007]) );
  XOR U289 ( .A(in[1394]), .B(in[114]), .Z(n173) );
  XNOR U290 ( .A(in[1074]), .B(in[754]), .Z(n172) );
  XNOR U291 ( .A(n173), .B(n172), .Z(n174) );
  XOR U292 ( .A(in[434]), .B(n174), .Z(n1419) );
  XOR U293 ( .A(in[1523]), .B(in[563]), .Z(n176) );
  XNOR U294 ( .A(in[883]), .B(in[243]), .Z(n175) );
  XNOR U295 ( .A(n176), .B(n175), .Z(n177) );
  XOR U296 ( .A(in[1203]), .B(n177), .Z(n1362) );
  XNOR U297 ( .A(n1419), .B(n1362), .Z(n3786) );
  XNOR U298 ( .A(in[179]), .B(n3786), .Z(n1334) );
  XOR U299 ( .A(in[148]), .B(in[1428]), .Z(n179) );
  XNOR U300 ( .A(in[1108]), .B(in[788]), .Z(n178) );
  XNOR U301 ( .A(n179), .B(n178), .Z(n180) );
  XOR U302 ( .A(in[468]), .B(n180), .Z(n518) );
  XOR U303 ( .A(in[979]), .B(in[19]), .Z(n182) );
  XNOR U304 ( .A(in[1299]), .B(in[339]), .Z(n181) );
  XNOR U305 ( .A(n182), .B(n181), .Z(n183) );
  XNOR U306 ( .A(in[659]), .B(n183), .Z(n1245) );
  XNOR U307 ( .A(n518), .B(n1245), .Z(n4123) );
  XNOR U308 ( .A(in[1364]), .B(n4123), .Z(n1729) );
  XOR U309 ( .A(in[1372]), .B(in[732]), .Z(n185) );
  XNOR U310 ( .A(in[92]), .B(in[412]), .Z(n184) );
  XNOR U311 ( .A(n185), .B(n184), .Z(n186) );
  XOR U312 ( .A(in[1052]), .B(n186), .Z(n890) );
  XOR U313 ( .A(in[1563]), .B(in[603]), .Z(n188) );
  XNOR U314 ( .A(in[923]), .B(in[283]), .Z(n187) );
  XNOR U315 ( .A(n188), .B(n187), .Z(n189) );
  XOR U316 ( .A(in[1243]), .B(n189), .Z(n620) );
  XNOR U317 ( .A(n890), .B(n620), .Z(n3900) );
  XNOR U318 ( .A(in[988]), .B(n3900), .Z(n1726) );
  NAND U319 ( .A(n1729), .B(n1726), .Z(n190) );
  XNOR U320 ( .A(n1334), .B(n190), .Z(out[1008]) );
  XOR U321 ( .A(in[1395]), .B(in[115]), .Z(n192) );
  XNOR U322 ( .A(in[1075]), .B(in[755]), .Z(n191) );
  XNOR U323 ( .A(n192), .B(n191), .Z(n193) );
  XOR U324 ( .A(in[435]), .B(n193), .Z(n1423) );
  XOR U325 ( .A(in[1524]), .B(in[564]), .Z(n195) );
  XNOR U326 ( .A(in[884]), .B(in[244]), .Z(n194) );
  XNOR U327 ( .A(n195), .B(n194), .Z(n196) );
  XOR U328 ( .A(in[1204]), .B(n196), .Z(n1366) );
  XNOR U329 ( .A(n1423), .B(n1366), .Z(n3790) );
  XNOR U330 ( .A(in[180]), .B(n3790), .Z(n1338) );
  XOR U331 ( .A(in[340]), .B(in[660]), .Z(n198) );
  XNOR U332 ( .A(in[20]), .B(in[1300]), .Z(n197) );
  XNOR U333 ( .A(n198), .B(n197), .Z(n199) );
  XOR U334 ( .A(in[980]), .B(n199), .Z(n1248) );
  XOR U335 ( .A(in[149]), .B(in[1429]), .Z(n201) );
  XNOR U336 ( .A(in[1109]), .B(in[789]), .Z(n200) );
  XNOR U337 ( .A(n201), .B(n200), .Z(n202) );
  XNOR U338 ( .A(in[469]), .B(n202), .Z(n533) );
  XNOR U339 ( .A(n1248), .B(n533), .Z(n4126) );
  XNOR U340 ( .A(in[1365]), .B(n4126), .Z(n1733) );
  XOR U341 ( .A(in[1373]), .B(in[733]), .Z(n204) );
  XNOR U342 ( .A(in[93]), .B(in[413]), .Z(n203) );
  XNOR U343 ( .A(n204), .B(n203), .Z(n205) );
  XOR U344 ( .A(in[1053]), .B(n205), .Z(n903) );
  XOR U345 ( .A(in[1564]), .B(in[604]), .Z(n207) );
  XNOR U346 ( .A(in[924]), .B(in[284]), .Z(n206) );
  XNOR U347 ( .A(n207), .B(n206), .Z(n208) );
  XOR U348 ( .A(in[1244]), .B(n208), .Z(n635) );
  XNOR U349 ( .A(n903), .B(n635), .Z(n3902) );
  XNOR U350 ( .A(in[989]), .B(n3902), .Z(n1730) );
  NAND U351 ( .A(n1733), .B(n1730), .Z(n209) );
  XNOR U352 ( .A(n1338), .B(n209), .Z(out[1009]) );
  XOR U353 ( .A(in[1339]), .B(in[59]), .Z(n211) );
  XNOR U354 ( .A(in[699]), .B(in[379]), .Z(n210) );
  XNOR U355 ( .A(n211), .B(n210), .Z(n212) );
  XOR U356 ( .A(in[1019]), .B(n212), .Z(n861) );
  XOR U357 ( .A(in[1530]), .B(in[570]), .Z(n214) );
  XNOR U358 ( .A(in[1210]), .B(in[250]), .Z(n213) );
  XNOR U359 ( .A(n214), .B(n213), .Z(n215) );
  XOR U360 ( .A(in[890]), .B(n215), .Z(n327) );
  XNOR U361 ( .A(n861), .B(n327), .Z(n3592) );
  XNOR U362 ( .A(in[635]), .B(n3592), .Z(n2550) );
  XOR U363 ( .A(in[161]), .B(in[1441]), .Z(n217) );
  XNOR U364 ( .A(in[801]), .B(in[1121]), .Z(n216) );
  XNOR U365 ( .A(n217), .B(n216), .Z(n218) );
  XOR U366 ( .A(in[481]), .B(n218), .Z(n454) );
  XOR U367 ( .A(in[1570]), .B(in[610]), .Z(n220) );
  XNOR U368 ( .A(in[930]), .B(in[290]), .Z(n219) );
  XNOR U369 ( .A(n220), .B(n219), .Z(n221) );
  XNOR U370 ( .A(in[1250]), .B(n221), .Z(n337) );
  XNOR U371 ( .A(n454), .B(n337), .Z(n3689) );
  XNOR U372 ( .A(in[226]), .B(n3689), .Z(n2831) );
  XOR U373 ( .A(in[1510]), .B(in[550]), .Z(n223) );
  XNOR U374 ( .A(in[870]), .B(in[230]), .Z(n222) );
  XNOR U375 ( .A(n223), .B(n222), .Z(n224) );
  XOR U376 ( .A(in[1190]), .B(n224), .Z(n1309) );
  XOR U377 ( .A(in[1061]), .B(in[421]), .Z(n226) );
  XNOR U378 ( .A(in[741]), .B(in[1381]), .Z(n225) );
  XNOR U379 ( .A(n226), .B(n225), .Z(n227) );
  XOR U380 ( .A(in[101]), .B(n227), .Z(n373) );
  XNOR U381 ( .A(n1309), .B(n373), .Z(n3730) );
  XNOR U382 ( .A(in[1446]), .B(n3730), .Z(n2828) );
  NAND U383 ( .A(n2831), .B(n2828), .Z(n228) );
  XNOR U384 ( .A(n2550), .B(n228), .Z(out[100]) );
  XOR U385 ( .A(in[1396]), .B(in[116]), .Z(n230) );
  XNOR U386 ( .A(in[1076]), .B(in[756]), .Z(n229) );
  XNOR U387 ( .A(n230), .B(n229), .Z(n231) );
  XOR U388 ( .A(in[436]), .B(n231), .Z(n1428) );
  XOR U389 ( .A(in[1525]), .B(in[565]), .Z(n233) );
  XNOR U390 ( .A(in[885]), .B(in[245]), .Z(n232) );
  XNOR U391 ( .A(n233), .B(n232), .Z(n234) );
  XOR U392 ( .A(in[1205]), .B(n234), .Z(n1370) );
  XNOR U393 ( .A(n1428), .B(n1370), .Z(n3794) );
  XNOR U394 ( .A(in[181]), .B(n3794), .Z(n1342) );
  XOR U395 ( .A(in[341]), .B(in[661]), .Z(n236) );
  XNOR U396 ( .A(in[21]), .B(in[1301]), .Z(n235) );
  XNOR U397 ( .A(n236), .B(n235), .Z(n237) );
  XOR U398 ( .A(in[981]), .B(n237), .Z(n1251) );
  XOR U399 ( .A(in[150]), .B(in[1430]), .Z(n239) );
  XNOR U400 ( .A(in[1110]), .B(in[790]), .Z(n238) );
  XNOR U401 ( .A(n239), .B(n238), .Z(n240) );
  XNOR U402 ( .A(in[470]), .B(n240), .Z(n548) );
  XNOR U403 ( .A(n1251), .B(n548), .Z(n4129) );
  XNOR U404 ( .A(in[1366]), .B(n4129), .Z(n1737) );
  XOR U405 ( .A(in[1374]), .B(in[734]), .Z(n242) );
  XNOR U406 ( .A(in[94]), .B(in[414]), .Z(n241) );
  XNOR U407 ( .A(n242), .B(n241), .Z(n243) );
  XOR U408 ( .A(in[1054]), .B(n243), .Z(n916) );
  XOR U409 ( .A(in[1565]), .B(in[605]), .Z(n245) );
  XNOR U410 ( .A(in[925]), .B(in[285]), .Z(n244) );
  XNOR U411 ( .A(n245), .B(n244), .Z(n246) );
  XOR U412 ( .A(in[1245]), .B(n246), .Z(n650) );
  XNOR U413 ( .A(n916), .B(n650), .Z(n3904) );
  XNOR U414 ( .A(in[990]), .B(n3904), .Z(n1734) );
  NAND U415 ( .A(n1737), .B(n1734), .Z(n247) );
  XNOR U416 ( .A(n1342), .B(n247), .Z(out[1010]) );
  XOR U417 ( .A(in[1526]), .B(in[566]), .Z(n249) );
  XNOR U418 ( .A(in[886]), .B(in[246]), .Z(n248) );
  XNOR U419 ( .A(n249), .B(n248), .Z(n250) );
  XOR U420 ( .A(in[1206]), .B(n250), .Z(n1374) );
  XOR U421 ( .A(in[1397]), .B(in[117]), .Z(n252) );
  XNOR U422 ( .A(in[1077]), .B(in[757]), .Z(n251) );
  XNOR U423 ( .A(n252), .B(n251), .Z(n253) );
  XOR U424 ( .A(in[437]), .B(n253), .Z(n1432) );
  XNOR U425 ( .A(n1374), .B(n1432), .Z(n3804) );
  XNOR U426 ( .A(in[182]), .B(n3804), .Z(n1346) );
  XOR U427 ( .A(in[151]), .B(in[1431]), .Z(n255) );
  XNOR U428 ( .A(in[1111]), .B(in[791]), .Z(n254) );
  XNOR U429 ( .A(n255), .B(n254), .Z(n256) );
  XOR U430 ( .A(in[471]), .B(n256), .Z(n563) );
  XOR U431 ( .A(in[342]), .B(in[662]), .Z(n258) );
  XNOR U432 ( .A(in[22]), .B(in[1302]), .Z(n257) );
  XNOR U433 ( .A(n258), .B(n257), .Z(n259) );
  XNOR U434 ( .A(in[982]), .B(n259), .Z(n1254) );
  XNOR U435 ( .A(n563), .B(n1254), .Z(n4132) );
  XNOR U436 ( .A(in[1367]), .B(n4132), .Z(n1741) );
  XOR U437 ( .A(in[1375]), .B(in[735]), .Z(n261) );
  XNOR U438 ( .A(in[95]), .B(in[415]), .Z(n260) );
  XNOR U439 ( .A(n261), .B(n260), .Z(n262) );
  XOR U440 ( .A(in[1055]), .B(n262), .Z(n929) );
  XOR U441 ( .A(in[1566]), .B(in[606]), .Z(n264) );
  XNOR U442 ( .A(in[926]), .B(in[286]), .Z(n263) );
  XNOR U443 ( .A(n264), .B(n263), .Z(n265) );
  XOR U444 ( .A(in[1246]), .B(n265), .Z(n665) );
  XNOR U445 ( .A(n929), .B(n665), .Z(n3906) );
  XNOR U446 ( .A(in[991]), .B(n3906), .Z(n1738) );
  NAND U447 ( .A(n1741), .B(n1738), .Z(n266) );
  XNOR U448 ( .A(n1346), .B(n266), .Z(out[1011]) );
  XOR U449 ( .A(in[1527]), .B(in[567]), .Z(n268) );
  XNOR U450 ( .A(in[887]), .B(in[247]), .Z(n267) );
  XNOR U451 ( .A(n268), .B(n267), .Z(n269) );
  XOR U452 ( .A(in[1207]), .B(n269), .Z(n1378) );
  XOR U453 ( .A(in[1398]), .B(in[118]), .Z(n271) );
  XNOR U454 ( .A(in[1078]), .B(in[758]), .Z(n270) );
  XNOR U455 ( .A(n271), .B(n270), .Z(n272) );
  XOR U456 ( .A(in[438]), .B(n272), .Z(n1436) );
  XNOR U457 ( .A(n1378), .B(n1436), .Z(n3808) );
  XNOR U458 ( .A(in[183]), .B(n3808), .Z(n1351) );
  XOR U459 ( .A(in[343]), .B(in[663]), .Z(n274) );
  XNOR U460 ( .A(in[23]), .B(in[1303]), .Z(n273) );
  XNOR U461 ( .A(n274), .B(n273), .Z(n275) );
  XOR U462 ( .A(in[983]), .B(n275), .Z(n1257) );
  XOR U463 ( .A(in[152]), .B(in[1432]), .Z(n277) );
  XNOR U464 ( .A(in[1112]), .B(in[792]), .Z(n276) );
  XNOR U465 ( .A(n277), .B(n276), .Z(n278) );
  XNOR U466 ( .A(in[472]), .B(n278), .Z(n589) );
  XNOR U467 ( .A(n1257), .B(n589), .Z(n4135) );
  XNOR U468 ( .A(in[1368]), .B(n4135), .Z(n1745) );
  XOR U469 ( .A(in[1376]), .B(in[736]), .Z(n280) );
  XNOR U470 ( .A(in[96]), .B(in[416]), .Z(n279) );
  XNOR U471 ( .A(n280), .B(n279), .Z(n281) );
  XOR U472 ( .A(in[1056]), .B(n281), .Z(n944) );
  XOR U473 ( .A(in[1567]), .B(in[607]), .Z(n283) );
  XNOR U474 ( .A(in[927]), .B(in[287]), .Z(n282) );
  XNOR U475 ( .A(n283), .B(n282), .Z(n284) );
  XOR U476 ( .A(in[1247]), .B(n284), .Z(n680) );
  XNOR U477 ( .A(n944), .B(n680), .Z(n3908) );
  XNOR U478 ( .A(in[992]), .B(n3908), .Z(n1742) );
  NAND U479 ( .A(n1745), .B(n1742), .Z(n285) );
  XNOR U480 ( .A(n1351), .B(n285), .Z(out[1012]) );
  XOR U481 ( .A(in[1528]), .B(in[568]), .Z(n287) );
  XNOR U482 ( .A(in[888]), .B(in[248]), .Z(n286) );
  XNOR U483 ( .A(n287), .B(n286), .Z(n288) );
  XOR U484 ( .A(in[1208]), .B(n288), .Z(n1382) );
  XOR U485 ( .A(in[1399]), .B(in[119]), .Z(n290) );
  XNOR U486 ( .A(in[1079]), .B(in[759]), .Z(n289) );
  XNOR U487 ( .A(n290), .B(n289), .Z(n291) );
  XOR U488 ( .A(in[439]), .B(n291), .Z(n1440) );
  XNOR U489 ( .A(n1382), .B(n1440), .Z(n3812) );
  XNOR U490 ( .A(in[184]), .B(n3812), .Z(n1355) );
  XOR U491 ( .A(in[153]), .B(in[1433]), .Z(n293) );
  XNOR U492 ( .A(in[1113]), .B(in[793]), .Z(n292) );
  XNOR U493 ( .A(n293), .B(n292), .Z(n294) );
  XOR U494 ( .A(in[473]), .B(n294), .Z(n604) );
  XOR U495 ( .A(in[344]), .B(in[664]), .Z(n296) );
  XNOR U496 ( .A(in[24]), .B(in[1304]), .Z(n295) );
  XNOR U497 ( .A(n296), .B(n295), .Z(n297) );
  XNOR U498 ( .A(in[984]), .B(n297), .Z(n1260) );
  XNOR U499 ( .A(n604), .B(n1260), .Z(n4138) );
  XNOR U500 ( .A(in[1369]), .B(n4138), .Z(n1749) );
  XOR U501 ( .A(in[1377]), .B(in[737]), .Z(n299) );
  XNOR U502 ( .A(in[97]), .B(in[417]), .Z(n298) );
  XNOR U503 ( .A(n299), .B(n298), .Z(n300) );
  XOR U504 ( .A(in[1057]), .B(n300), .Z(n959) );
  XOR U505 ( .A(in[1568]), .B(in[608]), .Z(n302) );
  XNOR U506 ( .A(in[928]), .B(in[288]), .Z(n301) );
  XNOR U507 ( .A(n302), .B(n301), .Z(n303) );
  XOR U508 ( .A(in[1248]), .B(n303), .Z(n695) );
  XNOR U509 ( .A(n959), .B(n695), .Z(n3910) );
  XNOR U510 ( .A(in[993]), .B(n3910), .Z(n1746) );
  NAND U511 ( .A(n1749), .B(n1746), .Z(n304) );
  XNOR U512 ( .A(n1355), .B(n304), .Z(out[1013]) );
  XOR U513 ( .A(in[1529]), .B(in[569]), .Z(n306) );
  XNOR U514 ( .A(in[889]), .B(in[249]), .Z(n305) );
  XNOR U515 ( .A(n306), .B(n305), .Z(n307) );
  XOR U516 ( .A(in[1209]), .B(n307), .Z(n1386) );
  XOR U517 ( .A(in[1400]), .B(in[120]), .Z(n309) );
  XNOR U518 ( .A(in[1080]), .B(in[760]), .Z(n308) );
  XNOR U519 ( .A(n309), .B(n308), .Z(n310) );
  XOR U520 ( .A(in[440]), .B(n310), .Z(n1444) );
  XNOR U521 ( .A(n1386), .B(n1444), .Z(n3816) );
  XNOR U522 ( .A(in[185]), .B(n3816), .Z(n1359) );
  XOR U523 ( .A(in[345]), .B(in[665]), .Z(n312) );
  XNOR U524 ( .A(in[25]), .B(in[1305]), .Z(n311) );
  XNOR U525 ( .A(n312), .B(n311), .Z(n313) );
  XOR U526 ( .A(in[985]), .B(n313), .Z(n1263) );
  XOR U527 ( .A(in[154]), .B(in[1434]), .Z(n315) );
  XNOR U528 ( .A(in[1114]), .B(in[794]), .Z(n314) );
  XNOR U529 ( .A(n315), .B(n314), .Z(n316) );
  XNOR U530 ( .A(in[474]), .B(n316), .Z(n619) );
  XNOR U531 ( .A(n1263), .B(n619), .Z(n4141) );
  XNOR U532 ( .A(in[1370]), .B(n4141), .Z(n1754) );
  XOR U533 ( .A(in[1569]), .B(in[609]), .Z(n318) );
  XNOR U534 ( .A(in[929]), .B(in[289]), .Z(n317) );
  XNOR U535 ( .A(n318), .B(n317), .Z(n319) );
  XOR U536 ( .A(in[1249]), .B(n319), .Z(n710) );
  XOR U537 ( .A(in[1378]), .B(in[738]), .Z(n321) );
  XNOR U538 ( .A(in[98]), .B(in[418]), .Z(n320) );
  XNOR U539 ( .A(n321), .B(n320), .Z(n322) );
  XOR U540 ( .A(in[1058]), .B(n322), .Z(n974) );
  XNOR U541 ( .A(n710), .B(n974), .Z(n3912) );
  XNOR U542 ( .A(in[994]), .B(n3912), .Z(n1751) );
  NAND U543 ( .A(n1754), .B(n1751), .Z(n323) );
  XNOR U544 ( .A(n1359), .B(n323), .Z(out[1014]) );
  XOR U545 ( .A(in[1401]), .B(in[121]), .Z(n325) );
  XNOR U546 ( .A(in[1081]), .B(in[761]), .Z(n324) );
  XNOR U547 ( .A(n325), .B(n324), .Z(n326) );
  XOR U548 ( .A(in[441]), .B(n326), .Z(n1448) );
  XNOR U549 ( .A(n327), .B(n1448), .Z(n3538) );
  XNOR U550 ( .A(in[186]), .B(n3538), .Z(n1363) );
  XOR U551 ( .A(in[155]), .B(in[1435]), .Z(n329) );
  XNOR U552 ( .A(in[1115]), .B(in[795]), .Z(n328) );
  XNOR U553 ( .A(n329), .B(n328), .Z(n330) );
  XOR U554 ( .A(in[475]), .B(n330), .Z(n634) );
  XOR U555 ( .A(in[346]), .B(in[666]), .Z(n332) );
  XNOR U556 ( .A(in[26]), .B(in[1306]), .Z(n331) );
  XNOR U557 ( .A(n332), .B(n331), .Z(n333) );
  XNOR U558 ( .A(in[986]), .B(n333), .Z(n1266) );
  XNOR U559 ( .A(n634), .B(n1266), .Z(n4148) );
  XNOR U560 ( .A(in[1371]), .B(n4148), .Z(n1758) );
  XOR U561 ( .A(in[1379]), .B(in[739]), .Z(n335) );
  XNOR U562 ( .A(in[99]), .B(in[419]), .Z(n334) );
  XNOR U563 ( .A(n335), .B(n334), .Z(n336) );
  XNOR U564 ( .A(in[1059]), .B(n336), .Z(n989) );
  XNOR U565 ( .A(n337), .B(n989), .Z(n3914) );
  XNOR U566 ( .A(in[995]), .B(n3914), .Z(n1755) );
  NAND U567 ( .A(n1758), .B(n1755), .Z(n338) );
  XNOR U568 ( .A(n1363), .B(n338), .Z(out[1015]) );
  XOR U569 ( .A(in[1402]), .B(in[122]), .Z(n340) );
  XNOR U570 ( .A(in[1082]), .B(in[762]), .Z(n339) );
  XNOR U571 ( .A(n340), .B(n339), .Z(n341) );
  XOR U572 ( .A(in[442]), .B(n341), .Z(n1452) );
  XOR U573 ( .A(in[1531]), .B(in[571]), .Z(n343) );
  XNOR U574 ( .A(in[1211]), .B(in[251]), .Z(n342) );
  XNOR U575 ( .A(n343), .B(n342), .Z(n344) );
  XOR U576 ( .A(in[891]), .B(n344), .Z(n416) );
  XNOR U577 ( .A(n1452), .B(n416), .Z(n3542) );
  XNOR U578 ( .A(in[187]), .B(n3542), .Z(n1367) );
  XOR U579 ( .A(in[156]), .B(in[1436]), .Z(n346) );
  XNOR U580 ( .A(in[1116]), .B(in[796]), .Z(n345) );
  XNOR U581 ( .A(n346), .B(n345), .Z(n347) );
  XOR U582 ( .A(in[476]), .B(n347), .Z(n649) );
  XOR U583 ( .A(in[347]), .B(in[667]), .Z(n349) );
  XNOR U584 ( .A(in[27]), .B(in[1307]), .Z(n348) );
  XNOR U585 ( .A(n349), .B(n348), .Z(n350) );
  XNOR U586 ( .A(in[987]), .B(n350), .Z(n1269) );
  XNOR U587 ( .A(n649), .B(n1269), .Z(n4151) );
  XNOR U588 ( .A(in[1372]), .B(n4151), .Z(n1762) );
  XOR U589 ( .A(in[1060]), .B(in[420]), .Z(n352) );
  XNOR U590 ( .A(in[740]), .B(in[1380]), .Z(n351) );
  XNOR U591 ( .A(n352), .B(n351), .Z(n353) );
  XOR U592 ( .A(in[100]), .B(n353), .Z(n1004) );
  XOR U593 ( .A(in[1571]), .B(in[611]), .Z(n355) );
  XNOR U594 ( .A(in[931]), .B(in[291]), .Z(n354) );
  XNOR U595 ( .A(n355), .B(n354), .Z(n356) );
  XOR U596 ( .A(in[1251]), .B(n356), .Z(n420) );
  XNOR U597 ( .A(n1004), .B(n420), .Z(n3916) );
  XNOR U598 ( .A(in[996]), .B(n3916), .Z(n1759) );
  NAND U599 ( .A(n1762), .B(n1759), .Z(n357) );
  XNOR U600 ( .A(n1367), .B(n357), .Z(out[1016]) );
  XOR U601 ( .A(in[1403]), .B(in[123]), .Z(n359) );
  XNOR U602 ( .A(in[1083]), .B(in[763]), .Z(n358) );
  XNOR U603 ( .A(n359), .B(n358), .Z(n360) );
  XOR U604 ( .A(in[443]), .B(n360), .Z(n1456) );
  XOR U605 ( .A(in[1532]), .B(in[572]), .Z(n362) );
  XNOR U606 ( .A(in[1212]), .B(in[252]), .Z(n361) );
  XNOR U607 ( .A(n362), .B(n361), .Z(n363) );
  XOR U608 ( .A(in[892]), .B(n363), .Z(n581) );
  XNOR U609 ( .A(n1456), .B(n581), .Z(n3546) );
  XNOR U610 ( .A(in[188]), .B(n3546), .Z(n1371) );
  XOR U611 ( .A(in[157]), .B(in[1437]), .Z(n365) );
  XNOR U612 ( .A(in[1117]), .B(in[797]), .Z(n364) );
  XNOR U613 ( .A(n365), .B(n364), .Z(n366) );
  XOR U614 ( .A(in[477]), .B(n366), .Z(n664) );
  XOR U615 ( .A(in[348]), .B(in[668]), .Z(n368) );
  XNOR U616 ( .A(in[28]), .B(in[1308]), .Z(n367) );
  XNOR U617 ( .A(n368), .B(n367), .Z(n369) );
  XNOR U618 ( .A(in[988]), .B(n369), .Z(n1272) );
  XNOR U619 ( .A(n664), .B(n1272), .Z(n4154) );
  XNOR U620 ( .A(in[1373]), .B(n4154), .Z(n1766) );
  XOR U621 ( .A(in[1572]), .B(in[612]), .Z(n371) );
  XNOR U622 ( .A(in[932]), .B(in[292]), .Z(n370) );
  XNOR U623 ( .A(n371), .B(n370), .Z(n372) );
  XOR U624 ( .A(in[1252]), .B(n372), .Z(n583) );
  XNOR U625 ( .A(n373), .B(n583), .Z(n3918) );
  XNOR U626 ( .A(in[997]), .B(n3918), .Z(n1763) );
  NAND U627 ( .A(n1766), .B(n1763), .Z(n374) );
  XNOR U628 ( .A(n1371), .B(n374), .Z(out[1017]) );
  XOR U629 ( .A(in[1404]), .B(in[124]), .Z(n376) );
  XNOR U630 ( .A(in[1084]), .B(in[764]), .Z(n375) );
  XNOR U631 ( .A(n376), .B(n375), .Z(n377) );
  XOR U632 ( .A(in[444]), .B(n377), .Z(n1460) );
  XOR U633 ( .A(in[1533]), .B(in[573]), .Z(n379) );
  XNOR U634 ( .A(in[1213]), .B(in[253]), .Z(n378) );
  XNOR U635 ( .A(n379), .B(n378), .Z(n380) );
  XOR U636 ( .A(in[893]), .B(n380), .Z(n740) );
  XNOR U637 ( .A(n1460), .B(n740), .Z(n3550) );
  XNOR U638 ( .A(in[189]), .B(n3550), .Z(n1375) );
  XOR U639 ( .A(in[158]), .B(in[1438]), .Z(n382) );
  XNOR U640 ( .A(in[1118]), .B(in[798]), .Z(n381) );
  XNOR U641 ( .A(n382), .B(n381), .Z(n383) );
  XOR U642 ( .A(in[478]), .B(n383), .Z(n679) );
  XOR U643 ( .A(in[349]), .B(in[669]), .Z(n385) );
  XNOR U644 ( .A(in[29]), .B(in[1309]), .Z(n384) );
  XNOR U645 ( .A(n385), .B(n384), .Z(n386) );
  XNOR U646 ( .A(in[989]), .B(n386), .Z(n1276) );
  XNOR U647 ( .A(n679), .B(n1276), .Z(n4157) );
  XNOR U648 ( .A(in[1374]), .B(n4157), .Z(n1770) );
  XOR U649 ( .A(in[1062]), .B(in[422]), .Z(n388) );
  XNOR U650 ( .A(in[742]), .B(in[1382]), .Z(n387) );
  XNOR U651 ( .A(n388), .B(n387), .Z(n389) );
  XOR U652 ( .A(in[102]), .B(n389), .Z(n424) );
  XOR U653 ( .A(in[1573]), .B(in[613]), .Z(n391) );
  XNOR U654 ( .A(in[933]), .B(in[293]), .Z(n390) );
  XNOR U655 ( .A(n391), .B(n390), .Z(n392) );
  XOR U656 ( .A(in[1253]), .B(n392), .Z(n742) );
  XNOR U657 ( .A(n424), .B(n742), .Z(n3924) );
  XNOR U658 ( .A(in[998]), .B(n3924), .Z(n1767) );
  NAND U659 ( .A(n1770), .B(n1767), .Z(n393) );
  XNOR U660 ( .A(n1375), .B(n393), .Z(out[1018]) );
  XOR U661 ( .A(in[1405]), .B(in[125]), .Z(n395) );
  XNOR U662 ( .A(in[1085]), .B(in[765]), .Z(n394) );
  XNOR U663 ( .A(n395), .B(n394), .Z(n396) );
  XOR U664 ( .A(in[445]), .B(n396), .Z(n1464) );
  XOR U665 ( .A(in[1534]), .B(in[894]), .Z(n398) );
  XNOR U666 ( .A(in[574]), .B(in[1214]), .Z(n397) );
  XNOR U667 ( .A(n398), .B(n397), .Z(n399) );
  XOR U668 ( .A(in[254]), .B(n399), .Z(n877) );
  XNOR U669 ( .A(n1464), .B(n877), .Z(n3554) );
  XNOR U670 ( .A(in[190]), .B(n3554), .Z(n1379) );
  XOR U671 ( .A(in[1439]), .B(in[479]), .Z(n401) );
  XNOR U672 ( .A(in[799]), .B(in[159]), .Z(n400) );
  XNOR U673 ( .A(n401), .B(n400), .Z(n402) );
  XOR U674 ( .A(in[1119]), .B(n402), .Z(n694) );
  XOR U675 ( .A(in[350]), .B(in[670]), .Z(n404) );
  XNOR U676 ( .A(in[30]), .B(in[1310]), .Z(n403) );
  XNOR U677 ( .A(n404), .B(n403), .Z(n405) );
  XNOR U678 ( .A(in[990]), .B(n405), .Z(n1279) );
  XNOR U679 ( .A(n694), .B(n1279), .Z(n4160) );
  XNOR U680 ( .A(in[1375]), .B(n4160), .Z(n1774) );
  XOR U681 ( .A(in[1063]), .B(in[423]), .Z(n407) );
  XNOR U682 ( .A(in[743]), .B(in[1383]), .Z(n406) );
  XNOR U683 ( .A(n407), .B(n406), .Z(n408) );
  XOR U684 ( .A(in[103]), .B(n408), .Z(n587) );
  XOR U685 ( .A(in[1574]), .B(in[614]), .Z(n410) );
  XNOR U686 ( .A(in[934]), .B(in[294]), .Z(n409) );
  XNOR U687 ( .A(n410), .B(n409), .Z(n411) );
  XOR U688 ( .A(in[1254]), .B(n411), .Z(n786) );
  XNOR U689 ( .A(n587), .B(n786), .Z(n3926) );
  XNOR U690 ( .A(in[999]), .B(n3926), .Z(n1771) );
  NAND U691 ( .A(n1774), .B(n1771), .Z(n412) );
  XNOR U692 ( .A(n1379), .B(n412), .Z(out[1019]) );
  XOR U693 ( .A(in[1340]), .B(in[60]), .Z(n414) );
  XNOR U694 ( .A(in[700]), .B(in[380]), .Z(n413) );
  XNOR U695 ( .A(n414), .B(n413), .Z(n415) );
  XOR U696 ( .A(in[1020]), .B(n415), .Z(n871) );
  XNOR U697 ( .A(n416), .B(n871), .Z(n3596) );
  XNOR U698 ( .A(in[636]), .B(n3596), .Z(n2552) );
  XOR U699 ( .A(in[162]), .B(in[1442]), .Z(n418) );
  XNOR U700 ( .A(in[802]), .B(in[1122]), .Z(n417) );
  XNOR U701 ( .A(n418), .B(n417), .Z(n419) );
  XNOR U702 ( .A(in[482]), .B(n419), .Z(n471) );
  XNOR U703 ( .A(n420), .B(n471), .Z(n3693) );
  XNOR U704 ( .A(in[227]), .B(n3693), .Z(n2845) );
  XOR U705 ( .A(in[1511]), .B(in[551]), .Z(n422) );
  XNOR U706 ( .A(in[871]), .B(in[231]), .Z(n421) );
  XNOR U707 ( .A(n422), .B(n421), .Z(n423) );
  XOR U708 ( .A(in[1191]), .B(n423), .Z(n1313) );
  XNOR U709 ( .A(n424), .B(n1313), .Z(n3734) );
  XNOR U710 ( .A(in[1447]), .B(n3734), .Z(n2842) );
  NAND U711 ( .A(n2845), .B(n2842), .Z(n425) );
  XNOR U712 ( .A(n2552), .B(n425), .Z(out[101]) );
  XOR U713 ( .A(in[1406]), .B(in[126]), .Z(n427) );
  XNOR U714 ( .A(in[1086]), .B(in[766]), .Z(n426) );
  XNOR U715 ( .A(n427), .B(n426), .Z(n428) );
  XOR U716 ( .A(in[446]), .B(n428), .Z(n1469) );
  XOR U717 ( .A(in[1535]), .B(in[575]), .Z(n430) );
  XNOR U718 ( .A(in[895]), .B(in[255]), .Z(n429) );
  XNOR U719 ( .A(n430), .B(n429), .Z(n431) );
  XOR U720 ( .A(in[1215]), .B(n431), .Z(n1024) );
  XNOR U721 ( .A(n1469), .B(n1024), .Z(n3558) );
  XNOR U722 ( .A(in[191]), .B(n3558), .Z(n1383) );
  XOR U723 ( .A(in[1440]), .B(in[480]), .Z(n433) );
  XNOR U724 ( .A(in[800]), .B(in[160]), .Z(n432) );
  XNOR U725 ( .A(n433), .B(n432), .Z(n434) );
  XOR U726 ( .A(in[1120]), .B(n434), .Z(n709) );
  XOR U727 ( .A(in[351]), .B(in[671]), .Z(n436) );
  XNOR U728 ( .A(in[31]), .B(in[1311]), .Z(n435) );
  XNOR U729 ( .A(n436), .B(n435), .Z(n437) );
  XNOR U730 ( .A(in[991]), .B(n437), .Z(n1282) );
  XNOR U731 ( .A(n709), .B(n1282), .Z(n4163) );
  XNOR U732 ( .A(in[1376]), .B(n4163), .Z(n1778) );
  XOR U733 ( .A(in[1064]), .B(in[424]), .Z(n439) );
  XNOR U734 ( .A(in[744]), .B(in[1384]), .Z(n438) );
  XNOR U735 ( .A(n439), .B(n438), .Z(n440) );
  XOR U736 ( .A(in[104]), .B(n440), .Z(n746) );
  XOR U737 ( .A(in[1575]), .B(in[615]), .Z(n442) );
  XNOR U738 ( .A(in[935]), .B(in[295]), .Z(n441) );
  XNOR U739 ( .A(n442), .B(n441), .Z(n443) );
  XOR U740 ( .A(in[1255]), .B(n443), .Z(n799) );
  XNOR U741 ( .A(n746), .B(n799), .Z(n3928) );
  XNOR U742 ( .A(in[1000]), .B(n3928), .Z(n1775) );
  NAND U743 ( .A(n1778), .B(n1775), .Z(n444) );
  XNOR U744 ( .A(n1383), .B(n444), .Z(out[1020]) );
  XOR U745 ( .A(in[1407]), .B(in[127]), .Z(n446) );
  XNOR U746 ( .A(in[1087]), .B(in[767]), .Z(n445) );
  XNOR U747 ( .A(n446), .B(n445), .Z(n447) );
  XOR U748 ( .A(in[447]), .B(n447), .Z(n1472) );
  XOR U749 ( .A(in[1472]), .B(in[512]), .Z(n449) );
  XNOR U750 ( .A(in[832]), .B(in[192]), .Z(n448) );
  XNOR U751 ( .A(n449), .B(n448), .Z(n450) );
  XOR U752 ( .A(in[1152]), .B(n450), .Z(n1091) );
  XNOR U753 ( .A(n1472), .B(n1091), .Z(n3562) );
  XNOR U754 ( .A(in[128]), .B(n3562), .Z(n1387) );
  XOR U755 ( .A(in[352]), .B(in[672]), .Z(n452) );
  XNOR U756 ( .A(in[32]), .B(in[1312]), .Z(n451) );
  XNOR U757 ( .A(n452), .B(n451), .Z(n453) );
  XNOR U758 ( .A(in[992]), .B(n453), .Z(n1285) );
  XNOR U759 ( .A(n454), .B(n1285), .Z(n4166) );
  XNOR U760 ( .A(in[1377]), .B(n4166), .Z(n1782) );
  XOR U761 ( .A(in[1065]), .B(in[425]), .Z(n456) );
  XNOR U762 ( .A(in[745]), .B(in[1385]), .Z(n455) );
  XNOR U763 ( .A(n456), .B(n455), .Z(n457) );
  XOR U764 ( .A(in[105]), .B(n457), .Z(n881) );
  XOR U765 ( .A(in[1576]), .B(in[616]), .Z(n459) );
  XNOR U766 ( .A(in[936]), .B(in[296]), .Z(n458) );
  XNOR U767 ( .A(n459), .B(n458), .Z(n460) );
  XOR U768 ( .A(in[1256]), .B(n460), .Z(n812) );
  XNOR U769 ( .A(n881), .B(n812), .Z(n3930) );
  XNOR U770 ( .A(in[1001]), .B(n3930), .Z(n1779) );
  NAND U771 ( .A(n1782), .B(n1779), .Z(n461) );
  XNOR U772 ( .A(n1387), .B(n461), .Z(out[1021]) );
  XOR U773 ( .A(in[1344]), .B(in[64]), .Z(n463) );
  XNOR U774 ( .A(in[1024]), .B(in[384]), .Z(n462) );
  XNOR U775 ( .A(n463), .B(n462), .Z(n464) );
  XOR U776 ( .A(in[704]), .B(n464), .Z(n1477) );
  XOR U777 ( .A(in[1473]), .B(in[513]), .Z(n466) );
  XNOR U778 ( .A(in[833]), .B(in[193]), .Z(n465) );
  XNOR U779 ( .A(n466), .B(n465), .Z(n467) );
  XOR U780 ( .A(in[1153]), .B(n467), .Z(n1144) );
  XNOR U781 ( .A(n1477), .B(n1144), .Z(n3566) );
  XNOR U782 ( .A(in[129]), .B(n3566), .Z(n1390) );
  XOR U783 ( .A(in[353]), .B(in[673]), .Z(n469) );
  XNOR U784 ( .A(in[33]), .B(in[1313]), .Z(n468) );
  XNOR U785 ( .A(n469), .B(n468), .Z(n470) );
  XOR U786 ( .A(in[993]), .B(n470), .Z(n1288) );
  XNOR U787 ( .A(n1288), .B(n471), .Z(n4169) );
  XNOR U788 ( .A(in[1378]), .B(n4169), .Z(n1786) );
  XOR U789 ( .A(in[1577]), .B(in[617]), .Z(n473) );
  XNOR U790 ( .A(in[937]), .B(in[297]), .Z(n472) );
  XNOR U791 ( .A(n473), .B(n472), .Z(n474) );
  XOR U792 ( .A(in[1257]), .B(n474), .Z(n825) );
  XNOR U793 ( .A(n475), .B(n825), .Z(n3932) );
  XNOR U794 ( .A(in[1002]), .B(n3932), .Z(n1783) );
  NAND U795 ( .A(n1786), .B(n1783), .Z(n476) );
  XNOR U796 ( .A(n1390), .B(n476), .Z(out[1022]) );
  XOR U797 ( .A(n3570), .B(in[130]), .Z(n1392) );
  XOR U798 ( .A(in[163]), .B(in[1443]), .Z(n478) );
  XNOR U799 ( .A(in[803]), .B(in[1123]), .Z(n477) );
  XNOR U800 ( .A(n478), .B(n477), .Z(n479) );
  XOR U801 ( .A(in[483]), .B(n479), .Z(n582) );
  XOR U802 ( .A(in[354]), .B(in[674]), .Z(n481) );
  XNOR U803 ( .A(in[34]), .B(in[1314]), .Z(n480) );
  XNOR U804 ( .A(n481), .B(n480), .Z(n482) );
  XNOR U805 ( .A(in[994]), .B(n482), .Z(n1291) );
  XNOR U806 ( .A(n582), .B(n1291), .Z(n4172) );
  XNOR U807 ( .A(in[1379]), .B(n4172), .Z(n1790) );
  XOR U808 ( .A(in[1578]), .B(in[618]), .Z(n484) );
  XNOR U809 ( .A(in[938]), .B(in[298]), .Z(n483) );
  XNOR U810 ( .A(n484), .B(n483), .Z(n485) );
  XOR U811 ( .A(in[1258]), .B(n485), .Z(n838) );
  XNOR U812 ( .A(n486), .B(n838), .Z(n3934) );
  XNOR U813 ( .A(in[1003]), .B(n3934), .Z(n1787) );
  NAND U814 ( .A(n1790), .B(n1787), .Z(n487) );
  XNOR U815 ( .A(n1392), .B(n487), .Z(out[1023]) );
  XNOR U816 ( .A(n489), .B(n488), .Z(n3625) );
  XNOR U817 ( .A(in[531]), .B(n3625), .Z(n1396) );
  XOR U818 ( .A(in[1346]), .B(in[66]), .Z(n491) );
  XNOR U819 ( .A(in[1026]), .B(in[386]), .Z(n490) );
  XNOR U820 ( .A(n491), .B(n490), .Z(n492) );
  XOR U821 ( .A(in[706]), .B(n492), .Z(n1485) );
  XOR U822 ( .A(in[1475]), .B(in[515]), .Z(n494) );
  XNOR U823 ( .A(in[835]), .B(in[195]), .Z(n493) );
  XNOR U824 ( .A(n494), .B(n493), .Z(n495) );
  XNOR U825 ( .A(in[1155]), .B(n495), .Z(n1196) );
  XNOR U826 ( .A(n1485), .B(n1196), .Z(n3574) );
  XNOR U827 ( .A(in[131]), .B(n3574), .Z(n4631) );
  XOR U828 ( .A(in[35]), .B(in[675]), .Z(n497) );
  XNOR U829 ( .A(in[355]), .B(in[1315]), .Z(n496) );
  XNOR U830 ( .A(n497), .B(n496), .Z(n498) );
  XOR U831 ( .A(in[995]), .B(n498), .Z(n1294) );
  XOR U832 ( .A(in[164]), .B(in[1444]), .Z(n500) );
  XNOR U833 ( .A(in[804]), .B(in[1124]), .Z(n499) );
  XNOR U834 ( .A(n500), .B(n499), .Z(n501) );
  XOR U835 ( .A(in[484]), .B(n501), .Z(n741) );
  XNOR U836 ( .A(n1294), .B(n741), .Z(n4175) );
  XNOR U837 ( .A(in[1380]), .B(n4175), .Z(n4628) );
  NAND U838 ( .A(n4631), .B(n4628), .Z(n502) );
  XNOR U839 ( .A(n1396), .B(n502), .Z(out[1024]) );
  XOR U840 ( .A(n504), .B(n503), .Z(n3629) );
  XNOR U841 ( .A(in[532]), .B(n3629), .Z(n1400) );
  XOR U842 ( .A(in[1347]), .B(in[67]), .Z(n506) );
  XNOR U843 ( .A(in[1027]), .B(in[387]), .Z(n505) );
  XNOR U844 ( .A(n506), .B(n505), .Z(n507) );
  XOR U845 ( .A(in[707]), .B(n507), .Z(n1489) );
  XOR U846 ( .A(in[1476]), .B(in[516]), .Z(n509) );
  XNOR U847 ( .A(in[836]), .B(in[196]), .Z(n508) );
  XNOR U848 ( .A(n509), .B(n508), .Z(n510) );
  XNOR U849 ( .A(in[1156]), .B(n510), .Z(n1199) );
  XNOR U850 ( .A(n1489), .B(n1199), .Z(n3582) );
  XNOR U851 ( .A(in[132]), .B(n3582), .Z(n4635) );
  XOR U852 ( .A(in[1445]), .B(in[165]), .Z(n512) );
  XNOR U853 ( .A(in[805]), .B(in[1125]), .Z(n511) );
  XNOR U854 ( .A(n512), .B(n511), .Z(n513) );
  XOR U855 ( .A(in[485]), .B(n513), .Z(n785) );
  XOR U856 ( .A(in[36]), .B(in[676]), .Z(n515) );
  XNOR U857 ( .A(in[356]), .B(in[1316]), .Z(n514) );
  XNOR U858 ( .A(n515), .B(n514), .Z(n516) );
  XOR U859 ( .A(in[996]), .B(n516), .Z(n1297) );
  XNOR U860 ( .A(n785), .B(n1297), .Z(n4182) );
  XNOR U861 ( .A(in[1381]), .B(n4182), .Z(n4632) );
  NAND U862 ( .A(n4635), .B(n4632), .Z(n517) );
  XNOR U863 ( .A(n1400), .B(n517), .Z(out[1025]) );
  XNOR U864 ( .A(n519), .B(n518), .Z(n3633) );
  XNOR U865 ( .A(in[533]), .B(n3633), .Z(n1404) );
  XOR U866 ( .A(in[1348]), .B(in[68]), .Z(n521) );
  XNOR U867 ( .A(in[1028]), .B(in[388]), .Z(n520) );
  XNOR U868 ( .A(n521), .B(n520), .Z(n522) );
  XOR U869 ( .A(in[708]), .B(n522), .Z(n1493) );
  XOR U870 ( .A(in[1477]), .B(in[517]), .Z(n524) );
  XNOR U871 ( .A(in[837]), .B(in[197]), .Z(n523) );
  XNOR U872 ( .A(n524), .B(n523), .Z(n525) );
  XNOR U873 ( .A(in[1157]), .B(n525), .Z(n1202) );
  XNOR U874 ( .A(n1493), .B(n1202), .Z(n3586) );
  XNOR U875 ( .A(in[133]), .B(n3586), .Z(n4639) );
  XOR U876 ( .A(in[37]), .B(in[677]), .Z(n527) );
  XNOR U877 ( .A(in[357]), .B(in[1317]), .Z(n526) );
  XNOR U878 ( .A(n527), .B(n526), .Z(n528) );
  XOR U879 ( .A(in[997]), .B(n528), .Z(n1300) );
  XOR U880 ( .A(in[166]), .B(in[806]), .Z(n530) );
  XNOR U881 ( .A(in[1126]), .B(in[486]), .Z(n529) );
  XNOR U882 ( .A(n530), .B(n529), .Z(n531) );
  XOR U883 ( .A(in[1446]), .B(n531), .Z(n798) );
  XNOR U884 ( .A(n1300), .B(n798), .Z(n4185) );
  XNOR U885 ( .A(in[1382]), .B(n4185), .Z(n4636) );
  NAND U886 ( .A(n4639), .B(n4636), .Z(n532) );
  XNOR U887 ( .A(n1404), .B(n532), .Z(out[1026]) );
  XOR U888 ( .A(n534), .B(n533), .Z(n3637) );
  XNOR U889 ( .A(in[534]), .B(n3637), .Z(n1408) );
  XOR U890 ( .A(in[1349]), .B(in[69]), .Z(n536) );
  XNOR U891 ( .A(in[1029]), .B(in[389]), .Z(n535) );
  XNOR U892 ( .A(n536), .B(n535), .Z(n537) );
  XOR U893 ( .A(in[709]), .B(n537), .Z(n1497) );
  XOR U894 ( .A(in[1478]), .B(in[518]), .Z(n539) );
  XNOR U895 ( .A(in[838]), .B(in[198]), .Z(n538) );
  XNOR U896 ( .A(n539), .B(n538), .Z(n540) );
  XNOR U897 ( .A(in[1158]), .B(n540), .Z(n1205) );
  XNOR U898 ( .A(n1497), .B(n1205), .Z(n3590) );
  XNOR U899 ( .A(in[134]), .B(n3590), .Z(n4643) );
  XOR U900 ( .A(in[38]), .B(in[678]), .Z(n542) );
  XNOR U901 ( .A(in[358]), .B(in[1318]), .Z(n541) );
  XNOR U902 ( .A(n542), .B(n541), .Z(n543) );
  XOR U903 ( .A(in[998]), .B(n543), .Z(n1304) );
  XOR U904 ( .A(in[167]), .B(in[807]), .Z(n545) );
  XNOR U905 ( .A(in[1127]), .B(in[487]), .Z(n544) );
  XNOR U906 ( .A(n545), .B(n544), .Z(n546) );
  XOR U907 ( .A(in[1447]), .B(n546), .Z(n811) );
  XNOR U908 ( .A(n1304), .B(n811), .Z(n3964) );
  XNOR U909 ( .A(in[1383]), .B(n3964), .Z(n4640) );
  NAND U910 ( .A(n4643), .B(n4640), .Z(n547) );
  XNOR U911 ( .A(n1408), .B(n547), .Z(out[1027]) );
  XOR U912 ( .A(n549), .B(n548), .Z(n3641) );
  XNOR U913 ( .A(in[535]), .B(n3641), .Z(n1412) );
  XOR U914 ( .A(in[1350]), .B(in[70]), .Z(n551) );
  XNOR U915 ( .A(in[1030]), .B(in[390]), .Z(n550) );
  XNOR U916 ( .A(n551), .B(n550), .Z(n552) );
  XOR U917 ( .A(in[710]), .B(n552), .Z(n1501) );
  XOR U918 ( .A(in[199]), .B(in[1479]), .Z(n554) );
  XNOR U919 ( .A(in[1159]), .B(in[839]), .Z(n553) );
  XNOR U920 ( .A(n554), .B(n553), .Z(n555) );
  XNOR U921 ( .A(in[519]), .B(n555), .Z(n1208) );
  XNOR U922 ( .A(n1501), .B(n1208), .Z(n3594) );
  XNOR U923 ( .A(in[135]), .B(n3594), .Z(n4647) );
  XOR U924 ( .A(in[39]), .B(in[679]), .Z(n557) );
  XNOR U925 ( .A(in[359]), .B(in[1319]), .Z(n556) );
  XNOR U926 ( .A(n557), .B(n556), .Z(n558) );
  XOR U927 ( .A(in[999]), .B(n558), .Z(n1308) );
  XOR U928 ( .A(in[168]), .B(in[1448]), .Z(n560) );
  XNOR U929 ( .A(in[1128]), .B(in[808]), .Z(n559) );
  XNOR U930 ( .A(n560), .B(n559), .Z(n561) );
  XOR U931 ( .A(in[488]), .B(n561), .Z(n824) );
  XNOR U932 ( .A(n1308), .B(n824), .Z(n3967) );
  XNOR U933 ( .A(in[1384]), .B(n3967), .Z(n4644) );
  NAND U934 ( .A(n4647), .B(n4644), .Z(n562) );
  XNOR U935 ( .A(n1412), .B(n562), .Z(out[1028]) );
  XNOR U936 ( .A(n564), .B(n563), .Z(n3645) );
  XNOR U937 ( .A(in[536]), .B(n3645), .Z(n1416) );
  XOR U938 ( .A(in[1351]), .B(in[711]), .Z(n566) );
  XNOR U939 ( .A(in[1031]), .B(in[391]), .Z(n565) );
  XNOR U940 ( .A(n566), .B(n565), .Z(n567) );
  XOR U941 ( .A(in[71]), .B(n567), .Z(n1505) );
  XOR U942 ( .A(in[1480]), .B(in[520]), .Z(n569) );
  XNOR U943 ( .A(in[840]), .B(in[200]), .Z(n568) );
  XNOR U944 ( .A(n569), .B(n568), .Z(n570) );
  XNOR U945 ( .A(in[1160]), .B(n570), .Z(n1213) );
  XNOR U946 ( .A(n1505), .B(n1213), .Z(n3598) );
  XNOR U947 ( .A(in[136]), .B(n3598), .Z(n4651) );
  XOR U948 ( .A(in[169]), .B(in[1449]), .Z(n572) );
  XNOR U949 ( .A(in[1129]), .B(in[809]), .Z(n571) );
  XNOR U950 ( .A(n572), .B(n571), .Z(n573) );
  XOR U951 ( .A(in[489]), .B(n573), .Z(n837) );
  XOR U952 ( .A(in[680]), .B(in[1320]), .Z(n575) );
  XNOR U953 ( .A(in[40]), .B(in[360]), .Z(n574) );
  XNOR U954 ( .A(n575), .B(n574), .Z(n576) );
  XOR U955 ( .A(in[1000]), .B(n576), .Z(n1312) );
  XNOR U956 ( .A(n837), .B(n1312), .Z(n3974) );
  XNOR U957 ( .A(in[1385]), .B(n3974), .Z(n4648) );
  NAND U958 ( .A(n4651), .B(n4648), .Z(n577) );
  XNOR U959 ( .A(n1416), .B(n577), .Z(out[1029]) );
  XOR U960 ( .A(in[1341]), .B(in[61]), .Z(n579) );
  XNOR U961 ( .A(in[701]), .B(in[381]), .Z(n578) );
  XNOR U962 ( .A(n579), .B(n578), .Z(n580) );
  XOR U963 ( .A(in[1021]), .B(n580), .Z(n894) );
  XNOR U964 ( .A(n581), .B(n894), .Z(n3600) );
  XNOR U965 ( .A(in[637]), .B(n3600), .Z(n2555) );
  XOR U966 ( .A(n583), .B(n582), .Z(n3697) );
  XNOR U967 ( .A(in[228]), .B(n3697), .Z(n2859) );
  XOR U968 ( .A(in[1512]), .B(in[552]), .Z(n585) );
  XNOR U969 ( .A(in[872]), .B(in[232]), .Z(n584) );
  XNOR U970 ( .A(n585), .B(n584), .Z(n586) );
  XOR U971 ( .A(in[1192]), .B(n586), .Z(n1317) );
  XNOR U972 ( .A(n587), .B(n1317), .Z(n3738) );
  XNOR U973 ( .A(in[1448]), .B(n3738), .Z(n2856) );
  NAND U974 ( .A(n2859), .B(n2856), .Z(n588) );
  XNOR U975 ( .A(n2555), .B(n588), .Z(out[102]) );
  XOR U976 ( .A(n590), .B(n589), .Z(n3649) );
  XNOR U977 ( .A(in[537]), .B(n3649), .Z(n1420) );
  XOR U978 ( .A(in[1352]), .B(in[712]), .Z(n592) );
  XNOR U979 ( .A(in[1032]), .B(in[392]), .Z(n591) );
  XNOR U980 ( .A(n592), .B(n591), .Z(n593) );
  XOR U981 ( .A(in[72]), .B(n593), .Z(n1510) );
  XOR U982 ( .A(in[1481]), .B(in[521]), .Z(n595) );
  XNOR U983 ( .A(in[841]), .B(in[201]), .Z(n594) );
  XNOR U984 ( .A(n595), .B(n594), .Z(n596) );
  XNOR U985 ( .A(in[1161]), .B(n596), .Z(n1216) );
  XNOR U986 ( .A(n1510), .B(n1216), .Z(n3602) );
  XNOR U987 ( .A(in[137]), .B(n3602), .Z(n4655) );
  XOR U988 ( .A(in[170]), .B(in[1450]), .Z(n598) );
  XNOR U989 ( .A(in[1130]), .B(in[810]), .Z(n597) );
  XNOR U990 ( .A(n598), .B(n597), .Z(n599) );
  XOR U991 ( .A(in[490]), .B(n599), .Z(n853) );
  XOR U992 ( .A(in[681]), .B(in[1321]), .Z(n601) );
  XNOR U993 ( .A(in[41]), .B(in[361]), .Z(n600) );
  XNOR U994 ( .A(n601), .B(n600), .Z(n602) );
  XOR U995 ( .A(in[1001]), .B(n602), .Z(n1316) );
  XNOR U996 ( .A(n853), .B(n1316), .Z(n3977) );
  XNOR U997 ( .A(in[1386]), .B(n3977), .Z(n4652) );
  NAND U998 ( .A(n4655), .B(n4652), .Z(n603) );
  XNOR U999 ( .A(n1420), .B(n603), .Z(out[1030]) );
  XNOR U1000 ( .A(n605), .B(n604), .Z(n3653) );
  XNOR U1001 ( .A(in[538]), .B(n3653), .Z(n1424) );
  XOR U1002 ( .A(in[1353]), .B(in[393]), .Z(n607) );
  XNOR U1003 ( .A(in[713]), .B(in[73]), .Z(n606) );
  XNOR U1004 ( .A(n607), .B(n606), .Z(n608) );
  XOR U1005 ( .A(in[1033]), .B(n608), .Z(n1514) );
  XOR U1006 ( .A(in[1482]), .B(in[522]), .Z(n610) );
  XNOR U1007 ( .A(in[842]), .B(in[202]), .Z(n609) );
  XNOR U1008 ( .A(n610), .B(n609), .Z(n611) );
  XNOR U1009 ( .A(in[1162]), .B(n611), .Z(n1219) );
  XNOR U1010 ( .A(n1514), .B(n1219), .Z(n3606) );
  XNOR U1011 ( .A(in[138]), .B(n3606), .Z(n4659) );
  XOR U1012 ( .A(in[811]), .B(in[491]), .Z(n613) );
  XNOR U1013 ( .A(in[1451]), .B(in[1131]), .Z(n612) );
  XNOR U1014 ( .A(n613), .B(n612), .Z(n614) );
  XOR U1015 ( .A(in[171]), .B(n614), .Z(n866) );
  XOR U1016 ( .A(in[682]), .B(in[1322]), .Z(n616) );
  XNOR U1017 ( .A(in[42]), .B(in[362]), .Z(n615) );
  XNOR U1018 ( .A(n616), .B(n615), .Z(n617) );
  XOR U1019 ( .A(in[1002]), .B(n617), .Z(n1321) );
  XNOR U1020 ( .A(n866), .B(n1321), .Z(n3980) );
  XNOR U1021 ( .A(in[1387]), .B(n3980), .Z(n4656) );
  NAND U1022 ( .A(n4659), .B(n4656), .Z(n618) );
  XNOR U1023 ( .A(n1424), .B(n618), .Z(out[1031]) );
  XOR U1024 ( .A(n620), .B(n619), .Z(n3657) );
  XNOR U1025 ( .A(in[539]), .B(n3657), .Z(n1429) );
  XOR U1026 ( .A(in[1483]), .B(in[523]), .Z(n622) );
  XNOR U1027 ( .A(in[843]), .B(in[203]), .Z(n621) );
  XNOR U1028 ( .A(n622), .B(n621), .Z(n623) );
  XOR U1029 ( .A(in[1163]), .B(n623), .Z(n1222) );
  XOR U1030 ( .A(in[1354]), .B(in[714]), .Z(n625) );
  XNOR U1031 ( .A(in[74]), .B(in[394]), .Z(n624) );
  XNOR U1032 ( .A(n625), .B(n624), .Z(n626) );
  XNOR U1033 ( .A(in[1034]), .B(n626), .Z(n1518) );
  XNOR U1034 ( .A(n1222), .B(n1518), .Z(n3610) );
  XNOR U1035 ( .A(n3610), .B(in[139]), .Z(n4663) );
  XOR U1036 ( .A(in[683]), .B(in[1323]), .Z(n628) );
  XNOR U1037 ( .A(in[43]), .B(in[363]), .Z(n627) );
  XNOR U1038 ( .A(n628), .B(n627), .Z(n629) );
  XOR U1039 ( .A(in[1003]), .B(n629), .Z(n1325) );
  XOR U1040 ( .A(in[812]), .B(in[492]), .Z(n631) );
  XNOR U1041 ( .A(in[1452]), .B(in[1132]), .Z(n630) );
  XNOR U1042 ( .A(n631), .B(n630), .Z(n632) );
  XOR U1043 ( .A(in[172]), .B(n632), .Z(n886) );
  XNOR U1044 ( .A(n1325), .B(n886), .Z(n3983) );
  XNOR U1045 ( .A(in[1388]), .B(n3983), .Z(n4660) );
  NAND U1046 ( .A(n4663), .B(n4660), .Z(n633) );
  XNOR U1047 ( .A(n1429), .B(n633), .Z(out[1032]) );
  XNOR U1048 ( .A(n635), .B(n634), .Z(n3661) );
  XNOR U1049 ( .A(in[540]), .B(n3661), .Z(n1433) );
  XOR U1050 ( .A(in[1355]), .B(in[715]), .Z(n637) );
  XNOR U1051 ( .A(in[1035]), .B(in[395]), .Z(n636) );
  XNOR U1052 ( .A(n637), .B(n636), .Z(n638) );
  XOR U1053 ( .A(in[75]), .B(n638), .Z(n1522) );
  XOR U1054 ( .A(in[1484]), .B(in[524]), .Z(n640) );
  XNOR U1055 ( .A(in[844]), .B(in[204]), .Z(n639) );
  XNOR U1056 ( .A(n640), .B(n639), .Z(n641) );
  XNOR U1057 ( .A(in[1164]), .B(n641), .Z(n1225) );
  XNOR U1058 ( .A(n1522), .B(n1225), .Z(n3614) );
  XNOR U1059 ( .A(in[140]), .B(n3614), .Z(n4667) );
  XOR U1060 ( .A(in[813]), .B(in[493]), .Z(n643) );
  XNOR U1061 ( .A(in[1453]), .B(in[1133]), .Z(n642) );
  XNOR U1062 ( .A(n643), .B(n642), .Z(n644) );
  XOR U1063 ( .A(in[173]), .B(n644), .Z(n899) );
  XOR U1064 ( .A(in[1324]), .B(in[44]), .Z(n646) );
  XNOR U1065 ( .A(in[684]), .B(in[364]), .Z(n645) );
  XNOR U1066 ( .A(n646), .B(n645), .Z(n647) );
  XOR U1067 ( .A(in[1004]), .B(n647), .Z(n1328) );
  XNOR U1068 ( .A(n899), .B(n1328), .Z(n3986) );
  XNOR U1069 ( .A(in[1389]), .B(n3986), .Z(n4664) );
  NAND U1070 ( .A(n4667), .B(n4664), .Z(n648) );
  XNOR U1071 ( .A(n1433), .B(n648), .Z(out[1033]) );
  XNOR U1072 ( .A(n650), .B(n649), .Z(n3669) );
  XNOR U1073 ( .A(in[541]), .B(n3669), .Z(n1437) );
  XOR U1074 ( .A(in[76]), .B(in[1036]), .Z(n652) );
  XNOR U1075 ( .A(in[716]), .B(in[396]), .Z(n651) );
  XNOR U1076 ( .A(n652), .B(n651), .Z(n653) );
  XOR U1077 ( .A(in[1356]), .B(n653), .Z(n1526) );
  XOR U1078 ( .A(in[1485]), .B(in[525]), .Z(n655) );
  XNOR U1079 ( .A(in[845]), .B(in[205]), .Z(n654) );
  XNOR U1080 ( .A(n655), .B(n654), .Z(n656) );
  XNOR U1081 ( .A(in[1165]), .B(n656), .Z(n1228) );
  XNOR U1082 ( .A(n1526), .B(n1228), .Z(n3618) );
  XNOR U1083 ( .A(in[141]), .B(n3618), .Z(n4675) );
  XOR U1084 ( .A(in[814]), .B(in[494]), .Z(n658) );
  XNOR U1085 ( .A(in[1454]), .B(in[1134]), .Z(n657) );
  XNOR U1086 ( .A(n658), .B(n657), .Z(n659) );
  XOR U1087 ( .A(in[174]), .B(n659), .Z(n912) );
  XOR U1088 ( .A(in[1325]), .B(in[45]), .Z(n661) );
  XNOR U1089 ( .A(in[685]), .B(in[365]), .Z(n660) );
  XNOR U1090 ( .A(n661), .B(n660), .Z(n662) );
  XOR U1091 ( .A(in[1005]), .B(n662), .Z(n1332) );
  XNOR U1092 ( .A(n912), .B(n1332), .Z(n3989) );
  XNOR U1093 ( .A(in[1390]), .B(n3989), .Z(n4672) );
  NAND U1094 ( .A(n4675), .B(n4672), .Z(n663) );
  XNOR U1095 ( .A(n1437), .B(n663), .Z(out[1034]) );
  XNOR U1096 ( .A(n665), .B(n664), .Z(n3673) );
  XNOR U1097 ( .A(in[542]), .B(n3673), .Z(n1441) );
  XOR U1098 ( .A(in[77]), .B(in[1037]), .Z(n667) );
  XNOR U1099 ( .A(in[717]), .B(in[397]), .Z(n666) );
  XNOR U1100 ( .A(n667), .B(n666), .Z(n668) );
  XOR U1101 ( .A(in[1357]), .B(n668), .Z(n1530) );
  XOR U1102 ( .A(in[1486]), .B(in[526]), .Z(n670) );
  XNOR U1103 ( .A(in[846]), .B(in[206]), .Z(n669) );
  XNOR U1104 ( .A(n670), .B(n669), .Z(n671) );
  XNOR U1105 ( .A(in[1166]), .B(n671), .Z(n1231) );
  XNOR U1106 ( .A(n1530), .B(n1231), .Z(n3626) );
  XNOR U1107 ( .A(in[142]), .B(n3626), .Z(n4679) );
  XOR U1108 ( .A(in[815]), .B(in[495]), .Z(n673) );
  XNOR U1109 ( .A(in[1455]), .B(in[1135]), .Z(n672) );
  XNOR U1110 ( .A(n673), .B(n672), .Z(n674) );
  XOR U1111 ( .A(in[175]), .B(n674), .Z(n925) );
  XOR U1112 ( .A(in[1326]), .B(in[46]), .Z(n676) );
  XNOR U1113 ( .A(in[686]), .B(in[366]), .Z(n675) );
  XNOR U1114 ( .A(n676), .B(n675), .Z(n677) );
  XOR U1115 ( .A(in[1006]), .B(n677), .Z(n1336) );
  XNOR U1116 ( .A(n925), .B(n1336), .Z(n3992) );
  XNOR U1117 ( .A(in[1391]), .B(n3992), .Z(n4676) );
  NAND U1118 ( .A(n4679), .B(n4676), .Z(n678) );
  XNOR U1119 ( .A(n1441), .B(n678), .Z(out[1035]) );
  XNOR U1120 ( .A(n680), .B(n679), .Z(n3677) );
  XNOR U1121 ( .A(in[543]), .B(n3677), .Z(n1445) );
  XOR U1122 ( .A(in[78]), .B(in[1038]), .Z(n682) );
  XNOR U1123 ( .A(in[718]), .B(in[398]), .Z(n681) );
  XNOR U1124 ( .A(n682), .B(n681), .Z(n683) );
  XOR U1125 ( .A(in[1358]), .B(n683), .Z(n1534) );
  XOR U1126 ( .A(in[1487]), .B(in[527]), .Z(n685) );
  XNOR U1127 ( .A(in[847]), .B(in[207]), .Z(n684) );
  XNOR U1128 ( .A(n685), .B(n684), .Z(n686) );
  XNOR U1129 ( .A(in[1167]), .B(n686), .Z(n1234) );
  XNOR U1130 ( .A(n1534), .B(n1234), .Z(n3630) );
  XNOR U1131 ( .A(in[143]), .B(n3630), .Z(n4683) );
  XOR U1132 ( .A(in[1327]), .B(in[47]), .Z(n688) );
  XNOR U1133 ( .A(in[687]), .B(in[367]), .Z(n687) );
  XNOR U1134 ( .A(n688), .B(n687), .Z(n689) );
  XOR U1135 ( .A(in[1007]), .B(n689), .Z(n1340) );
  XOR U1136 ( .A(in[816]), .B(in[496]), .Z(n691) );
  XNOR U1137 ( .A(in[1456]), .B(in[1136]), .Z(n690) );
  XNOR U1138 ( .A(n691), .B(n690), .Z(n692) );
  XOR U1139 ( .A(in[176]), .B(n692), .Z(n940) );
  XNOR U1140 ( .A(n1340), .B(n940), .Z(n3995) );
  XNOR U1141 ( .A(in[1392]), .B(n3995), .Z(n4680) );
  NAND U1142 ( .A(n4683), .B(n4680), .Z(n693) );
  XNOR U1143 ( .A(n1445), .B(n693), .Z(out[1036]) );
  XNOR U1144 ( .A(n695), .B(n694), .Z(n3681) );
  XNOR U1145 ( .A(in[544]), .B(n3681), .Z(n1449) );
  XOR U1146 ( .A(in[79]), .B(in[1039]), .Z(n697) );
  XNOR U1147 ( .A(in[719]), .B(in[399]), .Z(n696) );
  XNOR U1148 ( .A(n697), .B(n696), .Z(n698) );
  XOR U1149 ( .A(in[1359]), .B(n698), .Z(n1538) );
  XOR U1150 ( .A(in[1488]), .B(in[528]), .Z(n700) );
  XNOR U1151 ( .A(in[848]), .B(in[208]), .Z(n699) );
  XNOR U1152 ( .A(n700), .B(n699), .Z(n701) );
  XNOR U1153 ( .A(in[1168]), .B(n701), .Z(n1237) );
  XNOR U1154 ( .A(n1538), .B(n1237), .Z(n3634) );
  XNOR U1155 ( .A(in[144]), .B(n3634), .Z(n4687) );
  XOR U1156 ( .A(in[817]), .B(in[497]), .Z(n703) );
  XNOR U1157 ( .A(in[1457]), .B(in[1137]), .Z(n702) );
  XNOR U1158 ( .A(n703), .B(n702), .Z(n704) );
  XOR U1159 ( .A(in[177]), .B(n704), .Z(n955) );
  XOR U1160 ( .A(in[1328]), .B(in[48]), .Z(n706) );
  XNOR U1161 ( .A(in[688]), .B(in[368]), .Z(n705) );
  XNOR U1162 ( .A(n706), .B(n705), .Z(n707) );
  XOR U1163 ( .A(in[1008]), .B(n707), .Z(n1344) );
  XNOR U1164 ( .A(n955), .B(n1344), .Z(n3998) );
  XNOR U1165 ( .A(in[1393]), .B(n3998), .Z(n4684) );
  NAND U1166 ( .A(n4687), .B(n4684), .Z(n708) );
  XNOR U1167 ( .A(n1449), .B(n708), .Z(out[1037]) );
  XNOR U1168 ( .A(n710), .B(n709), .Z(n3685) );
  XNOR U1169 ( .A(in[545]), .B(n3685), .Z(n1453) );
  XOR U1170 ( .A(in[80]), .B(in[1040]), .Z(n712) );
  XNOR U1171 ( .A(in[720]), .B(in[400]), .Z(n711) );
  XNOR U1172 ( .A(n712), .B(n711), .Z(n713) );
  XOR U1173 ( .A(in[1360]), .B(n713), .Z(n1542) );
  XOR U1174 ( .A(in[1489]), .B(in[529]), .Z(n715) );
  XNOR U1175 ( .A(in[849]), .B(in[209]), .Z(n714) );
  XNOR U1176 ( .A(n715), .B(n714), .Z(n716) );
  XNOR U1177 ( .A(in[1169]), .B(n716), .Z(n1240) );
  XNOR U1178 ( .A(n1542), .B(n1240), .Z(n3638) );
  XNOR U1179 ( .A(in[145]), .B(n3638), .Z(n4691) );
  XOR U1180 ( .A(in[1329]), .B(in[49]), .Z(n718) );
  XNOR U1181 ( .A(in[689]), .B(in[369]), .Z(n717) );
  XNOR U1182 ( .A(n718), .B(n717), .Z(n719) );
  XOR U1183 ( .A(in[1009]), .B(n719), .Z(n1349) );
  XOR U1184 ( .A(in[818]), .B(in[498]), .Z(n721) );
  XNOR U1185 ( .A(in[1458]), .B(in[1138]), .Z(n720) );
  XNOR U1186 ( .A(n721), .B(n720), .Z(n722) );
  XOR U1187 ( .A(in[178]), .B(n722), .Z(n970) );
  XNOR U1188 ( .A(n1349), .B(n970), .Z(n4001) );
  XNOR U1189 ( .A(in[1394]), .B(n4001), .Z(n4688) );
  NAND U1190 ( .A(n4691), .B(n4688), .Z(n723) );
  XNOR U1191 ( .A(n1453), .B(n723), .Z(out[1038]) );
  XOR U1192 ( .A(n3689), .B(in[546]), .Z(n1457) );
  XOR U1193 ( .A(in[81]), .B(in[1041]), .Z(n725) );
  XNOR U1194 ( .A(in[721]), .B(in[401]), .Z(n724) );
  XNOR U1195 ( .A(n725), .B(n724), .Z(n726) );
  XOR U1196 ( .A(in[1361]), .B(n726), .Z(n1546) );
  XOR U1197 ( .A(in[1490]), .B(in[530]), .Z(n728) );
  XNOR U1198 ( .A(in[850]), .B(in[210]), .Z(n727) );
  XNOR U1199 ( .A(n728), .B(n727), .Z(n729) );
  XNOR U1200 ( .A(in[1170]), .B(n729), .Z(n1244) );
  XNOR U1201 ( .A(n1546), .B(n1244), .Z(n3642) );
  XNOR U1202 ( .A(in[146]), .B(n3642), .Z(n4695) );
  XOR U1203 ( .A(in[819]), .B(in[499]), .Z(n731) );
  XNOR U1204 ( .A(in[1459]), .B(in[1139]), .Z(n730) );
  XNOR U1205 ( .A(n731), .B(n730), .Z(n732) );
  XOR U1206 ( .A(in[179]), .B(n732), .Z(n985) );
  XOR U1207 ( .A(in[1330]), .B(in[50]), .Z(n734) );
  XNOR U1208 ( .A(in[690]), .B(in[370]), .Z(n733) );
  XNOR U1209 ( .A(n734), .B(n733), .Z(n735) );
  XOR U1210 ( .A(in[1010]), .B(n735), .Z(n1353) );
  XNOR U1211 ( .A(n985), .B(n1353), .Z(n4008) );
  XNOR U1212 ( .A(in[1395]), .B(n4008), .Z(n4692) );
  NAND U1213 ( .A(n4695), .B(n4692), .Z(n736) );
  XNOR U1214 ( .A(n1457), .B(n736), .Z(out[1039]) );
  XOR U1215 ( .A(in[1342]), .B(in[62]), .Z(n738) );
  XNOR U1216 ( .A(in[702]), .B(in[382]), .Z(n737) );
  XNOR U1217 ( .A(n738), .B(n737), .Z(n739) );
  XOR U1218 ( .A(in[1022]), .B(n739), .Z(n907) );
  XNOR U1219 ( .A(n740), .B(n907), .Z(n3604) );
  XNOR U1220 ( .A(in[638]), .B(n3604), .Z(n2557) );
  XOR U1221 ( .A(n742), .B(n741), .Z(n3701) );
  XNOR U1222 ( .A(in[229]), .B(n3701), .Z(n2873) );
  XOR U1223 ( .A(in[1513]), .B(in[553]), .Z(n744) );
  XNOR U1224 ( .A(in[873]), .B(in[233]), .Z(n743) );
  XNOR U1225 ( .A(n744), .B(n743), .Z(n745) );
  XOR U1226 ( .A(in[1193]), .B(n745), .Z(n1320) );
  XNOR U1227 ( .A(n746), .B(n1320), .Z(n3742) );
  XNOR U1228 ( .A(in[1449]), .B(n3742), .Z(n2870) );
  NAND U1229 ( .A(n2873), .B(n2870), .Z(n747) );
  XNOR U1230 ( .A(n2557), .B(n747), .Z(out[103]) );
  XOR U1231 ( .A(n3693), .B(in[547]), .Z(n1461) );
  XOR U1232 ( .A(in[1042]), .B(in[402]), .Z(n749) );
  XNOR U1233 ( .A(in[722]), .B(in[82]), .Z(n748) );
  XNOR U1234 ( .A(n749), .B(n748), .Z(n750) );
  XOR U1235 ( .A(in[1362]), .B(n750), .Z(n1551) );
  XOR U1236 ( .A(in[851]), .B(in[1171]), .Z(n752) );
  XNOR U1237 ( .A(in[1491]), .B(in[211]), .Z(n751) );
  XNOR U1238 ( .A(n752), .B(n751), .Z(n753) );
  XNOR U1239 ( .A(in[531]), .B(n753), .Z(n1247) );
  XNOR U1240 ( .A(n1551), .B(n1247), .Z(n3646) );
  XNOR U1241 ( .A(in[147]), .B(n3646), .Z(n4699) );
  XOR U1242 ( .A(in[820]), .B(in[500]), .Z(n755) );
  XNOR U1243 ( .A(in[1460]), .B(in[1140]), .Z(n754) );
  XNOR U1244 ( .A(n755), .B(n754), .Z(n756) );
  XOR U1245 ( .A(in[180]), .B(n756), .Z(n1000) );
  XOR U1246 ( .A(in[1331]), .B(in[51]), .Z(n758) );
  XNOR U1247 ( .A(in[691]), .B(in[371]), .Z(n757) );
  XNOR U1248 ( .A(n758), .B(n757), .Z(n759) );
  XOR U1249 ( .A(in[1011]), .B(n759), .Z(n1357) );
  XNOR U1250 ( .A(n1000), .B(n1357), .Z(n4011) );
  XNOR U1251 ( .A(in[1396]), .B(n4011), .Z(n4696) );
  NAND U1252 ( .A(n4699), .B(n4696), .Z(n760) );
  XNOR U1253 ( .A(n1461), .B(n760), .Z(out[1040]) );
  XOR U1254 ( .A(n3697), .B(in[548]), .Z(n1465) );
  XOR U1255 ( .A(in[83]), .B(in[1043]), .Z(n762) );
  XNOR U1256 ( .A(in[723]), .B(in[403]), .Z(n761) );
  XNOR U1257 ( .A(n762), .B(n761), .Z(n763) );
  XOR U1258 ( .A(in[1363]), .B(n763), .Z(n1555) );
  XOR U1259 ( .A(in[852]), .B(in[1172]), .Z(n765) );
  XNOR U1260 ( .A(in[1492]), .B(in[212]), .Z(n764) );
  XNOR U1261 ( .A(n765), .B(n764), .Z(n766) );
  XNOR U1262 ( .A(in[532]), .B(n766), .Z(n1250) );
  XNOR U1263 ( .A(n1555), .B(n1250), .Z(n3650) );
  XNOR U1264 ( .A(in[148]), .B(n3650), .Z(n4703) );
  XOR U1265 ( .A(in[1332]), .B(in[52]), .Z(n768) );
  XNOR U1266 ( .A(in[692]), .B(in[372]), .Z(n767) );
  XNOR U1267 ( .A(n768), .B(n767), .Z(n769) );
  XOR U1268 ( .A(in[1012]), .B(n769), .Z(n1361) );
  XOR U1269 ( .A(in[821]), .B(in[501]), .Z(n771) );
  XNOR U1270 ( .A(in[1461]), .B(in[1141]), .Z(n770) );
  XNOR U1271 ( .A(n771), .B(n770), .Z(n772) );
  XOR U1272 ( .A(in[181]), .B(n772), .Z(n1015) );
  XNOR U1273 ( .A(n1361), .B(n1015), .Z(n4014) );
  XNOR U1274 ( .A(in[1397]), .B(n4014), .Z(n4700) );
  NAND U1275 ( .A(n4703), .B(n4700), .Z(n773) );
  XNOR U1276 ( .A(n1465), .B(n773), .Z(out[1041]) );
  XOR U1277 ( .A(n3701), .B(in[549]), .Z(n1470) );
  XOR U1278 ( .A(in[853]), .B(in[1173]), .Z(n775) );
  XNOR U1279 ( .A(in[1493]), .B(in[213]), .Z(n774) );
  XNOR U1280 ( .A(n775), .B(n774), .Z(n776) );
  XNOR U1281 ( .A(in[533]), .B(n776), .Z(n1253) );
  XNOR U1282 ( .A(n777), .B(n1253), .Z(n3654) );
  XNOR U1283 ( .A(in[149]), .B(n3654), .Z(n4707) );
  XOR U1284 ( .A(in[822]), .B(in[502]), .Z(n779) );
  XNOR U1285 ( .A(in[1462]), .B(in[1142]), .Z(n778) );
  XNOR U1286 ( .A(n779), .B(n778), .Z(n780) );
  XOR U1287 ( .A(in[182]), .B(n780), .Z(n1029) );
  XOR U1288 ( .A(in[1333]), .B(in[53]), .Z(n782) );
  XNOR U1289 ( .A(in[693]), .B(in[373]), .Z(n781) );
  XNOR U1290 ( .A(n782), .B(n781), .Z(n783) );
  XOR U1291 ( .A(in[1013]), .B(n783), .Z(n1365) );
  XNOR U1292 ( .A(n1029), .B(n1365), .Z(n4017) );
  XNOR U1293 ( .A(in[1398]), .B(n4017), .Z(n4704) );
  NAND U1294 ( .A(n4707), .B(n4704), .Z(n784) );
  XNOR U1295 ( .A(n1470), .B(n784), .Z(out[1042]) );
  XNOR U1296 ( .A(n786), .B(n785), .Z(n3705) );
  XNOR U1297 ( .A(in[550]), .B(n3705), .Z(n1474) );
  XOR U1298 ( .A(in[854]), .B(in[1174]), .Z(n788) );
  XNOR U1299 ( .A(in[1494]), .B(in[214]), .Z(n787) );
  XNOR U1300 ( .A(n788), .B(n787), .Z(n789) );
  XNOR U1301 ( .A(in[534]), .B(n789), .Z(n1256) );
  XNOR U1302 ( .A(n790), .B(n1256), .Z(n3658) );
  XNOR U1303 ( .A(in[150]), .B(n3658), .Z(n4711) );
  XOR U1304 ( .A(in[823]), .B(in[503]), .Z(n792) );
  XNOR U1305 ( .A(in[1463]), .B(in[1143]), .Z(n791) );
  XNOR U1306 ( .A(n792), .B(n791), .Z(n793) );
  XOR U1307 ( .A(in[183]), .B(n793), .Z(n1040) );
  XOR U1308 ( .A(in[1334]), .B(in[54]), .Z(n795) );
  XNOR U1309 ( .A(in[694]), .B(in[374]), .Z(n794) );
  XNOR U1310 ( .A(n795), .B(n794), .Z(n796) );
  XOR U1311 ( .A(in[1014]), .B(n796), .Z(n1369) );
  XNOR U1312 ( .A(n1040), .B(n1369), .Z(n4020) );
  XNOR U1313 ( .A(in[1399]), .B(n4020), .Z(n4708) );
  NAND U1314 ( .A(n4711), .B(n4708), .Z(n797) );
  XNOR U1315 ( .A(n1474), .B(n797), .Z(out[1043]) );
  XNOR U1316 ( .A(n799), .B(n798), .Z(n3713) );
  XNOR U1317 ( .A(in[551]), .B(n3713), .Z(n1478) );
  XOR U1318 ( .A(in[855]), .B(in[1175]), .Z(n801) );
  XNOR U1319 ( .A(in[1495]), .B(in[215]), .Z(n800) );
  XNOR U1320 ( .A(n801), .B(n800), .Z(n802) );
  XNOR U1321 ( .A(in[535]), .B(n802), .Z(n1259) );
  XNOR U1322 ( .A(n803), .B(n1259), .Z(n3662) );
  XNOR U1323 ( .A(in[151]), .B(n3662), .Z(n4719) );
  XOR U1324 ( .A(in[824]), .B(in[504]), .Z(n805) );
  XNOR U1325 ( .A(in[1464]), .B(in[1144]), .Z(n804) );
  XNOR U1326 ( .A(n805), .B(n804), .Z(n806) );
  XOR U1327 ( .A(in[184]), .B(n806), .Z(n1045) );
  XOR U1328 ( .A(in[1335]), .B(in[55]), .Z(n808) );
  XNOR U1329 ( .A(in[695]), .B(in[375]), .Z(n807) );
  XNOR U1330 ( .A(n808), .B(n807), .Z(n809) );
  XOR U1331 ( .A(in[1015]), .B(n809), .Z(n1373) );
  XNOR U1332 ( .A(n1045), .B(n1373), .Z(n4023) );
  XNOR U1333 ( .A(in[1400]), .B(n4023), .Z(n4716) );
  NAND U1334 ( .A(n4719), .B(n4716), .Z(n810) );
  XNOR U1335 ( .A(n1478), .B(n810), .Z(out[1044]) );
  XNOR U1336 ( .A(n812), .B(n811), .Z(n3717) );
  XNOR U1337 ( .A(in[552]), .B(n3717), .Z(n1482) );
  XOR U1338 ( .A(in[856]), .B(in[1176]), .Z(n814) );
  XNOR U1339 ( .A(in[1496]), .B(in[216]), .Z(n813) );
  XNOR U1340 ( .A(n814), .B(n813), .Z(n815) );
  XNOR U1341 ( .A(in[536]), .B(n815), .Z(n1262) );
  XNOR U1342 ( .A(n816), .B(n1262), .Z(n3670) );
  XNOR U1343 ( .A(in[152]), .B(n3670), .Z(n4723) );
  XOR U1344 ( .A(in[1336]), .B(in[56]), .Z(n818) );
  XNOR U1345 ( .A(in[696]), .B(in[376]), .Z(n817) );
  XNOR U1346 ( .A(n818), .B(n817), .Z(n819) );
  XOR U1347 ( .A(in[1016]), .B(n819), .Z(n1377) );
  XOR U1348 ( .A(in[825]), .B(in[505]), .Z(n821) );
  XNOR U1349 ( .A(in[1465]), .B(in[1145]), .Z(n820) );
  XNOR U1350 ( .A(n821), .B(n820), .Z(n822) );
  XOR U1351 ( .A(in[185]), .B(n822), .Z(n1056) );
  XNOR U1352 ( .A(n1377), .B(n1056), .Z(n4026) );
  XNOR U1353 ( .A(in[1401]), .B(n4026), .Z(n4720) );
  NAND U1354 ( .A(n4723), .B(n4720), .Z(n823) );
  XNOR U1355 ( .A(n1482), .B(n823), .Z(out[1045]) );
  XNOR U1356 ( .A(n825), .B(n824), .Z(n3721) );
  XNOR U1357 ( .A(in[553]), .B(n3721), .Z(n1486) );
  XOR U1358 ( .A(in[857]), .B(in[1177]), .Z(n827) );
  XNOR U1359 ( .A(in[1497]), .B(in[217]), .Z(n826) );
  XNOR U1360 ( .A(n827), .B(n826), .Z(n828) );
  XNOR U1361 ( .A(in[537]), .B(n828), .Z(n1265) );
  XNOR U1362 ( .A(n829), .B(n1265), .Z(n3674) );
  XNOR U1363 ( .A(in[153]), .B(n3674), .Z(n4727) );
  XOR U1364 ( .A(in[1337]), .B(in[57]), .Z(n831) );
  XNOR U1365 ( .A(in[697]), .B(in[377]), .Z(n830) );
  XNOR U1366 ( .A(n831), .B(n830), .Z(n832) );
  XOR U1367 ( .A(in[1017]), .B(n832), .Z(n1381) );
  XOR U1368 ( .A(in[826]), .B(in[506]), .Z(n834) );
  XNOR U1369 ( .A(in[1466]), .B(in[1146]), .Z(n833) );
  XNOR U1370 ( .A(n834), .B(n833), .Z(n835) );
  XOR U1371 ( .A(in[186]), .B(n835), .Z(n1067) );
  XNOR U1372 ( .A(n1381), .B(n1067), .Z(n4029) );
  XNOR U1373 ( .A(in[1402]), .B(n4029), .Z(n4724) );
  NAND U1374 ( .A(n4727), .B(n4724), .Z(n836) );
  XNOR U1375 ( .A(n1486), .B(n836), .Z(out[1046]) );
  XNOR U1376 ( .A(n838), .B(n837), .Z(n3725) );
  XNOR U1377 ( .A(in[554]), .B(n3725), .Z(n1490) );
  XOR U1378 ( .A(in[858]), .B(in[1178]), .Z(n840) );
  XNOR U1379 ( .A(in[1498]), .B(in[218]), .Z(n839) );
  XNOR U1380 ( .A(n840), .B(n839), .Z(n841) );
  XNOR U1381 ( .A(in[538]), .B(n841), .Z(n1268) );
  XNOR U1382 ( .A(n842), .B(n1268), .Z(n3678) );
  XNOR U1383 ( .A(in[154]), .B(n3678), .Z(n4731) );
  XOR U1384 ( .A(in[1338]), .B(in[58]), .Z(n844) );
  XNOR U1385 ( .A(in[698]), .B(in[378]), .Z(n843) );
  XNOR U1386 ( .A(n844), .B(n843), .Z(n845) );
  XOR U1387 ( .A(in[1018]), .B(n845), .Z(n1385) );
  XOR U1388 ( .A(in[827]), .B(in[507]), .Z(n847) );
  XNOR U1389 ( .A(in[1467]), .B(in[1147]), .Z(n846) );
  XNOR U1390 ( .A(n847), .B(n846), .Z(n848) );
  XOR U1391 ( .A(in[187]), .B(n848), .Z(n1072) );
  XNOR U1392 ( .A(n1385), .B(n1072), .Z(n4032) );
  XNOR U1393 ( .A(in[1403]), .B(n4032), .Z(n4728) );
  NAND U1394 ( .A(n4731), .B(n4728), .Z(n849) );
  XNOR U1395 ( .A(n1490), .B(n849), .Z(out[1047]) );
  XOR U1396 ( .A(in[1579]), .B(in[619]), .Z(n851) );
  XNOR U1397 ( .A(in[939]), .B(in[299]), .Z(n850) );
  XNOR U1398 ( .A(n851), .B(n850), .Z(n852) );
  XOR U1399 ( .A(in[1259]), .B(n852), .Z(n1394) );
  XNOR U1400 ( .A(n853), .B(n1394), .Z(n3729) );
  XNOR U1401 ( .A(in[555]), .B(n3729), .Z(n1494) );
  XOR U1402 ( .A(in[859]), .B(in[1179]), .Z(n855) );
  XNOR U1403 ( .A(in[1499]), .B(in[219]), .Z(n854) );
  XNOR U1404 ( .A(n855), .B(n854), .Z(n856) );
  XNOR U1405 ( .A(in[539]), .B(n856), .Z(n1271) );
  XNOR U1406 ( .A(n857), .B(n1271), .Z(n3682) );
  XNOR U1407 ( .A(in[155]), .B(n3682), .Z(n4735) );
  XOR U1408 ( .A(in[828]), .B(in[508]), .Z(n859) );
  XNOR U1409 ( .A(in[1468]), .B(in[1148]), .Z(n858) );
  XNOR U1410 ( .A(n859), .B(n858), .Z(n860) );
  XOR U1411 ( .A(in[188]), .B(n860), .Z(n1077) );
  XNOR U1412 ( .A(n861), .B(n1077), .Z(n4035) );
  XNOR U1413 ( .A(in[1404]), .B(n4035), .Z(n4732) );
  NAND U1414 ( .A(n4735), .B(n4732), .Z(n862) );
  XNOR U1415 ( .A(n1494), .B(n862), .Z(out[1048]) );
  XOR U1416 ( .A(in[1580]), .B(in[620]), .Z(n864) );
  XNOR U1417 ( .A(in[940]), .B(in[300]), .Z(n863) );
  XNOR U1418 ( .A(n864), .B(n863), .Z(n865) );
  XOR U1419 ( .A(in[1260]), .B(n865), .Z(n1398) );
  XNOR U1420 ( .A(n866), .B(n1398), .Z(n3733) );
  XNOR U1421 ( .A(in[556]), .B(n3733), .Z(n1498) );
  XOR U1422 ( .A(in[860]), .B(in[1180]), .Z(n868) );
  XNOR U1423 ( .A(in[1500]), .B(in[220]), .Z(n867) );
  XNOR U1424 ( .A(n868), .B(n867), .Z(n869) );
  XNOR U1425 ( .A(in[540]), .B(n869), .Z(n1275) );
  XNOR U1426 ( .A(n870), .B(n1275), .Z(n3686) );
  XNOR U1427 ( .A(in[156]), .B(n3686), .Z(n4739) );
  XNOR U1428 ( .A(n872), .B(n871), .Z(n4042) );
  XNOR U1429 ( .A(in[1405]), .B(n4042), .Z(n4736) );
  NAND U1430 ( .A(n4739), .B(n4736), .Z(n873) );
  XNOR U1431 ( .A(n1498), .B(n873), .Z(out[1049]) );
  XOR U1432 ( .A(in[1343]), .B(in[63]), .Z(n875) );
  XNOR U1433 ( .A(in[703]), .B(in[383]), .Z(n874) );
  XNOR U1434 ( .A(n875), .B(n874), .Z(n876) );
  XOR U1435 ( .A(in[1023]), .B(n876), .Z(n920) );
  XNOR U1436 ( .A(n877), .B(n920), .Z(n3608) );
  XNOR U1437 ( .A(in[639]), .B(n3608), .Z(n2559) );
  XOR U1438 ( .A(in[230]), .B(n3705), .Z(n2889) );
  XOR U1439 ( .A(in[874]), .B(in[1194]), .Z(n879) );
  XNOR U1440 ( .A(in[1514]), .B(in[234]), .Z(n878) );
  XNOR U1441 ( .A(n879), .B(n878), .Z(n880) );
  XOR U1442 ( .A(in[554]), .B(n880), .Z(n1324) );
  XNOR U1443 ( .A(n881), .B(n1324), .Z(n3746) );
  XNOR U1444 ( .A(in[1450]), .B(n3746), .Z(n2886) );
  NAND U1445 ( .A(n2889), .B(n2886), .Z(n882) );
  XNOR U1446 ( .A(n2559), .B(n882), .Z(out[104]) );
  XOR U1447 ( .A(in[1581]), .B(in[621]), .Z(n884) );
  XNOR U1448 ( .A(in[941]), .B(in[301]), .Z(n883) );
  XNOR U1449 ( .A(n884), .B(n883), .Z(n885) );
  XOR U1450 ( .A(in[1261]), .B(n885), .Z(n1402) );
  XNOR U1451 ( .A(n886), .B(n1402), .Z(n3737) );
  XNOR U1452 ( .A(in[557]), .B(n3737), .Z(n1502) );
  XOR U1453 ( .A(in[861]), .B(in[1181]), .Z(n888) );
  XNOR U1454 ( .A(in[1501]), .B(in[221]), .Z(n887) );
  XNOR U1455 ( .A(n888), .B(n887), .Z(n889) );
  XNOR U1456 ( .A(in[541]), .B(n889), .Z(n1278) );
  XNOR U1457 ( .A(n890), .B(n1278), .Z(n3690) );
  XNOR U1458 ( .A(in[157]), .B(n3690), .Z(n4743) );
  XOR U1459 ( .A(in[830]), .B(in[510]), .Z(n892) );
  XNOR U1460 ( .A(in[1470]), .B(in[1150]), .Z(n891) );
  XNOR U1461 ( .A(n892), .B(n891), .Z(n893) );
  XOR U1462 ( .A(in[190]), .B(n893), .Z(n1083) );
  XNOR U1463 ( .A(n894), .B(n1083), .Z(n4045) );
  XNOR U1464 ( .A(in[1406]), .B(n4045), .Z(n4740) );
  NAND U1465 ( .A(n4743), .B(n4740), .Z(n895) );
  XNOR U1466 ( .A(n1502), .B(n895), .Z(out[1050]) );
  XOR U1467 ( .A(in[1582]), .B(in[622]), .Z(n897) );
  XNOR U1468 ( .A(in[942]), .B(in[302]), .Z(n896) );
  XNOR U1469 ( .A(n897), .B(n896), .Z(n898) );
  XOR U1470 ( .A(in[1262]), .B(n898), .Z(n1406) );
  XNOR U1471 ( .A(n899), .B(n1406), .Z(n3741) );
  XNOR U1472 ( .A(in[558]), .B(n3741), .Z(n1506) );
  XOR U1473 ( .A(in[862]), .B(in[1182]), .Z(n901) );
  XNOR U1474 ( .A(in[1502]), .B(in[222]), .Z(n900) );
  XNOR U1475 ( .A(n901), .B(n900), .Z(n902) );
  XNOR U1476 ( .A(in[542]), .B(n902), .Z(n1281) );
  XNOR U1477 ( .A(n903), .B(n1281), .Z(n3694) );
  XNOR U1478 ( .A(in[158]), .B(n3694), .Z(n4747) );
  XOR U1479 ( .A(in[831]), .B(in[511]), .Z(n905) );
  XNOR U1480 ( .A(in[1471]), .B(in[1151]), .Z(n904) );
  XNOR U1481 ( .A(n905), .B(n904), .Z(n906) );
  XOR U1482 ( .A(in[191]), .B(n906), .Z(n1088) );
  XNOR U1483 ( .A(n907), .B(n1088), .Z(n4048) );
  XNOR U1484 ( .A(in[1407]), .B(n4048), .Z(n4744) );
  NAND U1485 ( .A(n4747), .B(n4744), .Z(n908) );
  XNOR U1486 ( .A(n1506), .B(n908), .Z(out[1051]) );
  XOR U1487 ( .A(in[1583]), .B(in[623]), .Z(n910) );
  XNOR U1488 ( .A(in[943]), .B(in[303]), .Z(n909) );
  XNOR U1489 ( .A(n910), .B(n909), .Z(n911) );
  XOR U1490 ( .A(in[1263]), .B(n911), .Z(n1410) );
  XNOR U1491 ( .A(n912), .B(n1410), .Z(n3745) );
  XNOR U1492 ( .A(in[559]), .B(n3745), .Z(n1511) );
  XOR U1493 ( .A(in[863]), .B(in[1183]), .Z(n914) );
  XNOR U1494 ( .A(in[1503]), .B(in[223]), .Z(n913) );
  XNOR U1495 ( .A(n914), .B(n913), .Z(n915) );
  XNOR U1496 ( .A(in[543]), .B(n915), .Z(n1284) );
  XNOR U1497 ( .A(n916), .B(n1284), .Z(n3698) );
  XNOR U1498 ( .A(in[159]), .B(n3698), .Z(n4751) );
  XOR U1499 ( .A(in[768]), .B(in[1088]), .Z(n918) );
  XNOR U1500 ( .A(in[448]), .B(in[1408]), .Z(n917) );
  XNOR U1501 ( .A(n918), .B(n917), .Z(n919) );
  XOR U1502 ( .A(in[128]), .B(n919), .Z(n1096) );
  XNOR U1503 ( .A(n920), .B(n1096), .Z(n4051) );
  XNOR U1504 ( .A(in[1344]), .B(n4051), .Z(n4748) );
  NAND U1505 ( .A(n4751), .B(n4748), .Z(n921) );
  XNOR U1506 ( .A(n1511), .B(n921), .Z(out[1052]) );
  XOR U1507 ( .A(in[1584]), .B(in[624]), .Z(n923) );
  XNOR U1508 ( .A(in[944]), .B(in[304]), .Z(n922) );
  XNOR U1509 ( .A(n923), .B(n922), .Z(n924) );
  XOR U1510 ( .A(in[1264]), .B(n924), .Z(n1414) );
  XNOR U1511 ( .A(n925), .B(n1414), .Z(n3749) );
  XNOR U1512 ( .A(in[560]), .B(n3749), .Z(n1515) );
  XOR U1513 ( .A(in[224]), .B(in[864]), .Z(n927) );
  XNOR U1514 ( .A(in[1184]), .B(in[1504]), .Z(n926) );
  XNOR U1515 ( .A(n927), .B(n926), .Z(n928) );
  XNOR U1516 ( .A(in[544]), .B(n928), .Z(n1287) );
  XNOR U1517 ( .A(n929), .B(n1287), .Z(n3702) );
  XNOR U1518 ( .A(in[160]), .B(n3702), .Z(n4755) );
  XOR U1519 ( .A(in[1280]), .B(in[640]), .Z(n931) );
  XNOR U1520 ( .A(in[960]), .B(in[320]), .Z(n930) );
  XNOR U1521 ( .A(n931), .B(n930), .Z(n932) );
  XOR U1522 ( .A(in[0]), .B(n932), .Z(n1023) );
  XOR U1523 ( .A(in[769]), .B(in[1089]), .Z(n934) );
  XNOR U1524 ( .A(in[449]), .B(in[1409]), .Z(n933) );
  XNOR U1525 ( .A(n934), .B(n933), .Z(n935) );
  XOR U1526 ( .A(in[129]), .B(n935), .Z(n1101) );
  XNOR U1527 ( .A(n1023), .B(n1101), .Z(n4054) );
  XNOR U1528 ( .A(in[1345]), .B(n4054), .Z(n4752) );
  NAND U1529 ( .A(n4755), .B(n4752), .Z(n936) );
  XNOR U1530 ( .A(n1515), .B(n936), .Z(out[1053]) );
  XOR U1531 ( .A(in[1585]), .B(in[625]), .Z(n938) );
  XNOR U1532 ( .A(in[945]), .B(in[305]), .Z(n937) );
  XNOR U1533 ( .A(n938), .B(n937), .Z(n939) );
  XOR U1534 ( .A(in[1265]), .B(n939), .Z(n1418) );
  XNOR U1535 ( .A(n940), .B(n1418), .Z(n3757) );
  XNOR U1536 ( .A(in[561]), .B(n3757), .Z(n1519) );
  XOR U1537 ( .A(in[225]), .B(in[865]), .Z(n942) );
  XNOR U1538 ( .A(in[1185]), .B(in[1505]), .Z(n941) );
  XNOR U1539 ( .A(n942), .B(n941), .Z(n943) );
  XNOR U1540 ( .A(in[545]), .B(n943), .Z(n1290) );
  XNOR U1541 ( .A(n944), .B(n1290), .Z(n3706) );
  XNOR U1542 ( .A(in[161]), .B(n3706), .Z(n4763) );
  XOR U1543 ( .A(in[1]), .B(in[641]), .Z(n946) );
  XNOR U1544 ( .A(in[961]), .B(in[321]), .Z(n945) );
  XNOR U1545 ( .A(n946), .B(n945), .Z(n947) );
  XOR U1546 ( .A(in[1281]), .B(n947), .Z(n1090) );
  XOR U1547 ( .A(in[1090]), .B(in[450]), .Z(n949) );
  XNOR U1548 ( .A(in[130]), .B(in[770]), .Z(n948) );
  XNOR U1549 ( .A(n949), .B(n948), .Z(n950) );
  XOR U1550 ( .A(in[1410]), .B(n950), .Z(n1106) );
  XNOR U1551 ( .A(n1090), .B(n1106), .Z(n4057) );
  XNOR U1552 ( .A(in[1346]), .B(n4057), .Z(n4760) );
  NAND U1553 ( .A(n4763), .B(n4760), .Z(n951) );
  XNOR U1554 ( .A(n1519), .B(n951), .Z(out[1054]) );
  XOR U1555 ( .A(in[1586]), .B(in[626]), .Z(n953) );
  XNOR U1556 ( .A(in[946]), .B(in[306]), .Z(n952) );
  XNOR U1557 ( .A(n953), .B(n952), .Z(n954) );
  XOR U1558 ( .A(in[1266]), .B(n954), .Z(n1422) );
  XNOR U1559 ( .A(n955), .B(n1422), .Z(n3761) );
  XNOR U1560 ( .A(in[562]), .B(n3761), .Z(n1523) );
  XOR U1561 ( .A(in[1186]), .B(in[1506]), .Z(n957) );
  XNOR U1562 ( .A(in[546]), .B(in[866]), .Z(n956) );
  XNOR U1563 ( .A(n957), .B(n956), .Z(n958) );
  XNOR U1564 ( .A(in[226]), .B(n958), .Z(n1293) );
  XNOR U1565 ( .A(n959), .B(n1293), .Z(n3714) );
  XNOR U1566 ( .A(in[162]), .B(n3714), .Z(n4767) );
  XOR U1567 ( .A(in[771]), .B(in[1091]), .Z(n961) );
  XNOR U1568 ( .A(in[451]), .B(in[1411]), .Z(n960) );
  XNOR U1569 ( .A(n961), .B(n960), .Z(n962) );
  XOR U1570 ( .A(in[131]), .B(n962), .Z(n1111) );
  XOR U1571 ( .A(in[2]), .B(in[642]), .Z(n964) );
  XNOR U1572 ( .A(in[962]), .B(in[322]), .Z(n963) );
  XNOR U1573 ( .A(n964), .B(n963), .Z(n965) );
  XOR U1574 ( .A(in[1282]), .B(n965), .Z(n1143) );
  XNOR U1575 ( .A(n1111), .B(n1143), .Z(n4060) );
  XNOR U1576 ( .A(in[1347]), .B(n4060), .Z(n4764) );
  NAND U1577 ( .A(n4767), .B(n4764), .Z(n966) );
  XNOR U1578 ( .A(n1523), .B(n966), .Z(out[1055]) );
  XOR U1579 ( .A(in[1587]), .B(in[627]), .Z(n968) );
  XNOR U1580 ( .A(in[947]), .B(in[307]), .Z(n967) );
  XNOR U1581 ( .A(n968), .B(n967), .Z(n969) );
  XOR U1582 ( .A(in[1267]), .B(n969), .Z(n1427) );
  XNOR U1583 ( .A(n970), .B(n1427), .Z(n3765) );
  XNOR U1584 ( .A(in[563]), .B(n3765), .Z(n1527) );
  XOR U1585 ( .A(in[1187]), .B(in[1507]), .Z(n972) );
  XNOR U1586 ( .A(in[547]), .B(in[867]), .Z(n971) );
  XNOR U1587 ( .A(n972), .B(n971), .Z(n973) );
  XNOR U1588 ( .A(in[227]), .B(n973), .Z(n1296) );
  XNOR U1589 ( .A(n974), .B(n1296), .Z(n3718) );
  XNOR U1590 ( .A(in[163]), .B(n3718), .Z(n4771) );
  XOR U1591 ( .A(in[323]), .B(in[643]), .Z(n976) );
  XNOR U1592 ( .A(in[963]), .B(in[3]), .Z(n975) );
  XNOR U1593 ( .A(n976), .B(n975), .Z(n977) );
  XOR U1594 ( .A(in[1283]), .B(n977), .Z(n1189) );
  XOR U1595 ( .A(in[772]), .B(in[1092]), .Z(n979) );
  XNOR U1596 ( .A(in[452]), .B(in[1412]), .Z(n978) );
  XNOR U1597 ( .A(n979), .B(n978), .Z(n980) );
  XOR U1598 ( .A(in[132]), .B(n980), .Z(n1116) );
  XNOR U1599 ( .A(n1189), .B(n1116), .Z(n4063) );
  XNOR U1600 ( .A(in[1348]), .B(n4063), .Z(n4768) );
  NAND U1601 ( .A(n4771), .B(n4768), .Z(n981) );
  XNOR U1602 ( .A(n1527), .B(n981), .Z(out[1056]) );
  XOR U1603 ( .A(in[1588]), .B(in[628]), .Z(n983) );
  XNOR U1604 ( .A(in[948]), .B(in[308]), .Z(n982) );
  XNOR U1605 ( .A(n983), .B(n982), .Z(n984) );
  XOR U1606 ( .A(in[1268]), .B(n984), .Z(n1431) );
  XNOR U1607 ( .A(n985), .B(n1431), .Z(n3769) );
  XNOR U1608 ( .A(in[564]), .B(n3769), .Z(n1531) );
  XOR U1609 ( .A(in[1188]), .B(in[1508]), .Z(n987) );
  XNOR U1610 ( .A(in[548]), .B(in[868]), .Z(n986) );
  XNOR U1611 ( .A(n987), .B(n986), .Z(n988) );
  XOR U1612 ( .A(in[228]), .B(n988), .Z(n1299) );
  XNOR U1613 ( .A(n1299), .B(n989), .Z(n3722) );
  XNOR U1614 ( .A(in[164]), .B(n3722), .Z(n4775) );
  XOR U1615 ( .A(in[324]), .B(in[644]), .Z(n991) );
  XNOR U1616 ( .A(in[964]), .B(in[4]), .Z(n990) );
  XNOR U1617 ( .A(n991), .B(n990), .Z(n992) );
  XOR U1618 ( .A(in[1284]), .B(n992), .Z(n1197) );
  XOR U1619 ( .A(in[773]), .B(in[1093]), .Z(n994) );
  XNOR U1620 ( .A(in[453]), .B(in[1413]), .Z(n993) );
  XNOR U1621 ( .A(n994), .B(n993), .Z(n995) );
  XOR U1622 ( .A(in[133]), .B(n995), .Z(n1121) );
  XNOR U1623 ( .A(n1197), .B(n1121), .Z(n4066) );
  XNOR U1624 ( .A(in[1349]), .B(n4066), .Z(n4772) );
  NAND U1625 ( .A(n4775), .B(n4772), .Z(n996) );
  XNOR U1626 ( .A(n1531), .B(n996), .Z(out[1057]) );
  XOR U1627 ( .A(in[1589]), .B(in[629]), .Z(n998) );
  XNOR U1628 ( .A(in[949]), .B(in[309]), .Z(n997) );
  XNOR U1629 ( .A(n998), .B(n997), .Z(n999) );
  XOR U1630 ( .A(in[1269]), .B(n999), .Z(n1435) );
  XNOR U1631 ( .A(n1000), .B(n1435), .Z(n3773) );
  XNOR U1632 ( .A(in[565]), .B(n3773), .Z(n1535) );
  XOR U1633 ( .A(in[1189]), .B(in[1509]), .Z(n1002) );
  XNOR U1634 ( .A(in[549]), .B(in[869]), .Z(n1001) );
  XNOR U1635 ( .A(n1002), .B(n1001), .Z(n1003) );
  XNOR U1636 ( .A(in[229]), .B(n1003), .Z(n1303) );
  XNOR U1637 ( .A(n1004), .B(n1303), .Z(n3726) );
  XNOR U1638 ( .A(in[165]), .B(n3726), .Z(n4779) );
  XOR U1639 ( .A(in[774]), .B(in[1094]), .Z(n1006) );
  XNOR U1640 ( .A(in[454]), .B(in[1414]), .Z(n1005) );
  XNOR U1641 ( .A(n1006), .B(n1005), .Z(n1007) );
  XOR U1642 ( .A(in[134]), .B(n1007), .Z(n1126) );
  XOR U1643 ( .A(in[325]), .B(in[645]), .Z(n1009) );
  XNOR U1644 ( .A(in[965]), .B(in[5]), .Z(n1008) );
  XNOR U1645 ( .A(n1009), .B(n1008), .Z(n1010) );
  XOR U1646 ( .A(in[1285]), .B(n1010), .Z(n1200) );
  XNOR U1647 ( .A(n1126), .B(n1200), .Z(n4069) );
  XNOR U1648 ( .A(in[1350]), .B(n4069), .Z(n4776) );
  NAND U1649 ( .A(n4779), .B(n4776), .Z(n1011) );
  XNOR U1650 ( .A(n1535), .B(n1011), .Z(out[1058]) );
  XOR U1651 ( .A(in[1590]), .B(in[630]), .Z(n1013) );
  XNOR U1652 ( .A(in[950]), .B(in[310]), .Z(n1012) );
  XNOR U1653 ( .A(n1013), .B(n1012), .Z(n1014) );
  XOR U1654 ( .A(in[1270]), .B(n1014), .Z(n1439) );
  XNOR U1655 ( .A(n1015), .B(n1439), .Z(n3777) );
  XNOR U1656 ( .A(in[566]), .B(n3777), .Z(n1539) );
  XOR U1657 ( .A(in[166]), .B(n3730), .Z(n4783) );
  XOR U1658 ( .A(in[326]), .B(in[6]), .Z(n1017) );
  XNOR U1659 ( .A(in[966]), .B(in[646]), .Z(n1016) );
  XNOR U1660 ( .A(n1017), .B(n1016), .Z(n1018) );
  XOR U1661 ( .A(in[1286]), .B(n1018), .Z(n1203) );
  XOR U1662 ( .A(in[775]), .B(in[1095]), .Z(n1020) );
  XNOR U1663 ( .A(in[455]), .B(in[1415]), .Z(n1019) );
  XNOR U1664 ( .A(n1020), .B(n1019), .Z(n1021) );
  XOR U1665 ( .A(in[135]), .B(n1021), .Z(n1131) );
  XNOR U1666 ( .A(n1203), .B(n1131), .Z(n4080) );
  XNOR U1667 ( .A(in[1351]), .B(n4080), .Z(n4780) );
  NAND U1668 ( .A(n4783), .B(n4780), .Z(n1022) );
  XNOR U1669 ( .A(n1539), .B(n1022), .Z(out[1059]) );
  XNOR U1670 ( .A(n1024), .B(n1023), .Z(n3612) );
  XNOR U1671 ( .A(in[576]), .B(n3612), .Z(n2561) );
  XOR U1672 ( .A(in[231]), .B(n3713), .Z(n2903) );
  XNOR U1673 ( .A(in[1451]), .B(n3750), .Z(n2900) );
  NAND U1674 ( .A(n2903), .B(n2900), .Z(n1025) );
  XNOR U1675 ( .A(n2561), .B(n1025), .Z(out[105]) );
  XOR U1676 ( .A(in[1591]), .B(in[631]), .Z(n1027) );
  XNOR U1677 ( .A(in[951]), .B(in[311]), .Z(n1026) );
  XNOR U1678 ( .A(n1027), .B(n1026), .Z(n1028) );
  XOR U1679 ( .A(in[1271]), .B(n1028), .Z(n1443) );
  XNOR U1680 ( .A(n1029), .B(n1443), .Z(n3781) );
  XNOR U1681 ( .A(in[567]), .B(n3781), .Z(n1543) );
  XOR U1682 ( .A(in[167]), .B(n3734), .Z(n4787) );
  XOR U1683 ( .A(in[776]), .B(in[1096]), .Z(n1031) );
  XNOR U1684 ( .A(in[456]), .B(in[1416]), .Z(n1030) );
  XNOR U1685 ( .A(n1031), .B(n1030), .Z(n1032) );
  XOR U1686 ( .A(in[136]), .B(n1032), .Z(n1136) );
  XOR U1687 ( .A(in[327]), .B(in[7]), .Z(n1034) );
  XNOR U1688 ( .A(in[967]), .B(in[647]), .Z(n1033) );
  XNOR U1689 ( .A(n1034), .B(n1033), .Z(n1035) );
  XOR U1690 ( .A(in[1287]), .B(n1035), .Z(n1206) );
  XNOR U1691 ( .A(n1136), .B(n1206), .Z(n4083) );
  XNOR U1692 ( .A(in[1352]), .B(n4083), .Z(n4784) );
  NAND U1693 ( .A(n4787), .B(n4784), .Z(n1036) );
  XNOR U1694 ( .A(n1543), .B(n1036), .Z(out[1060]) );
  XOR U1695 ( .A(in[632]), .B(in[1592]), .Z(n1038) );
  XNOR U1696 ( .A(in[1272]), .B(in[312]), .Z(n1037) );
  XNOR U1697 ( .A(n1038), .B(n1037), .Z(n1039) );
  XOR U1698 ( .A(in[952]), .B(n1039), .Z(n1447) );
  XNOR U1699 ( .A(n1040), .B(n1447), .Z(n3785) );
  XNOR U1700 ( .A(in[568]), .B(n3785), .Z(n1547) );
  XOR U1701 ( .A(in[168]), .B(n3738), .Z(n4791) );
  XNOR U1702 ( .A(in[1353]), .B(n4086), .Z(n4788) );
  NAND U1703 ( .A(n4791), .B(n4788), .Z(n1041) );
  XNOR U1704 ( .A(n1547), .B(n1041), .Z(out[1061]) );
  XOR U1705 ( .A(in[633]), .B(in[1593]), .Z(n1043) );
  XNOR U1706 ( .A(in[1273]), .B(in[313]), .Z(n1042) );
  XNOR U1707 ( .A(n1043), .B(n1042), .Z(n1044) );
  XOR U1708 ( .A(in[953]), .B(n1044), .Z(n1451) );
  XNOR U1709 ( .A(n1045), .B(n1451), .Z(n3789) );
  XNOR U1710 ( .A(in[569]), .B(n3789), .Z(n1552) );
  XOR U1711 ( .A(in[169]), .B(n3742), .Z(n4795) );
  XOR U1712 ( .A(in[329]), .B(in[969]), .Z(n1047) );
  XNOR U1713 ( .A(in[9]), .B(in[649]), .Z(n1046) );
  XNOR U1714 ( .A(n1047), .B(n1046), .Z(n1048) );
  XOR U1715 ( .A(in[1289]), .B(n1048), .Z(n1214) );
  XOR U1716 ( .A(in[778]), .B(in[1098]), .Z(n1050) );
  XNOR U1717 ( .A(in[458]), .B(in[1418]), .Z(n1049) );
  XNOR U1718 ( .A(n1050), .B(n1049), .Z(n1051) );
  XOR U1719 ( .A(in[138]), .B(n1051), .Z(n1149) );
  XNOR U1720 ( .A(n1214), .B(n1149), .Z(n4089) );
  XNOR U1721 ( .A(in[1354]), .B(n4089), .Z(n4792) );
  NAND U1722 ( .A(n4795), .B(n4792), .Z(n1052) );
  XNOR U1723 ( .A(n1552), .B(n1052), .Z(out[1062]) );
  XOR U1724 ( .A(in[634]), .B(in[1594]), .Z(n1054) );
  XNOR U1725 ( .A(in[1274]), .B(in[314]), .Z(n1053) );
  XNOR U1726 ( .A(n1054), .B(n1053), .Z(n1055) );
  XOR U1727 ( .A(in[954]), .B(n1055), .Z(n1455) );
  XNOR U1728 ( .A(n1056), .B(n1455), .Z(n3793) );
  XNOR U1729 ( .A(in[570]), .B(n3793), .Z(n1556) );
  XOR U1730 ( .A(in[170]), .B(n3746), .Z(n4799) );
  XOR U1731 ( .A(in[1419]), .B(in[779]), .Z(n1058) );
  XNOR U1732 ( .A(in[1099]), .B(in[459]), .Z(n1057) );
  XNOR U1733 ( .A(n1058), .B(n1057), .Z(n1059) );
  XOR U1734 ( .A(in[139]), .B(n1059), .Z(n1154) );
  XOR U1735 ( .A(in[1290]), .B(in[650]), .Z(n1061) );
  XNOR U1736 ( .A(in[970]), .B(in[330]), .Z(n1060) );
  XNOR U1737 ( .A(n1061), .B(n1060), .Z(n1062) );
  XOR U1738 ( .A(in[10]), .B(n1062), .Z(n1217) );
  XNOR U1739 ( .A(n1154), .B(n1217), .Z(n4092) );
  XNOR U1740 ( .A(in[1355]), .B(n4092), .Z(n4796) );
  NAND U1741 ( .A(n4799), .B(n4796), .Z(n1063) );
  XNOR U1742 ( .A(n1556), .B(n1063), .Z(out[1063]) );
  XOR U1743 ( .A(in[955]), .B(in[1275]), .Z(n1065) );
  XNOR U1744 ( .A(in[1595]), .B(in[315]), .Z(n1064) );
  XNOR U1745 ( .A(n1065), .B(n1064), .Z(n1066) );
  XNOR U1746 ( .A(in[635]), .B(n1066), .Z(n1459) );
  XNOR U1747 ( .A(n1067), .B(n1459), .Z(n3803) );
  XNOR U1748 ( .A(in[571]), .B(n3803), .Z(n1558) );
  NOR U1749 ( .A(n1301), .B(n1696), .Z(n1068) );
  XNOR U1750 ( .A(n1558), .B(n1068), .Z(out[1064]) );
  XOR U1751 ( .A(in[956]), .B(in[1276]), .Z(n1070) );
  XNOR U1752 ( .A(in[1596]), .B(in[316]), .Z(n1069) );
  XNOR U1753 ( .A(n1070), .B(n1069), .Z(n1071) );
  XNOR U1754 ( .A(in[636]), .B(n1071), .Z(n1463) );
  XNOR U1755 ( .A(n1072), .B(n1463), .Z(n3807) );
  XNOR U1756 ( .A(in[572]), .B(n3807), .Z(n1560) );
  NOR U1757 ( .A(n1305), .B(n1700), .Z(n1073) );
  XNOR U1758 ( .A(n1560), .B(n1073), .Z(out[1065]) );
  XOR U1759 ( .A(in[957]), .B(in[1277]), .Z(n1075) );
  XNOR U1760 ( .A(in[1597]), .B(in[317]), .Z(n1074) );
  XNOR U1761 ( .A(n1075), .B(n1074), .Z(n1076) );
  XNOR U1762 ( .A(in[637]), .B(n1076), .Z(n1468) );
  XNOR U1763 ( .A(n1077), .B(n1468), .Z(n3811) );
  XNOR U1764 ( .A(in[573]), .B(n3811), .Z(n1562) );
  NOR U1765 ( .A(n1310), .B(n1704), .Z(n1078) );
  XNOR U1766 ( .A(n1562), .B(n1078), .Z(out[1066]) );
  XOR U1767 ( .A(in[574]), .B(n3815), .Z(n1564) );
  NOR U1768 ( .A(n1314), .B(n1708), .Z(n1079) );
  XNOR U1769 ( .A(n1564), .B(n1079), .Z(out[1067]) );
  XOR U1770 ( .A(in[959]), .B(in[1279]), .Z(n1081) );
  XNOR U1771 ( .A(in[1599]), .B(in[319]), .Z(n1080) );
  XNOR U1772 ( .A(n1081), .B(n1080), .Z(n1082) );
  XNOR U1773 ( .A(in[639]), .B(n1082), .Z(n1476) );
  XNOR U1774 ( .A(n1083), .B(n1476), .Z(n3537) );
  XNOR U1775 ( .A(in[575]), .B(n3537), .Z(n1566) );
  NOR U1776 ( .A(n1318), .B(n1713), .Z(n1084) );
  XNOR U1777 ( .A(n1566), .B(n1084), .Z(out[1068]) );
  XOR U1778 ( .A(in[896]), .B(in[1216]), .Z(n1086) );
  XNOR U1779 ( .A(in[1536]), .B(in[256]), .Z(n1085) );
  XNOR U1780 ( .A(n1086), .B(n1085), .Z(n1087) );
  XNOR U1781 ( .A(in[576]), .B(n1087), .Z(n1480) );
  XNOR U1782 ( .A(n1088), .B(n1480), .Z(n3541) );
  XNOR U1783 ( .A(in[512]), .B(n3541), .Z(n1568) );
  NOR U1784 ( .A(n1322), .B(n1717), .Z(n1089) );
  XNOR U1785 ( .A(n1568), .B(n1089), .Z(out[1069]) );
  XNOR U1786 ( .A(n1091), .B(n1090), .Z(n3616) );
  XNOR U1787 ( .A(in[577]), .B(n3616), .Z(n2563) );
  XOR U1788 ( .A(in[232]), .B(n3717), .Z(n2917) );
  XNOR U1789 ( .A(in[1452]), .B(n3758), .Z(n2914) );
  NAND U1790 ( .A(n2917), .B(n2914), .Z(n1092) );
  XNOR U1791 ( .A(n2563), .B(n1092), .Z(out[106]) );
  XOR U1792 ( .A(in[897]), .B(in[1217]), .Z(n1094) );
  XNOR U1793 ( .A(in[1537]), .B(in[257]), .Z(n1093) );
  XNOR U1794 ( .A(n1094), .B(n1093), .Z(n1095) );
  XNOR U1795 ( .A(in[577]), .B(n1095), .Z(n1484) );
  XNOR U1796 ( .A(n1096), .B(n1484), .Z(n3545) );
  XNOR U1797 ( .A(in[513]), .B(n3545), .Z(n1570) );
  NOR U1798 ( .A(n1326), .B(n1721), .Z(n1097) );
  XNOR U1799 ( .A(n1570), .B(n1097), .Z(out[1070]) );
  XOR U1800 ( .A(in[1538]), .B(in[578]), .Z(n1099) );
  XNOR U1801 ( .A(in[898]), .B(in[258]), .Z(n1098) );
  XNOR U1802 ( .A(n1099), .B(n1098), .Z(n1100) );
  XNOR U1803 ( .A(in[1218]), .B(n1100), .Z(n1488) );
  XNOR U1804 ( .A(n1101), .B(n1488), .Z(n3549) );
  XNOR U1805 ( .A(in[514]), .B(n3549), .Z(n1572) );
  NOR U1806 ( .A(n1330), .B(n1725), .Z(n1102) );
  XNOR U1807 ( .A(n1572), .B(n1102), .Z(out[1071]) );
  XOR U1808 ( .A(in[1539]), .B(in[579]), .Z(n1104) );
  XNOR U1809 ( .A(in[899]), .B(in[259]), .Z(n1103) );
  XNOR U1810 ( .A(n1104), .B(n1103), .Z(n1105) );
  XNOR U1811 ( .A(in[1219]), .B(n1105), .Z(n1492) );
  XNOR U1812 ( .A(n1106), .B(n1492), .Z(n3553) );
  XNOR U1813 ( .A(in[515]), .B(n3553), .Z(n1576) );
  NOR U1814 ( .A(n1334), .B(n1729), .Z(n1107) );
  XNOR U1815 ( .A(n1576), .B(n1107), .Z(out[1072]) );
  XOR U1816 ( .A(in[1540]), .B(in[580]), .Z(n1109) );
  XNOR U1817 ( .A(in[900]), .B(in[260]), .Z(n1108) );
  XNOR U1818 ( .A(n1109), .B(n1108), .Z(n1110) );
  XNOR U1819 ( .A(in[1220]), .B(n1110), .Z(n1496) );
  XNOR U1820 ( .A(n1111), .B(n1496), .Z(n3557) );
  XNOR U1821 ( .A(in[516]), .B(n3557), .Z(n1578) );
  NOR U1822 ( .A(n1338), .B(n1733), .Z(n1112) );
  XNOR U1823 ( .A(n1578), .B(n1112), .Z(out[1073]) );
  XOR U1824 ( .A(in[1541]), .B(in[581]), .Z(n1114) );
  XNOR U1825 ( .A(in[901]), .B(in[261]), .Z(n1113) );
  XNOR U1826 ( .A(n1114), .B(n1113), .Z(n1115) );
  XNOR U1827 ( .A(in[1221]), .B(n1115), .Z(n1500) );
  XNOR U1828 ( .A(n1116), .B(n1500), .Z(n3561) );
  XNOR U1829 ( .A(in[517]), .B(n3561), .Z(n1580) );
  NOR U1830 ( .A(n1342), .B(n1737), .Z(n1117) );
  XNOR U1831 ( .A(n1580), .B(n1117), .Z(out[1074]) );
  XOR U1832 ( .A(in[1542]), .B(in[582]), .Z(n1119) );
  XNOR U1833 ( .A(in[902]), .B(in[262]), .Z(n1118) );
  XNOR U1834 ( .A(n1119), .B(n1118), .Z(n1120) );
  XNOR U1835 ( .A(in[1222]), .B(n1120), .Z(n1504) );
  XNOR U1836 ( .A(n1121), .B(n1504), .Z(n3565) );
  XNOR U1837 ( .A(in[518]), .B(n3565), .Z(n1582) );
  NOR U1838 ( .A(n1346), .B(n1741), .Z(n1122) );
  XNOR U1839 ( .A(n1582), .B(n1122), .Z(out[1075]) );
  XOR U1840 ( .A(in[1543]), .B(in[583]), .Z(n1124) );
  XNOR U1841 ( .A(in[903]), .B(in[263]), .Z(n1123) );
  XNOR U1842 ( .A(n1124), .B(n1123), .Z(n1125) );
  XNOR U1843 ( .A(in[1223]), .B(n1125), .Z(n1509) );
  XNOR U1844 ( .A(n1126), .B(n1509), .Z(n3569) );
  XNOR U1845 ( .A(in[519]), .B(n3569), .Z(n1584) );
  NOR U1846 ( .A(n1351), .B(n1745), .Z(n1127) );
  XNOR U1847 ( .A(n1584), .B(n1127), .Z(out[1076]) );
  XOR U1848 ( .A(in[1544]), .B(in[584]), .Z(n1129) );
  XNOR U1849 ( .A(in[904]), .B(in[264]), .Z(n1128) );
  XNOR U1850 ( .A(n1129), .B(n1128), .Z(n1130) );
  XNOR U1851 ( .A(in[1224]), .B(n1130), .Z(n1513) );
  XNOR U1852 ( .A(n1131), .B(n1513), .Z(n3573) );
  XNOR U1853 ( .A(in[520]), .B(n3573), .Z(n1586) );
  NOR U1854 ( .A(n1355), .B(n1749), .Z(n1132) );
  XNOR U1855 ( .A(n1586), .B(n1132), .Z(out[1077]) );
  XOR U1856 ( .A(in[1545]), .B(in[585]), .Z(n1134) );
  XNOR U1857 ( .A(in[905]), .B(in[265]), .Z(n1133) );
  XNOR U1858 ( .A(n1134), .B(n1133), .Z(n1135) );
  XNOR U1859 ( .A(in[1225]), .B(n1135), .Z(n1517) );
  XNOR U1860 ( .A(n1136), .B(n1517), .Z(n3581) );
  XNOR U1861 ( .A(in[521]), .B(n3581), .Z(n1588) );
  NOR U1862 ( .A(n1359), .B(n1754), .Z(n1137) );
  XNOR U1863 ( .A(n1588), .B(n1137), .Z(out[1078]) );
  XOR U1864 ( .A(in[1546]), .B(in[586]), .Z(n1139) );
  XNOR U1865 ( .A(in[906]), .B(in[266]), .Z(n1138) );
  XNOR U1866 ( .A(n1139), .B(n1138), .Z(n1140) );
  XNOR U1867 ( .A(in[1226]), .B(n1140), .Z(n1521) );
  XNOR U1868 ( .A(n1141), .B(n1521), .Z(n3585) );
  XNOR U1869 ( .A(in[522]), .B(n3585), .Z(n1590) );
  NOR U1870 ( .A(n1363), .B(n1758), .Z(n1142) );
  XNOR U1871 ( .A(n1590), .B(n1142), .Z(out[1079]) );
  XNOR U1872 ( .A(n1144), .B(n1143), .Z(n3624) );
  XNOR U1873 ( .A(in[578]), .B(n3624), .Z(n2565) );
  XOR U1874 ( .A(in[233]), .B(n3721), .Z(n2931) );
  XNOR U1875 ( .A(in[1453]), .B(n3762), .Z(n2928) );
  NAND U1876 ( .A(n2931), .B(n2928), .Z(n1145) );
  XNOR U1877 ( .A(n2565), .B(n1145), .Z(out[107]) );
  XOR U1878 ( .A(in[1547]), .B(in[587]), .Z(n1147) );
  XNOR U1879 ( .A(in[907]), .B(in[267]), .Z(n1146) );
  XNOR U1880 ( .A(n1147), .B(n1146), .Z(n1148) );
  XNOR U1881 ( .A(in[1227]), .B(n1148), .Z(n1525) );
  XNOR U1882 ( .A(n1149), .B(n1525), .Z(n3589) );
  XNOR U1883 ( .A(in[523]), .B(n3589), .Z(n1592) );
  NOR U1884 ( .A(n1367), .B(n1762), .Z(n1150) );
  XNOR U1885 ( .A(n1592), .B(n1150), .Z(out[1080]) );
  XOR U1886 ( .A(in[1548]), .B(in[588]), .Z(n1152) );
  XNOR U1887 ( .A(in[908]), .B(in[268]), .Z(n1151) );
  XNOR U1888 ( .A(n1152), .B(n1151), .Z(n1153) );
  XNOR U1889 ( .A(in[1228]), .B(n1153), .Z(n1529) );
  XNOR U1890 ( .A(n1154), .B(n1529), .Z(n3593) );
  XNOR U1891 ( .A(in[524]), .B(n3593), .Z(n1594) );
  NOR U1892 ( .A(n1371), .B(n1766), .Z(n1155) );
  XNOR U1893 ( .A(n1594), .B(n1155), .Z(out[1081]) );
  XOR U1894 ( .A(in[1549]), .B(in[589]), .Z(n1157) );
  XNOR U1895 ( .A(in[909]), .B(in[269]), .Z(n1156) );
  XNOR U1896 ( .A(n1157), .B(n1156), .Z(n1158) );
  XNOR U1897 ( .A(in[1229]), .B(n1158), .Z(n1533) );
  XNOR U1898 ( .A(n1159), .B(n1533), .Z(n3597) );
  XNOR U1899 ( .A(in[525]), .B(n3597), .Z(n1597) );
  NOR U1900 ( .A(n1375), .B(n1770), .Z(n1160) );
  XNOR U1901 ( .A(n1597), .B(n1160), .Z(out[1082]) );
  XOR U1902 ( .A(in[1550]), .B(in[590]), .Z(n1162) );
  XNOR U1903 ( .A(in[910]), .B(in[270]), .Z(n1161) );
  XNOR U1904 ( .A(n1162), .B(n1161), .Z(n1163) );
  XOR U1905 ( .A(in[1230]), .B(n1163), .Z(n1537) );
  XNOR U1906 ( .A(n1537), .B(n1164), .Z(n3601) );
  XNOR U1907 ( .A(in[526]), .B(n3601), .Z(n1599) );
  NOR U1908 ( .A(n1379), .B(n1774), .Z(n1165) );
  XNOR U1909 ( .A(n1599), .B(n1165), .Z(out[1083]) );
  XOR U1910 ( .A(in[1551]), .B(in[591]), .Z(n1167) );
  XNOR U1911 ( .A(in[911]), .B(in[271]), .Z(n1166) );
  XNOR U1912 ( .A(n1167), .B(n1166), .Z(n1168) );
  XOR U1913 ( .A(in[1231]), .B(n1168), .Z(n1541) );
  XNOR U1914 ( .A(n1541), .B(n1169), .Z(n3605) );
  XNOR U1915 ( .A(in[527]), .B(n3605), .Z(n1601) );
  NOR U1916 ( .A(n1383), .B(n1778), .Z(n1170) );
  XNOR U1917 ( .A(n1601), .B(n1170), .Z(out[1084]) );
  XOR U1918 ( .A(in[1552]), .B(in[592]), .Z(n1172) );
  XNOR U1919 ( .A(in[912]), .B(in[272]), .Z(n1171) );
  XNOR U1920 ( .A(n1172), .B(n1171), .Z(n1173) );
  XNOR U1921 ( .A(in[1232]), .B(n1173), .Z(n1545) );
  XNOR U1922 ( .A(n1174), .B(n1545), .Z(n3609) );
  XNOR U1923 ( .A(in[528]), .B(n3609), .Z(n1603) );
  NOR U1924 ( .A(n1387), .B(n1782), .Z(n1175) );
  XNOR U1925 ( .A(n1603), .B(n1175), .Z(out[1085]) );
  XOR U1926 ( .A(in[1553]), .B(in[593]), .Z(n1177) );
  XNOR U1927 ( .A(in[913]), .B(in[273]), .Z(n1176) );
  XNOR U1928 ( .A(n1177), .B(n1176), .Z(n1178) );
  XNOR U1929 ( .A(in[1233]), .B(n1178), .Z(n1550) );
  XNOR U1930 ( .A(n1179), .B(n1550), .Z(n3613) );
  XNOR U1931 ( .A(in[529]), .B(n3613), .Z(n1605) );
  NOR U1932 ( .A(n1390), .B(n1786), .Z(n1180) );
  XNOR U1933 ( .A(n1605), .B(n1180), .Z(out[1086]) );
  XOR U1934 ( .A(in[1554]), .B(in[594]), .Z(n1182) );
  XNOR U1935 ( .A(in[914]), .B(in[274]), .Z(n1181) );
  XNOR U1936 ( .A(n1182), .B(n1181), .Z(n1183) );
  XOR U1937 ( .A(in[1234]), .B(n1183), .Z(n1554) );
  XNOR U1938 ( .A(n1554), .B(n1184), .Z(n3617) );
  XNOR U1939 ( .A(in[530]), .B(n3617), .Z(n1607) );
  NOR U1940 ( .A(n1392), .B(n1790), .Z(n1185) );
  XNOR U1941 ( .A(n1607), .B(n1185), .Z(out[1087]) );
  XOR U1942 ( .A(in[957]), .B(n3600), .Z(n1609) );
  NOR U1943 ( .A(n1396), .B(n4631), .Z(n1186) );
  XNOR U1944 ( .A(n1609), .B(n1186), .Z(out[1088]) );
  XOR U1945 ( .A(in[958]), .B(n3604), .Z(n1611) );
  NOR U1946 ( .A(n1400), .B(n4635), .Z(n1187) );
  XNOR U1947 ( .A(n1611), .B(n1187), .Z(out[1089]) );
  XOR U1948 ( .A(n1189), .B(n1188), .Z(n3628) );
  XNOR U1949 ( .A(in[579]), .B(n3628), .Z(n2567) );
  XOR U1950 ( .A(in[234]), .B(n3725), .Z(n2947) );
  XNOR U1951 ( .A(in[1454]), .B(n3766), .Z(n2944) );
  NAND U1952 ( .A(n2947), .B(n2944), .Z(n1190) );
  XNOR U1953 ( .A(n2567), .B(n1190), .Z(out[108]) );
  XOR U1954 ( .A(in[959]), .B(n3608), .Z(n1613) );
  NOR U1955 ( .A(n1404), .B(n4639), .Z(n1191) );
  XNOR U1956 ( .A(n1613), .B(n1191), .Z(out[1090]) );
  XOR U1957 ( .A(in[896]), .B(n3612), .Z(n1615) );
  NOR U1958 ( .A(n1408), .B(n4643), .Z(n1192) );
  XNOR U1959 ( .A(n1615), .B(n1192), .Z(out[1091]) );
  XOR U1960 ( .A(in[897]), .B(n3616), .Z(n1618) );
  NOR U1961 ( .A(n1412), .B(n4647), .Z(n1193) );
  XNOR U1962 ( .A(n1618), .B(n1193), .Z(out[1092]) );
  XOR U1963 ( .A(in[898]), .B(n3624), .Z(n1620) );
  NOR U1964 ( .A(n1416), .B(n4651), .Z(n1194) );
  XNOR U1965 ( .A(n1620), .B(n1194), .Z(out[1093]) );
  XOR U1966 ( .A(in[899]), .B(n3628), .Z(n1622) );
  NOR U1967 ( .A(n1420), .B(n4655), .Z(n1195) );
  XNOR U1968 ( .A(n1622), .B(n1195), .Z(out[1094]) );
  XNOR U1969 ( .A(n1197), .B(n1196), .Z(n3632) );
  XNOR U1970 ( .A(in[900]), .B(n3632), .Z(n1624) );
  NOR U1971 ( .A(n1424), .B(n4659), .Z(n1198) );
  XNOR U1972 ( .A(n1624), .B(n1198), .Z(out[1095]) );
  XNOR U1973 ( .A(n1200), .B(n1199), .Z(n3636) );
  XNOR U1974 ( .A(in[901]), .B(n3636), .Z(n1626) );
  NOR U1975 ( .A(n1429), .B(n4663), .Z(n1201) );
  XNOR U1976 ( .A(n1626), .B(n1201), .Z(out[1096]) );
  XNOR U1977 ( .A(n1203), .B(n1202), .Z(n3640) );
  XNOR U1978 ( .A(in[902]), .B(n3640), .Z(n1628) );
  NOR U1979 ( .A(n1433), .B(n4667), .Z(n1204) );
  XNOR U1980 ( .A(n1628), .B(n1204), .Z(out[1097]) );
  XNOR U1981 ( .A(n1206), .B(n1205), .Z(n3644) );
  XNOR U1982 ( .A(in[903]), .B(n3644), .Z(n1630) );
  NOR U1983 ( .A(n1437), .B(n4675), .Z(n1207) );
  XNOR U1984 ( .A(n1630), .B(n1207), .Z(out[1098]) );
  XNOR U1985 ( .A(n1209), .B(n1208), .Z(n3648) );
  XNOR U1986 ( .A(in[904]), .B(n3648), .Z(n1632) );
  NOR U1987 ( .A(n1441), .B(n4679), .Z(n1210) );
  XNOR U1988 ( .A(n1632), .B(n1210), .Z(out[1099]) );
  XOR U1989 ( .A(in[580]), .B(n3632), .Z(n2569) );
  XOR U1990 ( .A(in[235]), .B(n3729), .Z(n2971) );
  XNOR U1991 ( .A(in[1455]), .B(n3770), .Z(n2968) );
  NAND U1992 ( .A(n2971), .B(n2968), .Z(n1211) );
  XNOR U1993 ( .A(n2569), .B(n1211), .Z(out[109]) );
  XOR U1994 ( .A(in[200]), .B(n3573), .Z(n3921) );
  XNOR U1995 ( .A(in[1420]), .B(n3614), .Z(n3920) );
  XOR U1996 ( .A(n4120), .B(in[1043]), .Z(n2632) );
  NAND U1997 ( .A(n3920), .B(n2632), .Z(n1212) );
  XNOR U1998 ( .A(n3921), .B(n1212), .Z(out[10]) );
  XNOR U1999 ( .A(n1214), .B(n1213), .Z(n3652) );
  XNOR U2000 ( .A(in[905]), .B(n3652), .Z(n1634) );
  NOR U2001 ( .A(n1445), .B(n4683), .Z(n1215) );
  XNOR U2002 ( .A(n1634), .B(n1215), .Z(out[1100]) );
  XNOR U2003 ( .A(n1217), .B(n1216), .Z(n3656) );
  XNOR U2004 ( .A(in[906]), .B(n3656), .Z(n1636) );
  NOR U2005 ( .A(n1449), .B(n4687), .Z(n1218) );
  XNOR U2006 ( .A(n1636), .B(n1218), .Z(out[1101]) );
  XOR U2007 ( .A(n1220), .B(n1219), .Z(n3660) );
  XNOR U2008 ( .A(in[907]), .B(n3660), .Z(n1639) );
  NOR U2009 ( .A(n1453), .B(n4691), .Z(n1221) );
  XNOR U2010 ( .A(n1639), .B(n1221), .Z(out[1102]) );
  XOR U2011 ( .A(n1223), .B(n1222), .Z(n3668) );
  XNOR U2012 ( .A(in[908]), .B(n3668), .Z(n1641) );
  NOR U2013 ( .A(n1457), .B(n4695), .Z(n1224) );
  XNOR U2014 ( .A(n1641), .B(n1224), .Z(out[1103]) );
  XNOR U2015 ( .A(n1226), .B(n1225), .Z(n3672) );
  XNOR U2016 ( .A(in[909]), .B(n3672), .Z(n1643) );
  NOR U2017 ( .A(n1461), .B(n4699), .Z(n1227) );
  XNOR U2018 ( .A(n1643), .B(n1227), .Z(out[1104]) );
  XOR U2019 ( .A(n1229), .B(n1228), .Z(n3676) );
  XNOR U2020 ( .A(in[910]), .B(n3676), .Z(n1645) );
  NOR U2021 ( .A(n1465), .B(n4703), .Z(n1230) );
  XNOR U2022 ( .A(n1645), .B(n1230), .Z(out[1105]) );
  XOR U2023 ( .A(n1232), .B(n1231), .Z(n3680) );
  XNOR U2024 ( .A(in[911]), .B(n3680), .Z(n1647) );
  NOR U2025 ( .A(n1470), .B(n4707), .Z(n1233) );
  XNOR U2026 ( .A(n1647), .B(n1233), .Z(out[1106]) );
  XNOR U2027 ( .A(n1235), .B(n1234), .Z(n3684) );
  XNOR U2028 ( .A(in[912]), .B(n3684), .Z(n1649) );
  NOR U2029 ( .A(n1474), .B(n4711), .Z(n1236) );
  XNOR U2030 ( .A(n1649), .B(n1236), .Z(out[1107]) );
  XOR U2031 ( .A(n1238), .B(n1237), .Z(n3688) );
  XNOR U2032 ( .A(in[913]), .B(n3688), .Z(n1651) );
  NOR U2033 ( .A(n1478), .B(n4719), .Z(n1239) );
  XNOR U2034 ( .A(n1651), .B(n1239), .Z(out[1108]) );
  XNOR U2035 ( .A(n1241), .B(n1240), .Z(n3692) );
  XNOR U2036 ( .A(in[914]), .B(n3692), .Z(n1653) );
  NOR U2037 ( .A(n1482), .B(n4723), .Z(n1242) );
  XNOR U2038 ( .A(n1653), .B(n1242), .Z(out[1109]) );
  XOR U2039 ( .A(in[581]), .B(n3636), .Z(n2571) );
  XOR U2040 ( .A(in[236]), .B(n3733), .Z(n2995) );
  XNOR U2041 ( .A(in[1456]), .B(n3774), .Z(n2992) );
  NAND U2042 ( .A(n2995), .B(n2992), .Z(n1243) );
  XNOR U2043 ( .A(n2571), .B(n1243), .Z(out[110]) );
  XOR U2044 ( .A(n1245), .B(n1244), .Z(n3696) );
  XNOR U2045 ( .A(in[915]), .B(n3696), .Z(n1655) );
  NOR U2046 ( .A(n1486), .B(n4727), .Z(n1246) );
  XNOR U2047 ( .A(n1655), .B(n1246), .Z(out[1110]) );
  XNOR U2048 ( .A(n1248), .B(n1247), .Z(n3700) );
  XNOR U2049 ( .A(in[916]), .B(n3700), .Z(n1657) );
  NOR U2050 ( .A(n1490), .B(n4731), .Z(n1249) );
  XNOR U2051 ( .A(n1657), .B(n1249), .Z(out[1111]) );
  XNOR U2052 ( .A(n1251), .B(n1250), .Z(n3704) );
  XNOR U2053 ( .A(in[917]), .B(n3704), .Z(n1660) );
  NOR U2054 ( .A(n1494), .B(n4735), .Z(n1252) );
  XNOR U2055 ( .A(n1660), .B(n1252), .Z(out[1112]) );
  XOR U2056 ( .A(n1254), .B(n1253), .Z(n3712) );
  XNOR U2057 ( .A(in[918]), .B(n3712), .Z(n1662) );
  NOR U2058 ( .A(n1498), .B(n4739), .Z(n1255) );
  XNOR U2059 ( .A(n1662), .B(n1255), .Z(out[1113]) );
  XNOR U2060 ( .A(n1257), .B(n1256), .Z(n3716) );
  XNOR U2061 ( .A(in[919]), .B(n3716), .Z(n1664) );
  NOR U2062 ( .A(n1502), .B(n4743), .Z(n1258) );
  XNOR U2063 ( .A(n1664), .B(n1258), .Z(out[1114]) );
  XOR U2064 ( .A(n1260), .B(n1259), .Z(n3720) );
  XNOR U2065 ( .A(in[920]), .B(n3720), .Z(n1666) );
  NOR U2066 ( .A(n1506), .B(n4747), .Z(n1261) );
  XNOR U2067 ( .A(n1666), .B(n1261), .Z(out[1115]) );
  XNOR U2068 ( .A(n1263), .B(n1262), .Z(n3724) );
  XNOR U2069 ( .A(in[921]), .B(n3724), .Z(n1668) );
  NOR U2070 ( .A(n1511), .B(n4751), .Z(n1264) );
  XNOR U2071 ( .A(n1668), .B(n1264), .Z(out[1116]) );
  XOR U2072 ( .A(n1266), .B(n1265), .Z(n3728) );
  XNOR U2073 ( .A(in[922]), .B(n3728), .Z(n1670) );
  NOR U2074 ( .A(n1515), .B(n4755), .Z(n1267) );
  XNOR U2075 ( .A(n1670), .B(n1267), .Z(out[1117]) );
  XOR U2076 ( .A(n1269), .B(n1268), .Z(n3732) );
  XNOR U2077 ( .A(in[923]), .B(n3732), .Z(n1672) );
  NOR U2078 ( .A(n1519), .B(n4763), .Z(n1270) );
  XNOR U2079 ( .A(n1672), .B(n1270), .Z(out[1118]) );
  XOR U2080 ( .A(n1272), .B(n1271), .Z(n3736) );
  XNOR U2081 ( .A(in[924]), .B(n3736), .Z(n1674) );
  NOR U2082 ( .A(n1523), .B(n4767), .Z(n1273) );
  XNOR U2083 ( .A(n1674), .B(n1273), .Z(out[1119]) );
  XOR U2084 ( .A(in[582]), .B(n3640), .Z(n2573) );
  XOR U2085 ( .A(in[237]), .B(n3737), .Z(n3019) );
  XNOR U2086 ( .A(in[1457]), .B(n3778), .Z(n3016) );
  NAND U2087 ( .A(n3019), .B(n3016), .Z(n1274) );
  XNOR U2088 ( .A(n2573), .B(n1274), .Z(out[111]) );
  XOR U2089 ( .A(n1276), .B(n1275), .Z(n3740) );
  XNOR U2090 ( .A(in[925]), .B(n3740), .Z(n1676) );
  NOR U2091 ( .A(n1527), .B(n4771), .Z(n1277) );
  XNOR U2092 ( .A(n1676), .B(n1277), .Z(out[1120]) );
  XOR U2093 ( .A(n1279), .B(n1278), .Z(n3744) );
  XNOR U2094 ( .A(in[926]), .B(n3744), .Z(n1678) );
  NOR U2095 ( .A(n1531), .B(n4775), .Z(n1280) );
  XNOR U2096 ( .A(n1678), .B(n1280), .Z(out[1121]) );
  XOR U2097 ( .A(n1282), .B(n1281), .Z(n3748) );
  XNOR U2098 ( .A(in[927]), .B(n3748), .Z(n1681) );
  NOR U2099 ( .A(n1535), .B(n4779), .Z(n1283) );
  XNOR U2100 ( .A(n1681), .B(n1283), .Z(out[1122]) );
  XOR U2101 ( .A(n1285), .B(n1284), .Z(n3756) );
  XNOR U2102 ( .A(in[928]), .B(n3756), .Z(n1683) );
  NOR U2103 ( .A(n1539), .B(n4783), .Z(n1286) );
  XNOR U2104 ( .A(n1683), .B(n1286), .Z(out[1123]) );
  XNOR U2105 ( .A(n1288), .B(n1287), .Z(n3760) );
  XNOR U2106 ( .A(in[929]), .B(n3760), .Z(n1685) );
  NOR U2107 ( .A(n1543), .B(n4787), .Z(n1289) );
  XNOR U2108 ( .A(n1685), .B(n1289), .Z(out[1124]) );
  XOR U2109 ( .A(n1291), .B(n1290), .Z(n3764) );
  XNOR U2110 ( .A(in[930]), .B(n3764), .Z(n1687) );
  NOR U2111 ( .A(n1547), .B(n4791), .Z(n1292) );
  XNOR U2112 ( .A(n1687), .B(n1292), .Z(out[1125]) );
  XNOR U2113 ( .A(n1294), .B(n1293), .Z(n3768) );
  XNOR U2114 ( .A(in[931]), .B(n3768), .Z(n1689) );
  NOR U2115 ( .A(n1552), .B(n4795), .Z(n1295) );
  XNOR U2116 ( .A(n1689), .B(n1295), .Z(out[1126]) );
  XNOR U2117 ( .A(n1297), .B(n1296), .Z(n3772) );
  XNOR U2118 ( .A(in[932]), .B(n3772), .Z(n1691) );
  NOR U2119 ( .A(n1556), .B(n4799), .Z(n1298) );
  XNOR U2120 ( .A(n1691), .B(n1298), .Z(out[1127]) );
  XNOR U2121 ( .A(n1300), .B(n1299), .Z(n3776) );
  XNOR U2122 ( .A(in[933]), .B(n3776), .Z(n1694) );
  NAND U2123 ( .A(n1558), .B(n1301), .Z(n1302) );
  XNOR U2124 ( .A(n1694), .B(n1302), .Z(out[1128]) );
  XOR U2125 ( .A(n1304), .B(n1303), .Z(n3780) );
  XNOR U2126 ( .A(in[934]), .B(n3780), .Z(n1698) );
  NAND U2127 ( .A(n1560), .B(n1305), .Z(n1306) );
  XNOR U2128 ( .A(n1698), .B(n1306), .Z(out[1129]) );
  XOR U2129 ( .A(in[583]), .B(n3644), .Z(n2576) );
  XOR U2130 ( .A(in[238]), .B(n3741), .Z(n3043) );
  XNOR U2131 ( .A(in[1458]), .B(n3782), .Z(n3040) );
  NAND U2132 ( .A(n3043), .B(n3040), .Z(n1307) );
  XNOR U2133 ( .A(n2576), .B(n1307), .Z(out[112]) );
  XNOR U2134 ( .A(n1309), .B(n1308), .Z(n3784) );
  XNOR U2135 ( .A(in[935]), .B(n3784), .Z(n1702) );
  NAND U2136 ( .A(n1562), .B(n1310), .Z(n1311) );
  XNOR U2137 ( .A(n1702), .B(n1311), .Z(out[1130]) );
  XNOR U2138 ( .A(n1313), .B(n1312), .Z(n3788) );
  XNOR U2139 ( .A(in[936]), .B(n3788), .Z(n1706) );
  NAND U2140 ( .A(n1564), .B(n1314), .Z(n1315) );
  XNOR U2141 ( .A(n1706), .B(n1315), .Z(out[1131]) );
  XNOR U2142 ( .A(n1317), .B(n1316), .Z(n3792) );
  XNOR U2143 ( .A(in[937]), .B(n3792), .Z(n1711) );
  NAND U2144 ( .A(n1566), .B(n1318), .Z(n1319) );
  XNOR U2145 ( .A(n1711), .B(n1319), .Z(out[1132]) );
  XNOR U2146 ( .A(n1321), .B(n1320), .Z(n3802) );
  XNOR U2147 ( .A(in[938]), .B(n3802), .Z(n1715) );
  NAND U2148 ( .A(n1568), .B(n1322), .Z(n1323) );
  XNOR U2149 ( .A(n1715), .B(n1323), .Z(out[1133]) );
  XNOR U2150 ( .A(n1325), .B(n1324), .Z(n3806) );
  XNOR U2151 ( .A(in[939]), .B(n3806), .Z(n1719) );
  NAND U2152 ( .A(n1570), .B(n1326), .Z(n1327) );
  XNOR U2153 ( .A(n1719), .B(n1327), .Z(out[1134]) );
  XNOR U2154 ( .A(n1329), .B(n1328), .Z(n3810) );
  XNOR U2155 ( .A(in[940]), .B(n3810), .Z(n1723) );
  NAND U2156 ( .A(n1572), .B(n1330), .Z(n1331) );
  XNOR U2157 ( .A(n1723), .B(n1331), .Z(out[1135]) );
  XNOR U2158 ( .A(n1333), .B(n1332), .Z(n3814) );
  XNOR U2159 ( .A(in[941]), .B(n3814), .Z(n1727) );
  NAND U2160 ( .A(n1576), .B(n1334), .Z(n1335) );
  XNOR U2161 ( .A(n1727), .B(n1335), .Z(out[1136]) );
  XNOR U2162 ( .A(n1337), .B(n1336), .Z(n3536) );
  XNOR U2163 ( .A(in[942]), .B(n3536), .Z(n1731) );
  NAND U2164 ( .A(n1578), .B(n1338), .Z(n1339) );
  XNOR U2165 ( .A(n1731), .B(n1339), .Z(out[1137]) );
  XNOR U2166 ( .A(n1341), .B(n1340), .Z(n3540) );
  XNOR U2167 ( .A(in[943]), .B(n3540), .Z(n1735) );
  NAND U2168 ( .A(n1580), .B(n1342), .Z(n1343) );
  XNOR U2169 ( .A(n1735), .B(n1343), .Z(out[1138]) );
  XNOR U2170 ( .A(n1345), .B(n1344), .Z(n3544) );
  XNOR U2171 ( .A(in[944]), .B(n3544), .Z(n1739) );
  NAND U2172 ( .A(n1582), .B(n1346), .Z(n1347) );
  XNOR U2173 ( .A(n1739), .B(n1347), .Z(out[1139]) );
  XOR U2174 ( .A(in[584]), .B(n3648), .Z(n2578) );
  XOR U2175 ( .A(in[239]), .B(n3745), .Z(n3067) );
  XNOR U2176 ( .A(in[1459]), .B(n3786), .Z(n3064) );
  NAND U2177 ( .A(n3067), .B(n3064), .Z(n1348) );
  XNOR U2178 ( .A(n2578), .B(n1348), .Z(out[113]) );
  XNOR U2179 ( .A(n1350), .B(n1349), .Z(n3548) );
  XNOR U2180 ( .A(in[945]), .B(n3548), .Z(n1743) );
  NAND U2181 ( .A(n1584), .B(n1351), .Z(n1352) );
  XNOR U2182 ( .A(n1743), .B(n1352), .Z(out[1140]) );
  XNOR U2183 ( .A(n1354), .B(n1353), .Z(n3552) );
  XNOR U2184 ( .A(in[946]), .B(n3552), .Z(n1747) );
  NAND U2185 ( .A(n1586), .B(n1355), .Z(n1356) );
  XNOR U2186 ( .A(n1747), .B(n1356), .Z(out[1141]) );
  XNOR U2187 ( .A(n1358), .B(n1357), .Z(n3556) );
  XNOR U2188 ( .A(in[947]), .B(n3556), .Z(n1752) );
  NAND U2189 ( .A(n1588), .B(n1359), .Z(n1360) );
  XNOR U2190 ( .A(n1752), .B(n1360), .Z(out[1142]) );
  XNOR U2191 ( .A(n1362), .B(n1361), .Z(n3560) );
  XNOR U2192 ( .A(in[948]), .B(n3560), .Z(n1756) );
  NAND U2193 ( .A(n1590), .B(n1363), .Z(n1364) );
  XNOR U2194 ( .A(n1756), .B(n1364), .Z(out[1143]) );
  XNOR U2195 ( .A(n1366), .B(n1365), .Z(n3564) );
  XNOR U2196 ( .A(in[949]), .B(n3564), .Z(n1760) );
  NAND U2197 ( .A(n1592), .B(n1367), .Z(n1368) );
  XNOR U2198 ( .A(n1760), .B(n1368), .Z(out[1144]) );
  XNOR U2199 ( .A(n1370), .B(n1369), .Z(n3568) );
  XNOR U2200 ( .A(in[950]), .B(n3568), .Z(n1764) );
  NAND U2201 ( .A(n1594), .B(n1371), .Z(n1372) );
  XNOR U2202 ( .A(n1764), .B(n1372), .Z(out[1145]) );
  XNOR U2203 ( .A(n1374), .B(n1373), .Z(n3572) );
  XNOR U2204 ( .A(in[951]), .B(n3572), .Z(n1768) );
  NAND U2205 ( .A(n1597), .B(n1375), .Z(n1376) );
  XNOR U2206 ( .A(n1768), .B(n1376), .Z(out[1146]) );
  XNOR U2207 ( .A(n1378), .B(n1377), .Z(n3580) );
  XNOR U2208 ( .A(in[952]), .B(n3580), .Z(n1772) );
  NAND U2209 ( .A(n1599), .B(n1379), .Z(n1380) );
  XNOR U2210 ( .A(n1772), .B(n1380), .Z(out[1147]) );
  XNOR U2211 ( .A(n1382), .B(n1381), .Z(n3584) );
  XNOR U2212 ( .A(in[953]), .B(n3584), .Z(n1776) );
  NAND U2213 ( .A(n1601), .B(n1383), .Z(n1384) );
  XNOR U2214 ( .A(n1776), .B(n1384), .Z(out[1148]) );
  XNOR U2215 ( .A(n1386), .B(n1385), .Z(n3588) );
  XNOR U2216 ( .A(in[954]), .B(n3588), .Z(n1780) );
  NAND U2217 ( .A(n1603), .B(n1387), .Z(n1388) );
  XNOR U2218 ( .A(n1780), .B(n1388), .Z(out[1149]) );
  XOR U2219 ( .A(in[585]), .B(n3652), .Z(n2580) );
  XOR U2220 ( .A(in[240]), .B(n3749), .Z(n3093) );
  XNOR U2221 ( .A(in[1460]), .B(n3790), .Z(n3090) );
  NAND U2222 ( .A(n3093), .B(n3090), .Z(n1389) );
  XNOR U2223 ( .A(n2580), .B(n1389), .Z(out[114]) );
  XNOR U2224 ( .A(in[955]), .B(n3592), .Z(n1784) );
  NAND U2225 ( .A(n1605), .B(n1390), .Z(n1391) );
  XNOR U2226 ( .A(n1784), .B(n1391), .Z(out[1150]) );
  XNOR U2227 ( .A(in[956]), .B(n3596), .Z(n1788) );
  NAND U2228 ( .A(n1607), .B(n1392), .Z(n1393) );
  XNOR U2229 ( .A(n1788), .B(n1393), .Z(out[1151]) );
  XNOR U2230 ( .A(n1395), .B(n1394), .Z(n3936) );
  XNOR U2231 ( .A(in[1004]), .B(n3936), .Z(n4629) );
  NAND U2232 ( .A(n1609), .B(n1396), .Z(n1397) );
  XNOR U2233 ( .A(n4629), .B(n1397), .Z(out[1152]) );
  XNOR U2234 ( .A(n1399), .B(n1398), .Z(n3938) );
  XNOR U2235 ( .A(in[1005]), .B(n3938), .Z(n4633) );
  NAND U2236 ( .A(n1611), .B(n1400), .Z(n1401) );
  XNOR U2237 ( .A(n4633), .B(n1401), .Z(out[1153]) );
  XNOR U2238 ( .A(n1403), .B(n1402), .Z(n3940) );
  XNOR U2239 ( .A(in[1006]), .B(n3940), .Z(n4637) );
  NAND U2240 ( .A(n1613), .B(n1404), .Z(n1405) );
  XNOR U2241 ( .A(n4637), .B(n1405), .Z(out[1154]) );
  XNOR U2242 ( .A(n1407), .B(n1406), .Z(n3942) );
  XNOR U2243 ( .A(in[1007]), .B(n3942), .Z(n4641) );
  NAND U2244 ( .A(n1615), .B(n1408), .Z(n1409) );
  XNOR U2245 ( .A(n4641), .B(n1409), .Z(out[1155]) );
  XNOR U2246 ( .A(n1411), .B(n1410), .Z(n3948) );
  XNOR U2247 ( .A(in[1008]), .B(n3948), .Z(n4645) );
  NAND U2248 ( .A(n1618), .B(n1412), .Z(n1413) );
  XNOR U2249 ( .A(n4645), .B(n1413), .Z(out[1156]) );
  XNOR U2250 ( .A(n1415), .B(n1414), .Z(n3950) );
  XNOR U2251 ( .A(in[1009]), .B(n3950), .Z(n4649) );
  NAND U2252 ( .A(n1620), .B(n1416), .Z(n1417) );
  XNOR U2253 ( .A(n4649), .B(n1417), .Z(out[1157]) );
  XNOR U2254 ( .A(n1419), .B(n1418), .Z(n3952) );
  XNOR U2255 ( .A(in[1010]), .B(n3952), .Z(n4653) );
  NAND U2256 ( .A(n1622), .B(n1420), .Z(n1421) );
  XNOR U2257 ( .A(n4653), .B(n1421), .Z(out[1158]) );
  XNOR U2258 ( .A(n1423), .B(n1422), .Z(n3954) );
  XNOR U2259 ( .A(in[1011]), .B(n3954), .Z(n4657) );
  NAND U2260 ( .A(n1624), .B(n1424), .Z(n1425) );
  XNOR U2261 ( .A(n4657), .B(n1425), .Z(out[1159]) );
  XOR U2262 ( .A(in[586]), .B(n3656), .Z(n2582) );
  XOR U2263 ( .A(in[241]), .B(n3757), .Z(n3117) );
  XNOR U2264 ( .A(in[1461]), .B(n3794), .Z(n3114) );
  NAND U2265 ( .A(n3117), .B(n3114), .Z(n1426) );
  XNOR U2266 ( .A(n2582), .B(n1426), .Z(out[115]) );
  XNOR U2267 ( .A(n1428), .B(n1427), .Z(n3956) );
  XNOR U2268 ( .A(in[1012]), .B(n3956), .Z(n4661) );
  NAND U2269 ( .A(n1626), .B(n1429), .Z(n1430) );
  XNOR U2270 ( .A(n4661), .B(n1430), .Z(out[1160]) );
  XNOR U2271 ( .A(n1432), .B(n1431), .Z(n3958) );
  XNOR U2272 ( .A(in[1013]), .B(n3958), .Z(n4665) );
  NAND U2273 ( .A(n1628), .B(n1433), .Z(n1434) );
  XNOR U2274 ( .A(n4665), .B(n1434), .Z(out[1161]) );
  XNOR U2275 ( .A(n1436), .B(n1435), .Z(n3960) );
  XNOR U2276 ( .A(in[1014]), .B(n3960), .Z(n4673) );
  NAND U2277 ( .A(n1630), .B(n1437), .Z(n1438) );
  XNOR U2278 ( .A(n4673), .B(n1438), .Z(out[1162]) );
  XNOR U2279 ( .A(n1440), .B(n1439), .Z(n3962) );
  XNOR U2280 ( .A(in[1015]), .B(n3962), .Z(n4677) );
  NAND U2281 ( .A(n1632), .B(n1441), .Z(n1442) );
  XNOR U2282 ( .A(n4677), .B(n1442), .Z(out[1163]) );
  XNOR U2283 ( .A(n1444), .B(n1443), .Z(n3818) );
  XNOR U2284 ( .A(in[1016]), .B(n3818), .Z(n4681) );
  NAND U2285 ( .A(n1634), .B(n1445), .Z(n1446) );
  XNOR U2286 ( .A(n4681), .B(n1446), .Z(out[1164]) );
  XNOR U2287 ( .A(n1448), .B(n1447), .Z(n3820) );
  XNOR U2288 ( .A(in[1017]), .B(n3820), .Z(n4685) );
  NAND U2289 ( .A(n1636), .B(n1449), .Z(n1450) );
  XNOR U2290 ( .A(n4685), .B(n1450), .Z(out[1165]) );
  XNOR U2291 ( .A(n1452), .B(n1451), .Z(n3822) );
  XNOR U2292 ( .A(in[1018]), .B(n3822), .Z(n4689) );
  NAND U2293 ( .A(n1639), .B(n1453), .Z(n1454) );
  XNOR U2294 ( .A(n4689), .B(n1454), .Z(out[1166]) );
  XNOR U2295 ( .A(n1456), .B(n1455), .Z(n3824) );
  XNOR U2296 ( .A(in[1019]), .B(n3824), .Z(n4693) );
  NAND U2297 ( .A(n1641), .B(n1457), .Z(n1458) );
  XNOR U2298 ( .A(n4693), .B(n1458), .Z(out[1167]) );
  XOR U2299 ( .A(n1460), .B(n1459), .Z(n3826) );
  XNOR U2300 ( .A(in[1020]), .B(n3826), .Z(n4697) );
  NAND U2301 ( .A(n1643), .B(n1461), .Z(n1462) );
  XNOR U2302 ( .A(n4697), .B(n1462), .Z(out[1168]) );
  XOR U2303 ( .A(n1464), .B(n1463), .Z(n3828) );
  XNOR U2304 ( .A(in[1021]), .B(n3828), .Z(n4701) );
  NAND U2305 ( .A(n1645), .B(n1465), .Z(n1466) );
  XNOR U2306 ( .A(n4701), .B(n1466), .Z(out[1169]) );
  XOR U2307 ( .A(in[587]), .B(n3660), .Z(n2584) );
  XOR U2308 ( .A(in[242]), .B(n3761), .Z(n3141) );
  XNOR U2309 ( .A(in[1462]), .B(n3804), .Z(n3138) );
  NAND U2310 ( .A(n3141), .B(n3138), .Z(n1467) );
  XNOR U2311 ( .A(n2584), .B(n1467), .Z(out[116]) );
  XOR U2312 ( .A(n1469), .B(n1468), .Z(n3834) );
  XNOR U2313 ( .A(in[1022]), .B(n3834), .Z(n4705) );
  NAND U2314 ( .A(n1647), .B(n1470), .Z(n1471) );
  XNOR U2315 ( .A(n4705), .B(n1471), .Z(out[1170]) );
  XNOR U2316 ( .A(n1473), .B(n1472), .Z(n3836) );
  XNOR U2317 ( .A(in[1023]), .B(n3836), .Z(n4709) );
  NAND U2318 ( .A(n1649), .B(n1474), .Z(n1475) );
  XNOR U2319 ( .A(n4709), .B(n1475), .Z(out[1171]) );
  XOR U2320 ( .A(n1477), .B(n1476), .Z(n3838) );
  XNOR U2321 ( .A(in[960]), .B(n3838), .Z(n4717) );
  NAND U2322 ( .A(n1651), .B(n1478), .Z(n1479) );
  XNOR U2323 ( .A(n4717), .B(n1479), .Z(out[1172]) );
  XOR U2324 ( .A(n1481), .B(n1480), .Z(n3840) );
  XNOR U2325 ( .A(in[961]), .B(n3840), .Z(n4721) );
  NAND U2326 ( .A(n1653), .B(n1482), .Z(n1483) );
  XNOR U2327 ( .A(n4721), .B(n1483), .Z(out[1173]) );
  XOR U2328 ( .A(n1485), .B(n1484), .Z(n3842) );
  XNOR U2329 ( .A(in[962]), .B(n3842), .Z(n4725) );
  NAND U2330 ( .A(n1655), .B(n1486), .Z(n1487) );
  XNOR U2331 ( .A(n4725), .B(n1487), .Z(out[1174]) );
  XOR U2332 ( .A(n1489), .B(n1488), .Z(n3844) );
  XNOR U2333 ( .A(in[963]), .B(n3844), .Z(n4729) );
  NAND U2334 ( .A(n1657), .B(n1490), .Z(n1491) );
  XNOR U2335 ( .A(n4729), .B(n1491), .Z(out[1175]) );
  XOR U2336 ( .A(n1493), .B(n1492), .Z(n3846) );
  XNOR U2337 ( .A(in[964]), .B(n3846), .Z(n4733) );
  NAND U2338 ( .A(n1660), .B(n1494), .Z(n1495) );
  XNOR U2339 ( .A(n4733), .B(n1495), .Z(out[1176]) );
  XOR U2340 ( .A(n1497), .B(n1496), .Z(n3848) );
  XNOR U2341 ( .A(in[965]), .B(n3848), .Z(n4737) );
  NAND U2342 ( .A(n1662), .B(n1498), .Z(n1499) );
  XNOR U2343 ( .A(n4737), .B(n1499), .Z(out[1177]) );
  XOR U2344 ( .A(n1501), .B(n1500), .Z(n3850) );
  XNOR U2345 ( .A(in[966]), .B(n3850), .Z(n4741) );
  NAND U2346 ( .A(n1664), .B(n1502), .Z(n1503) );
  XNOR U2347 ( .A(n4741), .B(n1503), .Z(out[1178]) );
  XOR U2348 ( .A(n1505), .B(n1504), .Z(n3852) );
  XNOR U2349 ( .A(in[967]), .B(n3852), .Z(n4745) );
  NAND U2350 ( .A(n1666), .B(n1506), .Z(n1507) );
  XNOR U2351 ( .A(n4745), .B(n1507), .Z(out[1179]) );
  XOR U2352 ( .A(in[588]), .B(n3668), .Z(n2586) );
  XOR U2353 ( .A(in[243]), .B(n3765), .Z(n3165) );
  XNOR U2354 ( .A(in[1463]), .B(n3808), .Z(n3162) );
  NAND U2355 ( .A(n3165), .B(n3162), .Z(n1508) );
  XNOR U2356 ( .A(n2586), .B(n1508), .Z(out[117]) );
  XOR U2357 ( .A(n1510), .B(n1509), .Z(n3856) );
  XNOR U2358 ( .A(in[968]), .B(n3856), .Z(n4749) );
  NAND U2359 ( .A(n1668), .B(n1511), .Z(n1512) );
  XNOR U2360 ( .A(n4749), .B(n1512), .Z(out[1180]) );
  XOR U2361 ( .A(n1514), .B(n1513), .Z(n3858) );
  XNOR U2362 ( .A(in[969]), .B(n3858), .Z(n4753) );
  NAND U2363 ( .A(n1670), .B(n1515), .Z(n1516) );
  XNOR U2364 ( .A(n4753), .B(n1516), .Z(out[1181]) );
  XNOR U2365 ( .A(n1518), .B(n1517), .Z(n3860) );
  XNOR U2366 ( .A(in[970]), .B(n3860), .Z(n4761) );
  NAND U2367 ( .A(n1672), .B(n1519), .Z(n1520) );
  XNOR U2368 ( .A(n4761), .B(n1520), .Z(out[1182]) );
  XOR U2369 ( .A(n1522), .B(n1521), .Z(n3862) );
  XNOR U2370 ( .A(in[971]), .B(n3862), .Z(n4765) );
  NAND U2371 ( .A(n1674), .B(n1523), .Z(n1524) );
  XNOR U2372 ( .A(n4765), .B(n1524), .Z(out[1183]) );
  XOR U2373 ( .A(n1526), .B(n1525), .Z(n3864) );
  XNOR U2374 ( .A(in[972]), .B(n3864), .Z(n4769) );
  NAND U2375 ( .A(n1676), .B(n1527), .Z(n1528) );
  XNOR U2376 ( .A(n4769), .B(n1528), .Z(out[1184]) );
  XOR U2377 ( .A(n1530), .B(n1529), .Z(n3866) );
  XNOR U2378 ( .A(in[973]), .B(n3866), .Z(n4773) );
  NAND U2379 ( .A(n1678), .B(n1531), .Z(n1532) );
  XNOR U2380 ( .A(n4773), .B(n1532), .Z(out[1185]) );
  XOR U2381 ( .A(n1534), .B(n1533), .Z(n3868) );
  XNOR U2382 ( .A(in[974]), .B(n3868), .Z(n4777) );
  NAND U2383 ( .A(n1681), .B(n1535), .Z(n1536) );
  XNOR U2384 ( .A(n4777), .B(n1536), .Z(out[1186]) );
  XNOR U2385 ( .A(n1538), .B(n1537), .Z(n3870) );
  XNOR U2386 ( .A(in[975]), .B(n3870), .Z(n4781) );
  NAND U2387 ( .A(n1683), .B(n1539), .Z(n1540) );
  XNOR U2388 ( .A(n4781), .B(n1540), .Z(out[1187]) );
  XNOR U2389 ( .A(n1542), .B(n1541), .Z(n3872) );
  XNOR U2390 ( .A(in[976]), .B(n3872), .Z(n4785) );
  NAND U2391 ( .A(n1685), .B(n1543), .Z(n1544) );
  XNOR U2392 ( .A(n4785), .B(n1544), .Z(out[1188]) );
  XOR U2393 ( .A(n1546), .B(n1545), .Z(n3874) );
  XNOR U2394 ( .A(in[977]), .B(n3874), .Z(n4789) );
  NAND U2395 ( .A(n1687), .B(n1547), .Z(n1548) );
  XNOR U2396 ( .A(n4789), .B(n1548), .Z(out[1189]) );
  XOR U2397 ( .A(in[589]), .B(n3672), .Z(n2588) );
  XOR U2398 ( .A(in[244]), .B(n3769), .Z(n3189) );
  XNOR U2399 ( .A(in[1464]), .B(n3812), .Z(n3186) );
  NAND U2400 ( .A(n3189), .B(n3186), .Z(n1549) );
  XNOR U2401 ( .A(n2588), .B(n1549), .Z(out[118]) );
  XOR U2402 ( .A(n1551), .B(n1550), .Z(n3878) );
  XNOR U2403 ( .A(in[978]), .B(n3878), .Z(n4793) );
  NAND U2404 ( .A(n1689), .B(n1552), .Z(n1553) );
  XNOR U2405 ( .A(n4793), .B(n1553), .Z(out[1190]) );
  XNOR U2406 ( .A(n1555), .B(n1554), .Z(n3880) );
  XNOR U2407 ( .A(in[979]), .B(n3880), .Z(n4797) );
  NAND U2408 ( .A(n1691), .B(n1556), .Z(n1557) );
  XNOR U2409 ( .A(n4797), .B(n1557), .Z(out[1191]) );
  OR U2410 ( .A(n1694), .B(n1558), .Z(n1559) );
  XNOR U2411 ( .A(n1693), .B(n1559), .Z(out[1192]) );
  OR U2412 ( .A(n1698), .B(n1560), .Z(n1561) );
  XNOR U2413 ( .A(n1697), .B(n1561), .Z(out[1193]) );
  OR U2414 ( .A(n1702), .B(n1562), .Z(n1563) );
  XNOR U2415 ( .A(n1701), .B(n1563), .Z(out[1194]) );
  OR U2416 ( .A(n1706), .B(n1564), .Z(n1565) );
  XNOR U2417 ( .A(n1705), .B(n1565), .Z(out[1195]) );
  OR U2418 ( .A(n1711), .B(n1566), .Z(n1567) );
  XNOR U2419 ( .A(n1710), .B(n1567), .Z(out[1196]) );
  OR U2420 ( .A(n1715), .B(n1568), .Z(n1569) );
  XNOR U2421 ( .A(n1714), .B(n1569), .Z(out[1197]) );
  OR U2422 ( .A(n1719), .B(n1570), .Z(n1571) );
  XNOR U2423 ( .A(n1718), .B(n1571), .Z(out[1198]) );
  OR U2424 ( .A(n1723), .B(n1572), .Z(n1573) );
  XNOR U2425 ( .A(n1722), .B(n1573), .Z(out[1199]) );
  XOR U2426 ( .A(in[590]), .B(n3676), .Z(n2590) );
  XOR U2427 ( .A(in[245]), .B(n3773), .Z(n3213) );
  XNOR U2428 ( .A(in[1465]), .B(n3816), .Z(n3210) );
  NAND U2429 ( .A(n3213), .B(n3210), .Z(n1574) );
  XNOR U2430 ( .A(n2590), .B(n1574), .Z(out[119]) );
  XOR U2431 ( .A(in[201]), .B(n3581), .Z(n3945) );
  XNOR U2432 ( .A(in[1421]), .B(n3618), .Z(n3944) );
  XOR U2433 ( .A(in[1044]), .B(n4123), .Z(n2635) );
  NAND U2434 ( .A(n3944), .B(n2635), .Z(n1575) );
  XNOR U2435 ( .A(n3945), .B(n1575), .Z(out[11]) );
  OR U2436 ( .A(n1727), .B(n1576), .Z(n1577) );
  XNOR U2437 ( .A(n1726), .B(n1577), .Z(out[1200]) );
  OR U2438 ( .A(n1731), .B(n1578), .Z(n1579) );
  XNOR U2439 ( .A(n1730), .B(n1579), .Z(out[1201]) );
  OR U2440 ( .A(n1735), .B(n1580), .Z(n1581) );
  XNOR U2441 ( .A(n1734), .B(n1581), .Z(out[1202]) );
  OR U2442 ( .A(n1739), .B(n1582), .Z(n1583) );
  XNOR U2443 ( .A(n1738), .B(n1583), .Z(out[1203]) );
  OR U2444 ( .A(n1743), .B(n1584), .Z(n1585) );
  XNOR U2445 ( .A(n1742), .B(n1585), .Z(out[1204]) );
  OR U2446 ( .A(n1747), .B(n1586), .Z(n1587) );
  XNOR U2447 ( .A(n1746), .B(n1587), .Z(out[1205]) );
  OR U2448 ( .A(n1752), .B(n1588), .Z(n1589) );
  XNOR U2449 ( .A(n1751), .B(n1589), .Z(out[1206]) );
  OR U2450 ( .A(n1756), .B(n1590), .Z(n1591) );
  XNOR U2451 ( .A(n1755), .B(n1591), .Z(out[1207]) );
  OR U2452 ( .A(n1760), .B(n1592), .Z(n1593) );
  XNOR U2453 ( .A(n1759), .B(n1593), .Z(out[1208]) );
  OR U2454 ( .A(n1764), .B(n1594), .Z(n1595) );
  XNOR U2455 ( .A(n1763), .B(n1595), .Z(out[1209]) );
  XOR U2456 ( .A(in[591]), .B(n3680), .Z(n2592) );
  XOR U2457 ( .A(in[246]), .B(n3777), .Z(n3237) );
  XNOR U2458 ( .A(in[1466]), .B(n3538), .Z(n3234) );
  NAND U2459 ( .A(n3237), .B(n3234), .Z(n1596) );
  XNOR U2460 ( .A(n2592), .B(n1596), .Z(out[120]) );
  OR U2461 ( .A(n1768), .B(n1597), .Z(n1598) );
  XNOR U2462 ( .A(n1767), .B(n1598), .Z(out[1210]) );
  OR U2463 ( .A(n1772), .B(n1599), .Z(n1600) );
  XNOR U2464 ( .A(n1771), .B(n1600), .Z(out[1211]) );
  OR U2465 ( .A(n1776), .B(n1601), .Z(n1602) );
  XNOR U2466 ( .A(n1775), .B(n1602), .Z(out[1212]) );
  OR U2467 ( .A(n1780), .B(n1603), .Z(n1604) );
  XNOR U2468 ( .A(n1779), .B(n1604), .Z(out[1213]) );
  OR U2469 ( .A(n1784), .B(n1605), .Z(n1606) );
  XNOR U2470 ( .A(n1783), .B(n1606), .Z(out[1214]) );
  OR U2471 ( .A(n1788), .B(n1607), .Z(n1608) );
  XNOR U2472 ( .A(n1787), .B(n1608), .Z(out[1215]) );
  OR U2473 ( .A(n4629), .B(n1609), .Z(n1610) );
  XNOR U2474 ( .A(n4628), .B(n1610), .Z(out[1216]) );
  OR U2475 ( .A(n4633), .B(n1611), .Z(n1612) );
  XNOR U2476 ( .A(n4632), .B(n1612), .Z(out[1217]) );
  OR U2477 ( .A(n4637), .B(n1613), .Z(n1614) );
  XNOR U2478 ( .A(n4636), .B(n1614), .Z(out[1218]) );
  OR U2479 ( .A(n4641), .B(n1615), .Z(n1616) );
  XNOR U2480 ( .A(n4640), .B(n1616), .Z(out[1219]) );
  XOR U2481 ( .A(in[592]), .B(n3684), .Z(n2594) );
  XOR U2482 ( .A(in[247]), .B(n3781), .Z(n3269) );
  XNOR U2483 ( .A(in[1467]), .B(n3542), .Z(n3266) );
  NAND U2484 ( .A(n3269), .B(n3266), .Z(n1617) );
  XNOR U2485 ( .A(n2594), .B(n1617), .Z(out[121]) );
  OR U2486 ( .A(n4645), .B(n1618), .Z(n1619) );
  XNOR U2487 ( .A(n4644), .B(n1619), .Z(out[1220]) );
  OR U2488 ( .A(n4649), .B(n1620), .Z(n1621) );
  XNOR U2489 ( .A(n4648), .B(n1621), .Z(out[1221]) );
  OR U2490 ( .A(n4653), .B(n1622), .Z(n1623) );
  XNOR U2491 ( .A(n4652), .B(n1623), .Z(out[1222]) );
  OR U2492 ( .A(n4657), .B(n1624), .Z(n1625) );
  XNOR U2493 ( .A(n4656), .B(n1625), .Z(out[1223]) );
  OR U2494 ( .A(n4661), .B(n1626), .Z(n1627) );
  XNOR U2495 ( .A(n4660), .B(n1627), .Z(out[1224]) );
  OR U2496 ( .A(n4665), .B(n1628), .Z(n1629) );
  XNOR U2497 ( .A(n4664), .B(n1629), .Z(out[1225]) );
  OR U2498 ( .A(n4673), .B(n1630), .Z(n1631) );
  XNOR U2499 ( .A(n4672), .B(n1631), .Z(out[1226]) );
  OR U2500 ( .A(n4677), .B(n1632), .Z(n1633) );
  XNOR U2501 ( .A(n4676), .B(n1633), .Z(out[1227]) );
  OR U2502 ( .A(n4681), .B(n1634), .Z(n1635) );
  XNOR U2503 ( .A(n4680), .B(n1635), .Z(out[1228]) );
  OR U2504 ( .A(n4685), .B(n1636), .Z(n1637) );
  XNOR U2505 ( .A(n4684), .B(n1637), .Z(out[1229]) );
  XOR U2506 ( .A(in[593]), .B(n3688), .Z(n2597) );
  XOR U2507 ( .A(in[248]), .B(n3785), .Z(n3313) );
  XNOR U2508 ( .A(in[1468]), .B(n3546), .Z(n3310) );
  NAND U2509 ( .A(n3313), .B(n3310), .Z(n1638) );
  XNOR U2510 ( .A(n2597), .B(n1638), .Z(out[122]) );
  OR U2511 ( .A(n4689), .B(n1639), .Z(n1640) );
  XNOR U2512 ( .A(n4688), .B(n1640), .Z(out[1230]) );
  OR U2513 ( .A(n4693), .B(n1641), .Z(n1642) );
  XNOR U2514 ( .A(n4692), .B(n1642), .Z(out[1231]) );
  OR U2515 ( .A(n4697), .B(n1643), .Z(n1644) );
  XNOR U2516 ( .A(n4696), .B(n1644), .Z(out[1232]) );
  OR U2517 ( .A(n4701), .B(n1645), .Z(n1646) );
  XNOR U2518 ( .A(n4700), .B(n1646), .Z(out[1233]) );
  OR U2519 ( .A(n4705), .B(n1647), .Z(n1648) );
  XNOR U2520 ( .A(n4704), .B(n1648), .Z(out[1234]) );
  OR U2521 ( .A(n4709), .B(n1649), .Z(n1650) );
  XNOR U2522 ( .A(n4708), .B(n1650), .Z(out[1235]) );
  OR U2523 ( .A(n4717), .B(n1651), .Z(n1652) );
  XNOR U2524 ( .A(n4716), .B(n1652), .Z(out[1236]) );
  OR U2525 ( .A(n4721), .B(n1653), .Z(n1654) );
  XNOR U2526 ( .A(n4720), .B(n1654), .Z(out[1237]) );
  OR U2527 ( .A(n4725), .B(n1655), .Z(n1656) );
  XNOR U2528 ( .A(n4724), .B(n1656), .Z(out[1238]) );
  OR U2529 ( .A(n4729), .B(n1657), .Z(n1658) );
  XNOR U2530 ( .A(n4728), .B(n1658), .Z(out[1239]) );
  XOR U2531 ( .A(in[594]), .B(n3692), .Z(n2599) );
  XOR U2532 ( .A(in[249]), .B(n3789), .Z(n3357) );
  XNOR U2533 ( .A(in[1469]), .B(n3550), .Z(n3354) );
  NAND U2534 ( .A(n3357), .B(n3354), .Z(n1659) );
  XNOR U2535 ( .A(n2599), .B(n1659), .Z(out[123]) );
  OR U2536 ( .A(n4733), .B(n1660), .Z(n1661) );
  XNOR U2537 ( .A(n4732), .B(n1661), .Z(out[1240]) );
  OR U2538 ( .A(n4737), .B(n1662), .Z(n1663) );
  XNOR U2539 ( .A(n4736), .B(n1663), .Z(out[1241]) );
  OR U2540 ( .A(n4741), .B(n1664), .Z(n1665) );
  XNOR U2541 ( .A(n4740), .B(n1665), .Z(out[1242]) );
  OR U2542 ( .A(n4745), .B(n1666), .Z(n1667) );
  XNOR U2543 ( .A(n4744), .B(n1667), .Z(out[1243]) );
  OR U2544 ( .A(n4749), .B(n1668), .Z(n1669) );
  XNOR U2545 ( .A(n4748), .B(n1669), .Z(out[1244]) );
  OR U2546 ( .A(n4753), .B(n1670), .Z(n1671) );
  XNOR U2547 ( .A(n4752), .B(n1671), .Z(out[1245]) );
  OR U2548 ( .A(n4761), .B(n1672), .Z(n1673) );
  XNOR U2549 ( .A(n4760), .B(n1673), .Z(out[1246]) );
  OR U2550 ( .A(n4765), .B(n1674), .Z(n1675) );
  XNOR U2551 ( .A(n4764), .B(n1675), .Z(out[1247]) );
  OR U2552 ( .A(n4769), .B(n1676), .Z(n1677) );
  XNOR U2553 ( .A(n4768), .B(n1677), .Z(out[1248]) );
  OR U2554 ( .A(n4773), .B(n1678), .Z(n1679) );
  XNOR U2555 ( .A(n4772), .B(n1679), .Z(out[1249]) );
  XOR U2556 ( .A(in[595]), .B(n3696), .Z(n2601) );
  XOR U2557 ( .A(in[250]), .B(n3793), .Z(n3403) );
  XNOR U2558 ( .A(in[1470]), .B(n3554), .Z(n3400) );
  NAND U2559 ( .A(n3403), .B(n3400), .Z(n1680) );
  XNOR U2560 ( .A(n2601), .B(n1680), .Z(out[124]) );
  OR U2561 ( .A(n4777), .B(n1681), .Z(n1682) );
  XNOR U2562 ( .A(n4776), .B(n1682), .Z(out[1250]) );
  OR U2563 ( .A(n4781), .B(n1683), .Z(n1684) );
  XNOR U2564 ( .A(n4780), .B(n1684), .Z(out[1251]) );
  OR U2565 ( .A(n4785), .B(n1685), .Z(n1686) );
  XNOR U2566 ( .A(n4784), .B(n1686), .Z(out[1252]) );
  OR U2567 ( .A(n4789), .B(n1687), .Z(n1688) );
  XNOR U2568 ( .A(n4788), .B(n1688), .Z(out[1253]) );
  OR U2569 ( .A(n4793), .B(n1689), .Z(n1690) );
  XNOR U2570 ( .A(n4792), .B(n1690), .Z(out[1254]) );
  OR U2571 ( .A(n4797), .B(n1691), .Z(n1692) );
  XNOR U2572 ( .A(n4796), .B(n1692), .Z(out[1255]) );
  ANDN U2573 ( .B(n1694), .A(n1693), .Z(n1695) );
  XNOR U2574 ( .A(n1696), .B(n1695), .Z(out[1256]) );
  ANDN U2575 ( .B(n1698), .A(n1697), .Z(n1699) );
  XNOR U2576 ( .A(n1700), .B(n1699), .Z(out[1257]) );
  ANDN U2577 ( .B(n1702), .A(n1701), .Z(n1703) );
  XNOR U2578 ( .A(n1704), .B(n1703), .Z(out[1258]) );
  ANDN U2579 ( .B(n1706), .A(n1705), .Z(n1707) );
  XNOR U2580 ( .A(n1708), .B(n1707), .Z(out[1259]) );
  XOR U2581 ( .A(in[596]), .B(n3700), .Z(n2603) );
  XNOR U2582 ( .A(in[251]), .B(n3803), .Z(n3447) );
  XNOR U2583 ( .A(in[1471]), .B(n3558), .Z(n3444) );
  NAND U2584 ( .A(n3447), .B(n3444), .Z(n1709) );
  XNOR U2585 ( .A(n2603), .B(n1709), .Z(out[125]) );
  ANDN U2586 ( .B(n1711), .A(n1710), .Z(n1712) );
  XNOR U2587 ( .A(n1713), .B(n1712), .Z(out[1260]) );
  ANDN U2588 ( .B(n1715), .A(n1714), .Z(n1716) );
  XNOR U2589 ( .A(n1717), .B(n1716), .Z(out[1261]) );
  ANDN U2590 ( .B(n1719), .A(n1718), .Z(n1720) );
  XNOR U2591 ( .A(n1721), .B(n1720), .Z(out[1262]) );
  ANDN U2592 ( .B(n1723), .A(n1722), .Z(n1724) );
  XNOR U2593 ( .A(n1725), .B(n1724), .Z(out[1263]) );
  ANDN U2594 ( .B(n1727), .A(n1726), .Z(n1728) );
  XNOR U2595 ( .A(n1729), .B(n1728), .Z(out[1264]) );
  ANDN U2596 ( .B(n1731), .A(n1730), .Z(n1732) );
  XNOR U2597 ( .A(n1733), .B(n1732), .Z(out[1265]) );
  ANDN U2598 ( .B(n1735), .A(n1734), .Z(n1736) );
  XNOR U2599 ( .A(n1737), .B(n1736), .Z(out[1266]) );
  ANDN U2600 ( .B(n1739), .A(n1738), .Z(n1740) );
  XNOR U2601 ( .A(n1741), .B(n1740), .Z(out[1267]) );
  ANDN U2602 ( .B(n1743), .A(n1742), .Z(n1744) );
  XNOR U2603 ( .A(n1745), .B(n1744), .Z(out[1268]) );
  ANDN U2604 ( .B(n1747), .A(n1746), .Z(n1748) );
  XNOR U2605 ( .A(n1749), .B(n1748), .Z(out[1269]) );
  XOR U2606 ( .A(in[597]), .B(n3704), .Z(n2605) );
  XNOR U2607 ( .A(in[252]), .B(n3807), .Z(n3491) );
  XNOR U2608 ( .A(in[1408]), .B(n3562), .Z(n3488) );
  NAND U2609 ( .A(n3491), .B(n3488), .Z(n1750) );
  XNOR U2610 ( .A(n2605), .B(n1750), .Z(out[126]) );
  ANDN U2611 ( .B(n1752), .A(n1751), .Z(n1753) );
  XNOR U2612 ( .A(n1754), .B(n1753), .Z(out[1270]) );
  ANDN U2613 ( .B(n1756), .A(n1755), .Z(n1757) );
  XNOR U2614 ( .A(n1758), .B(n1757), .Z(out[1271]) );
  ANDN U2615 ( .B(n1760), .A(n1759), .Z(n1761) );
  XNOR U2616 ( .A(n1762), .B(n1761), .Z(out[1272]) );
  ANDN U2617 ( .B(n1764), .A(n1763), .Z(n1765) );
  XNOR U2618 ( .A(n1766), .B(n1765), .Z(out[1273]) );
  ANDN U2619 ( .B(n1768), .A(n1767), .Z(n1769) );
  XNOR U2620 ( .A(n1770), .B(n1769), .Z(out[1274]) );
  ANDN U2621 ( .B(n1772), .A(n1771), .Z(n1773) );
  XNOR U2622 ( .A(n1774), .B(n1773), .Z(out[1275]) );
  ANDN U2623 ( .B(n1776), .A(n1775), .Z(n1777) );
  XNOR U2624 ( .A(n1778), .B(n1777), .Z(out[1276]) );
  ANDN U2625 ( .B(n1780), .A(n1779), .Z(n1781) );
  XNOR U2626 ( .A(n1782), .B(n1781), .Z(out[1277]) );
  ANDN U2627 ( .B(n1784), .A(n1783), .Z(n1785) );
  XNOR U2628 ( .A(n1786), .B(n1785), .Z(out[1278]) );
  ANDN U2629 ( .B(n1788), .A(n1787), .Z(n1789) );
  XNOR U2630 ( .A(n1790), .B(n1789), .Z(out[1279]) );
  XOR U2631 ( .A(in[598]), .B(n3712), .Z(n2607) );
  XNOR U2632 ( .A(in[253]), .B(n3811), .Z(n3535) );
  XNOR U2633 ( .A(in[1409]), .B(n3566), .Z(n3532) );
  NAND U2634 ( .A(n3535), .B(n3532), .Z(n1791) );
  XNOR U2635 ( .A(n2607), .B(n1791), .Z(out[127]) );
  XNOR U2636 ( .A(in[50]), .B(n3952), .Z(n1934) );
  XOR U2637 ( .A(in[1536]), .B(n3612), .Z(n2206) );
  XNOR U2638 ( .A(in[1172]), .B(n3629), .Z(n2204) );
  NAND U2639 ( .A(n2206), .B(n2204), .Z(n1792) );
  XNOR U2640 ( .A(n1934), .B(n1792), .Z(out[1280]) );
  XNOR U2641 ( .A(in[51]), .B(n3954), .Z(n1936) );
  XOR U2642 ( .A(in[1537]), .B(n3616), .Z(n2211) );
  XNOR U2643 ( .A(in[1173]), .B(n3633), .Z(n2209) );
  NAND U2644 ( .A(n2211), .B(n2209), .Z(n1793) );
  XNOR U2645 ( .A(n1936), .B(n1793), .Z(out[1281]) );
  XNOR U2646 ( .A(in[52]), .B(n3956), .Z(n1939) );
  XOR U2647 ( .A(in[1538]), .B(n3624), .Z(n2217) );
  XNOR U2648 ( .A(in[1174]), .B(n3637), .Z(n2214) );
  NAND U2649 ( .A(n2217), .B(n2214), .Z(n1794) );
  XNOR U2650 ( .A(n1939), .B(n1794), .Z(out[1282]) );
  XNOR U2651 ( .A(in[53]), .B(n3958), .Z(n1941) );
  XOR U2652 ( .A(in[1539]), .B(n3628), .Z(n2220) );
  XNOR U2653 ( .A(in[1175]), .B(n3641), .Z(n2218) );
  NAND U2654 ( .A(n2220), .B(n2218), .Z(n1795) );
  XNOR U2655 ( .A(n1941), .B(n1795), .Z(out[1283]) );
  XNOR U2656 ( .A(in[54]), .B(n3960), .Z(n1943) );
  XNOR U2657 ( .A(in[1540]), .B(n3632), .Z(n2227) );
  XNOR U2658 ( .A(in[1176]), .B(n3645), .Z(n2224) );
  NAND U2659 ( .A(n2227), .B(n2224), .Z(n1796) );
  XNOR U2660 ( .A(n1943), .B(n1796), .Z(out[1284]) );
  XNOR U2661 ( .A(in[55]), .B(n3962), .Z(n1945) );
  XNOR U2662 ( .A(in[1541]), .B(n3636), .Z(n2231) );
  XNOR U2663 ( .A(in[1177]), .B(n3649), .Z(n2228) );
  NAND U2664 ( .A(n2231), .B(n2228), .Z(n1797) );
  XNOR U2665 ( .A(n1945), .B(n1797), .Z(out[1285]) );
  XNOR U2666 ( .A(in[56]), .B(n3818), .Z(n1947) );
  XNOR U2667 ( .A(in[1542]), .B(n3640), .Z(n2235) );
  XNOR U2668 ( .A(in[1178]), .B(n3653), .Z(n2232) );
  NAND U2669 ( .A(n2235), .B(n2232), .Z(n1798) );
  XNOR U2670 ( .A(n1947), .B(n1798), .Z(out[1286]) );
  XNOR U2671 ( .A(in[57]), .B(n3820), .Z(n1949) );
  XNOR U2672 ( .A(in[1543]), .B(n3644), .Z(n2238) );
  XNOR U2673 ( .A(in[1179]), .B(n3657), .Z(n2236) );
  NAND U2674 ( .A(n2238), .B(n2236), .Z(n1799) );
  XNOR U2675 ( .A(n1949), .B(n1799), .Z(out[1287]) );
  XNOR U2676 ( .A(in[58]), .B(n3822), .Z(n1951) );
  XNOR U2677 ( .A(in[1544]), .B(n3648), .Z(n2244) );
  XNOR U2678 ( .A(in[1180]), .B(n3661), .Z(n2241) );
  NAND U2679 ( .A(n2244), .B(n2241), .Z(n1800) );
  XNOR U2680 ( .A(n1951), .B(n1800), .Z(out[1288]) );
  XNOR U2681 ( .A(in[59]), .B(n3824), .Z(n1953) );
  XNOR U2682 ( .A(in[1545]), .B(n3652), .Z(n2248) );
  XNOR U2683 ( .A(in[1181]), .B(n3669), .Z(n2245) );
  NAND U2684 ( .A(n2248), .B(n2245), .Z(n1801) );
  XNOR U2685 ( .A(n1953), .B(n1801), .Z(out[1289]) );
  XNOR U2686 ( .A(in[665]), .B(n3892), .Z(n2610) );
  XNOR U2687 ( .A(in[599]), .B(n3716), .Z(n3579) );
  NAND U2688 ( .A(n3579), .B(n3577), .Z(n1802) );
  XNOR U2689 ( .A(n2610), .B(n1802), .Z(out[128]) );
  XNOR U2690 ( .A(in[60]), .B(n3826), .Z(n1955) );
  XNOR U2691 ( .A(in[1546]), .B(n3656), .Z(n2252) );
  XNOR U2692 ( .A(in[1182]), .B(n3673), .Z(n2249) );
  NAND U2693 ( .A(n2252), .B(n2249), .Z(n1803) );
  XNOR U2694 ( .A(n1955), .B(n1803), .Z(out[1290]) );
  XNOR U2695 ( .A(in[61]), .B(n3828), .Z(n1957) );
  XNOR U2696 ( .A(in[1547]), .B(n3660), .Z(n2256) );
  XNOR U2697 ( .A(in[1183]), .B(n3677), .Z(n2253) );
  NAND U2698 ( .A(n2256), .B(n2253), .Z(n1804) );
  XNOR U2699 ( .A(n1957), .B(n1804), .Z(out[1291]) );
  XNOR U2700 ( .A(in[62]), .B(n3834), .Z(n1960) );
  XNOR U2701 ( .A(in[1548]), .B(n3668), .Z(n2260) );
  XNOR U2702 ( .A(in[1184]), .B(n3681), .Z(n2257) );
  NAND U2703 ( .A(n2260), .B(n2257), .Z(n1805) );
  XNOR U2704 ( .A(n1960), .B(n1805), .Z(out[1292]) );
  XNOR U2705 ( .A(in[63]), .B(n3836), .Z(n1962) );
  XNOR U2706 ( .A(in[1549]), .B(n3672), .Z(n2264) );
  XNOR U2707 ( .A(in[1185]), .B(n3685), .Z(n2261) );
  NAND U2708 ( .A(n2264), .B(n2261), .Z(n1806) );
  XNOR U2709 ( .A(n1962), .B(n1806), .Z(out[1293]) );
  XNOR U2710 ( .A(in[0]), .B(n3838), .Z(n1964) );
  XNOR U2711 ( .A(in[1550]), .B(n3676), .Z(n2269) );
  XOR U2712 ( .A(n3689), .B(in[1186]), .Z(n2266) );
  NAND U2713 ( .A(n2269), .B(n2266), .Z(n1807) );
  XNOR U2714 ( .A(n1964), .B(n1807), .Z(out[1294]) );
  XNOR U2715 ( .A(in[1]), .B(n3840), .Z(n1966) );
  XNOR U2716 ( .A(in[1551]), .B(n3680), .Z(n2272) );
  XOR U2717 ( .A(n3693), .B(in[1187]), .Z(n2270) );
  NAND U2718 ( .A(n2272), .B(n2270), .Z(n1808) );
  XNOR U2719 ( .A(n1966), .B(n1808), .Z(out[1295]) );
  XNOR U2720 ( .A(in[2]), .B(n3842), .Z(n1968) );
  XNOR U2721 ( .A(in[1552]), .B(n3684), .Z(n2278) );
  XOR U2722 ( .A(n3697), .B(in[1188]), .Z(n2275) );
  NAND U2723 ( .A(n2278), .B(n2275), .Z(n1809) );
  XNOR U2724 ( .A(n1968), .B(n1809), .Z(out[1296]) );
  XNOR U2725 ( .A(in[3]), .B(n3844), .Z(n1970) );
  XNOR U2726 ( .A(in[1553]), .B(n3688), .Z(n2282) );
  XOR U2727 ( .A(n3701), .B(in[1189]), .Z(n2279) );
  NAND U2728 ( .A(n2282), .B(n2279), .Z(n1810) );
  XNOR U2729 ( .A(n1970), .B(n1810), .Z(out[1297]) );
  XNOR U2730 ( .A(in[4]), .B(n3846), .Z(n1972) );
  XNOR U2731 ( .A(in[1554]), .B(n3692), .Z(n2286) );
  XNOR U2732 ( .A(in[1190]), .B(n3705), .Z(n2283) );
  NAND U2733 ( .A(n2286), .B(n2283), .Z(n1811) );
  XNOR U2734 ( .A(n1972), .B(n1811), .Z(out[1298]) );
  XNOR U2735 ( .A(in[5]), .B(n3848), .Z(n1974) );
  XNOR U2736 ( .A(in[1555]), .B(n3696), .Z(n2290) );
  XNOR U2737 ( .A(in[1191]), .B(n3713), .Z(n2287) );
  NAND U2738 ( .A(n2290), .B(n2287), .Z(n1812) );
  XNOR U2739 ( .A(n1974), .B(n1812), .Z(out[1299]) );
  XNOR U2740 ( .A(in[666]), .B(n3894), .Z(n2612) );
  XNOR U2741 ( .A(in[600]), .B(n3720), .Z(n3623) );
  XOR U2742 ( .A(in[255]), .B(n3537), .Z(n3621) );
  NAND U2743 ( .A(n3623), .B(n3621), .Z(n1813) );
  XNOR U2744 ( .A(n2612), .B(n1813), .Z(out[129]) );
  XOR U2745 ( .A(in[202]), .B(n3585), .Z(n3971) );
  XNOR U2746 ( .A(in[1422]), .B(n3626), .Z(n3970) );
  XOR U2747 ( .A(in[1045]), .B(n4126), .Z(n2638) );
  NAND U2748 ( .A(n3970), .B(n2638), .Z(n1814) );
  XNOR U2749 ( .A(n3971), .B(n1814), .Z(out[12]) );
  XNOR U2750 ( .A(in[6]), .B(n3850), .Z(n1976) );
  XNOR U2751 ( .A(in[1556]), .B(n3700), .Z(n2294) );
  XNOR U2752 ( .A(in[1192]), .B(n3717), .Z(n2291) );
  NAND U2753 ( .A(n2294), .B(n2291), .Z(n1815) );
  XNOR U2754 ( .A(n1976), .B(n1815), .Z(out[1300]) );
  XNOR U2755 ( .A(in[7]), .B(n3852), .Z(n1978) );
  XNOR U2756 ( .A(in[1557]), .B(n3704), .Z(n2298) );
  XNOR U2757 ( .A(in[1193]), .B(n3721), .Z(n2295) );
  NAND U2758 ( .A(n2298), .B(n2295), .Z(n1816) );
  XNOR U2759 ( .A(n1978), .B(n1816), .Z(out[1301]) );
  XNOR U2760 ( .A(in[8]), .B(n3856), .Z(n1981) );
  XNOR U2761 ( .A(in[1558]), .B(n3712), .Z(n2302) );
  XNOR U2762 ( .A(in[1194]), .B(n3725), .Z(n2299) );
  NAND U2763 ( .A(n2302), .B(n2299), .Z(n1817) );
  XNOR U2764 ( .A(n1981), .B(n1817), .Z(out[1302]) );
  XNOR U2765 ( .A(in[9]), .B(n3858), .Z(n1983) );
  XNOR U2766 ( .A(in[1559]), .B(n3716), .Z(n2306) );
  XNOR U2767 ( .A(in[1195]), .B(n3729), .Z(n2303) );
  NAND U2768 ( .A(n2306), .B(n2303), .Z(n1818) );
  XNOR U2769 ( .A(n1983), .B(n1818), .Z(out[1303]) );
  XNOR U2770 ( .A(in[10]), .B(n3860), .Z(n1985) );
  XNOR U2771 ( .A(in[1560]), .B(n3720), .Z(n2311) );
  XNOR U2772 ( .A(in[1196]), .B(n3733), .Z(n2308) );
  NAND U2773 ( .A(n2311), .B(n2308), .Z(n1819) );
  XNOR U2774 ( .A(n1985), .B(n1819), .Z(out[1304]) );
  XNOR U2775 ( .A(in[11]), .B(n3862), .Z(n1987) );
  XNOR U2776 ( .A(in[1561]), .B(n3724), .Z(n2315) );
  XNOR U2777 ( .A(in[1197]), .B(n3737), .Z(n2312) );
  NAND U2778 ( .A(n2315), .B(n2312), .Z(n1820) );
  XNOR U2779 ( .A(n1987), .B(n1820), .Z(out[1305]) );
  XNOR U2780 ( .A(in[12]), .B(n3864), .Z(n1989) );
  XNOR U2781 ( .A(in[1562]), .B(n3728), .Z(n2319) );
  XNOR U2782 ( .A(in[1198]), .B(n3741), .Z(n2316) );
  NAND U2783 ( .A(n2319), .B(n2316), .Z(n1821) );
  XNOR U2784 ( .A(n1989), .B(n1821), .Z(out[1306]) );
  XNOR U2785 ( .A(in[13]), .B(n3866), .Z(n1991) );
  XNOR U2786 ( .A(in[1563]), .B(n3732), .Z(n2323) );
  XNOR U2787 ( .A(in[1199]), .B(n3745), .Z(n2320) );
  NAND U2788 ( .A(n2323), .B(n2320), .Z(n1822) );
  XNOR U2789 ( .A(n1991), .B(n1822), .Z(out[1307]) );
  XNOR U2790 ( .A(in[14]), .B(n3868), .Z(n1993) );
  XNOR U2791 ( .A(in[1564]), .B(n3736), .Z(n2327) );
  XNOR U2792 ( .A(in[1200]), .B(n3749), .Z(n2324) );
  NAND U2793 ( .A(n2327), .B(n2324), .Z(n1823) );
  XNOR U2794 ( .A(n1993), .B(n1823), .Z(out[1308]) );
  XNOR U2795 ( .A(in[15]), .B(n3870), .Z(n1995) );
  XNOR U2796 ( .A(in[1565]), .B(n3740), .Z(n2331) );
  XNOR U2797 ( .A(in[1201]), .B(n3757), .Z(n2328) );
  NAND U2798 ( .A(n2331), .B(n2328), .Z(n1824) );
  XNOR U2799 ( .A(n1995), .B(n1824), .Z(out[1309]) );
  XNOR U2800 ( .A(in[667]), .B(n3896), .Z(n2615) );
  XNOR U2801 ( .A(in[601]), .B(n3724), .Z(n3667) );
  XOR U2802 ( .A(in[192]), .B(n3541), .Z(n3664) );
  NAND U2803 ( .A(n3667), .B(n3664), .Z(n1825) );
  XNOR U2804 ( .A(n2615), .B(n1825), .Z(out[130]) );
  XNOR U2805 ( .A(in[16]), .B(n3872), .Z(n1997) );
  XNOR U2806 ( .A(in[1566]), .B(n3744), .Z(n2335) );
  XNOR U2807 ( .A(in[1202]), .B(n3761), .Z(n2332) );
  NAND U2808 ( .A(n2335), .B(n2332), .Z(n1826) );
  XNOR U2809 ( .A(n1997), .B(n1826), .Z(out[1310]) );
  XNOR U2810 ( .A(in[17]), .B(n3874), .Z(n1999) );
  XNOR U2811 ( .A(in[1567]), .B(n3748), .Z(n2338) );
  XNOR U2812 ( .A(in[1203]), .B(n3765), .Z(n2336) );
  NAND U2813 ( .A(n2338), .B(n2336), .Z(n1827) );
  XNOR U2814 ( .A(n1999), .B(n1827), .Z(out[1311]) );
  XNOR U2815 ( .A(in[18]), .B(n3878), .Z(n2002) );
  XNOR U2816 ( .A(in[1568]), .B(n3756), .Z(n2344) );
  XNOR U2817 ( .A(in[1204]), .B(n3769), .Z(n2341) );
  NAND U2818 ( .A(n2344), .B(n2341), .Z(n1828) );
  XNOR U2819 ( .A(n2002), .B(n1828), .Z(out[1312]) );
  XNOR U2820 ( .A(in[19]), .B(n3880), .Z(n2004) );
  XNOR U2821 ( .A(in[1569]), .B(n3760), .Z(n2348) );
  XNOR U2822 ( .A(in[1205]), .B(n3773), .Z(n2345) );
  NAND U2823 ( .A(n2348), .B(n2345), .Z(n1829) );
  XNOR U2824 ( .A(n2004), .B(n1829), .Z(out[1313]) );
  XNOR U2825 ( .A(in[20]), .B(n3882), .Z(n2006) );
  XNOR U2826 ( .A(in[1570]), .B(n3764), .Z(n2353) );
  XNOR U2827 ( .A(in[1206]), .B(n3777), .Z(n2350) );
  NAND U2828 ( .A(n2353), .B(n2350), .Z(n1830) );
  XNOR U2829 ( .A(n2006), .B(n1830), .Z(out[1314]) );
  XNOR U2830 ( .A(in[21]), .B(n3884), .Z(n2008) );
  XNOR U2831 ( .A(in[1571]), .B(n3768), .Z(n2357) );
  XNOR U2832 ( .A(in[1207]), .B(n3781), .Z(n2354) );
  NAND U2833 ( .A(n2357), .B(n2354), .Z(n1831) );
  XNOR U2834 ( .A(n2008), .B(n1831), .Z(out[1315]) );
  XNOR U2835 ( .A(in[22]), .B(n3886), .Z(n2010) );
  XNOR U2836 ( .A(in[1572]), .B(n3772), .Z(n2361) );
  XNOR U2837 ( .A(in[1208]), .B(n3785), .Z(n2358) );
  NAND U2838 ( .A(n2361), .B(n2358), .Z(n1832) );
  XNOR U2839 ( .A(n2010), .B(n1832), .Z(out[1316]) );
  XNOR U2840 ( .A(in[23]), .B(n3888), .Z(n2012) );
  XOR U2841 ( .A(in[1573]), .B(n3776), .Z(n2365) );
  XNOR U2842 ( .A(in[1209]), .B(n3789), .Z(n2362) );
  NAND U2843 ( .A(n2365), .B(n2362), .Z(n1833) );
  XNOR U2844 ( .A(n2012), .B(n1833), .Z(out[1317]) );
  XNOR U2845 ( .A(in[24]), .B(n3890), .Z(n2014) );
  XOR U2846 ( .A(in[1574]), .B(n3780), .Z(n2369) );
  XNOR U2847 ( .A(in[1210]), .B(n3793), .Z(n2366) );
  NAND U2848 ( .A(n2369), .B(n2366), .Z(n1834) );
  XNOR U2849 ( .A(n2014), .B(n1834), .Z(out[1318]) );
  XNOR U2850 ( .A(in[25]), .B(n3892), .Z(n2016) );
  XOR U2851 ( .A(in[1575]), .B(n3784), .Z(n2373) );
  XOR U2852 ( .A(in[1211]), .B(n3803), .Z(n2370) );
  NAND U2853 ( .A(n2373), .B(n2370), .Z(n1835) );
  XNOR U2854 ( .A(n2016), .B(n1835), .Z(out[1319]) );
  XNOR U2855 ( .A(in[668]), .B(n3900), .Z(n2617) );
  XNOR U2856 ( .A(in[602]), .B(n3728), .Z(n3711) );
  XOR U2857 ( .A(in[193]), .B(n3545), .Z(n3708) );
  NAND U2858 ( .A(n3711), .B(n3708), .Z(n1836) );
  XNOR U2859 ( .A(n2617), .B(n1836), .Z(out[131]) );
  XNOR U2860 ( .A(in[26]), .B(n3894), .Z(n2018) );
  XOR U2861 ( .A(in[1576]), .B(n3788), .Z(n2377) );
  XOR U2862 ( .A(in[1212]), .B(n3807), .Z(n2374) );
  NAND U2863 ( .A(n2377), .B(n2374), .Z(n1837) );
  XNOR U2864 ( .A(n2018), .B(n1837), .Z(out[1320]) );
  XNOR U2865 ( .A(in[27]), .B(n3896), .Z(n2020) );
  XOR U2866 ( .A(in[1577]), .B(n3792), .Z(n2381) );
  XOR U2867 ( .A(in[1213]), .B(n3811), .Z(n2378) );
  NAND U2868 ( .A(n2381), .B(n2378), .Z(n1838) );
  XNOR U2869 ( .A(n2020), .B(n1838), .Z(out[1321]) );
  XNOR U2870 ( .A(in[28]), .B(n3900), .Z(n2023) );
  XOR U2871 ( .A(in[1578]), .B(n3802), .Z(n2385) );
  XNOR U2872 ( .A(in[1214]), .B(n3815), .Z(n2382) );
  NAND U2873 ( .A(n2385), .B(n2382), .Z(n1839) );
  XNOR U2874 ( .A(n2023), .B(n1839), .Z(out[1322]) );
  XNOR U2875 ( .A(in[29]), .B(n3902), .Z(n2025) );
  XOR U2876 ( .A(in[1579]), .B(n3806), .Z(n2389) );
  XOR U2877 ( .A(in[1215]), .B(n3537), .Z(n2386) );
  NAND U2878 ( .A(n2389), .B(n2386), .Z(n1840) );
  XNOR U2879 ( .A(n2025), .B(n1840), .Z(out[1323]) );
  XNOR U2880 ( .A(in[30]), .B(n3904), .Z(n2027) );
  XOR U2881 ( .A(in[1580]), .B(n3810), .Z(n2394) );
  XOR U2882 ( .A(in[1152]), .B(n3541), .Z(n2391) );
  NAND U2883 ( .A(n2394), .B(n2391), .Z(n1841) );
  XNOR U2884 ( .A(n2027), .B(n1841), .Z(out[1324]) );
  XNOR U2885 ( .A(in[31]), .B(n3906), .Z(n2029) );
  XOR U2886 ( .A(in[1581]), .B(n3814), .Z(n2398) );
  XOR U2887 ( .A(in[1153]), .B(n3545), .Z(n2395) );
  NAND U2888 ( .A(n2398), .B(n2395), .Z(n1842) );
  XNOR U2889 ( .A(n2029), .B(n1842), .Z(out[1325]) );
  XNOR U2890 ( .A(in[32]), .B(n3908), .Z(n2031) );
  XOR U2891 ( .A(in[1582]), .B(n3536), .Z(n2402) );
  XOR U2892 ( .A(in[1154]), .B(n3549), .Z(n2399) );
  NAND U2893 ( .A(n2402), .B(n2399), .Z(n1843) );
  XNOR U2894 ( .A(n2031), .B(n1843), .Z(out[1326]) );
  XNOR U2895 ( .A(in[33]), .B(n3910), .Z(n2033) );
  XOR U2896 ( .A(in[1583]), .B(n3540), .Z(n2406) );
  XOR U2897 ( .A(in[1155]), .B(n3553), .Z(n2403) );
  NAND U2898 ( .A(n2406), .B(n2403), .Z(n1844) );
  XNOR U2899 ( .A(n2033), .B(n1844), .Z(out[1327]) );
  XNOR U2900 ( .A(in[34]), .B(n3912), .Z(n2035) );
  XOR U2901 ( .A(in[1584]), .B(n3544), .Z(n2410) );
  XOR U2902 ( .A(in[1156]), .B(n3557), .Z(n2407) );
  NAND U2903 ( .A(n2410), .B(n2407), .Z(n1845) );
  XNOR U2904 ( .A(n2035), .B(n1845), .Z(out[1328]) );
  XNOR U2905 ( .A(in[35]), .B(n3914), .Z(n2037) );
  XOR U2906 ( .A(in[1585]), .B(n3548), .Z(n2414) );
  XOR U2907 ( .A(in[1157]), .B(n3561), .Z(n2411) );
  NAND U2908 ( .A(n2414), .B(n2411), .Z(n1846) );
  XNOR U2909 ( .A(n2037), .B(n1846), .Z(out[1329]) );
  XNOR U2910 ( .A(in[669]), .B(n3902), .Z(n2620) );
  XNOR U2911 ( .A(in[603]), .B(n3732), .Z(n3755) );
  XOR U2912 ( .A(in[194]), .B(n3549), .Z(n3752) );
  NAND U2913 ( .A(n3755), .B(n3752), .Z(n1847) );
  XNOR U2914 ( .A(n2620), .B(n1847), .Z(out[132]) );
  XNOR U2915 ( .A(in[36]), .B(n3916), .Z(n2039) );
  XOR U2916 ( .A(in[1586]), .B(n3552), .Z(n2418) );
  XOR U2917 ( .A(in[1158]), .B(n3565), .Z(n2415) );
  NAND U2918 ( .A(n2418), .B(n2415), .Z(n1848) );
  XNOR U2919 ( .A(n2039), .B(n1848), .Z(out[1330]) );
  XNOR U2920 ( .A(in[37]), .B(n3918), .Z(n2041) );
  XOR U2921 ( .A(in[1587]), .B(n3556), .Z(n2422) );
  XOR U2922 ( .A(in[1159]), .B(n3569), .Z(n2419) );
  NAND U2923 ( .A(n2422), .B(n2419), .Z(n1849) );
  XNOR U2924 ( .A(n2041), .B(n1849), .Z(out[1331]) );
  XNOR U2925 ( .A(in[38]), .B(n3924), .Z(n2044) );
  XOR U2926 ( .A(in[1588]), .B(n3560), .Z(n2426) );
  XOR U2927 ( .A(in[1160]), .B(n3573), .Z(n2423) );
  NAND U2928 ( .A(n2426), .B(n2423), .Z(n1850) );
  XNOR U2929 ( .A(n2044), .B(n1850), .Z(out[1332]) );
  XNOR U2930 ( .A(in[39]), .B(n3926), .Z(n2046) );
  XOR U2931 ( .A(in[1589]), .B(n3564), .Z(n2430) );
  XOR U2932 ( .A(in[1161]), .B(n3581), .Z(n2427) );
  NAND U2933 ( .A(n2430), .B(n2427), .Z(n1851) );
  XNOR U2934 ( .A(n2046), .B(n1851), .Z(out[1333]) );
  XNOR U2935 ( .A(in[40]), .B(n3928), .Z(n2048) );
  XOR U2936 ( .A(in[1590]), .B(n3568), .Z(n2435) );
  XOR U2937 ( .A(in[1162]), .B(n3585), .Z(n2432) );
  NAND U2938 ( .A(n2435), .B(n2432), .Z(n1852) );
  XNOR U2939 ( .A(n2048), .B(n1852), .Z(out[1334]) );
  XNOR U2940 ( .A(in[41]), .B(n3930), .Z(n2050) );
  XOR U2941 ( .A(in[1591]), .B(n3572), .Z(n2439) );
  XOR U2942 ( .A(in[1163]), .B(n3589), .Z(n2436) );
  NAND U2943 ( .A(n2439), .B(n2436), .Z(n1853) );
  XNOR U2944 ( .A(n2050), .B(n1853), .Z(out[1335]) );
  XNOR U2945 ( .A(in[42]), .B(n3932), .Z(n2052) );
  XOR U2946 ( .A(in[1592]), .B(n3580), .Z(n2443) );
  XOR U2947 ( .A(in[1164]), .B(n3593), .Z(n2440) );
  NAND U2948 ( .A(n2443), .B(n2440), .Z(n1854) );
  XNOR U2949 ( .A(n2052), .B(n1854), .Z(out[1336]) );
  XNOR U2950 ( .A(in[43]), .B(n3934), .Z(n2054) );
  XOR U2951 ( .A(in[1593]), .B(n3584), .Z(n2447) );
  XOR U2952 ( .A(in[1165]), .B(n3597), .Z(n2444) );
  NAND U2953 ( .A(n2447), .B(n2444), .Z(n1855) );
  XNOR U2954 ( .A(n2054), .B(n1855), .Z(out[1337]) );
  XNOR U2955 ( .A(in[44]), .B(n3936), .Z(n2056) );
  XOR U2956 ( .A(in[1594]), .B(n3588), .Z(n2451) );
  XOR U2957 ( .A(in[1166]), .B(n3601), .Z(n2448) );
  NAND U2958 ( .A(n2451), .B(n2448), .Z(n1856) );
  XNOR U2959 ( .A(n2056), .B(n1856), .Z(out[1338]) );
  XNOR U2960 ( .A(in[45]), .B(n3938), .Z(n2058) );
  XOR U2961 ( .A(in[1595]), .B(n3592), .Z(n2455) );
  XOR U2962 ( .A(in[1167]), .B(n3605), .Z(n2452) );
  NAND U2963 ( .A(n2455), .B(n2452), .Z(n1857) );
  XNOR U2964 ( .A(n2058), .B(n1857), .Z(out[1339]) );
  XNOR U2965 ( .A(in[670]), .B(n3904), .Z(n2622) );
  XNOR U2966 ( .A(in[604]), .B(n3736), .Z(n3799) );
  XOR U2967 ( .A(in[195]), .B(n3553), .Z(n3796) );
  NAND U2968 ( .A(n3799), .B(n3796), .Z(n1858) );
  XNOR U2969 ( .A(n2622), .B(n1858), .Z(out[133]) );
  XNOR U2970 ( .A(in[46]), .B(n3940), .Z(n2060) );
  XOR U2971 ( .A(in[1596]), .B(n3596), .Z(n2459) );
  XOR U2972 ( .A(in[1168]), .B(n3609), .Z(n2456) );
  NAND U2973 ( .A(n2459), .B(n2456), .Z(n1859) );
  XNOR U2974 ( .A(n2060), .B(n1859), .Z(out[1340]) );
  XNOR U2975 ( .A(in[47]), .B(n3942), .Z(n2062) );
  XOR U2976 ( .A(in[1597]), .B(n3600), .Z(n2463) );
  XOR U2977 ( .A(in[1169]), .B(n3613), .Z(n2460) );
  NAND U2978 ( .A(n2463), .B(n2460), .Z(n1860) );
  XNOR U2979 ( .A(n2062), .B(n1860), .Z(out[1341]) );
  XNOR U2980 ( .A(in[48]), .B(n3948), .Z(n2065) );
  XOR U2981 ( .A(in[1598]), .B(n3604), .Z(n2467) );
  XOR U2982 ( .A(in[1170]), .B(n3617), .Z(n2464) );
  NAND U2983 ( .A(n2467), .B(n2464), .Z(n1861) );
  XNOR U2984 ( .A(n2065), .B(n1861), .Z(out[1342]) );
  XNOR U2985 ( .A(in[49]), .B(n3950), .Z(n2067) );
  XOR U2986 ( .A(in[1599]), .B(n3608), .Z(n2470) );
  XNOR U2987 ( .A(in[1171]), .B(n3625), .Z(n2468) );
  NAND U2988 ( .A(n2470), .B(n2468), .Z(n1862) );
  XNOR U2989 ( .A(n2067), .B(n1862), .Z(out[1343]) );
  XOR U2990 ( .A(in[427]), .B(n3980), .Z(n2069) );
  NOR U2991 ( .A(n1934), .B(n2206), .Z(n1863) );
  XNOR U2992 ( .A(n2069), .B(n1863), .Z(out[1344]) );
  XOR U2993 ( .A(in[428]), .B(n3983), .Z(n2071) );
  NOR U2994 ( .A(n1936), .B(n2211), .Z(n1864) );
  XNOR U2995 ( .A(n2071), .B(n1864), .Z(out[1345]) );
  XOR U2996 ( .A(in[429]), .B(n3986), .Z(n2073) );
  NOR U2997 ( .A(n1939), .B(n2217), .Z(n1865) );
  XNOR U2998 ( .A(n2073), .B(n1865), .Z(out[1346]) );
  XOR U2999 ( .A(in[430]), .B(n3989), .Z(n2075) );
  NOR U3000 ( .A(n1941), .B(n2220), .Z(n1866) );
  XNOR U3001 ( .A(n2075), .B(n1866), .Z(out[1347]) );
  XOR U3002 ( .A(in[431]), .B(n3992), .Z(n2077) );
  NOR U3003 ( .A(n1943), .B(n2227), .Z(n1867) );
  XNOR U3004 ( .A(n2077), .B(n1867), .Z(out[1348]) );
  XOR U3005 ( .A(in[432]), .B(n3995), .Z(n2079) );
  NOR U3006 ( .A(n1945), .B(n2231), .Z(n1868) );
  XNOR U3007 ( .A(n2079), .B(n1868), .Z(out[1349]) );
  XNOR U3008 ( .A(in[671]), .B(n3906), .Z(n2624) );
  XNOR U3009 ( .A(in[605]), .B(n3740), .Z(n3833) );
  XOR U3010 ( .A(in[196]), .B(n3557), .Z(n3830) );
  NAND U3011 ( .A(n3833), .B(n3830), .Z(n1869) );
  XNOR U3012 ( .A(n2624), .B(n1869), .Z(out[134]) );
  XOR U3013 ( .A(in[433]), .B(n3998), .Z(n2081) );
  NOR U3014 ( .A(n1947), .B(n2235), .Z(n1870) );
  XNOR U3015 ( .A(n2081), .B(n1870), .Z(out[1350]) );
  XOR U3016 ( .A(in[434]), .B(n4001), .Z(n2083) );
  NOR U3017 ( .A(n1949), .B(n2238), .Z(n1871) );
  XNOR U3018 ( .A(n2083), .B(n1871), .Z(out[1351]) );
  XOR U3019 ( .A(in[435]), .B(n4008), .Z(n2086) );
  NOR U3020 ( .A(n1951), .B(n2244), .Z(n1872) );
  XNOR U3021 ( .A(n2086), .B(n1872), .Z(out[1352]) );
  XOR U3022 ( .A(in[436]), .B(n4011), .Z(n2088) );
  NOR U3023 ( .A(n1953), .B(n2248), .Z(n1873) );
  XNOR U3024 ( .A(n2088), .B(n1873), .Z(out[1353]) );
  XOR U3025 ( .A(in[437]), .B(n4014), .Z(n2090) );
  NOR U3026 ( .A(n1955), .B(n2252), .Z(n1874) );
  XNOR U3027 ( .A(n2090), .B(n1874), .Z(out[1354]) );
  XOR U3028 ( .A(in[438]), .B(n4017), .Z(n2092) );
  NOR U3029 ( .A(n1957), .B(n2256), .Z(n1875) );
  XNOR U3030 ( .A(n2092), .B(n1875), .Z(out[1355]) );
  XOR U3031 ( .A(in[439]), .B(n4020), .Z(n2094) );
  NOR U3032 ( .A(n1960), .B(n2260), .Z(n1876) );
  XNOR U3033 ( .A(n2094), .B(n1876), .Z(out[1356]) );
  XOR U3034 ( .A(in[440]), .B(n4023), .Z(n2096) );
  NOR U3035 ( .A(n1962), .B(n2264), .Z(n1877) );
  XNOR U3036 ( .A(n2096), .B(n1877), .Z(out[1357]) );
  XOR U3037 ( .A(in[441]), .B(n4026), .Z(n2098) );
  NOR U3038 ( .A(n1964), .B(n2269), .Z(n1878) );
  XNOR U3039 ( .A(n2098), .B(n1878), .Z(out[1358]) );
  XOR U3040 ( .A(in[442]), .B(n4029), .Z(n2100) );
  NOR U3041 ( .A(n1966), .B(n2272), .Z(n1879) );
  XNOR U3042 ( .A(n2100), .B(n1879), .Z(out[1359]) );
  XNOR U3043 ( .A(in[672]), .B(n3908), .Z(n2626) );
  XNOR U3044 ( .A(in[606]), .B(n3744), .Z(n3855) );
  XOR U3045 ( .A(in[197]), .B(n3561), .Z(n4079) );
  NAND U3046 ( .A(n3855), .B(n4079), .Z(n1880) );
  XNOR U3047 ( .A(n2626), .B(n1880), .Z(out[135]) );
  XOR U3048 ( .A(in[443]), .B(n4032), .Z(n2102) );
  NOR U3049 ( .A(n1968), .B(n2278), .Z(n1881) );
  XNOR U3050 ( .A(n2102), .B(n1881), .Z(out[1360]) );
  XOR U3051 ( .A(in[444]), .B(n4035), .Z(n2104) );
  NOR U3052 ( .A(n1970), .B(n2282), .Z(n1882) );
  XNOR U3053 ( .A(n2104), .B(n1882), .Z(out[1361]) );
  XOR U3054 ( .A(in[445]), .B(n4042), .Z(n2107) );
  NOR U3055 ( .A(n1972), .B(n2286), .Z(n1883) );
  XNOR U3056 ( .A(n2107), .B(n1883), .Z(out[1362]) );
  XOR U3057 ( .A(in[446]), .B(n4045), .Z(n2109) );
  NOR U3058 ( .A(n1974), .B(n2290), .Z(n1884) );
  XNOR U3059 ( .A(n2109), .B(n1884), .Z(out[1363]) );
  XOR U3060 ( .A(in[447]), .B(n4048), .Z(n2111) );
  NOR U3061 ( .A(n1976), .B(n2294), .Z(n1885) );
  XNOR U3062 ( .A(n2111), .B(n1885), .Z(out[1364]) );
  XOR U3063 ( .A(in[384]), .B(n4051), .Z(n2113) );
  NOR U3064 ( .A(n1978), .B(n2298), .Z(n1886) );
  XNOR U3065 ( .A(n2113), .B(n1886), .Z(out[1365]) );
  XOR U3066 ( .A(in[385]), .B(n4054), .Z(n2115) );
  NOR U3067 ( .A(n1981), .B(n2302), .Z(n1887) );
  XNOR U3068 ( .A(n2115), .B(n1887), .Z(out[1366]) );
  XOR U3069 ( .A(in[386]), .B(n4057), .Z(n2117) );
  NOR U3070 ( .A(n1983), .B(n2306), .Z(n1888) );
  XNOR U3071 ( .A(n2117), .B(n1888), .Z(out[1367]) );
  XOR U3072 ( .A(in[387]), .B(n4060), .Z(n2119) );
  NOR U3073 ( .A(n1985), .B(n2311), .Z(n1889) );
  XNOR U3074 ( .A(n2119), .B(n1889), .Z(out[1368]) );
  XOR U3075 ( .A(in[388]), .B(n4063), .Z(n2121) );
  NOR U3076 ( .A(n1987), .B(n2315), .Z(n1890) );
  XNOR U3077 ( .A(n2121), .B(n1890), .Z(out[1369]) );
  XNOR U3078 ( .A(in[673]), .B(n3910), .Z(n2628) );
  XNOR U3079 ( .A(in[607]), .B(n3748), .Z(n3877) );
  XOR U3080 ( .A(in[198]), .B(n3565), .Z(n4363) );
  NAND U3081 ( .A(n3877), .B(n4363), .Z(n1891) );
  XNOR U3082 ( .A(n2628), .B(n1891), .Z(out[136]) );
  XOR U3083 ( .A(in[389]), .B(n4066), .Z(n2123) );
  NOR U3084 ( .A(n1989), .B(n2319), .Z(n1892) );
  XNOR U3085 ( .A(n2123), .B(n1892), .Z(out[1370]) );
  XOR U3086 ( .A(in[390]), .B(n4069), .Z(n2125) );
  NOR U3087 ( .A(n1991), .B(n2323), .Z(n1893) );
  XNOR U3088 ( .A(n2125), .B(n1893), .Z(out[1371]) );
  XOR U3089 ( .A(in[391]), .B(n4080), .Z(n2129) );
  NOR U3090 ( .A(n1993), .B(n2327), .Z(n1894) );
  XNOR U3091 ( .A(n2129), .B(n1894), .Z(out[1372]) );
  XOR U3092 ( .A(in[392]), .B(n4083), .Z(n2131) );
  NOR U3093 ( .A(n1995), .B(n2331), .Z(n1895) );
  XNOR U3094 ( .A(n2131), .B(n1895), .Z(out[1373]) );
  XOR U3095 ( .A(in[393]), .B(n4086), .Z(n2133) );
  NOR U3096 ( .A(n1997), .B(n2335), .Z(n1896) );
  XNOR U3097 ( .A(n2133), .B(n1896), .Z(out[1374]) );
  XOR U3098 ( .A(in[394]), .B(n4089), .Z(n2135) );
  NOR U3099 ( .A(n1999), .B(n2338), .Z(n1897) );
  XNOR U3100 ( .A(n2135), .B(n1897), .Z(out[1375]) );
  XOR U3101 ( .A(in[395]), .B(n4092), .Z(n2137) );
  NOR U3102 ( .A(n2002), .B(n2344), .Z(n1898) );
  XNOR U3103 ( .A(n2137), .B(n1898), .Z(out[1376]) );
  XNOR U3104 ( .A(n4095), .B(in[396]), .Z(n2139) );
  NOR U3105 ( .A(n2004), .B(n2348), .Z(n1899) );
  XNOR U3106 ( .A(n2139), .B(n1899), .Z(out[1377]) );
  XNOR U3107 ( .A(n4098), .B(in[397]), .Z(n2141) );
  NOR U3108 ( .A(n2006), .B(n2353), .Z(n1900) );
  XNOR U3109 ( .A(n2141), .B(n1900), .Z(out[1378]) );
  XNOR U3110 ( .A(n4101), .B(in[398]), .Z(n2143) );
  NOR U3111 ( .A(n2008), .B(n2357), .Z(n1901) );
  XNOR U3112 ( .A(n2143), .B(n1901), .Z(out[1379]) );
  XNOR U3113 ( .A(in[674]), .B(n3912), .Z(n2630) );
  XNOR U3114 ( .A(in[608]), .B(n3756), .Z(n3899) );
  XOR U3115 ( .A(in[199]), .B(n3569), .Z(n4807) );
  NAND U3116 ( .A(n3899), .B(n4807), .Z(n1902) );
  XNOR U3117 ( .A(n2630), .B(n1902), .Z(out[137]) );
  XNOR U3118 ( .A(n4104), .B(in[399]), .Z(n2145) );
  NOR U3119 ( .A(n2010), .B(n2361), .Z(n1903) );
  XNOR U3120 ( .A(n2145), .B(n1903), .Z(out[1380]) );
  XNOR U3121 ( .A(n4107), .B(in[400]), .Z(n2147) );
  NOR U3122 ( .A(n2012), .B(n2365), .Z(n1904) );
  XNOR U3123 ( .A(n2147), .B(n1904), .Z(out[1381]) );
  XNOR U3124 ( .A(n4114), .B(in[401]), .Z(n2150) );
  NOR U3125 ( .A(n2014), .B(n2369), .Z(n1905) );
  XNOR U3126 ( .A(n2150), .B(n1905), .Z(out[1382]) );
  XNOR U3127 ( .A(n4117), .B(in[402]), .Z(n2152) );
  NOR U3128 ( .A(n2016), .B(n2373), .Z(n1906) );
  XNOR U3129 ( .A(n2152), .B(n1906), .Z(out[1383]) );
  XNOR U3130 ( .A(n4120), .B(in[403]), .Z(n2154) );
  NOR U3131 ( .A(n2018), .B(n2377), .Z(n1907) );
  XNOR U3132 ( .A(n2154), .B(n1907), .Z(out[1384]) );
  XNOR U3133 ( .A(in[404]), .B(n4123), .Z(n2156) );
  NOR U3134 ( .A(n2020), .B(n2381), .Z(n1908) );
  XNOR U3135 ( .A(n2156), .B(n1908), .Z(out[1385]) );
  XNOR U3136 ( .A(in[405]), .B(n4126), .Z(n2158) );
  NOR U3137 ( .A(n2023), .B(n2385), .Z(n1909) );
  XNOR U3138 ( .A(n2158), .B(n1909), .Z(out[1386]) );
  XNOR U3139 ( .A(in[406]), .B(n4129), .Z(n2160) );
  NOR U3140 ( .A(n2025), .B(n2389), .Z(n1910) );
  XNOR U3141 ( .A(n2160), .B(n1910), .Z(out[1387]) );
  XNOR U3142 ( .A(in[407]), .B(n4132), .Z(n2162) );
  NOR U3143 ( .A(n2027), .B(n2394), .Z(n1911) );
  XNOR U3144 ( .A(n2162), .B(n1911), .Z(out[1388]) );
  XNOR U3145 ( .A(in[408]), .B(n4135), .Z(n2164) );
  NOR U3146 ( .A(n2029), .B(n2398), .Z(n1912) );
  XNOR U3147 ( .A(n2164), .B(n1912), .Z(out[1389]) );
  XNOR U3148 ( .A(in[675]), .B(n3914), .Z(n2633) );
  XNOR U3149 ( .A(in[609]), .B(n3760), .Z(n3923) );
  NAND U3150 ( .A(n3923), .B(n3921), .Z(n1913) );
  XNOR U3151 ( .A(n2633), .B(n1913), .Z(out[138]) );
  XNOR U3152 ( .A(in[409]), .B(n4138), .Z(n2166) );
  NOR U3153 ( .A(n2031), .B(n2402), .Z(n1914) );
  XNOR U3154 ( .A(n2166), .B(n1914), .Z(out[1390]) );
  XNOR U3155 ( .A(in[410]), .B(n4141), .Z(n2168) );
  NOR U3156 ( .A(n2033), .B(n2406), .Z(n1915) );
  XNOR U3157 ( .A(n2168), .B(n1915), .Z(out[1391]) );
  XNOR U3158 ( .A(in[411]), .B(n4148), .Z(n2171) );
  NOR U3159 ( .A(n2035), .B(n2410), .Z(n1916) );
  XNOR U3160 ( .A(n2171), .B(n1916), .Z(out[1392]) );
  XNOR U3161 ( .A(in[412]), .B(n4151), .Z(n2173) );
  NOR U3162 ( .A(n2037), .B(n2414), .Z(n1917) );
  XNOR U3163 ( .A(n2173), .B(n1917), .Z(out[1393]) );
  XNOR U3164 ( .A(in[413]), .B(n4154), .Z(n2175) );
  NOR U3165 ( .A(n2039), .B(n2418), .Z(n1918) );
  XNOR U3166 ( .A(n2175), .B(n1918), .Z(out[1394]) );
  XNOR U3167 ( .A(in[414]), .B(n4157), .Z(n2177) );
  NOR U3168 ( .A(n2041), .B(n2422), .Z(n1919) );
  XNOR U3169 ( .A(n2177), .B(n1919), .Z(out[1395]) );
  XNOR U3170 ( .A(in[415]), .B(n4160), .Z(n2179) );
  NOR U3171 ( .A(n2044), .B(n2426), .Z(n1920) );
  XNOR U3172 ( .A(n2179), .B(n1920), .Z(out[1396]) );
  XNOR U3173 ( .A(in[416]), .B(n4163), .Z(n2181) );
  NOR U3174 ( .A(n2046), .B(n2430), .Z(n1921) );
  XNOR U3175 ( .A(n2181), .B(n1921), .Z(out[1397]) );
  XNOR U3176 ( .A(in[417]), .B(n4166), .Z(n2183) );
  NOR U3177 ( .A(n2048), .B(n2435), .Z(n1922) );
  XNOR U3178 ( .A(n2183), .B(n1922), .Z(out[1398]) );
  XNOR U3179 ( .A(in[418]), .B(n4169), .Z(n2185) );
  NOR U3180 ( .A(n2050), .B(n2439), .Z(n1923) );
  XNOR U3181 ( .A(n2185), .B(n1923), .Z(out[1399]) );
  XNOR U3182 ( .A(in[676]), .B(n3916), .Z(n2636) );
  XNOR U3183 ( .A(in[610]), .B(n3764), .Z(n3947) );
  NAND U3184 ( .A(n3947), .B(n3945), .Z(n1924) );
  XNOR U3185 ( .A(n2636), .B(n1924), .Z(out[139]) );
  XOR U3186 ( .A(in[203]), .B(n3589), .Z(n4005) );
  XNOR U3187 ( .A(in[1423]), .B(n3630), .Z(n4004) );
  XOR U3188 ( .A(in[1046]), .B(n4129), .Z(n2641) );
  NAND U3189 ( .A(n4004), .B(n2641), .Z(n1925) );
  XNOR U3190 ( .A(n4005), .B(n1925), .Z(out[13]) );
  XNOR U3191 ( .A(in[419]), .B(n4172), .Z(n2187) );
  NOR U3192 ( .A(n2052), .B(n2443), .Z(n1926) );
  XNOR U3193 ( .A(n2187), .B(n1926), .Z(out[1400]) );
  XOR U3194 ( .A(in[420]), .B(n4175), .Z(n2189) );
  NOR U3195 ( .A(n2054), .B(n2447), .Z(n1927) );
  XNOR U3196 ( .A(n2189), .B(n1927), .Z(out[1401]) );
  XOR U3197 ( .A(in[421]), .B(n4182), .Z(n2192) );
  NOR U3198 ( .A(n2056), .B(n2451), .Z(n1928) );
  XNOR U3199 ( .A(n2192), .B(n1928), .Z(out[1402]) );
  XOR U3200 ( .A(in[422]), .B(n4185), .Z(n2194) );
  NOR U3201 ( .A(n2058), .B(n2455), .Z(n1929) );
  XNOR U3202 ( .A(n2194), .B(n1929), .Z(out[1403]) );
  XOR U3203 ( .A(in[423]), .B(n3964), .Z(n2196) );
  NOR U3204 ( .A(n2060), .B(n2459), .Z(n1930) );
  XNOR U3205 ( .A(n2196), .B(n1930), .Z(out[1404]) );
  XOR U3206 ( .A(in[424]), .B(n3967), .Z(n2198) );
  NOR U3207 ( .A(n2062), .B(n2463), .Z(n1931) );
  XNOR U3208 ( .A(n2198), .B(n1931), .Z(out[1405]) );
  XOR U3209 ( .A(in[425]), .B(n3974), .Z(n2200) );
  NOR U3210 ( .A(n2065), .B(n2467), .Z(n1932) );
  XNOR U3211 ( .A(n2200), .B(n1932), .Z(out[1406]) );
  XOR U3212 ( .A(in[426]), .B(n3977), .Z(n2202) );
  NOR U3213 ( .A(n2067), .B(n2470), .Z(n1933) );
  XNOR U3214 ( .A(n2202), .B(n1933), .Z(out[1407]) );
  XOR U3215 ( .A(in[789]), .B(n3654), .Z(n2205) );
  NAND U3216 ( .A(n2069), .B(n1934), .Z(n1935) );
  XNOR U3217 ( .A(n2205), .B(n1935), .Z(out[1408]) );
  XOR U3218 ( .A(in[790]), .B(n3658), .Z(n2210) );
  NAND U3219 ( .A(n2071), .B(n1936), .Z(n1937) );
  XNOR U3220 ( .A(n2210), .B(n1937), .Z(out[1409]) );
  XNOR U3221 ( .A(in[677]), .B(n3918), .Z(n2639) );
  XNOR U3222 ( .A(in[611]), .B(n3768), .Z(n3973) );
  NAND U3223 ( .A(n3973), .B(n3971), .Z(n1938) );
  XNOR U3224 ( .A(n2639), .B(n1938), .Z(out[140]) );
  XOR U3225 ( .A(in[791]), .B(n3662), .Z(n2215) );
  NAND U3226 ( .A(n2073), .B(n1939), .Z(n1940) );
  XNOR U3227 ( .A(n2215), .B(n1940), .Z(out[1410]) );
  XOR U3228 ( .A(in[792]), .B(n3670), .Z(n2219) );
  NAND U3229 ( .A(n2075), .B(n1941), .Z(n1942) );
  XNOR U3230 ( .A(n2219), .B(n1942), .Z(out[1411]) );
  XOR U3231 ( .A(in[793]), .B(n3674), .Z(n2225) );
  NAND U3232 ( .A(n2077), .B(n1943), .Z(n1944) );
  XNOR U3233 ( .A(n2225), .B(n1944), .Z(out[1412]) );
  XOR U3234 ( .A(in[794]), .B(n3678), .Z(n2229) );
  NAND U3235 ( .A(n2079), .B(n1945), .Z(n1946) );
  XNOR U3236 ( .A(n2229), .B(n1946), .Z(out[1413]) );
  XOR U3237 ( .A(in[795]), .B(n3682), .Z(n2233) );
  NAND U3238 ( .A(n2081), .B(n1947), .Z(n1948) );
  XNOR U3239 ( .A(n2233), .B(n1948), .Z(out[1414]) );
  XOR U3240 ( .A(in[796]), .B(n3686), .Z(n2237) );
  NAND U3241 ( .A(n2083), .B(n1949), .Z(n1950) );
  XNOR U3242 ( .A(n2237), .B(n1950), .Z(out[1415]) );
  XOR U3243 ( .A(in[797]), .B(n3690), .Z(n2242) );
  NAND U3244 ( .A(n2086), .B(n1951), .Z(n1952) );
  XNOR U3245 ( .A(n2242), .B(n1952), .Z(out[1416]) );
  XOR U3246 ( .A(in[798]), .B(n3694), .Z(n2246) );
  NAND U3247 ( .A(n2088), .B(n1953), .Z(n1954) );
  XNOR U3248 ( .A(n2246), .B(n1954), .Z(out[1417]) );
  XOR U3249 ( .A(in[799]), .B(n3698), .Z(n2250) );
  NAND U3250 ( .A(n2090), .B(n1955), .Z(n1956) );
  XNOR U3251 ( .A(n2250), .B(n1956), .Z(out[1418]) );
  XOR U3252 ( .A(in[800]), .B(n3702), .Z(n2254) );
  NAND U3253 ( .A(n2092), .B(n1957), .Z(n1958) );
  XNOR U3254 ( .A(n2254), .B(n1958), .Z(out[1419]) );
  XNOR U3255 ( .A(in[678]), .B(n3924), .Z(n2642) );
  XNOR U3256 ( .A(in[612]), .B(n3772), .Z(n4007) );
  NAND U3257 ( .A(n4007), .B(n4005), .Z(n1959) );
  XNOR U3258 ( .A(n2642), .B(n1959), .Z(out[141]) );
  XOR U3259 ( .A(in[801]), .B(n3706), .Z(n2258) );
  NAND U3260 ( .A(n2094), .B(n1960), .Z(n1961) );
  XNOR U3261 ( .A(n2258), .B(n1961), .Z(out[1420]) );
  XOR U3262 ( .A(in[802]), .B(n3714), .Z(n2262) );
  NAND U3263 ( .A(n2096), .B(n1962), .Z(n1963) );
  XNOR U3264 ( .A(n2262), .B(n1963), .Z(out[1421]) );
  XOR U3265 ( .A(in[803]), .B(n3718), .Z(n2267) );
  NAND U3266 ( .A(n2098), .B(n1964), .Z(n1965) );
  XNOR U3267 ( .A(n2267), .B(n1965), .Z(out[1422]) );
  XOR U3268 ( .A(in[804]), .B(n3722), .Z(n2271) );
  NAND U3269 ( .A(n2100), .B(n1966), .Z(n1967) );
  XNOR U3270 ( .A(n2271), .B(n1967), .Z(out[1423]) );
  XOR U3271 ( .A(in[805]), .B(n3726), .Z(n2276) );
  NAND U3272 ( .A(n2102), .B(n1968), .Z(n1969) );
  XNOR U3273 ( .A(n2276), .B(n1969), .Z(out[1424]) );
  XNOR U3274 ( .A(in[806]), .B(n3730), .Z(n2280) );
  NAND U3275 ( .A(n2104), .B(n1970), .Z(n1971) );
  XNOR U3276 ( .A(n2280), .B(n1971), .Z(out[1425]) );
  XNOR U3277 ( .A(in[807]), .B(n3734), .Z(n2284) );
  NAND U3278 ( .A(n2107), .B(n1972), .Z(n1973) );
  XNOR U3279 ( .A(n2284), .B(n1973), .Z(out[1426]) );
  XNOR U3280 ( .A(in[808]), .B(n3738), .Z(n2288) );
  NAND U3281 ( .A(n2109), .B(n1974), .Z(n1975) );
  XNOR U3282 ( .A(n2288), .B(n1975), .Z(out[1427]) );
  XNOR U3283 ( .A(in[809]), .B(n3742), .Z(n2292) );
  NAND U3284 ( .A(n2111), .B(n1976), .Z(n1977) );
  XNOR U3285 ( .A(n2292), .B(n1977), .Z(out[1428]) );
  XNOR U3286 ( .A(in[810]), .B(n3746), .Z(n2296) );
  NAND U3287 ( .A(n2113), .B(n1978), .Z(n1979) );
  XNOR U3288 ( .A(n2296), .B(n1979), .Z(out[1429]) );
  XNOR U3289 ( .A(in[679]), .B(n3926), .Z(n2646) );
  XOR U3290 ( .A(in[613]), .B(n3776), .Z(n4041) );
  XOR U3291 ( .A(in[204]), .B(n3593), .Z(n4039) );
  NAND U3292 ( .A(n4041), .B(n4039), .Z(n1980) );
  XNOR U3293 ( .A(n2646), .B(n1980), .Z(out[142]) );
  XNOR U3294 ( .A(in[811]), .B(n3750), .Z(n2300) );
  NAND U3295 ( .A(n2115), .B(n1981), .Z(n1982) );
  XNOR U3296 ( .A(n2300), .B(n1982), .Z(out[1430]) );
  XNOR U3297 ( .A(in[812]), .B(n3758), .Z(n2304) );
  NAND U3298 ( .A(n2117), .B(n1983), .Z(n1984) );
  XNOR U3299 ( .A(n2304), .B(n1984), .Z(out[1431]) );
  XNOR U3300 ( .A(in[813]), .B(n3762), .Z(n2309) );
  NAND U3301 ( .A(n2119), .B(n1985), .Z(n1986) );
  XNOR U3302 ( .A(n2309), .B(n1986), .Z(out[1432]) );
  XNOR U3303 ( .A(in[814]), .B(n3766), .Z(n2313) );
  NAND U3304 ( .A(n2121), .B(n1987), .Z(n1988) );
  XNOR U3305 ( .A(n2313), .B(n1988), .Z(out[1433]) );
  XNOR U3306 ( .A(in[815]), .B(n3770), .Z(n2317) );
  NAND U3307 ( .A(n2123), .B(n1989), .Z(n1990) );
  XNOR U3308 ( .A(n2317), .B(n1990), .Z(out[1434]) );
  XNOR U3309 ( .A(in[816]), .B(n3774), .Z(n2321) );
  NAND U3310 ( .A(n2125), .B(n1991), .Z(n1992) );
  XNOR U3311 ( .A(n2321), .B(n1992), .Z(out[1435]) );
  XNOR U3312 ( .A(in[817]), .B(n3778), .Z(n2325) );
  NAND U3313 ( .A(n2129), .B(n1993), .Z(n1994) );
  XNOR U3314 ( .A(n2325), .B(n1994), .Z(out[1436]) );
  XNOR U3315 ( .A(in[818]), .B(n3782), .Z(n2329) );
  NAND U3316 ( .A(n2131), .B(n1995), .Z(n1996) );
  XNOR U3317 ( .A(n2329), .B(n1996), .Z(out[1437]) );
  XNOR U3318 ( .A(in[819]), .B(n3786), .Z(n2333) );
  NAND U3319 ( .A(n2133), .B(n1997), .Z(n1998) );
  XNOR U3320 ( .A(n2333), .B(n1998), .Z(out[1438]) );
  XNOR U3321 ( .A(in[820]), .B(n3790), .Z(n2337) );
  NAND U3322 ( .A(n2135), .B(n1999), .Z(n2000) );
  XNOR U3323 ( .A(n2337), .B(n2000), .Z(out[1439]) );
  XNOR U3324 ( .A(in[680]), .B(n3928), .Z(n2649) );
  XOR U3325 ( .A(in[614]), .B(n3780), .Z(n4075) );
  XOR U3326 ( .A(in[205]), .B(n3597), .Z(n4073) );
  NAND U3327 ( .A(n4075), .B(n4073), .Z(n2001) );
  XNOR U3328 ( .A(n2649), .B(n2001), .Z(out[143]) );
  XNOR U3329 ( .A(in[821]), .B(n3794), .Z(n2342) );
  NAND U3330 ( .A(n2137), .B(n2002), .Z(n2003) );
  XNOR U3331 ( .A(n2342), .B(n2003), .Z(out[1440]) );
  XNOR U3332 ( .A(in[822]), .B(n3804), .Z(n2346) );
  NAND U3333 ( .A(n2139), .B(n2004), .Z(n2005) );
  XNOR U3334 ( .A(n2346), .B(n2005), .Z(out[1441]) );
  XNOR U3335 ( .A(in[823]), .B(n3808), .Z(n2351) );
  NAND U3336 ( .A(n2141), .B(n2006), .Z(n2007) );
  XNOR U3337 ( .A(n2351), .B(n2007), .Z(out[1442]) );
  XNOR U3338 ( .A(in[824]), .B(n3812), .Z(n2355) );
  NAND U3339 ( .A(n2143), .B(n2008), .Z(n2009) );
  XNOR U3340 ( .A(n2355), .B(n2009), .Z(out[1443]) );
  XNOR U3341 ( .A(in[825]), .B(n3816), .Z(n2359) );
  NAND U3342 ( .A(n2145), .B(n2010), .Z(n2011) );
  XNOR U3343 ( .A(n2359), .B(n2011), .Z(out[1444]) );
  XNOR U3344 ( .A(in[826]), .B(n3538), .Z(n2363) );
  NAND U3345 ( .A(n2147), .B(n2012), .Z(n2013) );
  XNOR U3346 ( .A(n2363), .B(n2013), .Z(out[1445]) );
  XNOR U3347 ( .A(in[827]), .B(n3542), .Z(n2367) );
  NAND U3348 ( .A(n2150), .B(n2014), .Z(n2015) );
  XNOR U3349 ( .A(n2367), .B(n2015), .Z(out[1446]) );
  XNOR U3350 ( .A(in[828]), .B(n3546), .Z(n2371) );
  NAND U3351 ( .A(n2152), .B(n2016), .Z(n2017) );
  XNOR U3352 ( .A(n2371), .B(n2017), .Z(out[1447]) );
  XNOR U3353 ( .A(in[829]), .B(n3550), .Z(n2375) );
  NAND U3354 ( .A(n2154), .B(n2018), .Z(n2019) );
  XNOR U3355 ( .A(n2375), .B(n2019), .Z(out[1448]) );
  XNOR U3356 ( .A(in[830]), .B(n3554), .Z(n2379) );
  NAND U3357 ( .A(n2156), .B(n2020), .Z(n2021) );
  XNOR U3358 ( .A(n2379), .B(n2021), .Z(out[1449]) );
  XNOR U3359 ( .A(in[681]), .B(n3930), .Z(n2652) );
  XOR U3360 ( .A(in[615]), .B(n3784), .Z(n4113) );
  XOR U3361 ( .A(in[206]), .B(n3601), .Z(n4111) );
  NAND U3362 ( .A(n4113), .B(n4111), .Z(n2022) );
  XNOR U3363 ( .A(n2652), .B(n2022), .Z(out[144]) );
  XNOR U3364 ( .A(in[831]), .B(n3558), .Z(n2383) );
  NAND U3365 ( .A(n2158), .B(n2023), .Z(n2024) );
  XNOR U3366 ( .A(n2383), .B(n2024), .Z(out[1450]) );
  XNOR U3367 ( .A(in[768]), .B(n3562), .Z(n2387) );
  NAND U3368 ( .A(n2160), .B(n2025), .Z(n2026) );
  XNOR U3369 ( .A(n2387), .B(n2026), .Z(out[1451]) );
  XNOR U3370 ( .A(in[769]), .B(n3566), .Z(n2392) );
  NAND U3371 ( .A(n2162), .B(n2027), .Z(n2028) );
  XNOR U3372 ( .A(n2392), .B(n2028), .Z(out[1452]) );
  XOR U3373 ( .A(n3570), .B(in[770]), .Z(n2396) );
  NAND U3374 ( .A(n2164), .B(n2029), .Z(n2030) );
  XNOR U3375 ( .A(n2396), .B(n2030), .Z(out[1453]) );
  XOR U3376 ( .A(n3574), .B(in[771]), .Z(n2400) );
  NAND U3377 ( .A(n2166), .B(n2031), .Z(n2032) );
  XNOR U3378 ( .A(n2400), .B(n2032), .Z(out[1454]) );
  XOR U3379 ( .A(n3582), .B(in[772]), .Z(n2404) );
  NAND U3380 ( .A(n2168), .B(n2033), .Z(n2034) );
  XNOR U3381 ( .A(n2404), .B(n2034), .Z(out[1455]) );
  XOR U3382 ( .A(n3586), .B(in[773]), .Z(n2408) );
  NAND U3383 ( .A(n2171), .B(n2035), .Z(n2036) );
  XNOR U3384 ( .A(n2408), .B(n2036), .Z(out[1456]) );
  XOR U3385 ( .A(n3590), .B(in[774]), .Z(n2412) );
  NAND U3386 ( .A(n2173), .B(n2037), .Z(n2038) );
  XNOR U3387 ( .A(n2412), .B(n2038), .Z(out[1457]) );
  XOR U3388 ( .A(n3594), .B(in[775]), .Z(n2416) );
  NAND U3389 ( .A(n2175), .B(n2039), .Z(n2040) );
  XNOR U3390 ( .A(n2416), .B(n2040), .Z(out[1458]) );
  XOR U3391 ( .A(n3598), .B(in[776]), .Z(n2420) );
  NAND U3392 ( .A(n2177), .B(n2041), .Z(n2042) );
  XNOR U3393 ( .A(n2420), .B(n2042), .Z(out[1459]) );
  XNOR U3394 ( .A(in[682]), .B(n3932), .Z(n2655) );
  XOR U3395 ( .A(in[616]), .B(n3788), .Z(n4147) );
  XOR U3396 ( .A(in[207]), .B(n3605), .Z(n4145) );
  NAND U3397 ( .A(n4147), .B(n4145), .Z(n2043) );
  XNOR U3398 ( .A(n2655), .B(n2043), .Z(out[145]) );
  XOR U3399 ( .A(in[777]), .B(n3602), .Z(n2424) );
  NAND U3400 ( .A(n2179), .B(n2044), .Z(n2045) );
  XNOR U3401 ( .A(n2424), .B(n2045), .Z(out[1460]) );
  XOR U3402 ( .A(n3606), .B(in[778]), .Z(n2428) );
  NAND U3403 ( .A(n2181), .B(n2046), .Z(n2047) );
  XNOR U3404 ( .A(n2428), .B(n2047), .Z(out[1461]) );
  XOR U3405 ( .A(n3610), .B(in[779]), .Z(n2433) );
  NAND U3406 ( .A(n2183), .B(n2048), .Z(n2049) );
  XNOR U3407 ( .A(n2433), .B(n2049), .Z(out[1462]) );
  XOR U3408 ( .A(in[780]), .B(n3614), .Z(n2437) );
  NAND U3409 ( .A(n2185), .B(n2050), .Z(n2051) );
  XNOR U3410 ( .A(n2437), .B(n2051), .Z(out[1463]) );
  XOR U3411 ( .A(in[781]), .B(n3618), .Z(n2441) );
  NAND U3412 ( .A(n2187), .B(n2052), .Z(n2053) );
  XNOR U3413 ( .A(n2441), .B(n2053), .Z(out[1464]) );
  XOR U3414 ( .A(in[782]), .B(n3626), .Z(n2445) );
  NAND U3415 ( .A(n2189), .B(n2054), .Z(n2055) );
  XNOR U3416 ( .A(n2445), .B(n2055), .Z(out[1465]) );
  XOR U3417 ( .A(in[783]), .B(n3630), .Z(n2449) );
  NAND U3418 ( .A(n2192), .B(n2056), .Z(n2057) );
  XNOR U3419 ( .A(n2449), .B(n2057), .Z(out[1466]) );
  XOR U3420 ( .A(in[784]), .B(n3634), .Z(n2453) );
  NAND U3421 ( .A(n2194), .B(n2058), .Z(n2059) );
  XNOR U3422 ( .A(n2453), .B(n2059), .Z(out[1467]) );
  XOR U3423 ( .A(in[785]), .B(n3638), .Z(n2457) );
  NAND U3424 ( .A(n2196), .B(n2060), .Z(n2061) );
  XNOR U3425 ( .A(n2457), .B(n2061), .Z(out[1468]) );
  XOR U3426 ( .A(in[786]), .B(n3642), .Z(n2461) );
  NAND U3427 ( .A(n2198), .B(n2062), .Z(n2063) );
  XNOR U3428 ( .A(n2461), .B(n2063), .Z(out[1469]) );
  XNOR U3429 ( .A(in[683]), .B(n3934), .Z(n2658) );
  XOR U3430 ( .A(in[617]), .B(n3792), .Z(n4181) );
  XOR U3431 ( .A(in[208]), .B(n3609), .Z(n4179) );
  NAND U3432 ( .A(n4181), .B(n4179), .Z(n2064) );
  XNOR U3433 ( .A(n2658), .B(n2064), .Z(out[146]) );
  XOR U3434 ( .A(in[787]), .B(n3646), .Z(n2465) );
  NAND U3435 ( .A(n2200), .B(n2065), .Z(n2066) );
  XNOR U3436 ( .A(n2465), .B(n2066), .Z(out[1470]) );
  XOR U3437 ( .A(in[788]), .B(n3650), .Z(n2469) );
  NAND U3438 ( .A(n2202), .B(n2067), .Z(n2068) );
  XNOR U3439 ( .A(n2469), .B(n2068), .Z(out[1471]) );
  OR U3440 ( .A(n2205), .B(n2069), .Z(n2070) );
  XNOR U3441 ( .A(n2204), .B(n2070), .Z(out[1472]) );
  OR U3442 ( .A(n2210), .B(n2071), .Z(n2072) );
  XNOR U3443 ( .A(n2209), .B(n2072), .Z(out[1473]) );
  OR U3444 ( .A(n2215), .B(n2073), .Z(n2074) );
  XNOR U3445 ( .A(n2214), .B(n2074), .Z(out[1474]) );
  OR U3446 ( .A(n2219), .B(n2075), .Z(n2076) );
  XNOR U3447 ( .A(n2218), .B(n2076), .Z(out[1475]) );
  OR U3448 ( .A(n2225), .B(n2077), .Z(n2078) );
  XNOR U3449 ( .A(n2224), .B(n2078), .Z(out[1476]) );
  OR U3450 ( .A(n2229), .B(n2079), .Z(n2080) );
  XNOR U3451 ( .A(n2228), .B(n2080), .Z(out[1477]) );
  OR U3452 ( .A(n2233), .B(n2081), .Z(n2082) );
  XNOR U3453 ( .A(n2232), .B(n2082), .Z(out[1478]) );
  OR U3454 ( .A(n2237), .B(n2083), .Z(n2084) );
  XNOR U3455 ( .A(n2236), .B(n2084), .Z(out[1479]) );
  XNOR U3456 ( .A(in[684]), .B(n3936), .Z(n2661) );
  XOR U3457 ( .A(in[618]), .B(n3802), .Z(n4207) );
  XOR U3458 ( .A(in[209]), .B(n3613), .Z(n4205) );
  NAND U3459 ( .A(n4207), .B(n4205), .Z(n2085) );
  XNOR U3460 ( .A(n2661), .B(n2085), .Z(out[147]) );
  OR U3461 ( .A(n2242), .B(n2086), .Z(n2087) );
  XNOR U3462 ( .A(n2241), .B(n2087), .Z(out[1480]) );
  OR U3463 ( .A(n2246), .B(n2088), .Z(n2089) );
  XNOR U3464 ( .A(n2245), .B(n2089), .Z(out[1481]) );
  OR U3465 ( .A(n2250), .B(n2090), .Z(n2091) );
  XNOR U3466 ( .A(n2249), .B(n2091), .Z(out[1482]) );
  OR U3467 ( .A(n2254), .B(n2092), .Z(n2093) );
  XNOR U3468 ( .A(n2253), .B(n2093), .Z(out[1483]) );
  OR U3469 ( .A(n2258), .B(n2094), .Z(n2095) );
  XNOR U3470 ( .A(n2257), .B(n2095), .Z(out[1484]) );
  OR U3471 ( .A(n2262), .B(n2096), .Z(n2097) );
  XNOR U3472 ( .A(n2261), .B(n2097), .Z(out[1485]) );
  OR U3473 ( .A(n2267), .B(n2098), .Z(n2099) );
  XNOR U3474 ( .A(n2266), .B(n2099), .Z(out[1486]) );
  OR U3475 ( .A(n2271), .B(n2100), .Z(n2101) );
  XNOR U3476 ( .A(n2270), .B(n2101), .Z(out[1487]) );
  OR U3477 ( .A(n2276), .B(n2102), .Z(n2103) );
  XNOR U3478 ( .A(n2275), .B(n2103), .Z(out[1488]) );
  OR U3479 ( .A(n2280), .B(n2104), .Z(n2105) );
  XNOR U3480 ( .A(n2279), .B(n2105), .Z(out[1489]) );
  XNOR U3481 ( .A(in[685]), .B(n3938), .Z(n2664) );
  XOR U3482 ( .A(in[619]), .B(n3806), .Z(n4231) );
  XOR U3483 ( .A(in[210]), .B(n3617), .Z(n4229) );
  NAND U3484 ( .A(n4231), .B(n4229), .Z(n2106) );
  XNOR U3485 ( .A(n2664), .B(n2106), .Z(out[148]) );
  OR U3486 ( .A(n2284), .B(n2107), .Z(n2108) );
  XNOR U3487 ( .A(n2283), .B(n2108), .Z(out[1490]) );
  OR U3488 ( .A(n2288), .B(n2109), .Z(n2110) );
  XNOR U3489 ( .A(n2287), .B(n2110), .Z(out[1491]) );
  OR U3490 ( .A(n2292), .B(n2111), .Z(n2112) );
  XNOR U3491 ( .A(n2291), .B(n2112), .Z(out[1492]) );
  OR U3492 ( .A(n2296), .B(n2113), .Z(n2114) );
  XNOR U3493 ( .A(n2295), .B(n2114), .Z(out[1493]) );
  OR U3494 ( .A(n2300), .B(n2115), .Z(n2116) );
  XNOR U3495 ( .A(n2299), .B(n2116), .Z(out[1494]) );
  OR U3496 ( .A(n2304), .B(n2117), .Z(n2118) );
  XNOR U3497 ( .A(n2303), .B(n2118), .Z(out[1495]) );
  OR U3498 ( .A(n2309), .B(n2119), .Z(n2120) );
  XNOR U3499 ( .A(n2308), .B(n2120), .Z(out[1496]) );
  OR U3500 ( .A(n2313), .B(n2121), .Z(n2122) );
  XNOR U3501 ( .A(n2312), .B(n2122), .Z(out[1497]) );
  OR U3502 ( .A(n2317), .B(n2123), .Z(n2124) );
  XNOR U3503 ( .A(n2316), .B(n2124), .Z(out[1498]) );
  OR U3504 ( .A(n2321), .B(n2125), .Z(n2126) );
  XNOR U3505 ( .A(n2320), .B(n2126), .Z(out[1499]) );
  XNOR U3506 ( .A(in[686]), .B(n3940), .Z(n2666) );
  XOR U3507 ( .A(in[620]), .B(n3810), .Z(n4255) );
  XNOR U3508 ( .A(in[211]), .B(n3625), .Z(n4253) );
  NAND U3509 ( .A(n4255), .B(n4253), .Z(n2127) );
  XNOR U3510 ( .A(n2666), .B(n2127), .Z(out[149]) );
  XNOR U3511 ( .A(in[1424]), .B(n3634), .Z(n4038) );
  XOR U3512 ( .A(in[1047]), .B(n4132), .Z(n2645) );
  NAND U3513 ( .A(n4038), .B(n2645), .Z(n2128) );
  XNOR U3514 ( .A(n4039), .B(n2128), .Z(out[14]) );
  OR U3515 ( .A(n2325), .B(n2129), .Z(n2130) );
  XNOR U3516 ( .A(n2324), .B(n2130), .Z(out[1500]) );
  OR U3517 ( .A(n2329), .B(n2131), .Z(n2132) );
  XNOR U3518 ( .A(n2328), .B(n2132), .Z(out[1501]) );
  OR U3519 ( .A(n2333), .B(n2133), .Z(n2134) );
  XNOR U3520 ( .A(n2332), .B(n2134), .Z(out[1502]) );
  OR U3521 ( .A(n2337), .B(n2135), .Z(n2136) );
  XNOR U3522 ( .A(n2336), .B(n2136), .Z(out[1503]) );
  OR U3523 ( .A(n2342), .B(n2137), .Z(n2138) );
  XNOR U3524 ( .A(n2341), .B(n2138), .Z(out[1504]) );
  OR U3525 ( .A(n2346), .B(n2139), .Z(n2140) );
  XNOR U3526 ( .A(n2345), .B(n2140), .Z(out[1505]) );
  OR U3527 ( .A(n2351), .B(n2141), .Z(n2142) );
  XNOR U3528 ( .A(n2350), .B(n2142), .Z(out[1506]) );
  OR U3529 ( .A(n2355), .B(n2143), .Z(n2144) );
  XNOR U3530 ( .A(n2354), .B(n2144), .Z(out[1507]) );
  OR U3531 ( .A(n2359), .B(n2145), .Z(n2146) );
  XNOR U3532 ( .A(n2358), .B(n2146), .Z(out[1508]) );
  OR U3533 ( .A(n2363), .B(n2147), .Z(n2148) );
  XNOR U3534 ( .A(n2362), .B(n2148), .Z(out[1509]) );
  XNOR U3535 ( .A(in[687]), .B(n3942), .Z(n2669) );
  XOR U3536 ( .A(in[621]), .B(n3814), .Z(n4279) );
  XNOR U3537 ( .A(in[212]), .B(n3629), .Z(n4277) );
  NAND U3538 ( .A(n4279), .B(n4277), .Z(n2149) );
  XNOR U3539 ( .A(n2669), .B(n2149), .Z(out[150]) );
  OR U3540 ( .A(n2367), .B(n2150), .Z(n2151) );
  XNOR U3541 ( .A(n2366), .B(n2151), .Z(out[1510]) );
  OR U3542 ( .A(n2371), .B(n2152), .Z(n2153) );
  XNOR U3543 ( .A(n2370), .B(n2153), .Z(out[1511]) );
  OR U3544 ( .A(n2375), .B(n2154), .Z(n2155) );
  XNOR U3545 ( .A(n2374), .B(n2155), .Z(out[1512]) );
  OR U3546 ( .A(n2379), .B(n2156), .Z(n2157) );
  XNOR U3547 ( .A(n2378), .B(n2157), .Z(out[1513]) );
  OR U3548 ( .A(n2383), .B(n2158), .Z(n2159) );
  XNOR U3549 ( .A(n2382), .B(n2159), .Z(out[1514]) );
  OR U3550 ( .A(n2387), .B(n2160), .Z(n2161) );
  XNOR U3551 ( .A(n2386), .B(n2161), .Z(out[1515]) );
  OR U3552 ( .A(n2392), .B(n2162), .Z(n2163) );
  XNOR U3553 ( .A(n2391), .B(n2163), .Z(out[1516]) );
  OR U3554 ( .A(n2396), .B(n2164), .Z(n2165) );
  XNOR U3555 ( .A(n2395), .B(n2165), .Z(out[1517]) );
  OR U3556 ( .A(n2400), .B(n2166), .Z(n2167) );
  XNOR U3557 ( .A(n2399), .B(n2167), .Z(out[1518]) );
  OR U3558 ( .A(n2404), .B(n2168), .Z(n2169) );
  XNOR U3559 ( .A(n2403), .B(n2169), .Z(out[1519]) );
  XNOR U3560 ( .A(in[688]), .B(n3948), .Z(n2672) );
  XOR U3561 ( .A(in[622]), .B(n3536), .Z(n4303) );
  XNOR U3562 ( .A(in[213]), .B(n3633), .Z(n4301) );
  NAND U3563 ( .A(n4303), .B(n4301), .Z(n2170) );
  XNOR U3564 ( .A(n2672), .B(n2170), .Z(out[151]) );
  OR U3565 ( .A(n2408), .B(n2171), .Z(n2172) );
  XNOR U3566 ( .A(n2407), .B(n2172), .Z(out[1520]) );
  OR U3567 ( .A(n2412), .B(n2173), .Z(n2174) );
  XNOR U3568 ( .A(n2411), .B(n2174), .Z(out[1521]) );
  OR U3569 ( .A(n2416), .B(n2175), .Z(n2176) );
  XNOR U3570 ( .A(n2415), .B(n2176), .Z(out[1522]) );
  OR U3571 ( .A(n2420), .B(n2177), .Z(n2178) );
  XNOR U3572 ( .A(n2419), .B(n2178), .Z(out[1523]) );
  OR U3573 ( .A(n2424), .B(n2179), .Z(n2180) );
  XNOR U3574 ( .A(n2423), .B(n2180), .Z(out[1524]) );
  OR U3575 ( .A(n2428), .B(n2181), .Z(n2182) );
  XNOR U3576 ( .A(n2427), .B(n2182), .Z(out[1525]) );
  OR U3577 ( .A(n2433), .B(n2183), .Z(n2184) );
  XNOR U3578 ( .A(n2432), .B(n2184), .Z(out[1526]) );
  OR U3579 ( .A(n2437), .B(n2185), .Z(n2186) );
  XNOR U3580 ( .A(n2436), .B(n2186), .Z(out[1527]) );
  OR U3581 ( .A(n2441), .B(n2187), .Z(n2188) );
  XNOR U3582 ( .A(n2440), .B(n2188), .Z(out[1528]) );
  OR U3583 ( .A(n2445), .B(n2189), .Z(n2190) );
  XNOR U3584 ( .A(n2444), .B(n2190), .Z(out[1529]) );
  XNOR U3585 ( .A(in[689]), .B(n3950), .Z(n2676) );
  XOR U3586 ( .A(in[623]), .B(n3540), .Z(n4327) );
  XNOR U3587 ( .A(in[214]), .B(n3637), .Z(n4325) );
  NAND U3588 ( .A(n4327), .B(n4325), .Z(n2191) );
  XNOR U3589 ( .A(n2676), .B(n2191), .Z(out[152]) );
  OR U3590 ( .A(n2449), .B(n2192), .Z(n2193) );
  XNOR U3591 ( .A(n2448), .B(n2193), .Z(out[1530]) );
  OR U3592 ( .A(n2453), .B(n2194), .Z(n2195) );
  XNOR U3593 ( .A(n2452), .B(n2195), .Z(out[1531]) );
  OR U3594 ( .A(n2457), .B(n2196), .Z(n2197) );
  XNOR U3595 ( .A(n2456), .B(n2197), .Z(out[1532]) );
  OR U3596 ( .A(n2461), .B(n2198), .Z(n2199) );
  XNOR U3597 ( .A(n2460), .B(n2199), .Z(out[1533]) );
  OR U3598 ( .A(n2465), .B(n2200), .Z(n2201) );
  XNOR U3599 ( .A(n2464), .B(n2201), .Z(out[1534]) );
  OR U3600 ( .A(n2469), .B(n2202), .Z(n2203) );
  XNOR U3601 ( .A(n2468), .B(n2203), .Z(out[1535]) );
  ANDN U3602 ( .B(n2205), .A(n2204), .Z(n2208) );
  XOR U3603 ( .A(n2206), .B(round_const[0]), .Z(n2207) );
  XNOR U3604 ( .A(n2208), .B(n2207), .Z(out[1536]) );
  ANDN U3605 ( .B(n2210), .A(n2209), .Z(n2213) );
  XOR U3606 ( .A(n2211), .B(round_const[1]), .Z(n2212) );
  XNOR U3607 ( .A(n2213), .B(n2212), .Z(out[1537]) );
  ANDN U3608 ( .B(n2215), .A(n2214), .Z(n2216) );
  XNOR U3609 ( .A(n2217), .B(n2216), .Z(out[1538]) );
  ANDN U3610 ( .B(n2219), .A(n2218), .Z(n2222) );
  XOR U3611 ( .A(n2220), .B(round_const_3), .Z(n2221) );
  XNOR U3612 ( .A(n2222), .B(n2221), .Z(out[1539]) );
  XNOR U3613 ( .A(in[690]), .B(n3952), .Z(n2679) );
  XOR U3614 ( .A(in[624]), .B(n3544), .Z(n4359) );
  XNOR U3615 ( .A(in[215]), .B(n3641), .Z(n4357) );
  NAND U3616 ( .A(n4359), .B(n4357), .Z(n2223) );
  XNOR U3617 ( .A(n2679), .B(n2223), .Z(out[153]) );
  ANDN U3618 ( .B(n2225), .A(n2224), .Z(n2226) );
  XNOR U3619 ( .A(n2227), .B(n2226), .Z(out[1540]) );
  ANDN U3620 ( .B(n2229), .A(n2228), .Z(n2230) );
  XNOR U3621 ( .A(n2231), .B(n2230), .Z(out[1541]) );
  ANDN U3622 ( .B(n2233), .A(n2232), .Z(n2234) );
  XNOR U3623 ( .A(n2235), .B(n2234), .Z(out[1542]) );
  ANDN U3624 ( .B(n2237), .A(n2236), .Z(n2240) );
  XOR U3625 ( .A(n2238), .B(round_const_7), .Z(n2239) );
  XNOR U3626 ( .A(n2240), .B(n2239), .Z(out[1543]) );
  ANDN U3627 ( .B(n2242), .A(n2241), .Z(n2243) );
  XNOR U3628 ( .A(n2244), .B(n2243), .Z(out[1544]) );
  ANDN U3629 ( .B(n2246), .A(n2245), .Z(n2247) );
  XNOR U3630 ( .A(n2248), .B(n2247), .Z(out[1545]) );
  ANDN U3631 ( .B(n2250), .A(n2249), .Z(n2251) );
  XNOR U3632 ( .A(n2252), .B(n2251), .Z(out[1546]) );
  ANDN U3633 ( .B(n2254), .A(n2253), .Z(n2255) );
  XNOR U3634 ( .A(n2256), .B(n2255), .Z(out[1547]) );
  ANDN U3635 ( .B(n2258), .A(n2257), .Z(n2259) );
  XNOR U3636 ( .A(n2260), .B(n2259), .Z(out[1548]) );
  ANDN U3637 ( .B(n2262), .A(n2261), .Z(n2263) );
  XNOR U3638 ( .A(n2264), .B(n2263), .Z(out[1549]) );
  XNOR U3639 ( .A(in[691]), .B(n3954), .Z(n2682) );
  XOR U3640 ( .A(in[625]), .B(n3548), .Z(n4407) );
  XNOR U3641 ( .A(in[216]), .B(n3645), .Z(n4405) );
  NAND U3642 ( .A(n4407), .B(n4405), .Z(n2265) );
  XNOR U3643 ( .A(n2682), .B(n2265), .Z(out[154]) );
  ANDN U3644 ( .B(n2267), .A(n2266), .Z(n2268) );
  XNOR U3645 ( .A(n2269), .B(n2268), .Z(out[1550]) );
  ANDN U3646 ( .B(n2271), .A(n2270), .Z(n2274) );
  XOR U3647 ( .A(n2272), .B(round_const_15), .Z(n2273) );
  XNOR U3648 ( .A(n2274), .B(n2273), .Z(out[1551]) );
  ANDN U3649 ( .B(n2276), .A(n2275), .Z(n2277) );
  XNOR U3650 ( .A(n2278), .B(n2277), .Z(out[1552]) );
  ANDN U3651 ( .B(n2280), .A(n2279), .Z(n2281) );
  XNOR U3652 ( .A(n2282), .B(n2281), .Z(out[1553]) );
  ANDN U3653 ( .B(n2284), .A(n2283), .Z(n2285) );
  XNOR U3654 ( .A(n2286), .B(n2285), .Z(out[1554]) );
  ANDN U3655 ( .B(n2288), .A(n2287), .Z(n2289) );
  XNOR U3656 ( .A(n2290), .B(n2289), .Z(out[1555]) );
  ANDN U3657 ( .B(n2292), .A(n2291), .Z(n2293) );
  XNOR U3658 ( .A(n2294), .B(n2293), .Z(out[1556]) );
  ANDN U3659 ( .B(n2296), .A(n2295), .Z(n2297) );
  XNOR U3660 ( .A(n2298), .B(n2297), .Z(out[1557]) );
  ANDN U3661 ( .B(n2300), .A(n2299), .Z(n2301) );
  XNOR U3662 ( .A(n2302), .B(n2301), .Z(out[1558]) );
  ANDN U3663 ( .B(n2304), .A(n2303), .Z(n2305) );
  XNOR U3664 ( .A(n2306), .B(n2305), .Z(out[1559]) );
  XNOR U3665 ( .A(in[692]), .B(n3956), .Z(n2685) );
  XOR U3666 ( .A(in[626]), .B(n3552), .Z(n4451) );
  XNOR U3667 ( .A(in[217]), .B(n3649), .Z(n4449) );
  NAND U3668 ( .A(n4451), .B(n4449), .Z(n2307) );
  XNOR U3669 ( .A(n2685), .B(n2307), .Z(out[155]) );
  ANDN U3670 ( .B(n2309), .A(n2308), .Z(n2310) );
  XNOR U3671 ( .A(n2311), .B(n2310), .Z(out[1560]) );
  ANDN U3672 ( .B(n2313), .A(n2312), .Z(n2314) );
  XNOR U3673 ( .A(n2315), .B(n2314), .Z(out[1561]) );
  ANDN U3674 ( .B(n2317), .A(n2316), .Z(n2318) );
  XNOR U3675 ( .A(n2319), .B(n2318), .Z(out[1562]) );
  ANDN U3676 ( .B(n2321), .A(n2320), .Z(n2322) );
  XNOR U3677 ( .A(n2323), .B(n2322), .Z(out[1563]) );
  ANDN U3678 ( .B(n2325), .A(n2324), .Z(n2326) );
  XNOR U3679 ( .A(n2327), .B(n2326), .Z(out[1564]) );
  ANDN U3680 ( .B(n2329), .A(n2328), .Z(n2330) );
  XNOR U3681 ( .A(n2331), .B(n2330), .Z(out[1565]) );
  ANDN U3682 ( .B(n2333), .A(n2332), .Z(n2334) );
  XNOR U3683 ( .A(n2335), .B(n2334), .Z(out[1566]) );
  ANDN U3684 ( .B(n2337), .A(n2336), .Z(n2340) );
  XOR U3685 ( .A(n2338), .B(round_const_31), .Z(n2339) );
  XNOR U3686 ( .A(n2340), .B(n2339), .Z(out[1567]) );
  ANDN U3687 ( .B(n2342), .A(n2341), .Z(n2343) );
  XNOR U3688 ( .A(n2344), .B(n2343), .Z(out[1568]) );
  ANDN U3689 ( .B(n2346), .A(n2345), .Z(n2347) );
  XNOR U3690 ( .A(n2348), .B(n2347), .Z(out[1569]) );
  XNOR U3691 ( .A(in[693]), .B(n3958), .Z(n2688) );
  XOR U3692 ( .A(in[627]), .B(n3556), .Z(n4495) );
  XNOR U3693 ( .A(in[218]), .B(n3653), .Z(n4492) );
  NAND U3694 ( .A(n4495), .B(n4492), .Z(n2349) );
  XNOR U3695 ( .A(n2688), .B(n2349), .Z(out[156]) );
  ANDN U3696 ( .B(n2351), .A(n2350), .Z(n2352) );
  XNOR U3697 ( .A(n2353), .B(n2352), .Z(out[1570]) );
  ANDN U3698 ( .B(n2355), .A(n2354), .Z(n2356) );
  XNOR U3699 ( .A(n2357), .B(n2356), .Z(out[1571]) );
  ANDN U3700 ( .B(n2359), .A(n2358), .Z(n2360) );
  XNOR U3701 ( .A(n2361), .B(n2360), .Z(out[1572]) );
  ANDN U3702 ( .B(n2363), .A(n2362), .Z(n2364) );
  XNOR U3703 ( .A(n2365), .B(n2364), .Z(out[1573]) );
  ANDN U3704 ( .B(n2367), .A(n2366), .Z(n2368) );
  XNOR U3705 ( .A(n2369), .B(n2368), .Z(out[1574]) );
  ANDN U3706 ( .B(n2371), .A(n2370), .Z(n2372) );
  XNOR U3707 ( .A(n2373), .B(n2372), .Z(out[1575]) );
  ANDN U3708 ( .B(n2375), .A(n2374), .Z(n2376) );
  XNOR U3709 ( .A(n2377), .B(n2376), .Z(out[1576]) );
  ANDN U3710 ( .B(n2379), .A(n2378), .Z(n2380) );
  XNOR U3711 ( .A(n2381), .B(n2380), .Z(out[1577]) );
  ANDN U3712 ( .B(n2383), .A(n2382), .Z(n2384) );
  XNOR U3713 ( .A(n2385), .B(n2384), .Z(out[1578]) );
  ANDN U3714 ( .B(n2387), .A(n2386), .Z(n2388) );
  XNOR U3715 ( .A(n2389), .B(n2388), .Z(out[1579]) );
  XNOR U3716 ( .A(in[694]), .B(n3960), .Z(n2690) );
  XOR U3717 ( .A(in[628]), .B(n3560), .Z(n4539) );
  XNOR U3718 ( .A(in[219]), .B(n3657), .Z(n4536) );
  NAND U3719 ( .A(n4539), .B(n4536), .Z(n2390) );
  XNOR U3720 ( .A(n2690), .B(n2390), .Z(out[157]) );
  ANDN U3721 ( .B(n2392), .A(n2391), .Z(n2393) );
  XNOR U3722 ( .A(n2394), .B(n2393), .Z(out[1580]) );
  ANDN U3723 ( .B(n2396), .A(n2395), .Z(n2397) );
  XNOR U3724 ( .A(n2398), .B(n2397), .Z(out[1581]) );
  ANDN U3725 ( .B(n2400), .A(n2399), .Z(n2401) );
  XNOR U3726 ( .A(n2402), .B(n2401), .Z(out[1582]) );
  ANDN U3727 ( .B(n2404), .A(n2403), .Z(n2405) );
  XNOR U3728 ( .A(n2406), .B(n2405), .Z(out[1583]) );
  ANDN U3729 ( .B(n2408), .A(n2407), .Z(n2409) );
  XNOR U3730 ( .A(n2410), .B(n2409), .Z(out[1584]) );
  ANDN U3731 ( .B(n2412), .A(n2411), .Z(n2413) );
  XNOR U3732 ( .A(n2414), .B(n2413), .Z(out[1585]) );
  ANDN U3733 ( .B(n2416), .A(n2415), .Z(n2417) );
  XNOR U3734 ( .A(n2418), .B(n2417), .Z(out[1586]) );
  ANDN U3735 ( .B(n2420), .A(n2419), .Z(n2421) );
  XNOR U3736 ( .A(n2422), .B(n2421), .Z(out[1587]) );
  ANDN U3737 ( .B(n2424), .A(n2423), .Z(n2425) );
  XNOR U3738 ( .A(n2426), .B(n2425), .Z(out[1588]) );
  ANDN U3739 ( .B(n2428), .A(n2427), .Z(n2429) );
  XNOR U3740 ( .A(n2430), .B(n2429), .Z(out[1589]) );
  XNOR U3741 ( .A(in[695]), .B(n3962), .Z(n2692) );
  XOR U3742 ( .A(in[629]), .B(n3564), .Z(n4583) );
  XNOR U3743 ( .A(in[220]), .B(n3661), .Z(n4580) );
  NAND U3744 ( .A(n4583), .B(n4580), .Z(n2431) );
  XNOR U3745 ( .A(n2692), .B(n2431), .Z(out[158]) );
  ANDN U3746 ( .B(n2433), .A(n2432), .Z(n2434) );
  XNOR U3747 ( .A(n2435), .B(n2434), .Z(out[1590]) );
  ANDN U3748 ( .B(n2437), .A(n2436), .Z(n2438) );
  XNOR U3749 ( .A(n2439), .B(n2438), .Z(out[1591]) );
  ANDN U3750 ( .B(n2441), .A(n2440), .Z(n2442) );
  XNOR U3751 ( .A(n2443), .B(n2442), .Z(out[1592]) );
  ANDN U3752 ( .B(n2445), .A(n2444), .Z(n2446) );
  XNOR U3753 ( .A(n2447), .B(n2446), .Z(out[1593]) );
  ANDN U3754 ( .B(n2449), .A(n2448), .Z(n2450) );
  XNOR U3755 ( .A(n2451), .B(n2450), .Z(out[1594]) );
  ANDN U3756 ( .B(n2453), .A(n2452), .Z(n2454) );
  XNOR U3757 ( .A(n2455), .B(n2454), .Z(out[1595]) );
  ANDN U3758 ( .B(n2457), .A(n2456), .Z(n2458) );
  XNOR U3759 ( .A(n2459), .B(n2458), .Z(out[1596]) );
  ANDN U3760 ( .B(n2461), .A(n2460), .Z(n2462) );
  XNOR U3761 ( .A(n2463), .B(n2462), .Z(out[1597]) );
  ANDN U3762 ( .B(n2465), .A(n2464), .Z(n2466) );
  XNOR U3763 ( .A(n2467), .B(n2466), .Z(out[1598]) );
  ANDN U3764 ( .B(n2469), .A(n2468), .Z(n2472) );
  XOR U3765 ( .A(n2470), .B(round_const_63), .Z(n2471) );
  XNOR U3766 ( .A(n2472), .B(n2471), .Z(out[1599]) );
  XNOR U3767 ( .A(in[696]), .B(n3818), .Z(n2694) );
  XOR U3768 ( .A(in[630]), .B(n3568), .Z(n4627) );
  XNOR U3769 ( .A(in[221]), .B(n3669), .Z(n4624) );
  NAND U3770 ( .A(n4627), .B(n4624), .Z(n2473) );
  XNOR U3771 ( .A(n2694), .B(n2473), .Z(out[159]) );
  XNOR U3772 ( .A(in[1425]), .B(n3638), .Z(n4072) );
  XOR U3773 ( .A(in[1048]), .B(n4135), .Z(n2648) );
  NAND U3774 ( .A(n4072), .B(n2648), .Z(n2474) );
  XNOR U3775 ( .A(n4073), .B(n2474), .Z(out[15]) );
  XNOR U3776 ( .A(in[697]), .B(n3820), .Z(n2696) );
  XOR U3777 ( .A(in[631]), .B(n3572), .Z(n4671) );
  XNOR U3778 ( .A(in[222]), .B(n3673), .Z(n4668) );
  NAND U3779 ( .A(n4671), .B(n4668), .Z(n2475) );
  XNOR U3780 ( .A(n2696), .B(n2475), .Z(out[160]) );
  XNOR U3781 ( .A(in[698]), .B(n3822), .Z(n2698) );
  XOR U3782 ( .A(in[632]), .B(n3580), .Z(n4715) );
  XNOR U3783 ( .A(in[223]), .B(n3677), .Z(n4712) );
  NAND U3784 ( .A(n4715), .B(n4712), .Z(n2476) );
  XNOR U3785 ( .A(n2698), .B(n2476), .Z(out[161]) );
  XNOR U3786 ( .A(in[699]), .B(n3824), .Z(n2702) );
  XOR U3787 ( .A(in[633]), .B(n3584), .Z(n4759) );
  XNOR U3788 ( .A(in[224]), .B(n3681), .Z(n4756) );
  NAND U3789 ( .A(n4759), .B(n4756), .Z(n2477) );
  XNOR U3790 ( .A(n2702), .B(n2477), .Z(out[162]) );
  XNOR U3791 ( .A(in[700]), .B(n3826), .Z(n2704) );
  XOR U3792 ( .A(in[634]), .B(n3588), .Z(n4803) );
  XNOR U3793 ( .A(in[225]), .B(n3685), .Z(n4800) );
  NAND U3794 ( .A(n4803), .B(n4800), .Z(n2478) );
  XNOR U3795 ( .A(n2704), .B(n2478), .Z(out[163]) );
  XOR U3796 ( .A(in[701]), .B(n3828), .Z(n2706) );
  NOR U3797 ( .A(n2550), .B(n2831), .Z(n2479) );
  XNOR U3798 ( .A(n2706), .B(n2479), .Z(out[164]) );
  XOR U3799 ( .A(in[702]), .B(n3834), .Z(n2708) );
  NOR U3800 ( .A(n2552), .B(n2845), .Z(n2480) );
  XNOR U3801 ( .A(n2708), .B(n2480), .Z(out[165]) );
  XOR U3802 ( .A(in[703]), .B(n3836), .Z(n2710) );
  NOR U3803 ( .A(n2555), .B(n2859), .Z(n2481) );
  XNOR U3804 ( .A(n2710), .B(n2481), .Z(out[166]) );
  XOR U3805 ( .A(in[640]), .B(n3838), .Z(n2712) );
  NOR U3806 ( .A(n2557), .B(n2873), .Z(n2482) );
  XNOR U3807 ( .A(n2712), .B(n2482), .Z(out[167]) );
  XOR U3808 ( .A(in[641]), .B(n3840), .Z(n2714) );
  NOR U3809 ( .A(n2559), .B(n2889), .Z(n2483) );
  XNOR U3810 ( .A(n2714), .B(n2483), .Z(out[168]) );
  XOR U3811 ( .A(in[642]), .B(n3842), .Z(n2716) );
  NOR U3812 ( .A(n2561), .B(n2903), .Z(n2484) );
  XNOR U3813 ( .A(n2716), .B(n2484), .Z(out[169]) );
  XNOR U3814 ( .A(in[1426]), .B(n3642), .Z(n4110) );
  XOR U3815 ( .A(in[1049]), .B(n4138), .Z(n2651) );
  NAND U3816 ( .A(n4110), .B(n2651), .Z(n2485) );
  XNOR U3817 ( .A(n4111), .B(n2485), .Z(out[16]) );
  XOR U3818 ( .A(in[643]), .B(n3844), .Z(n2718) );
  NOR U3819 ( .A(n2563), .B(n2917), .Z(n2486) );
  XNOR U3820 ( .A(n2718), .B(n2486), .Z(out[170]) );
  XOR U3821 ( .A(in[644]), .B(n3846), .Z(n2720) );
  NOR U3822 ( .A(n2565), .B(n2931), .Z(n2487) );
  XNOR U3823 ( .A(n2720), .B(n2487), .Z(out[171]) );
  XOR U3824 ( .A(in[645]), .B(n3848), .Z(n2726) );
  NOR U3825 ( .A(n2567), .B(n2947), .Z(n2488) );
  XNOR U3826 ( .A(n2726), .B(n2488), .Z(out[172]) );
  XOR U3827 ( .A(in[646]), .B(n3850), .Z(n2728) );
  NOR U3828 ( .A(n2569), .B(n2971), .Z(n2489) );
  XNOR U3829 ( .A(n2728), .B(n2489), .Z(out[173]) );
  XOR U3830 ( .A(in[647]), .B(n3852), .Z(n2730) );
  NOR U3831 ( .A(n2571), .B(n2995), .Z(n2490) );
  XNOR U3832 ( .A(n2730), .B(n2490), .Z(out[174]) );
  XOR U3833 ( .A(in[648]), .B(n3856), .Z(n2732) );
  NOR U3834 ( .A(n2573), .B(n3019), .Z(n2491) );
  XNOR U3835 ( .A(n2732), .B(n2491), .Z(out[175]) );
  XOR U3836 ( .A(in[649]), .B(n3858), .Z(n2734) );
  NOR U3837 ( .A(n2576), .B(n3043), .Z(n2492) );
  XNOR U3838 ( .A(n2734), .B(n2492), .Z(out[176]) );
  XOR U3839 ( .A(in[650]), .B(n3860), .Z(n2736) );
  NOR U3840 ( .A(n2578), .B(n3067), .Z(n2493) );
  XNOR U3841 ( .A(n2736), .B(n2493), .Z(out[177]) );
  XOR U3842 ( .A(in[651]), .B(n3862), .Z(n2738) );
  NOR U3843 ( .A(n2580), .B(n3093), .Z(n2494) );
  XNOR U3844 ( .A(n2738), .B(n2494), .Z(out[178]) );
  XOR U3845 ( .A(in[652]), .B(n3864), .Z(n2740) );
  NOR U3846 ( .A(n2582), .B(n3117), .Z(n2495) );
  XNOR U3847 ( .A(n2740), .B(n2495), .Z(out[179]) );
  XNOR U3848 ( .A(in[1427]), .B(n3646), .Z(n4144) );
  XOR U3849 ( .A(in[1050]), .B(n4141), .Z(n2654) );
  NAND U3850 ( .A(n4144), .B(n2654), .Z(n2496) );
  XNOR U3851 ( .A(n4145), .B(n2496), .Z(out[17]) );
  XOR U3852 ( .A(in[653]), .B(n3866), .Z(n2742) );
  NOR U3853 ( .A(n2584), .B(n3141), .Z(n2497) );
  XNOR U3854 ( .A(n2742), .B(n2497), .Z(out[180]) );
  XOR U3855 ( .A(in[654]), .B(n3868), .Z(n2744) );
  NOR U3856 ( .A(n2586), .B(n3165), .Z(n2498) );
  XNOR U3857 ( .A(n2744), .B(n2498), .Z(out[181]) );
  XOR U3858 ( .A(in[655]), .B(n3870), .Z(n2748) );
  NOR U3859 ( .A(n2588), .B(n3189), .Z(n2499) );
  XNOR U3860 ( .A(n2748), .B(n2499), .Z(out[182]) );
  XOR U3861 ( .A(in[656]), .B(n3872), .Z(n2750) );
  NOR U3862 ( .A(n2590), .B(n3213), .Z(n2500) );
  XNOR U3863 ( .A(n2750), .B(n2500), .Z(out[183]) );
  XOR U3864 ( .A(in[657]), .B(n3874), .Z(n2752) );
  NOR U3865 ( .A(n2592), .B(n3237), .Z(n2501) );
  XNOR U3866 ( .A(n2752), .B(n2501), .Z(out[184]) );
  XOR U3867 ( .A(in[658]), .B(n3878), .Z(n2754) );
  NOR U3868 ( .A(n2594), .B(n3269), .Z(n2502) );
  XNOR U3869 ( .A(n2754), .B(n2502), .Z(out[185]) );
  XOR U3870 ( .A(in[659]), .B(n3880), .Z(n2756) );
  NOR U3871 ( .A(n2597), .B(n3313), .Z(n2503) );
  XNOR U3872 ( .A(n2756), .B(n2503), .Z(out[186]) );
  XOR U3873 ( .A(in[660]), .B(n3882), .Z(n2758) );
  NOR U3874 ( .A(n2599), .B(n3357), .Z(n2504) );
  XNOR U3875 ( .A(n2758), .B(n2504), .Z(out[187]) );
  XOR U3876 ( .A(in[661]), .B(n3884), .Z(n2760) );
  NOR U3877 ( .A(n2601), .B(n3403), .Z(n2505) );
  XNOR U3878 ( .A(n2760), .B(n2505), .Z(out[188]) );
  XOR U3879 ( .A(in[662]), .B(n3886), .Z(n2762) );
  NOR U3880 ( .A(n2603), .B(n3447), .Z(n2506) );
  XNOR U3881 ( .A(n2762), .B(n2506), .Z(out[189]) );
  XNOR U3882 ( .A(in[1428]), .B(n3650), .Z(n4178) );
  XOR U3883 ( .A(in[1051]), .B(n4148), .Z(n2657) );
  NAND U3884 ( .A(n4178), .B(n2657), .Z(n2507) );
  XNOR U3885 ( .A(n4179), .B(n2507), .Z(out[18]) );
  XOR U3886 ( .A(in[663]), .B(n3888), .Z(n2764) );
  NOR U3887 ( .A(n2605), .B(n3491), .Z(n2508) );
  XNOR U3888 ( .A(n2764), .B(n2508), .Z(out[190]) );
  XOR U3889 ( .A(in[664]), .B(n3890), .Z(n2766) );
  NOR U3890 ( .A(n2607), .B(n3535), .Z(n2509) );
  XNOR U3891 ( .A(n2766), .B(n2509), .Z(out[191]) );
  OR U3892 ( .A(n2610), .B(n3579), .Z(n2510) );
  XNOR U3893 ( .A(n2609), .B(n2510), .Z(out[192]) );
  XOR U3894 ( .A(in[1034]), .B(n4089), .Z(n2613) );
  NOR U3895 ( .A(n2612), .B(n3623), .Z(n2511) );
  XNOR U3896 ( .A(n2613), .B(n2511), .Z(out[193]) );
  XOR U3897 ( .A(in[1035]), .B(n4092), .Z(n2724) );
  NOR U3898 ( .A(n2615), .B(n3667), .Z(n2512) );
  XNOR U3899 ( .A(n2724), .B(n2512), .Z(out[194]) );
  XNOR U3900 ( .A(n4095), .B(in[1036]), .Z(n2874) );
  NOR U3901 ( .A(n2617), .B(n3711), .Z(n2513) );
  XNOR U3902 ( .A(n2874), .B(n2513), .Z(out[195]) );
  XNOR U3903 ( .A(n4098), .B(in[1037]), .Z(n3068) );
  NOR U3904 ( .A(n2620), .B(n3755), .Z(n2514) );
  XNOR U3905 ( .A(n3068), .B(n2514), .Z(out[196]) );
  XNOR U3906 ( .A(n4101), .B(in[1038]), .Z(n3358) );
  NOR U3907 ( .A(n2622), .B(n3799), .Z(n2515) );
  XNOR U3908 ( .A(n3358), .B(n2515), .Z(out[197]) );
  XNOR U3909 ( .A(n4104), .B(in[1039]), .Z(n3800) );
  NOR U3910 ( .A(n2624), .B(n3833), .Z(n2516) );
  XNOR U3911 ( .A(n3800), .B(n2516), .Z(out[198]) );
  XNOR U3912 ( .A(n4107), .B(in[1040]), .Z(n4076) );
  NOR U3913 ( .A(n2626), .B(n3855), .Z(n2517) );
  XNOR U3914 ( .A(n4076), .B(n2517), .Z(out[199]) );
  XNOR U3915 ( .A(in[1429]), .B(n3654), .Z(n4204) );
  XOR U3916 ( .A(in[1052]), .B(n4151), .Z(n2660) );
  NAND U3917 ( .A(n4204), .B(n2660), .Z(n2518) );
  XNOR U3918 ( .A(n4205), .B(n2518), .Z(out[19]) );
  XNOR U3919 ( .A(n3574), .B(in[1411]), .Z(n3620) );
  NANDN U3920 ( .A(n2613), .B(n3620), .Z(n2519) );
  XNOR U3921 ( .A(n3621), .B(n2519), .Z(out[1]) );
  XNOR U3922 ( .A(n4114), .B(in[1041]), .Z(n4360) );
  NOR U3923 ( .A(n2628), .B(n3877), .Z(n2520) );
  XNOR U3924 ( .A(n4360), .B(n2520), .Z(out[200]) );
  XNOR U3925 ( .A(n4117), .B(in[1042]), .Z(n4804) );
  NOR U3926 ( .A(n2630), .B(n3899), .Z(n2521) );
  XNOR U3927 ( .A(n4804), .B(n2521), .Z(out[201]) );
  OR U3928 ( .A(n2633), .B(n3923), .Z(n2522) );
  XNOR U3929 ( .A(n2632), .B(n2522), .Z(out[202]) );
  OR U3930 ( .A(n2636), .B(n3947), .Z(n2523) );
  XNOR U3931 ( .A(n2635), .B(n2523), .Z(out[203]) );
  OR U3932 ( .A(n2639), .B(n3973), .Z(n2524) );
  XNOR U3933 ( .A(n2638), .B(n2524), .Z(out[204]) );
  OR U3934 ( .A(n2642), .B(n4007), .Z(n2525) );
  XNOR U3935 ( .A(n2641), .B(n2525), .Z(out[205]) );
  OR U3936 ( .A(n2646), .B(n4041), .Z(n2526) );
  XNOR U3937 ( .A(n2645), .B(n2526), .Z(out[206]) );
  OR U3938 ( .A(n2649), .B(n4075), .Z(n2527) );
  XNOR U3939 ( .A(n2648), .B(n2527), .Z(out[207]) );
  OR U3940 ( .A(n2652), .B(n4113), .Z(n2528) );
  XNOR U3941 ( .A(n2651), .B(n2528), .Z(out[208]) );
  OR U3942 ( .A(n2655), .B(n4147), .Z(n2529) );
  XNOR U3943 ( .A(n2654), .B(n2529), .Z(out[209]) );
  XNOR U3944 ( .A(in[1430]), .B(n3658), .Z(n4228) );
  XOR U3945 ( .A(in[1053]), .B(n4154), .Z(n2663) );
  NAND U3946 ( .A(n4228), .B(n2663), .Z(n2530) );
  XNOR U3947 ( .A(n4229), .B(n2530), .Z(out[20]) );
  OR U3948 ( .A(n2658), .B(n4181), .Z(n2531) );
  XNOR U3949 ( .A(n2657), .B(n2531), .Z(out[210]) );
  OR U3950 ( .A(n2661), .B(n4207), .Z(n2532) );
  XNOR U3951 ( .A(n2660), .B(n2532), .Z(out[211]) );
  OR U3952 ( .A(n2664), .B(n4231), .Z(n2533) );
  XNOR U3953 ( .A(n2663), .B(n2533), .Z(out[212]) );
  XNOR U3954 ( .A(in[1054]), .B(n4157), .Z(n2667) );
  NOR U3955 ( .A(n2666), .B(n4255), .Z(n2534) );
  XNOR U3956 ( .A(n2667), .B(n2534), .Z(out[213]) );
  XNOR U3957 ( .A(in[1055]), .B(n4160), .Z(n2670) );
  NOR U3958 ( .A(n2669), .B(n4279), .Z(n2535) );
  XNOR U3959 ( .A(n2670), .B(n2535), .Z(out[214]) );
  XNOR U3960 ( .A(in[1056]), .B(n4163), .Z(n2673) );
  NOR U3961 ( .A(n2672), .B(n4303), .Z(n2536) );
  XNOR U3962 ( .A(n2673), .B(n2536), .Z(out[215]) );
  XNOR U3963 ( .A(in[1057]), .B(n4166), .Z(n2677) );
  NOR U3964 ( .A(n2676), .B(n4327), .Z(n2537) );
  XNOR U3965 ( .A(n2677), .B(n2537), .Z(out[216]) );
  XNOR U3966 ( .A(in[1058]), .B(n4169), .Z(n2680) );
  NOR U3967 ( .A(n2679), .B(n4359), .Z(n2538) );
  XNOR U3968 ( .A(n2680), .B(n2538), .Z(out[217]) );
  XNOR U3969 ( .A(in[1059]), .B(n4172), .Z(n2683) );
  NOR U3970 ( .A(n2682), .B(n4407), .Z(n2539) );
  XNOR U3971 ( .A(n2683), .B(n2539), .Z(out[218]) );
  XOR U3972 ( .A(in[1060]), .B(n4175), .Z(n2686) );
  NOR U3973 ( .A(n2685), .B(n4451), .Z(n2540) );
  XNOR U3974 ( .A(n2686), .B(n2540), .Z(out[219]) );
  XNOR U3975 ( .A(in[1431]), .B(n3662), .Z(n4252) );
  NANDN U3976 ( .A(n2667), .B(n4252), .Z(n2541) );
  XNOR U3977 ( .A(n4253), .B(n2541), .Z(out[21]) );
  XOR U3978 ( .A(in[1061]), .B(n4182), .Z(n2700) );
  NOR U3979 ( .A(n2688), .B(n4495), .Z(n2542) );
  XNOR U3980 ( .A(n2700), .B(n2542), .Z(out[220]) );
  XOR U3981 ( .A(in[1062]), .B(n4185), .Z(n2722) );
  NOR U3982 ( .A(n2690), .B(n4539), .Z(n2543) );
  XNOR U3983 ( .A(n2722), .B(n2543), .Z(out[221]) );
  XOR U3984 ( .A(in[1063]), .B(n3964), .Z(n2746) );
  NOR U3985 ( .A(n2692), .B(n4583), .Z(n2544) );
  XNOR U3986 ( .A(n2746), .B(n2544), .Z(out[222]) );
  XOR U3987 ( .A(in[1064]), .B(n3967), .Z(n2768) );
  NOR U3988 ( .A(n2694), .B(n4627), .Z(n2545) );
  XNOR U3989 ( .A(n2768), .B(n2545), .Z(out[223]) );
  XOR U3990 ( .A(in[1065]), .B(n3974), .Z(n2780) );
  NOR U3991 ( .A(n2696), .B(n4671), .Z(n2546) );
  XNOR U3992 ( .A(n2780), .B(n2546), .Z(out[224]) );
  XOR U3993 ( .A(in[1066]), .B(n3977), .Z(n2792) );
  NOR U3994 ( .A(n2698), .B(n4715), .Z(n2547) );
  XNOR U3995 ( .A(n2792), .B(n2547), .Z(out[225]) );
  XOR U3996 ( .A(in[1067]), .B(n3980), .Z(n2804) );
  NOR U3997 ( .A(n2702), .B(n4759), .Z(n2548) );
  XNOR U3998 ( .A(n2804), .B(n2548), .Z(out[226]) );
  XOR U3999 ( .A(in[1068]), .B(n3983), .Z(n2816) );
  NOR U4000 ( .A(n2704), .B(n4803), .Z(n2549) );
  XNOR U4001 ( .A(n2816), .B(n2549), .Z(out[227]) );
  XNOR U4002 ( .A(in[1069]), .B(n3986), .Z(n2829) );
  NAND U4003 ( .A(n2706), .B(n2550), .Z(n2551) );
  XNOR U4004 ( .A(n2829), .B(n2551), .Z(out[228]) );
  XNOR U4005 ( .A(in[1070]), .B(n3989), .Z(n2843) );
  NAND U4006 ( .A(n2708), .B(n2552), .Z(n2553) );
  XNOR U4007 ( .A(n2843), .B(n2553), .Z(out[229]) );
  XNOR U4008 ( .A(in[1432]), .B(n3670), .Z(n4276) );
  NANDN U4009 ( .A(n2670), .B(n4276), .Z(n2554) );
  XNOR U4010 ( .A(n4277), .B(n2554), .Z(out[22]) );
  XNOR U4011 ( .A(in[1071]), .B(n3992), .Z(n2857) );
  NAND U4012 ( .A(n2710), .B(n2555), .Z(n2556) );
  XNOR U4013 ( .A(n2857), .B(n2556), .Z(out[230]) );
  XNOR U4014 ( .A(in[1072]), .B(n3995), .Z(n2871) );
  NAND U4015 ( .A(n2712), .B(n2557), .Z(n2558) );
  XNOR U4016 ( .A(n2871), .B(n2558), .Z(out[231]) );
  XNOR U4017 ( .A(in[1073]), .B(n3998), .Z(n2887) );
  NAND U4018 ( .A(n2714), .B(n2559), .Z(n2560) );
  XNOR U4019 ( .A(n2887), .B(n2560), .Z(out[232]) );
  XNOR U4020 ( .A(in[1074]), .B(n4001), .Z(n2901) );
  NAND U4021 ( .A(n2716), .B(n2561), .Z(n2562) );
  XNOR U4022 ( .A(n2901), .B(n2562), .Z(out[233]) );
  XNOR U4023 ( .A(in[1075]), .B(n4008), .Z(n2915) );
  NAND U4024 ( .A(n2718), .B(n2563), .Z(n2564) );
  XNOR U4025 ( .A(n2915), .B(n2564), .Z(out[234]) );
  XNOR U4026 ( .A(in[1076]), .B(n4011), .Z(n2929) );
  NAND U4027 ( .A(n2720), .B(n2565), .Z(n2566) );
  XNOR U4028 ( .A(n2929), .B(n2566), .Z(out[235]) );
  XNOR U4029 ( .A(in[1077]), .B(n4014), .Z(n2945) );
  NAND U4030 ( .A(n2726), .B(n2567), .Z(n2568) );
  XNOR U4031 ( .A(n2945), .B(n2568), .Z(out[236]) );
  XNOR U4032 ( .A(in[1078]), .B(n4017), .Z(n2969) );
  NAND U4033 ( .A(n2728), .B(n2569), .Z(n2570) );
  XNOR U4034 ( .A(n2969), .B(n2570), .Z(out[237]) );
  XNOR U4035 ( .A(in[1079]), .B(n4020), .Z(n2993) );
  NAND U4036 ( .A(n2730), .B(n2571), .Z(n2572) );
  XNOR U4037 ( .A(n2993), .B(n2572), .Z(out[238]) );
  XNOR U4038 ( .A(in[1080]), .B(n4023), .Z(n3017) );
  NAND U4039 ( .A(n2732), .B(n2573), .Z(n2574) );
  XNOR U4040 ( .A(n3017), .B(n2574), .Z(out[239]) );
  XNOR U4041 ( .A(in[1433]), .B(n3674), .Z(n4300) );
  NANDN U4042 ( .A(n2673), .B(n4300), .Z(n2575) );
  XNOR U4043 ( .A(n4301), .B(n2575), .Z(out[23]) );
  XNOR U4044 ( .A(in[1081]), .B(n4026), .Z(n3041) );
  NAND U4045 ( .A(n2734), .B(n2576), .Z(n2577) );
  XNOR U4046 ( .A(n3041), .B(n2577), .Z(out[240]) );
  XNOR U4047 ( .A(in[1082]), .B(n4029), .Z(n3065) );
  NAND U4048 ( .A(n2736), .B(n2578), .Z(n2579) );
  XNOR U4049 ( .A(n3065), .B(n2579), .Z(out[241]) );
  XNOR U4050 ( .A(in[1083]), .B(n4032), .Z(n3091) );
  NAND U4051 ( .A(n2738), .B(n2580), .Z(n2581) );
  XNOR U4052 ( .A(n3091), .B(n2581), .Z(out[242]) );
  XNOR U4053 ( .A(in[1084]), .B(n4035), .Z(n3115) );
  NAND U4054 ( .A(n2740), .B(n2582), .Z(n2583) );
  XNOR U4055 ( .A(n3115), .B(n2583), .Z(out[243]) );
  XNOR U4056 ( .A(in[1085]), .B(n4042), .Z(n3139) );
  NAND U4057 ( .A(n2742), .B(n2584), .Z(n2585) );
  XNOR U4058 ( .A(n3139), .B(n2585), .Z(out[244]) );
  XNOR U4059 ( .A(in[1086]), .B(n4045), .Z(n3163) );
  NAND U4060 ( .A(n2744), .B(n2586), .Z(n2587) );
  XNOR U4061 ( .A(n3163), .B(n2587), .Z(out[245]) );
  XNOR U4062 ( .A(in[1087]), .B(n4048), .Z(n3187) );
  NAND U4063 ( .A(n2748), .B(n2588), .Z(n2589) );
  XNOR U4064 ( .A(n3187), .B(n2589), .Z(out[246]) );
  XNOR U4065 ( .A(in[1024]), .B(n4051), .Z(n3211) );
  NAND U4066 ( .A(n2750), .B(n2590), .Z(n2591) );
  XNOR U4067 ( .A(n3211), .B(n2591), .Z(out[247]) );
  XNOR U4068 ( .A(in[1025]), .B(n4054), .Z(n3235) );
  NAND U4069 ( .A(n2752), .B(n2592), .Z(n2593) );
  XNOR U4070 ( .A(n3235), .B(n2593), .Z(out[248]) );
  XNOR U4071 ( .A(in[1026]), .B(n4057), .Z(n3267) );
  NAND U4072 ( .A(n2754), .B(n2594), .Z(n2595) );
  XNOR U4073 ( .A(n3267), .B(n2595), .Z(out[249]) );
  XNOR U4074 ( .A(in[1434]), .B(n3678), .Z(n4324) );
  NANDN U4075 ( .A(n2677), .B(n4324), .Z(n2596) );
  XNOR U4076 ( .A(n4325), .B(n2596), .Z(out[24]) );
  XNOR U4077 ( .A(in[1027]), .B(n4060), .Z(n3311) );
  NAND U4078 ( .A(n2756), .B(n2597), .Z(n2598) );
  XNOR U4079 ( .A(n3311), .B(n2598), .Z(out[250]) );
  XNOR U4080 ( .A(in[1028]), .B(n4063), .Z(n3355) );
  NAND U4081 ( .A(n2758), .B(n2599), .Z(n2600) );
  XNOR U4082 ( .A(n3355), .B(n2600), .Z(out[251]) );
  XNOR U4083 ( .A(in[1029]), .B(n4066), .Z(n3401) );
  NAND U4084 ( .A(n2760), .B(n2601), .Z(n2602) );
  XNOR U4085 ( .A(n3401), .B(n2602), .Z(out[252]) );
  XNOR U4086 ( .A(in[1030]), .B(n4069), .Z(n3445) );
  NAND U4087 ( .A(n2762), .B(n2603), .Z(n2604) );
  XNOR U4088 ( .A(n3445), .B(n2604), .Z(out[253]) );
  XNOR U4089 ( .A(in[1031]), .B(n4080), .Z(n3489) );
  NAND U4090 ( .A(n2764), .B(n2605), .Z(n2606) );
  XNOR U4091 ( .A(n3489), .B(n2606), .Z(out[254]) );
  XNOR U4092 ( .A(in[1032]), .B(n4083), .Z(n3533) );
  NAND U4093 ( .A(n2766), .B(n2607), .Z(n2608) );
  XNOR U4094 ( .A(n3533), .B(n2608), .Z(out[255]) );
  ANDN U4095 ( .B(n2610), .A(n2609), .Z(n2611) );
  XNOR U4096 ( .A(n3576), .B(n2611), .Z(out[256]) );
  AND U4097 ( .A(n2613), .B(n2612), .Z(n2614) );
  XNOR U4098 ( .A(n3620), .B(n2614), .Z(out[257]) );
  XOR U4099 ( .A(n3582), .B(in[1412]), .Z(n3665) );
  NAND U4100 ( .A(n2724), .B(n2615), .Z(n2616) );
  XNOR U4101 ( .A(n3665), .B(n2616), .Z(out[258]) );
  XOR U4102 ( .A(n3586), .B(in[1413]), .Z(n3709) );
  NAND U4103 ( .A(n2874), .B(n2617), .Z(n2618) );
  XNOR U4104 ( .A(n3709), .B(n2618), .Z(out[259]) );
  XNOR U4105 ( .A(in[1435]), .B(n3682), .Z(n4356) );
  NANDN U4106 ( .A(n2680), .B(n4356), .Z(n2619) );
  XNOR U4107 ( .A(n4357), .B(n2619), .Z(out[25]) );
  XOR U4108 ( .A(n3590), .B(in[1414]), .Z(n3753) );
  NAND U4109 ( .A(n3068), .B(n2620), .Z(n2621) );
  XNOR U4110 ( .A(n3753), .B(n2621), .Z(out[260]) );
  XOR U4111 ( .A(n3594), .B(in[1415]), .Z(n3797) );
  NAND U4112 ( .A(n3358), .B(n2622), .Z(n2623) );
  XNOR U4113 ( .A(n3797), .B(n2623), .Z(out[261]) );
  XOR U4114 ( .A(n3598), .B(in[1416]), .Z(n3831) );
  NAND U4115 ( .A(n3800), .B(n2624), .Z(n2625) );
  XNOR U4116 ( .A(n3831), .B(n2625), .Z(out[262]) );
  XOR U4117 ( .A(in[1417]), .B(n3602), .Z(n4077) );
  NAND U4118 ( .A(n4076), .B(n2626), .Z(n2627) );
  XNOR U4119 ( .A(n4077), .B(n2627), .Z(out[263]) );
  XOR U4120 ( .A(n3606), .B(in[1418]), .Z(n4361) );
  NAND U4121 ( .A(n4360), .B(n2628), .Z(n2629) );
  XNOR U4122 ( .A(n4361), .B(n2629), .Z(out[264]) );
  XOR U4123 ( .A(n3610), .B(in[1419]), .Z(n4805) );
  NAND U4124 ( .A(n4804), .B(n2630), .Z(n2631) );
  XNOR U4125 ( .A(n4805), .B(n2631), .Z(out[265]) );
  ANDN U4126 ( .B(n2633), .A(n2632), .Z(n2634) );
  XNOR U4127 ( .A(n3920), .B(n2634), .Z(out[266]) );
  ANDN U4128 ( .B(n2636), .A(n2635), .Z(n2637) );
  XNOR U4129 ( .A(n3944), .B(n2637), .Z(out[267]) );
  ANDN U4130 ( .B(n2639), .A(n2638), .Z(n2640) );
  XNOR U4131 ( .A(n3970), .B(n2640), .Z(out[268]) );
  ANDN U4132 ( .B(n2642), .A(n2641), .Z(n2643) );
  XNOR U4133 ( .A(n4004), .B(n2643), .Z(out[269]) );
  XNOR U4134 ( .A(in[1436]), .B(n3686), .Z(n4404) );
  NANDN U4135 ( .A(n2683), .B(n4404), .Z(n2644) );
  XNOR U4136 ( .A(n4405), .B(n2644), .Z(out[26]) );
  ANDN U4137 ( .B(n2646), .A(n2645), .Z(n2647) );
  XNOR U4138 ( .A(n4038), .B(n2647), .Z(out[270]) );
  ANDN U4139 ( .B(n2649), .A(n2648), .Z(n2650) );
  XNOR U4140 ( .A(n4072), .B(n2650), .Z(out[271]) );
  ANDN U4141 ( .B(n2652), .A(n2651), .Z(n2653) );
  XNOR U4142 ( .A(n4110), .B(n2653), .Z(out[272]) );
  ANDN U4143 ( .B(n2655), .A(n2654), .Z(n2656) );
  XNOR U4144 ( .A(n4144), .B(n2656), .Z(out[273]) );
  ANDN U4145 ( .B(n2658), .A(n2657), .Z(n2659) );
  XNOR U4146 ( .A(n4178), .B(n2659), .Z(out[274]) );
  ANDN U4147 ( .B(n2661), .A(n2660), .Z(n2662) );
  XNOR U4148 ( .A(n4204), .B(n2662), .Z(out[275]) );
  ANDN U4149 ( .B(n2664), .A(n2663), .Z(n2665) );
  XNOR U4150 ( .A(n4228), .B(n2665), .Z(out[276]) );
  AND U4151 ( .A(n2667), .B(n2666), .Z(n2668) );
  XNOR U4152 ( .A(n4252), .B(n2668), .Z(out[277]) );
  AND U4153 ( .A(n2670), .B(n2669), .Z(n2671) );
  XNOR U4154 ( .A(n4276), .B(n2671), .Z(out[278]) );
  AND U4155 ( .A(n2673), .B(n2672), .Z(n2674) );
  XNOR U4156 ( .A(n4300), .B(n2674), .Z(out[279]) );
  XNOR U4157 ( .A(in[1437]), .B(n3690), .Z(n4448) );
  NANDN U4158 ( .A(n2686), .B(n4448), .Z(n2675) );
  XNOR U4159 ( .A(n4449), .B(n2675), .Z(out[27]) );
  AND U4160 ( .A(n2677), .B(n2676), .Z(n2678) );
  XNOR U4161 ( .A(n4324), .B(n2678), .Z(out[280]) );
  AND U4162 ( .A(n2680), .B(n2679), .Z(n2681) );
  XNOR U4163 ( .A(n4356), .B(n2681), .Z(out[281]) );
  AND U4164 ( .A(n2683), .B(n2682), .Z(n2684) );
  XNOR U4165 ( .A(n4404), .B(n2684), .Z(out[282]) );
  AND U4166 ( .A(n2686), .B(n2685), .Z(n2687) );
  XNOR U4167 ( .A(n4448), .B(n2687), .Z(out[283]) );
  XOR U4168 ( .A(in[1438]), .B(n3694), .Z(n4493) );
  NAND U4169 ( .A(n2700), .B(n2688), .Z(n2689) );
  XNOR U4170 ( .A(n4493), .B(n2689), .Z(out[284]) );
  XOR U4171 ( .A(in[1439]), .B(n3698), .Z(n4537) );
  NAND U4172 ( .A(n2722), .B(n2690), .Z(n2691) );
  XNOR U4173 ( .A(n4537), .B(n2691), .Z(out[285]) );
  XOR U4174 ( .A(in[1440]), .B(n3702), .Z(n4581) );
  NAND U4175 ( .A(n2746), .B(n2692), .Z(n2693) );
  XNOR U4176 ( .A(n4581), .B(n2693), .Z(out[286]) );
  XOR U4177 ( .A(in[1441]), .B(n3706), .Z(n4625) );
  NAND U4178 ( .A(n2768), .B(n2694), .Z(n2695) );
  XNOR U4179 ( .A(n4625), .B(n2695), .Z(out[287]) );
  XOR U4180 ( .A(in[1442]), .B(n3714), .Z(n4669) );
  NAND U4181 ( .A(n2780), .B(n2696), .Z(n2697) );
  XNOR U4182 ( .A(n4669), .B(n2697), .Z(out[288]) );
  XOR U4183 ( .A(in[1443]), .B(n3718), .Z(n4713) );
  NAND U4184 ( .A(n2792), .B(n2698), .Z(n2699) );
  XNOR U4185 ( .A(n4713), .B(n2699), .Z(out[289]) );
  OR U4186 ( .A(n4493), .B(n2700), .Z(n2701) );
  XNOR U4187 ( .A(n4492), .B(n2701), .Z(out[28]) );
  XOR U4188 ( .A(in[1444]), .B(n3722), .Z(n4757) );
  NAND U4189 ( .A(n2804), .B(n2702), .Z(n2703) );
  XNOR U4190 ( .A(n4757), .B(n2703), .Z(out[290]) );
  XOR U4191 ( .A(in[1445]), .B(n3726), .Z(n4801) );
  NAND U4192 ( .A(n2816), .B(n2704), .Z(n2705) );
  XNOR U4193 ( .A(n4801), .B(n2705), .Z(out[291]) );
  OR U4194 ( .A(n2829), .B(n2706), .Z(n2707) );
  XNOR U4195 ( .A(n2828), .B(n2707), .Z(out[292]) );
  OR U4196 ( .A(n2843), .B(n2708), .Z(n2709) );
  XNOR U4197 ( .A(n2842), .B(n2709), .Z(out[293]) );
  OR U4198 ( .A(n2857), .B(n2710), .Z(n2711) );
  XNOR U4199 ( .A(n2856), .B(n2711), .Z(out[294]) );
  OR U4200 ( .A(n2871), .B(n2712), .Z(n2713) );
  XNOR U4201 ( .A(n2870), .B(n2713), .Z(out[295]) );
  OR U4202 ( .A(n2887), .B(n2714), .Z(n2715) );
  XNOR U4203 ( .A(n2886), .B(n2715), .Z(out[296]) );
  OR U4204 ( .A(n2901), .B(n2716), .Z(n2717) );
  XNOR U4205 ( .A(n2900), .B(n2717), .Z(out[297]) );
  OR U4206 ( .A(n2915), .B(n2718), .Z(n2719) );
  XNOR U4207 ( .A(n2914), .B(n2719), .Z(out[298]) );
  OR U4208 ( .A(n2929), .B(n2720), .Z(n2721) );
  XNOR U4209 ( .A(n2928), .B(n2721), .Z(out[299]) );
  OR U4210 ( .A(n4537), .B(n2722), .Z(n2723) );
  XNOR U4211 ( .A(n4536), .B(n2723), .Z(out[29]) );
  OR U4212 ( .A(n3665), .B(n2724), .Z(n2725) );
  XNOR U4213 ( .A(n3664), .B(n2725), .Z(out[2]) );
  OR U4214 ( .A(n2945), .B(n2726), .Z(n2727) );
  XNOR U4215 ( .A(n2944), .B(n2727), .Z(out[300]) );
  OR U4216 ( .A(n2969), .B(n2728), .Z(n2729) );
  XNOR U4217 ( .A(n2968), .B(n2729), .Z(out[301]) );
  OR U4218 ( .A(n2993), .B(n2730), .Z(n2731) );
  XNOR U4219 ( .A(n2992), .B(n2731), .Z(out[302]) );
  OR U4220 ( .A(n3017), .B(n2732), .Z(n2733) );
  XNOR U4221 ( .A(n3016), .B(n2733), .Z(out[303]) );
  OR U4222 ( .A(n3041), .B(n2734), .Z(n2735) );
  XNOR U4223 ( .A(n3040), .B(n2735), .Z(out[304]) );
  OR U4224 ( .A(n3065), .B(n2736), .Z(n2737) );
  XNOR U4225 ( .A(n3064), .B(n2737), .Z(out[305]) );
  OR U4226 ( .A(n3091), .B(n2738), .Z(n2739) );
  XNOR U4227 ( .A(n3090), .B(n2739), .Z(out[306]) );
  OR U4228 ( .A(n3115), .B(n2740), .Z(n2741) );
  XNOR U4229 ( .A(n3114), .B(n2741), .Z(out[307]) );
  OR U4230 ( .A(n3139), .B(n2742), .Z(n2743) );
  XNOR U4231 ( .A(n3138), .B(n2743), .Z(out[308]) );
  OR U4232 ( .A(n3163), .B(n2744), .Z(n2745) );
  XNOR U4233 ( .A(n3162), .B(n2745), .Z(out[309]) );
  OR U4234 ( .A(n4581), .B(n2746), .Z(n2747) );
  XNOR U4235 ( .A(n4580), .B(n2747), .Z(out[30]) );
  OR U4236 ( .A(n3187), .B(n2748), .Z(n2749) );
  XNOR U4237 ( .A(n3186), .B(n2749), .Z(out[310]) );
  OR U4238 ( .A(n3211), .B(n2750), .Z(n2751) );
  XNOR U4239 ( .A(n3210), .B(n2751), .Z(out[311]) );
  OR U4240 ( .A(n3235), .B(n2752), .Z(n2753) );
  XNOR U4241 ( .A(n3234), .B(n2753), .Z(out[312]) );
  OR U4242 ( .A(n3267), .B(n2754), .Z(n2755) );
  XNOR U4243 ( .A(n3266), .B(n2755), .Z(out[313]) );
  OR U4244 ( .A(n3311), .B(n2756), .Z(n2757) );
  XNOR U4245 ( .A(n3310), .B(n2757), .Z(out[314]) );
  OR U4246 ( .A(n3355), .B(n2758), .Z(n2759) );
  XNOR U4247 ( .A(n3354), .B(n2759), .Z(out[315]) );
  OR U4248 ( .A(n3401), .B(n2760), .Z(n2761) );
  XNOR U4249 ( .A(n3400), .B(n2761), .Z(out[316]) );
  OR U4250 ( .A(n3445), .B(n2762), .Z(n2763) );
  XNOR U4251 ( .A(n3444), .B(n2763), .Z(out[317]) );
  OR U4252 ( .A(n3489), .B(n2764), .Z(n2765) );
  XNOR U4253 ( .A(n3488), .B(n2765), .Z(out[318]) );
  OR U4254 ( .A(n3533), .B(n2766), .Z(n2767) );
  XNOR U4255 ( .A(n3532), .B(n2767), .Z(out[319]) );
  OR U4256 ( .A(n4625), .B(n2768), .Z(n2769) );
  XNOR U4257 ( .A(n4624), .B(n2769), .Z(out[31]) );
  XNOR U4258 ( .A(in[72]), .B(n4083), .Z(n2940) );
  XOR U4259 ( .A(in[1317]), .B(n3918), .Z(n3253) );
  XOR U4260 ( .A(in[1244]), .B(n3736), .Z(n3250) );
  NAND U4261 ( .A(n3253), .B(n3250), .Z(n2770) );
  XNOR U4262 ( .A(n2940), .B(n2770), .Z(out[320]) );
  XNOR U4263 ( .A(in[73]), .B(n4086), .Z(n2942) );
  XOR U4264 ( .A(in[1318]), .B(n3924), .Z(n3257) );
  XOR U4265 ( .A(in[1245]), .B(n3740), .Z(n3254) );
  NAND U4266 ( .A(n3257), .B(n3254), .Z(n2771) );
  XNOR U4267 ( .A(n2942), .B(n2771), .Z(out[321]) );
  XNOR U4268 ( .A(in[74]), .B(n4089), .Z(n2948) );
  XOR U4269 ( .A(in[1319]), .B(n3926), .Z(n3261) );
  XOR U4270 ( .A(in[1246]), .B(n3744), .Z(n3258) );
  NAND U4271 ( .A(n3261), .B(n3258), .Z(n2772) );
  XNOR U4272 ( .A(n2948), .B(n2772), .Z(out[322]) );
  XNOR U4273 ( .A(in[75]), .B(n4092), .Z(n2950) );
  XOR U4274 ( .A(in[1320]), .B(n3928), .Z(n3265) );
  XOR U4275 ( .A(in[1247]), .B(n3748), .Z(n3262) );
  NAND U4276 ( .A(n3265), .B(n3262), .Z(n2773) );
  XNOR U4277 ( .A(n2950), .B(n2773), .Z(out[323]) );
  XOR U4278 ( .A(n4095), .B(in[76]), .Z(n2952) );
  XOR U4279 ( .A(in[1321]), .B(n3930), .Z(n3273) );
  XOR U4280 ( .A(in[1248]), .B(n3756), .Z(n3270) );
  NAND U4281 ( .A(n3273), .B(n3270), .Z(n2774) );
  XNOR U4282 ( .A(n2952), .B(n2774), .Z(out[324]) );
  XOR U4283 ( .A(n4098), .B(in[77]), .Z(n2954) );
  XOR U4284 ( .A(in[1322]), .B(n3932), .Z(n3277) );
  XOR U4285 ( .A(in[1249]), .B(n3760), .Z(n3274) );
  NAND U4286 ( .A(n3277), .B(n3274), .Z(n2775) );
  XNOR U4287 ( .A(n2954), .B(n2775), .Z(out[325]) );
  XOR U4288 ( .A(n4101), .B(in[78]), .Z(n2956) );
  XOR U4289 ( .A(in[1323]), .B(n3934), .Z(n3281) );
  XOR U4290 ( .A(in[1250]), .B(n3764), .Z(n3278) );
  NAND U4291 ( .A(n3281), .B(n3278), .Z(n2776) );
  XNOR U4292 ( .A(n2956), .B(n2776), .Z(out[326]) );
  XOR U4293 ( .A(n4104), .B(in[79]), .Z(n2958) );
  XOR U4294 ( .A(in[1324]), .B(n3936), .Z(n3285) );
  XOR U4295 ( .A(in[1251]), .B(n3768), .Z(n3282) );
  NAND U4296 ( .A(n3285), .B(n3282), .Z(n2777) );
  XNOR U4297 ( .A(n2958), .B(n2777), .Z(out[327]) );
  XOR U4298 ( .A(n4107), .B(in[80]), .Z(n2960) );
  XOR U4299 ( .A(in[1325]), .B(n3938), .Z(n3289) );
  XOR U4300 ( .A(in[1252]), .B(n3772), .Z(n3286) );
  NAND U4301 ( .A(n3289), .B(n3286), .Z(n2778) );
  XNOR U4302 ( .A(n2960), .B(n2778), .Z(out[328]) );
  XOR U4303 ( .A(n4114), .B(in[81]), .Z(n2962) );
  XOR U4304 ( .A(in[1326]), .B(n3940), .Z(n3293) );
  XNOR U4305 ( .A(in[1253]), .B(n3776), .Z(n3290) );
  NAND U4306 ( .A(n3293), .B(n3290), .Z(n2779) );
  XNOR U4307 ( .A(n2962), .B(n2779), .Z(out[329]) );
  OR U4308 ( .A(n4669), .B(n2780), .Z(n2781) );
  XNOR U4309 ( .A(n4668), .B(n2781), .Z(out[32]) );
  XOR U4310 ( .A(n4117), .B(in[82]), .Z(n2964) );
  XOR U4311 ( .A(in[1327]), .B(n3942), .Z(n3297) );
  XNOR U4312 ( .A(in[1254]), .B(n3780), .Z(n3294) );
  NAND U4313 ( .A(n3297), .B(n3294), .Z(n2782) );
  XNOR U4314 ( .A(n2964), .B(n2782), .Z(out[330]) );
  XOR U4315 ( .A(n4120), .B(in[83]), .Z(n2966) );
  XOR U4316 ( .A(in[1328]), .B(n3948), .Z(n3301) );
  XNOR U4317 ( .A(in[1255]), .B(n3784), .Z(n3298) );
  NAND U4318 ( .A(n3301), .B(n3298), .Z(n2783) );
  XNOR U4319 ( .A(n2966), .B(n2783), .Z(out[331]) );
  XOR U4320 ( .A(in[84]), .B(n4123), .Z(n2972) );
  XOR U4321 ( .A(in[1329]), .B(n3950), .Z(n3305) );
  XNOR U4322 ( .A(in[1256]), .B(n3788), .Z(n3302) );
  NAND U4323 ( .A(n3305), .B(n3302), .Z(n2784) );
  XNOR U4324 ( .A(n2972), .B(n2784), .Z(out[332]) );
  XOR U4325 ( .A(in[85]), .B(n4126), .Z(n2974) );
  XOR U4326 ( .A(in[1330]), .B(n3952), .Z(n3309) );
  XNOR U4327 ( .A(in[1257]), .B(n3792), .Z(n3306) );
  NAND U4328 ( .A(n3309), .B(n3306), .Z(n2785) );
  XNOR U4329 ( .A(n2974), .B(n2785), .Z(out[333]) );
  XOR U4330 ( .A(in[86]), .B(n4129), .Z(n2976) );
  XOR U4331 ( .A(in[1331]), .B(n3954), .Z(n3317) );
  XNOR U4332 ( .A(in[1258]), .B(n3802), .Z(n3314) );
  NAND U4333 ( .A(n3317), .B(n3314), .Z(n2786) );
  XNOR U4334 ( .A(n2976), .B(n2786), .Z(out[334]) );
  XOR U4335 ( .A(in[87]), .B(n4132), .Z(n2978) );
  XOR U4336 ( .A(in[1332]), .B(n3956), .Z(n3321) );
  XNOR U4337 ( .A(in[1259]), .B(n3806), .Z(n3318) );
  NAND U4338 ( .A(n3321), .B(n3318), .Z(n2787) );
  XNOR U4339 ( .A(n2978), .B(n2787), .Z(out[335]) );
  XOR U4340 ( .A(in[88]), .B(n4135), .Z(n2980) );
  XOR U4341 ( .A(in[1333]), .B(n3958), .Z(n3325) );
  XNOR U4342 ( .A(in[1260]), .B(n3810), .Z(n3322) );
  NAND U4343 ( .A(n3325), .B(n3322), .Z(n2788) );
  XNOR U4344 ( .A(n2980), .B(n2788), .Z(out[336]) );
  XOR U4345 ( .A(in[89]), .B(n4138), .Z(n2982) );
  XOR U4346 ( .A(in[1334]), .B(n3960), .Z(n3329) );
  XNOR U4347 ( .A(in[1261]), .B(n3814), .Z(n3326) );
  NAND U4348 ( .A(n3329), .B(n3326), .Z(n2789) );
  XNOR U4349 ( .A(n2982), .B(n2789), .Z(out[337]) );
  XOR U4350 ( .A(in[90]), .B(n4141), .Z(n2984) );
  XOR U4351 ( .A(in[1335]), .B(n3962), .Z(n3333) );
  XNOR U4352 ( .A(in[1262]), .B(n3536), .Z(n3330) );
  NAND U4353 ( .A(n3333), .B(n3330), .Z(n2790) );
  XNOR U4354 ( .A(n2984), .B(n2790), .Z(out[338]) );
  XOR U4355 ( .A(in[91]), .B(n4148), .Z(n2986) );
  XOR U4356 ( .A(in[1336]), .B(n3818), .Z(n3337) );
  XNOR U4357 ( .A(in[1263]), .B(n3540), .Z(n3334) );
  NAND U4358 ( .A(n3337), .B(n3334), .Z(n2791) );
  XNOR U4359 ( .A(n2986), .B(n2791), .Z(out[339]) );
  OR U4360 ( .A(n4713), .B(n2792), .Z(n2793) );
  XNOR U4361 ( .A(n4712), .B(n2793), .Z(out[33]) );
  XOR U4362 ( .A(in[92]), .B(n4151), .Z(n2988) );
  XOR U4363 ( .A(in[1337]), .B(n3820), .Z(n3341) );
  XNOR U4364 ( .A(in[1264]), .B(n3544), .Z(n3338) );
  NAND U4365 ( .A(n3341), .B(n3338), .Z(n2794) );
  XNOR U4366 ( .A(n2988), .B(n2794), .Z(out[340]) );
  XOR U4367 ( .A(in[93]), .B(n4154), .Z(n2990) );
  XOR U4368 ( .A(in[1338]), .B(n3822), .Z(n3345) );
  XNOR U4369 ( .A(in[1265]), .B(n3548), .Z(n3342) );
  NAND U4370 ( .A(n3345), .B(n3342), .Z(n2795) );
  XNOR U4371 ( .A(n2990), .B(n2795), .Z(out[341]) );
  XOR U4372 ( .A(in[94]), .B(n4157), .Z(n2996) );
  XOR U4373 ( .A(in[1339]), .B(n3824), .Z(n3349) );
  XNOR U4374 ( .A(in[1266]), .B(n3552), .Z(n3346) );
  NAND U4375 ( .A(n3349), .B(n3346), .Z(n2796) );
  XNOR U4376 ( .A(n2996), .B(n2796), .Z(out[342]) );
  XOR U4377 ( .A(in[95]), .B(n4160), .Z(n2998) );
  XOR U4378 ( .A(in[1340]), .B(n3826), .Z(n3353) );
  XNOR U4379 ( .A(in[1267]), .B(n3556), .Z(n3350) );
  NAND U4380 ( .A(n3353), .B(n3350), .Z(n2797) );
  XNOR U4381 ( .A(n2998), .B(n2797), .Z(out[343]) );
  XOR U4382 ( .A(in[96]), .B(n4163), .Z(n3000) );
  XOR U4383 ( .A(in[1341]), .B(n3828), .Z(n3363) );
  XNOR U4384 ( .A(in[1268]), .B(n3560), .Z(n3360) );
  NAND U4385 ( .A(n3363), .B(n3360), .Z(n2798) );
  XNOR U4386 ( .A(n3000), .B(n2798), .Z(out[344]) );
  XOR U4387 ( .A(in[97]), .B(n4166), .Z(n3002) );
  XOR U4388 ( .A(in[1342]), .B(n3834), .Z(n3367) );
  XNOR U4389 ( .A(in[1269]), .B(n3564), .Z(n3364) );
  NAND U4390 ( .A(n3367), .B(n3364), .Z(n2799) );
  XNOR U4391 ( .A(n3002), .B(n2799), .Z(out[345]) );
  XOR U4392 ( .A(in[98]), .B(n4169), .Z(n3004) );
  XOR U4393 ( .A(in[1343]), .B(n3836), .Z(n3371) );
  XNOR U4394 ( .A(in[1270]), .B(n3568), .Z(n3368) );
  NAND U4395 ( .A(n3371), .B(n3368), .Z(n2800) );
  XNOR U4396 ( .A(n3004), .B(n2800), .Z(out[346]) );
  XOR U4397 ( .A(in[99]), .B(n4172), .Z(n3006) );
  XOR U4398 ( .A(in[1280]), .B(n3838), .Z(n3375) );
  XNOR U4399 ( .A(in[1271]), .B(n3572), .Z(n3372) );
  NAND U4400 ( .A(n3375), .B(n3372), .Z(n2801) );
  XNOR U4401 ( .A(n3006), .B(n2801), .Z(out[347]) );
  XNOR U4402 ( .A(in[100]), .B(n4175), .Z(n3008) );
  XOR U4403 ( .A(in[1281]), .B(n3840), .Z(n3379) );
  XNOR U4404 ( .A(in[1272]), .B(n3580), .Z(n3376) );
  NAND U4405 ( .A(n3379), .B(n3376), .Z(n2802) );
  XNOR U4406 ( .A(n3008), .B(n2802), .Z(out[348]) );
  XNOR U4407 ( .A(in[101]), .B(n4182), .Z(n3010) );
  XOR U4408 ( .A(in[1282]), .B(n3842), .Z(n3383) );
  XNOR U4409 ( .A(in[1273]), .B(n3584), .Z(n3380) );
  NAND U4410 ( .A(n3383), .B(n3380), .Z(n2803) );
  XNOR U4411 ( .A(n3010), .B(n2803), .Z(out[349]) );
  OR U4412 ( .A(n4757), .B(n2804), .Z(n2805) );
  XNOR U4413 ( .A(n4756), .B(n2805), .Z(out[34]) );
  XNOR U4414 ( .A(in[102]), .B(n4185), .Z(n3012) );
  XOR U4415 ( .A(in[1283]), .B(n3844), .Z(n3387) );
  XNOR U4416 ( .A(in[1274]), .B(n3588), .Z(n3384) );
  NAND U4417 ( .A(n3387), .B(n3384), .Z(n2806) );
  XNOR U4418 ( .A(n3012), .B(n2806), .Z(out[350]) );
  XNOR U4419 ( .A(in[103]), .B(n3964), .Z(n3014) );
  XOR U4420 ( .A(in[1284]), .B(n3846), .Z(n3391) );
  XNOR U4421 ( .A(in[1275]), .B(n3592), .Z(n3388) );
  NAND U4422 ( .A(n3391), .B(n3388), .Z(n2807) );
  XNOR U4423 ( .A(n3014), .B(n2807), .Z(out[351]) );
  XNOR U4424 ( .A(in[104]), .B(n3967), .Z(n3020) );
  XOR U4425 ( .A(in[1285]), .B(n3848), .Z(n3395) );
  XNOR U4426 ( .A(in[1276]), .B(n3596), .Z(n3392) );
  NAND U4427 ( .A(n3395), .B(n3392), .Z(n2808) );
  XNOR U4428 ( .A(n3020), .B(n2808), .Z(out[352]) );
  XNOR U4429 ( .A(in[105]), .B(n3974), .Z(n3022) );
  XOR U4430 ( .A(in[1286]), .B(n3850), .Z(n3399) );
  XNOR U4431 ( .A(in[1277]), .B(n3600), .Z(n3396) );
  NAND U4432 ( .A(n3399), .B(n3396), .Z(n2809) );
  XNOR U4433 ( .A(n3022), .B(n2809), .Z(out[353]) );
  XNOR U4434 ( .A(in[106]), .B(n3977), .Z(n3024) );
  XOR U4435 ( .A(in[1287]), .B(n3852), .Z(n3407) );
  XNOR U4436 ( .A(in[1278]), .B(n3604), .Z(n3404) );
  NAND U4437 ( .A(n3407), .B(n3404), .Z(n2810) );
  XNOR U4438 ( .A(n3024), .B(n2810), .Z(out[354]) );
  XNOR U4439 ( .A(in[107]), .B(n3980), .Z(n3026) );
  XOR U4440 ( .A(in[1288]), .B(n3856), .Z(n3411) );
  XNOR U4441 ( .A(in[1279]), .B(n3608), .Z(n3408) );
  NAND U4442 ( .A(n3411), .B(n3408), .Z(n2811) );
  XNOR U4443 ( .A(n3026), .B(n2811), .Z(out[355]) );
  XNOR U4444 ( .A(in[108]), .B(n3983), .Z(n3028) );
  XOR U4445 ( .A(in[1289]), .B(n3858), .Z(n3415) );
  XNOR U4446 ( .A(in[1216]), .B(n3612), .Z(n3412) );
  NAND U4447 ( .A(n3415), .B(n3412), .Z(n2812) );
  XNOR U4448 ( .A(n3028), .B(n2812), .Z(out[356]) );
  XNOR U4449 ( .A(in[109]), .B(n3986), .Z(n3030) );
  XOR U4450 ( .A(in[1290]), .B(n3860), .Z(n3419) );
  XNOR U4451 ( .A(in[1217]), .B(n3616), .Z(n3416) );
  NAND U4452 ( .A(n3419), .B(n3416), .Z(n2813) );
  XNOR U4453 ( .A(n3030), .B(n2813), .Z(out[357]) );
  XNOR U4454 ( .A(in[110]), .B(n3989), .Z(n3032) );
  XOR U4455 ( .A(in[1291]), .B(n3862), .Z(n3423) );
  XNOR U4456 ( .A(in[1218]), .B(n3624), .Z(n3420) );
  NAND U4457 ( .A(n3423), .B(n3420), .Z(n2814) );
  XNOR U4458 ( .A(n3032), .B(n2814), .Z(out[358]) );
  XNOR U4459 ( .A(in[111]), .B(n3992), .Z(n3034) );
  XOR U4460 ( .A(in[1292]), .B(n3864), .Z(n3427) );
  XNOR U4461 ( .A(in[1219]), .B(n3628), .Z(n3424) );
  NAND U4462 ( .A(n3427), .B(n3424), .Z(n2815) );
  XNOR U4463 ( .A(n3034), .B(n2815), .Z(out[359]) );
  OR U4464 ( .A(n4801), .B(n2816), .Z(n2817) );
  XNOR U4465 ( .A(n4800), .B(n2817), .Z(out[35]) );
  XNOR U4466 ( .A(in[112]), .B(n3995), .Z(n3036) );
  XOR U4467 ( .A(in[1293]), .B(n3866), .Z(n3431) );
  XOR U4468 ( .A(in[1220]), .B(n3632), .Z(n3428) );
  NAND U4469 ( .A(n3431), .B(n3428), .Z(n2818) );
  XNOR U4470 ( .A(n3036), .B(n2818), .Z(out[360]) );
  XNOR U4471 ( .A(in[113]), .B(n3998), .Z(n3038) );
  XOR U4472 ( .A(in[1294]), .B(n3868), .Z(n3435) );
  XOR U4473 ( .A(in[1221]), .B(n3636), .Z(n3432) );
  NAND U4474 ( .A(n3435), .B(n3432), .Z(n2819) );
  XNOR U4475 ( .A(n3038), .B(n2819), .Z(out[361]) );
  XNOR U4476 ( .A(in[114]), .B(n4001), .Z(n3044) );
  XOR U4477 ( .A(in[1295]), .B(n3870), .Z(n3439) );
  XOR U4478 ( .A(in[1222]), .B(n3640), .Z(n3436) );
  NAND U4479 ( .A(n3439), .B(n3436), .Z(n2820) );
  XNOR U4480 ( .A(n3044), .B(n2820), .Z(out[362]) );
  XNOR U4481 ( .A(in[115]), .B(n4008), .Z(n3046) );
  XOR U4482 ( .A(in[1296]), .B(n3872), .Z(n3443) );
  XOR U4483 ( .A(in[1223]), .B(n3644), .Z(n3440) );
  NAND U4484 ( .A(n3443), .B(n3440), .Z(n2821) );
  XNOR U4485 ( .A(n3046), .B(n2821), .Z(out[363]) );
  XNOR U4486 ( .A(in[116]), .B(n4011), .Z(n3048) );
  XOR U4487 ( .A(in[1297]), .B(n3874), .Z(n3451) );
  XOR U4488 ( .A(in[1224]), .B(n3648), .Z(n3448) );
  NAND U4489 ( .A(n3451), .B(n3448), .Z(n2822) );
  XNOR U4490 ( .A(n3048), .B(n2822), .Z(out[364]) );
  XNOR U4491 ( .A(in[117]), .B(n4014), .Z(n3050) );
  XOR U4492 ( .A(in[1298]), .B(n3878), .Z(n3455) );
  XOR U4493 ( .A(in[1225]), .B(n3652), .Z(n3452) );
  NAND U4494 ( .A(n3455), .B(n3452), .Z(n2823) );
  XNOR U4495 ( .A(n3050), .B(n2823), .Z(out[365]) );
  XNOR U4496 ( .A(in[118]), .B(n4017), .Z(n3052) );
  XOR U4497 ( .A(in[1299]), .B(n3880), .Z(n3459) );
  XOR U4498 ( .A(in[1226]), .B(n3656), .Z(n3456) );
  NAND U4499 ( .A(n3459), .B(n3456), .Z(n2824) );
  XNOR U4500 ( .A(n3052), .B(n2824), .Z(out[366]) );
  XNOR U4501 ( .A(in[119]), .B(n4020), .Z(n3054) );
  XOR U4502 ( .A(in[1300]), .B(n3882), .Z(n3463) );
  XOR U4503 ( .A(in[1227]), .B(n3660), .Z(n3460) );
  NAND U4504 ( .A(n3463), .B(n3460), .Z(n2825) );
  XNOR U4505 ( .A(n3054), .B(n2825), .Z(out[367]) );
  XNOR U4506 ( .A(in[120]), .B(n4023), .Z(n3056) );
  XOR U4507 ( .A(in[1301]), .B(n3884), .Z(n3467) );
  XOR U4508 ( .A(in[1228]), .B(n3668), .Z(n3464) );
  NAND U4509 ( .A(n3467), .B(n3464), .Z(n2826) );
  XNOR U4510 ( .A(n3056), .B(n2826), .Z(out[368]) );
  XNOR U4511 ( .A(in[121]), .B(n4026), .Z(n3058) );
  XOR U4512 ( .A(in[1302]), .B(n3886), .Z(n3471) );
  XOR U4513 ( .A(in[1229]), .B(n3672), .Z(n3468) );
  NAND U4514 ( .A(n3471), .B(n3468), .Z(n2827) );
  XNOR U4515 ( .A(n3058), .B(n2827), .Z(out[369]) );
  ANDN U4516 ( .B(n2829), .A(n2828), .Z(n2830) );
  XNOR U4517 ( .A(n2831), .B(n2830), .Z(out[36]) );
  XNOR U4518 ( .A(in[122]), .B(n4029), .Z(n3060) );
  XOR U4519 ( .A(in[1303]), .B(n3888), .Z(n3475) );
  XOR U4520 ( .A(in[1230]), .B(n3676), .Z(n3472) );
  NAND U4521 ( .A(n3475), .B(n3472), .Z(n2832) );
  XNOR U4522 ( .A(n3060), .B(n2832), .Z(out[370]) );
  XNOR U4523 ( .A(in[123]), .B(n4032), .Z(n3062) );
  XOR U4524 ( .A(in[1304]), .B(n3890), .Z(n3479) );
  XOR U4525 ( .A(in[1231]), .B(n3680), .Z(n3476) );
  NAND U4526 ( .A(n3479), .B(n3476), .Z(n2833) );
  XNOR U4527 ( .A(n3062), .B(n2833), .Z(out[371]) );
  XNOR U4528 ( .A(in[124]), .B(n4035), .Z(n3070) );
  XOR U4529 ( .A(in[1305]), .B(n3892), .Z(n3483) );
  XOR U4530 ( .A(in[1232]), .B(n3684), .Z(n3480) );
  NAND U4531 ( .A(n3483), .B(n3480), .Z(n2834) );
  XNOR U4532 ( .A(n3070), .B(n2834), .Z(out[372]) );
  XNOR U4533 ( .A(in[125]), .B(n4042), .Z(n3072) );
  XOR U4534 ( .A(in[1306]), .B(n3894), .Z(n3487) );
  XOR U4535 ( .A(in[1233]), .B(n3688), .Z(n3484) );
  NAND U4536 ( .A(n3487), .B(n3484), .Z(n2835) );
  XNOR U4537 ( .A(n3072), .B(n2835), .Z(out[373]) );
  XNOR U4538 ( .A(in[126]), .B(n4045), .Z(n3074) );
  XOR U4539 ( .A(in[1307]), .B(n3896), .Z(n3495) );
  XOR U4540 ( .A(in[1234]), .B(n3692), .Z(n3492) );
  NAND U4541 ( .A(n3495), .B(n3492), .Z(n2836) );
  XNOR U4542 ( .A(n3074), .B(n2836), .Z(out[374]) );
  XNOR U4543 ( .A(in[127]), .B(n4048), .Z(n3076) );
  XOR U4544 ( .A(in[1308]), .B(n3900), .Z(n3499) );
  XOR U4545 ( .A(in[1235]), .B(n3696), .Z(n3496) );
  NAND U4546 ( .A(n3499), .B(n3496), .Z(n2837) );
  XNOR U4547 ( .A(n3076), .B(n2837), .Z(out[375]) );
  XNOR U4548 ( .A(in[64]), .B(n4051), .Z(n3078) );
  XOR U4549 ( .A(in[1309]), .B(n3902), .Z(n3503) );
  XOR U4550 ( .A(in[1236]), .B(n3700), .Z(n3500) );
  NAND U4551 ( .A(n3503), .B(n3500), .Z(n2838) );
  XNOR U4552 ( .A(n3078), .B(n2838), .Z(out[376]) );
  XNOR U4553 ( .A(in[65]), .B(n4054), .Z(n3080) );
  XOR U4554 ( .A(in[1310]), .B(n3904), .Z(n3507) );
  XOR U4555 ( .A(in[1237]), .B(n3704), .Z(n3504) );
  NAND U4556 ( .A(n3507), .B(n3504), .Z(n2839) );
  XNOR U4557 ( .A(n3080), .B(n2839), .Z(out[377]) );
  XNOR U4558 ( .A(in[66]), .B(n4057), .Z(n3082) );
  XOR U4559 ( .A(in[1311]), .B(n3906), .Z(n3511) );
  XOR U4560 ( .A(in[1238]), .B(n3712), .Z(n3508) );
  NAND U4561 ( .A(n3511), .B(n3508), .Z(n2840) );
  XNOR U4562 ( .A(n3082), .B(n2840), .Z(out[378]) );
  XNOR U4563 ( .A(in[67]), .B(n4060), .Z(n3084) );
  XOR U4564 ( .A(in[1312]), .B(n3908), .Z(n3515) );
  XOR U4565 ( .A(in[1239]), .B(n3716), .Z(n3512) );
  NAND U4566 ( .A(n3515), .B(n3512), .Z(n2841) );
  XNOR U4567 ( .A(n3084), .B(n2841), .Z(out[379]) );
  ANDN U4568 ( .B(n2843), .A(n2842), .Z(n2844) );
  XNOR U4569 ( .A(n2845), .B(n2844), .Z(out[37]) );
  XNOR U4570 ( .A(in[68]), .B(n4063), .Z(n3086) );
  XOR U4571 ( .A(in[1313]), .B(n3910), .Z(n3519) );
  XOR U4572 ( .A(in[1240]), .B(n3720), .Z(n3516) );
  NAND U4573 ( .A(n3519), .B(n3516), .Z(n2846) );
  XNOR U4574 ( .A(n3086), .B(n2846), .Z(out[380]) );
  XNOR U4575 ( .A(in[69]), .B(n4066), .Z(n3088) );
  XOR U4576 ( .A(in[1314]), .B(n3912), .Z(n3523) );
  XOR U4577 ( .A(in[1241]), .B(n3724), .Z(n3520) );
  NAND U4578 ( .A(n3523), .B(n3520), .Z(n2847) );
  XNOR U4579 ( .A(n3088), .B(n2847), .Z(out[381]) );
  XNOR U4580 ( .A(in[70]), .B(n4069), .Z(n3094) );
  XOR U4581 ( .A(in[1315]), .B(n3914), .Z(n3527) );
  XOR U4582 ( .A(in[1242]), .B(n3728), .Z(n3524) );
  NAND U4583 ( .A(n3527), .B(n3524), .Z(n2848) );
  XNOR U4584 ( .A(n3094), .B(n2848), .Z(out[382]) );
  XNOR U4585 ( .A(in[71]), .B(n4080), .Z(n3096) );
  XOR U4586 ( .A(in[1316]), .B(n3916), .Z(n3531) );
  XOR U4587 ( .A(in[1243]), .B(n3732), .Z(n3528) );
  NAND U4588 ( .A(n3531), .B(n3528), .Z(n2849) );
  XNOR U4589 ( .A(n3096), .B(n2849), .Z(out[383]) );
  XOR U4590 ( .A(in[497]), .B(n3778), .Z(n3098) );
  NOR U4591 ( .A(n2940), .B(n3253), .Z(n2850) );
  XNOR U4592 ( .A(n3098), .B(n2850), .Z(out[384]) );
  XOR U4593 ( .A(in[498]), .B(n3782), .Z(n3100) );
  NOR U4594 ( .A(n2942), .B(n3257), .Z(n2851) );
  XNOR U4595 ( .A(n3100), .B(n2851), .Z(out[385]) );
  XOR U4596 ( .A(in[499]), .B(n3786), .Z(n3102) );
  NOR U4597 ( .A(n2948), .B(n3261), .Z(n2852) );
  XNOR U4598 ( .A(n3102), .B(n2852), .Z(out[386]) );
  XOR U4599 ( .A(in[500]), .B(n3790), .Z(n3104) );
  NOR U4600 ( .A(n2950), .B(n3265), .Z(n2853) );
  XNOR U4601 ( .A(n3104), .B(n2853), .Z(out[387]) );
  XOR U4602 ( .A(in[501]), .B(n3794), .Z(n3106) );
  NOR U4603 ( .A(n2952), .B(n3273), .Z(n2854) );
  XNOR U4604 ( .A(n3106), .B(n2854), .Z(out[388]) );
  XOR U4605 ( .A(in[502]), .B(n3804), .Z(n3108) );
  NOR U4606 ( .A(n2954), .B(n3277), .Z(n2855) );
  XNOR U4607 ( .A(n3108), .B(n2855), .Z(out[389]) );
  ANDN U4608 ( .B(n2857), .A(n2856), .Z(n2858) );
  XNOR U4609 ( .A(n2859), .B(n2858), .Z(out[38]) );
  XOR U4610 ( .A(in[503]), .B(n3808), .Z(n3110) );
  NOR U4611 ( .A(n2956), .B(n3281), .Z(n2860) );
  XNOR U4612 ( .A(n3110), .B(n2860), .Z(out[390]) );
  XOR U4613 ( .A(in[504]), .B(n3812), .Z(n3112) );
  NOR U4614 ( .A(n2958), .B(n3285), .Z(n2861) );
  XNOR U4615 ( .A(n3112), .B(n2861), .Z(out[391]) );
  XOR U4616 ( .A(in[505]), .B(n3816), .Z(n3118) );
  NOR U4617 ( .A(n2960), .B(n3289), .Z(n2862) );
  XNOR U4618 ( .A(n3118), .B(n2862), .Z(out[392]) );
  XOR U4619 ( .A(in[506]), .B(n3538), .Z(n3120) );
  NOR U4620 ( .A(n2962), .B(n3293), .Z(n2863) );
  XNOR U4621 ( .A(n3120), .B(n2863), .Z(out[393]) );
  XOR U4622 ( .A(in[507]), .B(n3542), .Z(n3122) );
  NOR U4623 ( .A(n2964), .B(n3297), .Z(n2864) );
  XNOR U4624 ( .A(n3122), .B(n2864), .Z(out[394]) );
  XOR U4625 ( .A(in[508]), .B(n3546), .Z(n3124) );
  NOR U4626 ( .A(n2966), .B(n3301), .Z(n2865) );
  XNOR U4627 ( .A(n3124), .B(n2865), .Z(out[395]) );
  XOR U4628 ( .A(in[509]), .B(n3550), .Z(n3126) );
  NOR U4629 ( .A(n2972), .B(n3305), .Z(n2866) );
  XNOR U4630 ( .A(n3126), .B(n2866), .Z(out[396]) );
  XOR U4631 ( .A(in[510]), .B(n3554), .Z(n3128) );
  NOR U4632 ( .A(n2974), .B(n3309), .Z(n2867) );
  XNOR U4633 ( .A(n3128), .B(n2867), .Z(out[397]) );
  XOR U4634 ( .A(in[511]), .B(n3558), .Z(n3130) );
  NOR U4635 ( .A(n2976), .B(n3317), .Z(n2868) );
  XNOR U4636 ( .A(n3130), .B(n2868), .Z(out[398]) );
  XOR U4637 ( .A(in[448]), .B(n3562), .Z(n3132) );
  NOR U4638 ( .A(n2978), .B(n3321), .Z(n2869) );
  XNOR U4639 ( .A(n3132), .B(n2869), .Z(out[399]) );
  ANDN U4640 ( .B(n2871), .A(n2870), .Z(n2872) );
  XNOR U4641 ( .A(n2873), .B(n2872), .Z(out[39]) );
  OR U4642 ( .A(n3709), .B(n2874), .Z(n2875) );
  XNOR U4643 ( .A(n3708), .B(n2875), .Z(out[3]) );
  XOR U4644 ( .A(in[449]), .B(n3566), .Z(n3134) );
  NOR U4645 ( .A(n2980), .B(n3325), .Z(n2876) );
  XNOR U4646 ( .A(n3134), .B(n2876), .Z(out[400]) );
  XNOR U4647 ( .A(n3570), .B(in[450]), .Z(n3136) );
  NOR U4648 ( .A(n2982), .B(n3329), .Z(n2877) );
  XNOR U4649 ( .A(n3136), .B(n2877), .Z(out[401]) );
  XNOR U4650 ( .A(n3574), .B(in[451]), .Z(n3142) );
  NOR U4651 ( .A(n2984), .B(n3333), .Z(n2878) );
  XNOR U4652 ( .A(n3142), .B(n2878), .Z(out[402]) );
  XNOR U4653 ( .A(n3582), .B(in[452]), .Z(n3144) );
  NOR U4654 ( .A(n2986), .B(n3337), .Z(n2879) );
  XNOR U4655 ( .A(n3144), .B(n2879), .Z(out[403]) );
  XNOR U4656 ( .A(n3586), .B(in[453]), .Z(n3146) );
  NOR U4657 ( .A(n2988), .B(n3341), .Z(n2880) );
  XNOR U4658 ( .A(n3146), .B(n2880), .Z(out[404]) );
  XNOR U4659 ( .A(n3590), .B(in[454]), .Z(n3148) );
  NOR U4660 ( .A(n2990), .B(n3345), .Z(n2881) );
  XNOR U4661 ( .A(n3148), .B(n2881), .Z(out[405]) );
  XNOR U4662 ( .A(n3594), .B(in[455]), .Z(n3150) );
  NOR U4663 ( .A(n2996), .B(n3349), .Z(n2882) );
  XNOR U4664 ( .A(n3150), .B(n2882), .Z(out[406]) );
  XNOR U4665 ( .A(n3598), .B(in[456]), .Z(n3152) );
  NOR U4666 ( .A(n2998), .B(n3353), .Z(n2883) );
  XNOR U4667 ( .A(n3152), .B(n2883), .Z(out[407]) );
  XNOR U4668 ( .A(in[457]), .B(n3602), .Z(n3154) );
  NOR U4669 ( .A(n3000), .B(n3363), .Z(n2884) );
  XNOR U4670 ( .A(n3154), .B(n2884), .Z(out[408]) );
  XNOR U4671 ( .A(n3606), .B(in[458]), .Z(n3156) );
  NOR U4672 ( .A(n3002), .B(n3367), .Z(n2885) );
  XNOR U4673 ( .A(n3156), .B(n2885), .Z(out[409]) );
  ANDN U4674 ( .B(n2887), .A(n2886), .Z(n2888) );
  XNOR U4675 ( .A(n2889), .B(n2888), .Z(out[40]) );
  XNOR U4676 ( .A(n3610), .B(in[459]), .Z(n3158) );
  NOR U4677 ( .A(n3004), .B(n3371), .Z(n2890) );
  XNOR U4678 ( .A(n3158), .B(n2890), .Z(out[410]) );
  XNOR U4679 ( .A(in[460]), .B(n3614), .Z(n3160) );
  NOR U4680 ( .A(n3006), .B(n3375), .Z(n2891) );
  XNOR U4681 ( .A(n3160), .B(n2891), .Z(out[411]) );
  XNOR U4682 ( .A(in[461]), .B(n3618), .Z(n3166) );
  NOR U4683 ( .A(n3008), .B(n3379), .Z(n2892) );
  XNOR U4684 ( .A(n3166), .B(n2892), .Z(out[412]) );
  XNOR U4685 ( .A(in[462]), .B(n3626), .Z(n3168) );
  NOR U4686 ( .A(n3010), .B(n3383), .Z(n2893) );
  XNOR U4687 ( .A(n3168), .B(n2893), .Z(out[413]) );
  XNOR U4688 ( .A(in[463]), .B(n3630), .Z(n3170) );
  NOR U4689 ( .A(n3012), .B(n3387), .Z(n2894) );
  XNOR U4690 ( .A(n3170), .B(n2894), .Z(out[414]) );
  XNOR U4691 ( .A(in[464]), .B(n3634), .Z(n3172) );
  NOR U4692 ( .A(n3014), .B(n3391), .Z(n2895) );
  XNOR U4693 ( .A(n3172), .B(n2895), .Z(out[415]) );
  XNOR U4694 ( .A(in[465]), .B(n3638), .Z(n3174) );
  NOR U4695 ( .A(n3020), .B(n3395), .Z(n2896) );
  XNOR U4696 ( .A(n3174), .B(n2896), .Z(out[416]) );
  XNOR U4697 ( .A(in[466]), .B(n3642), .Z(n3176) );
  NOR U4698 ( .A(n3022), .B(n3399), .Z(n2897) );
  XNOR U4699 ( .A(n3176), .B(n2897), .Z(out[417]) );
  XNOR U4700 ( .A(in[467]), .B(n3646), .Z(n3178) );
  NOR U4701 ( .A(n3024), .B(n3407), .Z(n2898) );
  XNOR U4702 ( .A(n3178), .B(n2898), .Z(out[418]) );
  XNOR U4703 ( .A(in[468]), .B(n3650), .Z(n3180) );
  NOR U4704 ( .A(n3026), .B(n3411), .Z(n2899) );
  XNOR U4705 ( .A(n3180), .B(n2899), .Z(out[419]) );
  ANDN U4706 ( .B(n2901), .A(n2900), .Z(n2902) );
  XNOR U4707 ( .A(n2903), .B(n2902), .Z(out[41]) );
  XNOR U4708 ( .A(in[469]), .B(n3654), .Z(n3182) );
  NOR U4709 ( .A(n3028), .B(n3415), .Z(n2904) );
  XNOR U4710 ( .A(n3182), .B(n2904), .Z(out[420]) );
  XNOR U4711 ( .A(in[470]), .B(n3658), .Z(n3184) );
  NOR U4712 ( .A(n3030), .B(n3419), .Z(n2905) );
  XNOR U4713 ( .A(n3184), .B(n2905), .Z(out[421]) );
  XNOR U4714 ( .A(in[471]), .B(n3662), .Z(n3190) );
  NOR U4715 ( .A(n3032), .B(n3423), .Z(n2906) );
  XNOR U4716 ( .A(n3190), .B(n2906), .Z(out[422]) );
  XNOR U4717 ( .A(in[472]), .B(n3670), .Z(n3192) );
  NOR U4718 ( .A(n3034), .B(n3427), .Z(n2907) );
  XNOR U4719 ( .A(n3192), .B(n2907), .Z(out[423]) );
  XNOR U4720 ( .A(in[473]), .B(n3674), .Z(n3194) );
  NOR U4721 ( .A(n3036), .B(n3431), .Z(n2908) );
  XNOR U4722 ( .A(n3194), .B(n2908), .Z(out[424]) );
  XNOR U4723 ( .A(in[474]), .B(n3678), .Z(n3196) );
  NOR U4724 ( .A(n3038), .B(n3435), .Z(n2909) );
  XNOR U4725 ( .A(n3196), .B(n2909), .Z(out[425]) );
  XNOR U4726 ( .A(in[475]), .B(n3682), .Z(n3198) );
  NOR U4727 ( .A(n3044), .B(n3439), .Z(n2910) );
  XNOR U4728 ( .A(n3198), .B(n2910), .Z(out[426]) );
  XNOR U4729 ( .A(in[476]), .B(n3686), .Z(n3200) );
  NOR U4730 ( .A(n3046), .B(n3443), .Z(n2911) );
  XNOR U4731 ( .A(n3200), .B(n2911), .Z(out[427]) );
  XNOR U4732 ( .A(in[477]), .B(n3690), .Z(n3202) );
  NOR U4733 ( .A(n3048), .B(n3451), .Z(n2912) );
  XNOR U4734 ( .A(n3202), .B(n2912), .Z(out[428]) );
  XNOR U4735 ( .A(in[478]), .B(n3694), .Z(n3204) );
  NOR U4736 ( .A(n3050), .B(n3455), .Z(n2913) );
  XNOR U4737 ( .A(n3204), .B(n2913), .Z(out[429]) );
  ANDN U4738 ( .B(n2915), .A(n2914), .Z(n2916) );
  XNOR U4739 ( .A(n2917), .B(n2916), .Z(out[42]) );
  XNOR U4740 ( .A(in[479]), .B(n3698), .Z(n3206) );
  NOR U4741 ( .A(n3052), .B(n3459), .Z(n2918) );
  XNOR U4742 ( .A(n3206), .B(n2918), .Z(out[430]) );
  XNOR U4743 ( .A(in[480]), .B(n3702), .Z(n3208) );
  NOR U4744 ( .A(n3054), .B(n3463), .Z(n2919) );
  XNOR U4745 ( .A(n3208), .B(n2919), .Z(out[431]) );
  XNOR U4746 ( .A(in[481]), .B(n3706), .Z(n3214) );
  NOR U4747 ( .A(n3056), .B(n3467), .Z(n2920) );
  XNOR U4748 ( .A(n3214), .B(n2920), .Z(out[432]) );
  XNOR U4749 ( .A(in[482]), .B(n3714), .Z(n3216) );
  NOR U4750 ( .A(n3058), .B(n3471), .Z(n2921) );
  XNOR U4751 ( .A(n3216), .B(n2921), .Z(out[433]) );
  XNOR U4752 ( .A(in[483]), .B(n3718), .Z(n3218) );
  NOR U4753 ( .A(n3060), .B(n3475), .Z(n2922) );
  XNOR U4754 ( .A(n3218), .B(n2922), .Z(out[434]) );
  XNOR U4755 ( .A(in[484]), .B(n3722), .Z(n3220) );
  NOR U4756 ( .A(n3062), .B(n3479), .Z(n2923) );
  XNOR U4757 ( .A(n3220), .B(n2923), .Z(out[435]) );
  XNOR U4758 ( .A(in[485]), .B(n3726), .Z(n3222) );
  NOR U4759 ( .A(n3070), .B(n3483), .Z(n2924) );
  XNOR U4760 ( .A(n3222), .B(n2924), .Z(out[436]) );
  XOR U4761 ( .A(in[486]), .B(n3730), .Z(n3224) );
  NOR U4762 ( .A(n3072), .B(n3487), .Z(n2925) );
  XNOR U4763 ( .A(n3224), .B(n2925), .Z(out[437]) );
  XOR U4764 ( .A(in[487]), .B(n3734), .Z(n3226) );
  NOR U4765 ( .A(n3074), .B(n3495), .Z(n2926) );
  XNOR U4766 ( .A(n3226), .B(n2926), .Z(out[438]) );
  XOR U4767 ( .A(in[488]), .B(n3738), .Z(n3228) );
  NOR U4768 ( .A(n3076), .B(n3499), .Z(n2927) );
  XNOR U4769 ( .A(n3228), .B(n2927), .Z(out[439]) );
  ANDN U4770 ( .B(n2929), .A(n2928), .Z(n2930) );
  XNOR U4771 ( .A(n2931), .B(n2930), .Z(out[43]) );
  XOR U4772 ( .A(in[489]), .B(n3742), .Z(n3230) );
  NOR U4773 ( .A(n3078), .B(n3503), .Z(n2932) );
  XNOR U4774 ( .A(n3230), .B(n2932), .Z(out[440]) );
  XOR U4775 ( .A(in[490]), .B(n3746), .Z(n3232) );
  NOR U4776 ( .A(n3080), .B(n3507), .Z(n2933) );
  XNOR U4777 ( .A(n3232), .B(n2933), .Z(out[441]) );
  XOR U4778 ( .A(in[491]), .B(n3750), .Z(n3238) );
  NOR U4779 ( .A(n3082), .B(n3511), .Z(n2934) );
  XNOR U4780 ( .A(n3238), .B(n2934), .Z(out[442]) );
  XOR U4781 ( .A(in[492]), .B(n3758), .Z(n3240) );
  NOR U4782 ( .A(n3084), .B(n3515), .Z(n2935) );
  XNOR U4783 ( .A(n3240), .B(n2935), .Z(out[443]) );
  XOR U4784 ( .A(in[493]), .B(n3762), .Z(n3242) );
  NOR U4785 ( .A(n3086), .B(n3519), .Z(n2936) );
  XNOR U4786 ( .A(n3242), .B(n2936), .Z(out[444]) );
  XOR U4787 ( .A(in[494]), .B(n3766), .Z(n3244) );
  NOR U4788 ( .A(n3088), .B(n3523), .Z(n2937) );
  XNOR U4789 ( .A(n3244), .B(n2937), .Z(out[445]) );
  XOR U4790 ( .A(in[495]), .B(n3770), .Z(n3246) );
  NOR U4791 ( .A(n3094), .B(n3527), .Z(n2938) );
  XNOR U4792 ( .A(n3246), .B(n2938), .Z(out[446]) );
  XOR U4793 ( .A(in[496]), .B(n3774), .Z(n3248) );
  NOR U4794 ( .A(n3096), .B(n3531), .Z(n2939) );
  XNOR U4795 ( .A(n3248), .B(n2939), .Z(out[447]) );
  XNOR U4796 ( .A(in[886]), .B(n3777), .Z(n3251) );
  NAND U4797 ( .A(n3098), .B(n2940), .Z(n2941) );
  XNOR U4798 ( .A(n3251), .B(n2941), .Z(out[448]) );
  XNOR U4799 ( .A(in[887]), .B(n3781), .Z(n3255) );
  NAND U4800 ( .A(n3100), .B(n2942), .Z(n2943) );
  XNOR U4801 ( .A(n3255), .B(n2943), .Z(out[449]) );
  ANDN U4802 ( .B(n2945), .A(n2944), .Z(n2946) );
  XNOR U4803 ( .A(n2947), .B(n2946), .Z(out[44]) );
  XNOR U4804 ( .A(in[888]), .B(n3785), .Z(n3259) );
  NAND U4805 ( .A(n3102), .B(n2948), .Z(n2949) );
  XNOR U4806 ( .A(n3259), .B(n2949), .Z(out[450]) );
  XNOR U4807 ( .A(in[889]), .B(n3789), .Z(n3263) );
  NAND U4808 ( .A(n3104), .B(n2950), .Z(n2951) );
  XNOR U4809 ( .A(n3263), .B(n2951), .Z(out[451]) );
  XNOR U4810 ( .A(in[890]), .B(n3793), .Z(n3271) );
  NAND U4811 ( .A(n3106), .B(n2952), .Z(n2953) );
  XNOR U4812 ( .A(n3271), .B(n2953), .Z(out[452]) );
  XOR U4813 ( .A(in[891]), .B(n3803), .Z(n3275) );
  NAND U4814 ( .A(n3108), .B(n2954), .Z(n2955) );
  XNOR U4815 ( .A(n3275), .B(n2955), .Z(out[453]) );
  XOR U4816 ( .A(in[892]), .B(n3807), .Z(n3279) );
  NAND U4817 ( .A(n3110), .B(n2956), .Z(n2957) );
  XNOR U4818 ( .A(n3279), .B(n2957), .Z(out[454]) );
  XOR U4819 ( .A(in[893]), .B(n3811), .Z(n3283) );
  NAND U4820 ( .A(n3112), .B(n2958), .Z(n2959) );
  XNOR U4821 ( .A(n3283), .B(n2959), .Z(out[455]) );
  XNOR U4822 ( .A(in[894]), .B(n3815), .Z(n3287) );
  NAND U4823 ( .A(n3118), .B(n2960), .Z(n2961) );
  XNOR U4824 ( .A(n3287), .B(n2961), .Z(out[456]) );
  XOR U4825 ( .A(in[895]), .B(n3537), .Z(n3291) );
  NAND U4826 ( .A(n3120), .B(n2962), .Z(n2963) );
  XNOR U4827 ( .A(n3291), .B(n2963), .Z(out[457]) );
  XOR U4828 ( .A(in[832]), .B(n3541), .Z(n3295) );
  NAND U4829 ( .A(n3122), .B(n2964), .Z(n2965) );
  XNOR U4830 ( .A(n3295), .B(n2965), .Z(out[458]) );
  XOR U4831 ( .A(in[833]), .B(n3545), .Z(n3299) );
  NAND U4832 ( .A(n3124), .B(n2966), .Z(n2967) );
  XNOR U4833 ( .A(n3299), .B(n2967), .Z(out[459]) );
  ANDN U4834 ( .B(n2969), .A(n2968), .Z(n2970) );
  XNOR U4835 ( .A(n2971), .B(n2970), .Z(out[45]) );
  XOR U4836 ( .A(in[834]), .B(n3549), .Z(n3303) );
  NAND U4837 ( .A(n3126), .B(n2972), .Z(n2973) );
  XNOR U4838 ( .A(n3303), .B(n2973), .Z(out[460]) );
  XOR U4839 ( .A(in[835]), .B(n3553), .Z(n3307) );
  NAND U4840 ( .A(n3128), .B(n2974), .Z(n2975) );
  XNOR U4841 ( .A(n3307), .B(n2975), .Z(out[461]) );
  XOR U4842 ( .A(in[836]), .B(n3557), .Z(n3315) );
  NAND U4843 ( .A(n3130), .B(n2976), .Z(n2977) );
  XNOR U4844 ( .A(n3315), .B(n2977), .Z(out[462]) );
  XOR U4845 ( .A(in[837]), .B(n3561), .Z(n3319) );
  NAND U4846 ( .A(n3132), .B(n2978), .Z(n2979) );
  XNOR U4847 ( .A(n3319), .B(n2979), .Z(out[463]) );
  XOR U4848 ( .A(in[838]), .B(n3565), .Z(n3323) );
  NAND U4849 ( .A(n3134), .B(n2980), .Z(n2981) );
  XNOR U4850 ( .A(n3323), .B(n2981), .Z(out[464]) );
  XOR U4851 ( .A(in[839]), .B(n3569), .Z(n3327) );
  NAND U4852 ( .A(n3136), .B(n2982), .Z(n2983) );
  XNOR U4853 ( .A(n3327), .B(n2983), .Z(out[465]) );
  XOR U4854 ( .A(in[840]), .B(n3573), .Z(n3331) );
  NAND U4855 ( .A(n3142), .B(n2984), .Z(n2985) );
  XNOR U4856 ( .A(n3331), .B(n2985), .Z(out[466]) );
  XOR U4857 ( .A(in[841]), .B(n3581), .Z(n3335) );
  NAND U4858 ( .A(n3144), .B(n2986), .Z(n2987) );
  XNOR U4859 ( .A(n3335), .B(n2987), .Z(out[467]) );
  XOR U4860 ( .A(in[842]), .B(n3585), .Z(n3339) );
  NAND U4861 ( .A(n3146), .B(n2988), .Z(n2989) );
  XNOR U4862 ( .A(n3339), .B(n2989), .Z(out[468]) );
  XOR U4863 ( .A(in[843]), .B(n3589), .Z(n3343) );
  NAND U4864 ( .A(n3148), .B(n2990), .Z(n2991) );
  XNOR U4865 ( .A(n3343), .B(n2991), .Z(out[469]) );
  ANDN U4866 ( .B(n2993), .A(n2992), .Z(n2994) );
  XNOR U4867 ( .A(n2995), .B(n2994), .Z(out[46]) );
  XOR U4868 ( .A(in[844]), .B(n3593), .Z(n3347) );
  NAND U4869 ( .A(n3150), .B(n2996), .Z(n2997) );
  XNOR U4870 ( .A(n3347), .B(n2997), .Z(out[470]) );
  XOR U4871 ( .A(in[845]), .B(n3597), .Z(n3351) );
  NAND U4872 ( .A(n3152), .B(n2998), .Z(n2999) );
  XNOR U4873 ( .A(n3351), .B(n2999), .Z(out[471]) );
  XOR U4874 ( .A(in[846]), .B(n3601), .Z(n3361) );
  NAND U4875 ( .A(n3154), .B(n3000), .Z(n3001) );
  XNOR U4876 ( .A(n3361), .B(n3001), .Z(out[472]) );
  XOR U4877 ( .A(in[847]), .B(n3605), .Z(n3365) );
  NAND U4878 ( .A(n3156), .B(n3002), .Z(n3003) );
  XNOR U4879 ( .A(n3365), .B(n3003), .Z(out[473]) );
  XOR U4880 ( .A(in[848]), .B(n3609), .Z(n3369) );
  NAND U4881 ( .A(n3158), .B(n3004), .Z(n3005) );
  XNOR U4882 ( .A(n3369), .B(n3005), .Z(out[474]) );
  XOR U4883 ( .A(in[849]), .B(n3613), .Z(n3373) );
  NAND U4884 ( .A(n3160), .B(n3006), .Z(n3007) );
  XNOR U4885 ( .A(n3373), .B(n3007), .Z(out[475]) );
  XOR U4886 ( .A(in[850]), .B(n3617), .Z(n3377) );
  NAND U4887 ( .A(n3166), .B(n3008), .Z(n3009) );
  XNOR U4888 ( .A(n3377), .B(n3009), .Z(out[476]) );
  XNOR U4889 ( .A(in[851]), .B(n3625), .Z(n3381) );
  NAND U4890 ( .A(n3168), .B(n3010), .Z(n3011) );
  XNOR U4891 ( .A(n3381), .B(n3011), .Z(out[477]) );
  XNOR U4892 ( .A(in[852]), .B(n3629), .Z(n3385) );
  NAND U4893 ( .A(n3170), .B(n3012), .Z(n3013) );
  XNOR U4894 ( .A(n3385), .B(n3013), .Z(out[478]) );
  XNOR U4895 ( .A(in[853]), .B(n3633), .Z(n3389) );
  NAND U4896 ( .A(n3172), .B(n3014), .Z(n3015) );
  XNOR U4897 ( .A(n3389), .B(n3015), .Z(out[479]) );
  ANDN U4898 ( .B(n3017), .A(n3016), .Z(n3018) );
  XNOR U4899 ( .A(n3019), .B(n3018), .Z(out[47]) );
  XNOR U4900 ( .A(in[854]), .B(n3637), .Z(n3393) );
  NAND U4901 ( .A(n3174), .B(n3020), .Z(n3021) );
  XNOR U4902 ( .A(n3393), .B(n3021), .Z(out[480]) );
  XNOR U4903 ( .A(in[855]), .B(n3641), .Z(n3397) );
  NAND U4904 ( .A(n3176), .B(n3022), .Z(n3023) );
  XNOR U4905 ( .A(n3397), .B(n3023), .Z(out[481]) );
  XNOR U4906 ( .A(in[856]), .B(n3645), .Z(n3405) );
  NAND U4907 ( .A(n3178), .B(n3024), .Z(n3025) );
  XNOR U4908 ( .A(n3405), .B(n3025), .Z(out[482]) );
  XNOR U4909 ( .A(in[857]), .B(n3649), .Z(n3409) );
  NAND U4910 ( .A(n3180), .B(n3026), .Z(n3027) );
  XNOR U4911 ( .A(n3409), .B(n3027), .Z(out[483]) );
  XNOR U4912 ( .A(in[858]), .B(n3653), .Z(n3413) );
  NAND U4913 ( .A(n3182), .B(n3028), .Z(n3029) );
  XNOR U4914 ( .A(n3413), .B(n3029), .Z(out[484]) );
  XNOR U4915 ( .A(in[859]), .B(n3657), .Z(n3417) );
  NAND U4916 ( .A(n3184), .B(n3030), .Z(n3031) );
  XNOR U4917 ( .A(n3417), .B(n3031), .Z(out[485]) );
  XNOR U4918 ( .A(in[860]), .B(n3661), .Z(n3421) );
  NAND U4919 ( .A(n3190), .B(n3032), .Z(n3033) );
  XNOR U4920 ( .A(n3421), .B(n3033), .Z(out[486]) );
  XNOR U4921 ( .A(in[861]), .B(n3669), .Z(n3425) );
  NAND U4922 ( .A(n3192), .B(n3034), .Z(n3035) );
  XNOR U4923 ( .A(n3425), .B(n3035), .Z(out[487]) );
  XNOR U4924 ( .A(in[862]), .B(n3673), .Z(n3429) );
  NAND U4925 ( .A(n3194), .B(n3036), .Z(n3037) );
  XNOR U4926 ( .A(n3429), .B(n3037), .Z(out[488]) );
  XNOR U4927 ( .A(in[863]), .B(n3677), .Z(n3433) );
  NAND U4928 ( .A(n3196), .B(n3038), .Z(n3039) );
  XNOR U4929 ( .A(n3433), .B(n3039), .Z(out[489]) );
  ANDN U4930 ( .B(n3041), .A(n3040), .Z(n3042) );
  XNOR U4931 ( .A(n3043), .B(n3042), .Z(out[48]) );
  XNOR U4932 ( .A(in[864]), .B(n3681), .Z(n3437) );
  NAND U4933 ( .A(n3198), .B(n3044), .Z(n3045) );
  XNOR U4934 ( .A(n3437), .B(n3045), .Z(out[490]) );
  XNOR U4935 ( .A(in[865]), .B(n3685), .Z(n3441) );
  NAND U4936 ( .A(n3200), .B(n3046), .Z(n3047) );
  XNOR U4937 ( .A(n3441), .B(n3047), .Z(out[491]) );
  XOR U4938 ( .A(n3689), .B(in[866]), .Z(n3449) );
  NAND U4939 ( .A(n3202), .B(n3048), .Z(n3049) );
  XNOR U4940 ( .A(n3449), .B(n3049), .Z(out[492]) );
  XOR U4941 ( .A(n3693), .B(in[867]), .Z(n3453) );
  NAND U4942 ( .A(n3204), .B(n3050), .Z(n3051) );
  XNOR U4943 ( .A(n3453), .B(n3051), .Z(out[493]) );
  XOR U4944 ( .A(n3697), .B(in[868]), .Z(n3457) );
  NAND U4945 ( .A(n3206), .B(n3052), .Z(n3053) );
  XNOR U4946 ( .A(n3457), .B(n3053), .Z(out[494]) );
  XOR U4947 ( .A(n3701), .B(in[869]), .Z(n3461) );
  NAND U4948 ( .A(n3208), .B(n3054), .Z(n3055) );
  XNOR U4949 ( .A(n3461), .B(n3055), .Z(out[495]) );
  XNOR U4950 ( .A(in[870]), .B(n3705), .Z(n3465) );
  NAND U4951 ( .A(n3214), .B(n3056), .Z(n3057) );
  XNOR U4952 ( .A(n3465), .B(n3057), .Z(out[496]) );
  XNOR U4953 ( .A(in[871]), .B(n3713), .Z(n3469) );
  NAND U4954 ( .A(n3216), .B(n3058), .Z(n3059) );
  XNOR U4955 ( .A(n3469), .B(n3059), .Z(out[497]) );
  XNOR U4956 ( .A(in[872]), .B(n3717), .Z(n3473) );
  NAND U4957 ( .A(n3218), .B(n3060), .Z(n3061) );
  XNOR U4958 ( .A(n3473), .B(n3061), .Z(out[498]) );
  XNOR U4959 ( .A(in[873]), .B(n3721), .Z(n3477) );
  NAND U4960 ( .A(n3220), .B(n3062), .Z(n3063) );
  XNOR U4961 ( .A(n3477), .B(n3063), .Z(out[499]) );
  ANDN U4962 ( .B(n3065), .A(n3064), .Z(n3066) );
  XNOR U4963 ( .A(n3067), .B(n3066), .Z(out[49]) );
  OR U4964 ( .A(n3753), .B(n3068), .Z(n3069) );
  XNOR U4965 ( .A(n3752), .B(n3069), .Z(out[4]) );
  XNOR U4966 ( .A(in[874]), .B(n3725), .Z(n3481) );
  NAND U4967 ( .A(n3222), .B(n3070), .Z(n3071) );
  XNOR U4968 ( .A(n3481), .B(n3071), .Z(out[500]) );
  XNOR U4969 ( .A(in[875]), .B(n3729), .Z(n3485) );
  NAND U4970 ( .A(n3224), .B(n3072), .Z(n3073) );
  XNOR U4971 ( .A(n3485), .B(n3073), .Z(out[501]) );
  XNOR U4972 ( .A(in[876]), .B(n3733), .Z(n3493) );
  NAND U4973 ( .A(n3226), .B(n3074), .Z(n3075) );
  XNOR U4974 ( .A(n3493), .B(n3075), .Z(out[502]) );
  XNOR U4975 ( .A(in[877]), .B(n3737), .Z(n3497) );
  NAND U4976 ( .A(n3228), .B(n3076), .Z(n3077) );
  XNOR U4977 ( .A(n3497), .B(n3077), .Z(out[503]) );
  XNOR U4978 ( .A(in[878]), .B(n3741), .Z(n3501) );
  NAND U4979 ( .A(n3230), .B(n3078), .Z(n3079) );
  XNOR U4980 ( .A(n3501), .B(n3079), .Z(out[504]) );
  XNOR U4981 ( .A(in[879]), .B(n3745), .Z(n3505) );
  NAND U4982 ( .A(n3232), .B(n3080), .Z(n3081) );
  XNOR U4983 ( .A(n3505), .B(n3081), .Z(out[505]) );
  XNOR U4984 ( .A(in[880]), .B(n3749), .Z(n3509) );
  NAND U4985 ( .A(n3238), .B(n3082), .Z(n3083) );
  XNOR U4986 ( .A(n3509), .B(n3083), .Z(out[506]) );
  XNOR U4987 ( .A(in[881]), .B(n3757), .Z(n3513) );
  NAND U4988 ( .A(n3240), .B(n3084), .Z(n3085) );
  XNOR U4989 ( .A(n3513), .B(n3085), .Z(out[507]) );
  XNOR U4990 ( .A(in[882]), .B(n3761), .Z(n3517) );
  NAND U4991 ( .A(n3242), .B(n3086), .Z(n3087) );
  XNOR U4992 ( .A(n3517), .B(n3087), .Z(out[508]) );
  XNOR U4993 ( .A(in[883]), .B(n3765), .Z(n3521) );
  NAND U4994 ( .A(n3244), .B(n3088), .Z(n3089) );
  XNOR U4995 ( .A(n3521), .B(n3089), .Z(out[509]) );
  ANDN U4996 ( .B(n3091), .A(n3090), .Z(n3092) );
  XNOR U4997 ( .A(n3093), .B(n3092), .Z(out[50]) );
  XNOR U4998 ( .A(in[884]), .B(n3769), .Z(n3525) );
  NAND U4999 ( .A(n3246), .B(n3094), .Z(n3095) );
  XNOR U5000 ( .A(n3525), .B(n3095), .Z(out[510]) );
  XNOR U5001 ( .A(in[885]), .B(n3773), .Z(n3529) );
  NAND U5002 ( .A(n3248), .B(n3096), .Z(n3097) );
  XNOR U5003 ( .A(n3529), .B(n3097), .Z(out[511]) );
  OR U5004 ( .A(n3251), .B(n3098), .Z(n3099) );
  XNOR U5005 ( .A(n3250), .B(n3099), .Z(out[512]) );
  OR U5006 ( .A(n3255), .B(n3100), .Z(n3101) );
  XNOR U5007 ( .A(n3254), .B(n3101), .Z(out[513]) );
  OR U5008 ( .A(n3259), .B(n3102), .Z(n3103) );
  XNOR U5009 ( .A(n3258), .B(n3103), .Z(out[514]) );
  OR U5010 ( .A(n3263), .B(n3104), .Z(n3105) );
  XNOR U5011 ( .A(n3262), .B(n3105), .Z(out[515]) );
  OR U5012 ( .A(n3271), .B(n3106), .Z(n3107) );
  XNOR U5013 ( .A(n3270), .B(n3107), .Z(out[516]) );
  OR U5014 ( .A(n3275), .B(n3108), .Z(n3109) );
  XNOR U5015 ( .A(n3274), .B(n3109), .Z(out[517]) );
  OR U5016 ( .A(n3279), .B(n3110), .Z(n3111) );
  XNOR U5017 ( .A(n3278), .B(n3111), .Z(out[518]) );
  OR U5018 ( .A(n3283), .B(n3112), .Z(n3113) );
  XNOR U5019 ( .A(n3282), .B(n3113), .Z(out[519]) );
  ANDN U5020 ( .B(n3115), .A(n3114), .Z(n3116) );
  XNOR U5021 ( .A(n3117), .B(n3116), .Z(out[51]) );
  OR U5022 ( .A(n3287), .B(n3118), .Z(n3119) );
  XNOR U5023 ( .A(n3286), .B(n3119), .Z(out[520]) );
  OR U5024 ( .A(n3291), .B(n3120), .Z(n3121) );
  XNOR U5025 ( .A(n3290), .B(n3121), .Z(out[521]) );
  OR U5026 ( .A(n3295), .B(n3122), .Z(n3123) );
  XNOR U5027 ( .A(n3294), .B(n3123), .Z(out[522]) );
  OR U5028 ( .A(n3299), .B(n3124), .Z(n3125) );
  XNOR U5029 ( .A(n3298), .B(n3125), .Z(out[523]) );
  OR U5030 ( .A(n3303), .B(n3126), .Z(n3127) );
  XNOR U5031 ( .A(n3302), .B(n3127), .Z(out[524]) );
  OR U5032 ( .A(n3307), .B(n3128), .Z(n3129) );
  XNOR U5033 ( .A(n3306), .B(n3129), .Z(out[525]) );
  OR U5034 ( .A(n3315), .B(n3130), .Z(n3131) );
  XNOR U5035 ( .A(n3314), .B(n3131), .Z(out[526]) );
  OR U5036 ( .A(n3319), .B(n3132), .Z(n3133) );
  XNOR U5037 ( .A(n3318), .B(n3133), .Z(out[527]) );
  OR U5038 ( .A(n3323), .B(n3134), .Z(n3135) );
  XNOR U5039 ( .A(n3322), .B(n3135), .Z(out[528]) );
  OR U5040 ( .A(n3327), .B(n3136), .Z(n3137) );
  XNOR U5041 ( .A(n3326), .B(n3137), .Z(out[529]) );
  ANDN U5042 ( .B(n3139), .A(n3138), .Z(n3140) );
  XNOR U5043 ( .A(n3141), .B(n3140), .Z(out[52]) );
  OR U5044 ( .A(n3331), .B(n3142), .Z(n3143) );
  XNOR U5045 ( .A(n3330), .B(n3143), .Z(out[530]) );
  OR U5046 ( .A(n3335), .B(n3144), .Z(n3145) );
  XNOR U5047 ( .A(n3334), .B(n3145), .Z(out[531]) );
  OR U5048 ( .A(n3339), .B(n3146), .Z(n3147) );
  XNOR U5049 ( .A(n3338), .B(n3147), .Z(out[532]) );
  OR U5050 ( .A(n3343), .B(n3148), .Z(n3149) );
  XNOR U5051 ( .A(n3342), .B(n3149), .Z(out[533]) );
  OR U5052 ( .A(n3347), .B(n3150), .Z(n3151) );
  XNOR U5053 ( .A(n3346), .B(n3151), .Z(out[534]) );
  OR U5054 ( .A(n3351), .B(n3152), .Z(n3153) );
  XNOR U5055 ( .A(n3350), .B(n3153), .Z(out[535]) );
  OR U5056 ( .A(n3361), .B(n3154), .Z(n3155) );
  XNOR U5057 ( .A(n3360), .B(n3155), .Z(out[536]) );
  OR U5058 ( .A(n3365), .B(n3156), .Z(n3157) );
  XNOR U5059 ( .A(n3364), .B(n3157), .Z(out[537]) );
  OR U5060 ( .A(n3369), .B(n3158), .Z(n3159) );
  XNOR U5061 ( .A(n3368), .B(n3159), .Z(out[538]) );
  OR U5062 ( .A(n3373), .B(n3160), .Z(n3161) );
  XNOR U5063 ( .A(n3372), .B(n3161), .Z(out[539]) );
  ANDN U5064 ( .B(n3163), .A(n3162), .Z(n3164) );
  XNOR U5065 ( .A(n3165), .B(n3164), .Z(out[53]) );
  OR U5066 ( .A(n3377), .B(n3166), .Z(n3167) );
  XNOR U5067 ( .A(n3376), .B(n3167), .Z(out[540]) );
  OR U5068 ( .A(n3381), .B(n3168), .Z(n3169) );
  XNOR U5069 ( .A(n3380), .B(n3169), .Z(out[541]) );
  OR U5070 ( .A(n3385), .B(n3170), .Z(n3171) );
  XNOR U5071 ( .A(n3384), .B(n3171), .Z(out[542]) );
  OR U5072 ( .A(n3389), .B(n3172), .Z(n3173) );
  XNOR U5073 ( .A(n3388), .B(n3173), .Z(out[543]) );
  OR U5074 ( .A(n3393), .B(n3174), .Z(n3175) );
  XNOR U5075 ( .A(n3392), .B(n3175), .Z(out[544]) );
  OR U5076 ( .A(n3397), .B(n3176), .Z(n3177) );
  XNOR U5077 ( .A(n3396), .B(n3177), .Z(out[545]) );
  OR U5078 ( .A(n3405), .B(n3178), .Z(n3179) );
  XNOR U5079 ( .A(n3404), .B(n3179), .Z(out[546]) );
  OR U5080 ( .A(n3409), .B(n3180), .Z(n3181) );
  XNOR U5081 ( .A(n3408), .B(n3181), .Z(out[547]) );
  OR U5082 ( .A(n3413), .B(n3182), .Z(n3183) );
  XNOR U5083 ( .A(n3412), .B(n3183), .Z(out[548]) );
  OR U5084 ( .A(n3417), .B(n3184), .Z(n3185) );
  XNOR U5085 ( .A(n3416), .B(n3185), .Z(out[549]) );
  ANDN U5086 ( .B(n3187), .A(n3186), .Z(n3188) );
  XNOR U5087 ( .A(n3189), .B(n3188), .Z(out[54]) );
  OR U5088 ( .A(n3421), .B(n3190), .Z(n3191) );
  XNOR U5089 ( .A(n3420), .B(n3191), .Z(out[550]) );
  OR U5090 ( .A(n3425), .B(n3192), .Z(n3193) );
  XNOR U5091 ( .A(n3424), .B(n3193), .Z(out[551]) );
  OR U5092 ( .A(n3429), .B(n3194), .Z(n3195) );
  XNOR U5093 ( .A(n3428), .B(n3195), .Z(out[552]) );
  OR U5094 ( .A(n3433), .B(n3196), .Z(n3197) );
  XNOR U5095 ( .A(n3432), .B(n3197), .Z(out[553]) );
  OR U5096 ( .A(n3437), .B(n3198), .Z(n3199) );
  XNOR U5097 ( .A(n3436), .B(n3199), .Z(out[554]) );
  OR U5098 ( .A(n3441), .B(n3200), .Z(n3201) );
  XNOR U5099 ( .A(n3440), .B(n3201), .Z(out[555]) );
  OR U5100 ( .A(n3449), .B(n3202), .Z(n3203) );
  XNOR U5101 ( .A(n3448), .B(n3203), .Z(out[556]) );
  OR U5102 ( .A(n3453), .B(n3204), .Z(n3205) );
  XNOR U5103 ( .A(n3452), .B(n3205), .Z(out[557]) );
  OR U5104 ( .A(n3457), .B(n3206), .Z(n3207) );
  XNOR U5105 ( .A(n3456), .B(n3207), .Z(out[558]) );
  OR U5106 ( .A(n3461), .B(n3208), .Z(n3209) );
  XNOR U5107 ( .A(n3460), .B(n3209), .Z(out[559]) );
  ANDN U5108 ( .B(n3211), .A(n3210), .Z(n3212) );
  XNOR U5109 ( .A(n3213), .B(n3212), .Z(out[55]) );
  OR U5110 ( .A(n3465), .B(n3214), .Z(n3215) );
  XNOR U5111 ( .A(n3464), .B(n3215), .Z(out[560]) );
  OR U5112 ( .A(n3469), .B(n3216), .Z(n3217) );
  XNOR U5113 ( .A(n3468), .B(n3217), .Z(out[561]) );
  OR U5114 ( .A(n3473), .B(n3218), .Z(n3219) );
  XNOR U5115 ( .A(n3472), .B(n3219), .Z(out[562]) );
  OR U5116 ( .A(n3477), .B(n3220), .Z(n3221) );
  XNOR U5117 ( .A(n3476), .B(n3221), .Z(out[563]) );
  OR U5118 ( .A(n3481), .B(n3222), .Z(n3223) );
  XNOR U5119 ( .A(n3480), .B(n3223), .Z(out[564]) );
  OR U5120 ( .A(n3485), .B(n3224), .Z(n3225) );
  XNOR U5121 ( .A(n3484), .B(n3225), .Z(out[565]) );
  OR U5122 ( .A(n3493), .B(n3226), .Z(n3227) );
  XNOR U5123 ( .A(n3492), .B(n3227), .Z(out[566]) );
  OR U5124 ( .A(n3497), .B(n3228), .Z(n3229) );
  XNOR U5125 ( .A(n3496), .B(n3229), .Z(out[567]) );
  OR U5126 ( .A(n3501), .B(n3230), .Z(n3231) );
  XNOR U5127 ( .A(n3500), .B(n3231), .Z(out[568]) );
  OR U5128 ( .A(n3505), .B(n3232), .Z(n3233) );
  XNOR U5129 ( .A(n3504), .B(n3233), .Z(out[569]) );
  ANDN U5130 ( .B(n3235), .A(n3234), .Z(n3236) );
  XNOR U5131 ( .A(n3237), .B(n3236), .Z(out[56]) );
  OR U5132 ( .A(n3509), .B(n3238), .Z(n3239) );
  XNOR U5133 ( .A(n3508), .B(n3239), .Z(out[570]) );
  OR U5134 ( .A(n3513), .B(n3240), .Z(n3241) );
  XNOR U5135 ( .A(n3512), .B(n3241), .Z(out[571]) );
  OR U5136 ( .A(n3517), .B(n3242), .Z(n3243) );
  XNOR U5137 ( .A(n3516), .B(n3243), .Z(out[572]) );
  OR U5138 ( .A(n3521), .B(n3244), .Z(n3245) );
  XNOR U5139 ( .A(n3520), .B(n3245), .Z(out[573]) );
  OR U5140 ( .A(n3525), .B(n3246), .Z(n3247) );
  XNOR U5141 ( .A(n3524), .B(n3247), .Z(out[574]) );
  OR U5142 ( .A(n3529), .B(n3248), .Z(n3249) );
  XNOR U5143 ( .A(n3528), .B(n3249), .Z(out[575]) );
  ANDN U5144 ( .B(n3251), .A(n3250), .Z(n3252) );
  XNOR U5145 ( .A(n3253), .B(n3252), .Z(out[576]) );
  ANDN U5146 ( .B(n3255), .A(n3254), .Z(n3256) );
  XNOR U5147 ( .A(n3257), .B(n3256), .Z(out[577]) );
  ANDN U5148 ( .B(n3259), .A(n3258), .Z(n3260) );
  XNOR U5149 ( .A(n3261), .B(n3260), .Z(out[578]) );
  ANDN U5150 ( .B(n3263), .A(n3262), .Z(n3264) );
  XNOR U5151 ( .A(n3265), .B(n3264), .Z(out[579]) );
  ANDN U5152 ( .B(n3267), .A(n3266), .Z(n3268) );
  XNOR U5153 ( .A(n3269), .B(n3268), .Z(out[57]) );
  ANDN U5154 ( .B(n3271), .A(n3270), .Z(n3272) );
  XNOR U5155 ( .A(n3273), .B(n3272), .Z(out[580]) );
  ANDN U5156 ( .B(n3275), .A(n3274), .Z(n3276) );
  XNOR U5157 ( .A(n3277), .B(n3276), .Z(out[581]) );
  ANDN U5158 ( .B(n3279), .A(n3278), .Z(n3280) );
  XNOR U5159 ( .A(n3281), .B(n3280), .Z(out[582]) );
  ANDN U5160 ( .B(n3283), .A(n3282), .Z(n3284) );
  XNOR U5161 ( .A(n3285), .B(n3284), .Z(out[583]) );
  ANDN U5162 ( .B(n3287), .A(n3286), .Z(n3288) );
  XNOR U5163 ( .A(n3289), .B(n3288), .Z(out[584]) );
  ANDN U5164 ( .B(n3291), .A(n3290), .Z(n3292) );
  XNOR U5165 ( .A(n3293), .B(n3292), .Z(out[585]) );
  ANDN U5166 ( .B(n3295), .A(n3294), .Z(n3296) );
  XNOR U5167 ( .A(n3297), .B(n3296), .Z(out[586]) );
  ANDN U5168 ( .B(n3299), .A(n3298), .Z(n3300) );
  XNOR U5169 ( .A(n3301), .B(n3300), .Z(out[587]) );
  ANDN U5170 ( .B(n3303), .A(n3302), .Z(n3304) );
  XNOR U5171 ( .A(n3305), .B(n3304), .Z(out[588]) );
  ANDN U5172 ( .B(n3307), .A(n3306), .Z(n3308) );
  XNOR U5173 ( .A(n3309), .B(n3308), .Z(out[589]) );
  ANDN U5174 ( .B(n3311), .A(n3310), .Z(n3312) );
  XNOR U5175 ( .A(n3313), .B(n3312), .Z(out[58]) );
  ANDN U5176 ( .B(n3315), .A(n3314), .Z(n3316) );
  XNOR U5177 ( .A(n3317), .B(n3316), .Z(out[590]) );
  ANDN U5178 ( .B(n3319), .A(n3318), .Z(n3320) );
  XNOR U5179 ( .A(n3321), .B(n3320), .Z(out[591]) );
  ANDN U5180 ( .B(n3323), .A(n3322), .Z(n3324) );
  XNOR U5181 ( .A(n3325), .B(n3324), .Z(out[592]) );
  ANDN U5182 ( .B(n3327), .A(n3326), .Z(n3328) );
  XNOR U5183 ( .A(n3329), .B(n3328), .Z(out[593]) );
  ANDN U5184 ( .B(n3331), .A(n3330), .Z(n3332) );
  XNOR U5185 ( .A(n3333), .B(n3332), .Z(out[594]) );
  ANDN U5186 ( .B(n3335), .A(n3334), .Z(n3336) );
  XNOR U5187 ( .A(n3337), .B(n3336), .Z(out[595]) );
  ANDN U5188 ( .B(n3339), .A(n3338), .Z(n3340) );
  XNOR U5189 ( .A(n3341), .B(n3340), .Z(out[596]) );
  ANDN U5190 ( .B(n3343), .A(n3342), .Z(n3344) );
  XNOR U5191 ( .A(n3345), .B(n3344), .Z(out[597]) );
  ANDN U5192 ( .B(n3347), .A(n3346), .Z(n3348) );
  XNOR U5193 ( .A(n3349), .B(n3348), .Z(out[598]) );
  ANDN U5194 ( .B(n3351), .A(n3350), .Z(n3352) );
  XNOR U5195 ( .A(n3353), .B(n3352), .Z(out[599]) );
  ANDN U5196 ( .B(n3355), .A(n3354), .Z(n3356) );
  XNOR U5197 ( .A(n3357), .B(n3356), .Z(out[59]) );
  OR U5198 ( .A(n3797), .B(n3358), .Z(n3359) );
  XNOR U5199 ( .A(n3796), .B(n3359), .Z(out[5]) );
  ANDN U5200 ( .B(n3361), .A(n3360), .Z(n3362) );
  XNOR U5201 ( .A(n3363), .B(n3362), .Z(out[600]) );
  ANDN U5202 ( .B(n3365), .A(n3364), .Z(n3366) );
  XNOR U5203 ( .A(n3367), .B(n3366), .Z(out[601]) );
  ANDN U5204 ( .B(n3369), .A(n3368), .Z(n3370) );
  XNOR U5205 ( .A(n3371), .B(n3370), .Z(out[602]) );
  ANDN U5206 ( .B(n3373), .A(n3372), .Z(n3374) );
  XNOR U5207 ( .A(n3375), .B(n3374), .Z(out[603]) );
  ANDN U5208 ( .B(n3377), .A(n3376), .Z(n3378) );
  XNOR U5209 ( .A(n3379), .B(n3378), .Z(out[604]) );
  ANDN U5210 ( .B(n3381), .A(n3380), .Z(n3382) );
  XNOR U5211 ( .A(n3383), .B(n3382), .Z(out[605]) );
  ANDN U5212 ( .B(n3385), .A(n3384), .Z(n3386) );
  XNOR U5213 ( .A(n3387), .B(n3386), .Z(out[606]) );
  ANDN U5214 ( .B(n3389), .A(n3388), .Z(n3390) );
  XNOR U5215 ( .A(n3391), .B(n3390), .Z(out[607]) );
  ANDN U5216 ( .B(n3393), .A(n3392), .Z(n3394) );
  XNOR U5217 ( .A(n3395), .B(n3394), .Z(out[608]) );
  ANDN U5218 ( .B(n3397), .A(n3396), .Z(n3398) );
  XNOR U5219 ( .A(n3399), .B(n3398), .Z(out[609]) );
  ANDN U5220 ( .B(n3401), .A(n3400), .Z(n3402) );
  XNOR U5221 ( .A(n3403), .B(n3402), .Z(out[60]) );
  ANDN U5222 ( .B(n3405), .A(n3404), .Z(n3406) );
  XNOR U5223 ( .A(n3407), .B(n3406), .Z(out[610]) );
  ANDN U5224 ( .B(n3409), .A(n3408), .Z(n3410) );
  XNOR U5225 ( .A(n3411), .B(n3410), .Z(out[611]) );
  ANDN U5226 ( .B(n3413), .A(n3412), .Z(n3414) );
  XNOR U5227 ( .A(n3415), .B(n3414), .Z(out[612]) );
  ANDN U5228 ( .B(n3417), .A(n3416), .Z(n3418) );
  XNOR U5229 ( .A(n3419), .B(n3418), .Z(out[613]) );
  ANDN U5230 ( .B(n3421), .A(n3420), .Z(n3422) );
  XNOR U5231 ( .A(n3423), .B(n3422), .Z(out[614]) );
  ANDN U5232 ( .B(n3425), .A(n3424), .Z(n3426) );
  XNOR U5233 ( .A(n3427), .B(n3426), .Z(out[615]) );
  ANDN U5234 ( .B(n3429), .A(n3428), .Z(n3430) );
  XNOR U5235 ( .A(n3431), .B(n3430), .Z(out[616]) );
  ANDN U5236 ( .B(n3433), .A(n3432), .Z(n3434) );
  XNOR U5237 ( .A(n3435), .B(n3434), .Z(out[617]) );
  ANDN U5238 ( .B(n3437), .A(n3436), .Z(n3438) );
  XNOR U5239 ( .A(n3439), .B(n3438), .Z(out[618]) );
  ANDN U5240 ( .B(n3441), .A(n3440), .Z(n3442) );
  XNOR U5241 ( .A(n3443), .B(n3442), .Z(out[619]) );
  ANDN U5242 ( .B(n3445), .A(n3444), .Z(n3446) );
  XNOR U5243 ( .A(n3447), .B(n3446), .Z(out[61]) );
  ANDN U5244 ( .B(n3449), .A(n3448), .Z(n3450) );
  XNOR U5245 ( .A(n3451), .B(n3450), .Z(out[620]) );
  ANDN U5246 ( .B(n3453), .A(n3452), .Z(n3454) );
  XNOR U5247 ( .A(n3455), .B(n3454), .Z(out[621]) );
  ANDN U5248 ( .B(n3457), .A(n3456), .Z(n3458) );
  XNOR U5249 ( .A(n3459), .B(n3458), .Z(out[622]) );
  ANDN U5250 ( .B(n3461), .A(n3460), .Z(n3462) );
  XNOR U5251 ( .A(n3463), .B(n3462), .Z(out[623]) );
  ANDN U5252 ( .B(n3465), .A(n3464), .Z(n3466) );
  XNOR U5253 ( .A(n3467), .B(n3466), .Z(out[624]) );
  ANDN U5254 ( .B(n3469), .A(n3468), .Z(n3470) );
  XNOR U5255 ( .A(n3471), .B(n3470), .Z(out[625]) );
  ANDN U5256 ( .B(n3473), .A(n3472), .Z(n3474) );
  XNOR U5257 ( .A(n3475), .B(n3474), .Z(out[626]) );
  ANDN U5258 ( .B(n3477), .A(n3476), .Z(n3478) );
  XNOR U5259 ( .A(n3479), .B(n3478), .Z(out[627]) );
  ANDN U5260 ( .B(n3481), .A(n3480), .Z(n3482) );
  XNOR U5261 ( .A(n3483), .B(n3482), .Z(out[628]) );
  ANDN U5262 ( .B(n3485), .A(n3484), .Z(n3486) );
  XNOR U5263 ( .A(n3487), .B(n3486), .Z(out[629]) );
  ANDN U5264 ( .B(n3489), .A(n3488), .Z(n3490) );
  XNOR U5265 ( .A(n3491), .B(n3490), .Z(out[62]) );
  ANDN U5266 ( .B(n3493), .A(n3492), .Z(n3494) );
  XNOR U5267 ( .A(n3495), .B(n3494), .Z(out[630]) );
  ANDN U5268 ( .B(n3497), .A(n3496), .Z(n3498) );
  XNOR U5269 ( .A(n3499), .B(n3498), .Z(out[631]) );
  ANDN U5270 ( .B(n3501), .A(n3500), .Z(n3502) );
  XNOR U5271 ( .A(n3503), .B(n3502), .Z(out[632]) );
  ANDN U5272 ( .B(n3505), .A(n3504), .Z(n3506) );
  XNOR U5273 ( .A(n3507), .B(n3506), .Z(out[633]) );
  ANDN U5274 ( .B(n3509), .A(n3508), .Z(n3510) );
  XNOR U5275 ( .A(n3511), .B(n3510), .Z(out[634]) );
  ANDN U5276 ( .B(n3513), .A(n3512), .Z(n3514) );
  XNOR U5277 ( .A(n3515), .B(n3514), .Z(out[635]) );
  ANDN U5278 ( .B(n3517), .A(n3516), .Z(n3518) );
  XNOR U5279 ( .A(n3519), .B(n3518), .Z(out[636]) );
  ANDN U5280 ( .B(n3521), .A(n3520), .Z(n3522) );
  XNOR U5281 ( .A(n3523), .B(n3522), .Z(out[637]) );
  ANDN U5282 ( .B(n3525), .A(n3524), .Z(n3526) );
  XNOR U5283 ( .A(n3527), .B(n3526), .Z(out[638]) );
  ANDN U5284 ( .B(n3529), .A(n3528), .Z(n3530) );
  XNOR U5285 ( .A(n3531), .B(n3530), .Z(out[639]) );
  ANDN U5286 ( .B(n3533), .A(n3532), .Z(n3534) );
  XNOR U5287 ( .A(n3535), .B(n3534), .Z(out[63]) );
  XNOR U5288 ( .A(in[302]), .B(n3536), .Z(n3965) );
  XNOR U5289 ( .A(in[1535]), .B(n3537), .Z(n4343) );
  XNOR U5290 ( .A(in[1146]), .B(n3538), .Z(n4340) );
  NAND U5291 ( .A(n4343), .B(n4340), .Z(n3539) );
  XNOR U5292 ( .A(n3965), .B(n3539), .Z(out[640]) );
  XNOR U5293 ( .A(in[303]), .B(n3540), .Z(n3968) );
  XNOR U5294 ( .A(in[1472]), .B(n3541), .Z(n4347) );
  XNOR U5295 ( .A(in[1147]), .B(n3542), .Z(n4344) );
  NAND U5296 ( .A(n4347), .B(n4344), .Z(n3543) );
  XNOR U5297 ( .A(n3968), .B(n3543), .Z(out[641]) );
  XNOR U5298 ( .A(in[304]), .B(n3544), .Z(n3975) );
  XNOR U5299 ( .A(in[1473]), .B(n3545), .Z(n4351) );
  XNOR U5300 ( .A(in[1148]), .B(n3546), .Z(n4348) );
  NAND U5301 ( .A(n4351), .B(n4348), .Z(n3547) );
  XNOR U5302 ( .A(n3975), .B(n3547), .Z(out[642]) );
  XNOR U5303 ( .A(in[305]), .B(n3548), .Z(n3978) );
  XNOR U5304 ( .A(in[1474]), .B(n3549), .Z(n4355) );
  XNOR U5305 ( .A(in[1149]), .B(n3550), .Z(n4352) );
  NAND U5306 ( .A(n4355), .B(n4352), .Z(n3551) );
  XNOR U5307 ( .A(n3978), .B(n3551), .Z(out[643]) );
  XNOR U5308 ( .A(in[306]), .B(n3552), .Z(n3981) );
  XNOR U5309 ( .A(in[1475]), .B(n3553), .Z(n4367) );
  XNOR U5310 ( .A(in[1150]), .B(n3554), .Z(n4364) );
  NAND U5311 ( .A(n4367), .B(n4364), .Z(n3555) );
  XNOR U5312 ( .A(n3981), .B(n3555), .Z(out[644]) );
  XNOR U5313 ( .A(in[307]), .B(n3556), .Z(n3984) );
  XNOR U5314 ( .A(in[1476]), .B(n3557), .Z(n4371) );
  XNOR U5315 ( .A(in[1151]), .B(n3558), .Z(n4368) );
  NAND U5316 ( .A(n4371), .B(n4368), .Z(n3559) );
  XNOR U5317 ( .A(n3984), .B(n3559), .Z(out[645]) );
  XNOR U5318 ( .A(in[308]), .B(n3560), .Z(n3987) );
  XNOR U5319 ( .A(in[1477]), .B(n3561), .Z(n4375) );
  XNOR U5320 ( .A(in[1088]), .B(n3562), .Z(n4372) );
  NAND U5321 ( .A(n4375), .B(n4372), .Z(n3563) );
  XNOR U5322 ( .A(n3987), .B(n3563), .Z(out[646]) );
  XNOR U5323 ( .A(in[309]), .B(n3564), .Z(n3990) );
  XNOR U5324 ( .A(in[1478]), .B(n3565), .Z(n4379) );
  XNOR U5325 ( .A(in[1089]), .B(n3566), .Z(n4376) );
  NAND U5326 ( .A(n4379), .B(n4376), .Z(n3567) );
  XNOR U5327 ( .A(n3990), .B(n3567), .Z(out[647]) );
  XNOR U5328 ( .A(in[310]), .B(n3568), .Z(n3993) );
  XNOR U5329 ( .A(in[1479]), .B(n3569), .Z(n4383) );
  XOR U5330 ( .A(n3570), .B(in[1090]), .Z(n4380) );
  NAND U5331 ( .A(n4383), .B(n4380), .Z(n3571) );
  XNOR U5332 ( .A(n3993), .B(n3571), .Z(out[648]) );
  XNOR U5333 ( .A(in[311]), .B(n3572), .Z(n3996) );
  XNOR U5334 ( .A(in[1480]), .B(n3573), .Z(n4387) );
  XOR U5335 ( .A(n3574), .B(in[1091]), .Z(n4384) );
  NAND U5336 ( .A(n4387), .B(n4384), .Z(n3575) );
  XNOR U5337 ( .A(n3996), .B(n3575), .Z(out[649]) );
  NOR U5338 ( .A(n3577), .B(n3576), .Z(n3578) );
  XNOR U5339 ( .A(n3579), .B(n3578), .Z(out[64]) );
  XNOR U5340 ( .A(in[312]), .B(n3580), .Z(n3999) );
  XNOR U5341 ( .A(in[1481]), .B(n3581), .Z(n4391) );
  XOR U5342 ( .A(n3582), .B(in[1092]), .Z(n4388) );
  NAND U5343 ( .A(n4391), .B(n4388), .Z(n3583) );
  XNOR U5344 ( .A(n3999), .B(n3583), .Z(out[650]) );
  XNOR U5345 ( .A(in[313]), .B(n3584), .Z(n4002) );
  XNOR U5346 ( .A(in[1482]), .B(n3585), .Z(n4395) );
  XOR U5347 ( .A(n3586), .B(in[1093]), .Z(n4392) );
  NAND U5348 ( .A(n4395), .B(n4392), .Z(n3587) );
  XNOR U5349 ( .A(n4002), .B(n3587), .Z(out[651]) );
  XNOR U5350 ( .A(in[314]), .B(n3588), .Z(n4009) );
  XNOR U5351 ( .A(in[1483]), .B(n3589), .Z(n4399) );
  XOR U5352 ( .A(n3590), .B(in[1094]), .Z(n4396) );
  NAND U5353 ( .A(n4399), .B(n4396), .Z(n3591) );
  XNOR U5354 ( .A(n4009), .B(n3591), .Z(out[652]) );
  XNOR U5355 ( .A(in[315]), .B(n3592), .Z(n4012) );
  XNOR U5356 ( .A(in[1484]), .B(n3593), .Z(n4403) );
  XOR U5357 ( .A(n3594), .B(in[1095]), .Z(n4400) );
  NAND U5358 ( .A(n4403), .B(n4400), .Z(n3595) );
  XNOR U5359 ( .A(n4012), .B(n3595), .Z(out[653]) );
  XNOR U5360 ( .A(in[316]), .B(n3596), .Z(n4015) );
  XNOR U5361 ( .A(in[1485]), .B(n3597), .Z(n4411) );
  XOR U5362 ( .A(n3598), .B(in[1096]), .Z(n4408) );
  NAND U5363 ( .A(n4411), .B(n4408), .Z(n3599) );
  XNOR U5364 ( .A(n4015), .B(n3599), .Z(out[654]) );
  XNOR U5365 ( .A(in[317]), .B(n3600), .Z(n4018) );
  XNOR U5366 ( .A(in[1486]), .B(n3601), .Z(n4415) );
  XOR U5367 ( .A(in[1097]), .B(n3602), .Z(n4412) );
  NAND U5368 ( .A(n4415), .B(n4412), .Z(n3603) );
  XNOR U5369 ( .A(n4018), .B(n3603), .Z(out[655]) );
  XNOR U5370 ( .A(in[318]), .B(n3604), .Z(n4021) );
  XNOR U5371 ( .A(in[1487]), .B(n3605), .Z(n4419) );
  XOR U5372 ( .A(n3606), .B(in[1098]), .Z(n4416) );
  NAND U5373 ( .A(n4419), .B(n4416), .Z(n3607) );
  XNOR U5374 ( .A(n4021), .B(n3607), .Z(out[656]) );
  XNOR U5375 ( .A(in[319]), .B(n3608), .Z(n4024) );
  XNOR U5376 ( .A(in[1488]), .B(n3609), .Z(n4423) );
  XOR U5377 ( .A(n3610), .B(in[1099]), .Z(n4420) );
  NAND U5378 ( .A(n4423), .B(n4420), .Z(n3611) );
  XNOR U5379 ( .A(n4024), .B(n3611), .Z(out[657]) );
  XNOR U5380 ( .A(in[256]), .B(n3612), .Z(n4027) );
  XNOR U5381 ( .A(in[1489]), .B(n3613), .Z(n4427) );
  XOR U5382 ( .A(in[1100]), .B(n3614), .Z(n4424) );
  NAND U5383 ( .A(n4427), .B(n4424), .Z(n3615) );
  XNOR U5384 ( .A(n4027), .B(n3615), .Z(out[658]) );
  XNOR U5385 ( .A(in[257]), .B(n3616), .Z(n4030) );
  XNOR U5386 ( .A(in[1490]), .B(n3617), .Z(n4431) );
  XOR U5387 ( .A(in[1101]), .B(n3618), .Z(n4428) );
  NAND U5388 ( .A(n4431), .B(n4428), .Z(n3619) );
  XNOR U5389 ( .A(n4030), .B(n3619), .Z(out[659]) );
  NOR U5390 ( .A(n3621), .B(n3620), .Z(n3622) );
  XNOR U5391 ( .A(n3623), .B(n3622), .Z(out[65]) );
  XNOR U5392 ( .A(in[258]), .B(n3624), .Z(n4033) );
  XOR U5393 ( .A(in[1491]), .B(n3625), .Z(n4435) );
  XOR U5394 ( .A(in[1102]), .B(n3626), .Z(n4432) );
  NAND U5395 ( .A(n4435), .B(n4432), .Z(n3627) );
  XNOR U5396 ( .A(n4033), .B(n3627), .Z(out[660]) );
  XNOR U5397 ( .A(in[259]), .B(n3628), .Z(n4036) );
  XOR U5398 ( .A(in[1492]), .B(n3629), .Z(n4439) );
  XOR U5399 ( .A(in[1103]), .B(n3630), .Z(n4436) );
  NAND U5400 ( .A(n4439), .B(n4436), .Z(n3631) );
  XNOR U5401 ( .A(n4036), .B(n3631), .Z(out[661]) );
  XOR U5402 ( .A(in[260]), .B(n3632), .Z(n4043) );
  XOR U5403 ( .A(in[1493]), .B(n3633), .Z(n4443) );
  XOR U5404 ( .A(in[1104]), .B(n3634), .Z(n4440) );
  NAND U5405 ( .A(n4443), .B(n4440), .Z(n3635) );
  XNOR U5406 ( .A(n4043), .B(n3635), .Z(out[662]) );
  XOR U5407 ( .A(in[261]), .B(n3636), .Z(n4046) );
  XOR U5408 ( .A(in[1494]), .B(n3637), .Z(n4447) );
  XOR U5409 ( .A(in[1105]), .B(n3638), .Z(n4444) );
  NAND U5410 ( .A(n4447), .B(n4444), .Z(n3639) );
  XNOR U5411 ( .A(n4046), .B(n3639), .Z(out[663]) );
  XOR U5412 ( .A(in[262]), .B(n3640), .Z(n4049) );
  XOR U5413 ( .A(in[1495]), .B(n3641), .Z(n4455) );
  XOR U5414 ( .A(in[1106]), .B(n3642), .Z(n4452) );
  NAND U5415 ( .A(n4455), .B(n4452), .Z(n3643) );
  XNOR U5416 ( .A(n4049), .B(n3643), .Z(out[664]) );
  XOR U5417 ( .A(in[263]), .B(n3644), .Z(n4052) );
  XOR U5418 ( .A(in[1496]), .B(n3645), .Z(n4459) );
  XOR U5419 ( .A(in[1107]), .B(n3646), .Z(n4456) );
  NAND U5420 ( .A(n4459), .B(n4456), .Z(n3647) );
  XNOR U5421 ( .A(n4052), .B(n3647), .Z(out[665]) );
  XOR U5422 ( .A(in[264]), .B(n3648), .Z(n4055) );
  XOR U5423 ( .A(in[1497]), .B(n3649), .Z(n4463) );
  XOR U5424 ( .A(in[1108]), .B(n3650), .Z(n4460) );
  NAND U5425 ( .A(n4463), .B(n4460), .Z(n3651) );
  XNOR U5426 ( .A(n4055), .B(n3651), .Z(out[666]) );
  XOR U5427 ( .A(in[265]), .B(n3652), .Z(n4058) );
  XOR U5428 ( .A(in[1498]), .B(n3653), .Z(n4467) );
  XOR U5429 ( .A(in[1109]), .B(n3654), .Z(n4464) );
  NAND U5430 ( .A(n4467), .B(n4464), .Z(n3655) );
  XNOR U5431 ( .A(n4058), .B(n3655), .Z(out[667]) );
  XOR U5432 ( .A(in[266]), .B(n3656), .Z(n4061) );
  XOR U5433 ( .A(in[1499]), .B(n3657), .Z(n4471) );
  XOR U5434 ( .A(in[1110]), .B(n3658), .Z(n4468) );
  NAND U5435 ( .A(n4471), .B(n4468), .Z(n3659) );
  XNOR U5436 ( .A(n4061), .B(n3659), .Z(out[668]) );
  XOR U5437 ( .A(in[267]), .B(n3660), .Z(n4064) );
  XOR U5438 ( .A(in[1500]), .B(n3661), .Z(n4475) );
  XOR U5439 ( .A(in[1111]), .B(n3662), .Z(n4472) );
  NAND U5440 ( .A(n4475), .B(n4472), .Z(n3663) );
  XNOR U5441 ( .A(n4064), .B(n3663), .Z(out[669]) );
  ANDN U5442 ( .B(n3665), .A(n3664), .Z(n3666) );
  XNOR U5443 ( .A(n3667), .B(n3666), .Z(out[66]) );
  XOR U5444 ( .A(in[268]), .B(n3668), .Z(n4067) );
  XOR U5445 ( .A(in[1501]), .B(n3669), .Z(n4479) );
  XOR U5446 ( .A(in[1112]), .B(n3670), .Z(n4476) );
  NAND U5447 ( .A(n4479), .B(n4476), .Z(n3671) );
  XNOR U5448 ( .A(n4067), .B(n3671), .Z(out[670]) );
  XOR U5449 ( .A(in[269]), .B(n3672), .Z(n4070) );
  XOR U5450 ( .A(in[1502]), .B(n3673), .Z(n4483) );
  XOR U5451 ( .A(in[1113]), .B(n3674), .Z(n4480) );
  NAND U5452 ( .A(n4483), .B(n4480), .Z(n3675) );
  XNOR U5453 ( .A(n4070), .B(n3675), .Z(out[671]) );
  XOR U5454 ( .A(in[270]), .B(n3676), .Z(n4081) );
  XOR U5455 ( .A(in[1503]), .B(n3677), .Z(n4487) );
  XOR U5456 ( .A(in[1114]), .B(n3678), .Z(n4484) );
  NAND U5457 ( .A(n4487), .B(n4484), .Z(n3679) );
  XNOR U5458 ( .A(n4081), .B(n3679), .Z(out[672]) );
  XOR U5459 ( .A(in[271]), .B(n3680), .Z(n4084) );
  XOR U5460 ( .A(in[1504]), .B(n3681), .Z(n4491) );
  XOR U5461 ( .A(in[1115]), .B(n3682), .Z(n4488) );
  NAND U5462 ( .A(n4491), .B(n4488), .Z(n3683) );
  XNOR U5463 ( .A(n4084), .B(n3683), .Z(out[673]) );
  XOR U5464 ( .A(in[272]), .B(n3684), .Z(n4087) );
  XOR U5465 ( .A(in[1505]), .B(n3685), .Z(n4499) );
  XOR U5466 ( .A(in[1116]), .B(n3686), .Z(n4496) );
  NAND U5467 ( .A(n4499), .B(n4496), .Z(n3687) );
  XNOR U5468 ( .A(n4087), .B(n3687), .Z(out[674]) );
  XOR U5469 ( .A(in[273]), .B(n3688), .Z(n4090) );
  XNOR U5470 ( .A(n3689), .B(in[1506]), .Z(n4503) );
  XOR U5471 ( .A(in[1117]), .B(n3690), .Z(n4500) );
  NAND U5472 ( .A(n4503), .B(n4500), .Z(n3691) );
  XNOR U5473 ( .A(n4090), .B(n3691), .Z(out[675]) );
  XOR U5474 ( .A(in[274]), .B(n3692), .Z(n4093) );
  XNOR U5475 ( .A(n3693), .B(in[1507]), .Z(n4507) );
  XOR U5476 ( .A(in[1118]), .B(n3694), .Z(n4504) );
  NAND U5477 ( .A(n4507), .B(n4504), .Z(n3695) );
  XNOR U5478 ( .A(n4093), .B(n3695), .Z(out[676]) );
  XOR U5479 ( .A(in[275]), .B(n3696), .Z(n4096) );
  XNOR U5480 ( .A(n3697), .B(in[1508]), .Z(n4511) );
  XOR U5481 ( .A(in[1119]), .B(n3698), .Z(n4508) );
  NAND U5482 ( .A(n4511), .B(n4508), .Z(n3699) );
  XNOR U5483 ( .A(n4096), .B(n3699), .Z(out[677]) );
  XOR U5484 ( .A(in[276]), .B(n3700), .Z(n4099) );
  XNOR U5485 ( .A(n3701), .B(in[1509]), .Z(n4515) );
  XOR U5486 ( .A(in[1120]), .B(n3702), .Z(n4512) );
  NAND U5487 ( .A(n4515), .B(n4512), .Z(n3703) );
  XNOR U5488 ( .A(n4099), .B(n3703), .Z(out[678]) );
  XOR U5489 ( .A(in[277]), .B(n3704), .Z(n4102) );
  XOR U5490 ( .A(in[1510]), .B(n3705), .Z(n4519) );
  XOR U5491 ( .A(in[1121]), .B(n3706), .Z(n4516) );
  NAND U5492 ( .A(n4519), .B(n4516), .Z(n3707) );
  XNOR U5493 ( .A(n4102), .B(n3707), .Z(out[679]) );
  ANDN U5494 ( .B(n3709), .A(n3708), .Z(n3710) );
  XNOR U5495 ( .A(n3711), .B(n3710), .Z(out[67]) );
  XOR U5496 ( .A(in[278]), .B(n3712), .Z(n4105) );
  XOR U5497 ( .A(in[1511]), .B(n3713), .Z(n4523) );
  XOR U5498 ( .A(in[1122]), .B(n3714), .Z(n4520) );
  NAND U5499 ( .A(n4523), .B(n4520), .Z(n3715) );
  XNOR U5500 ( .A(n4105), .B(n3715), .Z(out[680]) );
  XOR U5501 ( .A(in[279]), .B(n3716), .Z(n4108) );
  XOR U5502 ( .A(in[1512]), .B(n3717), .Z(n4527) );
  XOR U5503 ( .A(in[1123]), .B(n3718), .Z(n4524) );
  NAND U5504 ( .A(n4527), .B(n4524), .Z(n3719) );
  XNOR U5505 ( .A(n4108), .B(n3719), .Z(out[681]) );
  XOR U5506 ( .A(in[280]), .B(n3720), .Z(n4115) );
  XOR U5507 ( .A(in[1513]), .B(n3721), .Z(n4531) );
  XOR U5508 ( .A(in[1124]), .B(n3722), .Z(n4528) );
  NAND U5509 ( .A(n4531), .B(n4528), .Z(n3723) );
  XNOR U5510 ( .A(n4115), .B(n3723), .Z(out[682]) );
  XOR U5511 ( .A(in[281]), .B(n3724), .Z(n4118) );
  XOR U5512 ( .A(in[1514]), .B(n3725), .Z(n4535) );
  XOR U5513 ( .A(in[1125]), .B(n3726), .Z(n4532) );
  NAND U5514 ( .A(n4535), .B(n4532), .Z(n3727) );
  XNOR U5515 ( .A(n4118), .B(n3727), .Z(out[683]) );
  XOR U5516 ( .A(in[282]), .B(n3728), .Z(n4121) );
  XOR U5517 ( .A(in[1515]), .B(n3729), .Z(n4543) );
  XNOR U5518 ( .A(in[1126]), .B(n3730), .Z(n4540) );
  NAND U5519 ( .A(n4543), .B(n4540), .Z(n3731) );
  XNOR U5520 ( .A(n4121), .B(n3731), .Z(out[684]) );
  XOR U5521 ( .A(in[283]), .B(n3732), .Z(n4124) );
  XOR U5522 ( .A(in[1516]), .B(n3733), .Z(n4547) );
  XNOR U5523 ( .A(in[1127]), .B(n3734), .Z(n4544) );
  NAND U5524 ( .A(n4547), .B(n4544), .Z(n3735) );
  XNOR U5525 ( .A(n4124), .B(n3735), .Z(out[685]) );
  XOR U5526 ( .A(in[284]), .B(n3736), .Z(n4127) );
  XOR U5527 ( .A(in[1517]), .B(n3737), .Z(n4551) );
  XNOR U5528 ( .A(in[1128]), .B(n3738), .Z(n4548) );
  NAND U5529 ( .A(n4551), .B(n4548), .Z(n3739) );
  XNOR U5530 ( .A(n4127), .B(n3739), .Z(out[686]) );
  XOR U5531 ( .A(in[285]), .B(n3740), .Z(n4130) );
  XOR U5532 ( .A(in[1518]), .B(n3741), .Z(n4555) );
  XNOR U5533 ( .A(in[1129]), .B(n3742), .Z(n4552) );
  NAND U5534 ( .A(n4555), .B(n4552), .Z(n3743) );
  XNOR U5535 ( .A(n4130), .B(n3743), .Z(out[687]) );
  XOR U5536 ( .A(in[286]), .B(n3744), .Z(n4133) );
  XOR U5537 ( .A(in[1519]), .B(n3745), .Z(n4559) );
  XNOR U5538 ( .A(in[1130]), .B(n3746), .Z(n4556) );
  NAND U5539 ( .A(n4559), .B(n4556), .Z(n3747) );
  XNOR U5540 ( .A(n4133), .B(n3747), .Z(out[688]) );
  XOR U5541 ( .A(in[287]), .B(n3748), .Z(n4136) );
  XOR U5542 ( .A(in[1520]), .B(n3749), .Z(n4563) );
  XNOR U5543 ( .A(in[1131]), .B(n3750), .Z(n4560) );
  NAND U5544 ( .A(n4563), .B(n4560), .Z(n3751) );
  XNOR U5545 ( .A(n4136), .B(n3751), .Z(out[689]) );
  ANDN U5546 ( .B(n3753), .A(n3752), .Z(n3754) );
  XNOR U5547 ( .A(n3755), .B(n3754), .Z(out[68]) );
  XOR U5548 ( .A(in[288]), .B(n3756), .Z(n4139) );
  XOR U5549 ( .A(in[1521]), .B(n3757), .Z(n4567) );
  XNOR U5550 ( .A(in[1132]), .B(n3758), .Z(n4564) );
  NAND U5551 ( .A(n4567), .B(n4564), .Z(n3759) );
  XNOR U5552 ( .A(n4139), .B(n3759), .Z(out[690]) );
  XOR U5553 ( .A(in[289]), .B(n3760), .Z(n4142) );
  XOR U5554 ( .A(in[1522]), .B(n3761), .Z(n4571) );
  XNOR U5555 ( .A(in[1133]), .B(n3762), .Z(n4568) );
  NAND U5556 ( .A(n4571), .B(n4568), .Z(n3763) );
  XNOR U5557 ( .A(n4142), .B(n3763), .Z(out[691]) );
  XOR U5558 ( .A(in[290]), .B(n3764), .Z(n4149) );
  XOR U5559 ( .A(in[1523]), .B(n3765), .Z(n4575) );
  XNOR U5560 ( .A(in[1134]), .B(n3766), .Z(n4572) );
  NAND U5561 ( .A(n4575), .B(n4572), .Z(n3767) );
  XNOR U5562 ( .A(n4149), .B(n3767), .Z(out[692]) );
  XOR U5563 ( .A(in[291]), .B(n3768), .Z(n4152) );
  XOR U5564 ( .A(in[1524]), .B(n3769), .Z(n4579) );
  XNOR U5565 ( .A(in[1135]), .B(n3770), .Z(n4576) );
  NAND U5566 ( .A(n4579), .B(n4576), .Z(n3771) );
  XNOR U5567 ( .A(n4152), .B(n3771), .Z(out[693]) );
  XOR U5568 ( .A(in[292]), .B(n3772), .Z(n4155) );
  XOR U5569 ( .A(in[1525]), .B(n3773), .Z(n4587) );
  XNOR U5570 ( .A(in[1136]), .B(n3774), .Z(n4584) );
  NAND U5571 ( .A(n4587), .B(n4584), .Z(n3775) );
  XNOR U5572 ( .A(n4155), .B(n3775), .Z(out[694]) );
  XNOR U5573 ( .A(in[293]), .B(n3776), .Z(n4158) );
  XOR U5574 ( .A(in[1526]), .B(n3777), .Z(n4591) );
  XNOR U5575 ( .A(in[1137]), .B(n3778), .Z(n4588) );
  NAND U5576 ( .A(n4591), .B(n4588), .Z(n3779) );
  XNOR U5577 ( .A(n4158), .B(n3779), .Z(out[695]) );
  XNOR U5578 ( .A(in[294]), .B(n3780), .Z(n4161) );
  XOR U5579 ( .A(in[1527]), .B(n3781), .Z(n4595) );
  XNOR U5580 ( .A(in[1138]), .B(n3782), .Z(n4592) );
  NAND U5581 ( .A(n4595), .B(n4592), .Z(n3783) );
  XNOR U5582 ( .A(n4161), .B(n3783), .Z(out[696]) );
  XNOR U5583 ( .A(in[295]), .B(n3784), .Z(n4164) );
  XOR U5584 ( .A(in[1528]), .B(n3785), .Z(n4599) );
  XNOR U5585 ( .A(in[1139]), .B(n3786), .Z(n4596) );
  NAND U5586 ( .A(n4599), .B(n4596), .Z(n3787) );
  XNOR U5587 ( .A(n4164), .B(n3787), .Z(out[697]) );
  XNOR U5588 ( .A(in[296]), .B(n3788), .Z(n4167) );
  XOR U5589 ( .A(in[1529]), .B(n3789), .Z(n4603) );
  XNOR U5590 ( .A(in[1140]), .B(n3790), .Z(n4600) );
  NAND U5591 ( .A(n4603), .B(n4600), .Z(n3791) );
  XNOR U5592 ( .A(n4167), .B(n3791), .Z(out[698]) );
  XNOR U5593 ( .A(in[297]), .B(n3792), .Z(n4170) );
  XOR U5594 ( .A(in[1530]), .B(n3793), .Z(n4607) );
  XNOR U5595 ( .A(in[1141]), .B(n3794), .Z(n4604) );
  NAND U5596 ( .A(n4607), .B(n4604), .Z(n3795) );
  XNOR U5597 ( .A(n4170), .B(n3795), .Z(out[699]) );
  ANDN U5598 ( .B(n3797), .A(n3796), .Z(n3798) );
  XNOR U5599 ( .A(n3799), .B(n3798), .Z(out[69]) );
  OR U5600 ( .A(n3831), .B(n3800), .Z(n3801) );
  XNOR U5601 ( .A(n3830), .B(n3801), .Z(out[6]) );
  XNOR U5602 ( .A(in[298]), .B(n3802), .Z(n4173) );
  XNOR U5603 ( .A(in[1531]), .B(n3803), .Z(n4611) );
  XNOR U5604 ( .A(in[1142]), .B(n3804), .Z(n4608) );
  NAND U5605 ( .A(n4611), .B(n4608), .Z(n3805) );
  XNOR U5606 ( .A(n4173), .B(n3805), .Z(out[700]) );
  XNOR U5607 ( .A(in[299]), .B(n3806), .Z(n4176) );
  XNOR U5608 ( .A(in[1532]), .B(n3807), .Z(n4615) );
  XNOR U5609 ( .A(in[1143]), .B(n3808), .Z(n4612) );
  NAND U5610 ( .A(n4615), .B(n4612), .Z(n3809) );
  XNOR U5611 ( .A(n4176), .B(n3809), .Z(out[701]) );
  XNOR U5612 ( .A(in[300]), .B(n3810), .Z(n4183) );
  XNOR U5613 ( .A(in[1533]), .B(n3811), .Z(n4619) );
  XNOR U5614 ( .A(in[1144]), .B(n3812), .Z(n4616) );
  NAND U5615 ( .A(n4619), .B(n4616), .Z(n3813) );
  XNOR U5616 ( .A(n4183), .B(n3813), .Z(out[702]) );
  XNOR U5617 ( .A(in[301]), .B(n3814), .Z(n4186) );
  XOR U5618 ( .A(in[1534]), .B(n3815), .Z(n4623) );
  XNOR U5619 ( .A(in[1145]), .B(n3816), .Z(n4620) );
  NAND U5620 ( .A(n4623), .B(n4620), .Z(n3817) );
  XNOR U5621 ( .A(n4186), .B(n3817), .Z(out[703]) );
  XOR U5622 ( .A(in[376]), .B(n3818), .Z(n4188) );
  NOR U5623 ( .A(n3965), .B(n4343), .Z(n3819) );
  XNOR U5624 ( .A(n4188), .B(n3819), .Z(out[704]) );
  XOR U5625 ( .A(in[377]), .B(n3820), .Z(n4190) );
  NOR U5626 ( .A(n3968), .B(n4347), .Z(n3821) );
  XNOR U5627 ( .A(n4190), .B(n3821), .Z(out[705]) );
  XOR U5628 ( .A(in[378]), .B(n3822), .Z(n4192) );
  NOR U5629 ( .A(n3975), .B(n4351), .Z(n3823) );
  XNOR U5630 ( .A(n4192), .B(n3823), .Z(out[706]) );
  XOR U5631 ( .A(in[379]), .B(n3824), .Z(n4194) );
  NOR U5632 ( .A(n3978), .B(n4355), .Z(n3825) );
  XNOR U5633 ( .A(n4194), .B(n3825), .Z(out[707]) );
  XOR U5634 ( .A(in[380]), .B(n3826), .Z(n4196) );
  NOR U5635 ( .A(n3981), .B(n4367), .Z(n3827) );
  XNOR U5636 ( .A(n4196), .B(n3827), .Z(out[708]) );
  XOR U5637 ( .A(in[381]), .B(n3828), .Z(n4198) );
  NOR U5638 ( .A(n3984), .B(n4371), .Z(n3829) );
  XNOR U5639 ( .A(n4198), .B(n3829), .Z(out[709]) );
  ANDN U5640 ( .B(n3831), .A(n3830), .Z(n3832) );
  XNOR U5641 ( .A(n3833), .B(n3832), .Z(out[70]) );
  XOR U5642 ( .A(in[382]), .B(n3834), .Z(n4200) );
  NOR U5643 ( .A(n3987), .B(n4375), .Z(n3835) );
  XNOR U5644 ( .A(n4200), .B(n3835), .Z(out[710]) );
  XOR U5645 ( .A(in[383]), .B(n3836), .Z(n4202) );
  NOR U5646 ( .A(n3990), .B(n4379), .Z(n3837) );
  XNOR U5647 ( .A(n4202), .B(n3837), .Z(out[711]) );
  XOR U5648 ( .A(in[320]), .B(n3838), .Z(n4208) );
  NOR U5649 ( .A(n3993), .B(n4383), .Z(n3839) );
  XNOR U5650 ( .A(n4208), .B(n3839), .Z(out[712]) );
  XOR U5651 ( .A(in[321]), .B(n3840), .Z(n4210) );
  NOR U5652 ( .A(n3996), .B(n4387), .Z(n3841) );
  XNOR U5653 ( .A(n4210), .B(n3841), .Z(out[713]) );
  XOR U5654 ( .A(in[322]), .B(n3842), .Z(n4212) );
  NOR U5655 ( .A(n3999), .B(n4391), .Z(n3843) );
  XNOR U5656 ( .A(n4212), .B(n3843), .Z(out[714]) );
  XOR U5657 ( .A(in[323]), .B(n3844), .Z(n4214) );
  NOR U5658 ( .A(n4002), .B(n4395), .Z(n3845) );
  XNOR U5659 ( .A(n4214), .B(n3845), .Z(out[715]) );
  XOR U5660 ( .A(in[324]), .B(n3846), .Z(n4216) );
  NOR U5661 ( .A(n4009), .B(n4399), .Z(n3847) );
  XNOR U5662 ( .A(n4216), .B(n3847), .Z(out[716]) );
  XOR U5663 ( .A(in[325]), .B(n3848), .Z(n4218) );
  NOR U5664 ( .A(n4012), .B(n4403), .Z(n3849) );
  XNOR U5665 ( .A(n4218), .B(n3849), .Z(out[717]) );
  XOR U5666 ( .A(in[326]), .B(n3850), .Z(n4220) );
  NOR U5667 ( .A(n4015), .B(n4411), .Z(n3851) );
  XNOR U5668 ( .A(n4220), .B(n3851), .Z(out[718]) );
  XOR U5669 ( .A(in[327]), .B(n3852), .Z(n4222) );
  NOR U5670 ( .A(n4018), .B(n4415), .Z(n3853) );
  XNOR U5671 ( .A(n4222), .B(n3853), .Z(out[719]) );
  ANDN U5672 ( .B(n4077), .A(n4079), .Z(n3854) );
  XNOR U5673 ( .A(n3855), .B(n3854), .Z(out[71]) );
  XOR U5674 ( .A(in[328]), .B(n3856), .Z(n4224) );
  NOR U5675 ( .A(n4021), .B(n4419), .Z(n3857) );
  XNOR U5676 ( .A(n4224), .B(n3857), .Z(out[720]) );
  XOR U5677 ( .A(in[329]), .B(n3858), .Z(n4226) );
  NOR U5678 ( .A(n4024), .B(n4423), .Z(n3859) );
  XNOR U5679 ( .A(n4226), .B(n3859), .Z(out[721]) );
  XOR U5680 ( .A(in[330]), .B(n3860), .Z(n4232) );
  NOR U5681 ( .A(n4027), .B(n4427), .Z(n3861) );
  XNOR U5682 ( .A(n4232), .B(n3861), .Z(out[722]) );
  XOR U5683 ( .A(in[331]), .B(n3862), .Z(n4234) );
  NOR U5684 ( .A(n4030), .B(n4431), .Z(n3863) );
  XNOR U5685 ( .A(n4234), .B(n3863), .Z(out[723]) );
  XOR U5686 ( .A(in[332]), .B(n3864), .Z(n4236) );
  NOR U5687 ( .A(n4033), .B(n4435), .Z(n3865) );
  XNOR U5688 ( .A(n4236), .B(n3865), .Z(out[724]) );
  XOR U5689 ( .A(in[333]), .B(n3866), .Z(n4238) );
  NOR U5690 ( .A(n4036), .B(n4439), .Z(n3867) );
  XNOR U5691 ( .A(n4238), .B(n3867), .Z(out[725]) );
  XOR U5692 ( .A(in[334]), .B(n3868), .Z(n4240) );
  NOR U5693 ( .A(n4043), .B(n4443), .Z(n3869) );
  XNOR U5694 ( .A(n4240), .B(n3869), .Z(out[726]) );
  XOR U5695 ( .A(in[335]), .B(n3870), .Z(n4242) );
  NOR U5696 ( .A(n4046), .B(n4447), .Z(n3871) );
  XNOR U5697 ( .A(n4242), .B(n3871), .Z(out[727]) );
  XOR U5698 ( .A(in[336]), .B(n3872), .Z(n4244) );
  NOR U5699 ( .A(n4049), .B(n4455), .Z(n3873) );
  XNOR U5700 ( .A(n4244), .B(n3873), .Z(out[728]) );
  XOR U5701 ( .A(in[337]), .B(n3874), .Z(n4246) );
  NOR U5702 ( .A(n4052), .B(n4459), .Z(n3875) );
  XNOR U5703 ( .A(n4246), .B(n3875), .Z(out[729]) );
  ANDN U5704 ( .B(n4361), .A(n4363), .Z(n3876) );
  XNOR U5705 ( .A(n3877), .B(n3876), .Z(out[72]) );
  XOR U5706 ( .A(in[338]), .B(n3878), .Z(n4248) );
  NOR U5707 ( .A(n4055), .B(n4463), .Z(n3879) );
  XNOR U5708 ( .A(n4248), .B(n3879), .Z(out[730]) );
  XOR U5709 ( .A(in[339]), .B(n3880), .Z(n4250) );
  NOR U5710 ( .A(n4058), .B(n4467), .Z(n3881) );
  XNOR U5711 ( .A(n4250), .B(n3881), .Z(out[731]) );
  XOR U5712 ( .A(in[340]), .B(n3882), .Z(n4256) );
  NOR U5713 ( .A(n4061), .B(n4471), .Z(n3883) );
  XNOR U5714 ( .A(n4256), .B(n3883), .Z(out[732]) );
  XOR U5715 ( .A(in[341]), .B(n3884), .Z(n4258) );
  NOR U5716 ( .A(n4064), .B(n4475), .Z(n3885) );
  XNOR U5717 ( .A(n4258), .B(n3885), .Z(out[733]) );
  XOR U5718 ( .A(in[342]), .B(n3886), .Z(n4260) );
  NOR U5719 ( .A(n4067), .B(n4479), .Z(n3887) );
  XNOR U5720 ( .A(n4260), .B(n3887), .Z(out[734]) );
  XOR U5721 ( .A(in[343]), .B(n3888), .Z(n4262) );
  NOR U5722 ( .A(n4070), .B(n4483), .Z(n3889) );
  XNOR U5723 ( .A(n4262), .B(n3889), .Z(out[735]) );
  XOR U5724 ( .A(in[344]), .B(n3890), .Z(n4264) );
  NOR U5725 ( .A(n4081), .B(n4487), .Z(n3891) );
  XNOR U5726 ( .A(n4264), .B(n3891), .Z(out[736]) );
  XOR U5727 ( .A(in[345]), .B(n3892), .Z(n4266) );
  NOR U5728 ( .A(n4084), .B(n4491), .Z(n3893) );
  XNOR U5729 ( .A(n4266), .B(n3893), .Z(out[737]) );
  XOR U5730 ( .A(in[346]), .B(n3894), .Z(n4268) );
  NOR U5731 ( .A(n4087), .B(n4499), .Z(n3895) );
  XNOR U5732 ( .A(n4268), .B(n3895), .Z(out[738]) );
  XOR U5733 ( .A(in[347]), .B(n3896), .Z(n4270) );
  NOR U5734 ( .A(n4090), .B(n4503), .Z(n3897) );
  XNOR U5735 ( .A(n4270), .B(n3897), .Z(out[739]) );
  ANDN U5736 ( .B(n4805), .A(n4807), .Z(n3898) );
  XNOR U5737 ( .A(n3899), .B(n3898), .Z(out[73]) );
  XOR U5738 ( .A(in[348]), .B(n3900), .Z(n4272) );
  NOR U5739 ( .A(n4093), .B(n4507), .Z(n3901) );
  XNOR U5740 ( .A(n4272), .B(n3901), .Z(out[740]) );
  XOR U5741 ( .A(in[349]), .B(n3902), .Z(n4274) );
  NOR U5742 ( .A(n4096), .B(n4511), .Z(n3903) );
  XNOR U5743 ( .A(n4274), .B(n3903), .Z(out[741]) );
  XOR U5744 ( .A(in[350]), .B(n3904), .Z(n4280) );
  NOR U5745 ( .A(n4099), .B(n4515), .Z(n3905) );
  XNOR U5746 ( .A(n4280), .B(n3905), .Z(out[742]) );
  XOR U5747 ( .A(in[351]), .B(n3906), .Z(n4282) );
  NOR U5748 ( .A(n4102), .B(n4519), .Z(n3907) );
  XNOR U5749 ( .A(n4282), .B(n3907), .Z(out[743]) );
  XOR U5750 ( .A(in[352]), .B(n3908), .Z(n4284) );
  NOR U5751 ( .A(n4105), .B(n4523), .Z(n3909) );
  XNOR U5752 ( .A(n4284), .B(n3909), .Z(out[744]) );
  XOR U5753 ( .A(in[353]), .B(n3910), .Z(n4286) );
  NOR U5754 ( .A(n4108), .B(n4527), .Z(n3911) );
  XNOR U5755 ( .A(n4286), .B(n3911), .Z(out[745]) );
  XOR U5756 ( .A(in[354]), .B(n3912), .Z(n4288) );
  NOR U5757 ( .A(n4115), .B(n4531), .Z(n3913) );
  XNOR U5758 ( .A(n4288), .B(n3913), .Z(out[746]) );
  XOR U5759 ( .A(in[355]), .B(n3914), .Z(n4290) );
  NOR U5760 ( .A(n4118), .B(n4535), .Z(n3915) );
  XNOR U5761 ( .A(n4290), .B(n3915), .Z(out[747]) );
  XOR U5762 ( .A(in[356]), .B(n3916), .Z(n4292) );
  NOR U5763 ( .A(n4121), .B(n4543), .Z(n3917) );
  XNOR U5764 ( .A(n4292), .B(n3917), .Z(out[748]) );
  XOR U5765 ( .A(in[357]), .B(n3918), .Z(n4294) );
  NOR U5766 ( .A(n4124), .B(n4547), .Z(n3919) );
  XNOR U5767 ( .A(n4294), .B(n3919), .Z(out[749]) );
  NOR U5768 ( .A(n3921), .B(n3920), .Z(n3922) );
  XNOR U5769 ( .A(n3923), .B(n3922), .Z(out[74]) );
  XOR U5770 ( .A(in[358]), .B(n3924), .Z(n4296) );
  NOR U5771 ( .A(n4127), .B(n4551), .Z(n3925) );
  XNOR U5772 ( .A(n4296), .B(n3925), .Z(out[750]) );
  XOR U5773 ( .A(in[359]), .B(n3926), .Z(n4298) );
  NOR U5774 ( .A(n4130), .B(n4555), .Z(n3927) );
  XNOR U5775 ( .A(n4298), .B(n3927), .Z(out[751]) );
  XOR U5776 ( .A(in[360]), .B(n3928), .Z(n4304) );
  NOR U5777 ( .A(n4133), .B(n4559), .Z(n3929) );
  XNOR U5778 ( .A(n4304), .B(n3929), .Z(out[752]) );
  XOR U5779 ( .A(in[361]), .B(n3930), .Z(n4306) );
  NOR U5780 ( .A(n4136), .B(n4563), .Z(n3931) );
  XNOR U5781 ( .A(n4306), .B(n3931), .Z(out[753]) );
  XOR U5782 ( .A(in[362]), .B(n3932), .Z(n4308) );
  NOR U5783 ( .A(n4139), .B(n4567), .Z(n3933) );
  XNOR U5784 ( .A(n4308), .B(n3933), .Z(out[754]) );
  XOR U5785 ( .A(in[363]), .B(n3934), .Z(n4310) );
  NOR U5786 ( .A(n4142), .B(n4571), .Z(n3935) );
  XNOR U5787 ( .A(n4310), .B(n3935), .Z(out[755]) );
  XOR U5788 ( .A(in[364]), .B(n3936), .Z(n4312) );
  NOR U5789 ( .A(n4149), .B(n4575), .Z(n3937) );
  XNOR U5790 ( .A(n4312), .B(n3937), .Z(out[756]) );
  XOR U5791 ( .A(in[365]), .B(n3938), .Z(n4314) );
  NOR U5792 ( .A(n4152), .B(n4579), .Z(n3939) );
  XNOR U5793 ( .A(n4314), .B(n3939), .Z(out[757]) );
  XOR U5794 ( .A(in[366]), .B(n3940), .Z(n4316) );
  NOR U5795 ( .A(n4155), .B(n4587), .Z(n3941) );
  XNOR U5796 ( .A(n4316), .B(n3941), .Z(out[758]) );
  XOR U5797 ( .A(in[367]), .B(n3942), .Z(n4318) );
  NOR U5798 ( .A(n4158), .B(n4591), .Z(n3943) );
  XNOR U5799 ( .A(n4318), .B(n3943), .Z(out[759]) );
  NOR U5800 ( .A(n3945), .B(n3944), .Z(n3946) );
  XNOR U5801 ( .A(n3947), .B(n3946), .Z(out[75]) );
  XOR U5802 ( .A(in[368]), .B(n3948), .Z(n4320) );
  NOR U5803 ( .A(n4161), .B(n4595), .Z(n3949) );
  XNOR U5804 ( .A(n4320), .B(n3949), .Z(out[760]) );
  XOR U5805 ( .A(in[369]), .B(n3950), .Z(n4322) );
  NOR U5806 ( .A(n4164), .B(n4599), .Z(n3951) );
  XNOR U5807 ( .A(n4322), .B(n3951), .Z(out[761]) );
  XOR U5808 ( .A(in[370]), .B(n3952), .Z(n4328) );
  NOR U5809 ( .A(n4167), .B(n4603), .Z(n3953) );
  XNOR U5810 ( .A(n4328), .B(n3953), .Z(out[762]) );
  XOR U5811 ( .A(in[371]), .B(n3954), .Z(n4330) );
  NOR U5812 ( .A(n4170), .B(n4607), .Z(n3955) );
  XNOR U5813 ( .A(n4330), .B(n3955), .Z(out[763]) );
  XOR U5814 ( .A(in[372]), .B(n3956), .Z(n4332) );
  NOR U5815 ( .A(n4173), .B(n4611), .Z(n3957) );
  XNOR U5816 ( .A(n4332), .B(n3957), .Z(out[764]) );
  XOR U5817 ( .A(in[373]), .B(n3958), .Z(n4334) );
  NOR U5818 ( .A(n4176), .B(n4615), .Z(n3959) );
  XNOR U5819 ( .A(n4334), .B(n3959), .Z(out[765]) );
  XOR U5820 ( .A(in[374]), .B(n3960), .Z(n4336) );
  NOR U5821 ( .A(n4183), .B(n4619), .Z(n3961) );
  XNOR U5822 ( .A(n4336), .B(n3961), .Z(out[766]) );
  XOR U5823 ( .A(in[375]), .B(n3962), .Z(n4338) );
  NOR U5824 ( .A(n4186), .B(n4623), .Z(n3963) );
  XNOR U5825 ( .A(n4338), .B(n3963), .Z(out[767]) );
  XNOR U5826 ( .A(in[743]), .B(n3964), .Z(n4341) );
  NAND U5827 ( .A(n4188), .B(n3965), .Z(n3966) );
  XNOR U5828 ( .A(n4341), .B(n3966), .Z(out[768]) );
  XNOR U5829 ( .A(in[744]), .B(n3967), .Z(n4345) );
  NAND U5830 ( .A(n4190), .B(n3968), .Z(n3969) );
  XNOR U5831 ( .A(n4345), .B(n3969), .Z(out[769]) );
  NOR U5832 ( .A(n3971), .B(n3970), .Z(n3972) );
  XNOR U5833 ( .A(n3973), .B(n3972), .Z(out[76]) );
  XNOR U5834 ( .A(in[745]), .B(n3974), .Z(n4349) );
  NAND U5835 ( .A(n4192), .B(n3975), .Z(n3976) );
  XNOR U5836 ( .A(n4349), .B(n3976), .Z(out[770]) );
  XNOR U5837 ( .A(in[746]), .B(n3977), .Z(n4353) );
  NAND U5838 ( .A(n4194), .B(n3978), .Z(n3979) );
  XNOR U5839 ( .A(n4353), .B(n3979), .Z(out[771]) );
  XNOR U5840 ( .A(in[747]), .B(n3980), .Z(n4365) );
  NAND U5841 ( .A(n4196), .B(n3981), .Z(n3982) );
  XNOR U5842 ( .A(n4365), .B(n3982), .Z(out[772]) );
  XNOR U5843 ( .A(in[748]), .B(n3983), .Z(n4369) );
  NAND U5844 ( .A(n4198), .B(n3984), .Z(n3985) );
  XNOR U5845 ( .A(n4369), .B(n3985), .Z(out[773]) );
  XNOR U5846 ( .A(in[749]), .B(n3986), .Z(n4373) );
  NAND U5847 ( .A(n4200), .B(n3987), .Z(n3988) );
  XNOR U5848 ( .A(n4373), .B(n3988), .Z(out[774]) );
  XNOR U5849 ( .A(in[750]), .B(n3989), .Z(n4377) );
  NAND U5850 ( .A(n4202), .B(n3990), .Z(n3991) );
  XNOR U5851 ( .A(n4377), .B(n3991), .Z(out[775]) );
  XNOR U5852 ( .A(in[751]), .B(n3992), .Z(n4381) );
  NAND U5853 ( .A(n4208), .B(n3993), .Z(n3994) );
  XNOR U5854 ( .A(n4381), .B(n3994), .Z(out[776]) );
  XNOR U5855 ( .A(in[752]), .B(n3995), .Z(n4385) );
  NAND U5856 ( .A(n4210), .B(n3996), .Z(n3997) );
  XNOR U5857 ( .A(n4385), .B(n3997), .Z(out[777]) );
  XNOR U5858 ( .A(in[753]), .B(n3998), .Z(n4389) );
  NAND U5859 ( .A(n4212), .B(n3999), .Z(n4000) );
  XNOR U5860 ( .A(n4389), .B(n4000), .Z(out[778]) );
  XNOR U5861 ( .A(in[754]), .B(n4001), .Z(n4393) );
  NAND U5862 ( .A(n4214), .B(n4002), .Z(n4003) );
  XNOR U5863 ( .A(n4393), .B(n4003), .Z(out[779]) );
  NOR U5864 ( .A(n4005), .B(n4004), .Z(n4006) );
  XNOR U5865 ( .A(n4007), .B(n4006), .Z(out[77]) );
  XNOR U5866 ( .A(in[755]), .B(n4008), .Z(n4397) );
  NAND U5867 ( .A(n4216), .B(n4009), .Z(n4010) );
  XNOR U5868 ( .A(n4397), .B(n4010), .Z(out[780]) );
  XNOR U5869 ( .A(in[756]), .B(n4011), .Z(n4401) );
  NAND U5870 ( .A(n4218), .B(n4012), .Z(n4013) );
  XNOR U5871 ( .A(n4401), .B(n4013), .Z(out[781]) );
  XNOR U5872 ( .A(in[757]), .B(n4014), .Z(n4409) );
  NAND U5873 ( .A(n4220), .B(n4015), .Z(n4016) );
  XNOR U5874 ( .A(n4409), .B(n4016), .Z(out[782]) );
  XNOR U5875 ( .A(in[758]), .B(n4017), .Z(n4413) );
  NAND U5876 ( .A(n4222), .B(n4018), .Z(n4019) );
  XNOR U5877 ( .A(n4413), .B(n4019), .Z(out[783]) );
  XNOR U5878 ( .A(in[759]), .B(n4020), .Z(n4417) );
  NAND U5879 ( .A(n4224), .B(n4021), .Z(n4022) );
  XNOR U5880 ( .A(n4417), .B(n4022), .Z(out[784]) );
  XNOR U5881 ( .A(in[760]), .B(n4023), .Z(n4421) );
  NAND U5882 ( .A(n4226), .B(n4024), .Z(n4025) );
  XNOR U5883 ( .A(n4421), .B(n4025), .Z(out[785]) );
  XNOR U5884 ( .A(in[761]), .B(n4026), .Z(n4425) );
  NAND U5885 ( .A(n4232), .B(n4027), .Z(n4028) );
  XNOR U5886 ( .A(n4425), .B(n4028), .Z(out[786]) );
  XNOR U5887 ( .A(in[762]), .B(n4029), .Z(n4429) );
  NAND U5888 ( .A(n4234), .B(n4030), .Z(n4031) );
  XNOR U5889 ( .A(n4429), .B(n4031), .Z(out[787]) );
  XNOR U5890 ( .A(in[763]), .B(n4032), .Z(n4433) );
  NAND U5891 ( .A(n4236), .B(n4033), .Z(n4034) );
  XNOR U5892 ( .A(n4433), .B(n4034), .Z(out[788]) );
  XNOR U5893 ( .A(in[764]), .B(n4035), .Z(n4437) );
  NAND U5894 ( .A(n4238), .B(n4036), .Z(n4037) );
  XNOR U5895 ( .A(n4437), .B(n4037), .Z(out[789]) );
  NOR U5896 ( .A(n4039), .B(n4038), .Z(n4040) );
  XNOR U5897 ( .A(n4041), .B(n4040), .Z(out[78]) );
  XNOR U5898 ( .A(in[765]), .B(n4042), .Z(n4441) );
  NAND U5899 ( .A(n4240), .B(n4043), .Z(n4044) );
  XNOR U5900 ( .A(n4441), .B(n4044), .Z(out[790]) );
  XNOR U5901 ( .A(in[766]), .B(n4045), .Z(n4445) );
  NAND U5902 ( .A(n4242), .B(n4046), .Z(n4047) );
  XNOR U5903 ( .A(n4445), .B(n4047), .Z(out[791]) );
  XNOR U5904 ( .A(in[767]), .B(n4048), .Z(n4453) );
  NAND U5905 ( .A(n4244), .B(n4049), .Z(n4050) );
  XNOR U5906 ( .A(n4453), .B(n4050), .Z(out[792]) );
  XNOR U5907 ( .A(in[704]), .B(n4051), .Z(n4457) );
  NAND U5908 ( .A(n4246), .B(n4052), .Z(n4053) );
  XNOR U5909 ( .A(n4457), .B(n4053), .Z(out[793]) );
  XNOR U5910 ( .A(in[705]), .B(n4054), .Z(n4461) );
  NAND U5911 ( .A(n4248), .B(n4055), .Z(n4056) );
  XNOR U5912 ( .A(n4461), .B(n4056), .Z(out[794]) );
  XNOR U5913 ( .A(in[706]), .B(n4057), .Z(n4465) );
  NAND U5914 ( .A(n4250), .B(n4058), .Z(n4059) );
  XNOR U5915 ( .A(n4465), .B(n4059), .Z(out[795]) );
  XNOR U5916 ( .A(in[707]), .B(n4060), .Z(n4469) );
  NAND U5917 ( .A(n4256), .B(n4061), .Z(n4062) );
  XNOR U5918 ( .A(n4469), .B(n4062), .Z(out[796]) );
  XNOR U5919 ( .A(in[708]), .B(n4063), .Z(n4473) );
  NAND U5920 ( .A(n4258), .B(n4064), .Z(n4065) );
  XNOR U5921 ( .A(n4473), .B(n4065), .Z(out[797]) );
  XNOR U5922 ( .A(in[709]), .B(n4066), .Z(n4477) );
  NAND U5923 ( .A(n4260), .B(n4067), .Z(n4068) );
  XNOR U5924 ( .A(n4477), .B(n4068), .Z(out[798]) );
  XNOR U5925 ( .A(in[710]), .B(n4069), .Z(n4481) );
  NAND U5926 ( .A(n4262), .B(n4070), .Z(n4071) );
  XNOR U5927 ( .A(n4481), .B(n4071), .Z(out[799]) );
  NOR U5928 ( .A(n4073), .B(n4072), .Z(n4074) );
  XNOR U5929 ( .A(n4075), .B(n4074), .Z(out[79]) );
  OR U5930 ( .A(n4077), .B(n4076), .Z(n4078) );
  XNOR U5931 ( .A(n4079), .B(n4078), .Z(out[7]) );
  XNOR U5932 ( .A(in[711]), .B(n4080), .Z(n4485) );
  NAND U5933 ( .A(n4264), .B(n4081), .Z(n4082) );
  XNOR U5934 ( .A(n4485), .B(n4082), .Z(out[800]) );
  XNOR U5935 ( .A(in[712]), .B(n4083), .Z(n4489) );
  NAND U5936 ( .A(n4266), .B(n4084), .Z(n4085) );
  XNOR U5937 ( .A(n4489), .B(n4085), .Z(out[801]) );
  XNOR U5938 ( .A(in[713]), .B(n4086), .Z(n4497) );
  NAND U5939 ( .A(n4268), .B(n4087), .Z(n4088) );
  XNOR U5940 ( .A(n4497), .B(n4088), .Z(out[802]) );
  XNOR U5941 ( .A(in[714]), .B(n4089), .Z(n4501) );
  NAND U5942 ( .A(n4270), .B(n4090), .Z(n4091) );
  XNOR U5943 ( .A(n4501), .B(n4091), .Z(out[803]) );
  XNOR U5944 ( .A(in[715]), .B(n4092), .Z(n4505) );
  NAND U5945 ( .A(n4272), .B(n4093), .Z(n4094) );
  XNOR U5946 ( .A(n4505), .B(n4094), .Z(out[804]) );
  XOR U5947 ( .A(n4095), .B(in[716]), .Z(n4509) );
  NAND U5948 ( .A(n4274), .B(n4096), .Z(n4097) );
  XNOR U5949 ( .A(n4509), .B(n4097), .Z(out[805]) );
  XOR U5950 ( .A(n4098), .B(in[717]), .Z(n4513) );
  NAND U5951 ( .A(n4280), .B(n4099), .Z(n4100) );
  XNOR U5952 ( .A(n4513), .B(n4100), .Z(out[806]) );
  XOR U5953 ( .A(n4101), .B(in[718]), .Z(n4517) );
  NAND U5954 ( .A(n4282), .B(n4102), .Z(n4103) );
  XNOR U5955 ( .A(n4517), .B(n4103), .Z(out[807]) );
  XOR U5956 ( .A(n4104), .B(in[719]), .Z(n4521) );
  NAND U5957 ( .A(n4284), .B(n4105), .Z(n4106) );
  XNOR U5958 ( .A(n4521), .B(n4106), .Z(out[808]) );
  XOR U5959 ( .A(n4107), .B(in[720]), .Z(n4525) );
  NAND U5960 ( .A(n4286), .B(n4108), .Z(n4109) );
  XNOR U5961 ( .A(n4525), .B(n4109), .Z(out[809]) );
  NOR U5962 ( .A(n4111), .B(n4110), .Z(n4112) );
  XNOR U5963 ( .A(n4113), .B(n4112), .Z(out[80]) );
  XOR U5964 ( .A(n4114), .B(in[721]), .Z(n4529) );
  NAND U5965 ( .A(n4288), .B(n4115), .Z(n4116) );
  XNOR U5966 ( .A(n4529), .B(n4116), .Z(out[810]) );
  XOR U5967 ( .A(n4117), .B(in[722]), .Z(n4533) );
  NAND U5968 ( .A(n4290), .B(n4118), .Z(n4119) );
  XNOR U5969 ( .A(n4533), .B(n4119), .Z(out[811]) );
  XOR U5970 ( .A(n4120), .B(in[723]), .Z(n4541) );
  NAND U5971 ( .A(n4292), .B(n4121), .Z(n4122) );
  XNOR U5972 ( .A(n4541), .B(n4122), .Z(out[812]) );
  XOR U5973 ( .A(in[724]), .B(n4123), .Z(n4545) );
  NAND U5974 ( .A(n4294), .B(n4124), .Z(n4125) );
  XNOR U5975 ( .A(n4545), .B(n4125), .Z(out[813]) );
  XOR U5976 ( .A(in[725]), .B(n4126), .Z(n4549) );
  NAND U5977 ( .A(n4296), .B(n4127), .Z(n4128) );
  XNOR U5978 ( .A(n4549), .B(n4128), .Z(out[814]) );
  XOR U5979 ( .A(in[726]), .B(n4129), .Z(n4553) );
  NAND U5980 ( .A(n4298), .B(n4130), .Z(n4131) );
  XNOR U5981 ( .A(n4553), .B(n4131), .Z(out[815]) );
  XOR U5982 ( .A(in[727]), .B(n4132), .Z(n4557) );
  NAND U5983 ( .A(n4304), .B(n4133), .Z(n4134) );
  XNOR U5984 ( .A(n4557), .B(n4134), .Z(out[816]) );
  XOR U5985 ( .A(in[728]), .B(n4135), .Z(n4561) );
  NAND U5986 ( .A(n4306), .B(n4136), .Z(n4137) );
  XNOR U5987 ( .A(n4561), .B(n4137), .Z(out[817]) );
  XOR U5988 ( .A(in[729]), .B(n4138), .Z(n4565) );
  NAND U5989 ( .A(n4308), .B(n4139), .Z(n4140) );
  XNOR U5990 ( .A(n4565), .B(n4140), .Z(out[818]) );
  XOR U5991 ( .A(in[730]), .B(n4141), .Z(n4569) );
  NAND U5992 ( .A(n4310), .B(n4142), .Z(n4143) );
  XNOR U5993 ( .A(n4569), .B(n4143), .Z(out[819]) );
  NOR U5994 ( .A(n4145), .B(n4144), .Z(n4146) );
  XNOR U5995 ( .A(n4147), .B(n4146), .Z(out[81]) );
  XOR U5996 ( .A(in[731]), .B(n4148), .Z(n4573) );
  NAND U5997 ( .A(n4312), .B(n4149), .Z(n4150) );
  XNOR U5998 ( .A(n4573), .B(n4150), .Z(out[820]) );
  XOR U5999 ( .A(in[732]), .B(n4151), .Z(n4577) );
  NAND U6000 ( .A(n4314), .B(n4152), .Z(n4153) );
  XNOR U6001 ( .A(n4577), .B(n4153), .Z(out[821]) );
  XOR U6002 ( .A(in[733]), .B(n4154), .Z(n4585) );
  NAND U6003 ( .A(n4316), .B(n4155), .Z(n4156) );
  XNOR U6004 ( .A(n4585), .B(n4156), .Z(out[822]) );
  XOR U6005 ( .A(in[734]), .B(n4157), .Z(n4589) );
  NAND U6006 ( .A(n4318), .B(n4158), .Z(n4159) );
  XNOR U6007 ( .A(n4589), .B(n4159), .Z(out[823]) );
  XOR U6008 ( .A(in[735]), .B(n4160), .Z(n4593) );
  NAND U6009 ( .A(n4320), .B(n4161), .Z(n4162) );
  XNOR U6010 ( .A(n4593), .B(n4162), .Z(out[824]) );
  XOR U6011 ( .A(in[736]), .B(n4163), .Z(n4597) );
  NAND U6012 ( .A(n4322), .B(n4164), .Z(n4165) );
  XNOR U6013 ( .A(n4597), .B(n4165), .Z(out[825]) );
  XOR U6014 ( .A(in[737]), .B(n4166), .Z(n4601) );
  NAND U6015 ( .A(n4328), .B(n4167), .Z(n4168) );
  XNOR U6016 ( .A(n4601), .B(n4168), .Z(out[826]) );
  XOR U6017 ( .A(in[738]), .B(n4169), .Z(n4605) );
  NAND U6018 ( .A(n4330), .B(n4170), .Z(n4171) );
  XNOR U6019 ( .A(n4605), .B(n4171), .Z(out[827]) );
  XOR U6020 ( .A(in[739]), .B(n4172), .Z(n4609) );
  NAND U6021 ( .A(n4332), .B(n4173), .Z(n4174) );
  XNOR U6022 ( .A(n4609), .B(n4174), .Z(out[828]) );
  XNOR U6023 ( .A(in[740]), .B(n4175), .Z(n4613) );
  NAND U6024 ( .A(n4334), .B(n4176), .Z(n4177) );
  XNOR U6025 ( .A(n4613), .B(n4177), .Z(out[829]) );
  NOR U6026 ( .A(n4179), .B(n4178), .Z(n4180) );
  XNOR U6027 ( .A(n4181), .B(n4180), .Z(out[82]) );
  XNOR U6028 ( .A(in[741]), .B(n4182), .Z(n4617) );
  NAND U6029 ( .A(n4336), .B(n4183), .Z(n4184) );
  XNOR U6030 ( .A(n4617), .B(n4184), .Z(out[830]) );
  XNOR U6031 ( .A(in[742]), .B(n4185), .Z(n4621) );
  NAND U6032 ( .A(n4338), .B(n4186), .Z(n4187) );
  XNOR U6033 ( .A(n4621), .B(n4187), .Z(out[831]) );
  OR U6034 ( .A(n4341), .B(n4188), .Z(n4189) );
  XNOR U6035 ( .A(n4340), .B(n4189), .Z(out[832]) );
  OR U6036 ( .A(n4345), .B(n4190), .Z(n4191) );
  XNOR U6037 ( .A(n4344), .B(n4191), .Z(out[833]) );
  OR U6038 ( .A(n4349), .B(n4192), .Z(n4193) );
  XNOR U6039 ( .A(n4348), .B(n4193), .Z(out[834]) );
  OR U6040 ( .A(n4353), .B(n4194), .Z(n4195) );
  XNOR U6041 ( .A(n4352), .B(n4195), .Z(out[835]) );
  OR U6042 ( .A(n4365), .B(n4196), .Z(n4197) );
  XNOR U6043 ( .A(n4364), .B(n4197), .Z(out[836]) );
  OR U6044 ( .A(n4369), .B(n4198), .Z(n4199) );
  XNOR U6045 ( .A(n4368), .B(n4199), .Z(out[837]) );
  OR U6046 ( .A(n4373), .B(n4200), .Z(n4201) );
  XNOR U6047 ( .A(n4372), .B(n4201), .Z(out[838]) );
  OR U6048 ( .A(n4377), .B(n4202), .Z(n4203) );
  XNOR U6049 ( .A(n4376), .B(n4203), .Z(out[839]) );
  NOR U6050 ( .A(n4205), .B(n4204), .Z(n4206) );
  XNOR U6051 ( .A(n4207), .B(n4206), .Z(out[83]) );
  OR U6052 ( .A(n4381), .B(n4208), .Z(n4209) );
  XNOR U6053 ( .A(n4380), .B(n4209), .Z(out[840]) );
  OR U6054 ( .A(n4385), .B(n4210), .Z(n4211) );
  XNOR U6055 ( .A(n4384), .B(n4211), .Z(out[841]) );
  OR U6056 ( .A(n4389), .B(n4212), .Z(n4213) );
  XNOR U6057 ( .A(n4388), .B(n4213), .Z(out[842]) );
  OR U6058 ( .A(n4393), .B(n4214), .Z(n4215) );
  XNOR U6059 ( .A(n4392), .B(n4215), .Z(out[843]) );
  OR U6060 ( .A(n4397), .B(n4216), .Z(n4217) );
  XNOR U6061 ( .A(n4396), .B(n4217), .Z(out[844]) );
  OR U6062 ( .A(n4401), .B(n4218), .Z(n4219) );
  XNOR U6063 ( .A(n4400), .B(n4219), .Z(out[845]) );
  OR U6064 ( .A(n4409), .B(n4220), .Z(n4221) );
  XNOR U6065 ( .A(n4408), .B(n4221), .Z(out[846]) );
  OR U6066 ( .A(n4413), .B(n4222), .Z(n4223) );
  XNOR U6067 ( .A(n4412), .B(n4223), .Z(out[847]) );
  OR U6068 ( .A(n4417), .B(n4224), .Z(n4225) );
  XNOR U6069 ( .A(n4416), .B(n4225), .Z(out[848]) );
  OR U6070 ( .A(n4421), .B(n4226), .Z(n4227) );
  XNOR U6071 ( .A(n4420), .B(n4227), .Z(out[849]) );
  NOR U6072 ( .A(n4229), .B(n4228), .Z(n4230) );
  XNOR U6073 ( .A(n4231), .B(n4230), .Z(out[84]) );
  OR U6074 ( .A(n4425), .B(n4232), .Z(n4233) );
  XNOR U6075 ( .A(n4424), .B(n4233), .Z(out[850]) );
  OR U6076 ( .A(n4429), .B(n4234), .Z(n4235) );
  XNOR U6077 ( .A(n4428), .B(n4235), .Z(out[851]) );
  OR U6078 ( .A(n4433), .B(n4236), .Z(n4237) );
  XNOR U6079 ( .A(n4432), .B(n4237), .Z(out[852]) );
  OR U6080 ( .A(n4437), .B(n4238), .Z(n4239) );
  XNOR U6081 ( .A(n4436), .B(n4239), .Z(out[853]) );
  OR U6082 ( .A(n4441), .B(n4240), .Z(n4241) );
  XNOR U6083 ( .A(n4440), .B(n4241), .Z(out[854]) );
  OR U6084 ( .A(n4445), .B(n4242), .Z(n4243) );
  XNOR U6085 ( .A(n4444), .B(n4243), .Z(out[855]) );
  OR U6086 ( .A(n4453), .B(n4244), .Z(n4245) );
  XNOR U6087 ( .A(n4452), .B(n4245), .Z(out[856]) );
  OR U6088 ( .A(n4457), .B(n4246), .Z(n4247) );
  XNOR U6089 ( .A(n4456), .B(n4247), .Z(out[857]) );
  OR U6090 ( .A(n4461), .B(n4248), .Z(n4249) );
  XNOR U6091 ( .A(n4460), .B(n4249), .Z(out[858]) );
  OR U6092 ( .A(n4465), .B(n4250), .Z(n4251) );
  XNOR U6093 ( .A(n4464), .B(n4251), .Z(out[859]) );
  NOR U6094 ( .A(n4253), .B(n4252), .Z(n4254) );
  XNOR U6095 ( .A(n4255), .B(n4254), .Z(out[85]) );
  OR U6096 ( .A(n4469), .B(n4256), .Z(n4257) );
  XNOR U6097 ( .A(n4468), .B(n4257), .Z(out[860]) );
  OR U6098 ( .A(n4473), .B(n4258), .Z(n4259) );
  XNOR U6099 ( .A(n4472), .B(n4259), .Z(out[861]) );
  OR U6100 ( .A(n4477), .B(n4260), .Z(n4261) );
  XNOR U6101 ( .A(n4476), .B(n4261), .Z(out[862]) );
  OR U6102 ( .A(n4481), .B(n4262), .Z(n4263) );
  XNOR U6103 ( .A(n4480), .B(n4263), .Z(out[863]) );
  OR U6104 ( .A(n4485), .B(n4264), .Z(n4265) );
  XNOR U6105 ( .A(n4484), .B(n4265), .Z(out[864]) );
  OR U6106 ( .A(n4489), .B(n4266), .Z(n4267) );
  XNOR U6107 ( .A(n4488), .B(n4267), .Z(out[865]) );
  OR U6108 ( .A(n4497), .B(n4268), .Z(n4269) );
  XNOR U6109 ( .A(n4496), .B(n4269), .Z(out[866]) );
  OR U6110 ( .A(n4501), .B(n4270), .Z(n4271) );
  XNOR U6111 ( .A(n4500), .B(n4271), .Z(out[867]) );
  OR U6112 ( .A(n4505), .B(n4272), .Z(n4273) );
  XNOR U6113 ( .A(n4504), .B(n4273), .Z(out[868]) );
  OR U6114 ( .A(n4509), .B(n4274), .Z(n4275) );
  XNOR U6115 ( .A(n4508), .B(n4275), .Z(out[869]) );
  NOR U6116 ( .A(n4277), .B(n4276), .Z(n4278) );
  XNOR U6117 ( .A(n4279), .B(n4278), .Z(out[86]) );
  OR U6118 ( .A(n4513), .B(n4280), .Z(n4281) );
  XNOR U6119 ( .A(n4512), .B(n4281), .Z(out[870]) );
  OR U6120 ( .A(n4517), .B(n4282), .Z(n4283) );
  XNOR U6121 ( .A(n4516), .B(n4283), .Z(out[871]) );
  OR U6122 ( .A(n4521), .B(n4284), .Z(n4285) );
  XNOR U6123 ( .A(n4520), .B(n4285), .Z(out[872]) );
  OR U6124 ( .A(n4525), .B(n4286), .Z(n4287) );
  XNOR U6125 ( .A(n4524), .B(n4287), .Z(out[873]) );
  OR U6126 ( .A(n4529), .B(n4288), .Z(n4289) );
  XNOR U6127 ( .A(n4528), .B(n4289), .Z(out[874]) );
  OR U6128 ( .A(n4533), .B(n4290), .Z(n4291) );
  XNOR U6129 ( .A(n4532), .B(n4291), .Z(out[875]) );
  OR U6130 ( .A(n4541), .B(n4292), .Z(n4293) );
  XNOR U6131 ( .A(n4540), .B(n4293), .Z(out[876]) );
  OR U6132 ( .A(n4545), .B(n4294), .Z(n4295) );
  XNOR U6133 ( .A(n4544), .B(n4295), .Z(out[877]) );
  OR U6134 ( .A(n4549), .B(n4296), .Z(n4297) );
  XNOR U6135 ( .A(n4548), .B(n4297), .Z(out[878]) );
  OR U6136 ( .A(n4553), .B(n4298), .Z(n4299) );
  XNOR U6137 ( .A(n4552), .B(n4299), .Z(out[879]) );
  NOR U6138 ( .A(n4301), .B(n4300), .Z(n4302) );
  XNOR U6139 ( .A(n4303), .B(n4302), .Z(out[87]) );
  OR U6140 ( .A(n4557), .B(n4304), .Z(n4305) );
  XNOR U6141 ( .A(n4556), .B(n4305), .Z(out[880]) );
  OR U6142 ( .A(n4561), .B(n4306), .Z(n4307) );
  XNOR U6143 ( .A(n4560), .B(n4307), .Z(out[881]) );
  OR U6144 ( .A(n4565), .B(n4308), .Z(n4309) );
  XNOR U6145 ( .A(n4564), .B(n4309), .Z(out[882]) );
  OR U6146 ( .A(n4569), .B(n4310), .Z(n4311) );
  XNOR U6147 ( .A(n4568), .B(n4311), .Z(out[883]) );
  OR U6148 ( .A(n4573), .B(n4312), .Z(n4313) );
  XNOR U6149 ( .A(n4572), .B(n4313), .Z(out[884]) );
  OR U6150 ( .A(n4577), .B(n4314), .Z(n4315) );
  XNOR U6151 ( .A(n4576), .B(n4315), .Z(out[885]) );
  OR U6152 ( .A(n4585), .B(n4316), .Z(n4317) );
  XNOR U6153 ( .A(n4584), .B(n4317), .Z(out[886]) );
  OR U6154 ( .A(n4589), .B(n4318), .Z(n4319) );
  XNOR U6155 ( .A(n4588), .B(n4319), .Z(out[887]) );
  OR U6156 ( .A(n4593), .B(n4320), .Z(n4321) );
  XNOR U6157 ( .A(n4592), .B(n4321), .Z(out[888]) );
  OR U6158 ( .A(n4597), .B(n4322), .Z(n4323) );
  XNOR U6159 ( .A(n4596), .B(n4323), .Z(out[889]) );
  NOR U6160 ( .A(n4325), .B(n4324), .Z(n4326) );
  XNOR U6161 ( .A(n4327), .B(n4326), .Z(out[88]) );
  OR U6162 ( .A(n4601), .B(n4328), .Z(n4329) );
  XNOR U6163 ( .A(n4600), .B(n4329), .Z(out[890]) );
  OR U6164 ( .A(n4605), .B(n4330), .Z(n4331) );
  XNOR U6165 ( .A(n4604), .B(n4331), .Z(out[891]) );
  OR U6166 ( .A(n4609), .B(n4332), .Z(n4333) );
  XNOR U6167 ( .A(n4608), .B(n4333), .Z(out[892]) );
  OR U6168 ( .A(n4613), .B(n4334), .Z(n4335) );
  XNOR U6169 ( .A(n4612), .B(n4335), .Z(out[893]) );
  OR U6170 ( .A(n4617), .B(n4336), .Z(n4337) );
  XNOR U6171 ( .A(n4616), .B(n4337), .Z(out[894]) );
  OR U6172 ( .A(n4621), .B(n4338), .Z(n4339) );
  XNOR U6173 ( .A(n4620), .B(n4339), .Z(out[895]) );
  ANDN U6174 ( .B(n4341), .A(n4340), .Z(n4342) );
  XNOR U6175 ( .A(n4343), .B(n4342), .Z(out[896]) );
  ANDN U6176 ( .B(n4345), .A(n4344), .Z(n4346) );
  XNOR U6177 ( .A(n4347), .B(n4346), .Z(out[897]) );
  ANDN U6178 ( .B(n4349), .A(n4348), .Z(n4350) );
  XNOR U6179 ( .A(n4351), .B(n4350), .Z(out[898]) );
  ANDN U6180 ( .B(n4353), .A(n4352), .Z(n4354) );
  XNOR U6181 ( .A(n4355), .B(n4354), .Z(out[899]) );
  NOR U6182 ( .A(n4357), .B(n4356), .Z(n4358) );
  XNOR U6183 ( .A(n4359), .B(n4358), .Z(out[89]) );
  OR U6184 ( .A(n4361), .B(n4360), .Z(n4362) );
  XNOR U6185 ( .A(n4363), .B(n4362), .Z(out[8]) );
  ANDN U6186 ( .B(n4365), .A(n4364), .Z(n4366) );
  XNOR U6187 ( .A(n4367), .B(n4366), .Z(out[900]) );
  ANDN U6188 ( .B(n4369), .A(n4368), .Z(n4370) );
  XNOR U6189 ( .A(n4371), .B(n4370), .Z(out[901]) );
  ANDN U6190 ( .B(n4373), .A(n4372), .Z(n4374) );
  XNOR U6191 ( .A(n4375), .B(n4374), .Z(out[902]) );
  ANDN U6192 ( .B(n4377), .A(n4376), .Z(n4378) );
  XNOR U6193 ( .A(n4379), .B(n4378), .Z(out[903]) );
  ANDN U6194 ( .B(n4381), .A(n4380), .Z(n4382) );
  XNOR U6195 ( .A(n4383), .B(n4382), .Z(out[904]) );
  ANDN U6196 ( .B(n4385), .A(n4384), .Z(n4386) );
  XNOR U6197 ( .A(n4387), .B(n4386), .Z(out[905]) );
  ANDN U6198 ( .B(n4389), .A(n4388), .Z(n4390) );
  XNOR U6199 ( .A(n4391), .B(n4390), .Z(out[906]) );
  ANDN U6200 ( .B(n4393), .A(n4392), .Z(n4394) );
  XNOR U6201 ( .A(n4395), .B(n4394), .Z(out[907]) );
  ANDN U6202 ( .B(n4397), .A(n4396), .Z(n4398) );
  XNOR U6203 ( .A(n4399), .B(n4398), .Z(out[908]) );
  ANDN U6204 ( .B(n4401), .A(n4400), .Z(n4402) );
  XNOR U6205 ( .A(n4403), .B(n4402), .Z(out[909]) );
  NOR U6206 ( .A(n4405), .B(n4404), .Z(n4406) );
  XNOR U6207 ( .A(n4407), .B(n4406), .Z(out[90]) );
  ANDN U6208 ( .B(n4409), .A(n4408), .Z(n4410) );
  XNOR U6209 ( .A(n4411), .B(n4410), .Z(out[910]) );
  ANDN U6210 ( .B(n4413), .A(n4412), .Z(n4414) );
  XNOR U6211 ( .A(n4415), .B(n4414), .Z(out[911]) );
  ANDN U6212 ( .B(n4417), .A(n4416), .Z(n4418) );
  XNOR U6213 ( .A(n4419), .B(n4418), .Z(out[912]) );
  ANDN U6214 ( .B(n4421), .A(n4420), .Z(n4422) );
  XNOR U6215 ( .A(n4423), .B(n4422), .Z(out[913]) );
  ANDN U6216 ( .B(n4425), .A(n4424), .Z(n4426) );
  XNOR U6217 ( .A(n4427), .B(n4426), .Z(out[914]) );
  ANDN U6218 ( .B(n4429), .A(n4428), .Z(n4430) );
  XNOR U6219 ( .A(n4431), .B(n4430), .Z(out[915]) );
  ANDN U6220 ( .B(n4433), .A(n4432), .Z(n4434) );
  XNOR U6221 ( .A(n4435), .B(n4434), .Z(out[916]) );
  ANDN U6222 ( .B(n4437), .A(n4436), .Z(n4438) );
  XNOR U6223 ( .A(n4439), .B(n4438), .Z(out[917]) );
  ANDN U6224 ( .B(n4441), .A(n4440), .Z(n4442) );
  XNOR U6225 ( .A(n4443), .B(n4442), .Z(out[918]) );
  ANDN U6226 ( .B(n4445), .A(n4444), .Z(n4446) );
  XNOR U6227 ( .A(n4447), .B(n4446), .Z(out[919]) );
  NOR U6228 ( .A(n4449), .B(n4448), .Z(n4450) );
  XNOR U6229 ( .A(n4451), .B(n4450), .Z(out[91]) );
  ANDN U6230 ( .B(n4453), .A(n4452), .Z(n4454) );
  XNOR U6231 ( .A(n4455), .B(n4454), .Z(out[920]) );
  ANDN U6232 ( .B(n4457), .A(n4456), .Z(n4458) );
  XNOR U6233 ( .A(n4459), .B(n4458), .Z(out[921]) );
  ANDN U6234 ( .B(n4461), .A(n4460), .Z(n4462) );
  XNOR U6235 ( .A(n4463), .B(n4462), .Z(out[922]) );
  ANDN U6236 ( .B(n4465), .A(n4464), .Z(n4466) );
  XNOR U6237 ( .A(n4467), .B(n4466), .Z(out[923]) );
  ANDN U6238 ( .B(n4469), .A(n4468), .Z(n4470) );
  XNOR U6239 ( .A(n4471), .B(n4470), .Z(out[924]) );
  ANDN U6240 ( .B(n4473), .A(n4472), .Z(n4474) );
  XNOR U6241 ( .A(n4475), .B(n4474), .Z(out[925]) );
  ANDN U6242 ( .B(n4477), .A(n4476), .Z(n4478) );
  XNOR U6243 ( .A(n4479), .B(n4478), .Z(out[926]) );
  ANDN U6244 ( .B(n4481), .A(n4480), .Z(n4482) );
  XNOR U6245 ( .A(n4483), .B(n4482), .Z(out[927]) );
  ANDN U6246 ( .B(n4485), .A(n4484), .Z(n4486) );
  XNOR U6247 ( .A(n4487), .B(n4486), .Z(out[928]) );
  ANDN U6248 ( .B(n4489), .A(n4488), .Z(n4490) );
  XNOR U6249 ( .A(n4491), .B(n4490), .Z(out[929]) );
  ANDN U6250 ( .B(n4493), .A(n4492), .Z(n4494) );
  XNOR U6251 ( .A(n4495), .B(n4494), .Z(out[92]) );
  ANDN U6252 ( .B(n4497), .A(n4496), .Z(n4498) );
  XNOR U6253 ( .A(n4499), .B(n4498), .Z(out[930]) );
  ANDN U6254 ( .B(n4501), .A(n4500), .Z(n4502) );
  XNOR U6255 ( .A(n4503), .B(n4502), .Z(out[931]) );
  ANDN U6256 ( .B(n4505), .A(n4504), .Z(n4506) );
  XNOR U6257 ( .A(n4507), .B(n4506), .Z(out[932]) );
  ANDN U6258 ( .B(n4509), .A(n4508), .Z(n4510) );
  XNOR U6259 ( .A(n4511), .B(n4510), .Z(out[933]) );
  ANDN U6260 ( .B(n4513), .A(n4512), .Z(n4514) );
  XNOR U6261 ( .A(n4515), .B(n4514), .Z(out[934]) );
  ANDN U6262 ( .B(n4517), .A(n4516), .Z(n4518) );
  XNOR U6263 ( .A(n4519), .B(n4518), .Z(out[935]) );
  ANDN U6264 ( .B(n4521), .A(n4520), .Z(n4522) );
  XNOR U6265 ( .A(n4523), .B(n4522), .Z(out[936]) );
  ANDN U6266 ( .B(n4525), .A(n4524), .Z(n4526) );
  XNOR U6267 ( .A(n4527), .B(n4526), .Z(out[937]) );
  ANDN U6268 ( .B(n4529), .A(n4528), .Z(n4530) );
  XNOR U6269 ( .A(n4531), .B(n4530), .Z(out[938]) );
  ANDN U6270 ( .B(n4533), .A(n4532), .Z(n4534) );
  XNOR U6271 ( .A(n4535), .B(n4534), .Z(out[939]) );
  ANDN U6272 ( .B(n4537), .A(n4536), .Z(n4538) );
  XNOR U6273 ( .A(n4539), .B(n4538), .Z(out[93]) );
  ANDN U6274 ( .B(n4541), .A(n4540), .Z(n4542) );
  XNOR U6275 ( .A(n4543), .B(n4542), .Z(out[940]) );
  ANDN U6276 ( .B(n4545), .A(n4544), .Z(n4546) );
  XNOR U6277 ( .A(n4547), .B(n4546), .Z(out[941]) );
  ANDN U6278 ( .B(n4549), .A(n4548), .Z(n4550) );
  XNOR U6279 ( .A(n4551), .B(n4550), .Z(out[942]) );
  ANDN U6280 ( .B(n4553), .A(n4552), .Z(n4554) );
  XNOR U6281 ( .A(n4555), .B(n4554), .Z(out[943]) );
  ANDN U6282 ( .B(n4557), .A(n4556), .Z(n4558) );
  XNOR U6283 ( .A(n4559), .B(n4558), .Z(out[944]) );
  ANDN U6284 ( .B(n4561), .A(n4560), .Z(n4562) );
  XNOR U6285 ( .A(n4563), .B(n4562), .Z(out[945]) );
  ANDN U6286 ( .B(n4565), .A(n4564), .Z(n4566) );
  XNOR U6287 ( .A(n4567), .B(n4566), .Z(out[946]) );
  ANDN U6288 ( .B(n4569), .A(n4568), .Z(n4570) );
  XNOR U6289 ( .A(n4571), .B(n4570), .Z(out[947]) );
  ANDN U6290 ( .B(n4573), .A(n4572), .Z(n4574) );
  XNOR U6291 ( .A(n4575), .B(n4574), .Z(out[948]) );
  ANDN U6292 ( .B(n4577), .A(n4576), .Z(n4578) );
  XNOR U6293 ( .A(n4579), .B(n4578), .Z(out[949]) );
  ANDN U6294 ( .B(n4581), .A(n4580), .Z(n4582) );
  XNOR U6295 ( .A(n4583), .B(n4582), .Z(out[94]) );
  ANDN U6296 ( .B(n4585), .A(n4584), .Z(n4586) );
  XNOR U6297 ( .A(n4587), .B(n4586), .Z(out[950]) );
  ANDN U6298 ( .B(n4589), .A(n4588), .Z(n4590) );
  XNOR U6299 ( .A(n4591), .B(n4590), .Z(out[951]) );
  ANDN U6300 ( .B(n4593), .A(n4592), .Z(n4594) );
  XNOR U6301 ( .A(n4595), .B(n4594), .Z(out[952]) );
  ANDN U6302 ( .B(n4597), .A(n4596), .Z(n4598) );
  XNOR U6303 ( .A(n4599), .B(n4598), .Z(out[953]) );
  ANDN U6304 ( .B(n4601), .A(n4600), .Z(n4602) );
  XNOR U6305 ( .A(n4603), .B(n4602), .Z(out[954]) );
  ANDN U6306 ( .B(n4605), .A(n4604), .Z(n4606) );
  XNOR U6307 ( .A(n4607), .B(n4606), .Z(out[955]) );
  ANDN U6308 ( .B(n4609), .A(n4608), .Z(n4610) );
  XNOR U6309 ( .A(n4611), .B(n4610), .Z(out[956]) );
  ANDN U6310 ( .B(n4613), .A(n4612), .Z(n4614) );
  XNOR U6311 ( .A(n4615), .B(n4614), .Z(out[957]) );
  ANDN U6312 ( .B(n4617), .A(n4616), .Z(n4618) );
  XNOR U6313 ( .A(n4619), .B(n4618), .Z(out[958]) );
  ANDN U6314 ( .B(n4621), .A(n4620), .Z(n4622) );
  XNOR U6315 ( .A(n4623), .B(n4622), .Z(out[959]) );
  ANDN U6316 ( .B(n4625), .A(n4624), .Z(n4626) );
  XNOR U6317 ( .A(n4627), .B(n4626), .Z(out[95]) );
  ANDN U6318 ( .B(n4629), .A(n4628), .Z(n4630) );
  XNOR U6319 ( .A(n4631), .B(n4630), .Z(out[960]) );
  ANDN U6320 ( .B(n4633), .A(n4632), .Z(n4634) );
  XNOR U6321 ( .A(n4635), .B(n4634), .Z(out[961]) );
  ANDN U6322 ( .B(n4637), .A(n4636), .Z(n4638) );
  XNOR U6323 ( .A(n4639), .B(n4638), .Z(out[962]) );
  ANDN U6324 ( .B(n4641), .A(n4640), .Z(n4642) );
  XNOR U6325 ( .A(n4643), .B(n4642), .Z(out[963]) );
  ANDN U6326 ( .B(n4645), .A(n4644), .Z(n4646) );
  XNOR U6327 ( .A(n4647), .B(n4646), .Z(out[964]) );
  ANDN U6328 ( .B(n4649), .A(n4648), .Z(n4650) );
  XNOR U6329 ( .A(n4651), .B(n4650), .Z(out[965]) );
  ANDN U6330 ( .B(n4653), .A(n4652), .Z(n4654) );
  XNOR U6331 ( .A(n4655), .B(n4654), .Z(out[966]) );
  ANDN U6332 ( .B(n4657), .A(n4656), .Z(n4658) );
  XNOR U6333 ( .A(n4659), .B(n4658), .Z(out[967]) );
  ANDN U6334 ( .B(n4661), .A(n4660), .Z(n4662) );
  XNOR U6335 ( .A(n4663), .B(n4662), .Z(out[968]) );
  ANDN U6336 ( .B(n4665), .A(n4664), .Z(n4666) );
  XNOR U6337 ( .A(n4667), .B(n4666), .Z(out[969]) );
  ANDN U6338 ( .B(n4669), .A(n4668), .Z(n4670) );
  XNOR U6339 ( .A(n4671), .B(n4670), .Z(out[96]) );
  ANDN U6340 ( .B(n4673), .A(n4672), .Z(n4674) );
  XNOR U6341 ( .A(n4675), .B(n4674), .Z(out[970]) );
  ANDN U6342 ( .B(n4677), .A(n4676), .Z(n4678) );
  XNOR U6343 ( .A(n4679), .B(n4678), .Z(out[971]) );
  ANDN U6344 ( .B(n4681), .A(n4680), .Z(n4682) );
  XNOR U6345 ( .A(n4683), .B(n4682), .Z(out[972]) );
  ANDN U6346 ( .B(n4685), .A(n4684), .Z(n4686) );
  XNOR U6347 ( .A(n4687), .B(n4686), .Z(out[973]) );
  ANDN U6348 ( .B(n4689), .A(n4688), .Z(n4690) );
  XNOR U6349 ( .A(n4691), .B(n4690), .Z(out[974]) );
  ANDN U6350 ( .B(n4693), .A(n4692), .Z(n4694) );
  XNOR U6351 ( .A(n4695), .B(n4694), .Z(out[975]) );
  ANDN U6352 ( .B(n4697), .A(n4696), .Z(n4698) );
  XNOR U6353 ( .A(n4699), .B(n4698), .Z(out[976]) );
  ANDN U6354 ( .B(n4701), .A(n4700), .Z(n4702) );
  XNOR U6355 ( .A(n4703), .B(n4702), .Z(out[977]) );
  ANDN U6356 ( .B(n4705), .A(n4704), .Z(n4706) );
  XNOR U6357 ( .A(n4707), .B(n4706), .Z(out[978]) );
  ANDN U6358 ( .B(n4709), .A(n4708), .Z(n4710) );
  XNOR U6359 ( .A(n4711), .B(n4710), .Z(out[979]) );
  ANDN U6360 ( .B(n4713), .A(n4712), .Z(n4714) );
  XNOR U6361 ( .A(n4715), .B(n4714), .Z(out[97]) );
  ANDN U6362 ( .B(n4717), .A(n4716), .Z(n4718) );
  XNOR U6363 ( .A(n4719), .B(n4718), .Z(out[980]) );
  ANDN U6364 ( .B(n4721), .A(n4720), .Z(n4722) );
  XNOR U6365 ( .A(n4723), .B(n4722), .Z(out[981]) );
  ANDN U6366 ( .B(n4725), .A(n4724), .Z(n4726) );
  XNOR U6367 ( .A(n4727), .B(n4726), .Z(out[982]) );
  ANDN U6368 ( .B(n4729), .A(n4728), .Z(n4730) );
  XNOR U6369 ( .A(n4731), .B(n4730), .Z(out[983]) );
  ANDN U6370 ( .B(n4733), .A(n4732), .Z(n4734) );
  XNOR U6371 ( .A(n4735), .B(n4734), .Z(out[984]) );
  ANDN U6372 ( .B(n4737), .A(n4736), .Z(n4738) );
  XNOR U6373 ( .A(n4739), .B(n4738), .Z(out[985]) );
  ANDN U6374 ( .B(n4741), .A(n4740), .Z(n4742) );
  XNOR U6375 ( .A(n4743), .B(n4742), .Z(out[986]) );
  ANDN U6376 ( .B(n4745), .A(n4744), .Z(n4746) );
  XNOR U6377 ( .A(n4747), .B(n4746), .Z(out[987]) );
  ANDN U6378 ( .B(n4749), .A(n4748), .Z(n4750) );
  XNOR U6379 ( .A(n4751), .B(n4750), .Z(out[988]) );
  ANDN U6380 ( .B(n4753), .A(n4752), .Z(n4754) );
  XNOR U6381 ( .A(n4755), .B(n4754), .Z(out[989]) );
  ANDN U6382 ( .B(n4757), .A(n4756), .Z(n4758) );
  XNOR U6383 ( .A(n4759), .B(n4758), .Z(out[98]) );
  ANDN U6384 ( .B(n4761), .A(n4760), .Z(n4762) );
  XNOR U6385 ( .A(n4763), .B(n4762), .Z(out[990]) );
  ANDN U6386 ( .B(n4765), .A(n4764), .Z(n4766) );
  XNOR U6387 ( .A(n4767), .B(n4766), .Z(out[991]) );
  ANDN U6388 ( .B(n4769), .A(n4768), .Z(n4770) );
  XNOR U6389 ( .A(n4771), .B(n4770), .Z(out[992]) );
  ANDN U6390 ( .B(n4773), .A(n4772), .Z(n4774) );
  XNOR U6391 ( .A(n4775), .B(n4774), .Z(out[993]) );
  ANDN U6392 ( .B(n4777), .A(n4776), .Z(n4778) );
  XNOR U6393 ( .A(n4779), .B(n4778), .Z(out[994]) );
  ANDN U6394 ( .B(n4781), .A(n4780), .Z(n4782) );
  XNOR U6395 ( .A(n4783), .B(n4782), .Z(out[995]) );
  ANDN U6396 ( .B(n4785), .A(n4784), .Z(n4786) );
  XNOR U6397 ( .A(n4787), .B(n4786), .Z(out[996]) );
  ANDN U6398 ( .B(n4789), .A(n4788), .Z(n4790) );
  XNOR U6399 ( .A(n4791), .B(n4790), .Z(out[997]) );
  ANDN U6400 ( .B(n4793), .A(n4792), .Z(n4794) );
  XNOR U6401 ( .A(n4795), .B(n4794), .Z(out[998]) );
  ANDN U6402 ( .B(n4797), .A(n4796), .Z(n4798) );
  XNOR U6403 ( .A(n4799), .B(n4798), .Z(out[999]) );
  ANDN U6404 ( .B(n4801), .A(n4800), .Z(n4802) );
  XNOR U6405 ( .A(n4803), .B(n4802), .Z(out[99]) );
  OR U6406 ( .A(n4805), .B(n4804), .Z(n4806) );
  XNOR U6407 ( .A(n4807), .B(n4806), .Z(out[9]) );
endmodule


module sha3_seq_CC6 ( clk, rst, in, out );
  input [575:0] in;
  output [1599:0] out;
  input clk, rst;
  wire   init, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74,
         N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88,
         N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101,
         N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112,
         N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123,
         N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134,
         N135, N136, N137, N138, N139, N140, N141, N142, N143, N144, N145,
         N146, N147, N148, N149, N150, N151, N152, N153, N154, N155, N156,
         N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167,
         N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178,
         N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189,
         N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200,
         N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211,
         N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222,
         N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233,
         N234, N235, N236, N237, N238, N239, N240, N241, N242, N243, N244,
         N245, N246, N247, N248, N249, N250, N251, N252, N253, N254, N255,
         N256, N257, N258, N259, N260, N261, N262, N263, N264, N265, N266,
         N267, N268, N269, N270, N271, N272, N273, N274, N275, N276, N277,
         N278, N279, N280, N281, N282, N283, N284, N285, N286, N287, N288,
         N289, N290, N291, N292, N293, N294, N295, N296, N297, N298, N299,
         N300, N301, N302, N303, N304, N305, N306, N307, N308, N309, N310,
         N311, N312, N313, N314, N315, N316, N317, N318, N319, N320, N321,
         N322, N323, N324, N325, N326, N327, N328, N329, N330, N331, N332,
         N333, N334, N335, N336, N337, N338, N339, N340, N341, N342, N343,
         N344, N345, N346, N347, N348, N349, N350, N351, N352, N353, N354,
         N355, N356, N357, N358, N359, N360, N361, N362, N363, N364, N365,
         N366, N367, N368, N369, N370, N371, N372, N373, N374, N375, N376,
         N377, N378, N379, N380, N381, N382, N383, N384, N385, N386, N387,
         N388, N389, N390, N391, N392, N393, N394, N395, N396, N397, N398,
         N399, N400, N401, N402, N403, N404, N405, N406, N407, N408, N409,
         N410, N411, N412, N413, N414, N415, N416, N417, N418, N419, N420,
         N421, N422, N423, N424, N425, N426, N427, N428, N429, N430, N431,
         N432, N433, N434, N435, N436, N437, N438, N439, N440, N441, N442,
         N443, N444, N445, N446, N447, N448, N449, N450, N451, N452, N453,
         N454, N455, N456, N457, N458, N459, N460, N461, N462, N463, N464,
         N465, N466, N467, N468, N469, N470, N471, N472, N473, N474, N475,
         N476, N477, N478, N479, N480, N481, N482, N483, N484, N485, N486,
         N487, N488, N489, N490, N491, N492, N493, N494, N495, N496, N497,
         N498, N499, N500, N501, N502, N503, N504, N505, N506, N507, N508,
         N509, N510, N511, N512, N513, N514, N515, N516, N517, N518, N519,
         N520, N521, N522, N523, N524, N525, N526, N527, N528, N529, N530,
         N531, N532, N533, N534, N535, N536, N537, N538, N539, N540, N541,
         N542, N543, N544, N545, N546, N547, N548, N549, N550, N551, N552,
         N553, N554, N555, N556, N557, N558, N559, N560, N561, N562, N563,
         N564, N565, N566, N567, N568, N569, N570, N571, N572, N573, N574,
         N575, N576, N577, N578, N579, N580, N581, N582, N583, N584, N585,
         N586, N587, N588, N589, N590, N591, N592, N593, N594, N595, N596,
         N597, N598, N599, N600, N601, N602, N603, N604, N605, N606, N607,
         N608, N609, N610, N611, N612, N613, N614, N615, N616, N617, N618,
         N619, N620, N621, N622, N623, N624, N625, N626, N627, N628, N629,
         N630, N631, N632, N633, N634, N635, N636, N637, N638, N639, N640,
         N641, N642, N643, N644, N645, N646, N647, N648, N649, N650, N651,
         N652, N653, N654, N655, N656, N657, N658, N659, N660, N661, N662,
         N663, N664, N665, N666, N667, N668, N669, N670, N671, N672, N673,
         N674, N675, N676, N677, N678, N679, N680, N681, N682, N683, N684,
         N685, N686, N687, N688, N689, N690, N691, N692, N693, N694, N695,
         N696, N697, N698, N699, N700, N701, N702, N703, N704, N705, N706,
         N707, N708, N709, N710, N711, N712, N713, N714, N715, N716, N717,
         N718, N719, N720, N721, N722, N723, N724, N725, N726, N727, N728,
         N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739,
         N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750,
         N751, N752, N753, N754, N755, N756, N757, N758, N759, N760, N761,
         N762, N763, N764, N765, N766, N767, N768, N769, N770, N771, N772,
         N773, N774, N775, N776, N777, N778, N779, N780, N781, N782, N783,
         N784, N785, N786, N787, N788, N789, N790, N791, N792, N793, N794,
         N795, N796, N797, N798, N799, N800, N801, N802, N803, N804, N805,
         N806, N807, N808, N809, N810, N811, N812, N813, N814, N815, N816,
         N817, N818, N819, N820, N821, N822, N823, N824, N825, N826, N827,
         N828, N829, N830, N831, N832, N833, N834, N835, N836, N837, N838,
         N839, N840, N841, N842, N843, N844, N845, N846, N847, N848, N849,
         N850, N851, N852, N853, N854, N855, N856, N857, N858, N859, N860,
         N861, N862, N863, N864, N865, N866, N867, N868, N869, N870, N871,
         N872, N873, N874, N875, N876, N877, N878, N879, N880, N881, N882,
         N883, N884, N885, N886, N887, N888, N889, N890, N891, N892, N893,
         N894, N895, N896, N897, N898, N899, N900, N901, N902, N903, N904,
         N905, N906, N907, N908, N909, N910, N911, N912, N913, N914, N915,
         N916, N917, N918, N919, N920, N921, N922, N923, N924, N925, N926,
         N927, N928, N929, N930, N931, N932, N933, N934, N935, N936, N937,
         N938, N939, N940, N941, N942, N943, N944, N945, N946, N947, N948,
         N949, N950, N951, N952, N953, N954, N955, N956, N957, N958, N959,
         N960, N961, N962, N963, N964, N965, N966, N967, N968, N969, N970,
         N971, N972, N973, N974, N975, N976, N977, N978, N979, N980, N981,
         N982, N983, N984, N985, N986, N987, N988, N989, N990, N991, N992,
         N993, N994, N995, N996, N997, N998, N999, N1000, N1001, N1002, N1003,
         N1004, N1005, N1006, N1007, N1008, N1009, N1010, N1011, N1012, N1013,
         N1014, N1015, N1016, N1017, N1018, N1019, N1020, N1021, N1022, N1023,
         N1024, N1025, N1026, N1027, N1028, N1029, N1030, N1031, N1032, N1033,
         N1034, N1035, N1036, N1037, N1038, N1039, N1040, N1041, N1042, N1043,
         N1044, N1045, N1046, N1047, N1048, N1049, N1050, N1051, N1052, N1053,
         N1054, N1055, N1056, N1057, N1058, N1059, N1060, N1061, N1062, N1063,
         N1064, N1065, N1066, N1067, N1068, N1069, N1070, N1071, N1072, N1073,
         N1074, N1075, N1076, N1077, N1078, N1079, N1080, N1081, N1082, N1083,
         N1084, N1085, N1086, N1087, N1088, N1089, N1090, N1091, N1092, N1093,
         N1094, N1095, N1096, N1097, N1098, N1099, N1100, N1101, N1102, N1103,
         N1104, N1105, N1106, N1107, N1108, N1109, N1110, N1111, N1112, N1113,
         N1114, N1115, N1116, N1117, N1118, N1119, N1120, N1121, N1122, N1123,
         N1124, N1125, N1126, N1127, N1128, N1129, N1130, N1131, N1132, N1133,
         N1134, N1135, N1136, N1137, N1138, N1139, N1140, N1141, N1142, N1143,
         N1144, N1145, N1146, N1147, N1148, N1149, N1150, N1151, N1152, N1153,
         N1154, N1155, N1156, N1157, N1158, N1159, N1160, N1161, N1162, N1163,
         N1164, N1165, N1166, N1167, N1168, N1169, N1170, N1171, N1172, N1173,
         N1174, N1175, N1176, N1177, N1178, N1179, N1180, N1181, N1182, N1183,
         N1184, N1185, N1186, N1187, N1188, N1189, N1190, N1191, N1192, N1193,
         N1194, N1195, N1196, N1197, N1198, N1199, N1200, N1201, N1202, N1203,
         N1204, N1205, N1206, N1207, N1208, N1209, N1210, N1211, N1212, N1213,
         N1214, N1215, N1216, N1217, N1218, N1219, N1220, N1221, N1222, N1223,
         N1224, N1225, N1226, N1227, N1228, N1229, N1230, N1231, N1232, N1233,
         N1234, N1235, N1236, N1237, N1238, N1239, N1240, N1241, N1242, N1243,
         N1244, N1245, N1246, N1247, N1248, N1249, N1250, N1251, N1252, N1253,
         N1254, N1255, N1256, N1257, N1258, N1259, N1260, N1261, N1262, N1263,
         N1264, N1265, N1266, N1267, N1268, N1269, N1270, N1271, N1272, N1273,
         N1274, N1275, N1276, N1277, N1278, N1279, N1280, N1281, N1282, N1283,
         N1284, N1285, N1286, N1287, N1288, N1289, N1290, N1291, N1292, N1293,
         N1294, N1295, N1296, N1297, N1298, N1299, N1300, N1301, N1302, N1303,
         N1304, N1305, N1306, N1307, N1308, N1309, N1310, N1311, N1312, N1313,
         N1314, N1315, N1316, N1317, N1318, N1319, N1320, N1321, N1322, N1323,
         N1324, N1325, N1326, N1327, N1328, N1329, N1330, N1331, N1332, N1333,
         N1334, N1335, N1336, N1337, N1338, N1339, N1340, N1341, N1342, N1343,
         N1344, N1345, N1346, N1347, N1348, N1349, N1350, N1351, N1352, N1353,
         N1354, N1355, N1356, N1357, N1358, N1359, N1360, N1361, N1362, N1363,
         N1364, N1365, N1366, N1367, N1368, N1369, N1370, N1371, N1372, N1373,
         N1374, N1375, N1376, N1377, N1378, N1379, N1380, N1381, N1382, N1383,
         N1384, N1385, N1386, N1387, N1388, N1389, N1390, N1391, N1392, N1393,
         N1394, N1395, N1396, N1397, N1398, N1399, N1400, N1401, N1402, N1403,
         N1404, N1405, N1406, N1407, N1408, N1409, N1410, N1411, N1412, N1413,
         N1414, N1415, N1416, N1417, N1418, N1419, N1420, N1421, N1422, N1423,
         N1424, N1425, N1426, N1427, N1428, N1429, N1430, N1431, N1432, N1433,
         N1434, N1435, N1436, N1437, N1438, N1439, N1440, N1441, N1442, N1443,
         N1444, N1445, N1446, N1447, N1448, N1449, N1450, N1451, N1452, N1453,
         N1454, N1455, N1456, N1457, N1458, N1459, N1460, N1461, N1462, N1463,
         N1464, N1465, N1466, N1467, N1468, N1469, N1470, N1471, N1472, N1473,
         N1474, N1475, N1476, N1477, N1478, N1479, N1480, N1481, N1482, N1483,
         N1484, N1485, N1486, N1487, N1488, N1489, N1490, N1491, N1492, N1493,
         N1494, N1495, N1496, N1497, N1498, N1499, N1500, N1501, N1502, N1503,
         N1504, N1505, N1506, N1507, N1508, N1509, N1510, N1511, N1512, N1513,
         N1514, N1515, N1516, N1517, N1518, N1519, N1520, N1521, N1522, N1523,
         N1524, N1525, N1526, N1527, N1528, N1529, N1530, N1531, N1532, N1533,
         N1534, N1535, N1536, N1537, N1538, N1539, N1540, N1541, N1542, N1543,
         N1544, N1545, N1546, N1547, N1548, N1549, N1550, N1551, N1552, N1553,
         N1554, N1555, N1556, N1557, N1558, N1559, N1560, N1561, N1562, N1563,
         N1564, N1565, N1566, N1567, N1568, N1569, N1570, N1571, N1572, N1573,
         N1574, N1575, N1576, N1577, N1578, N1579, N1580, N1581, N1582, N1583,
         N1584, N1585, N1586, N1587, N1588, N1589, N1590, N1591, N1592, N1593,
         N1594, N1595, N1596, N1597, N1598, N1599, N1600, N1601, N1602, N1603,
         N1604, N1605, N1606, N1607, N1608, N1609, N1610, N1611,
         \round_in[3][1599] , \round_in[3][1598] , \round_in[3][1597] ,
         \round_in[3][1596] , \round_in[3][1595] , \round_in[3][1594] ,
         \round_in[3][1593] , \round_in[3][1592] , \round_in[3][1591] ,
         \round_in[3][1590] , \round_in[3][1589] , \round_in[3][1588] ,
         \round_in[3][1587] , \round_in[3][1586] , \round_in[3][1585] ,
         \round_in[3][1584] , \round_in[3][1583] , \round_in[3][1582] ,
         \round_in[3][1581] , \round_in[3][1580] , \round_in[3][1579] ,
         \round_in[3][1578] , \round_in[3][1577] , \round_in[3][1576] ,
         \round_in[3][1575] , \round_in[3][1574] , \round_in[3][1573] ,
         \round_in[3][1572] , \round_in[3][1571] , \round_in[3][1570] ,
         \round_in[3][1569] , \round_in[3][1568] , \round_in[3][1567] ,
         \round_in[3][1566] , \round_in[3][1565] , \round_in[3][1564] ,
         \round_in[3][1563] , \round_in[3][1562] , \round_in[3][1561] ,
         \round_in[3][1560] , \round_in[3][1559] , \round_in[3][1558] ,
         \round_in[3][1557] , \round_in[3][1556] , \round_in[3][1555] ,
         \round_in[3][1554] , \round_in[3][1553] , \round_in[3][1552] ,
         \round_in[3][1551] , \round_in[3][1550] , \round_in[3][1549] ,
         \round_in[3][1548] , \round_in[3][1547] , \round_in[3][1546] ,
         \round_in[3][1545] , \round_in[3][1544] , \round_in[3][1543] ,
         \round_in[3][1542] , \round_in[3][1541] , \round_in[3][1540] ,
         \round_in[3][1539] , \round_in[3][1538] , \round_in[3][1537] ,
         \round_in[3][1536] , \round_in[3][1535] , \round_in[3][1534] ,
         \round_in[3][1533] , \round_in[3][1532] , \round_in[3][1531] ,
         \round_in[3][1530] , \round_in[3][1529] , \round_in[3][1528] ,
         \round_in[3][1527] , \round_in[3][1526] , \round_in[3][1525] ,
         \round_in[3][1524] , \round_in[3][1523] , \round_in[3][1522] ,
         \round_in[3][1521] , \round_in[3][1520] , \round_in[3][1519] ,
         \round_in[3][1518] , \round_in[3][1517] , \round_in[3][1516] ,
         \round_in[3][1515] , \round_in[3][1514] , \round_in[3][1513] ,
         \round_in[3][1512] , \round_in[3][1511] , \round_in[3][1510] ,
         \round_in[3][1509] , \round_in[3][1508] , \round_in[3][1507] ,
         \round_in[3][1506] , \round_in[3][1505] , \round_in[3][1504] ,
         \round_in[3][1503] , \round_in[3][1502] , \round_in[3][1501] ,
         \round_in[3][1500] , \round_in[3][1499] , \round_in[3][1498] ,
         \round_in[3][1497] , \round_in[3][1496] , \round_in[3][1495] ,
         \round_in[3][1494] , \round_in[3][1493] , \round_in[3][1492] ,
         \round_in[3][1491] , \round_in[3][1490] , \round_in[3][1489] ,
         \round_in[3][1488] , \round_in[3][1487] , \round_in[3][1486] ,
         \round_in[3][1485] , \round_in[3][1484] , \round_in[3][1483] ,
         \round_in[3][1482] , \round_in[3][1481] , \round_in[3][1480] ,
         \round_in[3][1479] , \round_in[3][1478] , \round_in[3][1477] ,
         \round_in[3][1476] , \round_in[3][1475] , \round_in[3][1474] ,
         \round_in[3][1473] , \round_in[3][1472] , \round_in[3][1471] ,
         \round_in[3][1470] , \round_in[3][1469] , \round_in[3][1468] ,
         \round_in[3][1467] , \round_in[3][1466] , \round_in[3][1465] ,
         \round_in[3][1464] , \round_in[3][1463] , \round_in[3][1462] ,
         \round_in[3][1461] , \round_in[3][1460] , \round_in[3][1459] ,
         \round_in[3][1458] , \round_in[3][1457] , \round_in[3][1456] ,
         \round_in[3][1455] , \round_in[3][1454] , \round_in[3][1453] ,
         \round_in[3][1452] , \round_in[3][1451] , \round_in[3][1450] ,
         \round_in[3][1449] , \round_in[3][1448] , \round_in[3][1447] ,
         \round_in[3][1446] , \round_in[3][1445] , \round_in[3][1444] ,
         \round_in[3][1443] , \round_in[3][1442] , \round_in[3][1441] ,
         \round_in[3][1440] , \round_in[3][1439] , \round_in[3][1438] ,
         \round_in[3][1437] , \round_in[3][1436] , \round_in[3][1435] ,
         \round_in[3][1434] , \round_in[3][1433] , \round_in[3][1432] ,
         \round_in[3][1431] , \round_in[3][1430] , \round_in[3][1429] ,
         \round_in[3][1428] , \round_in[3][1427] , \round_in[3][1426] ,
         \round_in[3][1425] , \round_in[3][1424] , \round_in[3][1423] ,
         \round_in[3][1422] , \round_in[3][1421] , \round_in[3][1420] ,
         \round_in[3][1419] , \round_in[3][1418] , \round_in[3][1417] ,
         \round_in[3][1416] , \round_in[3][1415] , \round_in[3][1414] ,
         \round_in[3][1413] , \round_in[3][1412] , \round_in[3][1411] ,
         \round_in[3][1410] , \round_in[3][1409] , \round_in[3][1408] ,
         \round_in[3][1407] , \round_in[3][1406] , \round_in[3][1405] ,
         \round_in[3][1404] , \round_in[3][1403] , \round_in[3][1402] ,
         \round_in[3][1401] , \round_in[3][1400] , \round_in[3][1399] ,
         \round_in[3][1398] , \round_in[3][1397] , \round_in[3][1396] ,
         \round_in[3][1395] , \round_in[3][1394] , \round_in[3][1393] ,
         \round_in[3][1392] , \round_in[3][1391] , \round_in[3][1390] ,
         \round_in[3][1389] , \round_in[3][1388] , \round_in[3][1387] ,
         \round_in[3][1386] , \round_in[3][1385] , \round_in[3][1384] ,
         \round_in[3][1383] , \round_in[3][1382] , \round_in[3][1381] ,
         \round_in[3][1380] , \round_in[3][1379] , \round_in[3][1378] ,
         \round_in[3][1377] , \round_in[3][1376] , \round_in[3][1375] ,
         \round_in[3][1374] , \round_in[3][1373] , \round_in[3][1372] ,
         \round_in[3][1371] , \round_in[3][1370] , \round_in[3][1369] ,
         \round_in[3][1368] , \round_in[3][1367] , \round_in[3][1366] ,
         \round_in[3][1365] , \round_in[3][1364] , \round_in[3][1363] ,
         \round_in[3][1362] , \round_in[3][1361] , \round_in[3][1360] ,
         \round_in[3][1359] , \round_in[3][1358] , \round_in[3][1357] ,
         \round_in[3][1356] , \round_in[3][1355] , \round_in[3][1354] ,
         \round_in[3][1353] , \round_in[3][1352] , \round_in[3][1351] ,
         \round_in[3][1350] , \round_in[3][1349] , \round_in[3][1348] ,
         \round_in[3][1347] , \round_in[3][1346] , \round_in[3][1345] ,
         \round_in[3][1344] , \round_in[3][1343] , \round_in[3][1342] ,
         \round_in[3][1341] , \round_in[3][1340] , \round_in[3][1339] ,
         \round_in[3][1338] , \round_in[3][1337] , \round_in[3][1336] ,
         \round_in[3][1335] , \round_in[3][1334] , \round_in[3][1333] ,
         \round_in[3][1332] , \round_in[3][1331] , \round_in[3][1330] ,
         \round_in[3][1329] , \round_in[3][1328] , \round_in[3][1327] ,
         \round_in[3][1326] , \round_in[3][1325] , \round_in[3][1324] ,
         \round_in[3][1323] , \round_in[3][1322] , \round_in[3][1321] ,
         \round_in[3][1320] , \round_in[3][1319] , \round_in[3][1318] ,
         \round_in[3][1317] , \round_in[3][1316] , \round_in[3][1315] ,
         \round_in[3][1314] , \round_in[3][1313] , \round_in[3][1312] ,
         \round_in[3][1311] , \round_in[3][1310] , \round_in[3][1309] ,
         \round_in[3][1308] , \round_in[3][1307] , \round_in[3][1306] ,
         \round_in[3][1305] , \round_in[3][1304] , \round_in[3][1303] ,
         \round_in[3][1302] , \round_in[3][1301] , \round_in[3][1300] ,
         \round_in[3][1299] , \round_in[3][1298] , \round_in[3][1297] ,
         \round_in[3][1296] , \round_in[3][1295] , \round_in[3][1294] ,
         \round_in[3][1293] , \round_in[3][1292] , \round_in[3][1291] ,
         \round_in[3][1290] , \round_in[3][1289] , \round_in[3][1288] ,
         \round_in[3][1287] , \round_in[3][1286] , \round_in[3][1285] ,
         \round_in[3][1284] , \round_in[3][1283] , \round_in[3][1282] ,
         \round_in[3][1281] , \round_in[3][1280] , \round_in[3][1279] ,
         \round_in[3][1278] , \round_in[3][1277] , \round_in[3][1276] ,
         \round_in[3][1275] , \round_in[3][1274] , \round_in[3][1273] ,
         \round_in[3][1272] , \round_in[3][1271] , \round_in[3][1270] ,
         \round_in[3][1269] , \round_in[3][1268] , \round_in[3][1267] ,
         \round_in[3][1266] , \round_in[3][1265] , \round_in[3][1264] ,
         \round_in[3][1263] , \round_in[3][1262] , \round_in[3][1261] ,
         \round_in[3][1260] , \round_in[3][1259] , \round_in[3][1258] ,
         \round_in[3][1257] , \round_in[3][1256] , \round_in[3][1255] ,
         \round_in[3][1254] , \round_in[3][1253] , \round_in[3][1252] ,
         \round_in[3][1251] , \round_in[3][1250] , \round_in[3][1249] ,
         \round_in[3][1248] , \round_in[3][1247] , \round_in[3][1246] ,
         \round_in[3][1245] , \round_in[3][1244] , \round_in[3][1243] ,
         \round_in[3][1242] , \round_in[3][1241] , \round_in[3][1240] ,
         \round_in[3][1239] , \round_in[3][1238] , \round_in[3][1237] ,
         \round_in[3][1236] , \round_in[3][1235] , \round_in[3][1234] ,
         \round_in[3][1233] , \round_in[3][1232] , \round_in[3][1231] ,
         \round_in[3][1230] , \round_in[3][1229] , \round_in[3][1228] ,
         \round_in[3][1227] , \round_in[3][1226] , \round_in[3][1225] ,
         \round_in[3][1224] , \round_in[3][1223] , \round_in[3][1222] ,
         \round_in[3][1221] , \round_in[3][1220] , \round_in[3][1219] ,
         \round_in[3][1218] , \round_in[3][1217] , \round_in[3][1216] ,
         \round_in[3][1215] , \round_in[3][1214] , \round_in[3][1213] ,
         \round_in[3][1212] , \round_in[3][1211] , \round_in[3][1210] ,
         \round_in[3][1209] , \round_in[3][1208] , \round_in[3][1207] ,
         \round_in[3][1206] , \round_in[3][1205] , \round_in[3][1204] ,
         \round_in[3][1203] , \round_in[3][1202] , \round_in[3][1201] ,
         \round_in[3][1200] , \round_in[3][1199] , \round_in[3][1198] ,
         \round_in[3][1197] , \round_in[3][1196] , \round_in[3][1195] ,
         \round_in[3][1194] , \round_in[3][1193] , \round_in[3][1192] ,
         \round_in[3][1191] , \round_in[3][1190] , \round_in[3][1189] ,
         \round_in[3][1188] , \round_in[3][1187] , \round_in[3][1186] ,
         \round_in[3][1185] , \round_in[3][1184] , \round_in[3][1183] ,
         \round_in[3][1182] , \round_in[3][1181] , \round_in[3][1180] ,
         \round_in[3][1179] , \round_in[3][1178] , \round_in[3][1177] ,
         \round_in[3][1176] , \round_in[3][1175] , \round_in[3][1174] ,
         \round_in[3][1173] , \round_in[3][1172] , \round_in[3][1171] ,
         \round_in[3][1170] , \round_in[3][1169] , \round_in[3][1168] ,
         \round_in[3][1167] , \round_in[3][1166] , \round_in[3][1165] ,
         \round_in[3][1164] , \round_in[3][1163] , \round_in[3][1162] ,
         \round_in[3][1161] , \round_in[3][1160] , \round_in[3][1159] ,
         \round_in[3][1158] , \round_in[3][1157] , \round_in[3][1156] ,
         \round_in[3][1155] , \round_in[3][1154] , \round_in[3][1153] ,
         \round_in[3][1152] , \round_in[3][1151] , \round_in[3][1150] ,
         \round_in[3][1149] , \round_in[3][1148] , \round_in[3][1147] ,
         \round_in[3][1146] , \round_in[3][1145] , \round_in[3][1144] ,
         \round_in[3][1143] , \round_in[3][1142] , \round_in[3][1141] ,
         \round_in[3][1140] , \round_in[3][1139] , \round_in[3][1138] ,
         \round_in[3][1137] , \round_in[3][1136] , \round_in[3][1135] ,
         \round_in[3][1134] , \round_in[3][1133] , \round_in[3][1132] ,
         \round_in[3][1131] , \round_in[3][1130] , \round_in[3][1129] ,
         \round_in[3][1128] , \round_in[3][1127] , \round_in[3][1126] ,
         \round_in[3][1125] , \round_in[3][1124] , \round_in[3][1123] ,
         \round_in[3][1122] , \round_in[3][1121] , \round_in[3][1120] ,
         \round_in[3][1119] , \round_in[3][1118] , \round_in[3][1117] ,
         \round_in[3][1116] , \round_in[3][1115] , \round_in[3][1114] ,
         \round_in[3][1113] , \round_in[3][1112] , \round_in[3][1111] ,
         \round_in[3][1110] , \round_in[3][1109] , \round_in[3][1108] ,
         \round_in[3][1107] , \round_in[3][1106] , \round_in[3][1105] ,
         \round_in[3][1104] , \round_in[3][1103] , \round_in[3][1102] ,
         \round_in[3][1101] , \round_in[3][1100] , \round_in[3][1099] ,
         \round_in[3][1098] , \round_in[3][1097] , \round_in[3][1096] ,
         \round_in[3][1095] , \round_in[3][1094] , \round_in[3][1093] ,
         \round_in[3][1092] , \round_in[3][1091] , \round_in[3][1090] ,
         \round_in[3][1089] , \round_in[3][1088] , \round_in[3][1087] ,
         \round_in[3][1086] , \round_in[3][1085] , \round_in[3][1084] ,
         \round_in[3][1083] , \round_in[3][1082] , \round_in[3][1081] ,
         \round_in[3][1080] , \round_in[3][1079] , \round_in[3][1078] ,
         \round_in[3][1077] , \round_in[3][1076] , \round_in[3][1075] ,
         \round_in[3][1074] , \round_in[3][1073] , \round_in[3][1072] ,
         \round_in[3][1071] , \round_in[3][1070] , \round_in[3][1069] ,
         \round_in[3][1068] , \round_in[3][1067] , \round_in[3][1066] ,
         \round_in[3][1065] , \round_in[3][1064] , \round_in[3][1063] ,
         \round_in[3][1062] , \round_in[3][1061] , \round_in[3][1060] ,
         \round_in[3][1059] , \round_in[3][1058] , \round_in[3][1057] ,
         \round_in[3][1056] , \round_in[3][1055] , \round_in[3][1054] ,
         \round_in[3][1053] , \round_in[3][1052] , \round_in[3][1051] ,
         \round_in[3][1050] , \round_in[3][1049] , \round_in[3][1048] ,
         \round_in[3][1047] , \round_in[3][1046] , \round_in[3][1045] ,
         \round_in[3][1044] , \round_in[3][1043] , \round_in[3][1042] ,
         \round_in[3][1041] , \round_in[3][1040] , \round_in[3][1039] ,
         \round_in[3][1038] , \round_in[3][1037] , \round_in[3][1036] ,
         \round_in[3][1035] , \round_in[3][1034] , \round_in[3][1033] ,
         \round_in[3][1032] , \round_in[3][1031] , \round_in[3][1030] ,
         \round_in[3][1029] , \round_in[3][1028] , \round_in[3][1027] ,
         \round_in[3][1026] , \round_in[3][1025] , \round_in[3][1024] ,
         \round_in[3][1023] , \round_in[3][1022] , \round_in[3][1021] ,
         \round_in[3][1020] , \round_in[3][1019] , \round_in[3][1018] ,
         \round_in[3][1017] , \round_in[3][1016] , \round_in[3][1015] ,
         \round_in[3][1014] , \round_in[3][1013] , \round_in[3][1012] ,
         \round_in[3][1011] , \round_in[3][1010] , \round_in[3][1009] ,
         \round_in[3][1008] , \round_in[3][1007] , \round_in[3][1006] ,
         \round_in[3][1005] , \round_in[3][1004] , \round_in[3][1003] ,
         \round_in[3][1002] , \round_in[3][1001] , \round_in[3][1000] ,
         \round_in[3][999] , \round_in[3][998] , \round_in[3][997] ,
         \round_in[3][996] , \round_in[3][995] , \round_in[3][994] ,
         \round_in[3][993] , \round_in[3][992] , \round_in[3][991] ,
         \round_in[3][990] , \round_in[3][989] , \round_in[3][988] ,
         \round_in[3][987] , \round_in[3][986] , \round_in[3][985] ,
         \round_in[3][984] , \round_in[3][983] , \round_in[3][982] ,
         \round_in[3][981] , \round_in[3][980] , \round_in[3][979] ,
         \round_in[3][978] , \round_in[3][977] , \round_in[3][976] ,
         \round_in[3][975] , \round_in[3][974] , \round_in[3][973] ,
         \round_in[3][972] , \round_in[3][971] , \round_in[3][970] ,
         \round_in[3][969] , \round_in[3][968] , \round_in[3][967] ,
         \round_in[3][966] , \round_in[3][965] , \round_in[3][964] ,
         \round_in[3][963] , \round_in[3][962] , \round_in[3][961] ,
         \round_in[3][960] , \round_in[3][959] , \round_in[3][958] ,
         \round_in[3][957] , \round_in[3][956] , \round_in[3][955] ,
         \round_in[3][954] , \round_in[3][953] , \round_in[3][952] ,
         \round_in[3][951] , \round_in[3][950] , \round_in[3][949] ,
         \round_in[3][948] , \round_in[3][947] , \round_in[3][946] ,
         \round_in[3][945] , \round_in[3][944] , \round_in[3][943] ,
         \round_in[3][942] , \round_in[3][941] , \round_in[3][940] ,
         \round_in[3][939] , \round_in[3][938] , \round_in[3][937] ,
         \round_in[3][936] , \round_in[3][935] , \round_in[3][934] ,
         \round_in[3][933] , \round_in[3][932] , \round_in[3][931] ,
         \round_in[3][930] , \round_in[3][929] , \round_in[3][928] ,
         \round_in[3][927] , \round_in[3][926] , \round_in[3][925] ,
         \round_in[3][924] , \round_in[3][923] , \round_in[3][922] ,
         \round_in[3][921] , \round_in[3][920] , \round_in[3][919] ,
         \round_in[3][918] , \round_in[3][917] , \round_in[3][916] ,
         \round_in[3][915] , \round_in[3][914] , \round_in[3][913] ,
         \round_in[3][912] , \round_in[3][911] , \round_in[3][910] ,
         \round_in[3][909] , \round_in[3][908] , \round_in[3][907] ,
         \round_in[3][906] , \round_in[3][905] , \round_in[3][904] ,
         \round_in[3][903] , \round_in[3][902] , \round_in[3][901] ,
         \round_in[3][900] , \round_in[3][899] , \round_in[3][898] ,
         \round_in[3][897] , \round_in[3][896] , \round_in[3][895] ,
         \round_in[3][894] , \round_in[3][893] , \round_in[3][892] ,
         \round_in[3][891] , \round_in[3][890] , \round_in[3][889] ,
         \round_in[3][888] , \round_in[3][887] , \round_in[3][886] ,
         \round_in[3][885] , \round_in[3][884] , \round_in[3][883] ,
         \round_in[3][882] , \round_in[3][881] , \round_in[3][880] ,
         \round_in[3][879] , \round_in[3][878] , \round_in[3][877] ,
         \round_in[3][876] , \round_in[3][875] , \round_in[3][874] ,
         \round_in[3][873] , \round_in[3][872] , \round_in[3][871] ,
         \round_in[3][870] , \round_in[3][869] , \round_in[3][868] ,
         \round_in[3][867] , \round_in[3][866] , \round_in[3][865] ,
         \round_in[3][864] , \round_in[3][863] , \round_in[3][862] ,
         \round_in[3][861] , \round_in[3][860] , \round_in[3][859] ,
         \round_in[3][858] , \round_in[3][857] , \round_in[3][856] ,
         \round_in[3][855] , \round_in[3][854] , \round_in[3][853] ,
         \round_in[3][852] , \round_in[3][851] , \round_in[3][850] ,
         \round_in[3][849] , \round_in[3][848] , \round_in[3][847] ,
         \round_in[3][846] , \round_in[3][845] , \round_in[3][844] ,
         \round_in[3][843] , \round_in[3][842] , \round_in[3][841] ,
         \round_in[3][840] , \round_in[3][839] , \round_in[3][838] ,
         \round_in[3][837] , \round_in[3][836] , \round_in[3][835] ,
         \round_in[3][834] , \round_in[3][833] , \round_in[3][832] ,
         \round_in[3][831] , \round_in[3][830] , \round_in[3][829] ,
         \round_in[3][828] , \round_in[3][827] , \round_in[3][826] ,
         \round_in[3][825] , \round_in[3][824] , \round_in[3][823] ,
         \round_in[3][822] , \round_in[3][821] , \round_in[3][820] ,
         \round_in[3][819] , \round_in[3][818] , \round_in[3][817] ,
         \round_in[3][816] , \round_in[3][815] , \round_in[3][814] ,
         \round_in[3][813] , \round_in[3][812] , \round_in[3][811] ,
         \round_in[3][810] , \round_in[3][809] , \round_in[3][808] ,
         \round_in[3][807] , \round_in[3][806] , \round_in[3][805] ,
         \round_in[3][804] , \round_in[3][803] , \round_in[3][802] ,
         \round_in[3][801] , \round_in[3][800] , \round_in[3][799] ,
         \round_in[3][798] , \round_in[3][797] , \round_in[3][796] ,
         \round_in[3][795] , \round_in[3][794] , \round_in[3][793] ,
         \round_in[3][792] , \round_in[3][791] , \round_in[3][790] ,
         \round_in[3][789] , \round_in[3][788] , \round_in[3][787] ,
         \round_in[3][786] , \round_in[3][785] , \round_in[3][784] ,
         \round_in[3][783] , \round_in[3][782] , \round_in[3][781] ,
         \round_in[3][780] , \round_in[3][779] , \round_in[3][778] ,
         \round_in[3][777] , \round_in[3][776] , \round_in[3][775] ,
         \round_in[3][774] , \round_in[3][773] , \round_in[3][772] ,
         \round_in[3][771] , \round_in[3][770] , \round_in[3][769] ,
         \round_in[3][768] , \round_in[3][767] , \round_in[3][766] ,
         \round_in[3][765] , \round_in[3][764] , \round_in[3][763] ,
         \round_in[3][762] , \round_in[3][761] , \round_in[3][760] ,
         \round_in[3][759] , \round_in[3][758] , \round_in[3][757] ,
         \round_in[3][756] , \round_in[3][755] , \round_in[3][754] ,
         \round_in[3][753] , \round_in[3][752] , \round_in[3][751] ,
         \round_in[3][750] , \round_in[3][749] , \round_in[3][748] ,
         \round_in[3][747] , \round_in[3][746] , \round_in[3][745] ,
         \round_in[3][744] , \round_in[3][743] , \round_in[3][742] ,
         \round_in[3][741] , \round_in[3][740] , \round_in[3][739] ,
         \round_in[3][738] , \round_in[3][737] , \round_in[3][736] ,
         \round_in[3][735] , \round_in[3][734] , \round_in[3][733] ,
         \round_in[3][732] , \round_in[3][731] , \round_in[3][730] ,
         \round_in[3][729] , \round_in[3][728] , \round_in[3][727] ,
         \round_in[3][726] , \round_in[3][725] , \round_in[3][724] ,
         \round_in[3][723] , \round_in[3][722] , \round_in[3][721] ,
         \round_in[3][720] , \round_in[3][719] , \round_in[3][718] ,
         \round_in[3][717] , \round_in[3][716] , \round_in[3][715] ,
         \round_in[3][714] , \round_in[3][713] , \round_in[3][712] ,
         \round_in[3][711] , \round_in[3][710] , \round_in[3][709] ,
         \round_in[3][708] , \round_in[3][707] , \round_in[3][706] ,
         \round_in[3][705] , \round_in[3][704] , \round_in[3][703] ,
         \round_in[3][702] , \round_in[3][701] , \round_in[3][700] ,
         \round_in[3][699] , \round_in[3][698] , \round_in[3][697] ,
         \round_in[3][696] , \round_in[3][695] , \round_in[3][694] ,
         \round_in[3][693] , \round_in[3][692] , \round_in[3][691] ,
         \round_in[3][690] , \round_in[3][689] , \round_in[3][688] ,
         \round_in[3][687] , \round_in[3][686] , \round_in[3][685] ,
         \round_in[3][684] , \round_in[3][683] , \round_in[3][682] ,
         \round_in[3][681] , \round_in[3][680] , \round_in[3][679] ,
         \round_in[3][678] , \round_in[3][677] , \round_in[3][676] ,
         \round_in[3][675] , \round_in[3][674] , \round_in[3][673] ,
         \round_in[3][672] , \round_in[3][671] , \round_in[3][670] ,
         \round_in[3][669] , \round_in[3][668] , \round_in[3][667] ,
         \round_in[3][666] , \round_in[3][665] , \round_in[3][664] ,
         \round_in[3][663] , \round_in[3][662] , \round_in[3][661] ,
         \round_in[3][660] , \round_in[3][659] , \round_in[3][658] ,
         \round_in[3][657] , \round_in[3][656] , \round_in[3][655] ,
         \round_in[3][654] , \round_in[3][653] , \round_in[3][652] ,
         \round_in[3][651] , \round_in[3][650] , \round_in[3][649] ,
         \round_in[3][648] , \round_in[3][647] , \round_in[3][646] ,
         \round_in[3][645] , \round_in[3][644] , \round_in[3][643] ,
         \round_in[3][642] , \round_in[3][641] , \round_in[3][640] ,
         \round_in[3][639] , \round_in[3][638] , \round_in[3][637] ,
         \round_in[3][636] , \round_in[3][635] , \round_in[3][634] ,
         \round_in[3][633] , \round_in[3][632] , \round_in[3][631] ,
         \round_in[3][630] , \round_in[3][629] , \round_in[3][628] ,
         \round_in[3][627] , \round_in[3][626] , \round_in[3][625] ,
         \round_in[3][624] , \round_in[3][623] , \round_in[3][622] ,
         \round_in[3][621] , \round_in[3][620] , \round_in[3][619] ,
         \round_in[3][618] , \round_in[3][617] , \round_in[3][616] ,
         \round_in[3][615] , \round_in[3][614] , \round_in[3][613] ,
         \round_in[3][612] , \round_in[3][611] , \round_in[3][610] ,
         \round_in[3][609] , \round_in[3][608] , \round_in[3][607] ,
         \round_in[3][606] , \round_in[3][605] , \round_in[3][604] ,
         \round_in[3][603] , \round_in[3][602] , \round_in[3][601] ,
         \round_in[3][600] , \round_in[3][599] , \round_in[3][598] ,
         \round_in[3][597] , \round_in[3][596] , \round_in[3][595] ,
         \round_in[3][594] , \round_in[3][593] , \round_in[3][592] ,
         \round_in[3][591] , \round_in[3][590] , \round_in[3][589] ,
         \round_in[3][588] , \round_in[3][587] , \round_in[3][586] ,
         \round_in[3][585] , \round_in[3][584] , \round_in[3][583] ,
         \round_in[3][582] , \round_in[3][581] , \round_in[3][580] ,
         \round_in[3][579] , \round_in[3][578] , \round_in[3][577] ,
         \round_in[3][576] , \round_in[3][575] , \round_in[3][574] ,
         \round_in[3][573] , \round_in[3][572] , \round_in[3][571] ,
         \round_in[3][570] , \round_in[3][569] , \round_in[3][568] ,
         \round_in[3][567] , \round_in[3][566] , \round_in[3][565] ,
         \round_in[3][564] , \round_in[3][563] , \round_in[3][562] ,
         \round_in[3][561] , \round_in[3][560] , \round_in[3][559] ,
         \round_in[3][558] , \round_in[3][557] , \round_in[3][556] ,
         \round_in[3][555] , \round_in[3][554] , \round_in[3][553] ,
         \round_in[3][552] , \round_in[3][551] , \round_in[3][550] ,
         \round_in[3][549] , \round_in[3][548] , \round_in[3][547] ,
         \round_in[3][546] , \round_in[3][545] , \round_in[3][544] ,
         \round_in[3][543] , \round_in[3][542] , \round_in[3][541] ,
         \round_in[3][540] , \round_in[3][539] , \round_in[3][538] ,
         \round_in[3][537] , \round_in[3][536] , \round_in[3][535] ,
         \round_in[3][534] , \round_in[3][533] , \round_in[3][532] ,
         \round_in[3][531] , \round_in[3][530] , \round_in[3][529] ,
         \round_in[3][528] , \round_in[3][527] , \round_in[3][526] ,
         \round_in[3][525] , \round_in[3][524] , \round_in[3][523] ,
         \round_in[3][522] , \round_in[3][521] , \round_in[3][520] ,
         \round_in[3][519] , \round_in[3][518] , \round_in[3][517] ,
         \round_in[3][516] , \round_in[3][515] , \round_in[3][514] ,
         \round_in[3][513] , \round_in[3][512] , \round_in[3][511] ,
         \round_in[3][510] , \round_in[3][509] , \round_in[3][508] ,
         \round_in[3][507] , \round_in[3][506] , \round_in[3][505] ,
         \round_in[3][504] , \round_in[3][503] , \round_in[3][502] ,
         \round_in[3][501] , \round_in[3][500] , \round_in[3][499] ,
         \round_in[3][498] , \round_in[3][497] , \round_in[3][496] ,
         \round_in[3][495] , \round_in[3][494] , \round_in[3][493] ,
         \round_in[3][492] , \round_in[3][491] , \round_in[3][490] ,
         \round_in[3][489] , \round_in[3][488] , \round_in[3][487] ,
         \round_in[3][486] , \round_in[3][485] , \round_in[3][484] ,
         \round_in[3][483] , \round_in[3][482] , \round_in[3][481] ,
         \round_in[3][480] , \round_in[3][479] , \round_in[3][478] ,
         \round_in[3][477] , \round_in[3][476] , \round_in[3][475] ,
         \round_in[3][474] , \round_in[3][473] , \round_in[3][472] ,
         \round_in[3][471] , \round_in[3][470] , \round_in[3][469] ,
         \round_in[3][468] , \round_in[3][467] , \round_in[3][466] ,
         \round_in[3][465] , \round_in[3][464] , \round_in[3][463] ,
         \round_in[3][462] , \round_in[3][461] , \round_in[3][460] ,
         \round_in[3][459] , \round_in[3][458] , \round_in[3][457] ,
         \round_in[3][456] , \round_in[3][455] , \round_in[3][454] ,
         \round_in[3][453] , \round_in[3][452] , \round_in[3][451] ,
         \round_in[3][450] , \round_in[3][449] , \round_in[3][448] ,
         \round_in[3][447] , \round_in[3][446] , \round_in[3][445] ,
         \round_in[3][444] , \round_in[3][443] , \round_in[3][442] ,
         \round_in[3][441] , \round_in[3][440] , \round_in[3][439] ,
         \round_in[3][438] , \round_in[3][437] , \round_in[3][436] ,
         \round_in[3][435] , \round_in[3][434] , \round_in[3][433] ,
         \round_in[3][432] , \round_in[3][431] , \round_in[3][430] ,
         \round_in[3][429] , \round_in[3][428] , \round_in[3][427] ,
         \round_in[3][426] , \round_in[3][425] , \round_in[3][424] ,
         \round_in[3][423] , \round_in[3][422] , \round_in[3][421] ,
         \round_in[3][420] , \round_in[3][419] , \round_in[3][418] ,
         \round_in[3][417] , \round_in[3][416] , \round_in[3][415] ,
         \round_in[3][414] , \round_in[3][413] , \round_in[3][412] ,
         \round_in[3][411] , \round_in[3][410] , \round_in[3][409] ,
         \round_in[3][408] , \round_in[3][407] , \round_in[3][406] ,
         \round_in[3][405] , \round_in[3][404] , \round_in[3][403] ,
         \round_in[3][402] , \round_in[3][401] , \round_in[3][400] ,
         \round_in[3][399] , \round_in[3][398] , \round_in[3][397] ,
         \round_in[3][396] , \round_in[3][395] , \round_in[3][394] ,
         \round_in[3][393] , \round_in[3][392] , \round_in[3][391] ,
         \round_in[3][390] , \round_in[3][389] , \round_in[3][388] ,
         \round_in[3][387] , \round_in[3][386] , \round_in[3][385] ,
         \round_in[3][384] , \round_in[3][383] , \round_in[3][382] ,
         \round_in[3][381] , \round_in[3][380] , \round_in[3][379] ,
         \round_in[3][378] , \round_in[3][377] , \round_in[3][376] ,
         \round_in[3][375] , \round_in[3][374] , \round_in[3][373] ,
         \round_in[3][372] , \round_in[3][371] , \round_in[3][370] ,
         \round_in[3][369] , \round_in[3][368] , \round_in[3][367] ,
         \round_in[3][366] , \round_in[3][365] , \round_in[3][364] ,
         \round_in[3][363] , \round_in[3][362] , \round_in[3][361] ,
         \round_in[3][360] , \round_in[3][359] , \round_in[3][358] ,
         \round_in[3][357] , \round_in[3][356] , \round_in[3][355] ,
         \round_in[3][354] , \round_in[3][353] , \round_in[3][352] ,
         \round_in[3][351] , \round_in[3][350] , \round_in[3][349] ,
         \round_in[3][348] , \round_in[3][347] , \round_in[3][346] ,
         \round_in[3][345] , \round_in[3][344] , \round_in[3][343] ,
         \round_in[3][342] , \round_in[3][341] , \round_in[3][340] ,
         \round_in[3][339] , \round_in[3][338] , \round_in[3][337] ,
         \round_in[3][336] , \round_in[3][335] , \round_in[3][334] ,
         \round_in[3][333] , \round_in[3][332] , \round_in[3][331] ,
         \round_in[3][330] , \round_in[3][329] , \round_in[3][328] ,
         \round_in[3][327] , \round_in[3][326] , \round_in[3][325] ,
         \round_in[3][324] , \round_in[3][323] , \round_in[3][322] ,
         \round_in[3][321] , \round_in[3][320] , \round_in[3][319] ,
         \round_in[3][318] , \round_in[3][317] , \round_in[3][316] ,
         \round_in[3][315] , \round_in[3][314] , \round_in[3][313] ,
         \round_in[3][312] , \round_in[3][311] , \round_in[3][310] ,
         \round_in[3][309] , \round_in[3][308] , \round_in[3][307] ,
         \round_in[3][306] , \round_in[3][305] , \round_in[3][304] ,
         \round_in[3][303] , \round_in[3][302] , \round_in[3][301] ,
         \round_in[3][300] , \round_in[3][299] , \round_in[3][298] ,
         \round_in[3][297] , \round_in[3][296] , \round_in[3][295] ,
         \round_in[3][294] , \round_in[3][293] , \round_in[3][292] ,
         \round_in[3][291] , \round_in[3][290] , \round_in[3][289] ,
         \round_in[3][288] , \round_in[3][287] , \round_in[3][286] ,
         \round_in[3][285] , \round_in[3][284] , \round_in[3][283] ,
         \round_in[3][282] , \round_in[3][281] , \round_in[3][280] ,
         \round_in[3][279] , \round_in[3][278] , \round_in[3][277] ,
         \round_in[3][276] , \round_in[3][275] , \round_in[3][274] ,
         \round_in[3][273] , \round_in[3][272] , \round_in[3][271] ,
         \round_in[3][270] , \round_in[3][269] , \round_in[3][268] ,
         \round_in[3][267] , \round_in[3][266] , \round_in[3][265] ,
         \round_in[3][264] , \round_in[3][263] , \round_in[3][262] ,
         \round_in[3][261] , \round_in[3][260] , \round_in[3][259] ,
         \round_in[3][258] , \round_in[3][257] , \round_in[3][256] ,
         \round_in[3][255] , \round_in[3][254] , \round_in[3][253] ,
         \round_in[3][252] , \round_in[3][251] , \round_in[3][250] ,
         \round_in[3][249] , \round_in[3][248] , \round_in[3][247] ,
         \round_in[3][246] , \round_in[3][245] , \round_in[3][244] ,
         \round_in[3][243] , \round_in[3][242] , \round_in[3][241] ,
         \round_in[3][240] , \round_in[3][239] , \round_in[3][238] ,
         \round_in[3][237] , \round_in[3][236] , \round_in[3][235] ,
         \round_in[3][234] , \round_in[3][233] , \round_in[3][232] ,
         \round_in[3][231] , \round_in[3][230] , \round_in[3][229] ,
         \round_in[3][228] , \round_in[3][227] , \round_in[3][226] ,
         \round_in[3][225] , \round_in[3][224] , \round_in[3][223] ,
         \round_in[3][222] , \round_in[3][221] , \round_in[3][220] ,
         \round_in[3][219] , \round_in[3][218] , \round_in[3][217] ,
         \round_in[3][216] , \round_in[3][215] , \round_in[3][214] ,
         \round_in[3][213] , \round_in[3][212] , \round_in[3][211] ,
         \round_in[3][210] , \round_in[3][209] , \round_in[3][208] ,
         \round_in[3][207] , \round_in[3][206] , \round_in[3][205] ,
         \round_in[3][204] , \round_in[3][203] , \round_in[3][202] ,
         \round_in[3][201] , \round_in[3][200] , \round_in[3][199] ,
         \round_in[3][198] , \round_in[3][197] , \round_in[3][196] ,
         \round_in[3][195] , \round_in[3][194] , \round_in[3][193] ,
         \round_in[3][192] , \round_in[3][191] , \round_in[3][190] ,
         \round_in[3][189] , \round_in[3][188] , \round_in[3][187] ,
         \round_in[3][186] , \round_in[3][185] , \round_in[3][184] ,
         \round_in[3][183] , \round_in[3][182] , \round_in[3][181] ,
         \round_in[3][180] , \round_in[3][179] , \round_in[3][178] ,
         \round_in[3][177] , \round_in[3][176] , \round_in[3][175] ,
         \round_in[3][174] , \round_in[3][173] , \round_in[3][172] ,
         \round_in[3][171] , \round_in[3][170] , \round_in[3][169] ,
         \round_in[3][168] , \round_in[3][167] , \round_in[3][166] ,
         \round_in[3][165] , \round_in[3][164] , \round_in[3][163] ,
         \round_in[3][162] , \round_in[3][161] , \round_in[3][160] ,
         \round_in[3][159] , \round_in[3][158] , \round_in[3][157] ,
         \round_in[3][156] , \round_in[3][155] , \round_in[3][154] ,
         \round_in[3][153] , \round_in[3][152] , \round_in[3][151] ,
         \round_in[3][150] , \round_in[3][149] , \round_in[3][148] ,
         \round_in[3][147] , \round_in[3][146] , \round_in[3][145] ,
         \round_in[3][144] , \round_in[3][143] , \round_in[3][142] ,
         \round_in[3][141] , \round_in[3][140] , \round_in[3][139] ,
         \round_in[3][138] , \round_in[3][137] , \round_in[3][136] ,
         \round_in[3][135] , \round_in[3][134] , \round_in[3][133] ,
         \round_in[3][132] , \round_in[3][131] , \round_in[3][130] ,
         \round_in[3][129] , \round_in[3][128] , \round_in[3][127] ,
         \round_in[3][126] , \round_in[3][125] , \round_in[3][124] ,
         \round_in[3][123] , \round_in[3][122] , \round_in[3][121] ,
         \round_in[3][120] , \round_in[3][119] , \round_in[3][118] ,
         \round_in[3][117] , \round_in[3][116] , \round_in[3][115] ,
         \round_in[3][114] , \round_in[3][113] , \round_in[3][112] ,
         \round_in[3][111] , \round_in[3][110] , \round_in[3][109] ,
         \round_in[3][108] , \round_in[3][107] , \round_in[3][106] ,
         \round_in[3][105] , \round_in[3][104] , \round_in[3][103] ,
         \round_in[3][102] , \round_in[3][101] , \round_in[3][100] ,
         \round_in[3][99] , \round_in[3][98] , \round_in[3][97] ,
         \round_in[3][96] , \round_in[3][95] , \round_in[3][94] ,
         \round_in[3][93] , \round_in[3][92] , \round_in[3][91] ,
         \round_in[3][90] , \round_in[3][89] , \round_in[3][88] ,
         \round_in[3][87] , \round_in[3][86] , \round_in[3][85] ,
         \round_in[3][84] , \round_in[3][83] , \round_in[3][82] ,
         \round_in[3][81] , \round_in[3][80] , \round_in[3][79] ,
         \round_in[3][78] , \round_in[3][77] , \round_in[3][76] ,
         \round_in[3][75] , \round_in[3][74] , \round_in[3][73] ,
         \round_in[3][72] , \round_in[3][71] , \round_in[3][70] ,
         \round_in[3][69] , \round_in[3][68] , \round_in[3][67] ,
         \round_in[3][66] , \round_in[3][65] , \round_in[3][64] ,
         \round_in[3][63] , \round_in[3][62] , \round_in[3][61] ,
         \round_in[3][60] , \round_in[3][59] , \round_in[3][58] ,
         \round_in[3][57] , \round_in[3][56] , \round_in[3][55] ,
         \round_in[3][54] , \round_in[3][53] , \round_in[3][52] ,
         \round_in[3][51] , \round_in[3][50] , \round_in[3][49] ,
         \round_in[3][48] , \round_in[3][47] , \round_in[3][46] ,
         \round_in[3][45] , \round_in[3][44] , \round_in[3][43] ,
         \round_in[3][42] , \round_in[3][41] , \round_in[3][40] ,
         \round_in[3][39] , \round_in[3][38] , \round_in[3][37] ,
         \round_in[3][36] , \round_in[3][35] , \round_in[3][34] ,
         \round_in[3][33] , \round_in[3][32] , \round_in[3][31] ,
         \round_in[3][30] , \round_in[3][29] , \round_in[3][28] ,
         \round_in[3][27] , \round_in[3][26] , \round_in[3][25] ,
         \round_in[3][24] , \round_in[3][23] , \round_in[3][22] ,
         \round_in[3][21] , \round_in[3][20] , \round_in[3][19] ,
         \round_in[3][18] , \round_in[3][17] , \round_in[3][16] ,
         \round_in[3][15] , \round_in[3][14] , \round_in[3][13] ,
         \round_in[3][12] , \round_in[3][11] , \round_in[3][10] ,
         \round_in[3][9] , \round_in[3][8] , \round_in[3][7] ,
         \round_in[3][6] , \round_in[3][5] , \round_in[3][4] ,
         \round_in[3][3] , \round_in[3][2] , \round_in[3][1] ,
         \round_in[3][0] , \round_in[2][1599] , \round_in[2][1598] ,
         \round_in[2][1597] , \round_in[2][1596] , \round_in[2][1595] ,
         \round_in[2][1594] , \round_in[2][1593] , \round_in[2][1592] ,
         \round_in[2][1591] , \round_in[2][1590] , \round_in[2][1589] ,
         \round_in[2][1588] , \round_in[2][1587] , \round_in[2][1586] ,
         \round_in[2][1585] , \round_in[2][1584] , \round_in[2][1583] ,
         \round_in[2][1582] , \round_in[2][1581] , \round_in[2][1580] ,
         \round_in[2][1579] , \round_in[2][1578] , \round_in[2][1577] ,
         \round_in[2][1576] , \round_in[2][1575] , \round_in[2][1574] ,
         \round_in[2][1573] , \round_in[2][1572] , \round_in[2][1571] ,
         \round_in[2][1570] , \round_in[2][1569] , \round_in[2][1568] ,
         \round_in[2][1567] , \round_in[2][1566] , \round_in[2][1565] ,
         \round_in[2][1564] , \round_in[2][1563] , \round_in[2][1562] ,
         \round_in[2][1561] , \round_in[2][1560] , \round_in[2][1559] ,
         \round_in[2][1558] , \round_in[2][1557] , \round_in[2][1556] ,
         \round_in[2][1555] , \round_in[2][1554] , \round_in[2][1553] ,
         \round_in[2][1552] , \round_in[2][1551] , \round_in[2][1550] ,
         \round_in[2][1549] , \round_in[2][1548] , \round_in[2][1547] ,
         \round_in[2][1546] , \round_in[2][1545] , \round_in[2][1544] ,
         \round_in[2][1543] , \round_in[2][1542] , \round_in[2][1541] ,
         \round_in[2][1540] , \round_in[2][1539] , \round_in[2][1538] ,
         \round_in[2][1537] , \round_in[2][1536] , \round_in[2][1535] ,
         \round_in[2][1534] , \round_in[2][1533] , \round_in[2][1532] ,
         \round_in[2][1531] , \round_in[2][1530] , \round_in[2][1529] ,
         \round_in[2][1528] , \round_in[2][1527] , \round_in[2][1526] ,
         \round_in[2][1525] , \round_in[2][1524] , \round_in[2][1523] ,
         \round_in[2][1522] , \round_in[2][1521] , \round_in[2][1520] ,
         \round_in[2][1519] , \round_in[2][1518] , \round_in[2][1517] ,
         \round_in[2][1516] , \round_in[2][1515] , \round_in[2][1514] ,
         \round_in[2][1513] , \round_in[2][1512] , \round_in[2][1511] ,
         \round_in[2][1510] , \round_in[2][1509] , \round_in[2][1508] ,
         \round_in[2][1507] , \round_in[2][1506] , \round_in[2][1505] ,
         \round_in[2][1504] , \round_in[2][1503] , \round_in[2][1502] ,
         \round_in[2][1501] , \round_in[2][1500] , \round_in[2][1499] ,
         \round_in[2][1498] , \round_in[2][1497] , \round_in[2][1496] ,
         \round_in[2][1495] , \round_in[2][1494] , \round_in[2][1493] ,
         \round_in[2][1492] , \round_in[2][1491] , \round_in[2][1490] ,
         \round_in[2][1489] , \round_in[2][1488] , \round_in[2][1487] ,
         \round_in[2][1486] , \round_in[2][1485] , \round_in[2][1484] ,
         \round_in[2][1483] , \round_in[2][1482] , \round_in[2][1481] ,
         \round_in[2][1480] , \round_in[2][1479] , \round_in[2][1478] ,
         \round_in[2][1477] , \round_in[2][1476] , \round_in[2][1475] ,
         \round_in[2][1474] , \round_in[2][1473] , \round_in[2][1472] ,
         \round_in[2][1471] , \round_in[2][1470] , \round_in[2][1469] ,
         \round_in[2][1468] , \round_in[2][1467] , \round_in[2][1466] ,
         \round_in[2][1465] , \round_in[2][1464] , \round_in[2][1463] ,
         \round_in[2][1462] , \round_in[2][1461] , \round_in[2][1460] ,
         \round_in[2][1459] , \round_in[2][1458] , \round_in[2][1457] ,
         \round_in[2][1456] , \round_in[2][1455] , \round_in[2][1454] ,
         \round_in[2][1453] , \round_in[2][1452] , \round_in[2][1451] ,
         \round_in[2][1450] , \round_in[2][1449] , \round_in[2][1448] ,
         \round_in[2][1447] , \round_in[2][1446] , \round_in[2][1445] ,
         \round_in[2][1444] , \round_in[2][1443] , \round_in[2][1442] ,
         \round_in[2][1441] , \round_in[2][1440] , \round_in[2][1439] ,
         \round_in[2][1438] , \round_in[2][1437] , \round_in[2][1436] ,
         \round_in[2][1435] , \round_in[2][1434] , \round_in[2][1433] ,
         \round_in[2][1432] , \round_in[2][1431] , \round_in[2][1430] ,
         \round_in[2][1429] , \round_in[2][1428] , \round_in[2][1427] ,
         \round_in[2][1426] , \round_in[2][1425] , \round_in[2][1424] ,
         \round_in[2][1423] , \round_in[2][1422] , \round_in[2][1421] ,
         \round_in[2][1420] , \round_in[2][1419] , \round_in[2][1418] ,
         \round_in[2][1417] , \round_in[2][1416] , \round_in[2][1415] ,
         \round_in[2][1414] , \round_in[2][1413] , \round_in[2][1412] ,
         \round_in[2][1411] , \round_in[2][1410] , \round_in[2][1409] ,
         \round_in[2][1408] , \round_in[2][1407] , \round_in[2][1406] ,
         \round_in[2][1405] , \round_in[2][1404] , \round_in[2][1403] ,
         \round_in[2][1402] , \round_in[2][1401] , \round_in[2][1400] ,
         \round_in[2][1399] , \round_in[2][1398] , \round_in[2][1397] ,
         \round_in[2][1396] , \round_in[2][1395] , \round_in[2][1394] ,
         \round_in[2][1393] , \round_in[2][1392] , \round_in[2][1391] ,
         \round_in[2][1390] , \round_in[2][1389] , \round_in[2][1388] ,
         \round_in[2][1387] , \round_in[2][1386] , \round_in[2][1385] ,
         \round_in[2][1384] , \round_in[2][1383] , \round_in[2][1382] ,
         \round_in[2][1381] , \round_in[2][1380] , \round_in[2][1379] ,
         \round_in[2][1378] , \round_in[2][1377] , \round_in[2][1376] ,
         \round_in[2][1375] , \round_in[2][1374] , \round_in[2][1373] ,
         \round_in[2][1372] , \round_in[2][1371] , \round_in[2][1370] ,
         \round_in[2][1369] , \round_in[2][1368] , \round_in[2][1367] ,
         \round_in[2][1366] , \round_in[2][1365] , \round_in[2][1364] ,
         \round_in[2][1363] , \round_in[2][1362] , \round_in[2][1361] ,
         \round_in[2][1360] , \round_in[2][1359] , \round_in[2][1358] ,
         \round_in[2][1357] , \round_in[2][1356] , \round_in[2][1355] ,
         \round_in[2][1354] , \round_in[2][1353] , \round_in[2][1352] ,
         \round_in[2][1351] , \round_in[2][1350] , \round_in[2][1349] ,
         \round_in[2][1348] , \round_in[2][1347] , \round_in[2][1346] ,
         \round_in[2][1345] , \round_in[2][1344] , \round_in[2][1343] ,
         \round_in[2][1342] , \round_in[2][1341] , \round_in[2][1340] ,
         \round_in[2][1339] , \round_in[2][1338] , \round_in[2][1337] ,
         \round_in[2][1336] , \round_in[2][1335] , \round_in[2][1334] ,
         \round_in[2][1333] , \round_in[2][1332] , \round_in[2][1331] ,
         \round_in[2][1330] , \round_in[2][1329] , \round_in[2][1328] ,
         \round_in[2][1327] , \round_in[2][1326] , \round_in[2][1325] ,
         \round_in[2][1324] , \round_in[2][1323] , \round_in[2][1322] ,
         \round_in[2][1321] , \round_in[2][1320] , \round_in[2][1319] ,
         \round_in[2][1318] , \round_in[2][1317] , \round_in[2][1316] ,
         \round_in[2][1315] , \round_in[2][1314] , \round_in[2][1313] ,
         \round_in[2][1312] , \round_in[2][1311] , \round_in[2][1310] ,
         \round_in[2][1309] , \round_in[2][1308] , \round_in[2][1307] ,
         \round_in[2][1306] , \round_in[2][1305] , \round_in[2][1304] ,
         \round_in[2][1303] , \round_in[2][1302] , \round_in[2][1301] ,
         \round_in[2][1300] , \round_in[2][1299] , \round_in[2][1298] ,
         \round_in[2][1297] , \round_in[2][1296] , \round_in[2][1295] ,
         \round_in[2][1294] , \round_in[2][1293] , \round_in[2][1292] ,
         \round_in[2][1291] , \round_in[2][1290] , \round_in[2][1289] ,
         \round_in[2][1288] , \round_in[2][1287] , \round_in[2][1286] ,
         \round_in[2][1285] , \round_in[2][1284] , \round_in[2][1283] ,
         \round_in[2][1282] , \round_in[2][1281] , \round_in[2][1280] ,
         \round_in[2][1279] , \round_in[2][1278] , \round_in[2][1277] ,
         \round_in[2][1276] , \round_in[2][1275] , \round_in[2][1274] ,
         \round_in[2][1273] , \round_in[2][1272] , \round_in[2][1271] ,
         \round_in[2][1270] , \round_in[2][1269] , \round_in[2][1268] ,
         \round_in[2][1267] , \round_in[2][1266] , \round_in[2][1265] ,
         \round_in[2][1264] , \round_in[2][1263] , \round_in[2][1262] ,
         \round_in[2][1261] , \round_in[2][1260] , \round_in[2][1259] ,
         \round_in[2][1258] , \round_in[2][1257] , \round_in[2][1256] ,
         \round_in[2][1255] , \round_in[2][1254] , \round_in[2][1253] ,
         \round_in[2][1252] , \round_in[2][1251] , \round_in[2][1250] ,
         \round_in[2][1249] , \round_in[2][1248] , \round_in[2][1247] ,
         \round_in[2][1246] , \round_in[2][1245] , \round_in[2][1244] ,
         \round_in[2][1243] , \round_in[2][1242] , \round_in[2][1241] ,
         \round_in[2][1240] , \round_in[2][1239] , \round_in[2][1238] ,
         \round_in[2][1237] , \round_in[2][1236] , \round_in[2][1235] ,
         \round_in[2][1234] , \round_in[2][1233] , \round_in[2][1232] ,
         \round_in[2][1231] , \round_in[2][1230] , \round_in[2][1229] ,
         \round_in[2][1228] , \round_in[2][1227] , \round_in[2][1226] ,
         \round_in[2][1225] , \round_in[2][1224] , \round_in[2][1223] ,
         \round_in[2][1222] , \round_in[2][1221] , \round_in[2][1220] ,
         \round_in[2][1219] , \round_in[2][1218] , \round_in[2][1217] ,
         \round_in[2][1216] , \round_in[2][1215] , \round_in[2][1214] ,
         \round_in[2][1213] , \round_in[2][1212] , \round_in[2][1211] ,
         \round_in[2][1210] , \round_in[2][1209] , \round_in[2][1208] ,
         \round_in[2][1207] , \round_in[2][1206] , \round_in[2][1205] ,
         \round_in[2][1204] , \round_in[2][1203] , \round_in[2][1202] ,
         \round_in[2][1201] , \round_in[2][1200] , \round_in[2][1199] ,
         \round_in[2][1198] , \round_in[2][1197] , \round_in[2][1196] ,
         \round_in[2][1195] , \round_in[2][1194] , \round_in[2][1193] ,
         \round_in[2][1192] , \round_in[2][1191] , \round_in[2][1190] ,
         \round_in[2][1189] , \round_in[2][1188] , \round_in[2][1187] ,
         \round_in[2][1186] , \round_in[2][1185] , \round_in[2][1184] ,
         \round_in[2][1183] , \round_in[2][1182] , \round_in[2][1181] ,
         \round_in[2][1180] , \round_in[2][1179] , \round_in[2][1178] ,
         \round_in[2][1177] , \round_in[2][1176] , \round_in[2][1175] ,
         \round_in[2][1174] , \round_in[2][1173] , \round_in[2][1172] ,
         \round_in[2][1171] , \round_in[2][1170] , \round_in[2][1169] ,
         \round_in[2][1168] , \round_in[2][1167] , \round_in[2][1166] ,
         \round_in[2][1165] , \round_in[2][1164] , \round_in[2][1163] ,
         \round_in[2][1162] , \round_in[2][1161] , \round_in[2][1160] ,
         \round_in[2][1159] , \round_in[2][1158] , \round_in[2][1157] ,
         \round_in[2][1156] , \round_in[2][1155] , \round_in[2][1154] ,
         \round_in[2][1153] , \round_in[2][1152] , \round_in[2][1151] ,
         \round_in[2][1150] , \round_in[2][1149] , \round_in[2][1148] ,
         \round_in[2][1147] , \round_in[2][1146] , \round_in[2][1145] ,
         \round_in[2][1144] , \round_in[2][1143] , \round_in[2][1142] ,
         \round_in[2][1141] , \round_in[2][1140] , \round_in[2][1139] ,
         \round_in[2][1138] , \round_in[2][1137] , \round_in[2][1136] ,
         \round_in[2][1135] , \round_in[2][1134] , \round_in[2][1133] ,
         \round_in[2][1132] , \round_in[2][1131] , \round_in[2][1130] ,
         \round_in[2][1129] , \round_in[2][1128] , \round_in[2][1127] ,
         \round_in[2][1126] , \round_in[2][1125] , \round_in[2][1124] ,
         \round_in[2][1123] , \round_in[2][1122] , \round_in[2][1121] ,
         \round_in[2][1120] , \round_in[2][1119] , \round_in[2][1118] ,
         \round_in[2][1117] , \round_in[2][1116] , \round_in[2][1115] ,
         \round_in[2][1114] , \round_in[2][1113] , \round_in[2][1112] ,
         \round_in[2][1111] , \round_in[2][1110] , \round_in[2][1109] ,
         \round_in[2][1108] , \round_in[2][1107] , \round_in[2][1106] ,
         \round_in[2][1105] , \round_in[2][1104] , \round_in[2][1103] ,
         \round_in[2][1102] , \round_in[2][1101] , \round_in[2][1100] ,
         \round_in[2][1099] , \round_in[2][1098] , \round_in[2][1097] ,
         \round_in[2][1096] , \round_in[2][1095] , \round_in[2][1094] ,
         \round_in[2][1093] , \round_in[2][1092] , \round_in[2][1091] ,
         \round_in[2][1090] , \round_in[2][1089] , \round_in[2][1088] ,
         \round_in[2][1087] , \round_in[2][1086] , \round_in[2][1085] ,
         \round_in[2][1084] , \round_in[2][1083] , \round_in[2][1082] ,
         \round_in[2][1081] , \round_in[2][1080] , \round_in[2][1079] ,
         \round_in[2][1078] , \round_in[2][1077] , \round_in[2][1076] ,
         \round_in[2][1075] , \round_in[2][1074] , \round_in[2][1073] ,
         \round_in[2][1072] , \round_in[2][1071] , \round_in[2][1070] ,
         \round_in[2][1069] , \round_in[2][1068] , \round_in[2][1067] ,
         \round_in[2][1066] , \round_in[2][1065] , \round_in[2][1064] ,
         \round_in[2][1063] , \round_in[2][1062] , \round_in[2][1061] ,
         \round_in[2][1060] , \round_in[2][1059] , \round_in[2][1058] ,
         \round_in[2][1057] , \round_in[2][1056] , \round_in[2][1055] ,
         \round_in[2][1054] , \round_in[2][1053] , \round_in[2][1052] ,
         \round_in[2][1051] , \round_in[2][1050] , \round_in[2][1049] ,
         \round_in[2][1048] , \round_in[2][1047] , \round_in[2][1046] ,
         \round_in[2][1045] , \round_in[2][1044] , \round_in[2][1043] ,
         \round_in[2][1042] , \round_in[2][1041] , \round_in[2][1040] ,
         \round_in[2][1039] , \round_in[2][1038] , \round_in[2][1037] ,
         \round_in[2][1036] , \round_in[2][1035] , \round_in[2][1034] ,
         \round_in[2][1033] , \round_in[2][1032] , \round_in[2][1031] ,
         \round_in[2][1030] , \round_in[2][1029] , \round_in[2][1028] ,
         \round_in[2][1027] , \round_in[2][1026] , \round_in[2][1025] ,
         \round_in[2][1024] , \round_in[2][1023] , \round_in[2][1022] ,
         \round_in[2][1021] , \round_in[2][1020] , \round_in[2][1019] ,
         \round_in[2][1018] , \round_in[2][1017] , \round_in[2][1016] ,
         \round_in[2][1015] , \round_in[2][1014] , \round_in[2][1013] ,
         \round_in[2][1012] , \round_in[2][1011] , \round_in[2][1010] ,
         \round_in[2][1009] , \round_in[2][1008] , \round_in[2][1007] ,
         \round_in[2][1006] , \round_in[2][1005] , \round_in[2][1004] ,
         \round_in[2][1003] , \round_in[2][1002] , \round_in[2][1001] ,
         \round_in[2][1000] , \round_in[2][999] , \round_in[2][998] ,
         \round_in[2][997] , \round_in[2][996] , \round_in[2][995] ,
         \round_in[2][994] , \round_in[2][993] , \round_in[2][992] ,
         \round_in[2][991] , \round_in[2][990] , \round_in[2][989] ,
         \round_in[2][988] , \round_in[2][987] , \round_in[2][986] ,
         \round_in[2][985] , \round_in[2][984] , \round_in[2][983] ,
         \round_in[2][982] , \round_in[2][981] , \round_in[2][980] ,
         \round_in[2][979] , \round_in[2][978] , \round_in[2][977] ,
         \round_in[2][976] , \round_in[2][975] , \round_in[2][974] ,
         \round_in[2][973] , \round_in[2][972] , \round_in[2][971] ,
         \round_in[2][970] , \round_in[2][969] , \round_in[2][968] ,
         \round_in[2][967] , \round_in[2][966] , \round_in[2][965] ,
         \round_in[2][964] , \round_in[2][963] , \round_in[2][962] ,
         \round_in[2][961] , \round_in[2][960] , \round_in[2][959] ,
         \round_in[2][958] , \round_in[2][957] , \round_in[2][956] ,
         \round_in[2][955] , \round_in[2][954] , \round_in[2][953] ,
         \round_in[2][952] , \round_in[2][951] , \round_in[2][950] ,
         \round_in[2][949] , \round_in[2][948] , \round_in[2][947] ,
         \round_in[2][946] , \round_in[2][945] , \round_in[2][944] ,
         \round_in[2][943] , \round_in[2][942] , \round_in[2][941] ,
         \round_in[2][940] , \round_in[2][939] , \round_in[2][938] ,
         \round_in[2][937] , \round_in[2][936] , \round_in[2][935] ,
         \round_in[2][934] , \round_in[2][933] , \round_in[2][932] ,
         \round_in[2][931] , \round_in[2][930] , \round_in[2][929] ,
         \round_in[2][928] , \round_in[2][927] , \round_in[2][926] ,
         \round_in[2][925] , \round_in[2][924] , \round_in[2][923] ,
         \round_in[2][922] , \round_in[2][921] , \round_in[2][920] ,
         \round_in[2][919] , \round_in[2][918] , \round_in[2][917] ,
         \round_in[2][916] , \round_in[2][915] , \round_in[2][914] ,
         \round_in[2][913] , \round_in[2][912] , \round_in[2][911] ,
         \round_in[2][910] , \round_in[2][909] , \round_in[2][908] ,
         \round_in[2][907] , \round_in[2][906] , \round_in[2][905] ,
         \round_in[2][904] , \round_in[2][903] , \round_in[2][902] ,
         \round_in[2][901] , \round_in[2][900] , \round_in[2][899] ,
         \round_in[2][898] , \round_in[2][897] , \round_in[2][896] ,
         \round_in[2][895] , \round_in[2][894] , \round_in[2][893] ,
         \round_in[2][892] , \round_in[2][891] , \round_in[2][890] ,
         \round_in[2][889] , \round_in[2][888] , \round_in[2][887] ,
         \round_in[2][886] , \round_in[2][885] , \round_in[2][884] ,
         \round_in[2][883] , \round_in[2][882] , \round_in[2][881] ,
         \round_in[2][880] , \round_in[2][879] , \round_in[2][878] ,
         \round_in[2][877] , \round_in[2][876] , \round_in[2][875] ,
         \round_in[2][874] , \round_in[2][873] , \round_in[2][872] ,
         \round_in[2][871] , \round_in[2][870] , \round_in[2][869] ,
         \round_in[2][868] , \round_in[2][867] , \round_in[2][866] ,
         \round_in[2][865] , \round_in[2][864] , \round_in[2][863] ,
         \round_in[2][862] , \round_in[2][861] , \round_in[2][860] ,
         \round_in[2][859] , \round_in[2][858] , \round_in[2][857] ,
         \round_in[2][856] , \round_in[2][855] , \round_in[2][854] ,
         \round_in[2][853] , \round_in[2][852] , \round_in[2][851] ,
         \round_in[2][850] , \round_in[2][849] , \round_in[2][848] ,
         \round_in[2][847] , \round_in[2][846] , \round_in[2][845] ,
         \round_in[2][844] , \round_in[2][843] , \round_in[2][842] ,
         \round_in[2][841] , \round_in[2][840] , \round_in[2][839] ,
         \round_in[2][838] , \round_in[2][837] , \round_in[2][836] ,
         \round_in[2][835] , \round_in[2][834] , \round_in[2][833] ,
         \round_in[2][832] , \round_in[2][831] , \round_in[2][830] ,
         \round_in[2][829] , \round_in[2][828] , \round_in[2][827] ,
         \round_in[2][826] , \round_in[2][825] , \round_in[2][824] ,
         \round_in[2][823] , \round_in[2][822] , \round_in[2][821] ,
         \round_in[2][820] , \round_in[2][819] , \round_in[2][818] ,
         \round_in[2][817] , \round_in[2][816] , \round_in[2][815] ,
         \round_in[2][814] , \round_in[2][813] , \round_in[2][812] ,
         \round_in[2][811] , \round_in[2][810] , \round_in[2][809] ,
         \round_in[2][808] , \round_in[2][807] , \round_in[2][806] ,
         \round_in[2][805] , \round_in[2][804] , \round_in[2][803] ,
         \round_in[2][802] , \round_in[2][801] , \round_in[2][800] ,
         \round_in[2][799] , \round_in[2][798] , \round_in[2][797] ,
         \round_in[2][796] , \round_in[2][795] , \round_in[2][794] ,
         \round_in[2][793] , \round_in[2][792] , \round_in[2][791] ,
         \round_in[2][790] , \round_in[2][789] , \round_in[2][788] ,
         \round_in[2][787] , \round_in[2][786] , \round_in[2][785] ,
         \round_in[2][784] , \round_in[2][783] , \round_in[2][782] ,
         \round_in[2][781] , \round_in[2][780] , \round_in[2][779] ,
         \round_in[2][778] , \round_in[2][777] , \round_in[2][776] ,
         \round_in[2][775] , \round_in[2][774] , \round_in[2][773] ,
         \round_in[2][772] , \round_in[2][771] , \round_in[2][770] ,
         \round_in[2][769] , \round_in[2][768] , \round_in[2][767] ,
         \round_in[2][766] , \round_in[2][765] , \round_in[2][764] ,
         \round_in[2][763] , \round_in[2][762] , \round_in[2][761] ,
         \round_in[2][760] , \round_in[2][759] , \round_in[2][758] ,
         \round_in[2][757] , \round_in[2][756] , \round_in[2][755] ,
         \round_in[2][754] , \round_in[2][753] , \round_in[2][752] ,
         \round_in[2][751] , \round_in[2][750] , \round_in[2][749] ,
         \round_in[2][748] , \round_in[2][747] , \round_in[2][746] ,
         \round_in[2][745] , \round_in[2][744] , \round_in[2][743] ,
         \round_in[2][742] , \round_in[2][741] , \round_in[2][740] ,
         \round_in[2][739] , \round_in[2][738] , \round_in[2][737] ,
         \round_in[2][736] , \round_in[2][735] , \round_in[2][734] ,
         \round_in[2][733] , \round_in[2][732] , \round_in[2][731] ,
         \round_in[2][730] , \round_in[2][729] , \round_in[2][728] ,
         \round_in[2][727] , \round_in[2][726] , \round_in[2][725] ,
         \round_in[2][724] , \round_in[2][723] , \round_in[2][722] ,
         \round_in[2][721] , \round_in[2][720] , \round_in[2][719] ,
         \round_in[2][718] , \round_in[2][717] , \round_in[2][716] ,
         \round_in[2][715] , \round_in[2][714] , \round_in[2][713] ,
         \round_in[2][712] , \round_in[2][711] , \round_in[2][710] ,
         \round_in[2][709] , \round_in[2][708] , \round_in[2][707] ,
         \round_in[2][706] , \round_in[2][705] , \round_in[2][704] ,
         \round_in[2][703] , \round_in[2][702] , \round_in[2][701] ,
         \round_in[2][700] , \round_in[2][699] , \round_in[2][698] ,
         \round_in[2][697] , \round_in[2][696] , \round_in[2][695] ,
         \round_in[2][694] , \round_in[2][693] , \round_in[2][692] ,
         \round_in[2][691] , \round_in[2][690] , \round_in[2][689] ,
         \round_in[2][688] , \round_in[2][687] , \round_in[2][686] ,
         \round_in[2][685] , \round_in[2][684] , \round_in[2][683] ,
         \round_in[2][682] , \round_in[2][681] , \round_in[2][680] ,
         \round_in[2][679] , \round_in[2][678] , \round_in[2][677] ,
         \round_in[2][676] , \round_in[2][675] , \round_in[2][674] ,
         \round_in[2][673] , \round_in[2][672] , \round_in[2][671] ,
         \round_in[2][670] , \round_in[2][669] , \round_in[2][668] ,
         \round_in[2][667] , \round_in[2][666] , \round_in[2][665] ,
         \round_in[2][664] , \round_in[2][663] , \round_in[2][662] ,
         \round_in[2][661] , \round_in[2][660] , \round_in[2][659] ,
         \round_in[2][658] , \round_in[2][657] , \round_in[2][656] ,
         \round_in[2][655] , \round_in[2][654] , \round_in[2][653] ,
         \round_in[2][652] , \round_in[2][651] , \round_in[2][650] ,
         \round_in[2][649] , \round_in[2][648] , \round_in[2][647] ,
         \round_in[2][646] , \round_in[2][645] , \round_in[2][644] ,
         \round_in[2][643] , \round_in[2][642] , \round_in[2][641] ,
         \round_in[2][640] , \round_in[2][639] , \round_in[2][638] ,
         \round_in[2][637] , \round_in[2][636] , \round_in[2][635] ,
         \round_in[2][634] , \round_in[2][633] , \round_in[2][632] ,
         \round_in[2][631] , \round_in[2][630] , \round_in[2][629] ,
         \round_in[2][628] , \round_in[2][627] , \round_in[2][626] ,
         \round_in[2][625] , \round_in[2][624] , \round_in[2][623] ,
         \round_in[2][622] , \round_in[2][621] , \round_in[2][620] ,
         \round_in[2][619] , \round_in[2][618] , \round_in[2][617] ,
         \round_in[2][616] , \round_in[2][615] , \round_in[2][614] ,
         \round_in[2][613] , \round_in[2][612] , \round_in[2][611] ,
         \round_in[2][610] , \round_in[2][609] , \round_in[2][608] ,
         \round_in[2][607] , \round_in[2][606] , \round_in[2][605] ,
         \round_in[2][604] , \round_in[2][603] , \round_in[2][602] ,
         \round_in[2][601] , \round_in[2][600] , \round_in[2][599] ,
         \round_in[2][598] , \round_in[2][597] , \round_in[2][596] ,
         \round_in[2][595] , \round_in[2][594] , \round_in[2][593] ,
         \round_in[2][592] , \round_in[2][591] , \round_in[2][590] ,
         \round_in[2][589] , \round_in[2][588] , \round_in[2][587] ,
         \round_in[2][586] , \round_in[2][585] , \round_in[2][584] ,
         \round_in[2][583] , \round_in[2][582] , \round_in[2][581] ,
         \round_in[2][580] , \round_in[2][579] , \round_in[2][578] ,
         \round_in[2][577] , \round_in[2][576] , \round_in[2][575] ,
         \round_in[2][574] , \round_in[2][573] , \round_in[2][572] ,
         \round_in[2][571] , \round_in[2][570] , \round_in[2][569] ,
         \round_in[2][568] , \round_in[2][567] , \round_in[2][566] ,
         \round_in[2][565] , \round_in[2][564] , \round_in[2][563] ,
         \round_in[2][562] , \round_in[2][561] , \round_in[2][560] ,
         \round_in[2][559] , \round_in[2][558] , \round_in[2][557] ,
         \round_in[2][556] , \round_in[2][555] , \round_in[2][554] ,
         \round_in[2][553] , \round_in[2][552] , \round_in[2][551] ,
         \round_in[2][550] , \round_in[2][549] , \round_in[2][548] ,
         \round_in[2][547] , \round_in[2][546] , \round_in[2][545] ,
         \round_in[2][544] , \round_in[2][543] , \round_in[2][542] ,
         \round_in[2][541] , \round_in[2][540] , \round_in[2][539] ,
         \round_in[2][538] , \round_in[2][537] , \round_in[2][536] ,
         \round_in[2][535] , \round_in[2][534] , \round_in[2][533] ,
         \round_in[2][532] , \round_in[2][531] , \round_in[2][530] ,
         \round_in[2][529] , \round_in[2][528] , \round_in[2][527] ,
         \round_in[2][526] , \round_in[2][525] , \round_in[2][524] ,
         \round_in[2][523] , \round_in[2][522] , \round_in[2][521] ,
         \round_in[2][520] , \round_in[2][519] , \round_in[2][518] ,
         \round_in[2][517] , \round_in[2][516] , \round_in[2][515] ,
         \round_in[2][514] , \round_in[2][513] , \round_in[2][512] ,
         \round_in[2][511] , \round_in[2][510] , \round_in[2][509] ,
         \round_in[2][508] , \round_in[2][507] , \round_in[2][506] ,
         \round_in[2][505] , \round_in[2][504] , \round_in[2][503] ,
         \round_in[2][502] , \round_in[2][501] , \round_in[2][500] ,
         \round_in[2][499] , \round_in[2][498] , \round_in[2][497] ,
         \round_in[2][496] , \round_in[2][495] , \round_in[2][494] ,
         \round_in[2][493] , \round_in[2][492] , \round_in[2][491] ,
         \round_in[2][490] , \round_in[2][489] , \round_in[2][488] ,
         \round_in[2][487] , \round_in[2][486] , \round_in[2][485] ,
         \round_in[2][484] , \round_in[2][483] , \round_in[2][482] ,
         \round_in[2][481] , \round_in[2][480] , \round_in[2][479] ,
         \round_in[2][478] , \round_in[2][477] , \round_in[2][476] ,
         \round_in[2][475] , \round_in[2][474] , \round_in[2][473] ,
         \round_in[2][472] , \round_in[2][471] , \round_in[2][470] ,
         \round_in[2][469] , \round_in[2][468] , \round_in[2][467] ,
         \round_in[2][466] , \round_in[2][465] , \round_in[2][464] ,
         \round_in[2][463] , \round_in[2][462] , \round_in[2][461] ,
         \round_in[2][460] , \round_in[2][459] , \round_in[2][458] ,
         \round_in[2][457] , \round_in[2][456] , \round_in[2][455] ,
         \round_in[2][454] , \round_in[2][453] , \round_in[2][452] ,
         \round_in[2][451] , \round_in[2][450] , \round_in[2][449] ,
         \round_in[2][448] , \round_in[2][447] , \round_in[2][446] ,
         \round_in[2][445] , \round_in[2][444] , \round_in[2][443] ,
         \round_in[2][442] , \round_in[2][441] , \round_in[2][440] ,
         \round_in[2][439] , \round_in[2][438] , \round_in[2][437] ,
         \round_in[2][436] , \round_in[2][435] , \round_in[2][434] ,
         \round_in[2][433] , \round_in[2][432] , \round_in[2][431] ,
         \round_in[2][430] , \round_in[2][429] , \round_in[2][428] ,
         \round_in[2][427] , \round_in[2][426] , \round_in[2][425] ,
         \round_in[2][424] , \round_in[2][423] , \round_in[2][422] ,
         \round_in[2][421] , \round_in[2][420] , \round_in[2][419] ,
         \round_in[2][418] , \round_in[2][417] , \round_in[2][416] ,
         \round_in[2][415] , \round_in[2][414] , \round_in[2][413] ,
         \round_in[2][412] , \round_in[2][411] , \round_in[2][410] ,
         \round_in[2][409] , \round_in[2][408] , \round_in[2][407] ,
         \round_in[2][406] , \round_in[2][405] , \round_in[2][404] ,
         \round_in[2][403] , \round_in[2][402] , \round_in[2][401] ,
         \round_in[2][400] , \round_in[2][399] , \round_in[2][398] ,
         \round_in[2][397] , \round_in[2][396] , \round_in[2][395] ,
         \round_in[2][394] , \round_in[2][393] , \round_in[2][392] ,
         \round_in[2][391] , \round_in[2][390] , \round_in[2][389] ,
         \round_in[2][388] , \round_in[2][387] , \round_in[2][386] ,
         \round_in[2][385] , \round_in[2][384] , \round_in[2][383] ,
         \round_in[2][382] , \round_in[2][381] , \round_in[2][380] ,
         \round_in[2][379] , \round_in[2][378] , \round_in[2][377] ,
         \round_in[2][376] , \round_in[2][375] , \round_in[2][374] ,
         \round_in[2][373] , \round_in[2][372] , \round_in[2][371] ,
         \round_in[2][370] , \round_in[2][369] , \round_in[2][368] ,
         \round_in[2][367] , \round_in[2][366] , \round_in[2][365] ,
         \round_in[2][364] , \round_in[2][363] , \round_in[2][362] ,
         \round_in[2][361] , \round_in[2][360] , \round_in[2][359] ,
         \round_in[2][358] , \round_in[2][357] , \round_in[2][356] ,
         \round_in[2][355] , \round_in[2][354] , \round_in[2][353] ,
         \round_in[2][352] , \round_in[2][351] , \round_in[2][350] ,
         \round_in[2][349] , \round_in[2][348] , \round_in[2][347] ,
         \round_in[2][346] , \round_in[2][345] , \round_in[2][344] ,
         \round_in[2][343] , \round_in[2][342] , \round_in[2][341] ,
         \round_in[2][340] , \round_in[2][339] , \round_in[2][338] ,
         \round_in[2][337] , \round_in[2][336] , \round_in[2][335] ,
         \round_in[2][334] , \round_in[2][333] , \round_in[2][332] ,
         \round_in[2][331] , \round_in[2][330] , \round_in[2][329] ,
         \round_in[2][328] , \round_in[2][327] , \round_in[2][326] ,
         \round_in[2][325] , \round_in[2][324] , \round_in[2][323] ,
         \round_in[2][322] , \round_in[2][321] , \round_in[2][320] ,
         \round_in[2][319] , \round_in[2][318] , \round_in[2][317] ,
         \round_in[2][316] , \round_in[2][315] , \round_in[2][314] ,
         \round_in[2][313] , \round_in[2][312] , \round_in[2][311] ,
         \round_in[2][310] , \round_in[2][309] , \round_in[2][308] ,
         \round_in[2][307] , \round_in[2][306] , \round_in[2][305] ,
         \round_in[2][304] , \round_in[2][303] , \round_in[2][302] ,
         \round_in[2][301] , \round_in[2][300] , \round_in[2][299] ,
         \round_in[2][298] , \round_in[2][297] , \round_in[2][296] ,
         \round_in[2][295] , \round_in[2][294] , \round_in[2][293] ,
         \round_in[2][292] , \round_in[2][291] , \round_in[2][290] ,
         \round_in[2][289] , \round_in[2][288] , \round_in[2][287] ,
         \round_in[2][286] , \round_in[2][285] , \round_in[2][284] ,
         \round_in[2][283] , \round_in[2][282] , \round_in[2][281] ,
         \round_in[2][280] , \round_in[2][279] , \round_in[2][278] ,
         \round_in[2][277] , \round_in[2][276] , \round_in[2][275] ,
         \round_in[2][274] , \round_in[2][273] , \round_in[2][272] ,
         \round_in[2][271] , \round_in[2][270] , \round_in[2][269] ,
         \round_in[2][268] , \round_in[2][267] , \round_in[2][266] ,
         \round_in[2][265] , \round_in[2][264] , \round_in[2][263] ,
         \round_in[2][262] , \round_in[2][261] , \round_in[2][260] ,
         \round_in[2][259] , \round_in[2][258] , \round_in[2][257] ,
         \round_in[2][256] , \round_in[2][255] , \round_in[2][254] ,
         \round_in[2][253] , \round_in[2][252] , \round_in[2][251] ,
         \round_in[2][250] , \round_in[2][249] , \round_in[2][248] ,
         \round_in[2][247] , \round_in[2][246] , \round_in[2][245] ,
         \round_in[2][244] , \round_in[2][243] , \round_in[2][242] ,
         \round_in[2][241] , \round_in[2][240] , \round_in[2][239] ,
         \round_in[2][238] , \round_in[2][237] , \round_in[2][236] ,
         \round_in[2][235] , \round_in[2][234] , \round_in[2][233] ,
         \round_in[2][232] , \round_in[2][231] , \round_in[2][230] ,
         \round_in[2][229] , \round_in[2][228] , \round_in[2][227] ,
         \round_in[2][226] , \round_in[2][225] , \round_in[2][224] ,
         \round_in[2][223] , \round_in[2][222] , \round_in[2][221] ,
         \round_in[2][220] , \round_in[2][219] , \round_in[2][218] ,
         \round_in[2][217] , \round_in[2][216] , \round_in[2][215] ,
         \round_in[2][214] , \round_in[2][213] , \round_in[2][212] ,
         \round_in[2][211] , \round_in[2][210] , \round_in[2][209] ,
         \round_in[2][208] , \round_in[2][207] , \round_in[2][206] ,
         \round_in[2][205] , \round_in[2][204] , \round_in[2][203] ,
         \round_in[2][202] , \round_in[2][201] , \round_in[2][200] ,
         \round_in[2][199] , \round_in[2][198] , \round_in[2][197] ,
         \round_in[2][196] , \round_in[2][195] , \round_in[2][194] ,
         \round_in[2][193] , \round_in[2][192] , \round_in[2][191] ,
         \round_in[2][190] , \round_in[2][189] , \round_in[2][188] ,
         \round_in[2][187] , \round_in[2][186] , \round_in[2][185] ,
         \round_in[2][184] , \round_in[2][183] , \round_in[2][182] ,
         \round_in[2][181] , \round_in[2][180] , \round_in[2][179] ,
         \round_in[2][178] , \round_in[2][177] , \round_in[2][176] ,
         \round_in[2][175] , \round_in[2][174] , \round_in[2][173] ,
         \round_in[2][172] , \round_in[2][171] , \round_in[2][170] ,
         \round_in[2][169] , \round_in[2][168] , \round_in[2][167] ,
         \round_in[2][166] , \round_in[2][165] , \round_in[2][164] ,
         \round_in[2][163] , \round_in[2][162] , \round_in[2][161] ,
         \round_in[2][160] , \round_in[2][159] , \round_in[2][158] ,
         \round_in[2][157] , \round_in[2][156] , \round_in[2][155] ,
         \round_in[2][154] , \round_in[2][153] , \round_in[2][152] ,
         \round_in[2][151] , \round_in[2][150] , \round_in[2][149] ,
         \round_in[2][148] , \round_in[2][147] , \round_in[2][146] ,
         \round_in[2][145] , \round_in[2][144] , \round_in[2][143] ,
         \round_in[2][142] , \round_in[2][141] , \round_in[2][140] ,
         \round_in[2][139] , \round_in[2][138] , \round_in[2][137] ,
         \round_in[2][136] , \round_in[2][135] , \round_in[2][134] ,
         \round_in[2][133] , \round_in[2][132] , \round_in[2][131] ,
         \round_in[2][130] , \round_in[2][129] , \round_in[2][128] ,
         \round_in[2][127] , \round_in[2][126] , \round_in[2][125] ,
         \round_in[2][124] , \round_in[2][123] , \round_in[2][122] ,
         \round_in[2][121] , \round_in[2][120] , \round_in[2][119] ,
         \round_in[2][118] , \round_in[2][117] , \round_in[2][116] ,
         \round_in[2][115] , \round_in[2][114] , \round_in[2][113] ,
         \round_in[2][112] , \round_in[2][111] , \round_in[2][110] ,
         \round_in[2][109] , \round_in[2][108] , \round_in[2][107] ,
         \round_in[2][106] , \round_in[2][105] , \round_in[2][104] ,
         \round_in[2][103] , \round_in[2][102] , \round_in[2][101] ,
         \round_in[2][100] , \round_in[2][99] , \round_in[2][98] ,
         \round_in[2][97] , \round_in[2][96] , \round_in[2][95] ,
         \round_in[2][94] , \round_in[2][93] , \round_in[2][92] ,
         \round_in[2][91] , \round_in[2][90] , \round_in[2][89] ,
         \round_in[2][88] , \round_in[2][87] , \round_in[2][86] ,
         \round_in[2][85] , \round_in[2][84] , \round_in[2][83] ,
         \round_in[2][82] , \round_in[2][81] , \round_in[2][80] ,
         \round_in[2][79] , \round_in[2][78] , \round_in[2][77] ,
         \round_in[2][76] , \round_in[2][75] , \round_in[2][74] ,
         \round_in[2][73] , \round_in[2][72] , \round_in[2][71] ,
         \round_in[2][70] , \round_in[2][69] , \round_in[2][68] ,
         \round_in[2][67] , \round_in[2][66] , \round_in[2][65] ,
         \round_in[2][64] , \round_in[2][63] , \round_in[2][62] ,
         \round_in[2][61] , \round_in[2][60] , \round_in[2][59] ,
         \round_in[2][58] , \round_in[2][57] , \round_in[2][56] ,
         \round_in[2][55] , \round_in[2][54] , \round_in[2][53] ,
         \round_in[2][52] , \round_in[2][51] , \round_in[2][50] ,
         \round_in[2][49] , \round_in[2][48] , \round_in[2][47] ,
         \round_in[2][46] , \round_in[2][45] , \round_in[2][44] ,
         \round_in[2][43] , \round_in[2][42] , \round_in[2][41] ,
         \round_in[2][40] , \round_in[2][39] , \round_in[2][38] ,
         \round_in[2][37] , \round_in[2][36] , \round_in[2][35] ,
         \round_in[2][34] , \round_in[2][33] , \round_in[2][32] ,
         \round_in[2][31] , \round_in[2][30] , \round_in[2][29] ,
         \round_in[2][28] , \round_in[2][27] , \round_in[2][26] ,
         \round_in[2][25] , \round_in[2][24] , \round_in[2][23] ,
         \round_in[2][22] , \round_in[2][21] , \round_in[2][20] ,
         \round_in[2][19] , \round_in[2][18] , \round_in[2][17] ,
         \round_in[2][16] , \round_in[2][15] , \round_in[2][14] ,
         \round_in[2][13] , \round_in[2][12] , \round_in[2][11] ,
         \round_in[2][10] , \round_in[2][9] , \round_in[2][8] ,
         \round_in[2][7] , \round_in[2][6] , \round_in[2][5] ,
         \round_in[2][4] , \round_in[2][3] , \round_in[2][2] ,
         \round_in[2][1] , \round_in[2][0] , \round_in[1][1599] ,
         \round_in[1][1598] , \round_in[1][1597] , \round_in[1][1596] ,
         \round_in[1][1595] , \round_in[1][1594] , \round_in[1][1593] ,
         \round_in[1][1592] , \round_in[1][1591] , \round_in[1][1590] ,
         \round_in[1][1589] , \round_in[1][1588] , \round_in[1][1587] ,
         \round_in[1][1586] , \round_in[1][1585] , \round_in[1][1584] ,
         \round_in[1][1583] , \round_in[1][1582] , \round_in[1][1581] ,
         \round_in[1][1580] , \round_in[1][1579] , \round_in[1][1578] ,
         \round_in[1][1577] , \round_in[1][1576] , \round_in[1][1575] ,
         \round_in[1][1574] , \round_in[1][1573] , \round_in[1][1572] ,
         \round_in[1][1571] , \round_in[1][1570] , \round_in[1][1569] ,
         \round_in[1][1568] , \round_in[1][1567] , \round_in[1][1566] ,
         \round_in[1][1565] , \round_in[1][1564] , \round_in[1][1563] ,
         \round_in[1][1562] , \round_in[1][1561] , \round_in[1][1560] ,
         \round_in[1][1559] , \round_in[1][1558] , \round_in[1][1557] ,
         \round_in[1][1556] , \round_in[1][1555] , \round_in[1][1554] ,
         \round_in[1][1553] , \round_in[1][1552] , \round_in[1][1551] ,
         \round_in[1][1550] , \round_in[1][1549] , \round_in[1][1548] ,
         \round_in[1][1547] , \round_in[1][1546] , \round_in[1][1545] ,
         \round_in[1][1544] , \round_in[1][1543] , \round_in[1][1542] ,
         \round_in[1][1541] , \round_in[1][1540] , \round_in[1][1539] ,
         \round_in[1][1538] , \round_in[1][1537] , \round_in[1][1536] ,
         \round_in[1][1535] , \round_in[1][1534] , \round_in[1][1533] ,
         \round_in[1][1532] , \round_in[1][1531] , \round_in[1][1530] ,
         \round_in[1][1529] , \round_in[1][1528] , \round_in[1][1527] ,
         \round_in[1][1526] , \round_in[1][1525] , \round_in[1][1524] ,
         \round_in[1][1523] , \round_in[1][1522] , \round_in[1][1521] ,
         \round_in[1][1520] , \round_in[1][1519] , \round_in[1][1518] ,
         \round_in[1][1517] , \round_in[1][1516] , \round_in[1][1515] ,
         \round_in[1][1514] , \round_in[1][1513] , \round_in[1][1512] ,
         \round_in[1][1511] , \round_in[1][1510] , \round_in[1][1509] ,
         \round_in[1][1508] , \round_in[1][1507] , \round_in[1][1506] ,
         \round_in[1][1505] , \round_in[1][1504] , \round_in[1][1503] ,
         \round_in[1][1502] , \round_in[1][1501] , \round_in[1][1500] ,
         \round_in[1][1499] , \round_in[1][1498] , \round_in[1][1497] ,
         \round_in[1][1496] , \round_in[1][1495] , \round_in[1][1494] ,
         \round_in[1][1493] , \round_in[1][1492] , \round_in[1][1491] ,
         \round_in[1][1490] , \round_in[1][1489] , \round_in[1][1488] ,
         \round_in[1][1487] , \round_in[1][1486] , \round_in[1][1485] ,
         \round_in[1][1484] , \round_in[1][1483] , \round_in[1][1482] ,
         \round_in[1][1481] , \round_in[1][1480] , \round_in[1][1479] ,
         \round_in[1][1478] , \round_in[1][1477] , \round_in[1][1476] ,
         \round_in[1][1475] , \round_in[1][1474] , \round_in[1][1473] ,
         \round_in[1][1472] , \round_in[1][1471] , \round_in[1][1470] ,
         \round_in[1][1469] , \round_in[1][1468] , \round_in[1][1467] ,
         \round_in[1][1466] , \round_in[1][1465] , \round_in[1][1464] ,
         \round_in[1][1463] , \round_in[1][1462] , \round_in[1][1461] ,
         \round_in[1][1460] , \round_in[1][1459] , \round_in[1][1458] ,
         \round_in[1][1457] , \round_in[1][1456] , \round_in[1][1455] ,
         \round_in[1][1454] , \round_in[1][1453] , \round_in[1][1452] ,
         \round_in[1][1451] , \round_in[1][1450] , \round_in[1][1449] ,
         \round_in[1][1448] , \round_in[1][1447] , \round_in[1][1446] ,
         \round_in[1][1445] , \round_in[1][1444] , \round_in[1][1443] ,
         \round_in[1][1442] , \round_in[1][1441] , \round_in[1][1440] ,
         \round_in[1][1439] , \round_in[1][1438] , \round_in[1][1437] ,
         \round_in[1][1436] , \round_in[1][1435] , \round_in[1][1434] ,
         \round_in[1][1433] , \round_in[1][1432] , \round_in[1][1431] ,
         \round_in[1][1430] , \round_in[1][1429] , \round_in[1][1428] ,
         \round_in[1][1427] , \round_in[1][1426] , \round_in[1][1425] ,
         \round_in[1][1424] , \round_in[1][1423] , \round_in[1][1422] ,
         \round_in[1][1421] , \round_in[1][1420] , \round_in[1][1419] ,
         \round_in[1][1418] , \round_in[1][1417] , \round_in[1][1416] ,
         \round_in[1][1415] , \round_in[1][1414] , \round_in[1][1413] ,
         \round_in[1][1412] , \round_in[1][1411] , \round_in[1][1410] ,
         \round_in[1][1409] , \round_in[1][1408] , \round_in[1][1407] ,
         \round_in[1][1406] , \round_in[1][1405] , \round_in[1][1404] ,
         \round_in[1][1403] , \round_in[1][1402] , \round_in[1][1401] ,
         \round_in[1][1400] , \round_in[1][1399] , \round_in[1][1398] ,
         \round_in[1][1397] , \round_in[1][1396] , \round_in[1][1395] ,
         \round_in[1][1394] , \round_in[1][1393] , \round_in[1][1392] ,
         \round_in[1][1391] , \round_in[1][1390] , \round_in[1][1389] ,
         \round_in[1][1388] , \round_in[1][1387] , \round_in[1][1386] ,
         \round_in[1][1385] , \round_in[1][1384] , \round_in[1][1383] ,
         \round_in[1][1382] , \round_in[1][1381] , \round_in[1][1380] ,
         \round_in[1][1379] , \round_in[1][1378] , \round_in[1][1377] ,
         \round_in[1][1376] , \round_in[1][1375] , \round_in[1][1374] ,
         \round_in[1][1373] , \round_in[1][1372] , \round_in[1][1371] ,
         \round_in[1][1370] , \round_in[1][1369] , \round_in[1][1368] ,
         \round_in[1][1367] , \round_in[1][1366] , \round_in[1][1365] ,
         \round_in[1][1364] , \round_in[1][1363] , \round_in[1][1362] ,
         \round_in[1][1361] , \round_in[1][1360] , \round_in[1][1359] ,
         \round_in[1][1358] , \round_in[1][1357] , \round_in[1][1356] ,
         \round_in[1][1355] , \round_in[1][1354] , \round_in[1][1353] ,
         \round_in[1][1352] , \round_in[1][1351] , \round_in[1][1350] ,
         \round_in[1][1349] , \round_in[1][1348] , \round_in[1][1347] ,
         \round_in[1][1346] , \round_in[1][1345] , \round_in[1][1344] ,
         \round_in[1][1343] , \round_in[1][1342] , \round_in[1][1341] ,
         \round_in[1][1340] , \round_in[1][1339] , \round_in[1][1338] ,
         \round_in[1][1337] , \round_in[1][1336] , \round_in[1][1335] ,
         \round_in[1][1334] , \round_in[1][1333] , \round_in[1][1332] ,
         \round_in[1][1331] , \round_in[1][1330] , \round_in[1][1329] ,
         \round_in[1][1328] , \round_in[1][1327] , \round_in[1][1326] ,
         \round_in[1][1325] , \round_in[1][1324] , \round_in[1][1323] ,
         \round_in[1][1322] , \round_in[1][1321] , \round_in[1][1320] ,
         \round_in[1][1319] , \round_in[1][1318] , \round_in[1][1317] ,
         \round_in[1][1316] , \round_in[1][1315] , \round_in[1][1314] ,
         \round_in[1][1313] , \round_in[1][1312] , \round_in[1][1311] ,
         \round_in[1][1310] , \round_in[1][1309] , \round_in[1][1308] ,
         \round_in[1][1307] , \round_in[1][1306] , \round_in[1][1305] ,
         \round_in[1][1304] , \round_in[1][1303] , \round_in[1][1302] ,
         \round_in[1][1301] , \round_in[1][1300] , \round_in[1][1299] ,
         \round_in[1][1298] , \round_in[1][1297] , \round_in[1][1296] ,
         \round_in[1][1295] , \round_in[1][1294] , \round_in[1][1293] ,
         \round_in[1][1292] , \round_in[1][1291] , \round_in[1][1290] ,
         \round_in[1][1289] , \round_in[1][1288] , \round_in[1][1287] ,
         \round_in[1][1286] , \round_in[1][1285] , \round_in[1][1284] ,
         \round_in[1][1283] , \round_in[1][1282] , \round_in[1][1281] ,
         \round_in[1][1280] , \round_in[1][1279] , \round_in[1][1278] ,
         \round_in[1][1277] , \round_in[1][1276] , \round_in[1][1275] ,
         \round_in[1][1274] , \round_in[1][1273] , \round_in[1][1272] ,
         \round_in[1][1271] , \round_in[1][1270] , \round_in[1][1269] ,
         \round_in[1][1268] , \round_in[1][1267] , \round_in[1][1266] ,
         \round_in[1][1265] , \round_in[1][1264] , \round_in[1][1263] ,
         \round_in[1][1262] , \round_in[1][1261] , \round_in[1][1260] ,
         \round_in[1][1259] , \round_in[1][1258] , \round_in[1][1257] ,
         \round_in[1][1256] , \round_in[1][1255] , \round_in[1][1254] ,
         \round_in[1][1253] , \round_in[1][1252] , \round_in[1][1251] ,
         \round_in[1][1250] , \round_in[1][1249] , \round_in[1][1248] ,
         \round_in[1][1247] , \round_in[1][1246] , \round_in[1][1245] ,
         \round_in[1][1244] , \round_in[1][1243] , \round_in[1][1242] ,
         \round_in[1][1241] , \round_in[1][1240] , \round_in[1][1239] ,
         \round_in[1][1238] , \round_in[1][1237] , \round_in[1][1236] ,
         \round_in[1][1235] , \round_in[1][1234] , \round_in[1][1233] ,
         \round_in[1][1232] , \round_in[1][1231] , \round_in[1][1230] ,
         \round_in[1][1229] , \round_in[1][1228] , \round_in[1][1227] ,
         \round_in[1][1226] , \round_in[1][1225] , \round_in[1][1224] ,
         \round_in[1][1223] , \round_in[1][1222] , \round_in[1][1221] ,
         \round_in[1][1220] , \round_in[1][1219] , \round_in[1][1218] ,
         \round_in[1][1217] , \round_in[1][1216] , \round_in[1][1215] ,
         \round_in[1][1214] , \round_in[1][1213] , \round_in[1][1212] ,
         \round_in[1][1211] , \round_in[1][1210] , \round_in[1][1209] ,
         \round_in[1][1208] , \round_in[1][1207] , \round_in[1][1206] ,
         \round_in[1][1205] , \round_in[1][1204] , \round_in[1][1203] ,
         \round_in[1][1202] , \round_in[1][1201] , \round_in[1][1200] ,
         \round_in[1][1199] , \round_in[1][1198] , \round_in[1][1197] ,
         \round_in[1][1196] , \round_in[1][1195] , \round_in[1][1194] ,
         \round_in[1][1193] , \round_in[1][1192] , \round_in[1][1191] ,
         \round_in[1][1190] , \round_in[1][1189] , \round_in[1][1188] ,
         \round_in[1][1187] , \round_in[1][1186] , \round_in[1][1185] ,
         \round_in[1][1184] , \round_in[1][1183] , \round_in[1][1182] ,
         \round_in[1][1181] , \round_in[1][1180] , \round_in[1][1179] ,
         \round_in[1][1178] , \round_in[1][1177] , \round_in[1][1176] ,
         \round_in[1][1175] , \round_in[1][1174] , \round_in[1][1173] ,
         \round_in[1][1172] , \round_in[1][1171] , \round_in[1][1170] ,
         \round_in[1][1169] , \round_in[1][1168] , \round_in[1][1167] ,
         \round_in[1][1166] , \round_in[1][1165] , \round_in[1][1164] ,
         \round_in[1][1163] , \round_in[1][1162] , \round_in[1][1161] ,
         \round_in[1][1160] , \round_in[1][1159] , \round_in[1][1158] ,
         \round_in[1][1157] , \round_in[1][1156] , \round_in[1][1155] ,
         \round_in[1][1154] , \round_in[1][1153] , \round_in[1][1152] ,
         \round_in[1][1151] , \round_in[1][1150] , \round_in[1][1149] ,
         \round_in[1][1148] , \round_in[1][1147] , \round_in[1][1146] ,
         \round_in[1][1145] , \round_in[1][1144] , \round_in[1][1143] ,
         \round_in[1][1142] , \round_in[1][1141] , \round_in[1][1140] ,
         \round_in[1][1139] , \round_in[1][1138] , \round_in[1][1137] ,
         \round_in[1][1136] , \round_in[1][1135] , \round_in[1][1134] ,
         \round_in[1][1133] , \round_in[1][1132] , \round_in[1][1131] ,
         \round_in[1][1130] , \round_in[1][1129] , \round_in[1][1128] ,
         \round_in[1][1127] , \round_in[1][1126] , \round_in[1][1125] ,
         \round_in[1][1124] , \round_in[1][1123] , \round_in[1][1122] ,
         \round_in[1][1121] , \round_in[1][1120] , \round_in[1][1119] ,
         \round_in[1][1118] , \round_in[1][1117] , \round_in[1][1116] ,
         \round_in[1][1115] , \round_in[1][1114] , \round_in[1][1113] ,
         \round_in[1][1112] , \round_in[1][1111] , \round_in[1][1110] ,
         \round_in[1][1109] , \round_in[1][1108] , \round_in[1][1107] ,
         \round_in[1][1106] , \round_in[1][1105] , \round_in[1][1104] ,
         \round_in[1][1103] , \round_in[1][1102] , \round_in[1][1101] ,
         \round_in[1][1100] , \round_in[1][1099] , \round_in[1][1098] ,
         \round_in[1][1097] , \round_in[1][1096] , \round_in[1][1095] ,
         \round_in[1][1094] , \round_in[1][1093] , \round_in[1][1092] ,
         \round_in[1][1091] , \round_in[1][1090] , \round_in[1][1089] ,
         \round_in[1][1088] , \round_in[1][1087] , \round_in[1][1086] ,
         \round_in[1][1085] , \round_in[1][1084] , \round_in[1][1083] ,
         \round_in[1][1082] , \round_in[1][1081] , \round_in[1][1080] ,
         \round_in[1][1079] , \round_in[1][1078] , \round_in[1][1077] ,
         \round_in[1][1076] , \round_in[1][1075] , \round_in[1][1074] ,
         \round_in[1][1073] , \round_in[1][1072] , \round_in[1][1071] ,
         \round_in[1][1070] , \round_in[1][1069] , \round_in[1][1068] ,
         \round_in[1][1067] , \round_in[1][1066] , \round_in[1][1065] ,
         \round_in[1][1064] , \round_in[1][1063] , \round_in[1][1062] ,
         \round_in[1][1061] , \round_in[1][1060] , \round_in[1][1059] ,
         \round_in[1][1058] , \round_in[1][1057] , \round_in[1][1056] ,
         \round_in[1][1055] , \round_in[1][1054] , \round_in[1][1053] ,
         \round_in[1][1052] , \round_in[1][1051] , \round_in[1][1050] ,
         \round_in[1][1049] , \round_in[1][1048] , \round_in[1][1047] ,
         \round_in[1][1046] , \round_in[1][1045] , \round_in[1][1044] ,
         \round_in[1][1043] , \round_in[1][1042] , \round_in[1][1041] ,
         \round_in[1][1040] , \round_in[1][1039] , \round_in[1][1038] ,
         \round_in[1][1037] , \round_in[1][1036] , \round_in[1][1035] ,
         \round_in[1][1034] , \round_in[1][1033] , \round_in[1][1032] ,
         \round_in[1][1031] , \round_in[1][1030] , \round_in[1][1029] ,
         \round_in[1][1028] , \round_in[1][1027] , \round_in[1][1026] ,
         \round_in[1][1025] , \round_in[1][1024] , \round_in[1][1023] ,
         \round_in[1][1022] , \round_in[1][1021] , \round_in[1][1020] ,
         \round_in[1][1019] , \round_in[1][1018] , \round_in[1][1017] ,
         \round_in[1][1016] , \round_in[1][1015] , \round_in[1][1014] ,
         \round_in[1][1013] , \round_in[1][1012] , \round_in[1][1011] ,
         \round_in[1][1010] , \round_in[1][1009] , \round_in[1][1008] ,
         \round_in[1][1007] , \round_in[1][1006] , \round_in[1][1005] ,
         \round_in[1][1004] , \round_in[1][1003] , \round_in[1][1002] ,
         \round_in[1][1001] , \round_in[1][1000] , \round_in[1][999] ,
         \round_in[1][998] , \round_in[1][997] , \round_in[1][996] ,
         \round_in[1][995] , \round_in[1][994] , \round_in[1][993] ,
         \round_in[1][992] , \round_in[1][991] , \round_in[1][990] ,
         \round_in[1][989] , \round_in[1][988] , \round_in[1][987] ,
         \round_in[1][986] , \round_in[1][985] , \round_in[1][984] ,
         \round_in[1][983] , \round_in[1][982] , \round_in[1][981] ,
         \round_in[1][980] , \round_in[1][979] , \round_in[1][978] ,
         \round_in[1][977] , \round_in[1][976] , \round_in[1][975] ,
         \round_in[1][974] , \round_in[1][973] , \round_in[1][972] ,
         \round_in[1][971] , \round_in[1][970] , \round_in[1][969] ,
         \round_in[1][968] , \round_in[1][967] , \round_in[1][966] ,
         \round_in[1][965] , \round_in[1][964] , \round_in[1][963] ,
         \round_in[1][962] , \round_in[1][961] , \round_in[1][960] ,
         \round_in[1][959] , \round_in[1][958] , \round_in[1][957] ,
         \round_in[1][956] , \round_in[1][955] , \round_in[1][954] ,
         \round_in[1][953] , \round_in[1][952] , \round_in[1][951] ,
         \round_in[1][950] , \round_in[1][949] , \round_in[1][948] ,
         \round_in[1][947] , \round_in[1][946] , \round_in[1][945] ,
         \round_in[1][944] , \round_in[1][943] , \round_in[1][942] ,
         \round_in[1][941] , \round_in[1][940] , \round_in[1][939] ,
         \round_in[1][938] , \round_in[1][937] , \round_in[1][936] ,
         \round_in[1][935] , \round_in[1][934] , \round_in[1][933] ,
         \round_in[1][932] , \round_in[1][931] , \round_in[1][930] ,
         \round_in[1][929] , \round_in[1][928] , \round_in[1][927] ,
         \round_in[1][926] , \round_in[1][925] , \round_in[1][924] ,
         \round_in[1][923] , \round_in[1][922] , \round_in[1][921] ,
         \round_in[1][920] , \round_in[1][919] , \round_in[1][918] ,
         \round_in[1][917] , \round_in[1][916] , \round_in[1][915] ,
         \round_in[1][914] , \round_in[1][913] , \round_in[1][912] ,
         \round_in[1][911] , \round_in[1][910] , \round_in[1][909] ,
         \round_in[1][908] , \round_in[1][907] , \round_in[1][906] ,
         \round_in[1][905] , \round_in[1][904] , \round_in[1][903] ,
         \round_in[1][902] , \round_in[1][901] , \round_in[1][900] ,
         \round_in[1][899] , \round_in[1][898] , \round_in[1][897] ,
         \round_in[1][896] , \round_in[1][895] , \round_in[1][894] ,
         \round_in[1][893] , \round_in[1][892] , \round_in[1][891] ,
         \round_in[1][890] , \round_in[1][889] , \round_in[1][888] ,
         \round_in[1][887] , \round_in[1][886] , \round_in[1][885] ,
         \round_in[1][884] , \round_in[1][883] , \round_in[1][882] ,
         \round_in[1][881] , \round_in[1][880] , \round_in[1][879] ,
         \round_in[1][878] , \round_in[1][877] , \round_in[1][876] ,
         \round_in[1][875] , \round_in[1][874] , \round_in[1][873] ,
         \round_in[1][872] , \round_in[1][871] , \round_in[1][870] ,
         \round_in[1][869] , \round_in[1][868] , \round_in[1][867] ,
         \round_in[1][866] , \round_in[1][865] , \round_in[1][864] ,
         \round_in[1][863] , \round_in[1][862] , \round_in[1][861] ,
         \round_in[1][860] , \round_in[1][859] , \round_in[1][858] ,
         \round_in[1][857] , \round_in[1][856] , \round_in[1][855] ,
         \round_in[1][854] , \round_in[1][853] , \round_in[1][852] ,
         \round_in[1][851] , \round_in[1][850] , \round_in[1][849] ,
         \round_in[1][848] , \round_in[1][847] , \round_in[1][846] ,
         \round_in[1][845] , \round_in[1][844] , \round_in[1][843] ,
         \round_in[1][842] , \round_in[1][841] , \round_in[1][840] ,
         \round_in[1][839] , \round_in[1][838] , \round_in[1][837] ,
         \round_in[1][836] , \round_in[1][835] , \round_in[1][834] ,
         \round_in[1][833] , \round_in[1][832] , \round_in[1][831] ,
         \round_in[1][830] , \round_in[1][829] , \round_in[1][828] ,
         \round_in[1][827] , \round_in[1][826] , \round_in[1][825] ,
         \round_in[1][824] , \round_in[1][823] , \round_in[1][822] ,
         \round_in[1][821] , \round_in[1][820] , \round_in[1][819] ,
         \round_in[1][818] , \round_in[1][817] , \round_in[1][816] ,
         \round_in[1][815] , \round_in[1][814] , \round_in[1][813] ,
         \round_in[1][812] , \round_in[1][811] , \round_in[1][810] ,
         \round_in[1][809] , \round_in[1][808] , \round_in[1][807] ,
         \round_in[1][806] , \round_in[1][805] , \round_in[1][804] ,
         \round_in[1][803] , \round_in[1][802] , \round_in[1][801] ,
         \round_in[1][800] , \round_in[1][799] , \round_in[1][798] ,
         \round_in[1][797] , \round_in[1][796] , \round_in[1][795] ,
         \round_in[1][794] , \round_in[1][793] , \round_in[1][792] ,
         \round_in[1][791] , \round_in[1][790] , \round_in[1][789] ,
         \round_in[1][788] , \round_in[1][787] , \round_in[1][786] ,
         \round_in[1][785] , \round_in[1][784] , \round_in[1][783] ,
         \round_in[1][782] , \round_in[1][781] , \round_in[1][780] ,
         \round_in[1][779] , \round_in[1][778] , \round_in[1][777] ,
         \round_in[1][776] , \round_in[1][775] , \round_in[1][774] ,
         \round_in[1][773] , \round_in[1][772] , \round_in[1][771] ,
         \round_in[1][770] , \round_in[1][769] , \round_in[1][768] ,
         \round_in[1][767] , \round_in[1][766] , \round_in[1][765] ,
         \round_in[1][764] , \round_in[1][763] , \round_in[1][762] ,
         \round_in[1][761] , \round_in[1][760] , \round_in[1][759] ,
         \round_in[1][758] , \round_in[1][757] , \round_in[1][756] ,
         \round_in[1][755] , \round_in[1][754] , \round_in[1][753] ,
         \round_in[1][752] , \round_in[1][751] , \round_in[1][750] ,
         \round_in[1][749] , \round_in[1][748] , \round_in[1][747] ,
         \round_in[1][746] , \round_in[1][745] , \round_in[1][744] ,
         \round_in[1][743] , \round_in[1][742] , \round_in[1][741] ,
         \round_in[1][740] , \round_in[1][739] , \round_in[1][738] ,
         \round_in[1][737] , \round_in[1][736] , \round_in[1][735] ,
         \round_in[1][734] , \round_in[1][733] , \round_in[1][732] ,
         \round_in[1][731] , \round_in[1][730] , \round_in[1][729] ,
         \round_in[1][728] , \round_in[1][727] , \round_in[1][726] ,
         \round_in[1][725] , \round_in[1][724] , \round_in[1][723] ,
         \round_in[1][722] , \round_in[1][721] , \round_in[1][720] ,
         \round_in[1][719] , \round_in[1][718] , \round_in[1][717] ,
         \round_in[1][716] , \round_in[1][715] , \round_in[1][714] ,
         \round_in[1][713] , \round_in[1][712] , \round_in[1][711] ,
         \round_in[1][710] , \round_in[1][709] , \round_in[1][708] ,
         \round_in[1][707] , \round_in[1][706] , \round_in[1][705] ,
         \round_in[1][704] , \round_in[1][703] , \round_in[1][702] ,
         \round_in[1][701] , \round_in[1][700] , \round_in[1][699] ,
         \round_in[1][698] , \round_in[1][697] , \round_in[1][696] ,
         \round_in[1][695] , \round_in[1][694] , \round_in[1][693] ,
         \round_in[1][692] , \round_in[1][691] , \round_in[1][690] ,
         \round_in[1][689] , \round_in[1][688] , \round_in[1][687] ,
         \round_in[1][686] , \round_in[1][685] , \round_in[1][684] ,
         \round_in[1][683] , \round_in[1][682] , \round_in[1][681] ,
         \round_in[1][680] , \round_in[1][679] , \round_in[1][678] ,
         \round_in[1][677] , \round_in[1][676] , \round_in[1][675] ,
         \round_in[1][674] , \round_in[1][673] , \round_in[1][672] ,
         \round_in[1][671] , \round_in[1][670] , \round_in[1][669] ,
         \round_in[1][668] , \round_in[1][667] , \round_in[1][666] ,
         \round_in[1][665] , \round_in[1][664] , \round_in[1][663] ,
         \round_in[1][662] , \round_in[1][661] , \round_in[1][660] ,
         \round_in[1][659] , \round_in[1][658] , \round_in[1][657] ,
         \round_in[1][656] , \round_in[1][655] , \round_in[1][654] ,
         \round_in[1][653] , \round_in[1][652] , \round_in[1][651] ,
         \round_in[1][650] , \round_in[1][649] , \round_in[1][648] ,
         \round_in[1][647] , \round_in[1][646] , \round_in[1][645] ,
         \round_in[1][644] , \round_in[1][643] , \round_in[1][642] ,
         \round_in[1][641] , \round_in[1][640] , \round_in[1][639] ,
         \round_in[1][638] , \round_in[1][637] , \round_in[1][636] ,
         \round_in[1][635] , \round_in[1][634] , \round_in[1][633] ,
         \round_in[1][632] , \round_in[1][631] , \round_in[1][630] ,
         \round_in[1][629] , \round_in[1][628] , \round_in[1][627] ,
         \round_in[1][626] , \round_in[1][625] , \round_in[1][624] ,
         \round_in[1][623] , \round_in[1][622] , \round_in[1][621] ,
         \round_in[1][620] , \round_in[1][619] , \round_in[1][618] ,
         \round_in[1][617] , \round_in[1][616] , \round_in[1][615] ,
         \round_in[1][614] , \round_in[1][613] , \round_in[1][612] ,
         \round_in[1][611] , \round_in[1][610] , \round_in[1][609] ,
         \round_in[1][608] , \round_in[1][607] , \round_in[1][606] ,
         \round_in[1][605] , \round_in[1][604] , \round_in[1][603] ,
         \round_in[1][602] , \round_in[1][601] , \round_in[1][600] ,
         \round_in[1][599] , \round_in[1][598] , \round_in[1][597] ,
         \round_in[1][596] , \round_in[1][595] , \round_in[1][594] ,
         \round_in[1][593] , \round_in[1][592] , \round_in[1][591] ,
         \round_in[1][590] , \round_in[1][589] , \round_in[1][588] ,
         \round_in[1][587] , \round_in[1][586] , \round_in[1][585] ,
         \round_in[1][584] , \round_in[1][583] , \round_in[1][582] ,
         \round_in[1][581] , \round_in[1][580] , \round_in[1][579] ,
         \round_in[1][578] , \round_in[1][577] , \round_in[1][576] ,
         \round_in[1][575] , \round_in[1][574] , \round_in[1][573] ,
         \round_in[1][572] , \round_in[1][571] , \round_in[1][570] ,
         \round_in[1][569] , \round_in[1][568] , \round_in[1][567] ,
         \round_in[1][566] , \round_in[1][565] , \round_in[1][564] ,
         \round_in[1][563] , \round_in[1][562] , \round_in[1][561] ,
         \round_in[1][560] , \round_in[1][559] , \round_in[1][558] ,
         \round_in[1][557] , \round_in[1][556] , \round_in[1][555] ,
         \round_in[1][554] , \round_in[1][553] , \round_in[1][552] ,
         \round_in[1][551] , \round_in[1][550] , \round_in[1][549] ,
         \round_in[1][548] , \round_in[1][547] , \round_in[1][546] ,
         \round_in[1][545] , \round_in[1][544] , \round_in[1][543] ,
         \round_in[1][542] , \round_in[1][541] , \round_in[1][540] ,
         \round_in[1][539] , \round_in[1][538] , \round_in[1][537] ,
         \round_in[1][536] , \round_in[1][535] , \round_in[1][534] ,
         \round_in[1][533] , \round_in[1][532] , \round_in[1][531] ,
         \round_in[1][530] , \round_in[1][529] , \round_in[1][528] ,
         \round_in[1][527] , \round_in[1][526] , \round_in[1][525] ,
         \round_in[1][524] , \round_in[1][523] , \round_in[1][522] ,
         \round_in[1][521] , \round_in[1][520] , \round_in[1][519] ,
         \round_in[1][518] , \round_in[1][517] , \round_in[1][516] ,
         \round_in[1][515] , \round_in[1][514] , \round_in[1][513] ,
         \round_in[1][512] , \round_in[1][511] , \round_in[1][510] ,
         \round_in[1][509] , \round_in[1][508] , \round_in[1][507] ,
         \round_in[1][506] , \round_in[1][505] , \round_in[1][504] ,
         \round_in[1][503] , \round_in[1][502] , \round_in[1][501] ,
         \round_in[1][500] , \round_in[1][499] , \round_in[1][498] ,
         \round_in[1][497] , \round_in[1][496] , \round_in[1][495] ,
         \round_in[1][494] , \round_in[1][493] , \round_in[1][492] ,
         \round_in[1][491] , \round_in[1][490] , \round_in[1][489] ,
         \round_in[1][488] , \round_in[1][487] , \round_in[1][486] ,
         \round_in[1][485] , \round_in[1][484] , \round_in[1][483] ,
         \round_in[1][482] , \round_in[1][481] , \round_in[1][480] ,
         \round_in[1][479] , \round_in[1][478] , \round_in[1][477] ,
         \round_in[1][476] , \round_in[1][475] , \round_in[1][474] ,
         \round_in[1][473] , \round_in[1][472] , \round_in[1][471] ,
         \round_in[1][470] , \round_in[1][469] , \round_in[1][468] ,
         \round_in[1][467] , \round_in[1][466] , \round_in[1][465] ,
         \round_in[1][464] , \round_in[1][463] , \round_in[1][462] ,
         \round_in[1][461] , \round_in[1][460] , \round_in[1][459] ,
         \round_in[1][458] , \round_in[1][457] , \round_in[1][456] ,
         \round_in[1][455] , \round_in[1][454] , \round_in[1][453] ,
         \round_in[1][452] , \round_in[1][451] , \round_in[1][450] ,
         \round_in[1][449] , \round_in[1][448] , \round_in[1][447] ,
         \round_in[1][446] , \round_in[1][445] , \round_in[1][444] ,
         \round_in[1][443] , \round_in[1][442] , \round_in[1][441] ,
         \round_in[1][440] , \round_in[1][439] , \round_in[1][438] ,
         \round_in[1][437] , \round_in[1][436] , \round_in[1][435] ,
         \round_in[1][434] , \round_in[1][433] , \round_in[1][432] ,
         \round_in[1][431] , \round_in[1][430] , \round_in[1][429] ,
         \round_in[1][428] , \round_in[1][427] , \round_in[1][426] ,
         \round_in[1][425] , \round_in[1][424] , \round_in[1][423] ,
         \round_in[1][422] , \round_in[1][421] , \round_in[1][420] ,
         \round_in[1][419] , \round_in[1][418] , \round_in[1][417] ,
         \round_in[1][416] , \round_in[1][415] , \round_in[1][414] ,
         \round_in[1][413] , \round_in[1][412] , \round_in[1][411] ,
         \round_in[1][410] , \round_in[1][409] , \round_in[1][408] ,
         \round_in[1][407] , \round_in[1][406] , \round_in[1][405] ,
         \round_in[1][404] , \round_in[1][403] , \round_in[1][402] ,
         \round_in[1][401] , \round_in[1][400] , \round_in[1][399] ,
         \round_in[1][398] , \round_in[1][397] , \round_in[1][396] ,
         \round_in[1][395] , \round_in[1][394] , \round_in[1][393] ,
         \round_in[1][392] , \round_in[1][391] , \round_in[1][390] ,
         \round_in[1][389] , \round_in[1][388] , \round_in[1][387] ,
         \round_in[1][386] , \round_in[1][385] , \round_in[1][384] ,
         \round_in[1][383] , \round_in[1][382] , \round_in[1][381] ,
         \round_in[1][380] , \round_in[1][379] , \round_in[1][378] ,
         \round_in[1][377] , \round_in[1][376] , \round_in[1][375] ,
         \round_in[1][374] , \round_in[1][373] , \round_in[1][372] ,
         \round_in[1][371] , \round_in[1][370] , \round_in[1][369] ,
         \round_in[1][368] , \round_in[1][367] , \round_in[1][366] ,
         \round_in[1][365] , \round_in[1][364] , \round_in[1][363] ,
         \round_in[1][362] , \round_in[1][361] , \round_in[1][360] ,
         \round_in[1][359] , \round_in[1][358] , \round_in[1][357] ,
         \round_in[1][356] , \round_in[1][355] , \round_in[1][354] ,
         \round_in[1][353] , \round_in[1][352] , \round_in[1][351] ,
         \round_in[1][350] , \round_in[1][349] , \round_in[1][348] ,
         \round_in[1][347] , \round_in[1][346] , \round_in[1][345] ,
         \round_in[1][344] , \round_in[1][343] , \round_in[1][342] ,
         \round_in[1][341] , \round_in[1][340] , \round_in[1][339] ,
         \round_in[1][338] , \round_in[1][337] , \round_in[1][336] ,
         \round_in[1][335] , \round_in[1][334] , \round_in[1][333] ,
         \round_in[1][332] , \round_in[1][331] , \round_in[1][330] ,
         \round_in[1][329] , \round_in[1][328] , \round_in[1][327] ,
         \round_in[1][326] , \round_in[1][325] , \round_in[1][324] ,
         \round_in[1][323] , \round_in[1][322] , \round_in[1][321] ,
         \round_in[1][320] , \round_in[1][319] , \round_in[1][318] ,
         \round_in[1][317] , \round_in[1][316] , \round_in[1][315] ,
         \round_in[1][314] , \round_in[1][313] , \round_in[1][312] ,
         \round_in[1][311] , \round_in[1][310] , \round_in[1][309] ,
         \round_in[1][308] , \round_in[1][307] , \round_in[1][306] ,
         \round_in[1][305] , \round_in[1][304] , \round_in[1][303] ,
         \round_in[1][302] , \round_in[1][301] , \round_in[1][300] ,
         \round_in[1][299] , \round_in[1][298] , \round_in[1][297] ,
         \round_in[1][296] , \round_in[1][295] , \round_in[1][294] ,
         \round_in[1][293] , \round_in[1][292] , \round_in[1][291] ,
         \round_in[1][290] , \round_in[1][289] , \round_in[1][288] ,
         \round_in[1][287] , \round_in[1][286] , \round_in[1][285] ,
         \round_in[1][284] , \round_in[1][283] , \round_in[1][282] ,
         \round_in[1][281] , \round_in[1][280] , \round_in[1][279] ,
         \round_in[1][278] , \round_in[1][277] , \round_in[1][276] ,
         \round_in[1][275] , \round_in[1][274] , \round_in[1][273] ,
         \round_in[1][272] , \round_in[1][271] , \round_in[1][270] ,
         \round_in[1][269] , \round_in[1][268] , \round_in[1][267] ,
         \round_in[1][266] , \round_in[1][265] , \round_in[1][264] ,
         \round_in[1][263] , \round_in[1][262] , \round_in[1][261] ,
         \round_in[1][260] , \round_in[1][259] , \round_in[1][258] ,
         \round_in[1][257] , \round_in[1][256] , \round_in[1][255] ,
         \round_in[1][254] , \round_in[1][253] , \round_in[1][252] ,
         \round_in[1][251] , \round_in[1][250] , \round_in[1][249] ,
         \round_in[1][248] , \round_in[1][247] , \round_in[1][246] ,
         \round_in[1][245] , \round_in[1][244] , \round_in[1][243] ,
         \round_in[1][242] , \round_in[1][241] , \round_in[1][240] ,
         \round_in[1][239] , \round_in[1][238] , \round_in[1][237] ,
         \round_in[1][236] , \round_in[1][235] , \round_in[1][234] ,
         \round_in[1][233] , \round_in[1][232] , \round_in[1][231] ,
         \round_in[1][230] , \round_in[1][229] , \round_in[1][228] ,
         \round_in[1][227] , \round_in[1][226] , \round_in[1][225] ,
         \round_in[1][224] , \round_in[1][223] , \round_in[1][222] ,
         \round_in[1][221] , \round_in[1][220] , \round_in[1][219] ,
         \round_in[1][218] , \round_in[1][217] , \round_in[1][216] ,
         \round_in[1][215] , \round_in[1][214] , \round_in[1][213] ,
         \round_in[1][212] , \round_in[1][211] , \round_in[1][210] ,
         \round_in[1][209] , \round_in[1][208] , \round_in[1][207] ,
         \round_in[1][206] , \round_in[1][205] , \round_in[1][204] ,
         \round_in[1][203] , \round_in[1][202] , \round_in[1][201] ,
         \round_in[1][200] , \round_in[1][199] , \round_in[1][198] ,
         \round_in[1][197] , \round_in[1][196] , \round_in[1][195] ,
         \round_in[1][194] , \round_in[1][193] , \round_in[1][192] ,
         \round_in[1][191] , \round_in[1][190] , \round_in[1][189] ,
         \round_in[1][188] , \round_in[1][187] , \round_in[1][186] ,
         \round_in[1][185] , \round_in[1][184] , \round_in[1][183] ,
         \round_in[1][182] , \round_in[1][181] , \round_in[1][180] ,
         \round_in[1][179] , \round_in[1][178] , \round_in[1][177] ,
         \round_in[1][176] , \round_in[1][175] , \round_in[1][174] ,
         \round_in[1][173] , \round_in[1][172] , \round_in[1][171] ,
         \round_in[1][170] , \round_in[1][169] , \round_in[1][168] ,
         \round_in[1][167] , \round_in[1][166] , \round_in[1][165] ,
         \round_in[1][164] , \round_in[1][163] , \round_in[1][162] ,
         \round_in[1][161] , \round_in[1][160] , \round_in[1][159] ,
         \round_in[1][158] , \round_in[1][157] , \round_in[1][156] ,
         \round_in[1][155] , \round_in[1][154] , \round_in[1][153] ,
         \round_in[1][152] , \round_in[1][151] , \round_in[1][150] ,
         \round_in[1][149] , \round_in[1][148] , \round_in[1][147] ,
         \round_in[1][146] , \round_in[1][145] , \round_in[1][144] ,
         \round_in[1][143] , \round_in[1][142] , \round_in[1][141] ,
         \round_in[1][140] , \round_in[1][139] , \round_in[1][138] ,
         \round_in[1][137] , \round_in[1][136] , \round_in[1][135] ,
         \round_in[1][134] , \round_in[1][133] , \round_in[1][132] ,
         \round_in[1][131] , \round_in[1][130] , \round_in[1][129] ,
         \round_in[1][128] , \round_in[1][127] , \round_in[1][126] ,
         \round_in[1][125] , \round_in[1][124] , \round_in[1][123] ,
         \round_in[1][122] , \round_in[1][121] , \round_in[1][120] ,
         \round_in[1][119] , \round_in[1][118] , \round_in[1][117] ,
         \round_in[1][116] , \round_in[1][115] , \round_in[1][114] ,
         \round_in[1][113] , \round_in[1][112] , \round_in[1][111] ,
         \round_in[1][110] , \round_in[1][109] , \round_in[1][108] ,
         \round_in[1][107] , \round_in[1][106] , \round_in[1][105] ,
         \round_in[1][104] , \round_in[1][103] , \round_in[1][102] ,
         \round_in[1][101] , \round_in[1][100] , \round_in[1][99] ,
         \round_in[1][98] , \round_in[1][97] , \round_in[1][96] ,
         \round_in[1][95] , \round_in[1][94] , \round_in[1][93] ,
         \round_in[1][92] , \round_in[1][91] , \round_in[1][90] ,
         \round_in[1][89] , \round_in[1][88] , \round_in[1][87] ,
         \round_in[1][86] , \round_in[1][85] , \round_in[1][84] ,
         \round_in[1][83] , \round_in[1][82] , \round_in[1][81] ,
         \round_in[1][80] , \round_in[1][79] , \round_in[1][78] ,
         \round_in[1][77] , \round_in[1][76] , \round_in[1][75] ,
         \round_in[1][74] , \round_in[1][73] , \round_in[1][72] ,
         \round_in[1][71] , \round_in[1][70] , \round_in[1][69] ,
         \round_in[1][68] , \round_in[1][67] , \round_in[1][66] ,
         \round_in[1][65] , \round_in[1][64] , \round_in[1][63] ,
         \round_in[1][62] , \round_in[1][61] , \round_in[1][60] ,
         \round_in[1][59] , \round_in[1][58] , \round_in[1][57] ,
         \round_in[1][56] , \round_in[1][55] , \round_in[1][54] ,
         \round_in[1][53] , \round_in[1][52] , \round_in[1][51] ,
         \round_in[1][50] , \round_in[1][49] , \round_in[1][48] ,
         \round_in[1][47] , \round_in[1][46] , \round_in[1][45] ,
         \round_in[1][44] , \round_in[1][43] , \round_in[1][42] ,
         \round_in[1][41] , \round_in[1][40] , \round_in[1][39] ,
         \round_in[1][38] , \round_in[1][37] , \round_in[1][36] ,
         \round_in[1][35] , \round_in[1][34] , \round_in[1][33] ,
         \round_in[1][32] , \round_in[1][31] , \round_in[1][30] ,
         \round_in[1][29] , \round_in[1][28] , \round_in[1][27] ,
         \round_in[1][26] , \round_in[1][25] , \round_in[1][24] ,
         \round_in[1][23] , \round_in[1][22] , \round_in[1][21] ,
         \round_in[1][20] , \round_in[1][19] , \round_in[1][18] ,
         \round_in[1][17] , \round_in[1][16] , \round_in[1][15] ,
         \round_in[1][14] , \round_in[1][13] , \round_in[1][12] ,
         \round_in[1][11] , \round_in[1][10] , \round_in[1][9] ,
         \round_in[1][8] , \round_in[1][7] , \round_in[1][6] ,
         \round_in[1][5] , \round_in[1][4] , \round_in[1][3] ,
         \round_in[1][2] , \round_in[1][1] , \round_in[1][0] ,
         \round_in[0][1599] , \round_in[0][1598] , \round_in[0][1597] ,
         \round_in[0][1596] , \round_in[0][1595] , \round_in[0][1594] ,
         \round_in[0][1593] , \round_in[0][1592] , \round_in[0][1591] ,
         \round_in[0][1590] , \round_in[0][1589] , \round_in[0][1588] ,
         \round_in[0][1587] , \round_in[0][1586] , \round_in[0][1585] ,
         \round_in[0][1584] , \round_in[0][1583] , \round_in[0][1582] ,
         \round_in[0][1581] , \round_in[0][1580] , \round_in[0][1579] ,
         \round_in[0][1578] , \round_in[0][1577] , \round_in[0][1576] ,
         \round_in[0][1575] , \round_in[0][1574] , \round_in[0][1573] ,
         \round_in[0][1572] , \round_in[0][1571] , \round_in[0][1570] ,
         \round_in[0][1569] , \round_in[0][1568] , \round_in[0][1567] ,
         \round_in[0][1566] , \round_in[0][1565] , \round_in[0][1564] ,
         \round_in[0][1563] , \round_in[0][1562] , \round_in[0][1561] ,
         \round_in[0][1560] , \round_in[0][1559] , \round_in[0][1558] ,
         \round_in[0][1557] , \round_in[0][1556] , \round_in[0][1555] ,
         \round_in[0][1554] , \round_in[0][1553] , \round_in[0][1552] ,
         \round_in[0][1551] , \round_in[0][1550] , \round_in[0][1549] ,
         \round_in[0][1548] , \round_in[0][1547] , \round_in[0][1546] ,
         \round_in[0][1545] , \round_in[0][1544] , \round_in[0][1543] ,
         \round_in[0][1542] , \round_in[0][1541] , \round_in[0][1540] ,
         \round_in[0][1539] , \round_in[0][1538] , \round_in[0][1537] ,
         \round_in[0][1536] , \round_in[0][1535] , \round_in[0][1534] ,
         \round_in[0][1533] , \round_in[0][1532] , \round_in[0][1531] ,
         \round_in[0][1530] , \round_in[0][1529] , \round_in[0][1528] ,
         \round_in[0][1527] , \round_in[0][1526] , \round_in[0][1525] ,
         \round_in[0][1524] , \round_in[0][1523] , \round_in[0][1522] ,
         \round_in[0][1521] , \round_in[0][1520] , \round_in[0][1519] ,
         \round_in[0][1518] , \round_in[0][1517] , \round_in[0][1516] ,
         \round_in[0][1515] , \round_in[0][1514] , \round_in[0][1513] ,
         \round_in[0][1512] , \round_in[0][1511] , \round_in[0][1510] ,
         \round_in[0][1509] , \round_in[0][1508] , \round_in[0][1507] ,
         \round_in[0][1506] , \round_in[0][1505] , \round_in[0][1504] ,
         \round_in[0][1503] , \round_in[0][1502] , \round_in[0][1501] ,
         \round_in[0][1500] , \round_in[0][1499] , \round_in[0][1498] ,
         \round_in[0][1497] , \round_in[0][1496] , \round_in[0][1495] ,
         \round_in[0][1494] , \round_in[0][1493] , \round_in[0][1492] ,
         \round_in[0][1491] , \round_in[0][1490] , \round_in[0][1489] ,
         \round_in[0][1488] , \round_in[0][1487] , \round_in[0][1486] ,
         \round_in[0][1485] , \round_in[0][1484] , \round_in[0][1483] ,
         \round_in[0][1482] , \round_in[0][1481] , \round_in[0][1480] ,
         \round_in[0][1479] , \round_in[0][1478] , \round_in[0][1477] ,
         \round_in[0][1476] , \round_in[0][1475] , \round_in[0][1474] ,
         \round_in[0][1473] , \round_in[0][1472] , \round_in[0][1471] ,
         \round_in[0][1470] , \round_in[0][1469] , \round_in[0][1468] ,
         \round_in[0][1467] , \round_in[0][1466] , \round_in[0][1465] ,
         \round_in[0][1464] , \round_in[0][1463] , \round_in[0][1462] ,
         \round_in[0][1461] , \round_in[0][1460] , \round_in[0][1459] ,
         \round_in[0][1458] , \round_in[0][1457] , \round_in[0][1456] ,
         \round_in[0][1455] , \round_in[0][1454] , \round_in[0][1453] ,
         \round_in[0][1452] , \round_in[0][1451] , \round_in[0][1450] ,
         \round_in[0][1449] , \round_in[0][1448] , \round_in[0][1447] ,
         \round_in[0][1446] , \round_in[0][1445] , \round_in[0][1444] ,
         \round_in[0][1443] , \round_in[0][1442] , \round_in[0][1441] ,
         \round_in[0][1440] , \round_in[0][1439] , \round_in[0][1438] ,
         \round_in[0][1437] , \round_in[0][1436] , \round_in[0][1435] ,
         \round_in[0][1434] , \round_in[0][1433] , \round_in[0][1432] ,
         \round_in[0][1431] , \round_in[0][1430] , \round_in[0][1429] ,
         \round_in[0][1428] , \round_in[0][1427] , \round_in[0][1426] ,
         \round_in[0][1425] , \round_in[0][1424] , \round_in[0][1423] ,
         \round_in[0][1422] , \round_in[0][1421] , \round_in[0][1420] ,
         \round_in[0][1419] , \round_in[0][1418] , \round_in[0][1417] ,
         \round_in[0][1416] , \round_in[0][1415] , \round_in[0][1414] ,
         \round_in[0][1413] , \round_in[0][1412] , \round_in[0][1411] ,
         \round_in[0][1410] , \round_in[0][1409] , \round_in[0][1408] ,
         \round_in[0][1407] , \round_in[0][1406] , \round_in[0][1405] ,
         \round_in[0][1404] , \round_in[0][1403] , \round_in[0][1402] ,
         \round_in[0][1401] , \round_in[0][1400] , \round_in[0][1399] ,
         \round_in[0][1398] , \round_in[0][1397] , \round_in[0][1396] ,
         \round_in[0][1395] , \round_in[0][1394] , \round_in[0][1393] ,
         \round_in[0][1392] , \round_in[0][1391] , \round_in[0][1390] ,
         \round_in[0][1389] , \round_in[0][1388] , \round_in[0][1387] ,
         \round_in[0][1386] , \round_in[0][1385] , \round_in[0][1384] ,
         \round_in[0][1383] , \round_in[0][1382] , \round_in[0][1381] ,
         \round_in[0][1380] , \round_in[0][1379] , \round_in[0][1378] ,
         \round_in[0][1377] , \round_in[0][1376] , \round_in[0][1375] ,
         \round_in[0][1374] , \round_in[0][1373] , \round_in[0][1372] ,
         \round_in[0][1371] , \round_in[0][1370] , \round_in[0][1369] ,
         \round_in[0][1368] , \round_in[0][1367] , \round_in[0][1366] ,
         \round_in[0][1365] , \round_in[0][1364] , \round_in[0][1363] ,
         \round_in[0][1362] , \round_in[0][1361] , \round_in[0][1360] ,
         \round_in[0][1359] , \round_in[0][1358] , \round_in[0][1357] ,
         \round_in[0][1356] , \round_in[0][1355] , \round_in[0][1354] ,
         \round_in[0][1353] , \round_in[0][1352] , \round_in[0][1351] ,
         \round_in[0][1350] , \round_in[0][1349] , \round_in[0][1348] ,
         \round_in[0][1347] , \round_in[0][1346] , \round_in[0][1345] ,
         \round_in[0][1344] , \round_in[0][1343] , \round_in[0][1342] ,
         \round_in[0][1341] , \round_in[0][1340] , \round_in[0][1339] ,
         \round_in[0][1338] , \round_in[0][1337] , \round_in[0][1336] ,
         \round_in[0][1335] , \round_in[0][1334] , \round_in[0][1333] ,
         \round_in[0][1332] , \round_in[0][1331] , \round_in[0][1330] ,
         \round_in[0][1329] , \round_in[0][1328] , \round_in[0][1327] ,
         \round_in[0][1326] , \round_in[0][1325] , \round_in[0][1324] ,
         \round_in[0][1323] , \round_in[0][1322] , \round_in[0][1321] ,
         \round_in[0][1320] , \round_in[0][1319] , \round_in[0][1318] ,
         \round_in[0][1317] , \round_in[0][1316] , \round_in[0][1315] ,
         \round_in[0][1314] , \round_in[0][1313] , \round_in[0][1312] ,
         \round_in[0][1311] , \round_in[0][1310] , \round_in[0][1309] ,
         \round_in[0][1308] , \round_in[0][1307] , \round_in[0][1306] ,
         \round_in[0][1305] , \round_in[0][1304] , \round_in[0][1303] ,
         \round_in[0][1302] , \round_in[0][1301] , \round_in[0][1300] ,
         \round_in[0][1299] , \round_in[0][1298] , \round_in[0][1297] ,
         \round_in[0][1296] , \round_in[0][1295] , \round_in[0][1294] ,
         \round_in[0][1293] , \round_in[0][1292] , \round_in[0][1291] ,
         \round_in[0][1290] , \round_in[0][1289] , \round_in[0][1288] ,
         \round_in[0][1287] , \round_in[0][1286] , \round_in[0][1285] ,
         \round_in[0][1284] , \round_in[0][1283] , \round_in[0][1282] ,
         \round_in[0][1281] , \round_in[0][1280] , \round_in[0][1279] ,
         \round_in[0][1278] , \round_in[0][1277] , \round_in[0][1276] ,
         \round_in[0][1275] , \round_in[0][1274] , \round_in[0][1273] ,
         \round_in[0][1272] , \round_in[0][1271] , \round_in[0][1270] ,
         \round_in[0][1269] , \round_in[0][1268] , \round_in[0][1267] ,
         \round_in[0][1266] , \round_in[0][1265] , \round_in[0][1264] ,
         \round_in[0][1263] , \round_in[0][1262] , \round_in[0][1261] ,
         \round_in[0][1260] , \round_in[0][1259] , \round_in[0][1258] ,
         \round_in[0][1257] , \round_in[0][1256] , \round_in[0][1255] ,
         \round_in[0][1254] , \round_in[0][1253] , \round_in[0][1252] ,
         \round_in[0][1251] , \round_in[0][1250] , \round_in[0][1249] ,
         \round_in[0][1248] , \round_in[0][1247] , \round_in[0][1246] ,
         \round_in[0][1245] , \round_in[0][1244] , \round_in[0][1243] ,
         \round_in[0][1242] , \round_in[0][1241] , \round_in[0][1240] ,
         \round_in[0][1239] , \round_in[0][1238] , \round_in[0][1237] ,
         \round_in[0][1236] , \round_in[0][1235] , \round_in[0][1234] ,
         \round_in[0][1233] , \round_in[0][1232] , \round_in[0][1231] ,
         \round_in[0][1230] , \round_in[0][1229] , \round_in[0][1228] ,
         \round_in[0][1227] , \round_in[0][1226] , \round_in[0][1225] ,
         \round_in[0][1224] , \round_in[0][1223] , \round_in[0][1222] ,
         \round_in[0][1221] , \round_in[0][1220] , \round_in[0][1219] ,
         \round_in[0][1218] , \round_in[0][1217] , \round_in[0][1216] ,
         \round_in[0][1215] , \round_in[0][1214] , \round_in[0][1213] ,
         \round_in[0][1212] , \round_in[0][1211] , \round_in[0][1210] ,
         \round_in[0][1209] , \round_in[0][1208] , \round_in[0][1207] ,
         \round_in[0][1206] , \round_in[0][1205] , \round_in[0][1204] ,
         \round_in[0][1203] , \round_in[0][1202] , \round_in[0][1201] ,
         \round_in[0][1200] , \round_in[0][1199] , \round_in[0][1198] ,
         \round_in[0][1197] , \round_in[0][1196] , \round_in[0][1195] ,
         \round_in[0][1194] , \round_in[0][1193] , \round_in[0][1192] ,
         \round_in[0][1191] , \round_in[0][1190] , \round_in[0][1189] ,
         \round_in[0][1188] , \round_in[0][1187] , \round_in[0][1186] ,
         \round_in[0][1185] , \round_in[0][1184] , \round_in[0][1183] ,
         \round_in[0][1182] , \round_in[0][1181] , \round_in[0][1180] ,
         \round_in[0][1179] , \round_in[0][1178] , \round_in[0][1177] ,
         \round_in[0][1176] , \round_in[0][1175] , \round_in[0][1174] ,
         \round_in[0][1173] , \round_in[0][1172] , \round_in[0][1171] ,
         \round_in[0][1170] , \round_in[0][1169] , \round_in[0][1168] ,
         \round_in[0][1167] , \round_in[0][1166] , \round_in[0][1165] ,
         \round_in[0][1164] , \round_in[0][1163] , \round_in[0][1162] ,
         \round_in[0][1161] , \round_in[0][1160] , \round_in[0][1159] ,
         \round_in[0][1158] , \round_in[0][1157] , \round_in[0][1156] ,
         \round_in[0][1155] , \round_in[0][1154] , \round_in[0][1153] ,
         \round_in[0][1152] , \round_in[0][1151] , \round_in[0][1150] ,
         \round_in[0][1149] , \round_in[0][1148] , \round_in[0][1147] ,
         \round_in[0][1146] , \round_in[0][1145] , \round_in[0][1144] ,
         \round_in[0][1143] , \round_in[0][1142] , \round_in[0][1141] ,
         \round_in[0][1140] , \round_in[0][1139] , \round_in[0][1138] ,
         \round_in[0][1137] , \round_in[0][1136] , \round_in[0][1135] ,
         \round_in[0][1134] , \round_in[0][1133] , \round_in[0][1132] ,
         \round_in[0][1131] , \round_in[0][1130] , \round_in[0][1129] ,
         \round_in[0][1128] , \round_in[0][1127] , \round_in[0][1126] ,
         \round_in[0][1125] , \round_in[0][1124] , \round_in[0][1123] ,
         \round_in[0][1122] , \round_in[0][1121] , \round_in[0][1120] ,
         \round_in[0][1119] , \round_in[0][1118] , \round_in[0][1117] ,
         \round_in[0][1116] , \round_in[0][1115] , \round_in[0][1114] ,
         \round_in[0][1113] , \round_in[0][1112] , \round_in[0][1111] ,
         \round_in[0][1110] , \round_in[0][1109] , \round_in[0][1108] ,
         \round_in[0][1107] , \round_in[0][1106] , \round_in[0][1105] ,
         \round_in[0][1104] , \round_in[0][1103] , \round_in[0][1102] ,
         \round_in[0][1101] , \round_in[0][1100] , \round_in[0][1099] ,
         \round_in[0][1098] , \round_in[0][1097] , \round_in[0][1096] ,
         \round_in[0][1095] , \round_in[0][1094] , \round_in[0][1093] ,
         \round_in[0][1092] , \round_in[0][1091] , \round_in[0][1090] ,
         \round_in[0][1089] , \round_in[0][1088] , \round_in[0][1087] ,
         \round_in[0][1086] , \round_in[0][1085] , \round_in[0][1084] ,
         \round_in[0][1083] , \round_in[0][1082] , \round_in[0][1081] ,
         \round_in[0][1080] , \round_in[0][1079] , \round_in[0][1078] ,
         \round_in[0][1077] , \round_in[0][1076] , \round_in[0][1075] ,
         \round_in[0][1074] , \round_in[0][1073] , \round_in[0][1072] ,
         \round_in[0][1071] , \round_in[0][1070] , \round_in[0][1069] ,
         \round_in[0][1068] , \round_in[0][1067] , \round_in[0][1066] ,
         \round_in[0][1065] , \round_in[0][1064] , \round_in[0][1063] ,
         \round_in[0][1062] , \round_in[0][1061] , \round_in[0][1060] ,
         \round_in[0][1059] , \round_in[0][1058] , \round_in[0][1057] ,
         \round_in[0][1056] , \round_in[0][1055] , \round_in[0][1054] ,
         \round_in[0][1053] , \round_in[0][1052] , \round_in[0][1051] ,
         \round_in[0][1050] , \round_in[0][1049] , \round_in[0][1048] ,
         \round_in[0][1047] , \round_in[0][1046] , \round_in[0][1045] ,
         \round_in[0][1044] , \round_in[0][1043] , \round_in[0][1042] ,
         \round_in[0][1041] , \round_in[0][1040] , \round_in[0][1039] ,
         \round_in[0][1038] , \round_in[0][1037] , \round_in[0][1036] ,
         \round_in[0][1035] , \round_in[0][1034] , \round_in[0][1033] ,
         \round_in[0][1032] , \round_in[0][1031] , \round_in[0][1030] ,
         \round_in[0][1029] , \round_in[0][1028] , \round_in[0][1027] ,
         \round_in[0][1026] , \round_in[0][1025] , \round_in[0][1024] ,
         \round_in[0][1023] , \round_in[0][1022] , \round_in[0][1021] ,
         \round_in[0][1020] , \round_in[0][1019] , \round_in[0][1018] ,
         \round_in[0][1017] , \round_in[0][1016] , \round_in[0][1015] ,
         \round_in[0][1014] , \round_in[0][1013] , \round_in[0][1012] ,
         \round_in[0][1011] , \round_in[0][1010] , \round_in[0][1009] ,
         \round_in[0][1008] , \round_in[0][1007] , \round_in[0][1006] ,
         \round_in[0][1005] , \round_in[0][1004] , \round_in[0][1003] ,
         \round_in[0][1002] , \round_in[0][1001] , \round_in[0][1000] ,
         \round_in[0][999] , \round_in[0][998] , \round_in[0][997] ,
         \round_in[0][996] , \round_in[0][995] , \round_in[0][994] ,
         \round_in[0][993] , \round_in[0][992] , \round_in[0][991] ,
         \round_in[0][990] , \round_in[0][989] , \round_in[0][988] ,
         \round_in[0][987] , \round_in[0][986] , \round_in[0][985] ,
         \round_in[0][984] , \round_in[0][983] , \round_in[0][982] ,
         \round_in[0][981] , \round_in[0][980] , \round_in[0][979] ,
         \round_in[0][978] , \round_in[0][977] , \round_in[0][976] ,
         \round_in[0][975] , \round_in[0][974] , \round_in[0][973] ,
         \round_in[0][972] , \round_in[0][971] , \round_in[0][970] ,
         \round_in[0][969] , \round_in[0][968] , \round_in[0][967] ,
         \round_in[0][966] , \round_in[0][965] , \round_in[0][964] ,
         \round_in[0][963] , \round_in[0][962] , \round_in[0][961] ,
         \round_in[0][960] , \round_in[0][959] , \round_in[0][958] ,
         \round_in[0][957] , \round_in[0][956] , \round_in[0][955] ,
         \round_in[0][954] , \round_in[0][953] , \round_in[0][952] ,
         \round_in[0][951] , \round_in[0][950] , \round_in[0][949] ,
         \round_in[0][948] , \round_in[0][947] , \round_in[0][946] ,
         \round_in[0][945] , \round_in[0][944] , \round_in[0][943] ,
         \round_in[0][942] , \round_in[0][941] , \round_in[0][940] ,
         \round_in[0][939] , \round_in[0][938] , \round_in[0][937] ,
         \round_in[0][936] , \round_in[0][935] , \round_in[0][934] ,
         \round_in[0][933] , \round_in[0][932] , \round_in[0][931] ,
         \round_in[0][930] , \round_in[0][929] , \round_in[0][928] ,
         \round_in[0][927] , \round_in[0][926] , \round_in[0][925] ,
         \round_in[0][924] , \round_in[0][923] , \round_in[0][922] ,
         \round_in[0][921] , \round_in[0][920] , \round_in[0][919] ,
         \round_in[0][918] , \round_in[0][917] , \round_in[0][916] ,
         \round_in[0][915] , \round_in[0][914] , \round_in[0][913] ,
         \round_in[0][912] , \round_in[0][911] , \round_in[0][910] ,
         \round_in[0][909] , \round_in[0][908] , \round_in[0][907] ,
         \round_in[0][906] , \round_in[0][905] , \round_in[0][904] ,
         \round_in[0][903] , \round_in[0][902] , \round_in[0][901] ,
         \round_in[0][900] , \round_in[0][899] , \round_in[0][898] ,
         \round_in[0][897] , \round_in[0][896] , \round_in[0][895] ,
         \round_in[0][894] , \round_in[0][893] , \round_in[0][892] ,
         \round_in[0][891] , \round_in[0][890] , \round_in[0][889] ,
         \round_in[0][888] , \round_in[0][887] , \round_in[0][886] ,
         \round_in[0][885] , \round_in[0][884] , \round_in[0][883] ,
         \round_in[0][882] , \round_in[0][881] , \round_in[0][880] ,
         \round_in[0][879] , \round_in[0][878] , \round_in[0][877] ,
         \round_in[0][876] , \round_in[0][875] , \round_in[0][874] ,
         \round_in[0][873] , \round_in[0][872] , \round_in[0][871] ,
         \round_in[0][870] , \round_in[0][869] , \round_in[0][868] ,
         \round_in[0][867] , \round_in[0][866] , \round_in[0][865] ,
         \round_in[0][864] , \round_in[0][863] , \round_in[0][862] ,
         \round_in[0][861] , \round_in[0][860] , \round_in[0][859] ,
         \round_in[0][858] , \round_in[0][857] , \round_in[0][856] ,
         \round_in[0][855] , \round_in[0][854] , \round_in[0][853] ,
         \round_in[0][852] , \round_in[0][851] , \round_in[0][850] ,
         \round_in[0][849] , \round_in[0][848] , \round_in[0][847] ,
         \round_in[0][846] , \round_in[0][845] , \round_in[0][844] ,
         \round_in[0][843] , \round_in[0][842] , \round_in[0][841] ,
         \round_in[0][840] , \round_in[0][839] , \round_in[0][838] ,
         \round_in[0][837] , \round_in[0][836] , \round_in[0][835] ,
         \round_in[0][834] , \round_in[0][833] , \round_in[0][832] ,
         \round_in[0][831] , \round_in[0][830] , \round_in[0][829] ,
         \round_in[0][828] , \round_in[0][827] , \round_in[0][826] ,
         \round_in[0][825] , \round_in[0][824] , \round_in[0][823] ,
         \round_in[0][822] , \round_in[0][821] , \round_in[0][820] ,
         \round_in[0][819] , \round_in[0][818] , \round_in[0][817] ,
         \round_in[0][816] , \round_in[0][815] , \round_in[0][814] ,
         \round_in[0][813] , \round_in[0][812] , \round_in[0][811] ,
         \round_in[0][810] , \round_in[0][809] , \round_in[0][808] ,
         \round_in[0][807] , \round_in[0][806] , \round_in[0][805] ,
         \round_in[0][804] , \round_in[0][803] , \round_in[0][802] ,
         \round_in[0][801] , \round_in[0][800] , \round_in[0][799] ,
         \round_in[0][798] , \round_in[0][797] , \round_in[0][796] ,
         \round_in[0][795] , \round_in[0][794] , \round_in[0][793] ,
         \round_in[0][792] , \round_in[0][791] , \round_in[0][790] ,
         \round_in[0][789] , \round_in[0][788] , \round_in[0][787] ,
         \round_in[0][786] , \round_in[0][785] , \round_in[0][784] ,
         \round_in[0][783] , \round_in[0][782] , \round_in[0][781] ,
         \round_in[0][780] , \round_in[0][779] , \round_in[0][778] ,
         \round_in[0][777] , \round_in[0][776] , \round_in[0][775] ,
         \round_in[0][774] , \round_in[0][773] , \round_in[0][772] ,
         \round_in[0][771] , \round_in[0][770] , \round_in[0][769] ,
         \round_in[0][768] , \round_in[0][767] , \round_in[0][766] ,
         \round_in[0][765] , \round_in[0][764] , \round_in[0][763] ,
         \round_in[0][762] , \round_in[0][761] , \round_in[0][760] ,
         \round_in[0][759] , \round_in[0][758] , \round_in[0][757] ,
         \round_in[0][756] , \round_in[0][755] , \round_in[0][754] ,
         \round_in[0][753] , \round_in[0][752] , \round_in[0][751] ,
         \round_in[0][750] , \round_in[0][749] , \round_in[0][748] ,
         \round_in[0][747] , \round_in[0][746] , \round_in[0][745] ,
         \round_in[0][744] , \round_in[0][743] , \round_in[0][742] ,
         \round_in[0][741] , \round_in[0][740] , \round_in[0][739] ,
         \round_in[0][738] , \round_in[0][737] , \round_in[0][736] ,
         \round_in[0][735] , \round_in[0][734] , \round_in[0][733] ,
         \round_in[0][732] , \round_in[0][731] , \round_in[0][730] ,
         \round_in[0][729] , \round_in[0][728] , \round_in[0][727] ,
         \round_in[0][726] , \round_in[0][725] , \round_in[0][724] ,
         \round_in[0][723] , \round_in[0][722] , \round_in[0][721] ,
         \round_in[0][720] , \round_in[0][719] , \round_in[0][718] ,
         \round_in[0][717] , \round_in[0][716] , \round_in[0][715] ,
         \round_in[0][714] , \round_in[0][713] , \round_in[0][712] ,
         \round_in[0][711] , \round_in[0][710] , \round_in[0][709] ,
         \round_in[0][708] , \round_in[0][707] , \round_in[0][706] ,
         \round_in[0][705] , \round_in[0][704] , \round_in[0][703] ,
         \round_in[0][702] , \round_in[0][701] , \round_in[0][700] ,
         \round_in[0][699] , \round_in[0][698] , \round_in[0][697] ,
         \round_in[0][696] , \round_in[0][695] , \round_in[0][694] ,
         \round_in[0][693] , \round_in[0][692] , \round_in[0][691] ,
         \round_in[0][690] , \round_in[0][689] , \round_in[0][688] ,
         \round_in[0][687] , \round_in[0][686] , \round_in[0][685] ,
         \round_in[0][684] , \round_in[0][683] , \round_in[0][682] ,
         \round_in[0][681] , \round_in[0][680] , \round_in[0][679] ,
         \round_in[0][678] , \round_in[0][677] , \round_in[0][676] ,
         \round_in[0][675] , \round_in[0][674] , \round_in[0][673] ,
         \round_in[0][672] , \round_in[0][671] , \round_in[0][670] ,
         \round_in[0][669] , \round_in[0][668] , \round_in[0][667] ,
         \round_in[0][666] , \round_in[0][665] , \round_in[0][664] ,
         \round_in[0][663] , \round_in[0][662] , \round_in[0][661] ,
         \round_in[0][660] , \round_in[0][659] , \round_in[0][658] ,
         \round_in[0][657] , \round_in[0][656] , \round_in[0][655] ,
         \round_in[0][654] , \round_in[0][653] , \round_in[0][652] ,
         \round_in[0][651] , \round_in[0][650] , \round_in[0][649] ,
         \round_in[0][648] , \round_in[0][647] , \round_in[0][646] ,
         \round_in[0][645] , \round_in[0][644] , \round_in[0][643] ,
         \round_in[0][642] , \round_in[0][641] , \round_in[0][640] ,
         \round_in[0][639] , \round_in[0][638] , \round_in[0][637] ,
         \round_in[0][636] , \round_in[0][635] , \round_in[0][634] ,
         \round_in[0][633] , \round_in[0][632] , \round_in[0][631] ,
         \round_in[0][630] , \round_in[0][629] , \round_in[0][628] ,
         \round_in[0][627] , \round_in[0][626] , \round_in[0][625] ,
         \round_in[0][624] , \round_in[0][623] , \round_in[0][622] ,
         \round_in[0][621] , \round_in[0][620] , \round_in[0][619] ,
         \round_in[0][618] , \round_in[0][617] , \round_in[0][616] ,
         \round_in[0][615] , \round_in[0][614] , \round_in[0][613] ,
         \round_in[0][612] , \round_in[0][611] , \round_in[0][610] ,
         \round_in[0][609] , \round_in[0][608] , \round_in[0][607] ,
         \round_in[0][606] , \round_in[0][605] , \round_in[0][604] ,
         \round_in[0][603] , \round_in[0][602] , \round_in[0][601] ,
         \round_in[0][600] , \round_in[0][599] , \round_in[0][598] ,
         \round_in[0][597] , \round_in[0][596] , \round_in[0][595] ,
         \round_in[0][594] , \round_in[0][593] , \round_in[0][592] ,
         \round_in[0][591] , \round_in[0][590] , \round_in[0][589] ,
         \round_in[0][588] , \round_in[0][587] , \round_in[0][586] ,
         \round_in[0][585] , \round_in[0][584] , \round_in[0][583] ,
         \round_in[0][582] , \round_in[0][581] , \round_in[0][580] ,
         \round_in[0][579] , \round_in[0][578] , \round_in[0][577] ,
         \round_in[0][576] , \round_in[0][575] , \round_in[0][574] ,
         \round_in[0][573] , \round_in[0][572] , \round_in[0][571] ,
         \round_in[0][570] , \round_in[0][569] , \round_in[0][568] ,
         \round_in[0][567] , \round_in[0][566] , \round_in[0][565] ,
         \round_in[0][564] , \round_in[0][563] , \round_in[0][562] ,
         \round_in[0][561] , \round_in[0][560] , \round_in[0][559] ,
         \round_in[0][558] , \round_in[0][557] , \round_in[0][556] ,
         \round_in[0][555] , \round_in[0][554] , \round_in[0][553] ,
         \round_in[0][552] , \round_in[0][551] , \round_in[0][550] ,
         \round_in[0][549] , \round_in[0][548] , \round_in[0][547] ,
         \round_in[0][546] , \round_in[0][545] , \round_in[0][544] ,
         \round_in[0][543] , \round_in[0][542] , \round_in[0][541] ,
         \round_in[0][540] , \round_in[0][539] , \round_in[0][538] ,
         \round_in[0][537] , \round_in[0][536] , \round_in[0][535] ,
         \round_in[0][534] , \round_in[0][533] , \round_in[0][532] ,
         \round_in[0][531] , \round_in[0][530] , \round_in[0][529] ,
         \round_in[0][528] , \round_in[0][527] , \round_in[0][526] ,
         \round_in[0][525] , \round_in[0][524] , \round_in[0][523] ,
         \round_in[0][522] , \round_in[0][521] , \round_in[0][520] ,
         \round_in[0][519] , \round_in[0][518] , \round_in[0][517] ,
         \round_in[0][516] , \round_in[0][515] , \round_in[0][514] ,
         \round_in[0][513] , \round_in[0][512] , \round_in[0][511] ,
         \round_in[0][510] , \round_in[0][509] , \round_in[0][508] ,
         \round_in[0][507] , \round_in[0][506] , \round_in[0][505] ,
         \round_in[0][504] , \round_in[0][503] , \round_in[0][502] ,
         \round_in[0][501] , \round_in[0][500] , \round_in[0][499] ,
         \round_in[0][498] , \round_in[0][497] , \round_in[0][496] ,
         \round_in[0][495] , \round_in[0][494] , \round_in[0][493] ,
         \round_in[0][492] , \round_in[0][491] , \round_in[0][490] ,
         \round_in[0][489] , \round_in[0][488] , \round_in[0][487] ,
         \round_in[0][486] , \round_in[0][485] , \round_in[0][484] ,
         \round_in[0][483] , \round_in[0][482] , \round_in[0][481] ,
         \round_in[0][480] , \round_in[0][479] , \round_in[0][478] ,
         \round_in[0][477] , \round_in[0][476] , \round_in[0][475] ,
         \round_in[0][474] , \round_in[0][473] , \round_in[0][472] ,
         \round_in[0][471] , \round_in[0][470] , \round_in[0][469] ,
         \round_in[0][468] , \round_in[0][467] , \round_in[0][466] ,
         \round_in[0][465] , \round_in[0][464] , \round_in[0][463] ,
         \round_in[0][462] , \round_in[0][461] , \round_in[0][460] ,
         \round_in[0][459] , \round_in[0][458] , \round_in[0][457] ,
         \round_in[0][456] , \round_in[0][455] , \round_in[0][454] ,
         \round_in[0][453] , \round_in[0][452] , \round_in[0][451] ,
         \round_in[0][450] , \round_in[0][449] , \round_in[0][448] ,
         \round_in[0][447] , \round_in[0][446] , \round_in[0][445] ,
         \round_in[0][444] , \round_in[0][443] , \round_in[0][442] ,
         \round_in[0][441] , \round_in[0][440] , \round_in[0][439] ,
         \round_in[0][438] , \round_in[0][437] , \round_in[0][436] ,
         \round_in[0][435] , \round_in[0][434] , \round_in[0][433] ,
         \round_in[0][432] , \round_in[0][431] , \round_in[0][430] ,
         \round_in[0][429] , \round_in[0][428] , \round_in[0][427] ,
         \round_in[0][426] , \round_in[0][425] , \round_in[0][424] ,
         \round_in[0][423] , \round_in[0][422] , \round_in[0][421] ,
         \round_in[0][420] , \round_in[0][419] , \round_in[0][418] ,
         \round_in[0][417] , \round_in[0][416] , \round_in[0][415] ,
         \round_in[0][414] , \round_in[0][413] , \round_in[0][412] ,
         \round_in[0][411] , \round_in[0][410] , \round_in[0][409] ,
         \round_in[0][408] , \round_in[0][407] , \round_in[0][406] ,
         \round_in[0][405] , \round_in[0][404] , \round_in[0][403] ,
         \round_in[0][402] , \round_in[0][401] , \round_in[0][400] ,
         \round_in[0][399] , \round_in[0][398] , \round_in[0][397] ,
         \round_in[0][396] , \round_in[0][395] , \round_in[0][394] ,
         \round_in[0][393] , \round_in[0][392] , \round_in[0][391] ,
         \round_in[0][390] , \round_in[0][389] , \round_in[0][388] ,
         \round_in[0][387] , \round_in[0][386] , \round_in[0][385] ,
         \round_in[0][384] , \round_in[0][383] , \round_in[0][382] ,
         \round_in[0][381] , \round_in[0][380] , \round_in[0][379] ,
         \round_in[0][378] , \round_in[0][377] , \round_in[0][376] ,
         \round_in[0][375] , \round_in[0][374] , \round_in[0][373] ,
         \round_in[0][372] , \round_in[0][371] , \round_in[0][370] ,
         \round_in[0][369] , \round_in[0][368] , \round_in[0][367] ,
         \round_in[0][366] , \round_in[0][365] , \round_in[0][364] ,
         \round_in[0][363] , \round_in[0][362] , \round_in[0][361] ,
         \round_in[0][360] , \round_in[0][359] , \round_in[0][358] ,
         \round_in[0][357] , \round_in[0][356] , \round_in[0][355] ,
         \round_in[0][354] , \round_in[0][353] , \round_in[0][352] ,
         \round_in[0][351] , \round_in[0][350] , \round_in[0][349] ,
         \round_in[0][348] , \round_in[0][347] , \round_in[0][346] ,
         \round_in[0][345] , \round_in[0][344] , \round_in[0][343] ,
         \round_in[0][342] , \round_in[0][341] , \round_in[0][340] ,
         \round_in[0][339] , \round_in[0][338] , \round_in[0][337] ,
         \round_in[0][336] , \round_in[0][335] , \round_in[0][334] ,
         \round_in[0][333] , \round_in[0][332] , \round_in[0][331] ,
         \round_in[0][330] , \round_in[0][329] , \round_in[0][328] ,
         \round_in[0][327] , \round_in[0][326] , \round_in[0][325] ,
         \round_in[0][324] , \round_in[0][323] , \round_in[0][322] ,
         \round_in[0][321] , \round_in[0][320] , \round_in[0][319] ,
         \round_in[0][318] , \round_in[0][317] , \round_in[0][316] ,
         \round_in[0][315] , \round_in[0][314] , \round_in[0][313] ,
         \round_in[0][312] , \round_in[0][311] , \round_in[0][310] ,
         \round_in[0][309] , \round_in[0][308] , \round_in[0][307] ,
         \round_in[0][306] , \round_in[0][305] , \round_in[0][304] ,
         \round_in[0][303] , \round_in[0][302] , \round_in[0][301] ,
         \round_in[0][300] , \round_in[0][299] , \round_in[0][298] ,
         \round_in[0][297] , \round_in[0][296] , \round_in[0][295] ,
         \round_in[0][294] , \round_in[0][293] , \round_in[0][292] ,
         \round_in[0][291] , \round_in[0][290] , \round_in[0][289] ,
         \round_in[0][288] , \round_in[0][287] , \round_in[0][286] ,
         \round_in[0][285] , \round_in[0][284] , \round_in[0][283] ,
         \round_in[0][282] , \round_in[0][281] , \round_in[0][280] ,
         \round_in[0][279] , \round_in[0][278] , \round_in[0][277] ,
         \round_in[0][276] , \round_in[0][275] , \round_in[0][274] ,
         \round_in[0][273] , \round_in[0][272] , \round_in[0][271] ,
         \round_in[0][270] , \round_in[0][269] , \round_in[0][268] ,
         \round_in[0][267] , \round_in[0][266] , \round_in[0][265] ,
         \round_in[0][264] , \round_in[0][263] , \round_in[0][262] ,
         \round_in[0][261] , \round_in[0][260] , \round_in[0][259] ,
         \round_in[0][258] , \round_in[0][257] , \round_in[0][256] ,
         \round_in[0][255] , \round_in[0][254] , \round_in[0][253] ,
         \round_in[0][252] , \round_in[0][251] , \round_in[0][250] ,
         \round_in[0][249] , \round_in[0][248] , \round_in[0][247] ,
         \round_in[0][246] , \round_in[0][245] , \round_in[0][244] ,
         \round_in[0][243] , \round_in[0][242] , \round_in[0][241] ,
         \round_in[0][240] , \round_in[0][239] , \round_in[0][238] ,
         \round_in[0][237] , \round_in[0][236] , \round_in[0][235] ,
         \round_in[0][234] , \round_in[0][233] , \round_in[0][232] ,
         \round_in[0][231] , \round_in[0][230] , \round_in[0][229] ,
         \round_in[0][228] , \round_in[0][227] , \round_in[0][226] ,
         \round_in[0][225] , \round_in[0][224] , \round_in[0][223] ,
         \round_in[0][222] , \round_in[0][221] , \round_in[0][220] ,
         \round_in[0][219] , \round_in[0][218] , \round_in[0][217] ,
         \round_in[0][216] , \round_in[0][215] , \round_in[0][214] ,
         \round_in[0][213] , \round_in[0][212] , \round_in[0][211] ,
         \round_in[0][210] , \round_in[0][209] , \round_in[0][208] ,
         \round_in[0][207] , \round_in[0][206] , \round_in[0][205] ,
         \round_in[0][204] , \round_in[0][203] , \round_in[0][202] ,
         \round_in[0][201] , \round_in[0][200] , \round_in[0][199] ,
         \round_in[0][198] , \round_in[0][197] , \round_in[0][196] ,
         \round_in[0][195] , \round_in[0][194] , \round_in[0][193] ,
         \round_in[0][192] , \round_in[0][191] , \round_in[0][190] ,
         \round_in[0][189] , \round_in[0][188] , \round_in[0][187] ,
         \round_in[0][186] , \round_in[0][185] , \round_in[0][184] ,
         \round_in[0][183] , \round_in[0][182] , \round_in[0][181] ,
         \round_in[0][180] , \round_in[0][179] , \round_in[0][178] ,
         \round_in[0][177] , \round_in[0][176] , \round_in[0][175] ,
         \round_in[0][174] , \round_in[0][173] , \round_in[0][172] ,
         \round_in[0][171] , \round_in[0][170] , \round_in[0][169] ,
         \round_in[0][168] , \round_in[0][167] , \round_in[0][166] ,
         \round_in[0][165] , \round_in[0][164] , \round_in[0][163] ,
         \round_in[0][162] , \round_in[0][161] , \round_in[0][160] ,
         \round_in[0][159] , \round_in[0][158] , \round_in[0][157] ,
         \round_in[0][156] , \round_in[0][155] , \round_in[0][154] ,
         \round_in[0][153] , \round_in[0][152] , \round_in[0][151] ,
         \round_in[0][150] , \round_in[0][149] , \round_in[0][148] ,
         \round_in[0][147] , \round_in[0][146] , \round_in[0][145] ,
         \round_in[0][144] , \round_in[0][143] , \round_in[0][142] ,
         \round_in[0][141] , \round_in[0][140] , \round_in[0][139] ,
         \round_in[0][138] , \round_in[0][137] , \round_in[0][136] ,
         \round_in[0][135] , \round_in[0][134] , \round_in[0][133] ,
         \round_in[0][132] , \round_in[0][131] , \round_in[0][130] ,
         \round_in[0][129] , \round_in[0][128] , \round_in[0][127] ,
         \round_in[0][126] , \round_in[0][125] , \round_in[0][124] ,
         \round_in[0][123] , \round_in[0][122] , \round_in[0][121] ,
         \round_in[0][120] , \round_in[0][119] , \round_in[0][118] ,
         \round_in[0][117] , \round_in[0][116] , \round_in[0][115] ,
         \round_in[0][114] , \round_in[0][113] , \round_in[0][112] ,
         \round_in[0][111] , \round_in[0][110] , \round_in[0][109] ,
         \round_in[0][108] , \round_in[0][107] , \round_in[0][106] ,
         \round_in[0][105] , \round_in[0][104] , \round_in[0][103] ,
         \round_in[0][102] , \round_in[0][101] , \round_in[0][100] ,
         \round_in[0][99] , \round_in[0][98] , \round_in[0][97] ,
         \round_in[0][96] , \round_in[0][95] , \round_in[0][94] ,
         \round_in[0][93] , \round_in[0][92] , \round_in[0][91] ,
         \round_in[0][90] , \round_in[0][89] , \round_in[0][88] ,
         \round_in[0][87] , \round_in[0][86] , \round_in[0][85] ,
         \round_in[0][84] , \round_in[0][83] , \round_in[0][82] ,
         \round_in[0][81] , \round_in[0][80] , \round_in[0][79] ,
         \round_in[0][78] , \round_in[0][77] , \round_in[0][76] ,
         \round_in[0][75] , \round_in[0][74] , \round_in[0][73] ,
         \round_in[0][72] , \round_in[0][71] , \round_in[0][70] ,
         \round_in[0][69] , \round_in[0][68] , \round_in[0][67] ,
         \round_in[0][66] , \round_in[0][65] , \round_in[0][64] ,
         \round_in[0][63] , \round_in[0][62] , \round_in[0][61] ,
         \round_in[0][60] , \round_in[0][59] , \round_in[0][58] ,
         \round_in[0][57] , \round_in[0][56] , \round_in[0][55] ,
         \round_in[0][54] , \round_in[0][53] , \round_in[0][52] ,
         \round_in[0][51] , \round_in[0][50] , \round_in[0][49] ,
         \round_in[0][48] , \round_in[0][47] , \round_in[0][46] ,
         \round_in[0][45] , \round_in[0][44] , \round_in[0][43] ,
         \round_in[0][42] , \round_in[0][41] , \round_in[0][40] ,
         \round_in[0][39] , \round_in[0][38] , \round_in[0][37] ,
         \round_in[0][36] , \round_in[0][35] , \round_in[0][34] ,
         \round_in[0][33] , \round_in[0][32] , \round_in[0][31] ,
         \round_in[0][30] , \round_in[0][29] , \round_in[0][28] ,
         \round_in[0][27] , \round_in[0][26] , \round_in[0][25] ,
         \round_in[0][24] , \round_in[0][23] , \round_in[0][22] ,
         \round_in[0][21] , \round_in[0][20] , \round_in[0][19] ,
         \round_in[0][18] , \round_in[0][17] , \round_in[0][16] ,
         \round_in[0][15] , \round_in[0][14] , \round_in[0][13] ,
         \round_in[0][12] , \round_in[0][11] , \round_in[0][10] ,
         \round_in[0][9] , \round_in[0][8] , \round_in[0][7] ,
         \round_in[0][6] , \round_in[0][5] , \round_in[0][4] ,
         \round_in[0][3] , \round_in[0][2] , \round_in[0][1] ,
         \round_in[0][0] , \rc[3][63] , \rc[3][31] , \rc[3][15] , \rc[3][3] ,
         \rc[3][1] , \rc[2][0] , \rc[1][7] , \RCONST[0].rconst_/N67 ,
         \RCONST[0].rconst_/N56 , \RCONST[0].rconst_/N48 ,
         \RCONST[0].rconst_/N25 , \RCONST[0].rconst_/N17 ,
         \RCONST[1].rconst_/N68 , \RCONST[1].rconst_/N49 ,
         \RCONST[1].rconst_/N26 , \RCONST[1].rconst_/N15 ,
         \RCONST[2].rconst_/N62 , \RCONST[2].rconst_/N57 ,
         \RCONST[2].rconst_/N47 , \RCONST[2].rconst_/N28 ,
         \RCONST[2].rconst_/N18 , \RCONST[3].rconst_/N10 , n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916;
  wire   [5:0] rc_i;
  wire   [1599:0] round_reg;

  round_2 \ROUND[0].round_  ( .in({\round_in[0][1599] , \round_in[0][1598] , 
        \round_in[0][1597] , \round_in[0][1596] , \round_in[0][1595] , 
        \round_in[0][1594] , \round_in[0][1593] , \round_in[0][1592] , 
        \round_in[0][1591] , \round_in[0][1590] , \round_in[0][1589] , 
        \round_in[0][1588] , \round_in[0][1587] , \round_in[0][1586] , 
        \round_in[0][1585] , \round_in[0][1584] , \round_in[0][1583] , 
        \round_in[0][1582] , \round_in[0][1581] , \round_in[0][1580] , 
        \round_in[0][1579] , \round_in[0][1578] , \round_in[0][1577] , 
        \round_in[0][1576] , \round_in[0][1575] , \round_in[0][1574] , 
        \round_in[0][1573] , \round_in[0][1572] , \round_in[0][1571] , 
        \round_in[0][1570] , \round_in[0][1569] , \round_in[0][1568] , 
        \round_in[0][1567] , \round_in[0][1566] , \round_in[0][1565] , 
        \round_in[0][1564] , \round_in[0][1563] , \round_in[0][1562] , 
        \round_in[0][1561] , \round_in[0][1560] , \round_in[0][1559] , 
        \round_in[0][1558] , \round_in[0][1557] , \round_in[0][1556] , 
        \round_in[0][1555] , \round_in[0][1554] , \round_in[0][1553] , 
        \round_in[0][1552] , \round_in[0][1551] , \round_in[0][1550] , 
        \round_in[0][1549] , \round_in[0][1548] , \round_in[0][1547] , 
        \round_in[0][1546] , \round_in[0][1545] , \round_in[0][1544] , 
        \round_in[0][1543] , \round_in[0][1542] , \round_in[0][1541] , 
        \round_in[0][1540] , \round_in[0][1539] , \round_in[0][1538] , 
        \round_in[0][1537] , \round_in[0][1536] , \round_in[0][1535] , 
        \round_in[0][1534] , \round_in[0][1533] , \round_in[0][1532] , 
        \round_in[0][1531] , \round_in[0][1530] , \round_in[0][1529] , 
        \round_in[0][1528] , \round_in[0][1527] , \round_in[0][1526] , 
        \round_in[0][1525] , \round_in[0][1524] , \round_in[0][1523] , 
        \round_in[0][1522] , \round_in[0][1521] , \round_in[0][1520] , 
        \round_in[0][1519] , \round_in[0][1518] , \round_in[0][1517] , 
        \round_in[0][1516] , \round_in[0][1515] , \round_in[0][1514] , 
        \round_in[0][1513] , \round_in[0][1512] , \round_in[0][1511] , 
        \round_in[0][1510] , \round_in[0][1509] , \round_in[0][1508] , 
        \round_in[0][1507] , \round_in[0][1506] , \round_in[0][1505] , 
        \round_in[0][1504] , \round_in[0][1503] , \round_in[0][1502] , 
        \round_in[0][1501] , \round_in[0][1500] , \round_in[0][1499] , 
        \round_in[0][1498] , \round_in[0][1497] , \round_in[0][1496] , 
        \round_in[0][1495] , \round_in[0][1494] , \round_in[0][1493] , 
        \round_in[0][1492] , \round_in[0][1491] , \round_in[0][1490] , 
        \round_in[0][1489] , \round_in[0][1488] , \round_in[0][1487] , 
        \round_in[0][1486] , \round_in[0][1485] , \round_in[0][1484] , 
        \round_in[0][1483] , \round_in[0][1482] , \round_in[0][1481] , 
        \round_in[0][1480] , \round_in[0][1479] , \round_in[0][1478] , 
        \round_in[0][1477] , \round_in[0][1476] , \round_in[0][1475] , 
        \round_in[0][1474] , \round_in[0][1473] , \round_in[0][1472] , 
        \round_in[0][1471] , \round_in[0][1470] , \round_in[0][1469] , 
        \round_in[0][1468] , \round_in[0][1467] , \round_in[0][1466] , 
        \round_in[0][1465] , \round_in[0][1464] , \round_in[0][1463] , 
        \round_in[0][1462] , \round_in[0][1461] , \round_in[0][1460] , 
        \round_in[0][1459] , \round_in[0][1458] , \round_in[0][1457] , 
        \round_in[0][1456] , \round_in[0][1455] , \round_in[0][1454] , 
        \round_in[0][1453] , \round_in[0][1452] , \round_in[0][1451] , 
        \round_in[0][1450] , \round_in[0][1449] , \round_in[0][1448] , 
        \round_in[0][1447] , \round_in[0][1446] , \round_in[0][1445] , 
        \round_in[0][1444] , \round_in[0][1443] , \round_in[0][1442] , 
        \round_in[0][1441] , \round_in[0][1440] , \round_in[0][1439] , 
        \round_in[0][1438] , \round_in[0][1437] , \round_in[0][1436] , 
        \round_in[0][1435] , \round_in[0][1434] , \round_in[0][1433] , 
        \round_in[0][1432] , \round_in[0][1431] , \round_in[0][1430] , 
        \round_in[0][1429] , \round_in[0][1428] , \round_in[0][1427] , 
        \round_in[0][1426] , \round_in[0][1425] , \round_in[0][1424] , 
        \round_in[0][1423] , \round_in[0][1422] , \round_in[0][1421] , 
        \round_in[0][1420] , \round_in[0][1419] , \round_in[0][1418] , 
        \round_in[0][1417] , \round_in[0][1416] , \round_in[0][1415] , 
        \round_in[0][1414] , \round_in[0][1413] , \round_in[0][1412] , 
        \round_in[0][1411] , \round_in[0][1410] , \round_in[0][1409] , 
        \round_in[0][1408] , \round_in[0][1407] , \round_in[0][1406] , 
        \round_in[0][1405] , \round_in[0][1404] , \round_in[0][1403] , 
        \round_in[0][1402] , \round_in[0][1401] , \round_in[0][1400] , 
        \round_in[0][1399] , \round_in[0][1398] , \round_in[0][1397] , 
        \round_in[0][1396] , \round_in[0][1395] , \round_in[0][1394] , 
        \round_in[0][1393] , \round_in[0][1392] , \round_in[0][1391] , 
        \round_in[0][1390] , \round_in[0][1389] , \round_in[0][1388] , 
        \round_in[0][1387] , \round_in[0][1386] , \round_in[0][1385] , 
        \round_in[0][1384] , \round_in[0][1383] , \round_in[0][1382] , 
        \round_in[0][1381] , \round_in[0][1380] , \round_in[0][1379] , 
        \round_in[0][1378] , \round_in[0][1377] , \round_in[0][1376] , 
        \round_in[0][1375] , \round_in[0][1374] , \round_in[0][1373] , 
        \round_in[0][1372] , \round_in[0][1371] , \round_in[0][1370] , 
        \round_in[0][1369] , \round_in[0][1368] , \round_in[0][1367] , 
        \round_in[0][1366] , \round_in[0][1365] , \round_in[0][1364] , 
        \round_in[0][1363] , \round_in[0][1362] , \round_in[0][1361] , 
        \round_in[0][1360] , \round_in[0][1359] , \round_in[0][1358] , 
        \round_in[0][1357] , \round_in[0][1356] , \round_in[0][1355] , 
        \round_in[0][1354] , \round_in[0][1353] , \round_in[0][1352] , 
        \round_in[0][1351] , \round_in[0][1350] , \round_in[0][1349] , 
        \round_in[0][1348] , \round_in[0][1347] , \round_in[0][1346] , 
        \round_in[0][1345] , \round_in[0][1344] , \round_in[0][1343] , 
        \round_in[0][1342] , \round_in[0][1341] , \round_in[0][1340] , 
        \round_in[0][1339] , \round_in[0][1338] , \round_in[0][1337] , 
        \round_in[0][1336] , \round_in[0][1335] , \round_in[0][1334] , 
        \round_in[0][1333] , \round_in[0][1332] , \round_in[0][1331] , 
        \round_in[0][1330] , \round_in[0][1329] , \round_in[0][1328] , 
        \round_in[0][1327] , \round_in[0][1326] , \round_in[0][1325] , 
        \round_in[0][1324] , \round_in[0][1323] , \round_in[0][1322] , 
        \round_in[0][1321] , \round_in[0][1320] , \round_in[0][1319] , 
        \round_in[0][1318] , \round_in[0][1317] , \round_in[0][1316] , 
        \round_in[0][1315] , \round_in[0][1314] , \round_in[0][1313] , 
        \round_in[0][1312] , \round_in[0][1311] , \round_in[0][1310] , 
        \round_in[0][1309] , \round_in[0][1308] , \round_in[0][1307] , 
        \round_in[0][1306] , \round_in[0][1305] , \round_in[0][1304] , 
        \round_in[0][1303] , \round_in[0][1302] , \round_in[0][1301] , 
        \round_in[0][1300] , \round_in[0][1299] , \round_in[0][1298] , 
        \round_in[0][1297] , \round_in[0][1296] , \round_in[0][1295] , 
        \round_in[0][1294] , \round_in[0][1293] , \round_in[0][1292] , 
        \round_in[0][1291] , \round_in[0][1290] , \round_in[0][1289] , 
        \round_in[0][1288] , \round_in[0][1287] , \round_in[0][1286] , 
        \round_in[0][1285] , \round_in[0][1284] , \round_in[0][1283] , 
        \round_in[0][1282] , \round_in[0][1281] , \round_in[0][1280] , 
        \round_in[0][1279] , \round_in[0][1278] , \round_in[0][1277] , 
        \round_in[0][1276] , \round_in[0][1275] , \round_in[0][1274] , 
        \round_in[0][1273] , \round_in[0][1272] , \round_in[0][1271] , 
        \round_in[0][1270] , \round_in[0][1269] , \round_in[0][1268] , 
        \round_in[0][1267] , \round_in[0][1266] , \round_in[0][1265] , 
        \round_in[0][1264] , \round_in[0][1263] , \round_in[0][1262] , 
        \round_in[0][1261] , \round_in[0][1260] , \round_in[0][1259] , 
        \round_in[0][1258] , \round_in[0][1257] , \round_in[0][1256] , 
        \round_in[0][1255] , \round_in[0][1254] , \round_in[0][1253] , 
        \round_in[0][1252] , \round_in[0][1251] , \round_in[0][1250] , 
        \round_in[0][1249] , \round_in[0][1248] , \round_in[0][1247] , 
        \round_in[0][1246] , \round_in[0][1245] , \round_in[0][1244] , 
        \round_in[0][1243] , \round_in[0][1242] , \round_in[0][1241] , 
        \round_in[0][1240] , \round_in[0][1239] , \round_in[0][1238] , 
        \round_in[0][1237] , \round_in[0][1236] , \round_in[0][1235] , 
        \round_in[0][1234] , \round_in[0][1233] , \round_in[0][1232] , 
        \round_in[0][1231] , \round_in[0][1230] , \round_in[0][1229] , 
        \round_in[0][1228] , \round_in[0][1227] , \round_in[0][1226] , 
        \round_in[0][1225] , \round_in[0][1224] , \round_in[0][1223] , 
        \round_in[0][1222] , \round_in[0][1221] , \round_in[0][1220] , 
        \round_in[0][1219] , \round_in[0][1218] , \round_in[0][1217] , 
        \round_in[0][1216] , \round_in[0][1215] , \round_in[0][1214] , 
        \round_in[0][1213] , \round_in[0][1212] , \round_in[0][1211] , 
        \round_in[0][1210] , \round_in[0][1209] , \round_in[0][1208] , 
        \round_in[0][1207] , \round_in[0][1206] , \round_in[0][1205] , 
        \round_in[0][1204] , \round_in[0][1203] , \round_in[0][1202] , 
        \round_in[0][1201] , \round_in[0][1200] , \round_in[0][1199] , 
        \round_in[0][1198] , \round_in[0][1197] , \round_in[0][1196] , 
        \round_in[0][1195] , \round_in[0][1194] , \round_in[0][1193] , 
        \round_in[0][1192] , \round_in[0][1191] , \round_in[0][1190] , 
        \round_in[0][1189] , \round_in[0][1188] , \round_in[0][1187] , 
        \round_in[0][1186] , \round_in[0][1185] , \round_in[0][1184] , 
        \round_in[0][1183] , \round_in[0][1182] , \round_in[0][1181] , 
        \round_in[0][1180] , \round_in[0][1179] , \round_in[0][1178] , 
        \round_in[0][1177] , \round_in[0][1176] , \round_in[0][1175] , 
        \round_in[0][1174] , \round_in[0][1173] , \round_in[0][1172] , 
        \round_in[0][1171] , \round_in[0][1170] , \round_in[0][1169] , 
        \round_in[0][1168] , \round_in[0][1167] , \round_in[0][1166] , 
        \round_in[0][1165] , \round_in[0][1164] , \round_in[0][1163] , 
        \round_in[0][1162] , \round_in[0][1161] , \round_in[0][1160] , 
        \round_in[0][1159] , \round_in[0][1158] , \round_in[0][1157] , 
        \round_in[0][1156] , \round_in[0][1155] , \round_in[0][1154] , 
        \round_in[0][1153] , \round_in[0][1152] , \round_in[0][1151] , 
        \round_in[0][1150] , \round_in[0][1149] , \round_in[0][1148] , 
        \round_in[0][1147] , \round_in[0][1146] , \round_in[0][1145] , 
        \round_in[0][1144] , \round_in[0][1143] , \round_in[0][1142] , 
        \round_in[0][1141] , \round_in[0][1140] , \round_in[0][1139] , 
        \round_in[0][1138] , \round_in[0][1137] , \round_in[0][1136] , 
        \round_in[0][1135] , \round_in[0][1134] , \round_in[0][1133] , 
        \round_in[0][1132] , \round_in[0][1131] , \round_in[0][1130] , 
        \round_in[0][1129] , \round_in[0][1128] , \round_in[0][1127] , 
        \round_in[0][1126] , \round_in[0][1125] , \round_in[0][1124] , 
        \round_in[0][1123] , \round_in[0][1122] , \round_in[0][1121] , 
        \round_in[0][1120] , \round_in[0][1119] , \round_in[0][1118] , 
        \round_in[0][1117] , \round_in[0][1116] , \round_in[0][1115] , 
        \round_in[0][1114] , \round_in[0][1113] , \round_in[0][1112] , 
        \round_in[0][1111] , \round_in[0][1110] , \round_in[0][1109] , 
        \round_in[0][1108] , \round_in[0][1107] , \round_in[0][1106] , 
        \round_in[0][1105] , \round_in[0][1104] , \round_in[0][1103] , 
        \round_in[0][1102] , \round_in[0][1101] , \round_in[0][1100] , 
        \round_in[0][1099] , \round_in[0][1098] , \round_in[0][1097] , 
        \round_in[0][1096] , \round_in[0][1095] , \round_in[0][1094] , 
        \round_in[0][1093] , \round_in[0][1092] , \round_in[0][1091] , 
        \round_in[0][1090] , \round_in[0][1089] , \round_in[0][1088] , 
        \round_in[0][1087] , \round_in[0][1086] , \round_in[0][1085] , 
        \round_in[0][1084] , \round_in[0][1083] , \round_in[0][1082] , 
        \round_in[0][1081] , \round_in[0][1080] , \round_in[0][1079] , 
        \round_in[0][1078] , \round_in[0][1077] , \round_in[0][1076] , 
        \round_in[0][1075] , \round_in[0][1074] , \round_in[0][1073] , 
        \round_in[0][1072] , \round_in[0][1071] , \round_in[0][1070] , 
        \round_in[0][1069] , \round_in[0][1068] , \round_in[0][1067] , 
        \round_in[0][1066] , \round_in[0][1065] , \round_in[0][1064] , 
        \round_in[0][1063] , \round_in[0][1062] , \round_in[0][1061] , 
        \round_in[0][1060] , \round_in[0][1059] , \round_in[0][1058] , 
        \round_in[0][1057] , \round_in[0][1056] , \round_in[0][1055] , 
        \round_in[0][1054] , \round_in[0][1053] , \round_in[0][1052] , 
        \round_in[0][1051] , \round_in[0][1050] , \round_in[0][1049] , 
        \round_in[0][1048] , \round_in[0][1047] , \round_in[0][1046] , 
        \round_in[0][1045] , \round_in[0][1044] , \round_in[0][1043] , 
        \round_in[0][1042] , \round_in[0][1041] , \round_in[0][1040] , 
        \round_in[0][1039] , \round_in[0][1038] , \round_in[0][1037] , 
        \round_in[0][1036] , \round_in[0][1035] , \round_in[0][1034] , 
        \round_in[0][1033] , \round_in[0][1032] , \round_in[0][1031] , 
        \round_in[0][1030] , \round_in[0][1029] , \round_in[0][1028] , 
        \round_in[0][1027] , \round_in[0][1026] , \round_in[0][1025] , 
        \round_in[0][1024] , \round_in[0][1023] , \round_in[0][1022] , 
        \round_in[0][1021] , \round_in[0][1020] , \round_in[0][1019] , 
        \round_in[0][1018] , \round_in[0][1017] , \round_in[0][1016] , 
        \round_in[0][1015] , \round_in[0][1014] , \round_in[0][1013] , 
        \round_in[0][1012] , \round_in[0][1011] , \round_in[0][1010] , 
        \round_in[0][1009] , \round_in[0][1008] , \round_in[0][1007] , 
        \round_in[0][1006] , \round_in[0][1005] , \round_in[0][1004] , 
        \round_in[0][1003] , \round_in[0][1002] , \round_in[0][1001] , 
        \round_in[0][1000] , \round_in[0][999] , \round_in[0][998] , 
        \round_in[0][997] , \round_in[0][996] , \round_in[0][995] , 
        \round_in[0][994] , \round_in[0][993] , \round_in[0][992] , 
        \round_in[0][991] , \round_in[0][990] , \round_in[0][989] , 
        \round_in[0][988] , \round_in[0][987] , \round_in[0][986] , 
        \round_in[0][985] , \round_in[0][984] , \round_in[0][983] , 
        \round_in[0][982] , \round_in[0][981] , \round_in[0][980] , 
        \round_in[0][979] , \round_in[0][978] , \round_in[0][977] , 
        \round_in[0][976] , \round_in[0][975] , \round_in[0][974] , 
        \round_in[0][973] , \round_in[0][972] , \round_in[0][971] , 
        \round_in[0][970] , \round_in[0][969] , \round_in[0][968] , 
        \round_in[0][967] , \round_in[0][966] , \round_in[0][965] , 
        \round_in[0][964] , \round_in[0][963] , \round_in[0][962] , 
        \round_in[0][961] , \round_in[0][960] , \round_in[0][959] , 
        \round_in[0][958] , \round_in[0][957] , \round_in[0][956] , 
        \round_in[0][955] , \round_in[0][954] , \round_in[0][953] , 
        \round_in[0][952] , \round_in[0][951] , \round_in[0][950] , 
        \round_in[0][949] , \round_in[0][948] , \round_in[0][947] , 
        \round_in[0][946] , \round_in[0][945] , \round_in[0][944] , 
        \round_in[0][943] , \round_in[0][942] , \round_in[0][941] , 
        \round_in[0][940] , \round_in[0][939] , \round_in[0][938] , 
        \round_in[0][937] , \round_in[0][936] , \round_in[0][935] , 
        \round_in[0][934] , \round_in[0][933] , \round_in[0][932] , 
        \round_in[0][931] , \round_in[0][930] , \round_in[0][929] , 
        \round_in[0][928] , \round_in[0][927] , \round_in[0][926] , 
        \round_in[0][925] , \round_in[0][924] , \round_in[0][923] , 
        \round_in[0][922] , \round_in[0][921] , \round_in[0][920] , 
        \round_in[0][919] , \round_in[0][918] , \round_in[0][917] , 
        \round_in[0][916] , \round_in[0][915] , \round_in[0][914] , 
        \round_in[0][913] , \round_in[0][912] , \round_in[0][911] , 
        \round_in[0][910] , \round_in[0][909] , \round_in[0][908] , 
        \round_in[0][907] , \round_in[0][906] , \round_in[0][905] , 
        \round_in[0][904] , \round_in[0][903] , \round_in[0][902] , 
        \round_in[0][901] , \round_in[0][900] , \round_in[0][899] , 
        \round_in[0][898] , \round_in[0][897] , \round_in[0][896] , 
        \round_in[0][895] , \round_in[0][894] , \round_in[0][893] , 
        \round_in[0][892] , \round_in[0][891] , \round_in[0][890] , 
        \round_in[0][889] , \round_in[0][888] , \round_in[0][887] , 
        \round_in[0][886] , \round_in[0][885] , \round_in[0][884] , 
        \round_in[0][883] , \round_in[0][882] , \round_in[0][881] , 
        \round_in[0][880] , \round_in[0][879] , \round_in[0][878] , 
        \round_in[0][877] , \round_in[0][876] , \round_in[0][875] , 
        \round_in[0][874] , \round_in[0][873] , \round_in[0][872] , 
        \round_in[0][871] , \round_in[0][870] , \round_in[0][869] , 
        \round_in[0][868] , \round_in[0][867] , \round_in[0][866] , 
        \round_in[0][865] , \round_in[0][864] , \round_in[0][863] , 
        \round_in[0][862] , \round_in[0][861] , \round_in[0][860] , 
        \round_in[0][859] , \round_in[0][858] , \round_in[0][857] , 
        \round_in[0][856] , \round_in[0][855] , \round_in[0][854] , 
        \round_in[0][853] , \round_in[0][852] , \round_in[0][851] , 
        \round_in[0][850] , \round_in[0][849] , \round_in[0][848] , 
        \round_in[0][847] , \round_in[0][846] , \round_in[0][845] , 
        \round_in[0][844] , \round_in[0][843] , \round_in[0][842] , 
        \round_in[0][841] , \round_in[0][840] , \round_in[0][839] , 
        \round_in[0][838] , \round_in[0][837] , \round_in[0][836] , 
        \round_in[0][835] , \round_in[0][834] , \round_in[0][833] , 
        \round_in[0][832] , \round_in[0][831] , \round_in[0][830] , 
        \round_in[0][829] , \round_in[0][828] , \round_in[0][827] , 
        \round_in[0][826] , \round_in[0][825] , \round_in[0][824] , 
        \round_in[0][823] , \round_in[0][822] , \round_in[0][821] , 
        \round_in[0][820] , \round_in[0][819] , \round_in[0][818] , 
        \round_in[0][817] , \round_in[0][816] , \round_in[0][815] , 
        \round_in[0][814] , \round_in[0][813] , \round_in[0][812] , 
        \round_in[0][811] , \round_in[0][810] , \round_in[0][809] , 
        \round_in[0][808] , \round_in[0][807] , \round_in[0][806] , 
        \round_in[0][805] , \round_in[0][804] , \round_in[0][803] , 
        \round_in[0][802] , \round_in[0][801] , \round_in[0][800] , 
        \round_in[0][799] , \round_in[0][798] , \round_in[0][797] , 
        \round_in[0][796] , \round_in[0][795] , \round_in[0][794] , 
        \round_in[0][793] , \round_in[0][792] , \round_in[0][791] , 
        \round_in[0][790] , \round_in[0][789] , \round_in[0][788] , 
        \round_in[0][787] , \round_in[0][786] , \round_in[0][785] , 
        \round_in[0][784] , \round_in[0][783] , \round_in[0][782] , 
        \round_in[0][781] , \round_in[0][780] , \round_in[0][779] , 
        \round_in[0][778] , \round_in[0][777] , \round_in[0][776] , 
        \round_in[0][775] , \round_in[0][774] , \round_in[0][773] , 
        \round_in[0][772] , \round_in[0][771] , \round_in[0][770] , 
        \round_in[0][769] , \round_in[0][768] , \round_in[0][767] , 
        \round_in[0][766] , \round_in[0][765] , \round_in[0][764] , 
        \round_in[0][763] , \round_in[0][762] , \round_in[0][761] , 
        \round_in[0][760] , \round_in[0][759] , \round_in[0][758] , 
        \round_in[0][757] , \round_in[0][756] , \round_in[0][755] , 
        \round_in[0][754] , \round_in[0][753] , \round_in[0][752] , 
        \round_in[0][751] , \round_in[0][750] , \round_in[0][749] , 
        \round_in[0][748] , \round_in[0][747] , \round_in[0][746] , 
        \round_in[0][745] , \round_in[0][744] , \round_in[0][743] , 
        \round_in[0][742] , \round_in[0][741] , \round_in[0][740] , 
        \round_in[0][739] , \round_in[0][738] , \round_in[0][737] , 
        \round_in[0][736] , \round_in[0][735] , \round_in[0][734] , 
        \round_in[0][733] , \round_in[0][732] , \round_in[0][731] , 
        \round_in[0][730] , \round_in[0][729] , \round_in[0][728] , 
        \round_in[0][727] , \round_in[0][726] , \round_in[0][725] , 
        \round_in[0][724] , \round_in[0][723] , \round_in[0][722] , 
        \round_in[0][721] , \round_in[0][720] , \round_in[0][719] , 
        \round_in[0][718] , \round_in[0][717] , \round_in[0][716] , 
        \round_in[0][715] , \round_in[0][714] , \round_in[0][713] , 
        \round_in[0][712] , \round_in[0][711] , \round_in[0][710] , 
        \round_in[0][709] , \round_in[0][708] , \round_in[0][707] , 
        \round_in[0][706] , \round_in[0][705] , \round_in[0][704] , 
        \round_in[0][703] , \round_in[0][702] , \round_in[0][701] , 
        \round_in[0][700] , \round_in[0][699] , \round_in[0][698] , 
        \round_in[0][697] , \round_in[0][696] , \round_in[0][695] , 
        \round_in[0][694] , \round_in[0][693] , \round_in[0][692] , 
        \round_in[0][691] , \round_in[0][690] , \round_in[0][689] , 
        \round_in[0][688] , \round_in[0][687] , \round_in[0][686] , 
        \round_in[0][685] , \round_in[0][684] , \round_in[0][683] , 
        \round_in[0][682] , \round_in[0][681] , \round_in[0][680] , 
        \round_in[0][679] , \round_in[0][678] , \round_in[0][677] , 
        \round_in[0][676] , \round_in[0][675] , \round_in[0][674] , 
        \round_in[0][673] , \round_in[0][672] , \round_in[0][671] , 
        \round_in[0][670] , \round_in[0][669] , \round_in[0][668] , 
        \round_in[0][667] , \round_in[0][666] , \round_in[0][665] , 
        \round_in[0][664] , \round_in[0][663] , \round_in[0][662] , 
        \round_in[0][661] , \round_in[0][660] , \round_in[0][659] , 
        \round_in[0][658] , \round_in[0][657] , \round_in[0][656] , 
        \round_in[0][655] , \round_in[0][654] , \round_in[0][653] , 
        \round_in[0][652] , \round_in[0][651] , \round_in[0][650] , 
        \round_in[0][649] , \round_in[0][648] , \round_in[0][647] , 
        \round_in[0][646] , \round_in[0][645] , \round_in[0][644] , 
        \round_in[0][643] , \round_in[0][642] , \round_in[0][641] , 
        \round_in[0][640] , \round_in[0][639] , \round_in[0][638] , 
        \round_in[0][637] , \round_in[0][636] , \round_in[0][635] , 
        \round_in[0][634] , \round_in[0][633] , \round_in[0][632] , 
        \round_in[0][631] , \round_in[0][630] , \round_in[0][629] , 
        \round_in[0][628] , \round_in[0][627] , \round_in[0][626] , 
        \round_in[0][625] , \round_in[0][624] , \round_in[0][623] , 
        \round_in[0][622] , \round_in[0][621] , \round_in[0][620] , 
        \round_in[0][619] , \round_in[0][618] , \round_in[0][617] , 
        \round_in[0][616] , \round_in[0][615] , \round_in[0][614] , 
        \round_in[0][613] , \round_in[0][612] , \round_in[0][611] , 
        \round_in[0][610] , \round_in[0][609] , \round_in[0][608] , 
        \round_in[0][607] , \round_in[0][606] , \round_in[0][605] , 
        \round_in[0][604] , \round_in[0][603] , \round_in[0][602] , 
        \round_in[0][601] , \round_in[0][600] , \round_in[0][599] , 
        \round_in[0][598] , \round_in[0][597] , \round_in[0][596] , 
        \round_in[0][595] , \round_in[0][594] , \round_in[0][593] , 
        \round_in[0][592] , \round_in[0][591] , \round_in[0][590] , 
        \round_in[0][589] , \round_in[0][588] , \round_in[0][587] , 
        \round_in[0][586] , \round_in[0][585] , \round_in[0][584] , 
        \round_in[0][583] , \round_in[0][582] , \round_in[0][581] , 
        \round_in[0][580] , \round_in[0][579] , \round_in[0][578] , 
        \round_in[0][577] , \round_in[0][576] , \round_in[0][575] , 
        \round_in[0][574] , \round_in[0][573] , \round_in[0][572] , 
        \round_in[0][571] , \round_in[0][570] , \round_in[0][569] , 
        \round_in[0][568] , \round_in[0][567] , \round_in[0][566] , 
        \round_in[0][565] , \round_in[0][564] , \round_in[0][563] , 
        \round_in[0][562] , \round_in[0][561] , \round_in[0][560] , 
        \round_in[0][559] , \round_in[0][558] , \round_in[0][557] , 
        \round_in[0][556] , \round_in[0][555] , \round_in[0][554] , 
        \round_in[0][553] , \round_in[0][552] , \round_in[0][551] , 
        \round_in[0][550] , \round_in[0][549] , \round_in[0][548] , 
        \round_in[0][547] , \round_in[0][546] , \round_in[0][545] , 
        \round_in[0][544] , \round_in[0][543] , \round_in[0][542] , 
        \round_in[0][541] , \round_in[0][540] , \round_in[0][539] , 
        \round_in[0][538] , \round_in[0][537] , \round_in[0][536] , 
        \round_in[0][535] , \round_in[0][534] , \round_in[0][533] , 
        \round_in[0][532] , \round_in[0][531] , \round_in[0][530] , 
        \round_in[0][529] , \round_in[0][528] , \round_in[0][527] , 
        \round_in[0][526] , \round_in[0][525] , \round_in[0][524] , 
        \round_in[0][523] , \round_in[0][522] , \round_in[0][521] , 
        \round_in[0][520] , \round_in[0][519] , \round_in[0][518] , 
        \round_in[0][517] , \round_in[0][516] , \round_in[0][515] , 
        \round_in[0][514] , \round_in[0][513] , \round_in[0][512] , 
        \round_in[0][511] , \round_in[0][510] , \round_in[0][509] , 
        \round_in[0][508] , \round_in[0][507] , \round_in[0][506] , 
        \round_in[0][505] , \round_in[0][504] , \round_in[0][503] , 
        \round_in[0][502] , \round_in[0][501] , \round_in[0][500] , 
        \round_in[0][499] , \round_in[0][498] , \round_in[0][497] , 
        \round_in[0][496] , \round_in[0][495] , \round_in[0][494] , 
        \round_in[0][493] , \round_in[0][492] , \round_in[0][491] , 
        \round_in[0][490] , \round_in[0][489] , \round_in[0][488] , 
        \round_in[0][487] , \round_in[0][486] , \round_in[0][485] , 
        \round_in[0][484] , \round_in[0][483] , \round_in[0][482] , 
        \round_in[0][481] , \round_in[0][480] , \round_in[0][479] , 
        \round_in[0][478] , \round_in[0][477] , \round_in[0][476] , 
        \round_in[0][475] , \round_in[0][474] , \round_in[0][473] , 
        \round_in[0][472] , \round_in[0][471] , \round_in[0][470] , 
        \round_in[0][469] , \round_in[0][468] , \round_in[0][467] , 
        \round_in[0][466] , \round_in[0][465] , \round_in[0][464] , 
        \round_in[0][463] , \round_in[0][462] , \round_in[0][461] , 
        \round_in[0][460] , \round_in[0][459] , \round_in[0][458] , 
        \round_in[0][457] , \round_in[0][456] , \round_in[0][455] , 
        \round_in[0][454] , \round_in[0][453] , \round_in[0][452] , 
        \round_in[0][451] , \round_in[0][450] , \round_in[0][449] , 
        \round_in[0][448] , \round_in[0][447] , \round_in[0][446] , 
        \round_in[0][445] , \round_in[0][444] , \round_in[0][443] , 
        \round_in[0][442] , \round_in[0][441] , \round_in[0][440] , 
        \round_in[0][439] , \round_in[0][438] , \round_in[0][437] , 
        \round_in[0][436] , \round_in[0][435] , \round_in[0][434] , 
        \round_in[0][433] , \round_in[0][432] , \round_in[0][431] , 
        \round_in[0][430] , \round_in[0][429] , \round_in[0][428] , 
        \round_in[0][427] , \round_in[0][426] , \round_in[0][425] , 
        \round_in[0][424] , \round_in[0][423] , \round_in[0][422] , 
        \round_in[0][421] , \round_in[0][420] , \round_in[0][419] , 
        \round_in[0][418] , \round_in[0][417] , \round_in[0][416] , 
        \round_in[0][415] , \round_in[0][414] , \round_in[0][413] , 
        \round_in[0][412] , \round_in[0][411] , \round_in[0][410] , 
        \round_in[0][409] , \round_in[0][408] , \round_in[0][407] , 
        \round_in[0][406] , \round_in[0][405] , \round_in[0][404] , 
        \round_in[0][403] , \round_in[0][402] , \round_in[0][401] , 
        \round_in[0][400] , \round_in[0][399] , \round_in[0][398] , 
        \round_in[0][397] , \round_in[0][396] , \round_in[0][395] , 
        \round_in[0][394] , \round_in[0][393] , \round_in[0][392] , 
        \round_in[0][391] , \round_in[0][390] , \round_in[0][389] , 
        \round_in[0][388] , \round_in[0][387] , \round_in[0][386] , 
        \round_in[0][385] , \round_in[0][384] , \round_in[0][383] , 
        \round_in[0][382] , \round_in[0][381] , \round_in[0][380] , 
        \round_in[0][379] , \round_in[0][378] , \round_in[0][377] , 
        \round_in[0][376] , \round_in[0][375] , \round_in[0][374] , 
        \round_in[0][373] , \round_in[0][372] , \round_in[0][371] , 
        \round_in[0][370] , \round_in[0][369] , \round_in[0][368] , 
        \round_in[0][367] , \round_in[0][366] , \round_in[0][365] , 
        \round_in[0][364] , \round_in[0][363] , \round_in[0][362] , 
        \round_in[0][361] , \round_in[0][360] , \round_in[0][359] , 
        \round_in[0][358] , \round_in[0][357] , \round_in[0][356] , 
        \round_in[0][355] , \round_in[0][354] , \round_in[0][353] , 
        \round_in[0][352] , \round_in[0][351] , \round_in[0][350] , 
        \round_in[0][349] , \round_in[0][348] , \round_in[0][347] , 
        \round_in[0][346] , \round_in[0][345] , \round_in[0][344] , 
        \round_in[0][343] , \round_in[0][342] , \round_in[0][341] , 
        \round_in[0][340] , \round_in[0][339] , \round_in[0][338] , 
        \round_in[0][337] , \round_in[0][336] , \round_in[0][335] , 
        \round_in[0][334] , \round_in[0][333] , \round_in[0][332] , 
        \round_in[0][331] , \round_in[0][330] , \round_in[0][329] , 
        \round_in[0][328] , \round_in[0][327] , \round_in[0][326] , 
        \round_in[0][325] , \round_in[0][324] , \round_in[0][323] , 
        \round_in[0][322] , \round_in[0][321] , \round_in[0][320] , 
        \round_in[0][319] , \round_in[0][318] , \round_in[0][317] , 
        \round_in[0][316] , \round_in[0][315] , \round_in[0][314] , 
        \round_in[0][313] , \round_in[0][312] , \round_in[0][311] , 
        \round_in[0][310] , \round_in[0][309] , \round_in[0][308] , 
        \round_in[0][307] , \round_in[0][306] , \round_in[0][305] , 
        \round_in[0][304] , \round_in[0][303] , \round_in[0][302] , 
        \round_in[0][301] , \round_in[0][300] , \round_in[0][299] , 
        \round_in[0][298] , \round_in[0][297] , \round_in[0][296] , 
        \round_in[0][295] , \round_in[0][294] , \round_in[0][293] , 
        \round_in[0][292] , \round_in[0][291] , \round_in[0][290] , 
        \round_in[0][289] , \round_in[0][288] , \round_in[0][287] , 
        \round_in[0][286] , \round_in[0][285] , \round_in[0][284] , 
        \round_in[0][283] , \round_in[0][282] , \round_in[0][281] , 
        \round_in[0][280] , \round_in[0][279] , \round_in[0][278] , 
        \round_in[0][277] , \round_in[0][276] , \round_in[0][275] , 
        \round_in[0][274] , \round_in[0][273] , \round_in[0][272] , 
        \round_in[0][271] , \round_in[0][270] , \round_in[0][269] , 
        \round_in[0][268] , \round_in[0][267] , \round_in[0][266] , 
        \round_in[0][265] , \round_in[0][264] , \round_in[0][263] , 
        \round_in[0][262] , \round_in[0][261] , \round_in[0][260] , 
        \round_in[0][259] , \round_in[0][258] , \round_in[0][257] , 
        \round_in[0][256] , \round_in[0][255] , \round_in[0][254] , 
        \round_in[0][253] , \round_in[0][252] , \round_in[0][251] , 
        \round_in[0][250] , \round_in[0][249] , \round_in[0][248] , 
        \round_in[0][247] , \round_in[0][246] , \round_in[0][245] , 
        \round_in[0][244] , \round_in[0][243] , \round_in[0][242] , 
        \round_in[0][241] , \round_in[0][240] , \round_in[0][239] , 
        \round_in[0][238] , \round_in[0][237] , \round_in[0][236] , 
        \round_in[0][235] , \round_in[0][234] , \round_in[0][233] , 
        \round_in[0][232] , \round_in[0][231] , \round_in[0][230] , 
        \round_in[0][229] , \round_in[0][228] , \round_in[0][227] , 
        \round_in[0][226] , \round_in[0][225] , \round_in[0][224] , 
        \round_in[0][223] , \round_in[0][222] , \round_in[0][221] , 
        \round_in[0][220] , \round_in[0][219] , \round_in[0][218] , 
        \round_in[0][217] , \round_in[0][216] , \round_in[0][215] , 
        \round_in[0][214] , \round_in[0][213] , \round_in[0][212] , 
        \round_in[0][211] , \round_in[0][210] , \round_in[0][209] , 
        \round_in[0][208] , \round_in[0][207] , \round_in[0][206] , 
        \round_in[0][205] , \round_in[0][204] , \round_in[0][203] , 
        \round_in[0][202] , \round_in[0][201] , \round_in[0][200] , 
        \round_in[0][199] , \round_in[0][198] , \round_in[0][197] , 
        \round_in[0][196] , \round_in[0][195] , \round_in[0][194] , 
        \round_in[0][193] , \round_in[0][192] , \round_in[0][191] , 
        \round_in[0][190] , \round_in[0][189] , \round_in[0][188] , 
        \round_in[0][187] , \round_in[0][186] , \round_in[0][185] , 
        \round_in[0][184] , \round_in[0][183] , \round_in[0][182] , 
        \round_in[0][181] , \round_in[0][180] , \round_in[0][179] , 
        \round_in[0][178] , \round_in[0][177] , \round_in[0][176] , 
        \round_in[0][175] , \round_in[0][174] , \round_in[0][173] , 
        \round_in[0][172] , \round_in[0][171] , \round_in[0][170] , 
        \round_in[0][169] , \round_in[0][168] , \round_in[0][167] , 
        \round_in[0][166] , \round_in[0][165] , \round_in[0][164] , 
        \round_in[0][163] , \round_in[0][162] , \round_in[0][161] , 
        \round_in[0][160] , \round_in[0][159] , \round_in[0][158] , 
        \round_in[0][157] , \round_in[0][156] , \round_in[0][155] , 
        \round_in[0][154] , \round_in[0][153] , \round_in[0][152] , 
        \round_in[0][151] , \round_in[0][150] , \round_in[0][149] , 
        \round_in[0][148] , \round_in[0][147] , \round_in[0][146] , 
        \round_in[0][145] , \round_in[0][144] , \round_in[0][143] , 
        \round_in[0][142] , \round_in[0][141] , \round_in[0][140] , 
        \round_in[0][139] , \round_in[0][138] , \round_in[0][137] , 
        \round_in[0][136] , \round_in[0][135] , \round_in[0][134] , 
        \round_in[0][133] , \round_in[0][132] , \round_in[0][131] , 
        \round_in[0][130] , \round_in[0][129] , \round_in[0][128] , 
        \round_in[0][127] , \round_in[0][126] , \round_in[0][125] , 
        \round_in[0][124] , \round_in[0][123] , \round_in[0][122] , 
        \round_in[0][121] , \round_in[0][120] , \round_in[0][119] , 
        \round_in[0][118] , \round_in[0][117] , \round_in[0][116] , 
        \round_in[0][115] , \round_in[0][114] , \round_in[0][113] , 
        \round_in[0][112] , \round_in[0][111] , \round_in[0][110] , 
        \round_in[0][109] , \round_in[0][108] , \round_in[0][107] , 
        \round_in[0][106] , \round_in[0][105] , \round_in[0][104] , 
        \round_in[0][103] , \round_in[0][102] , \round_in[0][101] , 
        \round_in[0][100] , \round_in[0][99] , \round_in[0][98] , 
        \round_in[0][97] , \round_in[0][96] , \round_in[0][95] , 
        \round_in[0][94] , \round_in[0][93] , \round_in[0][92] , 
        \round_in[0][91] , \round_in[0][90] , \round_in[0][89] , 
        \round_in[0][88] , \round_in[0][87] , \round_in[0][86] , 
        \round_in[0][85] , \round_in[0][84] , \round_in[0][83] , 
        \round_in[0][82] , \round_in[0][81] , \round_in[0][80] , 
        \round_in[0][79] , \round_in[0][78] , \round_in[0][77] , 
        \round_in[0][76] , \round_in[0][75] , \round_in[0][74] , 
        \round_in[0][73] , \round_in[0][72] , \round_in[0][71] , 
        \round_in[0][70] , \round_in[0][69] , \round_in[0][68] , 
        \round_in[0][67] , \round_in[0][66] , \round_in[0][65] , 
        \round_in[0][64] , \round_in[0][63] , \round_in[0][62] , 
        \round_in[0][61] , \round_in[0][60] , \round_in[0][59] , 
        \round_in[0][58] , \round_in[0][57] , \round_in[0][56] , 
        \round_in[0][55] , \round_in[0][54] , \round_in[0][53] , 
        \round_in[0][52] , \round_in[0][51] , \round_in[0][50] , 
        \round_in[0][49] , \round_in[0][48] , \round_in[0][47] , 
        \round_in[0][46] , \round_in[0][45] , \round_in[0][44] , 
        \round_in[0][43] , \round_in[0][42] , \round_in[0][41] , 
        \round_in[0][40] , \round_in[0][39] , \round_in[0][38] , 
        \round_in[0][37] , \round_in[0][36] , \round_in[0][35] , 
        \round_in[0][34] , \round_in[0][33] , \round_in[0][32] , 
        \round_in[0][31] , \round_in[0][30] , \round_in[0][29] , 
        \round_in[0][28] , \round_in[0][27] , \round_in[0][26] , 
        \round_in[0][25] , \round_in[0][24] , \round_in[0][23] , 
        \round_in[0][22] , \round_in[0][21] , \round_in[0][20] , 
        \round_in[0][19] , \round_in[0][18] , \round_in[0][17] , 
        \round_in[0][16] , \round_in[0][15] , \round_in[0][14] , 
        \round_in[0][13] , \round_in[0][12] , \round_in[0][11] , 
        \round_in[0][10] , \round_in[0][9] , \round_in[0][8] , 
        \round_in[0][7] , \round_in[0][6] , \round_in[0][5] , \round_in[0][4] , 
        \round_in[0][3] , \round_in[0][2] , \round_in[0][1] , \round_in[0][0] }), .round_const({\RCONST[0].rconst_/N67 , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, \RCONST[0].rconst_/N56 , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        \RCONST[0].rconst_/N48 , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        \rc[2][0] , 1'b0, 1'b0, 1'b0, \RCONST[0].rconst_/N25 , 1'b0, 
        \RCONST[0].rconst_/N17 , \rc[3][15] }), .out({\round_in[1][1599] , 
        \round_in[1][1598] , \round_in[1][1597] , \round_in[1][1596] , 
        \round_in[1][1595] , \round_in[1][1594] , \round_in[1][1593] , 
        \round_in[1][1592] , \round_in[1][1591] , \round_in[1][1590] , 
        \round_in[1][1589] , \round_in[1][1588] , \round_in[1][1587] , 
        \round_in[1][1586] , \round_in[1][1585] , \round_in[1][1584] , 
        \round_in[1][1583] , \round_in[1][1582] , \round_in[1][1581] , 
        \round_in[1][1580] , \round_in[1][1579] , \round_in[1][1578] , 
        \round_in[1][1577] , \round_in[1][1576] , \round_in[1][1575] , 
        \round_in[1][1574] , \round_in[1][1573] , \round_in[1][1572] , 
        \round_in[1][1571] , \round_in[1][1570] , \round_in[1][1569] , 
        \round_in[1][1568] , \round_in[1][1567] , \round_in[1][1566] , 
        \round_in[1][1565] , \round_in[1][1564] , \round_in[1][1563] , 
        \round_in[1][1562] , \round_in[1][1561] , \round_in[1][1560] , 
        \round_in[1][1559] , \round_in[1][1558] , \round_in[1][1557] , 
        \round_in[1][1556] , \round_in[1][1555] , \round_in[1][1554] , 
        \round_in[1][1553] , \round_in[1][1552] , \round_in[1][1551] , 
        \round_in[1][1550] , \round_in[1][1549] , \round_in[1][1548] , 
        \round_in[1][1547] , \round_in[1][1546] , \round_in[1][1545] , 
        \round_in[1][1544] , \round_in[1][1543] , \round_in[1][1542] , 
        \round_in[1][1541] , \round_in[1][1540] , \round_in[1][1539] , 
        \round_in[1][1538] , \round_in[1][1537] , \round_in[1][1536] , 
        \round_in[1][1535] , \round_in[1][1534] , \round_in[1][1533] , 
        \round_in[1][1532] , \round_in[1][1531] , \round_in[1][1530] , 
        \round_in[1][1529] , \round_in[1][1528] , \round_in[1][1527] , 
        \round_in[1][1526] , \round_in[1][1525] , \round_in[1][1524] , 
        \round_in[1][1523] , \round_in[1][1522] , \round_in[1][1521] , 
        \round_in[1][1520] , \round_in[1][1519] , \round_in[1][1518] , 
        \round_in[1][1517] , \round_in[1][1516] , \round_in[1][1515] , 
        \round_in[1][1514] , \round_in[1][1513] , \round_in[1][1512] , 
        \round_in[1][1511] , \round_in[1][1510] , \round_in[1][1509] , 
        \round_in[1][1508] , \round_in[1][1507] , \round_in[1][1506] , 
        \round_in[1][1505] , \round_in[1][1504] , \round_in[1][1503] , 
        \round_in[1][1502] , \round_in[1][1501] , \round_in[1][1500] , 
        \round_in[1][1499] , \round_in[1][1498] , \round_in[1][1497] , 
        \round_in[1][1496] , \round_in[1][1495] , \round_in[1][1494] , 
        \round_in[1][1493] , \round_in[1][1492] , \round_in[1][1491] , 
        \round_in[1][1490] , \round_in[1][1489] , \round_in[1][1488] , 
        \round_in[1][1487] , \round_in[1][1486] , \round_in[1][1485] , 
        \round_in[1][1484] , \round_in[1][1483] , \round_in[1][1482] , 
        \round_in[1][1481] , \round_in[1][1480] , \round_in[1][1479] , 
        \round_in[1][1478] , \round_in[1][1477] , \round_in[1][1476] , 
        \round_in[1][1475] , \round_in[1][1474] , \round_in[1][1473] , 
        \round_in[1][1472] , \round_in[1][1471] , \round_in[1][1470] , 
        \round_in[1][1469] , \round_in[1][1468] , \round_in[1][1467] , 
        \round_in[1][1466] , \round_in[1][1465] , \round_in[1][1464] , 
        \round_in[1][1463] , \round_in[1][1462] , \round_in[1][1461] , 
        \round_in[1][1460] , \round_in[1][1459] , \round_in[1][1458] , 
        \round_in[1][1457] , \round_in[1][1456] , \round_in[1][1455] , 
        \round_in[1][1454] , \round_in[1][1453] , \round_in[1][1452] , 
        \round_in[1][1451] , \round_in[1][1450] , \round_in[1][1449] , 
        \round_in[1][1448] , \round_in[1][1447] , \round_in[1][1446] , 
        \round_in[1][1445] , \round_in[1][1444] , \round_in[1][1443] , 
        \round_in[1][1442] , \round_in[1][1441] , \round_in[1][1440] , 
        \round_in[1][1439] , \round_in[1][1438] , \round_in[1][1437] , 
        \round_in[1][1436] , \round_in[1][1435] , \round_in[1][1434] , 
        \round_in[1][1433] , \round_in[1][1432] , \round_in[1][1431] , 
        \round_in[1][1430] , \round_in[1][1429] , \round_in[1][1428] , 
        \round_in[1][1427] , \round_in[1][1426] , \round_in[1][1425] , 
        \round_in[1][1424] , \round_in[1][1423] , \round_in[1][1422] , 
        \round_in[1][1421] , \round_in[1][1420] , \round_in[1][1419] , 
        \round_in[1][1418] , \round_in[1][1417] , \round_in[1][1416] , 
        \round_in[1][1415] , \round_in[1][1414] , \round_in[1][1413] , 
        \round_in[1][1412] , \round_in[1][1411] , \round_in[1][1410] , 
        \round_in[1][1409] , \round_in[1][1408] , \round_in[1][1407] , 
        \round_in[1][1406] , \round_in[1][1405] , \round_in[1][1404] , 
        \round_in[1][1403] , \round_in[1][1402] , \round_in[1][1401] , 
        \round_in[1][1400] , \round_in[1][1399] , \round_in[1][1398] , 
        \round_in[1][1397] , \round_in[1][1396] , \round_in[1][1395] , 
        \round_in[1][1394] , \round_in[1][1393] , \round_in[1][1392] , 
        \round_in[1][1391] , \round_in[1][1390] , \round_in[1][1389] , 
        \round_in[1][1388] , \round_in[1][1387] , \round_in[1][1386] , 
        \round_in[1][1385] , \round_in[1][1384] , \round_in[1][1383] , 
        \round_in[1][1382] , \round_in[1][1381] , \round_in[1][1380] , 
        \round_in[1][1379] , \round_in[1][1378] , \round_in[1][1377] , 
        \round_in[1][1376] , \round_in[1][1375] , \round_in[1][1374] , 
        \round_in[1][1373] , \round_in[1][1372] , \round_in[1][1371] , 
        \round_in[1][1370] , \round_in[1][1369] , \round_in[1][1368] , 
        \round_in[1][1367] , \round_in[1][1366] , \round_in[1][1365] , 
        \round_in[1][1364] , \round_in[1][1363] , \round_in[1][1362] , 
        \round_in[1][1361] , \round_in[1][1360] , \round_in[1][1359] , 
        \round_in[1][1358] , \round_in[1][1357] , \round_in[1][1356] , 
        \round_in[1][1355] , \round_in[1][1354] , \round_in[1][1353] , 
        \round_in[1][1352] , \round_in[1][1351] , \round_in[1][1350] , 
        \round_in[1][1349] , \round_in[1][1348] , \round_in[1][1347] , 
        \round_in[1][1346] , \round_in[1][1345] , \round_in[1][1344] , 
        \round_in[1][1343] , \round_in[1][1342] , \round_in[1][1341] , 
        \round_in[1][1340] , \round_in[1][1339] , \round_in[1][1338] , 
        \round_in[1][1337] , \round_in[1][1336] , \round_in[1][1335] , 
        \round_in[1][1334] , \round_in[1][1333] , \round_in[1][1332] , 
        \round_in[1][1331] , \round_in[1][1330] , \round_in[1][1329] , 
        \round_in[1][1328] , \round_in[1][1327] , \round_in[1][1326] , 
        \round_in[1][1325] , \round_in[1][1324] , \round_in[1][1323] , 
        \round_in[1][1322] , \round_in[1][1321] , \round_in[1][1320] , 
        \round_in[1][1319] , \round_in[1][1318] , \round_in[1][1317] , 
        \round_in[1][1316] , \round_in[1][1315] , \round_in[1][1314] , 
        \round_in[1][1313] , \round_in[1][1312] , \round_in[1][1311] , 
        \round_in[1][1310] , \round_in[1][1309] , \round_in[1][1308] , 
        \round_in[1][1307] , \round_in[1][1306] , \round_in[1][1305] , 
        \round_in[1][1304] , \round_in[1][1303] , \round_in[1][1302] , 
        \round_in[1][1301] , \round_in[1][1300] , \round_in[1][1299] , 
        \round_in[1][1298] , \round_in[1][1297] , \round_in[1][1296] , 
        \round_in[1][1295] , \round_in[1][1294] , \round_in[1][1293] , 
        \round_in[1][1292] , \round_in[1][1291] , \round_in[1][1290] , 
        \round_in[1][1289] , \round_in[1][1288] , \round_in[1][1287] , 
        \round_in[1][1286] , \round_in[1][1285] , \round_in[1][1284] , 
        \round_in[1][1283] , \round_in[1][1282] , \round_in[1][1281] , 
        \round_in[1][1280] , \round_in[1][1279] , \round_in[1][1278] , 
        \round_in[1][1277] , \round_in[1][1276] , \round_in[1][1275] , 
        \round_in[1][1274] , \round_in[1][1273] , \round_in[1][1272] , 
        \round_in[1][1271] , \round_in[1][1270] , \round_in[1][1269] , 
        \round_in[1][1268] , \round_in[1][1267] , \round_in[1][1266] , 
        \round_in[1][1265] , \round_in[1][1264] , \round_in[1][1263] , 
        \round_in[1][1262] , \round_in[1][1261] , \round_in[1][1260] , 
        \round_in[1][1259] , \round_in[1][1258] , \round_in[1][1257] , 
        \round_in[1][1256] , \round_in[1][1255] , \round_in[1][1254] , 
        \round_in[1][1253] , \round_in[1][1252] , \round_in[1][1251] , 
        \round_in[1][1250] , \round_in[1][1249] , \round_in[1][1248] , 
        \round_in[1][1247] , \round_in[1][1246] , \round_in[1][1245] , 
        \round_in[1][1244] , \round_in[1][1243] , \round_in[1][1242] , 
        \round_in[1][1241] , \round_in[1][1240] , \round_in[1][1239] , 
        \round_in[1][1238] , \round_in[1][1237] , \round_in[1][1236] , 
        \round_in[1][1235] , \round_in[1][1234] , \round_in[1][1233] , 
        \round_in[1][1232] , \round_in[1][1231] , \round_in[1][1230] , 
        \round_in[1][1229] , \round_in[1][1228] , \round_in[1][1227] , 
        \round_in[1][1226] , \round_in[1][1225] , \round_in[1][1224] , 
        \round_in[1][1223] , \round_in[1][1222] , \round_in[1][1221] , 
        \round_in[1][1220] , \round_in[1][1219] , \round_in[1][1218] , 
        \round_in[1][1217] , \round_in[1][1216] , \round_in[1][1215] , 
        \round_in[1][1214] , \round_in[1][1213] , \round_in[1][1212] , 
        \round_in[1][1211] , \round_in[1][1210] , \round_in[1][1209] , 
        \round_in[1][1208] , \round_in[1][1207] , \round_in[1][1206] , 
        \round_in[1][1205] , \round_in[1][1204] , \round_in[1][1203] , 
        \round_in[1][1202] , \round_in[1][1201] , \round_in[1][1200] , 
        \round_in[1][1199] , \round_in[1][1198] , \round_in[1][1197] , 
        \round_in[1][1196] , \round_in[1][1195] , \round_in[1][1194] , 
        \round_in[1][1193] , \round_in[1][1192] , \round_in[1][1191] , 
        \round_in[1][1190] , \round_in[1][1189] , \round_in[1][1188] , 
        \round_in[1][1187] , \round_in[1][1186] , \round_in[1][1185] , 
        \round_in[1][1184] , \round_in[1][1183] , \round_in[1][1182] , 
        \round_in[1][1181] , \round_in[1][1180] , \round_in[1][1179] , 
        \round_in[1][1178] , \round_in[1][1177] , \round_in[1][1176] , 
        \round_in[1][1175] , \round_in[1][1174] , \round_in[1][1173] , 
        \round_in[1][1172] , \round_in[1][1171] , \round_in[1][1170] , 
        \round_in[1][1169] , \round_in[1][1168] , \round_in[1][1167] , 
        \round_in[1][1166] , \round_in[1][1165] , \round_in[1][1164] , 
        \round_in[1][1163] , \round_in[1][1162] , \round_in[1][1161] , 
        \round_in[1][1160] , \round_in[1][1159] , \round_in[1][1158] , 
        \round_in[1][1157] , \round_in[1][1156] , \round_in[1][1155] , 
        \round_in[1][1154] , \round_in[1][1153] , \round_in[1][1152] , 
        \round_in[1][1151] , \round_in[1][1150] , \round_in[1][1149] , 
        \round_in[1][1148] , \round_in[1][1147] , \round_in[1][1146] , 
        \round_in[1][1145] , \round_in[1][1144] , \round_in[1][1143] , 
        \round_in[1][1142] , \round_in[1][1141] , \round_in[1][1140] , 
        \round_in[1][1139] , \round_in[1][1138] , \round_in[1][1137] , 
        \round_in[1][1136] , \round_in[1][1135] , \round_in[1][1134] , 
        \round_in[1][1133] , \round_in[1][1132] , \round_in[1][1131] , 
        \round_in[1][1130] , \round_in[1][1129] , \round_in[1][1128] , 
        \round_in[1][1127] , \round_in[1][1126] , \round_in[1][1125] , 
        \round_in[1][1124] , \round_in[1][1123] , \round_in[1][1122] , 
        \round_in[1][1121] , \round_in[1][1120] , \round_in[1][1119] , 
        \round_in[1][1118] , \round_in[1][1117] , \round_in[1][1116] , 
        \round_in[1][1115] , \round_in[1][1114] , \round_in[1][1113] , 
        \round_in[1][1112] , \round_in[1][1111] , \round_in[1][1110] , 
        \round_in[1][1109] , \round_in[1][1108] , \round_in[1][1107] , 
        \round_in[1][1106] , \round_in[1][1105] , \round_in[1][1104] , 
        \round_in[1][1103] , \round_in[1][1102] , \round_in[1][1101] , 
        \round_in[1][1100] , \round_in[1][1099] , \round_in[1][1098] , 
        \round_in[1][1097] , \round_in[1][1096] , \round_in[1][1095] , 
        \round_in[1][1094] , \round_in[1][1093] , \round_in[1][1092] , 
        \round_in[1][1091] , \round_in[1][1090] , \round_in[1][1089] , 
        \round_in[1][1088] , \round_in[1][1087] , \round_in[1][1086] , 
        \round_in[1][1085] , \round_in[1][1084] , \round_in[1][1083] , 
        \round_in[1][1082] , \round_in[1][1081] , \round_in[1][1080] , 
        \round_in[1][1079] , \round_in[1][1078] , \round_in[1][1077] , 
        \round_in[1][1076] , \round_in[1][1075] , \round_in[1][1074] , 
        \round_in[1][1073] , \round_in[1][1072] , \round_in[1][1071] , 
        \round_in[1][1070] , \round_in[1][1069] , \round_in[1][1068] , 
        \round_in[1][1067] , \round_in[1][1066] , \round_in[1][1065] , 
        \round_in[1][1064] , \round_in[1][1063] , \round_in[1][1062] , 
        \round_in[1][1061] , \round_in[1][1060] , \round_in[1][1059] , 
        \round_in[1][1058] , \round_in[1][1057] , \round_in[1][1056] , 
        \round_in[1][1055] , \round_in[1][1054] , \round_in[1][1053] , 
        \round_in[1][1052] , \round_in[1][1051] , \round_in[1][1050] , 
        \round_in[1][1049] , \round_in[1][1048] , \round_in[1][1047] , 
        \round_in[1][1046] , \round_in[1][1045] , \round_in[1][1044] , 
        \round_in[1][1043] , \round_in[1][1042] , \round_in[1][1041] , 
        \round_in[1][1040] , \round_in[1][1039] , \round_in[1][1038] , 
        \round_in[1][1037] , \round_in[1][1036] , \round_in[1][1035] , 
        \round_in[1][1034] , \round_in[1][1033] , \round_in[1][1032] , 
        \round_in[1][1031] , \round_in[1][1030] , \round_in[1][1029] , 
        \round_in[1][1028] , \round_in[1][1027] , \round_in[1][1026] , 
        \round_in[1][1025] , \round_in[1][1024] , \round_in[1][1023] , 
        \round_in[1][1022] , \round_in[1][1021] , \round_in[1][1020] , 
        \round_in[1][1019] , \round_in[1][1018] , \round_in[1][1017] , 
        \round_in[1][1016] , \round_in[1][1015] , \round_in[1][1014] , 
        \round_in[1][1013] , \round_in[1][1012] , \round_in[1][1011] , 
        \round_in[1][1010] , \round_in[1][1009] , \round_in[1][1008] , 
        \round_in[1][1007] , \round_in[1][1006] , \round_in[1][1005] , 
        \round_in[1][1004] , \round_in[1][1003] , \round_in[1][1002] , 
        \round_in[1][1001] , \round_in[1][1000] , \round_in[1][999] , 
        \round_in[1][998] , \round_in[1][997] , \round_in[1][996] , 
        \round_in[1][995] , \round_in[1][994] , \round_in[1][993] , 
        \round_in[1][992] , \round_in[1][991] , \round_in[1][990] , 
        \round_in[1][989] , \round_in[1][988] , \round_in[1][987] , 
        \round_in[1][986] , \round_in[1][985] , \round_in[1][984] , 
        \round_in[1][983] , \round_in[1][982] , \round_in[1][981] , 
        \round_in[1][980] , \round_in[1][979] , \round_in[1][978] , 
        \round_in[1][977] , \round_in[1][976] , \round_in[1][975] , 
        \round_in[1][974] , \round_in[1][973] , \round_in[1][972] , 
        \round_in[1][971] , \round_in[1][970] , \round_in[1][969] , 
        \round_in[1][968] , \round_in[1][967] , \round_in[1][966] , 
        \round_in[1][965] , \round_in[1][964] , \round_in[1][963] , 
        \round_in[1][962] , \round_in[1][961] , \round_in[1][960] , 
        \round_in[1][959] , \round_in[1][958] , \round_in[1][957] , 
        \round_in[1][956] , \round_in[1][955] , \round_in[1][954] , 
        \round_in[1][953] , \round_in[1][952] , \round_in[1][951] , 
        \round_in[1][950] , \round_in[1][949] , \round_in[1][948] , 
        \round_in[1][947] , \round_in[1][946] , \round_in[1][945] , 
        \round_in[1][944] , \round_in[1][943] , \round_in[1][942] , 
        \round_in[1][941] , \round_in[1][940] , \round_in[1][939] , 
        \round_in[1][938] , \round_in[1][937] , \round_in[1][936] , 
        \round_in[1][935] , \round_in[1][934] , \round_in[1][933] , 
        \round_in[1][932] , \round_in[1][931] , \round_in[1][930] , 
        \round_in[1][929] , \round_in[1][928] , \round_in[1][927] , 
        \round_in[1][926] , \round_in[1][925] , \round_in[1][924] , 
        \round_in[1][923] , \round_in[1][922] , \round_in[1][921] , 
        \round_in[1][920] , \round_in[1][919] , \round_in[1][918] , 
        \round_in[1][917] , \round_in[1][916] , \round_in[1][915] , 
        \round_in[1][914] , \round_in[1][913] , \round_in[1][912] , 
        \round_in[1][911] , \round_in[1][910] , \round_in[1][909] , 
        \round_in[1][908] , \round_in[1][907] , \round_in[1][906] , 
        \round_in[1][905] , \round_in[1][904] , \round_in[1][903] , 
        \round_in[1][902] , \round_in[1][901] , \round_in[1][900] , 
        \round_in[1][899] , \round_in[1][898] , \round_in[1][897] , 
        \round_in[1][896] , \round_in[1][895] , \round_in[1][894] , 
        \round_in[1][893] , \round_in[1][892] , \round_in[1][891] , 
        \round_in[1][890] , \round_in[1][889] , \round_in[1][888] , 
        \round_in[1][887] , \round_in[1][886] , \round_in[1][885] , 
        \round_in[1][884] , \round_in[1][883] , \round_in[1][882] , 
        \round_in[1][881] , \round_in[1][880] , \round_in[1][879] , 
        \round_in[1][878] , \round_in[1][877] , \round_in[1][876] , 
        \round_in[1][875] , \round_in[1][874] , \round_in[1][873] , 
        \round_in[1][872] , \round_in[1][871] , \round_in[1][870] , 
        \round_in[1][869] , \round_in[1][868] , \round_in[1][867] , 
        \round_in[1][866] , \round_in[1][865] , \round_in[1][864] , 
        \round_in[1][863] , \round_in[1][862] , \round_in[1][861] , 
        \round_in[1][860] , \round_in[1][859] , \round_in[1][858] , 
        \round_in[1][857] , \round_in[1][856] , \round_in[1][855] , 
        \round_in[1][854] , \round_in[1][853] , \round_in[1][852] , 
        \round_in[1][851] , \round_in[1][850] , \round_in[1][849] , 
        \round_in[1][848] , \round_in[1][847] , \round_in[1][846] , 
        \round_in[1][845] , \round_in[1][844] , \round_in[1][843] , 
        \round_in[1][842] , \round_in[1][841] , \round_in[1][840] , 
        \round_in[1][839] , \round_in[1][838] , \round_in[1][837] , 
        \round_in[1][836] , \round_in[1][835] , \round_in[1][834] , 
        \round_in[1][833] , \round_in[1][832] , \round_in[1][831] , 
        \round_in[1][830] , \round_in[1][829] , \round_in[1][828] , 
        \round_in[1][827] , \round_in[1][826] , \round_in[1][825] , 
        \round_in[1][824] , \round_in[1][823] , \round_in[1][822] , 
        \round_in[1][821] , \round_in[1][820] , \round_in[1][819] , 
        \round_in[1][818] , \round_in[1][817] , \round_in[1][816] , 
        \round_in[1][815] , \round_in[1][814] , \round_in[1][813] , 
        \round_in[1][812] , \round_in[1][811] , \round_in[1][810] , 
        \round_in[1][809] , \round_in[1][808] , \round_in[1][807] , 
        \round_in[1][806] , \round_in[1][805] , \round_in[1][804] , 
        \round_in[1][803] , \round_in[1][802] , \round_in[1][801] , 
        \round_in[1][800] , \round_in[1][799] , \round_in[1][798] , 
        \round_in[1][797] , \round_in[1][796] , \round_in[1][795] , 
        \round_in[1][794] , \round_in[1][793] , \round_in[1][792] , 
        \round_in[1][791] , \round_in[1][790] , \round_in[1][789] , 
        \round_in[1][788] , \round_in[1][787] , \round_in[1][786] , 
        \round_in[1][785] , \round_in[1][784] , \round_in[1][783] , 
        \round_in[1][782] , \round_in[1][781] , \round_in[1][780] , 
        \round_in[1][779] , \round_in[1][778] , \round_in[1][777] , 
        \round_in[1][776] , \round_in[1][775] , \round_in[1][774] , 
        \round_in[1][773] , \round_in[1][772] , \round_in[1][771] , 
        \round_in[1][770] , \round_in[1][769] , \round_in[1][768] , 
        \round_in[1][767] , \round_in[1][766] , \round_in[1][765] , 
        \round_in[1][764] , \round_in[1][763] , \round_in[1][762] , 
        \round_in[1][761] , \round_in[1][760] , \round_in[1][759] , 
        \round_in[1][758] , \round_in[1][757] , \round_in[1][756] , 
        \round_in[1][755] , \round_in[1][754] , \round_in[1][753] , 
        \round_in[1][752] , \round_in[1][751] , \round_in[1][750] , 
        \round_in[1][749] , \round_in[1][748] , \round_in[1][747] , 
        \round_in[1][746] , \round_in[1][745] , \round_in[1][744] , 
        \round_in[1][743] , \round_in[1][742] , \round_in[1][741] , 
        \round_in[1][740] , \round_in[1][739] , \round_in[1][738] , 
        \round_in[1][737] , \round_in[1][736] , \round_in[1][735] , 
        \round_in[1][734] , \round_in[1][733] , \round_in[1][732] , 
        \round_in[1][731] , \round_in[1][730] , \round_in[1][729] , 
        \round_in[1][728] , \round_in[1][727] , \round_in[1][726] , 
        \round_in[1][725] , \round_in[1][724] , \round_in[1][723] , 
        \round_in[1][722] , \round_in[1][721] , \round_in[1][720] , 
        \round_in[1][719] , \round_in[1][718] , \round_in[1][717] , 
        \round_in[1][716] , \round_in[1][715] , \round_in[1][714] , 
        \round_in[1][713] , \round_in[1][712] , \round_in[1][711] , 
        \round_in[1][710] , \round_in[1][709] , \round_in[1][708] , 
        \round_in[1][707] , \round_in[1][706] , \round_in[1][705] , 
        \round_in[1][704] , \round_in[1][703] , \round_in[1][702] , 
        \round_in[1][701] , \round_in[1][700] , \round_in[1][699] , 
        \round_in[1][698] , \round_in[1][697] , \round_in[1][696] , 
        \round_in[1][695] , \round_in[1][694] , \round_in[1][693] , 
        \round_in[1][692] , \round_in[1][691] , \round_in[1][690] , 
        \round_in[1][689] , \round_in[1][688] , \round_in[1][687] , 
        \round_in[1][686] , \round_in[1][685] , \round_in[1][684] , 
        \round_in[1][683] , \round_in[1][682] , \round_in[1][681] , 
        \round_in[1][680] , \round_in[1][679] , \round_in[1][678] , 
        \round_in[1][677] , \round_in[1][676] , \round_in[1][675] , 
        \round_in[1][674] , \round_in[1][673] , \round_in[1][672] , 
        \round_in[1][671] , \round_in[1][670] , \round_in[1][669] , 
        \round_in[1][668] , \round_in[1][667] , \round_in[1][666] , 
        \round_in[1][665] , \round_in[1][664] , \round_in[1][663] , 
        \round_in[1][662] , \round_in[1][661] , \round_in[1][660] , 
        \round_in[1][659] , \round_in[1][658] , \round_in[1][657] , 
        \round_in[1][656] , \round_in[1][655] , \round_in[1][654] , 
        \round_in[1][653] , \round_in[1][652] , \round_in[1][651] , 
        \round_in[1][650] , \round_in[1][649] , \round_in[1][648] , 
        \round_in[1][647] , \round_in[1][646] , \round_in[1][645] , 
        \round_in[1][644] , \round_in[1][643] , \round_in[1][642] , 
        \round_in[1][641] , \round_in[1][640] , \round_in[1][639] , 
        \round_in[1][638] , \round_in[1][637] , \round_in[1][636] , 
        \round_in[1][635] , \round_in[1][634] , \round_in[1][633] , 
        \round_in[1][632] , \round_in[1][631] , \round_in[1][630] , 
        \round_in[1][629] , \round_in[1][628] , \round_in[1][627] , 
        \round_in[1][626] , \round_in[1][625] , \round_in[1][624] , 
        \round_in[1][623] , \round_in[1][622] , \round_in[1][621] , 
        \round_in[1][620] , \round_in[1][619] , \round_in[1][618] , 
        \round_in[1][617] , \round_in[1][616] , \round_in[1][615] , 
        \round_in[1][614] , \round_in[1][613] , \round_in[1][612] , 
        \round_in[1][611] , \round_in[1][610] , \round_in[1][609] , 
        \round_in[1][608] , \round_in[1][607] , \round_in[1][606] , 
        \round_in[1][605] , \round_in[1][604] , \round_in[1][603] , 
        \round_in[1][602] , \round_in[1][601] , \round_in[1][600] , 
        \round_in[1][599] , \round_in[1][598] , \round_in[1][597] , 
        \round_in[1][596] , \round_in[1][595] , \round_in[1][594] , 
        \round_in[1][593] , \round_in[1][592] , \round_in[1][591] , 
        \round_in[1][590] , \round_in[1][589] , \round_in[1][588] , 
        \round_in[1][587] , \round_in[1][586] , \round_in[1][585] , 
        \round_in[1][584] , \round_in[1][583] , \round_in[1][582] , 
        \round_in[1][581] , \round_in[1][580] , \round_in[1][579] , 
        \round_in[1][578] , \round_in[1][577] , \round_in[1][576] , 
        \round_in[1][575] , \round_in[1][574] , \round_in[1][573] , 
        \round_in[1][572] , \round_in[1][571] , \round_in[1][570] , 
        \round_in[1][569] , \round_in[1][568] , \round_in[1][567] , 
        \round_in[1][566] , \round_in[1][565] , \round_in[1][564] , 
        \round_in[1][563] , \round_in[1][562] , \round_in[1][561] , 
        \round_in[1][560] , \round_in[1][559] , \round_in[1][558] , 
        \round_in[1][557] , \round_in[1][556] , \round_in[1][555] , 
        \round_in[1][554] , \round_in[1][553] , \round_in[1][552] , 
        \round_in[1][551] , \round_in[1][550] , \round_in[1][549] , 
        \round_in[1][548] , \round_in[1][547] , \round_in[1][546] , 
        \round_in[1][545] , \round_in[1][544] , \round_in[1][543] , 
        \round_in[1][542] , \round_in[1][541] , \round_in[1][540] , 
        \round_in[1][539] , \round_in[1][538] , \round_in[1][537] , 
        \round_in[1][536] , \round_in[1][535] , \round_in[1][534] , 
        \round_in[1][533] , \round_in[1][532] , \round_in[1][531] , 
        \round_in[1][530] , \round_in[1][529] , \round_in[1][528] , 
        \round_in[1][527] , \round_in[1][526] , \round_in[1][525] , 
        \round_in[1][524] , \round_in[1][523] , \round_in[1][522] , 
        \round_in[1][521] , \round_in[1][520] , \round_in[1][519] , 
        \round_in[1][518] , \round_in[1][517] , \round_in[1][516] , 
        \round_in[1][515] , \round_in[1][514] , \round_in[1][513] , 
        \round_in[1][512] , \round_in[1][511] , \round_in[1][510] , 
        \round_in[1][509] , \round_in[1][508] , \round_in[1][507] , 
        \round_in[1][506] , \round_in[1][505] , \round_in[1][504] , 
        \round_in[1][503] , \round_in[1][502] , \round_in[1][501] , 
        \round_in[1][500] , \round_in[1][499] , \round_in[1][498] , 
        \round_in[1][497] , \round_in[1][496] , \round_in[1][495] , 
        \round_in[1][494] , \round_in[1][493] , \round_in[1][492] , 
        \round_in[1][491] , \round_in[1][490] , \round_in[1][489] , 
        \round_in[1][488] , \round_in[1][487] , \round_in[1][486] , 
        \round_in[1][485] , \round_in[1][484] , \round_in[1][483] , 
        \round_in[1][482] , \round_in[1][481] , \round_in[1][480] , 
        \round_in[1][479] , \round_in[1][478] , \round_in[1][477] , 
        \round_in[1][476] , \round_in[1][475] , \round_in[1][474] , 
        \round_in[1][473] , \round_in[1][472] , \round_in[1][471] , 
        \round_in[1][470] , \round_in[1][469] , \round_in[1][468] , 
        \round_in[1][467] , \round_in[1][466] , \round_in[1][465] , 
        \round_in[1][464] , \round_in[1][463] , \round_in[1][462] , 
        \round_in[1][461] , \round_in[1][460] , \round_in[1][459] , 
        \round_in[1][458] , \round_in[1][457] , \round_in[1][456] , 
        \round_in[1][455] , \round_in[1][454] , \round_in[1][453] , 
        \round_in[1][452] , \round_in[1][451] , \round_in[1][450] , 
        \round_in[1][449] , \round_in[1][448] , \round_in[1][447] , 
        \round_in[1][446] , \round_in[1][445] , \round_in[1][444] , 
        \round_in[1][443] , \round_in[1][442] , \round_in[1][441] , 
        \round_in[1][440] , \round_in[1][439] , \round_in[1][438] , 
        \round_in[1][437] , \round_in[1][436] , \round_in[1][435] , 
        \round_in[1][434] , \round_in[1][433] , \round_in[1][432] , 
        \round_in[1][431] , \round_in[1][430] , \round_in[1][429] , 
        \round_in[1][428] , \round_in[1][427] , \round_in[1][426] , 
        \round_in[1][425] , \round_in[1][424] , \round_in[1][423] , 
        \round_in[1][422] , \round_in[1][421] , \round_in[1][420] , 
        \round_in[1][419] , \round_in[1][418] , \round_in[1][417] , 
        \round_in[1][416] , \round_in[1][415] , \round_in[1][414] , 
        \round_in[1][413] , \round_in[1][412] , \round_in[1][411] , 
        \round_in[1][410] , \round_in[1][409] , \round_in[1][408] , 
        \round_in[1][407] , \round_in[1][406] , \round_in[1][405] , 
        \round_in[1][404] , \round_in[1][403] , \round_in[1][402] , 
        \round_in[1][401] , \round_in[1][400] , \round_in[1][399] , 
        \round_in[1][398] , \round_in[1][397] , \round_in[1][396] , 
        \round_in[1][395] , \round_in[1][394] , \round_in[1][393] , 
        \round_in[1][392] , \round_in[1][391] , \round_in[1][390] , 
        \round_in[1][389] , \round_in[1][388] , \round_in[1][387] , 
        \round_in[1][386] , \round_in[1][385] , \round_in[1][384] , 
        \round_in[1][383] , \round_in[1][382] , \round_in[1][381] , 
        \round_in[1][380] , \round_in[1][379] , \round_in[1][378] , 
        \round_in[1][377] , \round_in[1][376] , \round_in[1][375] , 
        \round_in[1][374] , \round_in[1][373] , \round_in[1][372] , 
        \round_in[1][371] , \round_in[1][370] , \round_in[1][369] , 
        \round_in[1][368] , \round_in[1][367] , \round_in[1][366] , 
        \round_in[1][365] , \round_in[1][364] , \round_in[1][363] , 
        \round_in[1][362] , \round_in[1][361] , \round_in[1][360] , 
        \round_in[1][359] , \round_in[1][358] , \round_in[1][357] , 
        \round_in[1][356] , \round_in[1][355] , \round_in[1][354] , 
        \round_in[1][353] , \round_in[1][352] , \round_in[1][351] , 
        \round_in[1][350] , \round_in[1][349] , \round_in[1][348] , 
        \round_in[1][347] , \round_in[1][346] , \round_in[1][345] , 
        \round_in[1][344] , \round_in[1][343] , \round_in[1][342] , 
        \round_in[1][341] , \round_in[1][340] , \round_in[1][339] , 
        \round_in[1][338] , \round_in[1][337] , \round_in[1][336] , 
        \round_in[1][335] , \round_in[1][334] , \round_in[1][333] , 
        \round_in[1][332] , \round_in[1][331] , \round_in[1][330] , 
        \round_in[1][329] , \round_in[1][328] , \round_in[1][327] , 
        \round_in[1][326] , \round_in[1][325] , \round_in[1][324] , 
        \round_in[1][323] , \round_in[1][322] , \round_in[1][321] , 
        \round_in[1][320] , \round_in[1][319] , \round_in[1][318] , 
        \round_in[1][317] , \round_in[1][316] , \round_in[1][315] , 
        \round_in[1][314] , \round_in[1][313] , \round_in[1][312] , 
        \round_in[1][311] , \round_in[1][310] , \round_in[1][309] , 
        \round_in[1][308] , \round_in[1][307] , \round_in[1][306] , 
        \round_in[1][305] , \round_in[1][304] , \round_in[1][303] , 
        \round_in[1][302] , \round_in[1][301] , \round_in[1][300] , 
        \round_in[1][299] , \round_in[1][298] , \round_in[1][297] , 
        \round_in[1][296] , \round_in[1][295] , \round_in[1][294] , 
        \round_in[1][293] , \round_in[1][292] , \round_in[1][291] , 
        \round_in[1][290] , \round_in[1][289] , \round_in[1][288] , 
        \round_in[1][287] , \round_in[1][286] , \round_in[1][285] , 
        \round_in[1][284] , \round_in[1][283] , \round_in[1][282] , 
        \round_in[1][281] , \round_in[1][280] , \round_in[1][279] , 
        \round_in[1][278] , \round_in[1][277] , \round_in[1][276] , 
        \round_in[1][275] , \round_in[1][274] , \round_in[1][273] , 
        \round_in[1][272] , \round_in[1][271] , \round_in[1][270] , 
        \round_in[1][269] , \round_in[1][268] , \round_in[1][267] , 
        \round_in[1][266] , \round_in[1][265] , \round_in[1][264] , 
        \round_in[1][263] , \round_in[1][262] , \round_in[1][261] , 
        \round_in[1][260] , \round_in[1][259] , \round_in[1][258] , 
        \round_in[1][257] , \round_in[1][256] , \round_in[1][255] , 
        \round_in[1][254] , \round_in[1][253] , \round_in[1][252] , 
        \round_in[1][251] , \round_in[1][250] , \round_in[1][249] , 
        \round_in[1][248] , \round_in[1][247] , \round_in[1][246] , 
        \round_in[1][245] , \round_in[1][244] , \round_in[1][243] , 
        \round_in[1][242] , \round_in[1][241] , \round_in[1][240] , 
        \round_in[1][239] , \round_in[1][238] , \round_in[1][237] , 
        \round_in[1][236] , \round_in[1][235] , \round_in[1][234] , 
        \round_in[1][233] , \round_in[1][232] , \round_in[1][231] , 
        \round_in[1][230] , \round_in[1][229] , \round_in[1][228] , 
        \round_in[1][227] , \round_in[1][226] , \round_in[1][225] , 
        \round_in[1][224] , \round_in[1][223] , \round_in[1][222] , 
        \round_in[1][221] , \round_in[1][220] , \round_in[1][219] , 
        \round_in[1][218] , \round_in[1][217] , \round_in[1][216] , 
        \round_in[1][215] , \round_in[1][214] , \round_in[1][213] , 
        \round_in[1][212] , \round_in[1][211] , \round_in[1][210] , 
        \round_in[1][209] , \round_in[1][208] , \round_in[1][207] , 
        \round_in[1][206] , \round_in[1][205] , \round_in[1][204] , 
        \round_in[1][203] , \round_in[1][202] , \round_in[1][201] , 
        \round_in[1][200] , \round_in[1][199] , \round_in[1][198] , 
        \round_in[1][197] , \round_in[1][196] , \round_in[1][195] , 
        \round_in[1][194] , \round_in[1][193] , \round_in[1][192] , 
        \round_in[1][191] , \round_in[1][190] , \round_in[1][189] , 
        \round_in[1][188] , \round_in[1][187] , \round_in[1][186] , 
        \round_in[1][185] , \round_in[1][184] , \round_in[1][183] , 
        \round_in[1][182] , \round_in[1][181] , \round_in[1][180] , 
        \round_in[1][179] , \round_in[1][178] , \round_in[1][177] , 
        \round_in[1][176] , \round_in[1][175] , \round_in[1][174] , 
        \round_in[1][173] , \round_in[1][172] , \round_in[1][171] , 
        \round_in[1][170] , \round_in[1][169] , \round_in[1][168] , 
        \round_in[1][167] , \round_in[1][166] , \round_in[1][165] , 
        \round_in[1][164] , \round_in[1][163] , \round_in[1][162] , 
        \round_in[1][161] , \round_in[1][160] , \round_in[1][159] , 
        \round_in[1][158] , \round_in[1][157] , \round_in[1][156] , 
        \round_in[1][155] , \round_in[1][154] , \round_in[1][153] , 
        \round_in[1][152] , \round_in[1][151] , \round_in[1][150] , 
        \round_in[1][149] , \round_in[1][148] , \round_in[1][147] , 
        \round_in[1][146] , \round_in[1][145] , \round_in[1][144] , 
        \round_in[1][143] , \round_in[1][142] , \round_in[1][141] , 
        \round_in[1][140] , \round_in[1][139] , \round_in[1][138] , 
        \round_in[1][137] , \round_in[1][136] , \round_in[1][135] , 
        \round_in[1][134] , \round_in[1][133] , \round_in[1][132] , 
        \round_in[1][131] , \round_in[1][130] , \round_in[1][129] , 
        \round_in[1][128] , \round_in[1][127] , \round_in[1][126] , 
        \round_in[1][125] , \round_in[1][124] , \round_in[1][123] , 
        \round_in[1][122] , \round_in[1][121] , \round_in[1][120] , 
        \round_in[1][119] , \round_in[1][118] , \round_in[1][117] , 
        \round_in[1][116] , \round_in[1][115] , \round_in[1][114] , 
        \round_in[1][113] , \round_in[1][112] , \round_in[1][111] , 
        \round_in[1][110] , \round_in[1][109] , \round_in[1][108] , 
        \round_in[1][107] , \round_in[1][106] , \round_in[1][105] , 
        \round_in[1][104] , \round_in[1][103] , \round_in[1][102] , 
        \round_in[1][101] , \round_in[1][100] , \round_in[1][99] , 
        \round_in[1][98] , \round_in[1][97] , \round_in[1][96] , 
        \round_in[1][95] , \round_in[1][94] , \round_in[1][93] , 
        \round_in[1][92] , \round_in[1][91] , \round_in[1][90] , 
        \round_in[1][89] , \round_in[1][88] , \round_in[1][87] , 
        \round_in[1][86] , \round_in[1][85] , \round_in[1][84] , 
        \round_in[1][83] , \round_in[1][82] , \round_in[1][81] , 
        \round_in[1][80] , \round_in[1][79] , \round_in[1][78] , 
        \round_in[1][77] , \round_in[1][76] , \round_in[1][75] , 
        \round_in[1][74] , \round_in[1][73] , \round_in[1][72] , 
        \round_in[1][71] , \round_in[1][70] , \round_in[1][69] , 
        \round_in[1][68] , \round_in[1][67] , \round_in[1][66] , 
        \round_in[1][65] , \round_in[1][64] , \round_in[1][63] , 
        \round_in[1][62] , \round_in[1][61] , \round_in[1][60] , 
        \round_in[1][59] , \round_in[1][58] , \round_in[1][57] , 
        \round_in[1][56] , \round_in[1][55] , \round_in[1][54] , 
        \round_in[1][53] , \round_in[1][52] , \round_in[1][51] , 
        \round_in[1][50] , \round_in[1][49] , \round_in[1][48] , 
        \round_in[1][47] , \round_in[1][46] , \round_in[1][45] , 
        \round_in[1][44] , \round_in[1][43] , \round_in[1][42] , 
        \round_in[1][41] , \round_in[1][40] , \round_in[1][39] , 
        \round_in[1][38] , \round_in[1][37] , \round_in[1][36] , 
        \round_in[1][35] , \round_in[1][34] , \round_in[1][33] , 
        \round_in[1][32] , \round_in[1][31] , \round_in[1][30] , 
        \round_in[1][29] , \round_in[1][28] , \round_in[1][27] , 
        \round_in[1][26] , \round_in[1][25] , \round_in[1][24] , 
        \round_in[1][23] , \round_in[1][22] , \round_in[1][21] , 
        \round_in[1][20] , \round_in[1][19] , \round_in[1][18] , 
        \round_in[1][17] , \round_in[1][16] , \round_in[1][15] , 
        \round_in[1][14] , \round_in[1][13] , \round_in[1][12] , 
        \round_in[1][11] , \round_in[1][10] , \round_in[1][9] , 
        \round_in[1][8] , \round_in[1][7] , \round_in[1][6] , \round_in[1][5] , 
        \round_in[1][4] , \round_in[1][3] , \round_in[1][2] , \round_in[1][1] , 
        \round_in[1][0] }) );
  round_5 \ROUND[1].round_  ( .in({\round_in[1][1599] , \round_in[1][1598] , 
        \round_in[1][1597] , \round_in[1][1596] , \round_in[1][1595] , 
        \round_in[1][1594] , \round_in[1][1593] , \round_in[1][1592] , 
        \round_in[1][1591] , \round_in[1][1590] , \round_in[1][1589] , 
        \round_in[1][1588] , \round_in[1][1587] , \round_in[1][1586] , 
        \round_in[1][1585] , \round_in[1][1584] , \round_in[1][1583] , 
        \round_in[1][1582] , \round_in[1][1581] , \round_in[1][1580] , 
        \round_in[1][1579] , \round_in[1][1578] , \round_in[1][1577] , 
        \round_in[1][1576] , \round_in[1][1575] , \round_in[1][1574] , 
        \round_in[1][1573] , \round_in[1][1572] , \round_in[1][1571] , 
        \round_in[1][1570] , \round_in[1][1569] , \round_in[1][1568] , 
        \round_in[1][1567] , \round_in[1][1566] , \round_in[1][1565] , 
        \round_in[1][1564] , \round_in[1][1563] , \round_in[1][1562] , 
        \round_in[1][1561] , \round_in[1][1560] , \round_in[1][1559] , 
        \round_in[1][1558] , \round_in[1][1557] , \round_in[1][1556] , 
        \round_in[1][1555] , \round_in[1][1554] , \round_in[1][1553] , 
        \round_in[1][1552] , \round_in[1][1551] , \round_in[1][1550] , 
        \round_in[1][1549] , \round_in[1][1548] , \round_in[1][1547] , 
        \round_in[1][1546] , \round_in[1][1545] , \round_in[1][1544] , 
        \round_in[1][1543] , \round_in[1][1542] , \round_in[1][1541] , 
        \round_in[1][1540] , \round_in[1][1539] , \round_in[1][1538] , 
        \round_in[1][1537] , \round_in[1][1536] , \round_in[1][1535] , 
        \round_in[1][1534] , \round_in[1][1533] , \round_in[1][1532] , 
        \round_in[1][1531] , \round_in[1][1530] , \round_in[1][1529] , 
        \round_in[1][1528] , \round_in[1][1527] , \round_in[1][1526] , 
        \round_in[1][1525] , \round_in[1][1524] , \round_in[1][1523] , 
        \round_in[1][1522] , \round_in[1][1521] , \round_in[1][1520] , 
        \round_in[1][1519] , \round_in[1][1518] , \round_in[1][1517] , 
        \round_in[1][1516] , \round_in[1][1515] , \round_in[1][1514] , 
        \round_in[1][1513] , \round_in[1][1512] , \round_in[1][1511] , 
        \round_in[1][1510] , \round_in[1][1509] , \round_in[1][1508] , 
        \round_in[1][1507] , \round_in[1][1506] , \round_in[1][1505] , 
        \round_in[1][1504] , \round_in[1][1503] , \round_in[1][1502] , 
        \round_in[1][1501] , \round_in[1][1500] , \round_in[1][1499] , 
        \round_in[1][1498] , \round_in[1][1497] , \round_in[1][1496] , 
        \round_in[1][1495] , \round_in[1][1494] , \round_in[1][1493] , 
        \round_in[1][1492] , \round_in[1][1491] , \round_in[1][1490] , 
        \round_in[1][1489] , \round_in[1][1488] , \round_in[1][1487] , 
        \round_in[1][1486] , \round_in[1][1485] , \round_in[1][1484] , 
        \round_in[1][1483] , \round_in[1][1482] , \round_in[1][1481] , 
        \round_in[1][1480] , \round_in[1][1479] , \round_in[1][1478] , 
        \round_in[1][1477] , \round_in[1][1476] , \round_in[1][1475] , 
        \round_in[1][1474] , \round_in[1][1473] , \round_in[1][1472] , 
        \round_in[1][1471] , \round_in[1][1470] , \round_in[1][1469] , 
        \round_in[1][1468] , \round_in[1][1467] , \round_in[1][1466] , 
        \round_in[1][1465] , \round_in[1][1464] , \round_in[1][1463] , 
        \round_in[1][1462] , \round_in[1][1461] , \round_in[1][1460] , 
        \round_in[1][1459] , \round_in[1][1458] , \round_in[1][1457] , 
        \round_in[1][1456] , \round_in[1][1455] , \round_in[1][1454] , 
        \round_in[1][1453] , \round_in[1][1452] , \round_in[1][1451] , 
        \round_in[1][1450] , \round_in[1][1449] , \round_in[1][1448] , 
        \round_in[1][1447] , \round_in[1][1446] , \round_in[1][1445] , 
        \round_in[1][1444] , \round_in[1][1443] , \round_in[1][1442] , 
        \round_in[1][1441] , \round_in[1][1440] , \round_in[1][1439] , 
        \round_in[1][1438] , \round_in[1][1437] , \round_in[1][1436] , 
        \round_in[1][1435] , \round_in[1][1434] , \round_in[1][1433] , 
        \round_in[1][1432] , \round_in[1][1431] , \round_in[1][1430] , 
        \round_in[1][1429] , \round_in[1][1428] , \round_in[1][1427] , 
        \round_in[1][1426] , \round_in[1][1425] , \round_in[1][1424] , 
        \round_in[1][1423] , \round_in[1][1422] , \round_in[1][1421] , 
        \round_in[1][1420] , \round_in[1][1419] , \round_in[1][1418] , 
        \round_in[1][1417] , \round_in[1][1416] , \round_in[1][1415] , 
        \round_in[1][1414] , \round_in[1][1413] , \round_in[1][1412] , 
        \round_in[1][1411] , \round_in[1][1410] , \round_in[1][1409] , 
        \round_in[1][1408] , \round_in[1][1407] , \round_in[1][1406] , 
        \round_in[1][1405] , \round_in[1][1404] , \round_in[1][1403] , 
        \round_in[1][1402] , \round_in[1][1401] , \round_in[1][1400] , 
        \round_in[1][1399] , \round_in[1][1398] , \round_in[1][1397] , 
        \round_in[1][1396] , \round_in[1][1395] , \round_in[1][1394] , 
        \round_in[1][1393] , \round_in[1][1392] , \round_in[1][1391] , 
        \round_in[1][1390] , \round_in[1][1389] , \round_in[1][1388] , 
        \round_in[1][1387] , \round_in[1][1386] , \round_in[1][1385] , 
        \round_in[1][1384] , \round_in[1][1383] , \round_in[1][1382] , 
        \round_in[1][1381] , \round_in[1][1380] , \round_in[1][1379] , 
        \round_in[1][1378] , \round_in[1][1377] , \round_in[1][1376] , 
        \round_in[1][1375] , \round_in[1][1374] , \round_in[1][1373] , 
        \round_in[1][1372] , \round_in[1][1371] , \round_in[1][1370] , 
        \round_in[1][1369] , \round_in[1][1368] , \round_in[1][1367] , 
        \round_in[1][1366] , \round_in[1][1365] , \round_in[1][1364] , 
        \round_in[1][1363] , \round_in[1][1362] , \round_in[1][1361] , 
        \round_in[1][1360] , \round_in[1][1359] , \round_in[1][1358] , 
        \round_in[1][1357] , \round_in[1][1356] , \round_in[1][1355] , 
        \round_in[1][1354] , \round_in[1][1353] , \round_in[1][1352] , 
        \round_in[1][1351] , \round_in[1][1350] , \round_in[1][1349] , 
        \round_in[1][1348] , \round_in[1][1347] , \round_in[1][1346] , 
        \round_in[1][1345] , \round_in[1][1344] , \round_in[1][1343] , 
        \round_in[1][1342] , \round_in[1][1341] , \round_in[1][1340] , 
        \round_in[1][1339] , \round_in[1][1338] , \round_in[1][1337] , 
        \round_in[1][1336] , \round_in[1][1335] , \round_in[1][1334] , 
        \round_in[1][1333] , \round_in[1][1332] , \round_in[1][1331] , 
        \round_in[1][1330] , \round_in[1][1329] , \round_in[1][1328] , 
        \round_in[1][1327] , \round_in[1][1326] , \round_in[1][1325] , 
        \round_in[1][1324] , \round_in[1][1323] , \round_in[1][1322] , 
        \round_in[1][1321] , \round_in[1][1320] , \round_in[1][1319] , 
        \round_in[1][1318] , \round_in[1][1317] , \round_in[1][1316] , 
        \round_in[1][1315] , \round_in[1][1314] , \round_in[1][1313] , 
        \round_in[1][1312] , \round_in[1][1311] , \round_in[1][1310] , 
        \round_in[1][1309] , \round_in[1][1308] , \round_in[1][1307] , 
        \round_in[1][1306] , \round_in[1][1305] , \round_in[1][1304] , 
        \round_in[1][1303] , \round_in[1][1302] , \round_in[1][1301] , 
        \round_in[1][1300] , \round_in[1][1299] , \round_in[1][1298] , 
        \round_in[1][1297] , \round_in[1][1296] , \round_in[1][1295] , 
        \round_in[1][1294] , \round_in[1][1293] , \round_in[1][1292] , 
        \round_in[1][1291] , \round_in[1][1290] , \round_in[1][1289] , 
        \round_in[1][1288] , \round_in[1][1287] , \round_in[1][1286] , 
        \round_in[1][1285] , \round_in[1][1284] , \round_in[1][1283] , 
        \round_in[1][1282] , \round_in[1][1281] , \round_in[1][1280] , 
        \round_in[1][1279] , \round_in[1][1278] , \round_in[1][1277] , 
        \round_in[1][1276] , \round_in[1][1275] , \round_in[1][1274] , 
        \round_in[1][1273] , \round_in[1][1272] , \round_in[1][1271] , 
        \round_in[1][1270] , \round_in[1][1269] , \round_in[1][1268] , 
        \round_in[1][1267] , \round_in[1][1266] , \round_in[1][1265] , 
        \round_in[1][1264] , \round_in[1][1263] , \round_in[1][1262] , 
        \round_in[1][1261] , \round_in[1][1260] , \round_in[1][1259] , 
        \round_in[1][1258] , \round_in[1][1257] , \round_in[1][1256] , 
        \round_in[1][1255] , \round_in[1][1254] , \round_in[1][1253] , 
        \round_in[1][1252] , \round_in[1][1251] , \round_in[1][1250] , 
        \round_in[1][1249] , \round_in[1][1248] , \round_in[1][1247] , 
        \round_in[1][1246] , \round_in[1][1245] , \round_in[1][1244] , 
        \round_in[1][1243] , \round_in[1][1242] , \round_in[1][1241] , 
        \round_in[1][1240] , \round_in[1][1239] , \round_in[1][1238] , 
        \round_in[1][1237] , \round_in[1][1236] , \round_in[1][1235] , 
        \round_in[1][1234] , \round_in[1][1233] , \round_in[1][1232] , 
        \round_in[1][1231] , \round_in[1][1230] , \round_in[1][1229] , 
        \round_in[1][1228] , \round_in[1][1227] , \round_in[1][1226] , 
        \round_in[1][1225] , \round_in[1][1224] , \round_in[1][1223] , 
        \round_in[1][1222] , \round_in[1][1221] , \round_in[1][1220] , 
        \round_in[1][1219] , \round_in[1][1218] , \round_in[1][1217] , 
        \round_in[1][1216] , \round_in[1][1215] , \round_in[1][1214] , 
        \round_in[1][1213] , \round_in[1][1212] , \round_in[1][1211] , 
        \round_in[1][1210] , \round_in[1][1209] , \round_in[1][1208] , 
        \round_in[1][1207] , \round_in[1][1206] , \round_in[1][1205] , 
        \round_in[1][1204] , \round_in[1][1203] , \round_in[1][1202] , 
        \round_in[1][1201] , \round_in[1][1200] , \round_in[1][1199] , 
        \round_in[1][1198] , \round_in[1][1197] , \round_in[1][1196] , 
        \round_in[1][1195] , \round_in[1][1194] , \round_in[1][1193] , 
        \round_in[1][1192] , \round_in[1][1191] , \round_in[1][1190] , 
        \round_in[1][1189] , \round_in[1][1188] , \round_in[1][1187] , 
        \round_in[1][1186] , \round_in[1][1185] , \round_in[1][1184] , 
        \round_in[1][1183] , \round_in[1][1182] , \round_in[1][1181] , 
        \round_in[1][1180] , \round_in[1][1179] , \round_in[1][1178] , 
        \round_in[1][1177] , \round_in[1][1176] , \round_in[1][1175] , 
        \round_in[1][1174] , \round_in[1][1173] , \round_in[1][1172] , 
        \round_in[1][1171] , \round_in[1][1170] , \round_in[1][1169] , 
        \round_in[1][1168] , \round_in[1][1167] , \round_in[1][1166] , 
        \round_in[1][1165] , \round_in[1][1164] , \round_in[1][1163] , 
        \round_in[1][1162] , \round_in[1][1161] , \round_in[1][1160] , 
        \round_in[1][1159] , \round_in[1][1158] , \round_in[1][1157] , 
        \round_in[1][1156] , \round_in[1][1155] , \round_in[1][1154] , 
        \round_in[1][1153] , \round_in[1][1152] , \round_in[1][1151] , 
        \round_in[1][1150] , \round_in[1][1149] , \round_in[1][1148] , 
        \round_in[1][1147] , \round_in[1][1146] , \round_in[1][1145] , 
        \round_in[1][1144] , \round_in[1][1143] , \round_in[1][1142] , 
        \round_in[1][1141] , \round_in[1][1140] , \round_in[1][1139] , 
        \round_in[1][1138] , \round_in[1][1137] , \round_in[1][1136] , 
        \round_in[1][1135] , \round_in[1][1134] , \round_in[1][1133] , 
        \round_in[1][1132] , \round_in[1][1131] , \round_in[1][1130] , 
        \round_in[1][1129] , \round_in[1][1128] , \round_in[1][1127] , 
        \round_in[1][1126] , \round_in[1][1125] , \round_in[1][1124] , 
        \round_in[1][1123] , \round_in[1][1122] , \round_in[1][1121] , 
        \round_in[1][1120] , \round_in[1][1119] , \round_in[1][1118] , 
        \round_in[1][1117] , \round_in[1][1116] , \round_in[1][1115] , 
        \round_in[1][1114] , \round_in[1][1113] , \round_in[1][1112] , 
        \round_in[1][1111] , \round_in[1][1110] , \round_in[1][1109] , 
        \round_in[1][1108] , \round_in[1][1107] , \round_in[1][1106] , 
        \round_in[1][1105] , \round_in[1][1104] , \round_in[1][1103] , 
        \round_in[1][1102] , \round_in[1][1101] , \round_in[1][1100] , 
        \round_in[1][1099] , \round_in[1][1098] , \round_in[1][1097] , 
        \round_in[1][1096] , \round_in[1][1095] , \round_in[1][1094] , 
        \round_in[1][1093] , \round_in[1][1092] , \round_in[1][1091] , 
        \round_in[1][1090] , \round_in[1][1089] , \round_in[1][1088] , 
        \round_in[1][1087] , \round_in[1][1086] , \round_in[1][1085] , 
        \round_in[1][1084] , \round_in[1][1083] , \round_in[1][1082] , 
        \round_in[1][1081] , \round_in[1][1080] , \round_in[1][1079] , 
        \round_in[1][1078] , \round_in[1][1077] , \round_in[1][1076] , 
        \round_in[1][1075] , \round_in[1][1074] , \round_in[1][1073] , 
        \round_in[1][1072] , \round_in[1][1071] , \round_in[1][1070] , 
        \round_in[1][1069] , \round_in[1][1068] , \round_in[1][1067] , 
        \round_in[1][1066] , \round_in[1][1065] , \round_in[1][1064] , 
        \round_in[1][1063] , \round_in[1][1062] , \round_in[1][1061] , 
        \round_in[1][1060] , \round_in[1][1059] , \round_in[1][1058] , 
        \round_in[1][1057] , \round_in[1][1056] , \round_in[1][1055] , 
        \round_in[1][1054] , \round_in[1][1053] , \round_in[1][1052] , 
        \round_in[1][1051] , \round_in[1][1050] , \round_in[1][1049] , 
        \round_in[1][1048] , \round_in[1][1047] , \round_in[1][1046] , 
        \round_in[1][1045] , \round_in[1][1044] , \round_in[1][1043] , 
        \round_in[1][1042] , \round_in[1][1041] , \round_in[1][1040] , 
        \round_in[1][1039] , \round_in[1][1038] , \round_in[1][1037] , 
        \round_in[1][1036] , \round_in[1][1035] , \round_in[1][1034] , 
        \round_in[1][1033] , \round_in[1][1032] , \round_in[1][1031] , 
        \round_in[1][1030] , \round_in[1][1029] , \round_in[1][1028] , 
        \round_in[1][1027] , \round_in[1][1026] , \round_in[1][1025] , 
        \round_in[1][1024] , \round_in[1][1023] , \round_in[1][1022] , 
        \round_in[1][1021] , \round_in[1][1020] , \round_in[1][1019] , 
        \round_in[1][1018] , \round_in[1][1017] , \round_in[1][1016] , 
        \round_in[1][1015] , \round_in[1][1014] , \round_in[1][1013] , 
        \round_in[1][1012] , \round_in[1][1011] , \round_in[1][1010] , 
        \round_in[1][1009] , \round_in[1][1008] , \round_in[1][1007] , 
        \round_in[1][1006] , \round_in[1][1005] , \round_in[1][1004] , 
        \round_in[1][1003] , \round_in[1][1002] , \round_in[1][1001] , 
        \round_in[1][1000] , \round_in[1][999] , \round_in[1][998] , 
        \round_in[1][997] , \round_in[1][996] , \round_in[1][995] , 
        \round_in[1][994] , \round_in[1][993] , \round_in[1][992] , 
        \round_in[1][991] , \round_in[1][990] , \round_in[1][989] , 
        \round_in[1][988] , \round_in[1][987] , \round_in[1][986] , 
        \round_in[1][985] , \round_in[1][984] , \round_in[1][983] , 
        \round_in[1][982] , \round_in[1][981] , \round_in[1][980] , 
        \round_in[1][979] , \round_in[1][978] , \round_in[1][977] , 
        \round_in[1][976] , \round_in[1][975] , \round_in[1][974] , 
        \round_in[1][973] , \round_in[1][972] , \round_in[1][971] , 
        \round_in[1][970] , \round_in[1][969] , \round_in[1][968] , 
        \round_in[1][967] , \round_in[1][966] , \round_in[1][965] , 
        \round_in[1][964] , \round_in[1][963] , \round_in[1][962] , 
        \round_in[1][961] , \round_in[1][960] , \round_in[1][959] , 
        \round_in[1][958] , \round_in[1][957] , \round_in[1][956] , 
        \round_in[1][955] , \round_in[1][954] , \round_in[1][953] , 
        \round_in[1][952] , \round_in[1][951] , \round_in[1][950] , 
        \round_in[1][949] , \round_in[1][948] , \round_in[1][947] , 
        \round_in[1][946] , \round_in[1][945] , \round_in[1][944] , 
        \round_in[1][943] , \round_in[1][942] , \round_in[1][941] , 
        \round_in[1][940] , \round_in[1][939] , \round_in[1][938] , 
        \round_in[1][937] , \round_in[1][936] , \round_in[1][935] , 
        \round_in[1][934] , \round_in[1][933] , \round_in[1][932] , 
        \round_in[1][931] , \round_in[1][930] , \round_in[1][929] , 
        \round_in[1][928] , \round_in[1][927] , \round_in[1][926] , 
        \round_in[1][925] , \round_in[1][924] , \round_in[1][923] , 
        \round_in[1][922] , \round_in[1][921] , \round_in[1][920] , 
        \round_in[1][919] , \round_in[1][918] , \round_in[1][917] , 
        \round_in[1][916] , \round_in[1][915] , \round_in[1][914] , 
        \round_in[1][913] , \round_in[1][912] , \round_in[1][911] , 
        \round_in[1][910] , \round_in[1][909] , \round_in[1][908] , 
        \round_in[1][907] , \round_in[1][906] , \round_in[1][905] , 
        \round_in[1][904] , \round_in[1][903] , \round_in[1][902] , 
        \round_in[1][901] , \round_in[1][900] , \round_in[1][899] , 
        \round_in[1][898] , \round_in[1][897] , \round_in[1][896] , 
        \round_in[1][895] , \round_in[1][894] , \round_in[1][893] , 
        \round_in[1][892] , \round_in[1][891] , \round_in[1][890] , 
        \round_in[1][889] , \round_in[1][888] , \round_in[1][887] , 
        \round_in[1][886] , \round_in[1][885] , \round_in[1][884] , 
        \round_in[1][883] , \round_in[1][882] , \round_in[1][881] , 
        \round_in[1][880] , \round_in[1][879] , \round_in[1][878] , 
        \round_in[1][877] , \round_in[1][876] , \round_in[1][875] , 
        \round_in[1][874] , \round_in[1][873] , \round_in[1][872] , 
        \round_in[1][871] , \round_in[1][870] , \round_in[1][869] , 
        \round_in[1][868] , \round_in[1][867] , \round_in[1][866] , 
        \round_in[1][865] , \round_in[1][864] , \round_in[1][863] , 
        \round_in[1][862] , \round_in[1][861] , \round_in[1][860] , 
        \round_in[1][859] , \round_in[1][858] , \round_in[1][857] , 
        \round_in[1][856] , \round_in[1][855] , \round_in[1][854] , 
        \round_in[1][853] , \round_in[1][852] , \round_in[1][851] , 
        \round_in[1][850] , \round_in[1][849] , \round_in[1][848] , 
        \round_in[1][847] , \round_in[1][846] , \round_in[1][845] , 
        \round_in[1][844] , \round_in[1][843] , \round_in[1][842] , 
        \round_in[1][841] , \round_in[1][840] , \round_in[1][839] , 
        \round_in[1][838] , \round_in[1][837] , \round_in[1][836] , 
        \round_in[1][835] , \round_in[1][834] , \round_in[1][833] , 
        \round_in[1][832] , \round_in[1][831] , \round_in[1][830] , 
        \round_in[1][829] , \round_in[1][828] , \round_in[1][827] , 
        \round_in[1][826] , \round_in[1][825] , \round_in[1][824] , 
        \round_in[1][823] , \round_in[1][822] , \round_in[1][821] , 
        \round_in[1][820] , \round_in[1][819] , \round_in[1][818] , 
        \round_in[1][817] , \round_in[1][816] , \round_in[1][815] , 
        \round_in[1][814] , \round_in[1][813] , \round_in[1][812] , 
        \round_in[1][811] , \round_in[1][810] , \round_in[1][809] , 
        \round_in[1][808] , \round_in[1][807] , \round_in[1][806] , 
        \round_in[1][805] , \round_in[1][804] , \round_in[1][803] , 
        \round_in[1][802] , \round_in[1][801] , \round_in[1][800] , 
        \round_in[1][799] , \round_in[1][798] , \round_in[1][797] , 
        \round_in[1][796] , \round_in[1][795] , \round_in[1][794] , 
        \round_in[1][793] , \round_in[1][792] , \round_in[1][791] , 
        \round_in[1][790] , \round_in[1][789] , \round_in[1][788] , 
        \round_in[1][787] , \round_in[1][786] , \round_in[1][785] , 
        \round_in[1][784] , \round_in[1][783] , \round_in[1][782] , 
        \round_in[1][781] , \round_in[1][780] , \round_in[1][779] , 
        \round_in[1][778] , \round_in[1][777] , \round_in[1][776] , 
        \round_in[1][775] , \round_in[1][774] , \round_in[1][773] , 
        \round_in[1][772] , \round_in[1][771] , \round_in[1][770] , 
        \round_in[1][769] , \round_in[1][768] , \round_in[1][767] , 
        \round_in[1][766] , \round_in[1][765] , \round_in[1][764] , 
        \round_in[1][763] , \round_in[1][762] , \round_in[1][761] , 
        \round_in[1][760] , \round_in[1][759] , \round_in[1][758] , 
        \round_in[1][757] , \round_in[1][756] , \round_in[1][755] , 
        \round_in[1][754] , \round_in[1][753] , \round_in[1][752] , 
        \round_in[1][751] , \round_in[1][750] , \round_in[1][749] , 
        \round_in[1][748] , \round_in[1][747] , \round_in[1][746] , 
        \round_in[1][745] , \round_in[1][744] , \round_in[1][743] , 
        \round_in[1][742] , \round_in[1][741] , \round_in[1][740] , 
        \round_in[1][739] , \round_in[1][738] , \round_in[1][737] , 
        \round_in[1][736] , \round_in[1][735] , \round_in[1][734] , 
        \round_in[1][733] , \round_in[1][732] , \round_in[1][731] , 
        \round_in[1][730] , \round_in[1][729] , \round_in[1][728] , 
        \round_in[1][727] , \round_in[1][726] , \round_in[1][725] , 
        \round_in[1][724] , \round_in[1][723] , \round_in[1][722] , 
        \round_in[1][721] , \round_in[1][720] , \round_in[1][719] , 
        \round_in[1][718] , \round_in[1][717] , \round_in[1][716] , 
        \round_in[1][715] , \round_in[1][714] , \round_in[1][713] , 
        \round_in[1][712] , \round_in[1][711] , \round_in[1][710] , 
        \round_in[1][709] , \round_in[1][708] , \round_in[1][707] , 
        \round_in[1][706] , \round_in[1][705] , \round_in[1][704] , 
        \round_in[1][703] , \round_in[1][702] , \round_in[1][701] , 
        \round_in[1][700] , \round_in[1][699] , \round_in[1][698] , 
        \round_in[1][697] , \round_in[1][696] , \round_in[1][695] , 
        \round_in[1][694] , \round_in[1][693] , \round_in[1][692] , 
        \round_in[1][691] , \round_in[1][690] , \round_in[1][689] , 
        \round_in[1][688] , \round_in[1][687] , \round_in[1][686] , 
        \round_in[1][685] , \round_in[1][684] , \round_in[1][683] , 
        \round_in[1][682] , \round_in[1][681] , \round_in[1][680] , 
        \round_in[1][679] , \round_in[1][678] , \round_in[1][677] , 
        \round_in[1][676] , \round_in[1][675] , \round_in[1][674] , 
        \round_in[1][673] , \round_in[1][672] , \round_in[1][671] , 
        \round_in[1][670] , \round_in[1][669] , \round_in[1][668] , 
        \round_in[1][667] , \round_in[1][666] , \round_in[1][665] , 
        \round_in[1][664] , \round_in[1][663] , \round_in[1][662] , 
        \round_in[1][661] , \round_in[1][660] , \round_in[1][659] , 
        \round_in[1][658] , \round_in[1][657] , \round_in[1][656] , 
        \round_in[1][655] , \round_in[1][654] , \round_in[1][653] , 
        \round_in[1][652] , \round_in[1][651] , \round_in[1][650] , 
        \round_in[1][649] , \round_in[1][648] , \round_in[1][647] , 
        \round_in[1][646] , \round_in[1][645] , \round_in[1][644] , 
        \round_in[1][643] , \round_in[1][642] , \round_in[1][641] , 
        \round_in[1][640] , \round_in[1][639] , \round_in[1][638] , 
        \round_in[1][637] , \round_in[1][636] , \round_in[1][635] , 
        \round_in[1][634] , \round_in[1][633] , \round_in[1][632] , 
        \round_in[1][631] , \round_in[1][630] , \round_in[1][629] , 
        \round_in[1][628] , \round_in[1][627] , \round_in[1][626] , 
        \round_in[1][625] , \round_in[1][624] , \round_in[1][623] , 
        \round_in[1][622] , \round_in[1][621] , \round_in[1][620] , 
        \round_in[1][619] , \round_in[1][618] , \round_in[1][617] , 
        \round_in[1][616] , \round_in[1][615] , \round_in[1][614] , 
        \round_in[1][613] , \round_in[1][612] , \round_in[1][611] , 
        \round_in[1][610] , \round_in[1][609] , \round_in[1][608] , 
        \round_in[1][607] , \round_in[1][606] , \round_in[1][605] , 
        \round_in[1][604] , \round_in[1][603] , \round_in[1][602] , 
        \round_in[1][601] , \round_in[1][600] , \round_in[1][599] , 
        \round_in[1][598] , \round_in[1][597] , \round_in[1][596] , 
        \round_in[1][595] , \round_in[1][594] , \round_in[1][593] , 
        \round_in[1][592] , \round_in[1][591] , \round_in[1][590] , 
        \round_in[1][589] , \round_in[1][588] , \round_in[1][587] , 
        \round_in[1][586] , \round_in[1][585] , \round_in[1][584] , 
        \round_in[1][583] , \round_in[1][582] , \round_in[1][581] , 
        \round_in[1][580] , \round_in[1][579] , \round_in[1][578] , 
        \round_in[1][577] , \round_in[1][576] , \round_in[1][575] , 
        \round_in[1][574] , \round_in[1][573] , \round_in[1][572] , 
        \round_in[1][571] , \round_in[1][570] , \round_in[1][569] , 
        \round_in[1][568] , \round_in[1][567] , \round_in[1][566] , 
        \round_in[1][565] , \round_in[1][564] , \round_in[1][563] , 
        \round_in[1][562] , \round_in[1][561] , \round_in[1][560] , 
        \round_in[1][559] , \round_in[1][558] , \round_in[1][557] , 
        \round_in[1][556] , \round_in[1][555] , \round_in[1][554] , 
        \round_in[1][553] , \round_in[1][552] , \round_in[1][551] , 
        \round_in[1][550] , \round_in[1][549] , \round_in[1][548] , 
        \round_in[1][547] , \round_in[1][546] , \round_in[1][545] , 
        \round_in[1][544] , \round_in[1][543] , \round_in[1][542] , 
        \round_in[1][541] , \round_in[1][540] , \round_in[1][539] , 
        \round_in[1][538] , \round_in[1][537] , \round_in[1][536] , 
        \round_in[1][535] , \round_in[1][534] , \round_in[1][533] , 
        \round_in[1][532] , \round_in[1][531] , \round_in[1][530] , 
        \round_in[1][529] , \round_in[1][528] , \round_in[1][527] , 
        \round_in[1][526] , \round_in[1][525] , \round_in[1][524] , 
        \round_in[1][523] , \round_in[1][522] , \round_in[1][521] , 
        \round_in[1][520] , \round_in[1][519] , \round_in[1][518] , 
        \round_in[1][517] , \round_in[1][516] , \round_in[1][515] , 
        \round_in[1][514] , \round_in[1][513] , \round_in[1][512] , 
        \round_in[1][511] , \round_in[1][510] , \round_in[1][509] , 
        \round_in[1][508] , \round_in[1][507] , \round_in[1][506] , 
        \round_in[1][505] , \round_in[1][504] , \round_in[1][503] , 
        \round_in[1][502] , \round_in[1][501] , \round_in[1][500] , 
        \round_in[1][499] , \round_in[1][498] , \round_in[1][497] , 
        \round_in[1][496] , \round_in[1][495] , \round_in[1][494] , 
        \round_in[1][493] , \round_in[1][492] , \round_in[1][491] , 
        \round_in[1][490] , \round_in[1][489] , \round_in[1][488] , 
        \round_in[1][487] , \round_in[1][486] , \round_in[1][485] , 
        \round_in[1][484] , \round_in[1][483] , \round_in[1][482] , 
        \round_in[1][481] , \round_in[1][480] , \round_in[1][479] , 
        \round_in[1][478] , \round_in[1][477] , \round_in[1][476] , 
        \round_in[1][475] , \round_in[1][474] , \round_in[1][473] , 
        \round_in[1][472] , \round_in[1][471] , \round_in[1][470] , 
        \round_in[1][469] , \round_in[1][468] , \round_in[1][467] , 
        \round_in[1][466] , \round_in[1][465] , \round_in[1][464] , 
        \round_in[1][463] , \round_in[1][462] , \round_in[1][461] , 
        \round_in[1][460] , \round_in[1][459] , \round_in[1][458] , 
        \round_in[1][457] , \round_in[1][456] , \round_in[1][455] , 
        \round_in[1][454] , \round_in[1][453] , \round_in[1][452] , 
        \round_in[1][451] , \round_in[1][450] , \round_in[1][449] , 
        \round_in[1][448] , \round_in[1][447] , \round_in[1][446] , 
        \round_in[1][445] , \round_in[1][444] , \round_in[1][443] , 
        \round_in[1][442] , \round_in[1][441] , \round_in[1][440] , 
        \round_in[1][439] , \round_in[1][438] , \round_in[1][437] , 
        \round_in[1][436] , \round_in[1][435] , \round_in[1][434] , 
        \round_in[1][433] , \round_in[1][432] , \round_in[1][431] , 
        \round_in[1][430] , \round_in[1][429] , \round_in[1][428] , 
        \round_in[1][427] , \round_in[1][426] , \round_in[1][425] , 
        \round_in[1][424] , \round_in[1][423] , \round_in[1][422] , 
        \round_in[1][421] , \round_in[1][420] , \round_in[1][419] , 
        \round_in[1][418] , \round_in[1][417] , \round_in[1][416] , 
        \round_in[1][415] , \round_in[1][414] , \round_in[1][413] , 
        \round_in[1][412] , \round_in[1][411] , \round_in[1][410] , 
        \round_in[1][409] , \round_in[1][408] , \round_in[1][407] , 
        \round_in[1][406] , \round_in[1][405] , \round_in[1][404] , 
        \round_in[1][403] , \round_in[1][402] , \round_in[1][401] , 
        \round_in[1][400] , \round_in[1][399] , \round_in[1][398] , 
        \round_in[1][397] , \round_in[1][396] , \round_in[1][395] , 
        \round_in[1][394] , \round_in[1][393] , \round_in[1][392] , 
        \round_in[1][391] , \round_in[1][390] , \round_in[1][389] , 
        \round_in[1][388] , \round_in[1][387] , \round_in[1][386] , 
        \round_in[1][385] , \round_in[1][384] , \round_in[1][383] , 
        \round_in[1][382] , \round_in[1][381] , \round_in[1][380] , 
        \round_in[1][379] , \round_in[1][378] , \round_in[1][377] , 
        \round_in[1][376] , \round_in[1][375] , \round_in[1][374] , 
        \round_in[1][373] , \round_in[1][372] , \round_in[1][371] , 
        \round_in[1][370] , \round_in[1][369] , \round_in[1][368] , 
        \round_in[1][367] , \round_in[1][366] , \round_in[1][365] , 
        \round_in[1][364] , \round_in[1][363] , \round_in[1][362] , 
        \round_in[1][361] , \round_in[1][360] , \round_in[1][359] , 
        \round_in[1][358] , \round_in[1][357] , \round_in[1][356] , 
        \round_in[1][355] , \round_in[1][354] , \round_in[1][353] , 
        \round_in[1][352] , \round_in[1][351] , \round_in[1][350] , 
        \round_in[1][349] , \round_in[1][348] , \round_in[1][347] , 
        \round_in[1][346] , \round_in[1][345] , \round_in[1][344] , 
        \round_in[1][343] , \round_in[1][342] , \round_in[1][341] , 
        \round_in[1][340] , \round_in[1][339] , \round_in[1][338] , 
        \round_in[1][337] , \round_in[1][336] , \round_in[1][335] , 
        \round_in[1][334] , \round_in[1][333] , \round_in[1][332] , 
        \round_in[1][331] , \round_in[1][330] , \round_in[1][329] , 
        \round_in[1][328] , \round_in[1][327] , \round_in[1][326] , 
        \round_in[1][325] , \round_in[1][324] , \round_in[1][323] , 
        \round_in[1][322] , \round_in[1][321] , \round_in[1][320] , 
        \round_in[1][319] , \round_in[1][318] , \round_in[1][317] , 
        \round_in[1][316] , \round_in[1][315] , \round_in[1][314] , 
        \round_in[1][313] , \round_in[1][312] , \round_in[1][311] , 
        \round_in[1][310] , \round_in[1][309] , \round_in[1][308] , 
        \round_in[1][307] , \round_in[1][306] , \round_in[1][305] , 
        \round_in[1][304] , \round_in[1][303] , \round_in[1][302] , 
        \round_in[1][301] , \round_in[1][300] , \round_in[1][299] , 
        \round_in[1][298] , \round_in[1][297] , \round_in[1][296] , 
        \round_in[1][295] , \round_in[1][294] , \round_in[1][293] , 
        \round_in[1][292] , \round_in[1][291] , \round_in[1][290] , 
        \round_in[1][289] , \round_in[1][288] , \round_in[1][287] , 
        \round_in[1][286] , \round_in[1][285] , \round_in[1][284] , 
        \round_in[1][283] , \round_in[1][282] , \round_in[1][281] , 
        \round_in[1][280] , \round_in[1][279] , \round_in[1][278] , 
        \round_in[1][277] , \round_in[1][276] , \round_in[1][275] , 
        \round_in[1][274] , \round_in[1][273] , \round_in[1][272] , 
        \round_in[1][271] , \round_in[1][270] , \round_in[1][269] , 
        \round_in[1][268] , \round_in[1][267] , \round_in[1][266] , 
        \round_in[1][265] , \round_in[1][264] , \round_in[1][263] , 
        \round_in[1][262] , \round_in[1][261] , \round_in[1][260] , 
        \round_in[1][259] , \round_in[1][258] , \round_in[1][257] , 
        \round_in[1][256] , \round_in[1][255] , \round_in[1][254] , 
        \round_in[1][253] , \round_in[1][252] , \round_in[1][251] , 
        \round_in[1][250] , \round_in[1][249] , \round_in[1][248] , 
        \round_in[1][247] , \round_in[1][246] , \round_in[1][245] , 
        \round_in[1][244] , \round_in[1][243] , \round_in[1][242] , 
        \round_in[1][241] , \round_in[1][240] , \round_in[1][239] , 
        \round_in[1][238] , \round_in[1][237] , \round_in[1][236] , 
        \round_in[1][235] , \round_in[1][234] , \round_in[1][233] , 
        \round_in[1][232] , \round_in[1][231] , \round_in[1][230] , 
        \round_in[1][229] , \round_in[1][228] , \round_in[1][227] , 
        \round_in[1][226] , \round_in[1][225] , \round_in[1][224] , 
        \round_in[1][223] , \round_in[1][222] , \round_in[1][221] , 
        \round_in[1][220] , \round_in[1][219] , \round_in[1][218] , 
        \round_in[1][217] , \round_in[1][216] , \round_in[1][215] , 
        \round_in[1][214] , \round_in[1][213] , \round_in[1][212] , 
        \round_in[1][211] , \round_in[1][210] , \round_in[1][209] , 
        \round_in[1][208] , \round_in[1][207] , \round_in[1][206] , 
        \round_in[1][205] , \round_in[1][204] , \round_in[1][203] , 
        \round_in[1][202] , \round_in[1][201] , \round_in[1][200] , 
        \round_in[1][199] , \round_in[1][198] , \round_in[1][197] , 
        \round_in[1][196] , \round_in[1][195] , \round_in[1][194] , 
        \round_in[1][193] , \round_in[1][192] , \round_in[1][191] , 
        \round_in[1][190] , \round_in[1][189] , \round_in[1][188] , 
        \round_in[1][187] , \round_in[1][186] , \round_in[1][185] , 
        \round_in[1][184] , \round_in[1][183] , \round_in[1][182] , 
        \round_in[1][181] , \round_in[1][180] , \round_in[1][179] , 
        \round_in[1][178] , \round_in[1][177] , \round_in[1][176] , 
        \round_in[1][175] , \round_in[1][174] , \round_in[1][173] , 
        \round_in[1][172] , \round_in[1][171] , \round_in[1][170] , 
        \round_in[1][169] , \round_in[1][168] , \round_in[1][167] , 
        \round_in[1][166] , \round_in[1][165] , \round_in[1][164] , 
        \round_in[1][163] , \round_in[1][162] , \round_in[1][161] , 
        \round_in[1][160] , \round_in[1][159] , \round_in[1][158] , 
        \round_in[1][157] , \round_in[1][156] , \round_in[1][155] , 
        \round_in[1][154] , \round_in[1][153] , \round_in[1][152] , 
        \round_in[1][151] , \round_in[1][150] , \round_in[1][149] , 
        \round_in[1][148] , \round_in[1][147] , \round_in[1][146] , 
        \round_in[1][145] , \round_in[1][144] , \round_in[1][143] , 
        \round_in[1][142] , \round_in[1][141] , \round_in[1][140] , 
        \round_in[1][139] , \round_in[1][138] , \round_in[1][137] , 
        \round_in[1][136] , \round_in[1][135] , \round_in[1][134] , 
        \round_in[1][133] , \round_in[1][132] , \round_in[1][131] , 
        \round_in[1][130] , \round_in[1][129] , \round_in[1][128] , 
        \round_in[1][127] , \round_in[1][126] , \round_in[1][125] , 
        \round_in[1][124] , \round_in[1][123] , \round_in[1][122] , 
        \round_in[1][121] , \round_in[1][120] , \round_in[1][119] , 
        \round_in[1][118] , \round_in[1][117] , \round_in[1][116] , 
        \round_in[1][115] , \round_in[1][114] , \round_in[1][113] , 
        \round_in[1][112] , \round_in[1][111] , \round_in[1][110] , 
        \round_in[1][109] , \round_in[1][108] , \round_in[1][107] , 
        \round_in[1][106] , \round_in[1][105] , \round_in[1][104] , 
        \round_in[1][103] , \round_in[1][102] , \round_in[1][101] , 
        \round_in[1][100] , \round_in[1][99] , \round_in[1][98] , 
        \round_in[1][97] , \round_in[1][96] , \round_in[1][95] , 
        \round_in[1][94] , \round_in[1][93] , \round_in[1][92] , 
        \round_in[1][91] , \round_in[1][90] , \round_in[1][89] , 
        \round_in[1][88] , \round_in[1][87] , \round_in[1][86] , 
        \round_in[1][85] , \round_in[1][84] , \round_in[1][83] , 
        \round_in[1][82] , \round_in[1][81] , \round_in[1][80] , 
        \round_in[1][79] , \round_in[1][78] , \round_in[1][77] , 
        \round_in[1][76] , \round_in[1][75] , \round_in[1][74] , 
        \round_in[1][73] , \round_in[1][72] , \round_in[1][71] , 
        \round_in[1][70] , \round_in[1][69] , \round_in[1][68] , 
        \round_in[1][67] , \round_in[1][66] , \round_in[1][65] , 
        \round_in[1][64] , \round_in[1][63] , \round_in[1][62] , 
        \round_in[1][61] , \round_in[1][60] , \round_in[1][59] , 
        \round_in[1][58] , \round_in[1][57] , \round_in[1][56] , 
        \round_in[1][55] , \round_in[1][54] , \round_in[1][53] , 
        \round_in[1][52] , \round_in[1][51] , \round_in[1][50] , 
        \round_in[1][49] , \round_in[1][48] , \round_in[1][47] , 
        \round_in[1][46] , \round_in[1][45] , \round_in[1][44] , 
        \round_in[1][43] , \round_in[1][42] , \round_in[1][41] , 
        \round_in[1][40] , \round_in[1][39] , \round_in[1][38] , 
        \round_in[1][37] , \round_in[1][36] , \round_in[1][35] , 
        \round_in[1][34] , \round_in[1][33] , \round_in[1][32] , 
        \round_in[1][31] , \round_in[1][30] , \round_in[1][29] , 
        \round_in[1][28] , \round_in[1][27] , \round_in[1][26] , 
        \round_in[1][25] , \round_in[1][24] , \round_in[1][23] , 
        \round_in[1][22] , \round_in[1][21] , \round_in[1][20] , 
        \round_in[1][19] , \round_in[1][18] , \round_in[1][17] , 
        \round_in[1][16] , \round_in[1][15] , \round_in[1][14] , 
        \round_in[1][13] , \round_in[1][12] , \round_in[1][11] , 
        \round_in[1][10] , \round_in[1][9] , \round_in[1][8] , 
        \round_in[1][7] , \round_in[1][6] , \round_in[1][5] , \round_in[1][4] , 
        \round_in[1][3] , \round_in[1][2] , \round_in[1][1] , \round_in[1][0] }), .round_const({\RCONST[1].rconst_/N68 , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, rc_i[1], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \RCONST[1].rconst_/N49 , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \rc[1][7] , 1'b0, 1'b0, 1'b0, 
        \RCONST[1].rconst_/N26 , 1'b0, \RCONST[1].rconst_/N15 , 
        \RCONST[3].rconst_/N10 }), .out({\round_in[2][1599] , 
        \round_in[2][1598] , \round_in[2][1597] , \round_in[2][1596] , 
        \round_in[2][1595] , \round_in[2][1594] , \round_in[2][1593] , 
        \round_in[2][1592] , \round_in[2][1591] , \round_in[2][1590] , 
        \round_in[2][1589] , \round_in[2][1588] , \round_in[2][1587] , 
        \round_in[2][1586] , \round_in[2][1585] , \round_in[2][1584] , 
        \round_in[2][1583] , \round_in[2][1582] , \round_in[2][1581] , 
        \round_in[2][1580] , \round_in[2][1579] , \round_in[2][1578] , 
        \round_in[2][1577] , \round_in[2][1576] , \round_in[2][1575] , 
        \round_in[2][1574] , \round_in[2][1573] , \round_in[2][1572] , 
        \round_in[2][1571] , \round_in[2][1570] , \round_in[2][1569] , 
        \round_in[2][1568] , \round_in[2][1567] , \round_in[2][1566] , 
        \round_in[2][1565] , \round_in[2][1564] , \round_in[2][1563] , 
        \round_in[2][1562] , \round_in[2][1561] , \round_in[2][1560] , 
        \round_in[2][1559] , \round_in[2][1558] , \round_in[2][1557] , 
        \round_in[2][1556] , \round_in[2][1555] , \round_in[2][1554] , 
        \round_in[2][1553] , \round_in[2][1552] , \round_in[2][1551] , 
        \round_in[2][1550] , \round_in[2][1549] , \round_in[2][1548] , 
        \round_in[2][1547] , \round_in[2][1546] , \round_in[2][1545] , 
        \round_in[2][1544] , \round_in[2][1543] , \round_in[2][1542] , 
        \round_in[2][1541] , \round_in[2][1540] , \round_in[2][1539] , 
        \round_in[2][1538] , \round_in[2][1537] , \round_in[2][1536] , 
        \round_in[2][1535] , \round_in[2][1534] , \round_in[2][1533] , 
        \round_in[2][1532] , \round_in[2][1531] , \round_in[2][1530] , 
        \round_in[2][1529] , \round_in[2][1528] , \round_in[2][1527] , 
        \round_in[2][1526] , \round_in[2][1525] , \round_in[2][1524] , 
        \round_in[2][1523] , \round_in[2][1522] , \round_in[2][1521] , 
        \round_in[2][1520] , \round_in[2][1519] , \round_in[2][1518] , 
        \round_in[2][1517] , \round_in[2][1516] , \round_in[2][1515] , 
        \round_in[2][1514] , \round_in[2][1513] , \round_in[2][1512] , 
        \round_in[2][1511] , \round_in[2][1510] , \round_in[2][1509] , 
        \round_in[2][1508] , \round_in[2][1507] , \round_in[2][1506] , 
        \round_in[2][1505] , \round_in[2][1504] , \round_in[2][1503] , 
        \round_in[2][1502] , \round_in[2][1501] , \round_in[2][1500] , 
        \round_in[2][1499] , \round_in[2][1498] , \round_in[2][1497] , 
        \round_in[2][1496] , \round_in[2][1495] , \round_in[2][1494] , 
        \round_in[2][1493] , \round_in[2][1492] , \round_in[2][1491] , 
        \round_in[2][1490] , \round_in[2][1489] , \round_in[2][1488] , 
        \round_in[2][1487] , \round_in[2][1486] , \round_in[2][1485] , 
        \round_in[2][1484] , \round_in[2][1483] , \round_in[2][1482] , 
        \round_in[2][1481] , \round_in[2][1480] , \round_in[2][1479] , 
        \round_in[2][1478] , \round_in[2][1477] , \round_in[2][1476] , 
        \round_in[2][1475] , \round_in[2][1474] , \round_in[2][1473] , 
        \round_in[2][1472] , \round_in[2][1471] , \round_in[2][1470] , 
        \round_in[2][1469] , \round_in[2][1468] , \round_in[2][1467] , 
        \round_in[2][1466] , \round_in[2][1465] , \round_in[2][1464] , 
        \round_in[2][1463] , \round_in[2][1462] , \round_in[2][1461] , 
        \round_in[2][1460] , \round_in[2][1459] , \round_in[2][1458] , 
        \round_in[2][1457] , \round_in[2][1456] , \round_in[2][1455] , 
        \round_in[2][1454] , \round_in[2][1453] , \round_in[2][1452] , 
        \round_in[2][1451] , \round_in[2][1450] , \round_in[2][1449] , 
        \round_in[2][1448] , \round_in[2][1447] , \round_in[2][1446] , 
        \round_in[2][1445] , \round_in[2][1444] , \round_in[2][1443] , 
        \round_in[2][1442] , \round_in[2][1441] , \round_in[2][1440] , 
        \round_in[2][1439] , \round_in[2][1438] , \round_in[2][1437] , 
        \round_in[2][1436] , \round_in[2][1435] , \round_in[2][1434] , 
        \round_in[2][1433] , \round_in[2][1432] , \round_in[2][1431] , 
        \round_in[2][1430] , \round_in[2][1429] , \round_in[2][1428] , 
        \round_in[2][1427] , \round_in[2][1426] , \round_in[2][1425] , 
        \round_in[2][1424] , \round_in[2][1423] , \round_in[2][1422] , 
        \round_in[2][1421] , \round_in[2][1420] , \round_in[2][1419] , 
        \round_in[2][1418] , \round_in[2][1417] , \round_in[2][1416] , 
        \round_in[2][1415] , \round_in[2][1414] , \round_in[2][1413] , 
        \round_in[2][1412] , \round_in[2][1411] , \round_in[2][1410] , 
        \round_in[2][1409] , \round_in[2][1408] , \round_in[2][1407] , 
        \round_in[2][1406] , \round_in[2][1405] , \round_in[2][1404] , 
        \round_in[2][1403] , \round_in[2][1402] , \round_in[2][1401] , 
        \round_in[2][1400] , \round_in[2][1399] , \round_in[2][1398] , 
        \round_in[2][1397] , \round_in[2][1396] , \round_in[2][1395] , 
        \round_in[2][1394] , \round_in[2][1393] , \round_in[2][1392] , 
        \round_in[2][1391] , \round_in[2][1390] , \round_in[2][1389] , 
        \round_in[2][1388] , \round_in[2][1387] , \round_in[2][1386] , 
        \round_in[2][1385] , \round_in[2][1384] , \round_in[2][1383] , 
        \round_in[2][1382] , \round_in[2][1381] , \round_in[2][1380] , 
        \round_in[2][1379] , \round_in[2][1378] , \round_in[2][1377] , 
        \round_in[2][1376] , \round_in[2][1375] , \round_in[2][1374] , 
        \round_in[2][1373] , \round_in[2][1372] , \round_in[2][1371] , 
        \round_in[2][1370] , \round_in[2][1369] , \round_in[2][1368] , 
        \round_in[2][1367] , \round_in[2][1366] , \round_in[2][1365] , 
        \round_in[2][1364] , \round_in[2][1363] , \round_in[2][1362] , 
        \round_in[2][1361] , \round_in[2][1360] , \round_in[2][1359] , 
        \round_in[2][1358] , \round_in[2][1357] , \round_in[2][1356] , 
        \round_in[2][1355] , \round_in[2][1354] , \round_in[2][1353] , 
        \round_in[2][1352] , \round_in[2][1351] , \round_in[2][1350] , 
        \round_in[2][1349] , \round_in[2][1348] , \round_in[2][1347] , 
        \round_in[2][1346] , \round_in[2][1345] , \round_in[2][1344] , 
        \round_in[2][1343] , \round_in[2][1342] , \round_in[2][1341] , 
        \round_in[2][1340] , \round_in[2][1339] , \round_in[2][1338] , 
        \round_in[2][1337] , \round_in[2][1336] , \round_in[2][1335] , 
        \round_in[2][1334] , \round_in[2][1333] , \round_in[2][1332] , 
        \round_in[2][1331] , \round_in[2][1330] , \round_in[2][1329] , 
        \round_in[2][1328] , \round_in[2][1327] , \round_in[2][1326] , 
        \round_in[2][1325] , \round_in[2][1324] , \round_in[2][1323] , 
        \round_in[2][1322] , \round_in[2][1321] , \round_in[2][1320] , 
        \round_in[2][1319] , \round_in[2][1318] , \round_in[2][1317] , 
        \round_in[2][1316] , \round_in[2][1315] , \round_in[2][1314] , 
        \round_in[2][1313] , \round_in[2][1312] , \round_in[2][1311] , 
        \round_in[2][1310] , \round_in[2][1309] , \round_in[2][1308] , 
        \round_in[2][1307] , \round_in[2][1306] , \round_in[2][1305] , 
        \round_in[2][1304] , \round_in[2][1303] , \round_in[2][1302] , 
        \round_in[2][1301] , \round_in[2][1300] , \round_in[2][1299] , 
        \round_in[2][1298] , \round_in[2][1297] , \round_in[2][1296] , 
        \round_in[2][1295] , \round_in[2][1294] , \round_in[2][1293] , 
        \round_in[2][1292] , \round_in[2][1291] , \round_in[2][1290] , 
        \round_in[2][1289] , \round_in[2][1288] , \round_in[2][1287] , 
        \round_in[2][1286] , \round_in[2][1285] , \round_in[2][1284] , 
        \round_in[2][1283] , \round_in[2][1282] , \round_in[2][1281] , 
        \round_in[2][1280] , \round_in[2][1279] , \round_in[2][1278] , 
        \round_in[2][1277] , \round_in[2][1276] , \round_in[2][1275] , 
        \round_in[2][1274] , \round_in[2][1273] , \round_in[2][1272] , 
        \round_in[2][1271] , \round_in[2][1270] , \round_in[2][1269] , 
        \round_in[2][1268] , \round_in[2][1267] , \round_in[2][1266] , 
        \round_in[2][1265] , \round_in[2][1264] , \round_in[2][1263] , 
        \round_in[2][1262] , \round_in[2][1261] , \round_in[2][1260] , 
        \round_in[2][1259] , \round_in[2][1258] , \round_in[2][1257] , 
        \round_in[2][1256] , \round_in[2][1255] , \round_in[2][1254] , 
        \round_in[2][1253] , \round_in[2][1252] , \round_in[2][1251] , 
        \round_in[2][1250] , \round_in[2][1249] , \round_in[2][1248] , 
        \round_in[2][1247] , \round_in[2][1246] , \round_in[2][1245] , 
        \round_in[2][1244] , \round_in[2][1243] , \round_in[2][1242] , 
        \round_in[2][1241] , \round_in[2][1240] , \round_in[2][1239] , 
        \round_in[2][1238] , \round_in[2][1237] , \round_in[2][1236] , 
        \round_in[2][1235] , \round_in[2][1234] , \round_in[2][1233] , 
        \round_in[2][1232] , \round_in[2][1231] , \round_in[2][1230] , 
        \round_in[2][1229] , \round_in[2][1228] , \round_in[2][1227] , 
        \round_in[2][1226] , \round_in[2][1225] , \round_in[2][1224] , 
        \round_in[2][1223] , \round_in[2][1222] , \round_in[2][1221] , 
        \round_in[2][1220] , \round_in[2][1219] , \round_in[2][1218] , 
        \round_in[2][1217] , \round_in[2][1216] , \round_in[2][1215] , 
        \round_in[2][1214] , \round_in[2][1213] , \round_in[2][1212] , 
        \round_in[2][1211] , \round_in[2][1210] , \round_in[2][1209] , 
        \round_in[2][1208] , \round_in[2][1207] , \round_in[2][1206] , 
        \round_in[2][1205] , \round_in[2][1204] , \round_in[2][1203] , 
        \round_in[2][1202] , \round_in[2][1201] , \round_in[2][1200] , 
        \round_in[2][1199] , \round_in[2][1198] , \round_in[2][1197] , 
        \round_in[2][1196] , \round_in[2][1195] , \round_in[2][1194] , 
        \round_in[2][1193] , \round_in[2][1192] , \round_in[2][1191] , 
        \round_in[2][1190] , \round_in[2][1189] , \round_in[2][1188] , 
        \round_in[2][1187] , \round_in[2][1186] , \round_in[2][1185] , 
        \round_in[2][1184] , \round_in[2][1183] , \round_in[2][1182] , 
        \round_in[2][1181] , \round_in[2][1180] , \round_in[2][1179] , 
        \round_in[2][1178] , \round_in[2][1177] , \round_in[2][1176] , 
        \round_in[2][1175] , \round_in[2][1174] , \round_in[2][1173] , 
        \round_in[2][1172] , \round_in[2][1171] , \round_in[2][1170] , 
        \round_in[2][1169] , \round_in[2][1168] , \round_in[2][1167] , 
        \round_in[2][1166] , \round_in[2][1165] , \round_in[2][1164] , 
        \round_in[2][1163] , \round_in[2][1162] , \round_in[2][1161] , 
        \round_in[2][1160] , \round_in[2][1159] , \round_in[2][1158] , 
        \round_in[2][1157] , \round_in[2][1156] , \round_in[2][1155] , 
        \round_in[2][1154] , \round_in[2][1153] , \round_in[2][1152] , 
        \round_in[2][1151] , \round_in[2][1150] , \round_in[2][1149] , 
        \round_in[2][1148] , \round_in[2][1147] , \round_in[2][1146] , 
        \round_in[2][1145] , \round_in[2][1144] , \round_in[2][1143] , 
        \round_in[2][1142] , \round_in[2][1141] , \round_in[2][1140] , 
        \round_in[2][1139] , \round_in[2][1138] , \round_in[2][1137] , 
        \round_in[2][1136] , \round_in[2][1135] , \round_in[2][1134] , 
        \round_in[2][1133] , \round_in[2][1132] , \round_in[2][1131] , 
        \round_in[2][1130] , \round_in[2][1129] , \round_in[2][1128] , 
        \round_in[2][1127] , \round_in[2][1126] , \round_in[2][1125] , 
        \round_in[2][1124] , \round_in[2][1123] , \round_in[2][1122] , 
        \round_in[2][1121] , \round_in[2][1120] , \round_in[2][1119] , 
        \round_in[2][1118] , \round_in[2][1117] , \round_in[2][1116] , 
        \round_in[2][1115] , \round_in[2][1114] , \round_in[2][1113] , 
        \round_in[2][1112] , \round_in[2][1111] , \round_in[2][1110] , 
        \round_in[2][1109] , \round_in[2][1108] , \round_in[2][1107] , 
        \round_in[2][1106] , \round_in[2][1105] , \round_in[2][1104] , 
        \round_in[2][1103] , \round_in[2][1102] , \round_in[2][1101] , 
        \round_in[2][1100] , \round_in[2][1099] , \round_in[2][1098] , 
        \round_in[2][1097] , \round_in[2][1096] , \round_in[2][1095] , 
        \round_in[2][1094] , \round_in[2][1093] , \round_in[2][1092] , 
        \round_in[2][1091] , \round_in[2][1090] , \round_in[2][1089] , 
        \round_in[2][1088] , \round_in[2][1087] , \round_in[2][1086] , 
        \round_in[2][1085] , \round_in[2][1084] , \round_in[2][1083] , 
        \round_in[2][1082] , \round_in[2][1081] , \round_in[2][1080] , 
        \round_in[2][1079] , \round_in[2][1078] , \round_in[2][1077] , 
        \round_in[2][1076] , \round_in[2][1075] , \round_in[2][1074] , 
        \round_in[2][1073] , \round_in[2][1072] , \round_in[2][1071] , 
        \round_in[2][1070] , \round_in[2][1069] , \round_in[2][1068] , 
        \round_in[2][1067] , \round_in[2][1066] , \round_in[2][1065] , 
        \round_in[2][1064] , \round_in[2][1063] , \round_in[2][1062] , 
        \round_in[2][1061] , \round_in[2][1060] , \round_in[2][1059] , 
        \round_in[2][1058] , \round_in[2][1057] , \round_in[2][1056] , 
        \round_in[2][1055] , \round_in[2][1054] , \round_in[2][1053] , 
        \round_in[2][1052] , \round_in[2][1051] , \round_in[2][1050] , 
        \round_in[2][1049] , \round_in[2][1048] , \round_in[2][1047] , 
        \round_in[2][1046] , \round_in[2][1045] , \round_in[2][1044] , 
        \round_in[2][1043] , \round_in[2][1042] , \round_in[2][1041] , 
        \round_in[2][1040] , \round_in[2][1039] , \round_in[2][1038] , 
        \round_in[2][1037] , \round_in[2][1036] , \round_in[2][1035] , 
        \round_in[2][1034] , \round_in[2][1033] , \round_in[2][1032] , 
        \round_in[2][1031] , \round_in[2][1030] , \round_in[2][1029] , 
        \round_in[2][1028] , \round_in[2][1027] , \round_in[2][1026] , 
        \round_in[2][1025] , \round_in[2][1024] , \round_in[2][1023] , 
        \round_in[2][1022] , \round_in[2][1021] , \round_in[2][1020] , 
        \round_in[2][1019] , \round_in[2][1018] , \round_in[2][1017] , 
        \round_in[2][1016] , \round_in[2][1015] , \round_in[2][1014] , 
        \round_in[2][1013] , \round_in[2][1012] , \round_in[2][1011] , 
        \round_in[2][1010] , \round_in[2][1009] , \round_in[2][1008] , 
        \round_in[2][1007] , \round_in[2][1006] , \round_in[2][1005] , 
        \round_in[2][1004] , \round_in[2][1003] , \round_in[2][1002] , 
        \round_in[2][1001] , \round_in[2][1000] , \round_in[2][999] , 
        \round_in[2][998] , \round_in[2][997] , \round_in[2][996] , 
        \round_in[2][995] , \round_in[2][994] , \round_in[2][993] , 
        \round_in[2][992] , \round_in[2][991] , \round_in[2][990] , 
        \round_in[2][989] , \round_in[2][988] , \round_in[2][987] , 
        \round_in[2][986] , \round_in[2][985] , \round_in[2][984] , 
        \round_in[2][983] , \round_in[2][982] , \round_in[2][981] , 
        \round_in[2][980] , \round_in[2][979] , \round_in[2][978] , 
        \round_in[2][977] , \round_in[2][976] , \round_in[2][975] , 
        \round_in[2][974] , \round_in[2][973] , \round_in[2][972] , 
        \round_in[2][971] , \round_in[2][970] , \round_in[2][969] , 
        \round_in[2][968] , \round_in[2][967] , \round_in[2][966] , 
        \round_in[2][965] , \round_in[2][964] , \round_in[2][963] , 
        \round_in[2][962] , \round_in[2][961] , \round_in[2][960] , 
        \round_in[2][959] , \round_in[2][958] , \round_in[2][957] , 
        \round_in[2][956] , \round_in[2][955] , \round_in[2][954] , 
        \round_in[2][953] , \round_in[2][952] , \round_in[2][951] , 
        \round_in[2][950] , \round_in[2][949] , \round_in[2][948] , 
        \round_in[2][947] , \round_in[2][946] , \round_in[2][945] , 
        \round_in[2][944] , \round_in[2][943] , \round_in[2][942] , 
        \round_in[2][941] , \round_in[2][940] , \round_in[2][939] , 
        \round_in[2][938] , \round_in[2][937] , \round_in[2][936] , 
        \round_in[2][935] , \round_in[2][934] , \round_in[2][933] , 
        \round_in[2][932] , \round_in[2][931] , \round_in[2][930] , 
        \round_in[2][929] , \round_in[2][928] , \round_in[2][927] , 
        \round_in[2][926] , \round_in[2][925] , \round_in[2][924] , 
        \round_in[2][923] , \round_in[2][922] , \round_in[2][921] , 
        \round_in[2][920] , \round_in[2][919] , \round_in[2][918] , 
        \round_in[2][917] , \round_in[2][916] , \round_in[2][915] , 
        \round_in[2][914] , \round_in[2][913] , \round_in[2][912] , 
        \round_in[2][911] , \round_in[2][910] , \round_in[2][909] , 
        \round_in[2][908] , \round_in[2][907] , \round_in[2][906] , 
        \round_in[2][905] , \round_in[2][904] , \round_in[2][903] , 
        \round_in[2][902] , \round_in[2][901] , \round_in[2][900] , 
        \round_in[2][899] , \round_in[2][898] , \round_in[2][897] , 
        \round_in[2][896] , \round_in[2][895] , \round_in[2][894] , 
        \round_in[2][893] , \round_in[2][892] , \round_in[2][891] , 
        \round_in[2][890] , \round_in[2][889] , \round_in[2][888] , 
        \round_in[2][887] , \round_in[2][886] , \round_in[2][885] , 
        \round_in[2][884] , \round_in[2][883] , \round_in[2][882] , 
        \round_in[2][881] , \round_in[2][880] , \round_in[2][879] , 
        \round_in[2][878] , \round_in[2][877] , \round_in[2][876] , 
        \round_in[2][875] , \round_in[2][874] , \round_in[2][873] , 
        \round_in[2][872] , \round_in[2][871] , \round_in[2][870] , 
        \round_in[2][869] , \round_in[2][868] , \round_in[2][867] , 
        \round_in[2][866] , \round_in[2][865] , \round_in[2][864] , 
        \round_in[2][863] , \round_in[2][862] , \round_in[2][861] , 
        \round_in[2][860] , \round_in[2][859] , \round_in[2][858] , 
        \round_in[2][857] , \round_in[2][856] , \round_in[2][855] , 
        \round_in[2][854] , \round_in[2][853] , \round_in[2][852] , 
        \round_in[2][851] , \round_in[2][850] , \round_in[2][849] , 
        \round_in[2][848] , \round_in[2][847] , \round_in[2][846] , 
        \round_in[2][845] , \round_in[2][844] , \round_in[2][843] , 
        \round_in[2][842] , \round_in[2][841] , \round_in[2][840] , 
        \round_in[2][839] , \round_in[2][838] , \round_in[2][837] , 
        \round_in[2][836] , \round_in[2][835] , \round_in[2][834] , 
        \round_in[2][833] , \round_in[2][832] , \round_in[2][831] , 
        \round_in[2][830] , \round_in[2][829] , \round_in[2][828] , 
        \round_in[2][827] , \round_in[2][826] , \round_in[2][825] , 
        \round_in[2][824] , \round_in[2][823] , \round_in[2][822] , 
        \round_in[2][821] , \round_in[2][820] , \round_in[2][819] , 
        \round_in[2][818] , \round_in[2][817] , \round_in[2][816] , 
        \round_in[2][815] , \round_in[2][814] , \round_in[2][813] , 
        \round_in[2][812] , \round_in[2][811] , \round_in[2][810] , 
        \round_in[2][809] , \round_in[2][808] , \round_in[2][807] , 
        \round_in[2][806] , \round_in[2][805] , \round_in[2][804] , 
        \round_in[2][803] , \round_in[2][802] , \round_in[2][801] , 
        \round_in[2][800] , \round_in[2][799] , \round_in[2][798] , 
        \round_in[2][797] , \round_in[2][796] , \round_in[2][795] , 
        \round_in[2][794] , \round_in[2][793] , \round_in[2][792] , 
        \round_in[2][791] , \round_in[2][790] , \round_in[2][789] , 
        \round_in[2][788] , \round_in[2][787] , \round_in[2][786] , 
        \round_in[2][785] , \round_in[2][784] , \round_in[2][783] , 
        \round_in[2][782] , \round_in[2][781] , \round_in[2][780] , 
        \round_in[2][779] , \round_in[2][778] , \round_in[2][777] , 
        \round_in[2][776] , \round_in[2][775] , \round_in[2][774] , 
        \round_in[2][773] , \round_in[2][772] , \round_in[2][771] , 
        \round_in[2][770] , \round_in[2][769] , \round_in[2][768] , 
        \round_in[2][767] , \round_in[2][766] , \round_in[2][765] , 
        \round_in[2][764] , \round_in[2][763] , \round_in[2][762] , 
        \round_in[2][761] , \round_in[2][760] , \round_in[2][759] , 
        \round_in[2][758] , \round_in[2][757] , \round_in[2][756] , 
        \round_in[2][755] , \round_in[2][754] , \round_in[2][753] , 
        \round_in[2][752] , \round_in[2][751] , \round_in[2][750] , 
        \round_in[2][749] , \round_in[2][748] , \round_in[2][747] , 
        \round_in[2][746] , \round_in[2][745] , \round_in[2][744] , 
        \round_in[2][743] , \round_in[2][742] , \round_in[2][741] , 
        \round_in[2][740] , \round_in[2][739] , \round_in[2][738] , 
        \round_in[2][737] , \round_in[2][736] , \round_in[2][735] , 
        \round_in[2][734] , \round_in[2][733] , \round_in[2][732] , 
        \round_in[2][731] , \round_in[2][730] , \round_in[2][729] , 
        \round_in[2][728] , \round_in[2][727] , \round_in[2][726] , 
        \round_in[2][725] , \round_in[2][724] , \round_in[2][723] , 
        \round_in[2][722] , \round_in[2][721] , \round_in[2][720] , 
        \round_in[2][719] , \round_in[2][718] , \round_in[2][717] , 
        \round_in[2][716] , \round_in[2][715] , \round_in[2][714] , 
        \round_in[2][713] , \round_in[2][712] , \round_in[2][711] , 
        \round_in[2][710] , \round_in[2][709] , \round_in[2][708] , 
        \round_in[2][707] , \round_in[2][706] , \round_in[2][705] , 
        \round_in[2][704] , \round_in[2][703] , \round_in[2][702] , 
        \round_in[2][701] , \round_in[2][700] , \round_in[2][699] , 
        \round_in[2][698] , \round_in[2][697] , \round_in[2][696] , 
        \round_in[2][695] , \round_in[2][694] , \round_in[2][693] , 
        \round_in[2][692] , \round_in[2][691] , \round_in[2][690] , 
        \round_in[2][689] , \round_in[2][688] , \round_in[2][687] , 
        \round_in[2][686] , \round_in[2][685] , \round_in[2][684] , 
        \round_in[2][683] , \round_in[2][682] , \round_in[2][681] , 
        \round_in[2][680] , \round_in[2][679] , \round_in[2][678] , 
        \round_in[2][677] , \round_in[2][676] , \round_in[2][675] , 
        \round_in[2][674] , \round_in[2][673] , \round_in[2][672] , 
        \round_in[2][671] , \round_in[2][670] , \round_in[2][669] , 
        \round_in[2][668] , \round_in[2][667] , \round_in[2][666] , 
        \round_in[2][665] , \round_in[2][664] , \round_in[2][663] , 
        \round_in[2][662] , \round_in[2][661] , \round_in[2][660] , 
        \round_in[2][659] , \round_in[2][658] , \round_in[2][657] , 
        \round_in[2][656] , \round_in[2][655] , \round_in[2][654] , 
        \round_in[2][653] , \round_in[2][652] , \round_in[2][651] , 
        \round_in[2][650] , \round_in[2][649] , \round_in[2][648] , 
        \round_in[2][647] , \round_in[2][646] , \round_in[2][645] , 
        \round_in[2][644] , \round_in[2][643] , \round_in[2][642] , 
        \round_in[2][641] , \round_in[2][640] , \round_in[2][639] , 
        \round_in[2][638] , \round_in[2][637] , \round_in[2][636] , 
        \round_in[2][635] , \round_in[2][634] , \round_in[2][633] , 
        \round_in[2][632] , \round_in[2][631] , \round_in[2][630] , 
        \round_in[2][629] , \round_in[2][628] , \round_in[2][627] , 
        \round_in[2][626] , \round_in[2][625] , \round_in[2][624] , 
        \round_in[2][623] , \round_in[2][622] , \round_in[2][621] , 
        \round_in[2][620] , \round_in[2][619] , \round_in[2][618] , 
        \round_in[2][617] , \round_in[2][616] , \round_in[2][615] , 
        \round_in[2][614] , \round_in[2][613] , \round_in[2][612] , 
        \round_in[2][611] , \round_in[2][610] , \round_in[2][609] , 
        \round_in[2][608] , \round_in[2][607] , \round_in[2][606] , 
        \round_in[2][605] , \round_in[2][604] , \round_in[2][603] , 
        \round_in[2][602] , \round_in[2][601] , \round_in[2][600] , 
        \round_in[2][599] , \round_in[2][598] , \round_in[2][597] , 
        \round_in[2][596] , \round_in[2][595] , \round_in[2][594] , 
        \round_in[2][593] , \round_in[2][592] , \round_in[2][591] , 
        \round_in[2][590] , \round_in[2][589] , \round_in[2][588] , 
        \round_in[2][587] , \round_in[2][586] , \round_in[2][585] , 
        \round_in[2][584] , \round_in[2][583] , \round_in[2][582] , 
        \round_in[2][581] , \round_in[2][580] , \round_in[2][579] , 
        \round_in[2][578] , \round_in[2][577] , \round_in[2][576] , 
        \round_in[2][575] , \round_in[2][574] , \round_in[2][573] , 
        \round_in[2][572] , \round_in[2][571] , \round_in[2][570] , 
        \round_in[2][569] , \round_in[2][568] , \round_in[2][567] , 
        \round_in[2][566] , \round_in[2][565] , \round_in[2][564] , 
        \round_in[2][563] , \round_in[2][562] , \round_in[2][561] , 
        \round_in[2][560] , \round_in[2][559] , \round_in[2][558] , 
        \round_in[2][557] , \round_in[2][556] , \round_in[2][555] , 
        \round_in[2][554] , \round_in[2][553] , \round_in[2][552] , 
        \round_in[2][551] , \round_in[2][550] , \round_in[2][549] , 
        \round_in[2][548] , \round_in[2][547] , \round_in[2][546] , 
        \round_in[2][545] , \round_in[2][544] , \round_in[2][543] , 
        \round_in[2][542] , \round_in[2][541] , \round_in[2][540] , 
        \round_in[2][539] , \round_in[2][538] , \round_in[2][537] , 
        \round_in[2][536] , \round_in[2][535] , \round_in[2][534] , 
        \round_in[2][533] , \round_in[2][532] , \round_in[2][531] , 
        \round_in[2][530] , \round_in[2][529] , \round_in[2][528] , 
        \round_in[2][527] , \round_in[2][526] , \round_in[2][525] , 
        \round_in[2][524] , \round_in[2][523] , \round_in[2][522] , 
        \round_in[2][521] , \round_in[2][520] , \round_in[2][519] , 
        \round_in[2][518] , \round_in[2][517] , \round_in[2][516] , 
        \round_in[2][515] , \round_in[2][514] , \round_in[2][513] , 
        \round_in[2][512] , \round_in[2][511] , \round_in[2][510] , 
        \round_in[2][509] , \round_in[2][508] , \round_in[2][507] , 
        \round_in[2][506] , \round_in[2][505] , \round_in[2][504] , 
        \round_in[2][503] , \round_in[2][502] , \round_in[2][501] , 
        \round_in[2][500] , \round_in[2][499] , \round_in[2][498] , 
        \round_in[2][497] , \round_in[2][496] , \round_in[2][495] , 
        \round_in[2][494] , \round_in[2][493] , \round_in[2][492] , 
        \round_in[2][491] , \round_in[2][490] , \round_in[2][489] , 
        \round_in[2][488] , \round_in[2][487] , \round_in[2][486] , 
        \round_in[2][485] , \round_in[2][484] , \round_in[2][483] , 
        \round_in[2][482] , \round_in[2][481] , \round_in[2][480] , 
        \round_in[2][479] , \round_in[2][478] , \round_in[2][477] , 
        \round_in[2][476] , \round_in[2][475] , \round_in[2][474] , 
        \round_in[2][473] , \round_in[2][472] , \round_in[2][471] , 
        \round_in[2][470] , \round_in[2][469] , \round_in[2][468] , 
        \round_in[2][467] , \round_in[2][466] , \round_in[2][465] , 
        \round_in[2][464] , \round_in[2][463] , \round_in[2][462] , 
        \round_in[2][461] , \round_in[2][460] , \round_in[2][459] , 
        \round_in[2][458] , \round_in[2][457] , \round_in[2][456] , 
        \round_in[2][455] , \round_in[2][454] , \round_in[2][453] , 
        \round_in[2][452] , \round_in[2][451] , \round_in[2][450] , 
        \round_in[2][449] , \round_in[2][448] , \round_in[2][447] , 
        \round_in[2][446] , \round_in[2][445] , \round_in[2][444] , 
        \round_in[2][443] , \round_in[2][442] , \round_in[2][441] , 
        \round_in[2][440] , \round_in[2][439] , \round_in[2][438] , 
        \round_in[2][437] , \round_in[2][436] , \round_in[2][435] , 
        \round_in[2][434] , \round_in[2][433] , \round_in[2][432] , 
        \round_in[2][431] , \round_in[2][430] , \round_in[2][429] , 
        \round_in[2][428] , \round_in[2][427] , \round_in[2][426] , 
        \round_in[2][425] , \round_in[2][424] , \round_in[2][423] , 
        \round_in[2][422] , \round_in[2][421] , \round_in[2][420] , 
        \round_in[2][419] , \round_in[2][418] , \round_in[2][417] , 
        \round_in[2][416] , \round_in[2][415] , \round_in[2][414] , 
        \round_in[2][413] , \round_in[2][412] , \round_in[2][411] , 
        \round_in[2][410] , \round_in[2][409] , \round_in[2][408] , 
        \round_in[2][407] , \round_in[2][406] , \round_in[2][405] , 
        \round_in[2][404] , \round_in[2][403] , \round_in[2][402] , 
        \round_in[2][401] , \round_in[2][400] , \round_in[2][399] , 
        \round_in[2][398] , \round_in[2][397] , \round_in[2][396] , 
        \round_in[2][395] , \round_in[2][394] , \round_in[2][393] , 
        \round_in[2][392] , \round_in[2][391] , \round_in[2][390] , 
        \round_in[2][389] , \round_in[2][388] , \round_in[2][387] , 
        \round_in[2][386] , \round_in[2][385] , \round_in[2][384] , 
        \round_in[2][383] , \round_in[2][382] , \round_in[2][381] , 
        \round_in[2][380] , \round_in[2][379] , \round_in[2][378] , 
        \round_in[2][377] , \round_in[2][376] , \round_in[2][375] , 
        \round_in[2][374] , \round_in[2][373] , \round_in[2][372] , 
        \round_in[2][371] , \round_in[2][370] , \round_in[2][369] , 
        \round_in[2][368] , \round_in[2][367] , \round_in[2][366] , 
        \round_in[2][365] , \round_in[2][364] , \round_in[2][363] , 
        \round_in[2][362] , \round_in[2][361] , \round_in[2][360] , 
        \round_in[2][359] , \round_in[2][358] , \round_in[2][357] , 
        \round_in[2][356] , \round_in[2][355] , \round_in[2][354] , 
        \round_in[2][353] , \round_in[2][352] , \round_in[2][351] , 
        \round_in[2][350] , \round_in[2][349] , \round_in[2][348] , 
        \round_in[2][347] , \round_in[2][346] , \round_in[2][345] , 
        \round_in[2][344] , \round_in[2][343] , \round_in[2][342] , 
        \round_in[2][341] , \round_in[2][340] , \round_in[2][339] , 
        \round_in[2][338] , \round_in[2][337] , \round_in[2][336] , 
        \round_in[2][335] , \round_in[2][334] , \round_in[2][333] , 
        \round_in[2][332] , \round_in[2][331] , \round_in[2][330] , 
        \round_in[2][329] , \round_in[2][328] , \round_in[2][327] , 
        \round_in[2][326] , \round_in[2][325] , \round_in[2][324] , 
        \round_in[2][323] , \round_in[2][322] , \round_in[2][321] , 
        \round_in[2][320] , \round_in[2][319] , \round_in[2][318] , 
        \round_in[2][317] , \round_in[2][316] , \round_in[2][315] , 
        \round_in[2][314] , \round_in[2][313] , \round_in[2][312] , 
        \round_in[2][311] , \round_in[2][310] , \round_in[2][309] , 
        \round_in[2][308] , \round_in[2][307] , \round_in[2][306] , 
        \round_in[2][305] , \round_in[2][304] , \round_in[2][303] , 
        \round_in[2][302] , \round_in[2][301] , \round_in[2][300] , 
        \round_in[2][299] , \round_in[2][298] , \round_in[2][297] , 
        \round_in[2][296] , \round_in[2][295] , \round_in[2][294] , 
        \round_in[2][293] , \round_in[2][292] , \round_in[2][291] , 
        \round_in[2][290] , \round_in[2][289] , \round_in[2][288] , 
        \round_in[2][287] , \round_in[2][286] , \round_in[2][285] , 
        \round_in[2][284] , \round_in[2][283] , \round_in[2][282] , 
        \round_in[2][281] , \round_in[2][280] , \round_in[2][279] , 
        \round_in[2][278] , \round_in[2][277] , \round_in[2][276] , 
        \round_in[2][275] , \round_in[2][274] , \round_in[2][273] , 
        \round_in[2][272] , \round_in[2][271] , \round_in[2][270] , 
        \round_in[2][269] , \round_in[2][268] , \round_in[2][267] , 
        \round_in[2][266] , \round_in[2][265] , \round_in[2][264] , 
        \round_in[2][263] , \round_in[2][262] , \round_in[2][261] , 
        \round_in[2][260] , \round_in[2][259] , \round_in[2][258] , 
        \round_in[2][257] , \round_in[2][256] , \round_in[2][255] , 
        \round_in[2][254] , \round_in[2][253] , \round_in[2][252] , 
        \round_in[2][251] , \round_in[2][250] , \round_in[2][249] , 
        \round_in[2][248] , \round_in[2][247] , \round_in[2][246] , 
        \round_in[2][245] , \round_in[2][244] , \round_in[2][243] , 
        \round_in[2][242] , \round_in[2][241] , \round_in[2][240] , 
        \round_in[2][239] , \round_in[2][238] , \round_in[2][237] , 
        \round_in[2][236] , \round_in[2][235] , \round_in[2][234] , 
        \round_in[2][233] , \round_in[2][232] , \round_in[2][231] , 
        \round_in[2][230] , \round_in[2][229] , \round_in[2][228] , 
        \round_in[2][227] , \round_in[2][226] , \round_in[2][225] , 
        \round_in[2][224] , \round_in[2][223] , \round_in[2][222] , 
        \round_in[2][221] , \round_in[2][220] , \round_in[2][219] , 
        \round_in[2][218] , \round_in[2][217] , \round_in[2][216] , 
        \round_in[2][215] , \round_in[2][214] , \round_in[2][213] , 
        \round_in[2][212] , \round_in[2][211] , \round_in[2][210] , 
        \round_in[2][209] , \round_in[2][208] , \round_in[2][207] , 
        \round_in[2][206] , \round_in[2][205] , \round_in[2][204] , 
        \round_in[2][203] , \round_in[2][202] , \round_in[2][201] , 
        \round_in[2][200] , \round_in[2][199] , \round_in[2][198] , 
        \round_in[2][197] , \round_in[2][196] , \round_in[2][195] , 
        \round_in[2][194] , \round_in[2][193] , \round_in[2][192] , 
        \round_in[2][191] , \round_in[2][190] , \round_in[2][189] , 
        \round_in[2][188] , \round_in[2][187] , \round_in[2][186] , 
        \round_in[2][185] , \round_in[2][184] , \round_in[2][183] , 
        \round_in[2][182] , \round_in[2][181] , \round_in[2][180] , 
        \round_in[2][179] , \round_in[2][178] , \round_in[2][177] , 
        \round_in[2][176] , \round_in[2][175] , \round_in[2][174] , 
        \round_in[2][173] , \round_in[2][172] , \round_in[2][171] , 
        \round_in[2][170] , \round_in[2][169] , \round_in[2][168] , 
        \round_in[2][167] , \round_in[2][166] , \round_in[2][165] , 
        \round_in[2][164] , \round_in[2][163] , \round_in[2][162] , 
        \round_in[2][161] , \round_in[2][160] , \round_in[2][159] , 
        \round_in[2][158] , \round_in[2][157] , \round_in[2][156] , 
        \round_in[2][155] , \round_in[2][154] , \round_in[2][153] , 
        \round_in[2][152] , \round_in[2][151] , \round_in[2][150] , 
        \round_in[2][149] , \round_in[2][148] , \round_in[2][147] , 
        \round_in[2][146] , \round_in[2][145] , \round_in[2][144] , 
        \round_in[2][143] , \round_in[2][142] , \round_in[2][141] , 
        \round_in[2][140] , \round_in[2][139] , \round_in[2][138] , 
        \round_in[2][137] , \round_in[2][136] , \round_in[2][135] , 
        \round_in[2][134] , \round_in[2][133] , \round_in[2][132] , 
        \round_in[2][131] , \round_in[2][130] , \round_in[2][129] , 
        \round_in[2][128] , \round_in[2][127] , \round_in[2][126] , 
        \round_in[2][125] , \round_in[2][124] , \round_in[2][123] , 
        \round_in[2][122] , \round_in[2][121] , \round_in[2][120] , 
        \round_in[2][119] , \round_in[2][118] , \round_in[2][117] , 
        \round_in[2][116] , \round_in[2][115] , \round_in[2][114] , 
        \round_in[2][113] , \round_in[2][112] , \round_in[2][111] , 
        \round_in[2][110] , \round_in[2][109] , \round_in[2][108] , 
        \round_in[2][107] , \round_in[2][106] , \round_in[2][105] , 
        \round_in[2][104] , \round_in[2][103] , \round_in[2][102] , 
        \round_in[2][101] , \round_in[2][100] , \round_in[2][99] , 
        \round_in[2][98] , \round_in[2][97] , \round_in[2][96] , 
        \round_in[2][95] , \round_in[2][94] , \round_in[2][93] , 
        \round_in[2][92] , \round_in[2][91] , \round_in[2][90] , 
        \round_in[2][89] , \round_in[2][88] , \round_in[2][87] , 
        \round_in[2][86] , \round_in[2][85] , \round_in[2][84] , 
        \round_in[2][83] , \round_in[2][82] , \round_in[2][81] , 
        \round_in[2][80] , \round_in[2][79] , \round_in[2][78] , 
        \round_in[2][77] , \round_in[2][76] , \round_in[2][75] , 
        \round_in[2][74] , \round_in[2][73] , \round_in[2][72] , 
        \round_in[2][71] , \round_in[2][70] , \round_in[2][69] , 
        \round_in[2][68] , \round_in[2][67] , \round_in[2][66] , 
        \round_in[2][65] , \round_in[2][64] , \round_in[2][63] , 
        \round_in[2][62] , \round_in[2][61] , \round_in[2][60] , 
        \round_in[2][59] , \round_in[2][58] , \round_in[2][57] , 
        \round_in[2][56] , \round_in[2][55] , \round_in[2][54] , 
        \round_in[2][53] , \round_in[2][52] , \round_in[2][51] , 
        \round_in[2][50] , \round_in[2][49] , \round_in[2][48] , 
        \round_in[2][47] , \round_in[2][46] , \round_in[2][45] , 
        \round_in[2][44] , \round_in[2][43] , \round_in[2][42] , 
        \round_in[2][41] , \round_in[2][40] , \round_in[2][39] , 
        \round_in[2][38] , \round_in[2][37] , \round_in[2][36] , 
        \round_in[2][35] , \round_in[2][34] , \round_in[2][33] , 
        \round_in[2][32] , \round_in[2][31] , \round_in[2][30] , 
        \round_in[2][29] , \round_in[2][28] , \round_in[2][27] , 
        \round_in[2][26] , \round_in[2][25] , \round_in[2][24] , 
        \round_in[2][23] , \round_in[2][22] , \round_in[2][21] , 
        \round_in[2][20] , \round_in[2][19] , \round_in[2][18] , 
        \round_in[2][17] , \round_in[2][16] , \round_in[2][15] , 
        \round_in[2][14] , \round_in[2][13] , \round_in[2][12] , 
        \round_in[2][11] , \round_in[2][10] , \round_in[2][9] , 
        \round_in[2][8] , \round_in[2][7] , \round_in[2][6] , \round_in[2][5] , 
        \round_in[2][4] , \round_in[2][3] , \round_in[2][2] , \round_in[2][1] , 
        \round_in[2][0] }) );
  round_4 \ROUND[2].round_  ( .in({\round_in[2][1599] , \round_in[2][1598] , 
        \round_in[2][1597] , \round_in[2][1596] , \round_in[2][1595] , 
        \round_in[2][1594] , \round_in[2][1593] , \round_in[2][1592] , 
        \round_in[2][1591] , \round_in[2][1590] , \round_in[2][1589] , 
        \round_in[2][1588] , \round_in[2][1587] , \round_in[2][1586] , 
        \round_in[2][1585] , \round_in[2][1584] , \round_in[2][1583] , 
        \round_in[2][1582] , \round_in[2][1581] , \round_in[2][1580] , 
        \round_in[2][1579] , \round_in[2][1578] , \round_in[2][1577] , 
        \round_in[2][1576] , \round_in[2][1575] , \round_in[2][1574] , 
        \round_in[2][1573] , \round_in[2][1572] , \round_in[2][1571] , 
        \round_in[2][1570] , \round_in[2][1569] , \round_in[2][1568] , 
        \round_in[2][1567] , \round_in[2][1566] , \round_in[2][1565] , 
        \round_in[2][1564] , \round_in[2][1563] , \round_in[2][1562] , 
        \round_in[2][1561] , \round_in[2][1560] , \round_in[2][1559] , 
        \round_in[2][1558] , \round_in[2][1557] , \round_in[2][1556] , 
        \round_in[2][1555] , \round_in[2][1554] , \round_in[2][1553] , 
        \round_in[2][1552] , \round_in[2][1551] , \round_in[2][1550] , 
        \round_in[2][1549] , \round_in[2][1548] , \round_in[2][1547] , 
        \round_in[2][1546] , \round_in[2][1545] , \round_in[2][1544] , 
        \round_in[2][1543] , \round_in[2][1542] , \round_in[2][1541] , 
        \round_in[2][1540] , \round_in[2][1539] , \round_in[2][1538] , 
        \round_in[2][1537] , \round_in[2][1536] , \round_in[2][1535] , 
        \round_in[2][1534] , \round_in[2][1533] , \round_in[2][1532] , 
        \round_in[2][1531] , \round_in[2][1530] , \round_in[2][1529] , 
        \round_in[2][1528] , \round_in[2][1527] , \round_in[2][1526] , 
        \round_in[2][1525] , \round_in[2][1524] , \round_in[2][1523] , 
        \round_in[2][1522] , \round_in[2][1521] , \round_in[2][1520] , 
        \round_in[2][1519] , \round_in[2][1518] , \round_in[2][1517] , 
        \round_in[2][1516] , \round_in[2][1515] , \round_in[2][1514] , 
        \round_in[2][1513] , \round_in[2][1512] , \round_in[2][1511] , 
        \round_in[2][1510] , \round_in[2][1509] , \round_in[2][1508] , 
        \round_in[2][1507] , \round_in[2][1506] , \round_in[2][1505] , 
        \round_in[2][1504] , \round_in[2][1503] , \round_in[2][1502] , 
        \round_in[2][1501] , \round_in[2][1500] , \round_in[2][1499] , 
        \round_in[2][1498] , \round_in[2][1497] , \round_in[2][1496] , 
        \round_in[2][1495] , \round_in[2][1494] , \round_in[2][1493] , 
        \round_in[2][1492] , \round_in[2][1491] , \round_in[2][1490] , 
        \round_in[2][1489] , \round_in[2][1488] , \round_in[2][1487] , 
        \round_in[2][1486] , \round_in[2][1485] , \round_in[2][1484] , 
        \round_in[2][1483] , \round_in[2][1482] , \round_in[2][1481] , 
        \round_in[2][1480] , \round_in[2][1479] , \round_in[2][1478] , 
        \round_in[2][1477] , \round_in[2][1476] , \round_in[2][1475] , 
        \round_in[2][1474] , \round_in[2][1473] , \round_in[2][1472] , 
        \round_in[2][1471] , \round_in[2][1470] , \round_in[2][1469] , 
        \round_in[2][1468] , \round_in[2][1467] , \round_in[2][1466] , 
        \round_in[2][1465] , \round_in[2][1464] , \round_in[2][1463] , 
        \round_in[2][1462] , \round_in[2][1461] , \round_in[2][1460] , 
        \round_in[2][1459] , \round_in[2][1458] , \round_in[2][1457] , 
        \round_in[2][1456] , \round_in[2][1455] , \round_in[2][1454] , 
        \round_in[2][1453] , \round_in[2][1452] , \round_in[2][1451] , 
        \round_in[2][1450] , \round_in[2][1449] , \round_in[2][1448] , 
        \round_in[2][1447] , \round_in[2][1446] , \round_in[2][1445] , 
        \round_in[2][1444] , \round_in[2][1443] , \round_in[2][1442] , 
        \round_in[2][1441] , \round_in[2][1440] , \round_in[2][1439] , 
        \round_in[2][1438] , \round_in[2][1437] , \round_in[2][1436] , 
        \round_in[2][1435] , \round_in[2][1434] , \round_in[2][1433] , 
        \round_in[2][1432] , \round_in[2][1431] , \round_in[2][1430] , 
        \round_in[2][1429] , \round_in[2][1428] , \round_in[2][1427] , 
        \round_in[2][1426] , \round_in[2][1425] , \round_in[2][1424] , 
        \round_in[2][1423] , \round_in[2][1422] , \round_in[2][1421] , 
        \round_in[2][1420] , \round_in[2][1419] , \round_in[2][1418] , 
        \round_in[2][1417] , \round_in[2][1416] , \round_in[2][1415] , 
        \round_in[2][1414] , \round_in[2][1413] , \round_in[2][1412] , 
        \round_in[2][1411] , \round_in[2][1410] , \round_in[2][1409] , 
        \round_in[2][1408] , \round_in[2][1407] , \round_in[2][1406] , 
        \round_in[2][1405] , \round_in[2][1404] , \round_in[2][1403] , 
        \round_in[2][1402] , \round_in[2][1401] , \round_in[2][1400] , 
        \round_in[2][1399] , \round_in[2][1398] , \round_in[2][1397] , 
        \round_in[2][1396] , \round_in[2][1395] , \round_in[2][1394] , 
        \round_in[2][1393] , \round_in[2][1392] , \round_in[2][1391] , 
        \round_in[2][1390] , \round_in[2][1389] , \round_in[2][1388] , 
        \round_in[2][1387] , \round_in[2][1386] , \round_in[2][1385] , 
        \round_in[2][1384] , \round_in[2][1383] , \round_in[2][1382] , 
        \round_in[2][1381] , \round_in[2][1380] , \round_in[2][1379] , 
        \round_in[2][1378] , \round_in[2][1377] , \round_in[2][1376] , 
        \round_in[2][1375] , \round_in[2][1374] , \round_in[2][1373] , 
        \round_in[2][1372] , \round_in[2][1371] , \round_in[2][1370] , 
        \round_in[2][1369] , \round_in[2][1368] , \round_in[2][1367] , 
        \round_in[2][1366] , \round_in[2][1365] , \round_in[2][1364] , 
        \round_in[2][1363] , \round_in[2][1362] , \round_in[2][1361] , 
        \round_in[2][1360] , \round_in[2][1359] , \round_in[2][1358] , 
        \round_in[2][1357] , \round_in[2][1356] , \round_in[2][1355] , 
        \round_in[2][1354] , \round_in[2][1353] , \round_in[2][1352] , 
        \round_in[2][1351] , \round_in[2][1350] , \round_in[2][1349] , 
        \round_in[2][1348] , \round_in[2][1347] , \round_in[2][1346] , 
        \round_in[2][1345] , \round_in[2][1344] , \round_in[2][1343] , 
        \round_in[2][1342] , \round_in[2][1341] , \round_in[2][1340] , 
        \round_in[2][1339] , \round_in[2][1338] , \round_in[2][1337] , 
        \round_in[2][1336] , \round_in[2][1335] , \round_in[2][1334] , 
        \round_in[2][1333] , \round_in[2][1332] , \round_in[2][1331] , 
        \round_in[2][1330] , \round_in[2][1329] , \round_in[2][1328] , 
        \round_in[2][1327] , \round_in[2][1326] , \round_in[2][1325] , 
        \round_in[2][1324] , \round_in[2][1323] , \round_in[2][1322] , 
        \round_in[2][1321] , \round_in[2][1320] , \round_in[2][1319] , 
        \round_in[2][1318] , \round_in[2][1317] , \round_in[2][1316] , 
        \round_in[2][1315] , \round_in[2][1314] , \round_in[2][1313] , 
        \round_in[2][1312] , \round_in[2][1311] , \round_in[2][1310] , 
        \round_in[2][1309] , \round_in[2][1308] , \round_in[2][1307] , 
        \round_in[2][1306] , \round_in[2][1305] , \round_in[2][1304] , 
        \round_in[2][1303] , \round_in[2][1302] , \round_in[2][1301] , 
        \round_in[2][1300] , \round_in[2][1299] , \round_in[2][1298] , 
        \round_in[2][1297] , \round_in[2][1296] , \round_in[2][1295] , 
        \round_in[2][1294] , \round_in[2][1293] , \round_in[2][1292] , 
        \round_in[2][1291] , \round_in[2][1290] , \round_in[2][1289] , 
        \round_in[2][1288] , \round_in[2][1287] , \round_in[2][1286] , 
        \round_in[2][1285] , \round_in[2][1284] , \round_in[2][1283] , 
        \round_in[2][1282] , \round_in[2][1281] , \round_in[2][1280] , 
        \round_in[2][1279] , \round_in[2][1278] , \round_in[2][1277] , 
        \round_in[2][1276] , \round_in[2][1275] , \round_in[2][1274] , 
        \round_in[2][1273] , \round_in[2][1272] , \round_in[2][1271] , 
        \round_in[2][1270] , \round_in[2][1269] , \round_in[2][1268] , 
        \round_in[2][1267] , \round_in[2][1266] , \round_in[2][1265] , 
        \round_in[2][1264] , \round_in[2][1263] , \round_in[2][1262] , 
        \round_in[2][1261] , \round_in[2][1260] , \round_in[2][1259] , 
        \round_in[2][1258] , \round_in[2][1257] , \round_in[2][1256] , 
        \round_in[2][1255] , \round_in[2][1254] , \round_in[2][1253] , 
        \round_in[2][1252] , \round_in[2][1251] , \round_in[2][1250] , 
        \round_in[2][1249] , \round_in[2][1248] , \round_in[2][1247] , 
        \round_in[2][1246] , \round_in[2][1245] , \round_in[2][1244] , 
        \round_in[2][1243] , \round_in[2][1242] , \round_in[2][1241] , 
        \round_in[2][1240] , \round_in[2][1239] , \round_in[2][1238] , 
        \round_in[2][1237] , \round_in[2][1236] , \round_in[2][1235] , 
        \round_in[2][1234] , \round_in[2][1233] , \round_in[2][1232] , 
        \round_in[2][1231] , \round_in[2][1230] , \round_in[2][1229] , 
        \round_in[2][1228] , \round_in[2][1227] , \round_in[2][1226] , 
        \round_in[2][1225] , \round_in[2][1224] , \round_in[2][1223] , 
        \round_in[2][1222] , \round_in[2][1221] , \round_in[2][1220] , 
        \round_in[2][1219] , \round_in[2][1218] , \round_in[2][1217] , 
        \round_in[2][1216] , \round_in[2][1215] , \round_in[2][1214] , 
        \round_in[2][1213] , \round_in[2][1212] , \round_in[2][1211] , 
        \round_in[2][1210] , \round_in[2][1209] , \round_in[2][1208] , 
        \round_in[2][1207] , \round_in[2][1206] , \round_in[2][1205] , 
        \round_in[2][1204] , \round_in[2][1203] , \round_in[2][1202] , 
        \round_in[2][1201] , \round_in[2][1200] , \round_in[2][1199] , 
        \round_in[2][1198] , \round_in[2][1197] , \round_in[2][1196] , 
        \round_in[2][1195] , \round_in[2][1194] , \round_in[2][1193] , 
        \round_in[2][1192] , \round_in[2][1191] , \round_in[2][1190] , 
        \round_in[2][1189] , \round_in[2][1188] , \round_in[2][1187] , 
        \round_in[2][1186] , \round_in[2][1185] , \round_in[2][1184] , 
        \round_in[2][1183] , \round_in[2][1182] , \round_in[2][1181] , 
        \round_in[2][1180] , \round_in[2][1179] , \round_in[2][1178] , 
        \round_in[2][1177] , \round_in[2][1176] , \round_in[2][1175] , 
        \round_in[2][1174] , \round_in[2][1173] , \round_in[2][1172] , 
        \round_in[2][1171] , \round_in[2][1170] , \round_in[2][1169] , 
        \round_in[2][1168] , \round_in[2][1167] , \round_in[2][1166] , 
        \round_in[2][1165] , \round_in[2][1164] , \round_in[2][1163] , 
        \round_in[2][1162] , \round_in[2][1161] , \round_in[2][1160] , 
        \round_in[2][1159] , \round_in[2][1158] , \round_in[2][1157] , 
        \round_in[2][1156] , \round_in[2][1155] , \round_in[2][1154] , 
        \round_in[2][1153] , \round_in[2][1152] , \round_in[2][1151] , 
        \round_in[2][1150] , \round_in[2][1149] , \round_in[2][1148] , 
        \round_in[2][1147] , \round_in[2][1146] , \round_in[2][1145] , 
        \round_in[2][1144] , \round_in[2][1143] , \round_in[2][1142] , 
        \round_in[2][1141] , \round_in[2][1140] , \round_in[2][1139] , 
        \round_in[2][1138] , \round_in[2][1137] , \round_in[2][1136] , 
        \round_in[2][1135] , \round_in[2][1134] , \round_in[2][1133] , 
        \round_in[2][1132] , \round_in[2][1131] , \round_in[2][1130] , 
        \round_in[2][1129] , \round_in[2][1128] , \round_in[2][1127] , 
        \round_in[2][1126] , \round_in[2][1125] , \round_in[2][1124] , 
        \round_in[2][1123] , \round_in[2][1122] , \round_in[2][1121] , 
        \round_in[2][1120] , \round_in[2][1119] , \round_in[2][1118] , 
        \round_in[2][1117] , \round_in[2][1116] , \round_in[2][1115] , 
        \round_in[2][1114] , \round_in[2][1113] , \round_in[2][1112] , 
        \round_in[2][1111] , \round_in[2][1110] , \round_in[2][1109] , 
        \round_in[2][1108] , \round_in[2][1107] , \round_in[2][1106] , 
        \round_in[2][1105] , \round_in[2][1104] , \round_in[2][1103] , 
        \round_in[2][1102] , \round_in[2][1101] , \round_in[2][1100] , 
        \round_in[2][1099] , \round_in[2][1098] , \round_in[2][1097] , 
        \round_in[2][1096] , \round_in[2][1095] , \round_in[2][1094] , 
        \round_in[2][1093] , \round_in[2][1092] , \round_in[2][1091] , 
        \round_in[2][1090] , \round_in[2][1089] , \round_in[2][1088] , 
        \round_in[2][1087] , \round_in[2][1086] , \round_in[2][1085] , 
        \round_in[2][1084] , \round_in[2][1083] , \round_in[2][1082] , 
        \round_in[2][1081] , \round_in[2][1080] , \round_in[2][1079] , 
        \round_in[2][1078] , \round_in[2][1077] , \round_in[2][1076] , 
        \round_in[2][1075] , \round_in[2][1074] , \round_in[2][1073] , 
        \round_in[2][1072] , \round_in[2][1071] , \round_in[2][1070] , 
        \round_in[2][1069] , \round_in[2][1068] , \round_in[2][1067] , 
        \round_in[2][1066] , \round_in[2][1065] , \round_in[2][1064] , 
        \round_in[2][1063] , \round_in[2][1062] , \round_in[2][1061] , 
        \round_in[2][1060] , \round_in[2][1059] , \round_in[2][1058] , 
        \round_in[2][1057] , \round_in[2][1056] , \round_in[2][1055] , 
        \round_in[2][1054] , \round_in[2][1053] , \round_in[2][1052] , 
        \round_in[2][1051] , \round_in[2][1050] , \round_in[2][1049] , 
        \round_in[2][1048] , \round_in[2][1047] , \round_in[2][1046] , 
        \round_in[2][1045] , \round_in[2][1044] , \round_in[2][1043] , 
        \round_in[2][1042] , \round_in[2][1041] , \round_in[2][1040] , 
        \round_in[2][1039] , \round_in[2][1038] , \round_in[2][1037] , 
        \round_in[2][1036] , \round_in[2][1035] , \round_in[2][1034] , 
        \round_in[2][1033] , \round_in[2][1032] , \round_in[2][1031] , 
        \round_in[2][1030] , \round_in[2][1029] , \round_in[2][1028] , 
        \round_in[2][1027] , \round_in[2][1026] , \round_in[2][1025] , 
        \round_in[2][1024] , \round_in[2][1023] , \round_in[2][1022] , 
        \round_in[2][1021] , \round_in[2][1020] , \round_in[2][1019] , 
        \round_in[2][1018] , \round_in[2][1017] , \round_in[2][1016] , 
        \round_in[2][1015] , \round_in[2][1014] , \round_in[2][1013] , 
        \round_in[2][1012] , \round_in[2][1011] , \round_in[2][1010] , 
        \round_in[2][1009] , \round_in[2][1008] , \round_in[2][1007] , 
        \round_in[2][1006] , \round_in[2][1005] , \round_in[2][1004] , 
        \round_in[2][1003] , \round_in[2][1002] , \round_in[2][1001] , 
        \round_in[2][1000] , \round_in[2][999] , \round_in[2][998] , 
        \round_in[2][997] , \round_in[2][996] , \round_in[2][995] , 
        \round_in[2][994] , \round_in[2][993] , \round_in[2][992] , 
        \round_in[2][991] , \round_in[2][990] , \round_in[2][989] , 
        \round_in[2][988] , \round_in[2][987] , \round_in[2][986] , 
        \round_in[2][985] , \round_in[2][984] , \round_in[2][983] , 
        \round_in[2][982] , \round_in[2][981] , \round_in[2][980] , 
        \round_in[2][979] , \round_in[2][978] , \round_in[2][977] , 
        \round_in[2][976] , \round_in[2][975] , \round_in[2][974] , 
        \round_in[2][973] , \round_in[2][972] , \round_in[2][971] , 
        \round_in[2][970] , \round_in[2][969] , \round_in[2][968] , 
        \round_in[2][967] , \round_in[2][966] , \round_in[2][965] , 
        \round_in[2][964] , \round_in[2][963] , \round_in[2][962] , 
        \round_in[2][961] , \round_in[2][960] , \round_in[2][959] , 
        \round_in[2][958] , \round_in[2][957] , \round_in[2][956] , 
        \round_in[2][955] , \round_in[2][954] , \round_in[2][953] , 
        \round_in[2][952] , \round_in[2][951] , \round_in[2][950] , 
        \round_in[2][949] , \round_in[2][948] , \round_in[2][947] , 
        \round_in[2][946] , \round_in[2][945] , \round_in[2][944] , 
        \round_in[2][943] , \round_in[2][942] , \round_in[2][941] , 
        \round_in[2][940] , \round_in[2][939] , \round_in[2][938] , 
        \round_in[2][937] , \round_in[2][936] , \round_in[2][935] , 
        \round_in[2][934] , \round_in[2][933] , \round_in[2][932] , 
        \round_in[2][931] , \round_in[2][930] , \round_in[2][929] , 
        \round_in[2][928] , \round_in[2][927] , \round_in[2][926] , 
        \round_in[2][925] , \round_in[2][924] , \round_in[2][923] , 
        \round_in[2][922] , \round_in[2][921] , \round_in[2][920] , 
        \round_in[2][919] , \round_in[2][918] , \round_in[2][917] , 
        \round_in[2][916] , \round_in[2][915] , \round_in[2][914] , 
        \round_in[2][913] , \round_in[2][912] , \round_in[2][911] , 
        \round_in[2][910] , \round_in[2][909] , \round_in[2][908] , 
        \round_in[2][907] , \round_in[2][906] , \round_in[2][905] , 
        \round_in[2][904] , \round_in[2][903] , \round_in[2][902] , 
        \round_in[2][901] , \round_in[2][900] , \round_in[2][899] , 
        \round_in[2][898] , \round_in[2][897] , \round_in[2][896] , 
        \round_in[2][895] , \round_in[2][894] , \round_in[2][893] , 
        \round_in[2][892] , \round_in[2][891] , \round_in[2][890] , 
        \round_in[2][889] , \round_in[2][888] , \round_in[2][887] , 
        \round_in[2][886] , \round_in[2][885] , \round_in[2][884] , 
        \round_in[2][883] , \round_in[2][882] , \round_in[2][881] , 
        \round_in[2][880] , \round_in[2][879] , \round_in[2][878] , 
        \round_in[2][877] , \round_in[2][876] , \round_in[2][875] , 
        \round_in[2][874] , \round_in[2][873] , \round_in[2][872] , 
        \round_in[2][871] , \round_in[2][870] , \round_in[2][869] , 
        \round_in[2][868] , \round_in[2][867] , \round_in[2][866] , 
        \round_in[2][865] , \round_in[2][864] , \round_in[2][863] , 
        \round_in[2][862] , \round_in[2][861] , \round_in[2][860] , 
        \round_in[2][859] , \round_in[2][858] , \round_in[2][857] , 
        \round_in[2][856] , \round_in[2][855] , \round_in[2][854] , 
        \round_in[2][853] , \round_in[2][852] , \round_in[2][851] , 
        \round_in[2][850] , \round_in[2][849] , \round_in[2][848] , 
        \round_in[2][847] , \round_in[2][846] , \round_in[2][845] , 
        \round_in[2][844] , \round_in[2][843] , \round_in[2][842] , 
        \round_in[2][841] , \round_in[2][840] , \round_in[2][839] , 
        \round_in[2][838] , \round_in[2][837] , \round_in[2][836] , 
        \round_in[2][835] , \round_in[2][834] , \round_in[2][833] , 
        \round_in[2][832] , \round_in[2][831] , \round_in[2][830] , 
        \round_in[2][829] , \round_in[2][828] , \round_in[2][827] , 
        \round_in[2][826] , \round_in[2][825] , \round_in[2][824] , 
        \round_in[2][823] , \round_in[2][822] , \round_in[2][821] , 
        \round_in[2][820] , \round_in[2][819] , \round_in[2][818] , 
        \round_in[2][817] , \round_in[2][816] , \round_in[2][815] , 
        \round_in[2][814] , \round_in[2][813] , \round_in[2][812] , 
        \round_in[2][811] , \round_in[2][810] , \round_in[2][809] , 
        \round_in[2][808] , \round_in[2][807] , \round_in[2][806] , 
        \round_in[2][805] , \round_in[2][804] , \round_in[2][803] , 
        \round_in[2][802] , \round_in[2][801] , \round_in[2][800] , 
        \round_in[2][799] , \round_in[2][798] , \round_in[2][797] , 
        \round_in[2][796] , \round_in[2][795] , \round_in[2][794] , 
        \round_in[2][793] , \round_in[2][792] , \round_in[2][791] , 
        \round_in[2][790] , \round_in[2][789] , \round_in[2][788] , 
        \round_in[2][787] , \round_in[2][786] , \round_in[2][785] , 
        \round_in[2][784] , \round_in[2][783] , \round_in[2][782] , 
        \round_in[2][781] , \round_in[2][780] , \round_in[2][779] , 
        \round_in[2][778] , \round_in[2][777] , \round_in[2][776] , 
        \round_in[2][775] , \round_in[2][774] , \round_in[2][773] , 
        \round_in[2][772] , \round_in[2][771] , \round_in[2][770] , 
        \round_in[2][769] , \round_in[2][768] , \round_in[2][767] , 
        \round_in[2][766] , \round_in[2][765] , \round_in[2][764] , 
        \round_in[2][763] , \round_in[2][762] , \round_in[2][761] , 
        \round_in[2][760] , \round_in[2][759] , \round_in[2][758] , 
        \round_in[2][757] , \round_in[2][756] , \round_in[2][755] , 
        \round_in[2][754] , \round_in[2][753] , \round_in[2][752] , 
        \round_in[2][751] , \round_in[2][750] , \round_in[2][749] , 
        \round_in[2][748] , \round_in[2][747] , \round_in[2][746] , 
        \round_in[2][745] , \round_in[2][744] , \round_in[2][743] , 
        \round_in[2][742] , \round_in[2][741] , \round_in[2][740] , 
        \round_in[2][739] , \round_in[2][738] , \round_in[2][737] , 
        \round_in[2][736] , \round_in[2][735] , \round_in[2][734] , 
        \round_in[2][733] , \round_in[2][732] , \round_in[2][731] , 
        \round_in[2][730] , \round_in[2][729] , \round_in[2][728] , 
        \round_in[2][727] , \round_in[2][726] , \round_in[2][725] , 
        \round_in[2][724] , \round_in[2][723] , \round_in[2][722] , 
        \round_in[2][721] , \round_in[2][720] , \round_in[2][719] , 
        \round_in[2][718] , \round_in[2][717] , \round_in[2][716] , 
        \round_in[2][715] , \round_in[2][714] , \round_in[2][713] , 
        \round_in[2][712] , \round_in[2][711] , \round_in[2][710] , 
        \round_in[2][709] , \round_in[2][708] , \round_in[2][707] , 
        \round_in[2][706] , \round_in[2][705] , \round_in[2][704] , 
        \round_in[2][703] , \round_in[2][702] , \round_in[2][701] , 
        \round_in[2][700] , \round_in[2][699] , \round_in[2][698] , 
        \round_in[2][697] , \round_in[2][696] , \round_in[2][695] , 
        \round_in[2][694] , \round_in[2][693] , \round_in[2][692] , 
        \round_in[2][691] , \round_in[2][690] , \round_in[2][689] , 
        \round_in[2][688] , \round_in[2][687] , \round_in[2][686] , 
        \round_in[2][685] , \round_in[2][684] , \round_in[2][683] , 
        \round_in[2][682] , \round_in[2][681] , \round_in[2][680] , 
        \round_in[2][679] , \round_in[2][678] , \round_in[2][677] , 
        \round_in[2][676] , \round_in[2][675] , \round_in[2][674] , 
        \round_in[2][673] , \round_in[2][672] , \round_in[2][671] , 
        \round_in[2][670] , \round_in[2][669] , \round_in[2][668] , 
        \round_in[2][667] , \round_in[2][666] , \round_in[2][665] , 
        \round_in[2][664] , \round_in[2][663] , \round_in[2][662] , 
        \round_in[2][661] , \round_in[2][660] , \round_in[2][659] , 
        \round_in[2][658] , \round_in[2][657] , \round_in[2][656] , 
        \round_in[2][655] , \round_in[2][654] , \round_in[2][653] , 
        \round_in[2][652] , \round_in[2][651] , \round_in[2][650] , 
        \round_in[2][649] , \round_in[2][648] , \round_in[2][647] , 
        \round_in[2][646] , \round_in[2][645] , \round_in[2][644] , 
        \round_in[2][643] , \round_in[2][642] , \round_in[2][641] , 
        \round_in[2][640] , \round_in[2][639] , \round_in[2][638] , 
        \round_in[2][637] , \round_in[2][636] , \round_in[2][635] , 
        \round_in[2][634] , \round_in[2][633] , \round_in[2][632] , 
        \round_in[2][631] , \round_in[2][630] , \round_in[2][629] , 
        \round_in[2][628] , \round_in[2][627] , \round_in[2][626] , 
        \round_in[2][625] , \round_in[2][624] , \round_in[2][623] , 
        \round_in[2][622] , \round_in[2][621] , \round_in[2][620] , 
        \round_in[2][619] , \round_in[2][618] , \round_in[2][617] , 
        \round_in[2][616] , \round_in[2][615] , \round_in[2][614] , 
        \round_in[2][613] , \round_in[2][612] , \round_in[2][611] , 
        \round_in[2][610] , \round_in[2][609] , \round_in[2][608] , 
        \round_in[2][607] , \round_in[2][606] , \round_in[2][605] , 
        \round_in[2][604] , \round_in[2][603] , \round_in[2][602] , 
        \round_in[2][601] , \round_in[2][600] , \round_in[2][599] , 
        \round_in[2][598] , \round_in[2][597] , \round_in[2][596] , 
        \round_in[2][595] , \round_in[2][594] , \round_in[2][593] , 
        \round_in[2][592] , \round_in[2][591] , \round_in[2][590] , 
        \round_in[2][589] , \round_in[2][588] , \round_in[2][587] , 
        \round_in[2][586] , \round_in[2][585] , \round_in[2][584] , 
        \round_in[2][583] , \round_in[2][582] , \round_in[2][581] , 
        \round_in[2][580] , \round_in[2][579] , \round_in[2][578] , 
        \round_in[2][577] , \round_in[2][576] , \round_in[2][575] , 
        \round_in[2][574] , \round_in[2][573] , \round_in[2][572] , 
        \round_in[2][571] , \round_in[2][570] , \round_in[2][569] , 
        \round_in[2][568] , \round_in[2][567] , \round_in[2][566] , 
        \round_in[2][565] , \round_in[2][564] , \round_in[2][563] , 
        \round_in[2][562] , \round_in[2][561] , \round_in[2][560] , 
        \round_in[2][559] , \round_in[2][558] , \round_in[2][557] , 
        \round_in[2][556] , \round_in[2][555] , \round_in[2][554] , 
        \round_in[2][553] , \round_in[2][552] , \round_in[2][551] , 
        \round_in[2][550] , \round_in[2][549] , \round_in[2][548] , 
        \round_in[2][547] , \round_in[2][546] , \round_in[2][545] , 
        \round_in[2][544] , \round_in[2][543] , \round_in[2][542] , 
        \round_in[2][541] , \round_in[2][540] , \round_in[2][539] , 
        \round_in[2][538] , \round_in[2][537] , \round_in[2][536] , 
        \round_in[2][535] , \round_in[2][534] , \round_in[2][533] , 
        \round_in[2][532] , \round_in[2][531] , \round_in[2][530] , 
        \round_in[2][529] , \round_in[2][528] , \round_in[2][527] , 
        \round_in[2][526] , \round_in[2][525] , \round_in[2][524] , 
        \round_in[2][523] , \round_in[2][522] , \round_in[2][521] , 
        \round_in[2][520] , \round_in[2][519] , \round_in[2][518] , 
        \round_in[2][517] , \round_in[2][516] , \round_in[2][515] , 
        \round_in[2][514] , \round_in[2][513] , \round_in[2][512] , 
        \round_in[2][511] , \round_in[2][510] , \round_in[2][509] , 
        \round_in[2][508] , \round_in[2][507] , \round_in[2][506] , 
        \round_in[2][505] , \round_in[2][504] , \round_in[2][503] , 
        \round_in[2][502] , \round_in[2][501] , \round_in[2][500] , 
        \round_in[2][499] , \round_in[2][498] , \round_in[2][497] , 
        \round_in[2][496] , \round_in[2][495] , \round_in[2][494] , 
        \round_in[2][493] , \round_in[2][492] , \round_in[2][491] , 
        \round_in[2][490] , \round_in[2][489] , \round_in[2][488] , 
        \round_in[2][487] , \round_in[2][486] , \round_in[2][485] , 
        \round_in[2][484] , \round_in[2][483] , \round_in[2][482] , 
        \round_in[2][481] , \round_in[2][480] , \round_in[2][479] , 
        \round_in[2][478] , \round_in[2][477] , \round_in[2][476] , 
        \round_in[2][475] , \round_in[2][474] , \round_in[2][473] , 
        \round_in[2][472] , \round_in[2][471] , \round_in[2][470] , 
        \round_in[2][469] , \round_in[2][468] , \round_in[2][467] , 
        \round_in[2][466] , \round_in[2][465] , \round_in[2][464] , 
        \round_in[2][463] , \round_in[2][462] , \round_in[2][461] , 
        \round_in[2][460] , \round_in[2][459] , \round_in[2][458] , 
        \round_in[2][457] , \round_in[2][456] , \round_in[2][455] , 
        \round_in[2][454] , \round_in[2][453] , \round_in[2][452] , 
        \round_in[2][451] , \round_in[2][450] , \round_in[2][449] , 
        \round_in[2][448] , \round_in[2][447] , \round_in[2][446] , 
        \round_in[2][445] , \round_in[2][444] , \round_in[2][443] , 
        \round_in[2][442] , \round_in[2][441] , \round_in[2][440] , 
        \round_in[2][439] , \round_in[2][438] , \round_in[2][437] , 
        \round_in[2][436] , \round_in[2][435] , \round_in[2][434] , 
        \round_in[2][433] , \round_in[2][432] , \round_in[2][431] , 
        \round_in[2][430] , \round_in[2][429] , \round_in[2][428] , 
        \round_in[2][427] , \round_in[2][426] , \round_in[2][425] , 
        \round_in[2][424] , \round_in[2][423] , \round_in[2][422] , 
        \round_in[2][421] , \round_in[2][420] , \round_in[2][419] , 
        \round_in[2][418] , \round_in[2][417] , \round_in[2][416] , 
        \round_in[2][415] , \round_in[2][414] , \round_in[2][413] , 
        \round_in[2][412] , \round_in[2][411] , \round_in[2][410] , 
        \round_in[2][409] , \round_in[2][408] , \round_in[2][407] , 
        \round_in[2][406] , \round_in[2][405] , \round_in[2][404] , 
        \round_in[2][403] , \round_in[2][402] , \round_in[2][401] , 
        \round_in[2][400] , \round_in[2][399] , \round_in[2][398] , 
        \round_in[2][397] , \round_in[2][396] , \round_in[2][395] , 
        \round_in[2][394] , \round_in[2][393] , \round_in[2][392] , 
        \round_in[2][391] , \round_in[2][390] , \round_in[2][389] , 
        \round_in[2][388] , \round_in[2][387] , \round_in[2][386] , 
        \round_in[2][385] , \round_in[2][384] , \round_in[2][383] , 
        \round_in[2][382] , \round_in[2][381] , \round_in[2][380] , 
        \round_in[2][379] , \round_in[2][378] , \round_in[2][377] , 
        \round_in[2][376] , \round_in[2][375] , \round_in[2][374] , 
        \round_in[2][373] , \round_in[2][372] , \round_in[2][371] , 
        \round_in[2][370] , \round_in[2][369] , \round_in[2][368] , 
        \round_in[2][367] , \round_in[2][366] , \round_in[2][365] , 
        \round_in[2][364] , \round_in[2][363] , \round_in[2][362] , 
        \round_in[2][361] , \round_in[2][360] , \round_in[2][359] , 
        \round_in[2][358] , \round_in[2][357] , \round_in[2][356] , 
        \round_in[2][355] , \round_in[2][354] , \round_in[2][353] , 
        \round_in[2][352] , \round_in[2][351] , \round_in[2][350] , 
        \round_in[2][349] , \round_in[2][348] , \round_in[2][347] , 
        \round_in[2][346] , \round_in[2][345] , \round_in[2][344] , 
        \round_in[2][343] , \round_in[2][342] , \round_in[2][341] , 
        \round_in[2][340] , \round_in[2][339] , \round_in[2][338] , 
        \round_in[2][337] , \round_in[2][336] , \round_in[2][335] , 
        \round_in[2][334] , \round_in[2][333] , \round_in[2][332] , 
        \round_in[2][331] , \round_in[2][330] , \round_in[2][329] , 
        \round_in[2][328] , \round_in[2][327] , \round_in[2][326] , 
        \round_in[2][325] , \round_in[2][324] , \round_in[2][323] , 
        \round_in[2][322] , \round_in[2][321] , \round_in[2][320] , 
        \round_in[2][319] , \round_in[2][318] , \round_in[2][317] , 
        \round_in[2][316] , \round_in[2][315] , \round_in[2][314] , 
        \round_in[2][313] , \round_in[2][312] , \round_in[2][311] , 
        \round_in[2][310] , \round_in[2][309] , \round_in[2][308] , 
        \round_in[2][307] , \round_in[2][306] , \round_in[2][305] , 
        \round_in[2][304] , \round_in[2][303] , \round_in[2][302] , 
        \round_in[2][301] , \round_in[2][300] , \round_in[2][299] , 
        \round_in[2][298] , \round_in[2][297] , \round_in[2][296] , 
        \round_in[2][295] , \round_in[2][294] , \round_in[2][293] , 
        \round_in[2][292] , \round_in[2][291] , \round_in[2][290] , 
        \round_in[2][289] , \round_in[2][288] , \round_in[2][287] , 
        \round_in[2][286] , \round_in[2][285] , \round_in[2][284] , 
        \round_in[2][283] , \round_in[2][282] , \round_in[2][281] , 
        \round_in[2][280] , \round_in[2][279] , \round_in[2][278] , 
        \round_in[2][277] , \round_in[2][276] , \round_in[2][275] , 
        \round_in[2][274] , \round_in[2][273] , \round_in[2][272] , 
        \round_in[2][271] , \round_in[2][270] , \round_in[2][269] , 
        \round_in[2][268] , \round_in[2][267] , \round_in[2][266] , 
        \round_in[2][265] , \round_in[2][264] , \round_in[2][263] , 
        \round_in[2][262] , \round_in[2][261] , \round_in[2][260] , 
        \round_in[2][259] , \round_in[2][258] , \round_in[2][257] , 
        \round_in[2][256] , \round_in[2][255] , \round_in[2][254] , 
        \round_in[2][253] , \round_in[2][252] , \round_in[2][251] , 
        \round_in[2][250] , \round_in[2][249] , \round_in[2][248] , 
        \round_in[2][247] , \round_in[2][246] , \round_in[2][245] , 
        \round_in[2][244] , \round_in[2][243] , \round_in[2][242] , 
        \round_in[2][241] , \round_in[2][240] , \round_in[2][239] , 
        \round_in[2][238] , \round_in[2][237] , \round_in[2][236] , 
        \round_in[2][235] , \round_in[2][234] , \round_in[2][233] , 
        \round_in[2][232] , \round_in[2][231] , \round_in[2][230] , 
        \round_in[2][229] , \round_in[2][228] , \round_in[2][227] , 
        \round_in[2][226] , \round_in[2][225] , \round_in[2][224] , 
        \round_in[2][223] , \round_in[2][222] , \round_in[2][221] , 
        \round_in[2][220] , \round_in[2][219] , \round_in[2][218] , 
        \round_in[2][217] , \round_in[2][216] , \round_in[2][215] , 
        \round_in[2][214] , \round_in[2][213] , \round_in[2][212] , 
        \round_in[2][211] , \round_in[2][210] , \round_in[2][209] , 
        \round_in[2][208] , \round_in[2][207] , \round_in[2][206] , 
        \round_in[2][205] , \round_in[2][204] , \round_in[2][203] , 
        \round_in[2][202] , \round_in[2][201] , \round_in[2][200] , 
        \round_in[2][199] , \round_in[2][198] , \round_in[2][197] , 
        \round_in[2][196] , \round_in[2][195] , \round_in[2][194] , 
        \round_in[2][193] , \round_in[2][192] , \round_in[2][191] , 
        \round_in[2][190] , \round_in[2][189] , \round_in[2][188] , 
        \round_in[2][187] , \round_in[2][186] , \round_in[2][185] , 
        \round_in[2][184] , \round_in[2][183] , \round_in[2][182] , 
        \round_in[2][181] , \round_in[2][180] , \round_in[2][179] , 
        \round_in[2][178] , \round_in[2][177] , \round_in[2][176] , 
        \round_in[2][175] , \round_in[2][174] , \round_in[2][173] , 
        \round_in[2][172] , \round_in[2][171] , \round_in[2][170] , 
        \round_in[2][169] , \round_in[2][168] , \round_in[2][167] , 
        \round_in[2][166] , \round_in[2][165] , \round_in[2][164] , 
        \round_in[2][163] , \round_in[2][162] , \round_in[2][161] , 
        \round_in[2][160] , \round_in[2][159] , \round_in[2][158] , 
        \round_in[2][157] , \round_in[2][156] , \round_in[2][155] , 
        \round_in[2][154] , \round_in[2][153] , \round_in[2][152] , 
        \round_in[2][151] , \round_in[2][150] , \round_in[2][149] , 
        \round_in[2][148] , \round_in[2][147] , \round_in[2][146] , 
        \round_in[2][145] , \round_in[2][144] , \round_in[2][143] , 
        \round_in[2][142] , \round_in[2][141] , \round_in[2][140] , 
        \round_in[2][139] , \round_in[2][138] , \round_in[2][137] , 
        \round_in[2][136] , \round_in[2][135] , \round_in[2][134] , 
        \round_in[2][133] , \round_in[2][132] , \round_in[2][131] , 
        \round_in[2][130] , \round_in[2][129] , \round_in[2][128] , 
        \round_in[2][127] , \round_in[2][126] , \round_in[2][125] , 
        \round_in[2][124] , \round_in[2][123] , \round_in[2][122] , 
        \round_in[2][121] , \round_in[2][120] , \round_in[2][119] , 
        \round_in[2][118] , \round_in[2][117] , \round_in[2][116] , 
        \round_in[2][115] , \round_in[2][114] , \round_in[2][113] , 
        \round_in[2][112] , \round_in[2][111] , \round_in[2][110] , 
        \round_in[2][109] , \round_in[2][108] , \round_in[2][107] , 
        \round_in[2][106] , \round_in[2][105] , \round_in[2][104] , 
        \round_in[2][103] , \round_in[2][102] , \round_in[2][101] , 
        \round_in[2][100] , \round_in[2][99] , \round_in[2][98] , 
        \round_in[2][97] , \round_in[2][96] , \round_in[2][95] , 
        \round_in[2][94] , \round_in[2][93] , \round_in[2][92] , 
        \round_in[2][91] , \round_in[2][90] , \round_in[2][89] , 
        \round_in[2][88] , \round_in[2][87] , \round_in[2][86] , 
        \round_in[2][85] , \round_in[2][84] , \round_in[2][83] , 
        \round_in[2][82] , \round_in[2][81] , \round_in[2][80] , 
        \round_in[2][79] , \round_in[2][78] , \round_in[2][77] , 
        \round_in[2][76] , \round_in[2][75] , \round_in[2][74] , 
        \round_in[2][73] , \round_in[2][72] , \round_in[2][71] , 
        \round_in[2][70] , \round_in[2][69] , \round_in[2][68] , 
        \round_in[2][67] , \round_in[2][66] , \round_in[2][65] , 
        \round_in[2][64] , \round_in[2][63] , \round_in[2][62] , 
        \round_in[2][61] , \round_in[2][60] , \round_in[2][59] , 
        \round_in[2][58] , \round_in[2][57] , \round_in[2][56] , 
        \round_in[2][55] , \round_in[2][54] , \round_in[2][53] , 
        \round_in[2][52] , \round_in[2][51] , \round_in[2][50] , 
        \round_in[2][49] , \round_in[2][48] , \round_in[2][47] , 
        \round_in[2][46] , \round_in[2][45] , \round_in[2][44] , 
        \round_in[2][43] , \round_in[2][42] , \round_in[2][41] , 
        \round_in[2][40] , \round_in[2][39] , \round_in[2][38] , 
        \round_in[2][37] , \round_in[2][36] , \round_in[2][35] , 
        \round_in[2][34] , \round_in[2][33] , \round_in[2][32] , 
        \round_in[2][31] , \round_in[2][30] , \round_in[2][29] , 
        \round_in[2][28] , \round_in[2][27] , \round_in[2][26] , 
        \round_in[2][25] , \round_in[2][24] , \round_in[2][23] , 
        \round_in[2][22] , \round_in[2][21] , \round_in[2][20] , 
        \round_in[2][19] , \round_in[2][18] , \round_in[2][17] , 
        \round_in[2][16] , \round_in[2][15] , \round_in[2][14] , 
        \round_in[2][13] , \round_in[2][12] , \round_in[2][11] , 
        \round_in[2][10] , \round_in[2][9] , \round_in[2][8] , 
        \round_in[2][7] , \round_in[2][6] , \round_in[2][5] , \round_in[2][4] , 
        \round_in[2][3] , \round_in[2][2] , \round_in[2][1] , \round_in[2][0] }), .round_const({\RCONST[2].rconst_/N62 , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, \RCONST[2].rconst_/N57 , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        \RCONST[2].rconst_/N47 , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        \RCONST[2].rconst_/N62 , 1'b0, 1'b0, 1'b0, \RCONST[2].rconst_/N28 , 
        1'b0, \RCONST[2].rconst_/N18 , \rc[2][0] }), .out({\round_in[3][1599] , 
        \round_in[3][1598] , \round_in[3][1597] , \round_in[3][1596] , 
        \round_in[3][1595] , \round_in[3][1594] , \round_in[3][1593] , 
        \round_in[3][1592] , \round_in[3][1591] , \round_in[3][1590] , 
        \round_in[3][1589] , \round_in[3][1588] , \round_in[3][1587] , 
        \round_in[3][1586] , \round_in[3][1585] , \round_in[3][1584] , 
        \round_in[3][1583] , \round_in[3][1582] , \round_in[3][1581] , 
        \round_in[3][1580] , \round_in[3][1579] , \round_in[3][1578] , 
        \round_in[3][1577] , \round_in[3][1576] , \round_in[3][1575] , 
        \round_in[3][1574] , \round_in[3][1573] , \round_in[3][1572] , 
        \round_in[3][1571] , \round_in[3][1570] , \round_in[3][1569] , 
        \round_in[3][1568] , \round_in[3][1567] , \round_in[3][1566] , 
        \round_in[3][1565] , \round_in[3][1564] , \round_in[3][1563] , 
        \round_in[3][1562] , \round_in[3][1561] , \round_in[3][1560] , 
        \round_in[3][1559] , \round_in[3][1558] , \round_in[3][1557] , 
        \round_in[3][1556] , \round_in[3][1555] , \round_in[3][1554] , 
        \round_in[3][1553] , \round_in[3][1552] , \round_in[3][1551] , 
        \round_in[3][1550] , \round_in[3][1549] , \round_in[3][1548] , 
        \round_in[3][1547] , \round_in[3][1546] , \round_in[3][1545] , 
        \round_in[3][1544] , \round_in[3][1543] , \round_in[3][1542] , 
        \round_in[3][1541] , \round_in[3][1540] , \round_in[3][1539] , 
        \round_in[3][1538] , \round_in[3][1537] , \round_in[3][1536] , 
        \round_in[3][1535] , \round_in[3][1534] , \round_in[3][1533] , 
        \round_in[3][1532] , \round_in[3][1531] , \round_in[3][1530] , 
        \round_in[3][1529] , \round_in[3][1528] , \round_in[3][1527] , 
        \round_in[3][1526] , \round_in[3][1525] , \round_in[3][1524] , 
        \round_in[3][1523] , \round_in[3][1522] , \round_in[3][1521] , 
        \round_in[3][1520] , \round_in[3][1519] , \round_in[3][1518] , 
        \round_in[3][1517] , \round_in[3][1516] , \round_in[3][1515] , 
        \round_in[3][1514] , \round_in[3][1513] , \round_in[3][1512] , 
        \round_in[3][1511] , \round_in[3][1510] , \round_in[3][1509] , 
        \round_in[3][1508] , \round_in[3][1507] , \round_in[3][1506] , 
        \round_in[3][1505] , \round_in[3][1504] , \round_in[3][1503] , 
        \round_in[3][1502] , \round_in[3][1501] , \round_in[3][1500] , 
        \round_in[3][1499] , \round_in[3][1498] , \round_in[3][1497] , 
        \round_in[3][1496] , \round_in[3][1495] , \round_in[3][1494] , 
        \round_in[3][1493] , \round_in[3][1492] , \round_in[3][1491] , 
        \round_in[3][1490] , \round_in[3][1489] , \round_in[3][1488] , 
        \round_in[3][1487] , \round_in[3][1486] , \round_in[3][1485] , 
        \round_in[3][1484] , \round_in[3][1483] , \round_in[3][1482] , 
        \round_in[3][1481] , \round_in[3][1480] , \round_in[3][1479] , 
        \round_in[3][1478] , \round_in[3][1477] , \round_in[3][1476] , 
        \round_in[3][1475] , \round_in[3][1474] , \round_in[3][1473] , 
        \round_in[3][1472] , \round_in[3][1471] , \round_in[3][1470] , 
        \round_in[3][1469] , \round_in[3][1468] , \round_in[3][1467] , 
        \round_in[3][1466] , \round_in[3][1465] , \round_in[3][1464] , 
        \round_in[3][1463] , \round_in[3][1462] , \round_in[3][1461] , 
        \round_in[3][1460] , \round_in[3][1459] , \round_in[3][1458] , 
        \round_in[3][1457] , \round_in[3][1456] , \round_in[3][1455] , 
        \round_in[3][1454] , \round_in[3][1453] , \round_in[3][1452] , 
        \round_in[3][1451] , \round_in[3][1450] , \round_in[3][1449] , 
        \round_in[3][1448] , \round_in[3][1447] , \round_in[3][1446] , 
        \round_in[3][1445] , \round_in[3][1444] , \round_in[3][1443] , 
        \round_in[3][1442] , \round_in[3][1441] , \round_in[3][1440] , 
        \round_in[3][1439] , \round_in[3][1438] , \round_in[3][1437] , 
        \round_in[3][1436] , \round_in[3][1435] , \round_in[3][1434] , 
        \round_in[3][1433] , \round_in[3][1432] , \round_in[3][1431] , 
        \round_in[3][1430] , \round_in[3][1429] , \round_in[3][1428] , 
        \round_in[3][1427] , \round_in[3][1426] , \round_in[3][1425] , 
        \round_in[3][1424] , \round_in[3][1423] , \round_in[3][1422] , 
        \round_in[3][1421] , \round_in[3][1420] , \round_in[3][1419] , 
        \round_in[3][1418] , \round_in[3][1417] , \round_in[3][1416] , 
        \round_in[3][1415] , \round_in[3][1414] , \round_in[3][1413] , 
        \round_in[3][1412] , \round_in[3][1411] , \round_in[3][1410] , 
        \round_in[3][1409] , \round_in[3][1408] , \round_in[3][1407] , 
        \round_in[3][1406] , \round_in[3][1405] , \round_in[3][1404] , 
        \round_in[3][1403] , \round_in[3][1402] , \round_in[3][1401] , 
        \round_in[3][1400] , \round_in[3][1399] , \round_in[3][1398] , 
        \round_in[3][1397] , \round_in[3][1396] , \round_in[3][1395] , 
        \round_in[3][1394] , \round_in[3][1393] , \round_in[3][1392] , 
        \round_in[3][1391] , \round_in[3][1390] , \round_in[3][1389] , 
        \round_in[3][1388] , \round_in[3][1387] , \round_in[3][1386] , 
        \round_in[3][1385] , \round_in[3][1384] , \round_in[3][1383] , 
        \round_in[3][1382] , \round_in[3][1381] , \round_in[3][1380] , 
        \round_in[3][1379] , \round_in[3][1378] , \round_in[3][1377] , 
        \round_in[3][1376] , \round_in[3][1375] , \round_in[3][1374] , 
        \round_in[3][1373] , \round_in[3][1372] , \round_in[3][1371] , 
        \round_in[3][1370] , \round_in[3][1369] , \round_in[3][1368] , 
        \round_in[3][1367] , \round_in[3][1366] , \round_in[3][1365] , 
        \round_in[3][1364] , \round_in[3][1363] , \round_in[3][1362] , 
        \round_in[3][1361] , \round_in[3][1360] , \round_in[3][1359] , 
        \round_in[3][1358] , \round_in[3][1357] , \round_in[3][1356] , 
        \round_in[3][1355] , \round_in[3][1354] , \round_in[3][1353] , 
        \round_in[3][1352] , \round_in[3][1351] , \round_in[3][1350] , 
        \round_in[3][1349] , \round_in[3][1348] , \round_in[3][1347] , 
        \round_in[3][1346] , \round_in[3][1345] , \round_in[3][1344] , 
        \round_in[3][1343] , \round_in[3][1342] , \round_in[3][1341] , 
        \round_in[3][1340] , \round_in[3][1339] , \round_in[3][1338] , 
        \round_in[3][1337] , \round_in[3][1336] , \round_in[3][1335] , 
        \round_in[3][1334] , \round_in[3][1333] , \round_in[3][1332] , 
        \round_in[3][1331] , \round_in[3][1330] , \round_in[3][1329] , 
        \round_in[3][1328] , \round_in[3][1327] , \round_in[3][1326] , 
        \round_in[3][1325] , \round_in[3][1324] , \round_in[3][1323] , 
        \round_in[3][1322] , \round_in[3][1321] , \round_in[3][1320] , 
        \round_in[3][1319] , \round_in[3][1318] , \round_in[3][1317] , 
        \round_in[3][1316] , \round_in[3][1315] , \round_in[3][1314] , 
        \round_in[3][1313] , \round_in[3][1312] , \round_in[3][1311] , 
        \round_in[3][1310] , \round_in[3][1309] , \round_in[3][1308] , 
        \round_in[3][1307] , \round_in[3][1306] , \round_in[3][1305] , 
        \round_in[3][1304] , \round_in[3][1303] , \round_in[3][1302] , 
        \round_in[3][1301] , \round_in[3][1300] , \round_in[3][1299] , 
        \round_in[3][1298] , \round_in[3][1297] , \round_in[3][1296] , 
        \round_in[3][1295] , \round_in[3][1294] , \round_in[3][1293] , 
        \round_in[3][1292] , \round_in[3][1291] , \round_in[3][1290] , 
        \round_in[3][1289] , \round_in[3][1288] , \round_in[3][1287] , 
        \round_in[3][1286] , \round_in[3][1285] , \round_in[3][1284] , 
        \round_in[3][1283] , \round_in[3][1282] , \round_in[3][1281] , 
        \round_in[3][1280] , \round_in[3][1279] , \round_in[3][1278] , 
        \round_in[3][1277] , \round_in[3][1276] , \round_in[3][1275] , 
        \round_in[3][1274] , \round_in[3][1273] , \round_in[3][1272] , 
        \round_in[3][1271] , \round_in[3][1270] , \round_in[3][1269] , 
        \round_in[3][1268] , \round_in[3][1267] , \round_in[3][1266] , 
        \round_in[3][1265] , \round_in[3][1264] , \round_in[3][1263] , 
        \round_in[3][1262] , \round_in[3][1261] , \round_in[3][1260] , 
        \round_in[3][1259] , \round_in[3][1258] , \round_in[3][1257] , 
        \round_in[3][1256] , \round_in[3][1255] , \round_in[3][1254] , 
        \round_in[3][1253] , \round_in[3][1252] , \round_in[3][1251] , 
        \round_in[3][1250] , \round_in[3][1249] , \round_in[3][1248] , 
        \round_in[3][1247] , \round_in[3][1246] , \round_in[3][1245] , 
        \round_in[3][1244] , \round_in[3][1243] , \round_in[3][1242] , 
        \round_in[3][1241] , \round_in[3][1240] , \round_in[3][1239] , 
        \round_in[3][1238] , \round_in[3][1237] , \round_in[3][1236] , 
        \round_in[3][1235] , \round_in[3][1234] , \round_in[3][1233] , 
        \round_in[3][1232] , \round_in[3][1231] , \round_in[3][1230] , 
        \round_in[3][1229] , \round_in[3][1228] , \round_in[3][1227] , 
        \round_in[3][1226] , \round_in[3][1225] , \round_in[3][1224] , 
        \round_in[3][1223] , \round_in[3][1222] , \round_in[3][1221] , 
        \round_in[3][1220] , \round_in[3][1219] , \round_in[3][1218] , 
        \round_in[3][1217] , \round_in[3][1216] , \round_in[3][1215] , 
        \round_in[3][1214] , \round_in[3][1213] , \round_in[3][1212] , 
        \round_in[3][1211] , \round_in[3][1210] , \round_in[3][1209] , 
        \round_in[3][1208] , \round_in[3][1207] , \round_in[3][1206] , 
        \round_in[3][1205] , \round_in[3][1204] , \round_in[3][1203] , 
        \round_in[3][1202] , \round_in[3][1201] , \round_in[3][1200] , 
        \round_in[3][1199] , \round_in[3][1198] , \round_in[3][1197] , 
        \round_in[3][1196] , \round_in[3][1195] , \round_in[3][1194] , 
        \round_in[3][1193] , \round_in[3][1192] , \round_in[3][1191] , 
        \round_in[3][1190] , \round_in[3][1189] , \round_in[3][1188] , 
        \round_in[3][1187] , \round_in[3][1186] , \round_in[3][1185] , 
        \round_in[3][1184] , \round_in[3][1183] , \round_in[3][1182] , 
        \round_in[3][1181] , \round_in[3][1180] , \round_in[3][1179] , 
        \round_in[3][1178] , \round_in[3][1177] , \round_in[3][1176] , 
        \round_in[3][1175] , \round_in[3][1174] , \round_in[3][1173] , 
        \round_in[3][1172] , \round_in[3][1171] , \round_in[3][1170] , 
        \round_in[3][1169] , \round_in[3][1168] , \round_in[3][1167] , 
        \round_in[3][1166] , \round_in[3][1165] , \round_in[3][1164] , 
        \round_in[3][1163] , \round_in[3][1162] , \round_in[3][1161] , 
        \round_in[3][1160] , \round_in[3][1159] , \round_in[3][1158] , 
        \round_in[3][1157] , \round_in[3][1156] , \round_in[3][1155] , 
        \round_in[3][1154] , \round_in[3][1153] , \round_in[3][1152] , 
        \round_in[3][1151] , \round_in[3][1150] , \round_in[3][1149] , 
        \round_in[3][1148] , \round_in[3][1147] , \round_in[3][1146] , 
        \round_in[3][1145] , \round_in[3][1144] , \round_in[3][1143] , 
        \round_in[3][1142] , \round_in[3][1141] , \round_in[3][1140] , 
        \round_in[3][1139] , \round_in[3][1138] , \round_in[3][1137] , 
        \round_in[3][1136] , \round_in[3][1135] , \round_in[3][1134] , 
        \round_in[3][1133] , \round_in[3][1132] , \round_in[3][1131] , 
        \round_in[3][1130] , \round_in[3][1129] , \round_in[3][1128] , 
        \round_in[3][1127] , \round_in[3][1126] , \round_in[3][1125] , 
        \round_in[3][1124] , \round_in[3][1123] , \round_in[3][1122] , 
        \round_in[3][1121] , \round_in[3][1120] , \round_in[3][1119] , 
        \round_in[3][1118] , \round_in[3][1117] , \round_in[3][1116] , 
        \round_in[3][1115] , \round_in[3][1114] , \round_in[3][1113] , 
        \round_in[3][1112] , \round_in[3][1111] , \round_in[3][1110] , 
        \round_in[3][1109] , \round_in[3][1108] , \round_in[3][1107] , 
        \round_in[3][1106] , \round_in[3][1105] , \round_in[3][1104] , 
        \round_in[3][1103] , \round_in[3][1102] , \round_in[3][1101] , 
        \round_in[3][1100] , \round_in[3][1099] , \round_in[3][1098] , 
        \round_in[3][1097] , \round_in[3][1096] , \round_in[3][1095] , 
        \round_in[3][1094] , \round_in[3][1093] , \round_in[3][1092] , 
        \round_in[3][1091] , \round_in[3][1090] , \round_in[3][1089] , 
        \round_in[3][1088] , \round_in[3][1087] , \round_in[3][1086] , 
        \round_in[3][1085] , \round_in[3][1084] , \round_in[3][1083] , 
        \round_in[3][1082] , \round_in[3][1081] , \round_in[3][1080] , 
        \round_in[3][1079] , \round_in[3][1078] , \round_in[3][1077] , 
        \round_in[3][1076] , \round_in[3][1075] , \round_in[3][1074] , 
        \round_in[3][1073] , \round_in[3][1072] , \round_in[3][1071] , 
        \round_in[3][1070] , \round_in[3][1069] , \round_in[3][1068] , 
        \round_in[3][1067] , \round_in[3][1066] , \round_in[3][1065] , 
        \round_in[3][1064] , \round_in[3][1063] , \round_in[3][1062] , 
        \round_in[3][1061] , \round_in[3][1060] , \round_in[3][1059] , 
        \round_in[3][1058] , \round_in[3][1057] , \round_in[3][1056] , 
        \round_in[3][1055] , \round_in[3][1054] , \round_in[3][1053] , 
        \round_in[3][1052] , \round_in[3][1051] , \round_in[3][1050] , 
        \round_in[3][1049] , \round_in[3][1048] , \round_in[3][1047] , 
        \round_in[3][1046] , \round_in[3][1045] , \round_in[3][1044] , 
        \round_in[3][1043] , \round_in[3][1042] , \round_in[3][1041] , 
        \round_in[3][1040] , \round_in[3][1039] , \round_in[3][1038] , 
        \round_in[3][1037] , \round_in[3][1036] , \round_in[3][1035] , 
        \round_in[3][1034] , \round_in[3][1033] , \round_in[3][1032] , 
        \round_in[3][1031] , \round_in[3][1030] , \round_in[3][1029] , 
        \round_in[3][1028] , \round_in[3][1027] , \round_in[3][1026] , 
        \round_in[3][1025] , \round_in[3][1024] , \round_in[3][1023] , 
        \round_in[3][1022] , \round_in[3][1021] , \round_in[3][1020] , 
        \round_in[3][1019] , \round_in[3][1018] , \round_in[3][1017] , 
        \round_in[3][1016] , \round_in[3][1015] , \round_in[3][1014] , 
        \round_in[3][1013] , \round_in[3][1012] , \round_in[3][1011] , 
        \round_in[3][1010] , \round_in[3][1009] , \round_in[3][1008] , 
        \round_in[3][1007] , \round_in[3][1006] , \round_in[3][1005] , 
        \round_in[3][1004] , \round_in[3][1003] , \round_in[3][1002] , 
        \round_in[3][1001] , \round_in[3][1000] , \round_in[3][999] , 
        \round_in[3][998] , \round_in[3][997] , \round_in[3][996] , 
        \round_in[3][995] , \round_in[3][994] , \round_in[3][993] , 
        \round_in[3][992] , \round_in[3][991] , \round_in[3][990] , 
        \round_in[3][989] , \round_in[3][988] , \round_in[3][987] , 
        \round_in[3][986] , \round_in[3][985] , \round_in[3][984] , 
        \round_in[3][983] , \round_in[3][982] , \round_in[3][981] , 
        \round_in[3][980] , \round_in[3][979] , \round_in[3][978] , 
        \round_in[3][977] , \round_in[3][976] , \round_in[3][975] , 
        \round_in[3][974] , \round_in[3][973] , \round_in[3][972] , 
        \round_in[3][971] , \round_in[3][970] , \round_in[3][969] , 
        \round_in[3][968] , \round_in[3][967] , \round_in[3][966] , 
        \round_in[3][965] , \round_in[3][964] , \round_in[3][963] , 
        \round_in[3][962] , \round_in[3][961] , \round_in[3][960] , 
        \round_in[3][959] , \round_in[3][958] , \round_in[3][957] , 
        \round_in[3][956] , \round_in[3][955] , \round_in[3][954] , 
        \round_in[3][953] , \round_in[3][952] , \round_in[3][951] , 
        \round_in[3][950] , \round_in[3][949] , \round_in[3][948] , 
        \round_in[3][947] , \round_in[3][946] , \round_in[3][945] , 
        \round_in[3][944] , \round_in[3][943] , \round_in[3][942] , 
        \round_in[3][941] , \round_in[3][940] , \round_in[3][939] , 
        \round_in[3][938] , \round_in[3][937] , \round_in[3][936] , 
        \round_in[3][935] , \round_in[3][934] , \round_in[3][933] , 
        \round_in[3][932] , \round_in[3][931] , \round_in[3][930] , 
        \round_in[3][929] , \round_in[3][928] , \round_in[3][927] , 
        \round_in[3][926] , \round_in[3][925] , \round_in[3][924] , 
        \round_in[3][923] , \round_in[3][922] , \round_in[3][921] , 
        \round_in[3][920] , \round_in[3][919] , \round_in[3][918] , 
        \round_in[3][917] , \round_in[3][916] , \round_in[3][915] , 
        \round_in[3][914] , \round_in[3][913] , \round_in[3][912] , 
        \round_in[3][911] , \round_in[3][910] , \round_in[3][909] , 
        \round_in[3][908] , \round_in[3][907] , \round_in[3][906] , 
        \round_in[3][905] , \round_in[3][904] , \round_in[3][903] , 
        \round_in[3][902] , \round_in[3][901] , \round_in[3][900] , 
        \round_in[3][899] , \round_in[3][898] , \round_in[3][897] , 
        \round_in[3][896] , \round_in[3][895] , \round_in[3][894] , 
        \round_in[3][893] , \round_in[3][892] , \round_in[3][891] , 
        \round_in[3][890] , \round_in[3][889] , \round_in[3][888] , 
        \round_in[3][887] , \round_in[3][886] , \round_in[3][885] , 
        \round_in[3][884] , \round_in[3][883] , \round_in[3][882] , 
        \round_in[3][881] , \round_in[3][880] , \round_in[3][879] , 
        \round_in[3][878] , \round_in[3][877] , \round_in[3][876] , 
        \round_in[3][875] , \round_in[3][874] , \round_in[3][873] , 
        \round_in[3][872] , \round_in[3][871] , \round_in[3][870] , 
        \round_in[3][869] , \round_in[3][868] , \round_in[3][867] , 
        \round_in[3][866] , \round_in[3][865] , \round_in[3][864] , 
        \round_in[3][863] , \round_in[3][862] , \round_in[3][861] , 
        \round_in[3][860] , \round_in[3][859] , \round_in[3][858] , 
        \round_in[3][857] , \round_in[3][856] , \round_in[3][855] , 
        \round_in[3][854] , \round_in[3][853] , \round_in[3][852] , 
        \round_in[3][851] , \round_in[3][850] , \round_in[3][849] , 
        \round_in[3][848] , \round_in[3][847] , \round_in[3][846] , 
        \round_in[3][845] , \round_in[3][844] , \round_in[3][843] , 
        \round_in[3][842] , \round_in[3][841] , \round_in[3][840] , 
        \round_in[3][839] , \round_in[3][838] , \round_in[3][837] , 
        \round_in[3][836] , \round_in[3][835] , \round_in[3][834] , 
        \round_in[3][833] , \round_in[3][832] , \round_in[3][831] , 
        \round_in[3][830] , \round_in[3][829] , \round_in[3][828] , 
        \round_in[3][827] , \round_in[3][826] , \round_in[3][825] , 
        \round_in[3][824] , \round_in[3][823] , \round_in[3][822] , 
        \round_in[3][821] , \round_in[3][820] , \round_in[3][819] , 
        \round_in[3][818] , \round_in[3][817] , \round_in[3][816] , 
        \round_in[3][815] , \round_in[3][814] , \round_in[3][813] , 
        \round_in[3][812] , \round_in[3][811] , \round_in[3][810] , 
        \round_in[3][809] , \round_in[3][808] , \round_in[3][807] , 
        \round_in[3][806] , \round_in[3][805] , \round_in[3][804] , 
        \round_in[3][803] , \round_in[3][802] , \round_in[3][801] , 
        \round_in[3][800] , \round_in[3][799] , \round_in[3][798] , 
        \round_in[3][797] , \round_in[3][796] , \round_in[3][795] , 
        \round_in[3][794] , \round_in[3][793] , \round_in[3][792] , 
        \round_in[3][791] , \round_in[3][790] , \round_in[3][789] , 
        \round_in[3][788] , \round_in[3][787] , \round_in[3][786] , 
        \round_in[3][785] , \round_in[3][784] , \round_in[3][783] , 
        \round_in[3][782] , \round_in[3][781] , \round_in[3][780] , 
        \round_in[3][779] , \round_in[3][778] , \round_in[3][777] , 
        \round_in[3][776] , \round_in[3][775] , \round_in[3][774] , 
        \round_in[3][773] , \round_in[3][772] , \round_in[3][771] , 
        \round_in[3][770] , \round_in[3][769] , \round_in[3][768] , 
        \round_in[3][767] , \round_in[3][766] , \round_in[3][765] , 
        \round_in[3][764] , \round_in[3][763] , \round_in[3][762] , 
        \round_in[3][761] , \round_in[3][760] , \round_in[3][759] , 
        \round_in[3][758] , \round_in[3][757] , \round_in[3][756] , 
        \round_in[3][755] , \round_in[3][754] , \round_in[3][753] , 
        \round_in[3][752] , \round_in[3][751] , \round_in[3][750] , 
        \round_in[3][749] , \round_in[3][748] , \round_in[3][747] , 
        \round_in[3][746] , \round_in[3][745] , \round_in[3][744] , 
        \round_in[3][743] , \round_in[3][742] , \round_in[3][741] , 
        \round_in[3][740] , \round_in[3][739] , \round_in[3][738] , 
        \round_in[3][737] , \round_in[3][736] , \round_in[3][735] , 
        \round_in[3][734] , \round_in[3][733] , \round_in[3][732] , 
        \round_in[3][731] , \round_in[3][730] , \round_in[3][729] , 
        \round_in[3][728] , \round_in[3][727] , \round_in[3][726] , 
        \round_in[3][725] , \round_in[3][724] , \round_in[3][723] , 
        \round_in[3][722] , \round_in[3][721] , \round_in[3][720] , 
        \round_in[3][719] , \round_in[3][718] , \round_in[3][717] , 
        \round_in[3][716] , \round_in[3][715] , \round_in[3][714] , 
        \round_in[3][713] , \round_in[3][712] , \round_in[3][711] , 
        \round_in[3][710] , \round_in[3][709] , \round_in[3][708] , 
        \round_in[3][707] , \round_in[3][706] , \round_in[3][705] , 
        \round_in[3][704] , \round_in[3][703] , \round_in[3][702] , 
        \round_in[3][701] , \round_in[3][700] , \round_in[3][699] , 
        \round_in[3][698] , \round_in[3][697] , \round_in[3][696] , 
        \round_in[3][695] , \round_in[3][694] , \round_in[3][693] , 
        \round_in[3][692] , \round_in[3][691] , \round_in[3][690] , 
        \round_in[3][689] , \round_in[3][688] , \round_in[3][687] , 
        \round_in[3][686] , \round_in[3][685] , \round_in[3][684] , 
        \round_in[3][683] , \round_in[3][682] , \round_in[3][681] , 
        \round_in[3][680] , \round_in[3][679] , \round_in[3][678] , 
        \round_in[3][677] , \round_in[3][676] , \round_in[3][675] , 
        \round_in[3][674] , \round_in[3][673] , \round_in[3][672] , 
        \round_in[3][671] , \round_in[3][670] , \round_in[3][669] , 
        \round_in[3][668] , \round_in[3][667] , \round_in[3][666] , 
        \round_in[3][665] , \round_in[3][664] , \round_in[3][663] , 
        \round_in[3][662] , \round_in[3][661] , \round_in[3][660] , 
        \round_in[3][659] , \round_in[3][658] , \round_in[3][657] , 
        \round_in[3][656] , \round_in[3][655] , \round_in[3][654] , 
        \round_in[3][653] , \round_in[3][652] , \round_in[3][651] , 
        \round_in[3][650] , \round_in[3][649] , \round_in[3][648] , 
        \round_in[3][647] , \round_in[3][646] , \round_in[3][645] , 
        \round_in[3][644] , \round_in[3][643] , \round_in[3][642] , 
        \round_in[3][641] , \round_in[3][640] , \round_in[3][639] , 
        \round_in[3][638] , \round_in[3][637] , \round_in[3][636] , 
        \round_in[3][635] , \round_in[3][634] , \round_in[3][633] , 
        \round_in[3][632] , \round_in[3][631] , \round_in[3][630] , 
        \round_in[3][629] , \round_in[3][628] , \round_in[3][627] , 
        \round_in[3][626] , \round_in[3][625] , \round_in[3][624] , 
        \round_in[3][623] , \round_in[3][622] , \round_in[3][621] , 
        \round_in[3][620] , \round_in[3][619] , \round_in[3][618] , 
        \round_in[3][617] , \round_in[3][616] , \round_in[3][615] , 
        \round_in[3][614] , \round_in[3][613] , \round_in[3][612] , 
        \round_in[3][611] , \round_in[3][610] , \round_in[3][609] , 
        \round_in[3][608] , \round_in[3][607] , \round_in[3][606] , 
        \round_in[3][605] , \round_in[3][604] , \round_in[3][603] , 
        \round_in[3][602] , \round_in[3][601] , \round_in[3][600] , 
        \round_in[3][599] , \round_in[3][598] , \round_in[3][597] , 
        \round_in[3][596] , \round_in[3][595] , \round_in[3][594] , 
        \round_in[3][593] , \round_in[3][592] , \round_in[3][591] , 
        \round_in[3][590] , \round_in[3][589] , \round_in[3][588] , 
        \round_in[3][587] , \round_in[3][586] , \round_in[3][585] , 
        \round_in[3][584] , \round_in[3][583] , \round_in[3][582] , 
        \round_in[3][581] , \round_in[3][580] , \round_in[3][579] , 
        \round_in[3][578] , \round_in[3][577] , \round_in[3][576] , 
        \round_in[3][575] , \round_in[3][574] , \round_in[3][573] , 
        \round_in[3][572] , \round_in[3][571] , \round_in[3][570] , 
        \round_in[3][569] , \round_in[3][568] , \round_in[3][567] , 
        \round_in[3][566] , \round_in[3][565] , \round_in[3][564] , 
        \round_in[3][563] , \round_in[3][562] , \round_in[3][561] , 
        \round_in[3][560] , \round_in[3][559] , \round_in[3][558] , 
        \round_in[3][557] , \round_in[3][556] , \round_in[3][555] , 
        \round_in[3][554] , \round_in[3][553] , \round_in[3][552] , 
        \round_in[3][551] , \round_in[3][550] , \round_in[3][549] , 
        \round_in[3][548] , \round_in[3][547] , \round_in[3][546] , 
        \round_in[3][545] , \round_in[3][544] , \round_in[3][543] , 
        \round_in[3][542] , \round_in[3][541] , \round_in[3][540] , 
        \round_in[3][539] , \round_in[3][538] , \round_in[3][537] , 
        \round_in[3][536] , \round_in[3][535] , \round_in[3][534] , 
        \round_in[3][533] , \round_in[3][532] , \round_in[3][531] , 
        \round_in[3][530] , \round_in[3][529] , \round_in[3][528] , 
        \round_in[3][527] , \round_in[3][526] , \round_in[3][525] , 
        \round_in[3][524] , \round_in[3][523] , \round_in[3][522] , 
        \round_in[3][521] , \round_in[3][520] , \round_in[3][519] , 
        \round_in[3][518] , \round_in[3][517] , \round_in[3][516] , 
        \round_in[3][515] , \round_in[3][514] , \round_in[3][513] , 
        \round_in[3][512] , \round_in[3][511] , \round_in[3][510] , 
        \round_in[3][509] , \round_in[3][508] , \round_in[3][507] , 
        \round_in[3][506] , \round_in[3][505] , \round_in[3][504] , 
        \round_in[3][503] , \round_in[3][502] , \round_in[3][501] , 
        \round_in[3][500] , \round_in[3][499] , \round_in[3][498] , 
        \round_in[3][497] , \round_in[3][496] , \round_in[3][495] , 
        \round_in[3][494] , \round_in[3][493] , \round_in[3][492] , 
        \round_in[3][491] , \round_in[3][490] , \round_in[3][489] , 
        \round_in[3][488] , \round_in[3][487] , \round_in[3][486] , 
        \round_in[3][485] , \round_in[3][484] , \round_in[3][483] , 
        \round_in[3][482] , \round_in[3][481] , \round_in[3][480] , 
        \round_in[3][479] , \round_in[3][478] , \round_in[3][477] , 
        \round_in[3][476] , \round_in[3][475] , \round_in[3][474] , 
        \round_in[3][473] , \round_in[3][472] , \round_in[3][471] , 
        \round_in[3][470] , \round_in[3][469] , \round_in[3][468] , 
        \round_in[3][467] , \round_in[3][466] , \round_in[3][465] , 
        \round_in[3][464] , \round_in[3][463] , \round_in[3][462] , 
        \round_in[3][461] , \round_in[3][460] , \round_in[3][459] , 
        \round_in[3][458] , \round_in[3][457] , \round_in[3][456] , 
        \round_in[3][455] , \round_in[3][454] , \round_in[3][453] , 
        \round_in[3][452] , \round_in[3][451] , \round_in[3][450] , 
        \round_in[3][449] , \round_in[3][448] , \round_in[3][447] , 
        \round_in[3][446] , \round_in[3][445] , \round_in[3][444] , 
        \round_in[3][443] , \round_in[3][442] , \round_in[3][441] , 
        \round_in[3][440] , \round_in[3][439] , \round_in[3][438] , 
        \round_in[3][437] , \round_in[3][436] , \round_in[3][435] , 
        \round_in[3][434] , \round_in[3][433] , \round_in[3][432] , 
        \round_in[3][431] , \round_in[3][430] , \round_in[3][429] , 
        \round_in[3][428] , \round_in[3][427] , \round_in[3][426] , 
        \round_in[3][425] , \round_in[3][424] , \round_in[3][423] , 
        \round_in[3][422] , \round_in[3][421] , \round_in[3][420] , 
        \round_in[3][419] , \round_in[3][418] , \round_in[3][417] , 
        \round_in[3][416] , \round_in[3][415] , \round_in[3][414] , 
        \round_in[3][413] , \round_in[3][412] , \round_in[3][411] , 
        \round_in[3][410] , \round_in[3][409] , \round_in[3][408] , 
        \round_in[3][407] , \round_in[3][406] , \round_in[3][405] , 
        \round_in[3][404] , \round_in[3][403] , \round_in[3][402] , 
        \round_in[3][401] , \round_in[3][400] , \round_in[3][399] , 
        \round_in[3][398] , \round_in[3][397] , \round_in[3][396] , 
        \round_in[3][395] , \round_in[3][394] , \round_in[3][393] , 
        \round_in[3][392] , \round_in[3][391] , \round_in[3][390] , 
        \round_in[3][389] , \round_in[3][388] , \round_in[3][387] , 
        \round_in[3][386] , \round_in[3][385] , \round_in[3][384] , 
        \round_in[3][383] , \round_in[3][382] , \round_in[3][381] , 
        \round_in[3][380] , \round_in[3][379] , \round_in[3][378] , 
        \round_in[3][377] , \round_in[3][376] , \round_in[3][375] , 
        \round_in[3][374] , \round_in[3][373] , \round_in[3][372] , 
        \round_in[3][371] , \round_in[3][370] , \round_in[3][369] , 
        \round_in[3][368] , \round_in[3][367] , \round_in[3][366] , 
        \round_in[3][365] , \round_in[3][364] , \round_in[3][363] , 
        \round_in[3][362] , \round_in[3][361] , \round_in[3][360] , 
        \round_in[3][359] , \round_in[3][358] , \round_in[3][357] , 
        \round_in[3][356] , \round_in[3][355] , \round_in[3][354] , 
        \round_in[3][353] , \round_in[3][352] , \round_in[3][351] , 
        \round_in[3][350] , \round_in[3][349] , \round_in[3][348] , 
        \round_in[3][347] , \round_in[3][346] , \round_in[3][345] , 
        \round_in[3][344] , \round_in[3][343] , \round_in[3][342] , 
        \round_in[3][341] , \round_in[3][340] , \round_in[3][339] , 
        \round_in[3][338] , \round_in[3][337] , \round_in[3][336] , 
        \round_in[3][335] , \round_in[3][334] , \round_in[3][333] , 
        \round_in[3][332] , \round_in[3][331] , \round_in[3][330] , 
        \round_in[3][329] , \round_in[3][328] , \round_in[3][327] , 
        \round_in[3][326] , \round_in[3][325] , \round_in[3][324] , 
        \round_in[3][323] , \round_in[3][322] , \round_in[3][321] , 
        \round_in[3][320] , \round_in[3][319] , \round_in[3][318] , 
        \round_in[3][317] , \round_in[3][316] , \round_in[3][315] , 
        \round_in[3][314] , \round_in[3][313] , \round_in[3][312] , 
        \round_in[3][311] , \round_in[3][310] , \round_in[3][309] , 
        \round_in[3][308] , \round_in[3][307] , \round_in[3][306] , 
        \round_in[3][305] , \round_in[3][304] , \round_in[3][303] , 
        \round_in[3][302] , \round_in[3][301] , \round_in[3][300] , 
        \round_in[3][299] , \round_in[3][298] , \round_in[3][297] , 
        \round_in[3][296] , \round_in[3][295] , \round_in[3][294] , 
        \round_in[3][293] , \round_in[3][292] , \round_in[3][291] , 
        \round_in[3][290] , \round_in[3][289] , \round_in[3][288] , 
        \round_in[3][287] , \round_in[3][286] , \round_in[3][285] , 
        \round_in[3][284] , \round_in[3][283] , \round_in[3][282] , 
        \round_in[3][281] , \round_in[3][280] , \round_in[3][279] , 
        \round_in[3][278] , \round_in[3][277] , \round_in[3][276] , 
        \round_in[3][275] , \round_in[3][274] , \round_in[3][273] , 
        \round_in[3][272] , \round_in[3][271] , \round_in[3][270] , 
        \round_in[3][269] , \round_in[3][268] , \round_in[3][267] , 
        \round_in[3][266] , \round_in[3][265] , \round_in[3][264] , 
        \round_in[3][263] , \round_in[3][262] , \round_in[3][261] , 
        \round_in[3][260] , \round_in[3][259] , \round_in[3][258] , 
        \round_in[3][257] , \round_in[3][256] , \round_in[3][255] , 
        \round_in[3][254] , \round_in[3][253] , \round_in[3][252] , 
        \round_in[3][251] , \round_in[3][250] , \round_in[3][249] , 
        \round_in[3][248] , \round_in[3][247] , \round_in[3][246] , 
        \round_in[3][245] , \round_in[3][244] , \round_in[3][243] , 
        \round_in[3][242] , \round_in[3][241] , \round_in[3][240] , 
        \round_in[3][239] , \round_in[3][238] , \round_in[3][237] , 
        \round_in[3][236] , \round_in[3][235] , \round_in[3][234] , 
        \round_in[3][233] , \round_in[3][232] , \round_in[3][231] , 
        \round_in[3][230] , \round_in[3][229] , \round_in[3][228] , 
        \round_in[3][227] , \round_in[3][226] , \round_in[3][225] , 
        \round_in[3][224] , \round_in[3][223] , \round_in[3][222] , 
        \round_in[3][221] , \round_in[3][220] , \round_in[3][219] , 
        \round_in[3][218] , \round_in[3][217] , \round_in[3][216] , 
        \round_in[3][215] , \round_in[3][214] , \round_in[3][213] , 
        \round_in[3][212] , \round_in[3][211] , \round_in[3][210] , 
        \round_in[3][209] , \round_in[3][208] , \round_in[3][207] , 
        \round_in[3][206] , \round_in[3][205] , \round_in[3][204] , 
        \round_in[3][203] , \round_in[3][202] , \round_in[3][201] , 
        \round_in[3][200] , \round_in[3][199] , \round_in[3][198] , 
        \round_in[3][197] , \round_in[3][196] , \round_in[3][195] , 
        \round_in[3][194] , \round_in[3][193] , \round_in[3][192] , 
        \round_in[3][191] , \round_in[3][190] , \round_in[3][189] , 
        \round_in[3][188] , \round_in[3][187] , \round_in[3][186] , 
        \round_in[3][185] , \round_in[3][184] , \round_in[3][183] , 
        \round_in[3][182] , \round_in[3][181] , \round_in[3][180] , 
        \round_in[3][179] , \round_in[3][178] , \round_in[3][177] , 
        \round_in[3][176] , \round_in[3][175] , \round_in[3][174] , 
        \round_in[3][173] , \round_in[3][172] , \round_in[3][171] , 
        \round_in[3][170] , \round_in[3][169] , \round_in[3][168] , 
        \round_in[3][167] , \round_in[3][166] , \round_in[3][165] , 
        \round_in[3][164] , \round_in[3][163] , \round_in[3][162] , 
        \round_in[3][161] , \round_in[3][160] , \round_in[3][159] , 
        \round_in[3][158] , \round_in[3][157] , \round_in[3][156] , 
        \round_in[3][155] , \round_in[3][154] , \round_in[3][153] , 
        \round_in[3][152] , \round_in[3][151] , \round_in[3][150] , 
        \round_in[3][149] , \round_in[3][148] , \round_in[3][147] , 
        \round_in[3][146] , \round_in[3][145] , \round_in[3][144] , 
        \round_in[3][143] , \round_in[3][142] , \round_in[3][141] , 
        \round_in[3][140] , \round_in[3][139] , \round_in[3][138] , 
        \round_in[3][137] , \round_in[3][136] , \round_in[3][135] , 
        \round_in[3][134] , \round_in[3][133] , \round_in[3][132] , 
        \round_in[3][131] , \round_in[3][130] , \round_in[3][129] , 
        \round_in[3][128] , \round_in[3][127] , \round_in[3][126] , 
        \round_in[3][125] , \round_in[3][124] , \round_in[3][123] , 
        \round_in[3][122] , \round_in[3][121] , \round_in[3][120] , 
        \round_in[3][119] , \round_in[3][118] , \round_in[3][117] , 
        \round_in[3][116] , \round_in[3][115] , \round_in[3][114] , 
        \round_in[3][113] , \round_in[3][112] , \round_in[3][111] , 
        \round_in[3][110] , \round_in[3][109] , \round_in[3][108] , 
        \round_in[3][107] , \round_in[3][106] , \round_in[3][105] , 
        \round_in[3][104] , \round_in[3][103] , \round_in[3][102] , 
        \round_in[3][101] , \round_in[3][100] , \round_in[3][99] , 
        \round_in[3][98] , \round_in[3][97] , \round_in[3][96] , 
        \round_in[3][95] , \round_in[3][94] , \round_in[3][93] , 
        \round_in[3][92] , \round_in[3][91] , \round_in[3][90] , 
        \round_in[3][89] , \round_in[3][88] , \round_in[3][87] , 
        \round_in[3][86] , \round_in[3][85] , \round_in[3][84] , 
        \round_in[3][83] , \round_in[3][82] , \round_in[3][81] , 
        \round_in[3][80] , \round_in[3][79] , \round_in[3][78] , 
        \round_in[3][77] , \round_in[3][76] , \round_in[3][75] , 
        \round_in[3][74] , \round_in[3][73] , \round_in[3][72] , 
        \round_in[3][71] , \round_in[3][70] , \round_in[3][69] , 
        \round_in[3][68] , \round_in[3][67] , \round_in[3][66] , 
        \round_in[3][65] , \round_in[3][64] , \round_in[3][63] , 
        \round_in[3][62] , \round_in[3][61] , \round_in[3][60] , 
        \round_in[3][59] , \round_in[3][58] , \round_in[3][57] , 
        \round_in[3][56] , \round_in[3][55] , \round_in[3][54] , 
        \round_in[3][53] , \round_in[3][52] , \round_in[3][51] , 
        \round_in[3][50] , \round_in[3][49] , \round_in[3][48] , 
        \round_in[3][47] , \round_in[3][46] , \round_in[3][45] , 
        \round_in[3][44] , \round_in[3][43] , \round_in[3][42] , 
        \round_in[3][41] , \round_in[3][40] , \round_in[3][39] , 
        \round_in[3][38] , \round_in[3][37] , \round_in[3][36] , 
        \round_in[3][35] , \round_in[3][34] , \round_in[3][33] , 
        \round_in[3][32] , \round_in[3][31] , \round_in[3][30] , 
        \round_in[3][29] , \round_in[3][28] , \round_in[3][27] , 
        \round_in[3][26] , \round_in[3][25] , \round_in[3][24] , 
        \round_in[3][23] , \round_in[3][22] , \round_in[3][21] , 
        \round_in[3][20] , \round_in[3][19] , \round_in[3][18] , 
        \round_in[3][17] , \round_in[3][16] , \round_in[3][15] , 
        \round_in[3][14] , \round_in[3][13] , \round_in[3][12] , 
        \round_in[3][11] , \round_in[3][10] , \round_in[3][9] , 
        \round_in[3][8] , \round_in[3][7] , \round_in[3][6] , \round_in[3][5] , 
        \round_in[3][4] , \round_in[3][3] , \round_in[3][2] , \round_in[3][1] , 
        \round_in[3][0] }) );
  round_3 \ROUND[3].round_  ( .in({\round_in[3][1599] , \round_in[3][1598] , 
        \round_in[3][1597] , \round_in[3][1596] , \round_in[3][1595] , 
        \round_in[3][1594] , \round_in[3][1593] , \round_in[3][1592] , 
        \round_in[3][1591] , \round_in[3][1590] , \round_in[3][1589] , 
        \round_in[3][1588] , \round_in[3][1587] , \round_in[3][1586] , 
        \round_in[3][1585] , \round_in[3][1584] , \round_in[3][1583] , 
        \round_in[3][1582] , \round_in[3][1581] , \round_in[3][1580] , 
        \round_in[3][1579] , \round_in[3][1578] , \round_in[3][1577] , 
        \round_in[3][1576] , \round_in[3][1575] , \round_in[3][1574] , 
        \round_in[3][1573] , \round_in[3][1572] , \round_in[3][1571] , 
        \round_in[3][1570] , \round_in[3][1569] , \round_in[3][1568] , 
        \round_in[3][1567] , \round_in[3][1566] , \round_in[3][1565] , 
        \round_in[3][1564] , \round_in[3][1563] , \round_in[3][1562] , 
        \round_in[3][1561] , \round_in[3][1560] , \round_in[3][1559] , 
        \round_in[3][1558] , \round_in[3][1557] , \round_in[3][1556] , 
        \round_in[3][1555] , \round_in[3][1554] , \round_in[3][1553] , 
        \round_in[3][1552] , \round_in[3][1551] , \round_in[3][1550] , 
        \round_in[3][1549] , \round_in[3][1548] , \round_in[3][1547] , 
        \round_in[3][1546] , \round_in[3][1545] , \round_in[3][1544] , 
        \round_in[3][1543] , \round_in[3][1542] , \round_in[3][1541] , 
        \round_in[3][1540] , \round_in[3][1539] , \round_in[3][1538] , 
        \round_in[3][1537] , \round_in[3][1536] , \round_in[3][1535] , 
        \round_in[3][1534] , \round_in[3][1533] , \round_in[3][1532] , 
        \round_in[3][1531] , \round_in[3][1530] , \round_in[3][1529] , 
        \round_in[3][1528] , \round_in[3][1527] , \round_in[3][1526] , 
        \round_in[3][1525] , \round_in[3][1524] , \round_in[3][1523] , 
        \round_in[3][1522] , \round_in[3][1521] , \round_in[3][1520] , 
        \round_in[3][1519] , \round_in[3][1518] , \round_in[3][1517] , 
        \round_in[3][1516] , \round_in[3][1515] , \round_in[3][1514] , 
        \round_in[3][1513] , \round_in[3][1512] , \round_in[3][1511] , 
        \round_in[3][1510] , \round_in[3][1509] , \round_in[3][1508] , 
        \round_in[3][1507] , \round_in[3][1506] , \round_in[3][1505] , 
        \round_in[3][1504] , \round_in[3][1503] , \round_in[3][1502] , 
        \round_in[3][1501] , \round_in[3][1500] , \round_in[3][1499] , 
        \round_in[3][1498] , \round_in[3][1497] , \round_in[3][1496] , 
        \round_in[3][1495] , \round_in[3][1494] , \round_in[3][1493] , 
        \round_in[3][1492] , \round_in[3][1491] , \round_in[3][1490] , 
        \round_in[3][1489] , \round_in[3][1488] , \round_in[3][1487] , 
        \round_in[3][1486] , \round_in[3][1485] , \round_in[3][1484] , 
        \round_in[3][1483] , \round_in[3][1482] , \round_in[3][1481] , 
        \round_in[3][1480] , \round_in[3][1479] , \round_in[3][1478] , 
        \round_in[3][1477] , \round_in[3][1476] , \round_in[3][1475] , 
        \round_in[3][1474] , \round_in[3][1473] , \round_in[3][1472] , 
        \round_in[3][1471] , \round_in[3][1470] , \round_in[3][1469] , 
        \round_in[3][1468] , \round_in[3][1467] , \round_in[3][1466] , 
        \round_in[3][1465] , \round_in[3][1464] , \round_in[3][1463] , 
        \round_in[3][1462] , \round_in[3][1461] , \round_in[3][1460] , 
        \round_in[3][1459] , \round_in[3][1458] , \round_in[3][1457] , 
        \round_in[3][1456] , \round_in[3][1455] , \round_in[3][1454] , 
        \round_in[3][1453] , \round_in[3][1452] , \round_in[3][1451] , 
        \round_in[3][1450] , \round_in[3][1449] , \round_in[3][1448] , 
        \round_in[3][1447] , \round_in[3][1446] , \round_in[3][1445] , 
        \round_in[3][1444] , \round_in[3][1443] , \round_in[3][1442] , 
        \round_in[3][1441] , \round_in[3][1440] , \round_in[3][1439] , 
        \round_in[3][1438] , \round_in[3][1437] , \round_in[3][1436] , 
        \round_in[3][1435] , \round_in[3][1434] , \round_in[3][1433] , 
        \round_in[3][1432] , \round_in[3][1431] , \round_in[3][1430] , 
        \round_in[3][1429] , \round_in[3][1428] , \round_in[3][1427] , 
        \round_in[3][1426] , \round_in[3][1425] , \round_in[3][1424] , 
        \round_in[3][1423] , \round_in[3][1422] , \round_in[3][1421] , 
        \round_in[3][1420] , \round_in[3][1419] , \round_in[3][1418] , 
        \round_in[3][1417] , \round_in[3][1416] , \round_in[3][1415] , 
        \round_in[3][1414] , \round_in[3][1413] , \round_in[3][1412] , 
        \round_in[3][1411] , \round_in[3][1410] , \round_in[3][1409] , 
        \round_in[3][1408] , \round_in[3][1407] , \round_in[3][1406] , 
        \round_in[3][1405] , \round_in[3][1404] , \round_in[3][1403] , 
        \round_in[3][1402] , \round_in[3][1401] , \round_in[3][1400] , 
        \round_in[3][1399] , \round_in[3][1398] , \round_in[3][1397] , 
        \round_in[3][1396] , \round_in[3][1395] , \round_in[3][1394] , 
        \round_in[3][1393] , \round_in[3][1392] , \round_in[3][1391] , 
        \round_in[3][1390] , \round_in[3][1389] , \round_in[3][1388] , 
        \round_in[3][1387] , \round_in[3][1386] , \round_in[3][1385] , 
        \round_in[3][1384] , \round_in[3][1383] , \round_in[3][1382] , 
        \round_in[3][1381] , \round_in[3][1380] , \round_in[3][1379] , 
        \round_in[3][1378] , \round_in[3][1377] , \round_in[3][1376] , 
        \round_in[3][1375] , \round_in[3][1374] , \round_in[3][1373] , 
        \round_in[3][1372] , \round_in[3][1371] , \round_in[3][1370] , 
        \round_in[3][1369] , \round_in[3][1368] , \round_in[3][1367] , 
        \round_in[3][1366] , \round_in[3][1365] , \round_in[3][1364] , 
        \round_in[3][1363] , \round_in[3][1362] , \round_in[3][1361] , 
        \round_in[3][1360] , \round_in[3][1359] , \round_in[3][1358] , 
        \round_in[3][1357] , \round_in[3][1356] , \round_in[3][1355] , 
        \round_in[3][1354] , \round_in[3][1353] , \round_in[3][1352] , 
        \round_in[3][1351] , \round_in[3][1350] , \round_in[3][1349] , 
        \round_in[3][1348] , \round_in[3][1347] , \round_in[3][1346] , 
        \round_in[3][1345] , \round_in[3][1344] , \round_in[3][1343] , 
        \round_in[3][1342] , \round_in[3][1341] , \round_in[3][1340] , 
        \round_in[3][1339] , \round_in[3][1338] , \round_in[3][1337] , 
        \round_in[3][1336] , \round_in[3][1335] , \round_in[3][1334] , 
        \round_in[3][1333] , \round_in[3][1332] , \round_in[3][1331] , 
        \round_in[3][1330] , \round_in[3][1329] , \round_in[3][1328] , 
        \round_in[3][1327] , \round_in[3][1326] , \round_in[3][1325] , 
        \round_in[3][1324] , \round_in[3][1323] , \round_in[3][1322] , 
        \round_in[3][1321] , \round_in[3][1320] , \round_in[3][1319] , 
        \round_in[3][1318] , \round_in[3][1317] , \round_in[3][1316] , 
        \round_in[3][1315] , \round_in[3][1314] , \round_in[3][1313] , 
        \round_in[3][1312] , \round_in[3][1311] , \round_in[3][1310] , 
        \round_in[3][1309] , \round_in[3][1308] , \round_in[3][1307] , 
        \round_in[3][1306] , \round_in[3][1305] , \round_in[3][1304] , 
        \round_in[3][1303] , \round_in[3][1302] , \round_in[3][1301] , 
        \round_in[3][1300] , \round_in[3][1299] , \round_in[3][1298] , 
        \round_in[3][1297] , \round_in[3][1296] , \round_in[3][1295] , 
        \round_in[3][1294] , \round_in[3][1293] , \round_in[3][1292] , 
        \round_in[3][1291] , \round_in[3][1290] , \round_in[3][1289] , 
        \round_in[3][1288] , \round_in[3][1287] , \round_in[3][1286] , 
        \round_in[3][1285] , \round_in[3][1284] , \round_in[3][1283] , 
        \round_in[3][1282] , \round_in[3][1281] , \round_in[3][1280] , 
        \round_in[3][1279] , \round_in[3][1278] , \round_in[3][1277] , 
        \round_in[3][1276] , \round_in[3][1275] , \round_in[3][1274] , 
        \round_in[3][1273] , \round_in[3][1272] , \round_in[3][1271] , 
        \round_in[3][1270] , \round_in[3][1269] , \round_in[3][1268] , 
        \round_in[3][1267] , \round_in[3][1266] , \round_in[3][1265] , 
        \round_in[3][1264] , \round_in[3][1263] , \round_in[3][1262] , 
        \round_in[3][1261] , \round_in[3][1260] , \round_in[3][1259] , 
        \round_in[3][1258] , \round_in[3][1257] , \round_in[3][1256] , 
        \round_in[3][1255] , \round_in[3][1254] , \round_in[3][1253] , 
        \round_in[3][1252] , \round_in[3][1251] , \round_in[3][1250] , 
        \round_in[3][1249] , \round_in[3][1248] , \round_in[3][1247] , 
        \round_in[3][1246] , \round_in[3][1245] , \round_in[3][1244] , 
        \round_in[3][1243] , \round_in[3][1242] , \round_in[3][1241] , 
        \round_in[3][1240] , \round_in[3][1239] , \round_in[3][1238] , 
        \round_in[3][1237] , \round_in[3][1236] , \round_in[3][1235] , 
        \round_in[3][1234] , \round_in[3][1233] , \round_in[3][1232] , 
        \round_in[3][1231] , \round_in[3][1230] , \round_in[3][1229] , 
        \round_in[3][1228] , \round_in[3][1227] , \round_in[3][1226] , 
        \round_in[3][1225] , \round_in[3][1224] , \round_in[3][1223] , 
        \round_in[3][1222] , \round_in[3][1221] , \round_in[3][1220] , 
        \round_in[3][1219] , \round_in[3][1218] , \round_in[3][1217] , 
        \round_in[3][1216] , \round_in[3][1215] , \round_in[3][1214] , 
        \round_in[3][1213] , \round_in[3][1212] , \round_in[3][1211] , 
        \round_in[3][1210] , \round_in[3][1209] , \round_in[3][1208] , 
        \round_in[3][1207] , \round_in[3][1206] , \round_in[3][1205] , 
        \round_in[3][1204] , \round_in[3][1203] , \round_in[3][1202] , 
        \round_in[3][1201] , \round_in[3][1200] , \round_in[3][1199] , 
        \round_in[3][1198] , \round_in[3][1197] , \round_in[3][1196] , 
        \round_in[3][1195] , \round_in[3][1194] , \round_in[3][1193] , 
        \round_in[3][1192] , \round_in[3][1191] , \round_in[3][1190] , 
        \round_in[3][1189] , \round_in[3][1188] , \round_in[3][1187] , 
        \round_in[3][1186] , \round_in[3][1185] , \round_in[3][1184] , 
        \round_in[3][1183] , \round_in[3][1182] , \round_in[3][1181] , 
        \round_in[3][1180] , \round_in[3][1179] , \round_in[3][1178] , 
        \round_in[3][1177] , \round_in[3][1176] , \round_in[3][1175] , 
        \round_in[3][1174] , \round_in[3][1173] , \round_in[3][1172] , 
        \round_in[3][1171] , \round_in[3][1170] , \round_in[3][1169] , 
        \round_in[3][1168] , \round_in[3][1167] , \round_in[3][1166] , 
        \round_in[3][1165] , \round_in[3][1164] , \round_in[3][1163] , 
        \round_in[3][1162] , \round_in[3][1161] , \round_in[3][1160] , 
        \round_in[3][1159] , \round_in[3][1158] , \round_in[3][1157] , 
        \round_in[3][1156] , \round_in[3][1155] , \round_in[3][1154] , 
        \round_in[3][1153] , \round_in[3][1152] , \round_in[3][1151] , 
        \round_in[3][1150] , \round_in[3][1149] , \round_in[3][1148] , 
        \round_in[3][1147] , \round_in[3][1146] , \round_in[3][1145] , 
        \round_in[3][1144] , \round_in[3][1143] , \round_in[3][1142] , 
        \round_in[3][1141] , \round_in[3][1140] , \round_in[3][1139] , 
        \round_in[3][1138] , \round_in[3][1137] , \round_in[3][1136] , 
        \round_in[3][1135] , \round_in[3][1134] , \round_in[3][1133] , 
        \round_in[3][1132] , \round_in[3][1131] , \round_in[3][1130] , 
        \round_in[3][1129] , \round_in[3][1128] , \round_in[3][1127] , 
        \round_in[3][1126] , \round_in[3][1125] , \round_in[3][1124] , 
        \round_in[3][1123] , \round_in[3][1122] , \round_in[3][1121] , 
        \round_in[3][1120] , \round_in[3][1119] , \round_in[3][1118] , 
        \round_in[3][1117] , \round_in[3][1116] , \round_in[3][1115] , 
        \round_in[3][1114] , \round_in[3][1113] , \round_in[3][1112] , 
        \round_in[3][1111] , \round_in[3][1110] , \round_in[3][1109] , 
        \round_in[3][1108] , \round_in[3][1107] , \round_in[3][1106] , 
        \round_in[3][1105] , \round_in[3][1104] , \round_in[3][1103] , 
        \round_in[3][1102] , \round_in[3][1101] , \round_in[3][1100] , 
        \round_in[3][1099] , \round_in[3][1098] , \round_in[3][1097] , 
        \round_in[3][1096] , \round_in[3][1095] , \round_in[3][1094] , 
        \round_in[3][1093] , \round_in[3][1092] , \round_in[3][1091] , 
        \round_in[3][1090] , \round_in[3][1089] , \round_in[3][1088] , 
        \round_in[3][1087] , \round_in[3][1086] , \round_in[3][1085] , 
        \round_in[3][1084] , \round_in[3][1083] , \round_in[3][1082] , 
        \round_in[3][1081] , \round_in[3][1080] , \round_in[3][1079] , 
        \round_in[3][1078] , \round_in[3][1077] , \round_in[3][1076] , 
        \round_in[3][1075] , \round_in[3][1074] , \round_in[3][1073] , 
        \round_in[3][1072] , \round_in[3][1071] , \round_in[3][1070] , 
        \round_in[3][1069] , \round_in[3][1068] , \round_in[3][1067] , 
        \round_in[3][1066] , \round_in[3][1065] , \round_in[3][1064] , 
        \round_in[3][1063] , \round_in[3][1062] , \round_in[3][1061] , 
        \round_in[3][1060] , \round_in[3][1059] , \round_in[3][1058] , 
        \round_in[3][1057] , \round_in[3][1056] , \round_in[3][1055] , 
        \round_in[3][1054] , \round_in[3][1053] , \round_in[3][1052] , 
        \round_in[3][1051] , \round_in[3][1050] , \round_in[3][1049] , 
        \round_in[3][1048] , \round_in[3][1047] , \round_in[3][1046] , 
        \round_in[3][1045] , \round_in[3][1044] , \round_in[3][1043] , 
        \round_in[3][1042] , \round_in[3][1041] , \round_in[3][1040] , 
        \round_in[3][1039] , \round_in[3][1038] , \round_in[3][1037] , 
        \round_in[3][1036] , \round_in[3][1035] , \round_in[3][1034] , 
        \round_in[3][1033] , \round_in[3][1032] , \round_in[3][1031] , 
        \round_in[3][1030] , \round_in[3][1029] , \round_in[3][1028] , 
        \round_in[3][1027] , \round_in[3][1026] , \round_in[3][1025] , 
        \round_in[3][1024] , \round_in[3][1023] , \round_in[3][1022] , 
        \round_in[3][1021] , \round_in[3][1020] , \round_in[3][1019] , 
        \round_in[3][1018] , \round_in[3][1017] , \round_in[3][1016] , 
        \round_in[3][1015] , \round_in[3][1014] , \round_in[3][1013] , 
        \round_in[3][1012] , \round_in[3][1011] , \round_in[3][1010] , 
        \round_in[3][1009] , \round_in[3][1008] , \round_in[3][1007] , 
        \round_in[3][1006] , \round_in[3][1005] , \round_in[3][1004] , 
        \round_in[3][1003] , \round_in[3][1002] , \round_in[3][1001] , 
        \round_in[3][1000] , \round_in[3][999] , \round_in[3][998] , 
        \round_in[3][997] , \round_in[3][996] , \round_in[3][995] , 
        \round_in[3][994] , \round_in[3][993] , \round_in[3][992] , 
        \round_in[3][991] , \round_in[3][990] , \round_in[3][989] , 
        \round_in[3][988] , \round_in[3][987] , \round_in[3][986] , 
        \round_in[3][985] , \round_in[3][984] , \round_in[3][983] , 
        \round_in[3][982] , \round_in[3][981] , \round_in[3][980] , 
        \round_in[3][979] , \round_in[3][978] , \round_in[3][977] , 
        \round_in[3][976] , \round_in[3][975] , \round_in[3][974] , 
        \round_in[3][973] , \round_in[3][972] , \round_in[3][971] , 
        \round_in[3][970] , \round_in[3][969] , \round_in[3][968] , 
        \round_in[3][967] , \round_in[3][966] , \round_in[3][965] , 
        \round_in[3][964] , \round_in[3][963] , \round_in[3][962] , 
        \round_in[3][961] , \round_in[3][960] , \round_in[3][959] , 
        \round_in[3][958] , \round_in[3][957] , \round_in[3][956] , 
        \round_in[3][955] , \round_in[3][954] , \round_in[3][953] , 
        \round_in[3][952] , \round_in[3][951] , \round_in[3][950] , 
        \round_in[3][949] , \round_in[3][948] , \round_in[3][947] , 
        \round_in[3][946] , \round_in[3][945] , \round_in[3][944] , 
        \round_in[3][943] , \round_in[3][942] , \round_in[3][941] , 
        \round_in[3][940] , \round_in[3][939] , \round_in[3][938] , 
        \round_in[3][937] , \round_in[3][936] , \round_in[3][935] , 
        \round_in[3][934] , \round_in[3][933] , \round_in[3][932] , 
        \round_in[3][931] , \round_in[3][930] , \round_in[3][929] , 
        \round_in[3][928] , \round_in[3][927] , \round_in[3][926] , 
        \round_in[3][925] , \round_in[3][924] , \round_in[3][923] , 
        \round_in[3][922] , \round_in[3][921] , \round_in[3][920] , 
        \round_in[3][919] , \round_in[3][918] , \round_in[3][917] , 
        \round_in[3][916] , \round_in[3][915] , \round_in[3][914] , 
        \round_in[3][913] , \round_in[3][912] , \round_in[3][911] , 
        \round_in[3][910] , \round_in[3][909] , \round_in[3][908] , 
        \round_in[3][907] , \round_in[3][906] , \round_in[3][905] , 
        \round_in[3][904] , \round_in[3][903] , \round_in[3][902] , 
        \round_in[3][901] , \round_in[3][900] , \round_in[3][899] , 
        \round_in[3][898] , \round_in[3][897] , \round_in[3][896] , 
        \round_in[3][895] , \round_in[3][894] , \round_in[3][893] , 
        \round_in[3][892] , \round_in[3][891] , \round_in[3][890] , 
        \round_in[3][889] , \round_in[3][888] , \round_in[3][887] , 
        \round_in[3][886] , \round_in[3][885] , \round_in[3][884] , 
        \round_in[3][883] , \round_in[3][882] , \round_in[3][881] , 
        \round_in[3][880] , \round_in[3][879] , \round_in[3][878] , 
        \round_in[3][877] , \round_in[3][876] , \round_in[3][875] , 
        \round_in[3][874] , \round_in[3][873] , \round_in[3][872] , 
        \round_in[3][871] , \round_in[3][870] , \round_in[3][869] , 
        \round_in[3][868] , \round_in[3][867] , \round_in[3][866] , 
        \round_in[3][865] , \round_in[3][864] , \round_in[3][863] , 
        \round_in[3][862] , \round_in[3][861] , \round_in[3][860] , 
        \round_in[3][859] , \round_in[3][858] , \round_in[3][857] , 
        \round_in[3][856] , \round_in[3][855] , \round_in[3][854] , 
        \round_in[3][853] , \round_in[3][852] , \round_in[3][851] , 
        \round_in[3][850] , \round_in[3][849] , \round_in[3][848] , 
        \round_in[3][847] , \round_in[3][846] , \round_in[3][845] , 
        \round_in[3][844] , \round_in[3][843] , \round_in[3][842] , 
        \round_in[3][841] , \round_in[3][840] , \round_in[3][839] , 
        \round_in[3][838] , \round_in[3][837] , \round_in[3][836] , 
        \round_in[3][835] , \round_in[3][834] , \round_in[3][833] , 
        \round_in[3][832] , \round_in[3][831] , \round_in[3][830] , 
        \round_in[3][829] , \round_in[3][828] , \round_in[3][827] , 
        \round_in[3][826] , \round_in[3][825] , \round_in[3][824] , 
        \round_in[3][823] , \round_in[3][822] , \round_in[3][821] , 
        \round_in[3][820] , \round_in[3][819] , \round_in[3][818] , 
        \round_in[3][817] , \round_in[3][816] , \round_in[3][815] , 
        \round_in[3][814] , \round_in[3][813] , \round_in[3][812] , 
        \round_in[3][811] , \round_in[3][810] , \round_in[3][809] , 
        \round_in[3][808] , \round_in[3][807] , \round_in[3][806] , 
        \round_in[3][805] , \round_in[3][804] , \round_in[3][803] , 
        \round_in[3][802] , \round_in[3][801] , \round_in[3][800] , 
        \round_in[3][799] , \round_in[3][798] , \round_in[3][797] , 
        \round_in[3][796] , \round_in[3][795] , \round_in[3][794] , 
        \round_in[3][793] , \round_in[3][792] , \round_in[3][791] , 
        \round_in[3][790] , \round_in[3][789] , \round_in[3][788] , 
        \round_in[3][787] , \round_in[3][786] , \round_in[3][785] , 
        \round_in[3][784] , \round_in[3][783] , \round_in[3][782] , 
        \round_in[3][781] , \round_in[3][780] , \round_in[3][779] , 
        \round_in[3][778] , \round_in[3][777] , \round_in[3][776] , 
        \round_in[3][775] , \round_in[3][774] , \round_in[3][773] , 
        \round_in[3][772] , \round_in[3][771] , \round_in[3][770] , 
        \round_in[3][769] , \round_in[3][768] , \round_in[3][767] , 
        \round_in[3][766] , \round_in[3][765] , \round_in[3][764] , 
        \round_in[3][763] , \round_in[3][762] , \round_in[3][761] , 
        \round_in[3][760] , \round_in[3][759] , \round_in[3][758] , 
        \round_in[3][757] , \round_in[3][756] , \round_in[3][755] , 
        \round_in[3][754] , \round_in[3][753] , \round_in[3][752] , 
        \round_in[3][751] , \round_in[3][750] , \round_in[3][749] , 
        \round_in[3][748] , \round_in[3][747] , \round_in[3][746] , 
        \round_in[3][745] , \round_in[3][744] , \round_in[3][743] , 
        \round_in[3][742] , \round_in[3][741] , \round_in[3][740] , 
        \round_in[3][739] , \round_in[3][738] , \round_in[3][737] , 
        \round_in[3][736] , \round_in[3][735] , \round_in[3][734] , 
        \round_in[3][733] , \round_in[3][732] , \round_in[3][731] , 
        \round_in[3][730] , \round_in[3][729] , \round_in[3][728] , 
        \round_in[3][727] , \round_in[3][726] , \round_in[3][725] , 
        \round_in[3][724] , \round_in[3][723] , \round_in[3][722] , 
        \round_in[3][721] , \round_in[3][720] , \round_in[3][719] , 
        \round_in[3][718] , \round_in[3][717] , \round_in[3][716] , 
        \round_in[3][715] , \round_in[3][714] , \round_in[3][713] , 
        \round_in[3][712] , \round_in[3][711] , \round_in[3][710] , 
        \round_in[3][709] , \round_in[3][708] , \round_in[3][707] , 
        \round_in[3][706] , \round_in[3][705] , \round_in[3][704] , 
        \round_in[3][703] , \round_in[3][702] , \round_in[3][701] , 
        \round_in[3][700] , \round_in[3][699] , \round_in[3][698] , 
        \round_in[3][697] , \round_in[3][696] , \round_in[3][695] , 
        \round_in[3][694] , \round_in[3][693] , \round_in[3][692] , 
        \round_in[3][691] , \round_in[3][690] , \round_in[3][689] , 
        \round_in[3][688] , \round_in[3][687] , \round_in[3][686] , 
        \round_in[3][685] , \round_in[3][684] , \round_in[3][683] , 
        \round_in[3][682] , \round_in[3][681] , \round_in[3][680] , 
        \round_in[3][679] , \round_in[3][678] , \round_in[3][677] , 
        \round_in[3][676] , \round_in[3][675] , \round_in[3][674] , 
        \round_in[3][673] , \round_in[3][672] , \round_in[3][671] , 
        \round_in[3][670] , \round_in[3][669] , \round_in[3][668] , 
        \round_in[3][667] , \round_in[3][666] , \round_in[3][665] , 
        \round_in[3][664] , \round_in[3][663] , \round_in[3][662] , 
        \round_in[3][661] , \round_in[3][660] , \round_in[3][659] , 
        \round_in[3][658] , \round_in[3][657] , \round_in[3][656] , 
        \round_in[3][655] , \round_in[3][654] , \round_in[3][653] , 
        \round_in[3][652] , \round_in[3][651] , \round_in[3][650] , 
        \round_in[3][649] , \round_in[3][648] , \round_in[3][647] , 
        \round_in[3][646] , \round_in[3][645] , \round_in[3][644] , 
        \round_in[3][643] , \round_in[3][642] , \round_in[3][641] , 
        \round_in[3][640] , \round_in[3][639] , \round_in[3][638] , 
        \round_in[3][637] , \round_in[3][636] , \round_in[3][635] , 
        \round_in[3][634] , \round_in[3][633] , \round_in[3][632] , 
        \round_in[3][631] , \round_in[3][630] , \round_in[3][629] , 
        \round_in[3][628] , \round_in[3][627] , \round_in[3][626] , 
        \round_in[3][625] , \round_in[3][624] , \round_in[3][623] , 
        \round_in[3][622] , \round_in[3][621] , \round_in[3][620] , 
        \round_in[3][619] , \round_in[3][618] , \round_in[3][617] , 
        \round_in[3][616] , \round_in[3][615] , \round_in[3][614] , 
        \round_in[3][613] , \round_in[3][612] , \round_in[3][611] , 
        \round_in[3][610] , \round_in[3][609] , \round_in[3][608] , 
        \round_in[3][607] , \round_in[3][606] , \round_in[3][605] , 
        \round_in[3][604] , \round_in[3][603] , \round_in[3][602] , 
        \round_in[3][601] , \round_in[3][600] , \round_in[3][599] , 
        \round_in[3][598] , \round_in[3][597] , \round_in[3][596] , 
        \round_in[3][595] , \round_in[3][594] , \round_in[3][593] , 
        \round_in[3][592] , \round_in[3][591] , \round_in[3][590] , 
        \round_in[3][589] , \round_in[3][588] , \round_in[3][587] , 
        \round_in[3][586] , \round_in[3][585] , \round_in[3][584] , 
        \round_in[3][583] , \round_in[3][582] , \round_in[3][581] , 
        \round_in[3][580] , \round_in[3][579] , \round_in[3][578] , 
        \round_in[3][577] , \round_in[3][576] , \round_in[3][575] , 
        \round_in[3][574] , \round_in[3][573] , \round_in[3][572] , 
        \round_in[3][571] , \round_in[3][570] , \round_in[3][569] , 
        \round_in[3][568] , \round_in[3][567] , \round_in[3][566] , 
        \round_in[3][565] , \round_in[3][564] , \round_in[3][563] , 
        \round_in[3][562] , \round_in[3][561] , \round_in[3][560] , 
        \round_in[3][559] , \round_in[3][558] , \round_in[3][557] , 
        \round_in[3][556] , \round_in[3][555] , \round_in[3][554] , 
        \round_in[3][553] , \round_in[3][552] , \round_in[3][551] , 
        \round_in[3][550] , \round_in[3][549] , \round_in[3][548] , 
        \round_in[3][547] , \round_in[3][546] , \round_in[3][545] , 
        \round_in[3][544] , \round_in[3][543] , \round_in[3][542] , 
        \round_in[3][541] , \round_in[3][540] , \round_in[3][539] , 
        \round_in[3][538] , \round_in[3][537] , \round_in[3][536] , 
        \round_in[3][535] , \round_in[3][534] , \round_in[3][533] , 
        \round_in[3][532] , \round_in[3][531] , \round_in[3][530] , 
        \round_in[3][529] , \round_in[3][528] , \round_in[3][527] , 
        \round_in[3][526] , \round_in[3][525] , \round_in[3][524] , 
        \round_in[3][523] , \round_in[3][522] , \round_in[3][521] , 
        \round_in[3][520] , \round_in[3][519] , \round_in[3][518] , 
        \round_in[3][517] , \round_in[3][516] , \round_in[3][515] , 
        \round_in[3][514] , \round_in[3][513] , \round_in[3][512] , 
        \round_in[3][511] , \round_in[3][510] , \round_in[3][509] , 
        \round_in[3][508] , \round_in[3][507] , \round_in[3][506] , 
        \round_in[3][505] , \round_in[3][504] , \round_in[3][503] , 
        \round_in[3][502] , \round_in[3][501] , \round_in[3][500] , 
        \round_in[3][499] , \round_in[3][498] , \round_in[3][497] , 
        \round_in[3][496] , \round_in[3][495] , \round_in[3][494] , 
        \round_in[3][493] , \round_in[3][492] , \round_in[3][491] , 
        \round_in[3][490] , \round_in[3][489] , \round_in[3][488] , 
        \round_in[3][487] , \round_in[3][486] , \round_in[3][485] , 
        \round_in[3][484] , \round_in[3][483] , \round_in[3][482] , 
        \round_in[3][481] , \round_in[3][480] , \round_in[3][479] , 
        \round_in[3][478] , \round_in[3][477] , \round_in[3][476] , 
        \round_in[3][475] , \round_in[3][474] , \round_in[3][473] , 
        \round_in[3][472] , \round_in[3][471] , \round_in[3][470] , 
        \round_in[3][469] , \round_in[3][468] , \round_in[3][467] , 
        \round_in[3][466] , \round_in[3][465] , \round_in[3][464] , 
        \round_in[3][463] , \round_in[3][462] , \round_in[3][461] , 
        \round_in[3][460] , \round_in[3][459] , \round_in[3][458] , 
        \round_in[3][457] , \round_in[3][456] , \round_in[3][455] , 
        \round_in[3][454] , \round_in[3][453] , \round_in[3][452] , 
        \round_in[3][451] , \round_in[3][450] , \round_in[3][449] , 
        \round_in[3][448] , \round_in[3][447] , \round_in[3][446] , 
        \round_in[3][445] , \round_in[3][444] , \round_in[3][443] , 
        \round_in[3][442] , \round_in[3][441] , \round_in[3][440] , 
        \round_in[3][439] , \round_in[3][438] , \round_in[3][437] , 
        \round_in[3][436] , \round_in[3][435] , \round_in[3][434] , 
        \round_in[3][433] , \round_in[3][432] , \round_in[3][431] , 
        \round_in[3][430] , \round_in[3][429] , \round_in[3][428] , 
        \round_in[3][427] , \round_in[3][426] , \round_in[3][425] , 
        \round_in[3][424] , \round_in[3][423] , \round_in[3][422] , 
        \round_in[3][421] , \round_in[3][420] , \round_in[3][419] , 
        \round_in[3][418] , \round_in[3][417] , \round_in[3][416] , 
        \round_in[3][415] , \round_in[3][414] , \round_in[3][413] , 
        \round_in[3][412] , \round_in[3][411] , \round_in[3][410] , 
        \round_in[3][409] , \round_in[3][408] , \round_in[3][407] , 
        \round_in[3][406] , \round_in[3][405] , \round_in[3][404] , 
        \round_in[3][403] , \round_in[3][402] , \round_in[3][401] , 
        \round_in[3][400] , \round_in[3][399] , \round_in[3][398] , 
        \round_in[3][397] , \round_in[3][396] , \round_in[3][395] , 
        \round_in[3][394] , \round_in[3][393] , \round_in[3][392] , 
        \round_in[3][391] , \round_in[3][390] , \round_in[3][389] , 
        \round_in[3][388] , \round_in[3][387] , \round_in[3][386] , 
        \round_in[3][385] , \round_in[3][384] , \round_in[3][383] , 
        \round_in[3][382] , \round_in[3][381] , \round_in[3][380] , 
        \round_in[3][379] , \round_in[3][378] , \round_in[3][377] , 
        \round_in[3][376] , \round_in[3][375] , \round_in[3][374] , 
        \round_in[3][373] , \round_in[3][372] , \round_in[3][371] , 
        \round_in[3][370] , \round_in[3][369] , \round_in[3][368] , 
        \round_in[3][367] , \round_in[3][366] , \round_in[3][365] , 
        \round_in[3][364] , \round_in[3][363] , \round_in[3][362] , 
        \round_in[3][361] , \round_in[3][360] , \round_in[3][359] , 
        \round_in[3][358] , \round_in[3][357] , \round_in[3][356] , 
        \round_in[3][355] , \round_in[3][354] , \round_in[3][353] , 
        \round_in[3][352] , \round_in[3][351] , \round_in[3][350] , 
        \round_in[3][349] , \round_in[3][348] , \round_in[3][347] , 
        \round_in[3][346] , \round_in[3][345] , \round_in[3][344] , 
        \round_in[3][343] , \round_in[3][342] , \round_in[3][341] , 
        \round_in[3][340] , \round_in[3][339] , \round_in[3][338] , 
        \round_in[3][337] , \round_in[3][336] , \round_in[3][335] , 
        \round_in[3][334] , \round_in[3][333] , \round_in[3][332] , 
        \round_in[3][331] , \round_in[3][330] , \round_in[3][329] , 
        \round_in[3][328] , \round_in[3][327] , \round_in[3][326] , 
        \round_in[3][325] , \round_in[3][324] , \round_in[3][323] , 
        \round_in[3][322] , \round_in[3][321] , \round_in[3][320] , 
        \round_in[3][319] , \round_in[3][318] , \round_in[3][317] , 
        \round_in[3][316] , \round_in[3][315] , \round_in[3][314] , 
        \round_in[3][313] , \round_in[3][312] , \round_in[3][311] , 
        \round_in[3][310] , \round_in[3][309] , \round_in[3][308] , 
        \round_in[3][307] , \round_in[3][306] , \round_in[3][305] , 
        \round_in[3][304] , \round_in[3][303] , \round_in[3][302] , 
        \round_in[3][301] , \round_in[3][300] , \round_in[3][299] , 
        \round_in[3][298] , \round_in[3][297] , \round_in[3][296] , 
        \round_in[3][295] , \round_in[3][294] , \round_in[3][293] , 
        \round_in[3][292] , \round_in[3][291] , \round_in[3][290] , 
        \round_in[3][289] , \round_in[3][288] , \round_in[3][287] , 
        \round_in[3][286] , \round_in[3][285] , \round_in[3][284] , 
        \round_in[3][283] , \round_in[3][282] , \round_in[3][281] , 
        \round_in[3][280] , \round_in[3][279] , \round_in[3][278] , 
        \round_in[3][277] , \round_in[3][276] , \round_in[3][275] , 
        \round_in[3][274] , \round_in[3][273] , \round_in[3][272] , 
        \round_in[3][271] , \round_in[3][270] , \round_in[3][269] , 
        \round_in[3][268] , \round_in[3][267] , \round_in[3][266] , 
        \round_in[3][265] , \round_in[3][264] , \round_in[3][263] , 
        \round_in[3][262] , \round_in[3][261] , \round_in[3][260] , 
        \round_in[3][259] , \round_in[3][258] , \round_in[3][257] , 
        \round_in[3][256] , \round_in[3][255] , \round_in[3][254] , 
        \round_in[3][253] , \round_in[3][252] , \round_in[3][251] , 
        \round_in[3][250] , \round_in[3][249] , \round_in[3][248] , 
        \round_in[3][247] , \round_in[3][246] , \round_in[3][245] , 
        \round_in[3][244] , \round_in[3][243] , \round_in[3][242] , 
        \round_in[3][241] , \round_in[3][240] , \round_in[3][239] , 
        \round_in[3][238] , \round_in[3][237] , \round_in[3][236] , 
        \round_in[3][235] , \round_in[3][234] , \round_in[3][233] , 
        \round_in[3][232] , \round_in[3][231] , \round_in[3][230] , 
        \round_in[3][229] , \round_in[3][228] , \round_in[3][227] , 
        \round_in[3][226] , \round_in[3][225] , \round_in[3][224] , 
        \round_in[3][223] , \round_in[3][222] , \round_in[3][221] , 
        \round_in[3][220] , \round_in[3][219] , \round_in[3][218] , 
        \round_in[3][217] , \round_in[3][216] , \round_in[3][215] , 
        \round_in[3][214] , \round_in[3][213] , \round_in[3][212] , 
        \round_in[3][211] , \round_in[3][210] , \round_in[3][209] , 
        \round_in[3][208] , \round_in[3][207] , \round_in[3][206] , 
        \round_in[3][205] , \round_in[3][204] , \round_in[3][203] , 
        \round_in[3][202] , \round_in[3][201] , \round_in[3][200] , 
        \round_in[3][199] , \round_in[3][198] , \round_in[3][197] , 
        \round_in[3][196] , \round_in[3][195] , \round_in[3][194] , 
        \round_in[3][193] , \round_in[3][192] , \round_in[3][191] , 
        \round_in[3][190] , \round_in[3][189] , \round_in[3][188] , 
        \round_in[3][187] , \round_in[3][186] , \round_in[3][185] , 
        \round_in[3][184] , \round_in[3][183] , \round_in[3][182] , 
        \round_in[3][181] , \round_in[3][180] , \round_in[3][179] , 
        \round_in[3][178] , \round_in[3][177] , \round_in[3][176] , 
        \round_in[3][175] , \round_in[3][174] , \round_in[3][173] , 
        \round_in[3][172] , \round_in[3][171] , \round_in[3][170] , 
        \round_in[3][169] , \round_in[3][168] , \round_in[3][167] , 
        \round_in[3][166] , \round_in[3][165] , \round_in[3][164] , 
        \round_in[3][163] , \round_in[3][162] , \round_in[3][161] , 
        \round_in[3][160] , \round_in[3][159] , \round_in[3][158] , 
        \round_in[3][157] , \round_in[3][156] , \round_in[3][155] , 
        \round_in[3][154] , \round_in[3][153] , \round_in[3][152] , 
        \round_in[3][151] , \round_in[3][150] , \round_in[3][149] , 
        \round_in[3][148] , \round_in[3][147] , \round_in[3][146] , 
        \round_in[3][145] , \round_in[3][144] , \round_in[3][143] , 
        \round_in[3][142] , \round_in[3][141] , \round_in[3][140] , 
        \round_in[3][139] , \round_in[3][138] , \round_in[3][137] , 
        \round_in[3][136] , \round_in[3][135] , \round_in[3][134] , 
        \round_in[3][133] , \round_in[3][132] , \round_in[3][131] , 
        \round_in[3][130] , \round_in[3][129] , \round_in[3][128] , 
        \round_in[3][127] , \round_in[3][126] , \round_in[3][125] , 
        \round_in[3][124] , \round_in[3][123] , \round_in[3][122] , 
        \round_in[3][121] , \round_in[3][120] , \round_in[3][119] , 
        \round_in[3][118] , \round_in[3][117] , \round_in[3][116] , 
        \round_in[3][115] , \round_in[3][114] , \round_in[3][113] , 
        \round_in[3][112] , \round_in[3][111] , \round_in[3][110] , 
        \round_in[3][109] , \round_in[3][108] , \round_in[3][107] , 
        \round_in[3][106] , \round_in[3][105] , \round_in[3][104] , 
        \round_in[3][103] , \round_in[3][102] , \round_in[3][101] , 
        \round_in[3][100] , \round_in[3][99] , \round_in[3][98] , 
        \round_in[3][97] , \round_in[3][96] , \round_in[3][95] , 
        \round_in[3][94] , \round_in[3][93] , \round_in[3][92] , 
        \round_in[3][91] , \round_in[3][90] , \round_in[3][89] , 
        \round_in[3][88] , \round_in[3][87] , \round_in[3][86] , 
        \round_in[3][85] , \round_in[3][84] , \round_in[3][83] , 
        \round_in[3][82] , \round_in[3][81] , \round_in[3][80] , 
        \round_in[3][79] , \round_in[3][78] , \round_in[3][77] , 
        \round_in[3][76] , \round_in[3][75] , \round_in[3][74] , 
        \round_in[3][73] , \round_in[3][72] , \round_in[3][71] , 
        \round_in[3][70] , \round_in[3][69] , \round_in[3][68] , 
        \round_in[3][67] , \round_in[3][66] , \round_in[3][65] , 
        \round_in[3][64] , \round_in[3][63] , \round_in[3][62] , 
        \round_in[3][61] , \round_in[3][60] , \round_in[3][59] , 
        \round_in[3][58] , \round_in[3][57] , \round_in[3][56] , 
        \round_in[3][55] , \round_in[3][54] , \round_in[3][53] , 
        \round_in[3][52] , \round_in[3][51] , \round_in[3][50] , 
        \round_in[3][49] , \round_in[3][48] , \round_in[3][47] , 
        \round_in[3][46] , \round_in[3][45] , \round_in[3][44] , 
        \round_in[3][43] , \round_in[3][42] , \round_in[3][41] , 
        \round_in[3][40] , \round_in[3][39] , \round_in[3][38] , 
        \round_in[3][37] , \round_in[3][36] , \round_in[3][35] , 
        \round_in[3][34] , \round_in[3][33] , \round_in[3][32] , 
        \round_in[3][31] , \round_in[3][30] , \round_in[3][29] , 
        \round_in[3][28] , \round_in[3][27] , \round_in[3][26] , 
        \round_in[3][25] , \round_in[3][24] , \round_in[3][23] , 
        \round_in[3][22] , \round_in[3][21] , \round_in[3][20] , 
        \round_in[3][19] , \round_in[3][18] , \round_in[3][17] , 
        \round_in[3][16] , \round_in[3][15] , \round_in[3][14] , 
        \round_in[3][13] , \round_in[3][12] , \round_in[3][11] , 
        \round_in[3][10] , \round_in[3][9] , \round_in[3][8] , 
        \round_in[3][7] , \round_in[3][6] , \round_in[3][5] , \round_in[3][4] , 
        \round_in[3][3] , \round_in[3][2] , \round_in[3][1] , \round_in[3][0] }), .round_const({\rc[3][63] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        \rc[3][31] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \rc[3][15] , 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \rc[3][3] , 1'b0, 
        \rc[3][1] , \RCONST[3].rconst_/N10 }), .out(out) );
  DFF init_reg ( .D(n2763), .CLK(clk), .RST(1'b0), .Q(init) );
  DFF \rc_i_reg[0]  ( .D(N6), .CLK(clk), .RST(1'b0), .Q(rc_i[0]) );
  DFF \rc_i_reg[1]  ( .D(N7), .CLK(clk), .RST(1'b0), .Q(rc_i[1]) );
  DFF \rc_i_reg[2]  ( .D(N8), .CLK(clk), .RST(1'b0), .Q(rc_i[2]) );
  DFF \rc_i_reg[3]  ( .D(N9), .CLK(clk), .RST(1'b0), .Q(rc_i[3]) );
  DFF \rc_i_reg[4]  ( .D(N10), .CLK(clk), .RST(1'b0), .Q(rc_i[4]) );
  DFF \rc_i_reg[5]  ( .D(N11), .CLK(clk), .RST(1'b0), .Q(rc_i[5]) );
  DFF \round_reg_reg[0]  ( .D(N12), .CLK(clk), .RST(1'b0), .Q(round_reg[0]) );
  DFF \round_reg_reg[1]  ( .D(N13), .CLK(clk), .RST(1'b0), .Q(round_reg[1]) );
  DFF \round_reg_reg[2]  ( .D(N14), .CLK(clk), .RST(1'b0), .Q(round_reg[2]) );
  DFF \round_reg_reg[3]  ( .D(N15), .CLK(clk), .RST(1'b0), .Q(round_reg[3]) );
  DFF \round_reg_reg[4]  ( .D(N16), .CLK(clk), .RST(1'b0), .Q(round_reg[4]) );
  DFF \round_reg_reg[5]  ( .D(N17), .CLK(clk), .RST(1'b0), .Q(round_reg[5]) );
  DFF \round_reg_reg[6]  ( .D(N18), .CLK(clk), .RST(1'b0), .Q(round_reg[6]) );
  DFF \round_reg_reg[7]  ( .D(N19), .CLK(clk), .RST(1'b0), .Q(round_reg[7]) );
  DFF \round_reg_reg[8]  ( .D(N20), .CLK(clk), .RST(1'b0), .Q(round_reg[8]) );
  DFF \round_reg_reg[9]  ( .D(N21), .CLK(clk), .RST(1'b0), .Q(round_reg[9]) );
  DFF \round_reg_reg[10]  ( .D(N22), .CLK(clk), .RST(1'b0), .Q(round_reg[10])
         );
  DFF \round_reg_reg[11]  ( .D(N23), .CLK(clk), .RST(1'b0), .Q(round_reg[11])
         );
  DFF \round_reg_reg[12]  ( .D(N24), .CLK(clk), .RST(1'b0), .Q(round_reg[12])
         );
  DFF \round_reg_reg[13]  ( .D(N25), .CLK(clk), .RST(1'b0), .Q(round_reg[13])
         );
  DFF \round_reg_reg[14]  ( .D(N26), .CLK(clk), .RST(1'b0), .Q(round_reg[14])
         );
  DFF \round_reg_reg[15]  ( .D(N27), .CLK(clk), .RST(1'b0), .Q(round_reg[15])
         );
  DFF \round_reg_reg[16]  ( .D(N28), .CLK(clk), .RST(1'b0), .Q(round_reg[16])
         );
  DFF \round_reg_reg[17]  ( .D(N29), .CLK(clk), .RST(1'b0), .Q(round_reg[17])
         );
  DFF \round_reg_reg[18]  ( .D(N30), .CLK(clk), .RST(1'b0), .Q(round_reg[18])
         );
  DFF \round_reg_reg[19]  ( .D(N31), .CLK(clk), .RST(1'b0), .Q(round_reg[19])
         );
  DFF \round_reg_reg[20]  ( .D(N32), .CLK(clk), .RST(1'b0), .Q(round_reg[20])
         );
  DFF \round_reg_reg[21]  ( .D(N33), .CLK(clk), .RST(1'b0), .Q(round_reg[21])
         );
  DFF \round_reg_reg[22]  ( .D(N34), .CLK(clk), .RST(1'b0), .Q(round_reg[22])
         );
  DFF \round_reg_reg[23]  ( .D(N35), .CLK(clk), .RST(1'b0), .Q(round_reg[23])
         );
  DFF \round_reg_reg[24]  ( .D(N36), .CLK(clk), .RST(1'b0), .Q(round_reg[24])
         );
  DFF \round_reg_reg[25]  ( .D(N37), .CLK(clk), .RST(1'b0), .Q(round_reg[25])
         );
  DFF \round_reg_reg[26]  ( .D(N38), .CLK(clk), .RST(1'b0), .Q(round_reg[26])
         );
  DFF \round_reg_reg[27]  ( .D(N39), .CLK(clk), .RST(1'b0), .Q(round_reg[27])
         );
  DFF \round_reg_reg[28]  ( .D(N40), .CLK(clk), .RST(1'b0), .Q(round_reg[28])
         );
  DFF \round_reg_reg[29]  ( .D(N41), .CLK(clk), .RST(1'b0), .Q(round_reg[29])
         );
  DFF \round_reg_reg[30]  ( .D(N42), .CLK(clk), .RST(1'b0), .Q(round_reg[30])
         );
  DFF \round_reg_reg[31]  ( .D(N43), .CLK(clk), .RST(1'b0), .Q(round_reg[31])
         );
  DFF \round_reg_reg[32]  ( .D(N44), .CLK(clk), .RST(1'b0), .Q(round_reg[32])
         );
  DFF \round_reg_reg[33]  ( .D(N45), .CLK(clk), .RST(1'b0), .Q(round_reg[33])
         );
  DFF \round_reg_reg[34]  ( .D(N46), .CLK(clk), .RST(1'b0), .Q(round_reg[34])
         );
  DFF \round_reg_reg[35]  ( .D(N47), .CLK(clk), .RST(1'b0), .Q(round_reg[35])
         );
  DFF \round_reg_reg[36]  ( .D(N48), .CLK(clk), .RST(1'b0), .Q(round_reg[36])
         );
  DFF \round_reg_reg[37]  ( .D(N49), .CLK(clk), .RST(1'b0), .Q(round_reg[37])
         );
  DFF \round_reg_reg[38]  ( .D(N50), .CLK(clk), .RST(1'b0), .Q(round_reg[38])
         );
  DFF \round_reg_reg[39]  ( .D(N51), .CLK(clk), .RST(1'b0), .Q(round_reg[39])
         );
  DFF \round_reg_reg[40]  ( .D(N52), .CLK(clk), .RST(1'b0), .Q(round_reg[40])
         );
  DFF \round_reg_reg[41]  ( .D(N53), .CLK(clk), .RST(1'b0), .Q(round_reg[41])
         );
  DFF \round_reg_reg[42]  ( .D(N54), .CLK(clk), .RST(1'b0), .Q(round_reg[42])
         );
  DFF \round_reg_reg[43]  ( .D(N55), .CLK(clk), .RST(1'b0), .Q(round_reg[43])
         );
  DFF \round_reg_reg[44]  ( .D(N56), .CLK(clk), .RST(1'b0), .Q(round_reg[44])
         );
  DFF \round_reg_reg[45]  ( .D(N57), .CLK(clk), .RST(1'b0), .Q(round_reg[45])
         );
  DFF \round_reg_reg[46]  ( .D(N58), .CLK(clk), .RST(1'b0), .Q(round_reg[46])
         );
  DFF \round_reg_reg[47]  ( .D(N59), .CLK(clk), .RST(1'b0), .Q(round_reg[47])
         );
  DFF \round_reg_reg[48]  ( .D(N60), .CLK(clk), .RST(1'b0), .Q(round_reg[48])
         );
  DFF \round_reg_reg[49]  ( .D(N61), .CLK(clk), .RST(1'b0), .Q(round_reg[49])
         );
  DFF \round_reg_reg[50]  ( .D(N62), .CLK(clk), .RST(1'b0), .Q(round_reg[50])
         );
  DFF \round_reg_reg[51]  ( .D(N63), .CLK(clk), .RST(1'b0), .Q(round_reg[51])
         );
  DFF \round_reg_reg[52]  ( .D(N64), .CLK(clk), .RST(1'b0), .Q(round_reg[52])
         );
  DFF \round_reg_reg[53]  ( .D(N65), .CLK(clk), .RST(1'b0), .Q(round_reg[53])
         );
  DFF \round_reg_reg[54]  ( .D(N66), .CLK(clk), .RST(1'b0), .Q(round_reg[54])
         );
  DFF \round_reg_reg[55]  ( .D(N67), .CLK(clk), .RST(1'b0), .Q(round_reg[55])
         );
  DFF \round_reg_reg[56]  ( .D(N68), .CLK(clk), .RST(1'b0), .Q(round_reg[56])
         );
  DFF \round_reg_reg[57]  ( .D(N69), .CLK(clk), .RST(1'b0), .Q(round_reg[57])
         );
  DFF \round_reg_reg[58]  ( .D(N70), .CLK(clk), .RST(1'b0), .Q(round_reg[58])
         );
  DFF \round_reg_reg[59]  ( .D(N71), .CLK(clk), .RST(1'b0), .Q(round_reg[59])
         );
  DFF \round_reg_reg[60]  ( .D(N72), .CLK(clk), .RST(1'b0), .Q(round_reg[60])
         );
  DFF \round_reg_reg[61]  ( .D(N73), .CLK(clk), .RST(1'b0), .Q(round_reg[61])
         );
  DFF \round_reg_reg[62]  ( .D(N74), .CLK(clk), .RST(1'b0), .Q(round_reg[62])
         );
  DFF \round_reg_reg[63]  ( .D(N75), .CLK(clk), .RST(1'b0), .Q(round_reg[63])
         );
  DFF \round_reg_reg[64]  ( .D(N76), .CLK(clk), .RST(1'b0), .Q(round_reg[64])
         );
  DFF \round_reg_reg[65]  ( .D(N77), .CLK(clk), .RST(1'b0), .Q(round_reg[65])
         );
  DFF \round_reg_reg[66]  ( .D(N78), .CLK(clk), .RST(1'b0), .Q(round_reg[66])
         );
  DFF \round_reg_reg[67]  ( .D(N79), .CLK(clk), .RST(1'b0), .Q(round_reg[67])
         );
  DFF \round_reg_reg[68]  ( .D(N80), .CLK(clk), .RST(1'b0), .Q(round_reg[68])
         );
  DFF \round_reg_reg[69]  ( .D(N81), .CLK(clk), .RST(1'b0), .Q(round_reg[69])
         );
  DFF \round_reg_reg[70]  ( .D(N82), .CLK(clk), .RST(1'b0), .Q(round_reg[70])
         );
  DFF \round_reg_reg[71]  ( .D(N83), .CLK(clk), .RST(1'b0), .Q(round_reg[71])
         );
  DFF \round_reg_reg[72]  ( .D(N84), .CLK(clk), .RST(1'b0), .Q(round_reg[72])
         );
  DFF \round_reg_reg[73]  ( .D(N85), .CLK(clk), .RST(1'b0), .Q(round_reg[73])
         );
  DFF \round_reg_reg[74]  ( .D(N86), .CLK(clk), .RST(1'b0), .Q(round_reg[74])
         );
  DFF \round_reg_reg[75]  ( .D(N87), .CLK(clk), .RST(1'b0), .Q(round_reg[75])
         );
  DFF \round_reg_reg[76]  ( .D(N88), .CLK(clk), .RST(1'b0), .Q(round_reg[76])
         );
  DFF \round_reg_reg[77]  ( .D(N89), .CLK(clk), .RST(1'b0), .Q(round_reg[77])
         );
  DFF \round_reg_reg[78]  ( .D(N90), .CLK(clk), .RST(1'b0), .Q(round_reg[78])
         );
  DFF \round_reg_reg[79]  ( .D(N91), .CLK(clk), .RST(1'b0), .Q(round_reg[79])
         );
  DFF \round_reg_reg[80]  ( .D(N92), .CLK(clk), .RST(1'b0), .Q(round_reg[80])
         );
  DFF \round_reg_reg[81]  ( .D(N93), .CLK(clk), .RST(1'b0), .Q(round_reg[81])
         );
  DFF \round_reg_reg[82]  ( .D(N94), .CLK(clk), .RST(1'b0), .Q(round_reg[82])
         );
  DFF \round_reg_reg[83]  ( .D(N95), .CLK(clk), .RST(1'b0), .Q(round_reg[83])
         );
  DFF \round_reg_reg[84]  ( .D(N96), .CLK(clk), .RST(1'b0), .Q(round_reg[84])
         );
  DFF \round_reg_reg[85]  ( .D(N97), .CLK(clk), .RST(1'b0), .Q(round_reg[85])
         );
  DFF \round_reg_reg[86]  ( .D(N98), .CLK(clk), .RST(1'b0), .Q(round_reg[86])
         );
  DFF \round_reg_reg[87]  ( .D(N99), .CLK(clk), .RST(1'b0), .Q(round_reg[87])
         );
  DFF \round_reg_reg[88]  ( .D(N100), .CLK(clk), .RST(1'b0), .Q(round_reg[88])
         );
  DFF \round_reg_reg[89]  ( .D(N101), .CLK(clk), .RST(1'b0), .Q(round_reg[89])
         );
  DFF \round_reg_reg[90]  ( .D(N102), .CLK(clk), .RST(1'b0), .Q(round_reg[90])
         );
  DFF \round_reg_reg[91]  ( .D(N103), .CLK(clk), .RST(1'b0), .Q(round_reg[91])
         );
  DFF \round_reg_reg[92]  ( .D(N104), .CLK(clk), .RST(1'b0), .Q(round_reg[92])
         );
  DFF \round_reg_reg[93]  ( .D(N105), .CLK(clk), .RST(1'b0), .Q(round_reg[93])
         );
  DFF \round_reg_reg[94]  ( .D(N106), .CLK(clk), .RST(1'b0), .Q(round_reg[94])
         );
  DFF \round_reg_reg[95]  ( .D(N107), .CLK(clk), .RST(1'b0), .Q(round_reg[95])
         );
  DFF \round_reg_reg[96]  ( .D(N108), .CLK(clk), .RST(1'b0), .Q(round_reg[96])
         );
  DFF \round_reg_reg[97]  ( .D(N109), .CLK(clk), .RST(1'b0), .Q(round_reg[97])
         );
  DFF \round_reg_reg[98]  ( .D(N110), .CLK(clk), .RST(1'b0), .Q(round_reg[98])
         );
  DFF \round_reg_reg[99]  ( .D(N111), .CLK(clk), .RST(1'b0), .Q(round_reg[99])
         );
  DFF \round_reg_reg[100]  ( .D(N112), .CLK(clk), .RST(1'b0), .Q(
        round_reg[100]) );
  DFF \round_reg_reg[101]  ( .D(N113), .CLK(clk), .RST(1'b0), .Q(
        round_reg[101]) );
  DFF \round_reg_reg[102]  ( .D(N114), .CLK(clk), .RST(1'b0), .Q(
        round_reg[102]) );
  DFF \round_reg_reg[103]  ( .D(N115), .CLK(clk), .RST(1'b0), .Q(
        round_reg[103]) );
  DFF \round_reg_reg[104]  ( .D(N116), .CLK(clk), .RST(1'b0), .Q(
        round_reg[104]) );
  DFF \round_reg_reg[105]  ( .D(N117), .CLK(clk), .RST(1'b0), .Q(
        round_reg[105]) );
  DFF \round_reg_reg[106]  ( .D(N118), .CLK(clk), .RST(1'b0), .Q(
        round_reg[106]) );
  DFF \round_reg_reg[107]  ( .D(N119), .CLK(clk), .RST(1'b0), .Q(
        round_reg[107]) );
  DFF \round_reg_reg[108]  ( .D(N120), .CLK(clk), .RST(1'b0), .Q(
        round_reg[108]) );
  DFF \round_reg_reg[109]  ( .D(N121), .CLK(clk), .RST(1'b0), .Q(
        round_reg[109]) );
  DFF \round_reg_reg[110]  ( .D(N122), .CLK(clk), .RST(1'b0), .Q(
        round_reg[110]) );
  DFF \round_reg_reg[111]  ( .D(N123), .CLK(clk), .RST(1'b0), .Q(
        round_reg[111]) );
  DFF \round_reg_reg[112]  ( .D(N124), .CLK(clk), .RST(1'b0), .Q(
        round_reg[112]) );
  DFF \round_reg_reg[113]  ( .D(N125), .CLK(clk), .RST(1'b0), .Q(
        round_reg[113]) );
  DFF \round_reg_reg[114]  ( .D(N126), .CLK(clk), .RST(1'b0), .Q(
        round_reg[114]) );
  DFF \round_reg_reg[115]  ( .D(N127), .CLK(clk), .RST(1'b0), .Q(
        round_reg[115]) );
  DFF \round_reg_reg[116]  ( .D(N128), .CLK(clk), .RST(1'b0), .Q(
        round_reg[116]) );
  DFF \round_reg_reg[117]  ( .D(N129), .CLK(clk), .RST(1'b0), .Q(
        round_reg[117]) );
  DFF \round_reg_reg[118]  ( .D(N130), .CLK(clk), .RST(1'b0), .Q(
        round_reg[118]) );
  DFF \round_reg_reg[119]  ( .D(N131), .CLK(clk), .RST(1'b0), .Q(
        round_reg[119]) );
  DFF \round_reg_reg[120]  ( .D(N132), .CLK(clk), .RST(1'b0), .Q(
        round_reg[120]) );
  DFF \round_reg_reg[121]  ( .D(N133), .CLK(clk), .RST(1'b0), .Q(
        round_reg[121]) );
  DFF \round_reg_reg[122]  ( .D(N134), .CLK(clk), .RST(1'b0), .Q(
        round_reg[122]) );
  DFF \round_reg_reg[123]  ( .D(N135), .CLK(clk), .RST(1'b0), .Q(
        round_reg[123]) );
  DFF \round_reg_reg[124]  ( .D(N136), .CLK(clk), .RST(1'b0), .Q(
        round_reg[124]) );
  DFF \round_reg_reg[125]  ( .D(N137), .CLK(clk), .RST(1'b0), .Q(
        round_reg[125]) );
  DFF \round_reg_reg[126]  ( .D(N138), .CLK(clk), .RST(1'b0), .Q(
        round_reg[126]) );
  DFF \round_reg_reg[127]  ( .D(N139), .CLK(clk), .RST(1'b0), .Q(
        round_reg[127]) );
  DFF \round_reg_reg[128]  ( .D(N140), .CLK(clk), .RST(1'b0), .Q(
        round_reg[128]) );
  DFF \round_reg_reg[129]  ( .D(N141), .CLK(clk), .RST(1'b0), .Q(
        round_reg[129]) );
  DFF \round_reg_reg[130]  ( .D(N142), .CLK(clk), .RST(1'b0), .Q(
        round_reg[130]) );
  DFF \round_reg_reg[131]  ( .D(N143), .CLK(clk), .RST(1'b0), .Q(
        round_reg[131]) );
  DFF \round_reg_reg[132]  ( .D(N144), .CLK(clk), .RST(1'b0), .Q(
        round_reg[132]) );
  DFF \round_reg_reg[133]  ( .D(N145), .CLK(clk), .RST(1'b0), .Q(
        round_reg[133]) );
  DFF \round_reg_reg[134]  ( .D(N146), .CLK(clk), .RST(1'b0), .Q(
        round_reg[134]) );
  DFF \round_reg_reg[135]  ( .D(N147), .CLK(clk), .RST(1'b0), .Q(
        round_reg[135]) );
  DFF \round_reg_reg[136]  ( .D(N148), .CLK(clk), .RST(1'b0), .Q(
        round_reg[136]) );
  DFF \round_reg_reg[137]  ( .D(N149), .CLK(clk), .RST(1'b0), .Q(
        round_reg[137]) );
  DFF \round_reg_reg[138]  ( .D(N150), .CLK(clk), .RST(1'b0), .Q(
        round_reg[138]) );
  DFF \round_reg_reg[139]  ( .D(N151), .CLK(clk), .RST(1'b0), .Q(
        round_reg[139]) );
  DFF \round_reg_reg[140]  ( .D(N152), .CLK(clk), .RST(1'b0), .Q(
        round_reg[140]) );
  DFF \round_reg_reg[141]  ( .D(N153), .CLK(clk), .RST(1'b0), .Q(
        round_reg[141]) );
  DFF \round_reg_reg[142]  ( .D(N154), .CLK(clk), .RST(1'b0), .Q(
        round_reg[142]) );
  DFF \round_reg_reg[143]  ( .D(N155), .CLK(clk), .RST(1'b0), .Q(
        round_reg[143]) );
  DFF \round_reg_reg[144]  ( .D(N156), .CLK(clk), .RST(1'b0), .Q(
        round_reg[144]) );
  DFF \round_reg_reg[145]  ( .D(N157), .CLK(clk), .RST(1'b0), .Q(
        round_reg[145]) );
  DFF \round_reg_reg[146]  ( .D(N158), .CLK(clk), .RST(1'b0), .Q(
        round_reg[146]) );
  DFF \round_reg_reg[147]  ( .D(N159), .CLK(clk), .RST(1'b0), .Q(
        round_reg[147]) );
  DFF \round_reg_reg[148]  ( .D(N160), .CLK(clk), .RST(1'b0), .Q(
        round_reg[148]) );
  DFF \round_reg_reg[149]  ( .D(N161), .CLK(clk), .RST(1'b0), .Q(
        round_reg[149]) );
  DFF \round_reg_reg[150]  ( .D(N162), .CLK(clk), .RST(1'b0), .Q(
        round_reg[150]) );
  DFF \round_reg_reg[151]  ( .D(N163), .CLK(clk), .RST(1'b0), .Q(
        round_reg[151]) );
  DFF \round_reg_reg[152]  ( .D(N164), .CLK(clk), .RST(1'b0), .Q(
        round_reg[152]) );
  DFF \round_reg_reg[153]  ( .D(N165), .CLK(clk), .RST(1'b0), .Q(
        round_reg[153]) );
  DFF \round_reg_reg[154]  ( .D(N166), .CLK(clk), .RST(1'b0), .Q(
        round_reg[154]) );
  DFF \round_reg_reg[155]  ( .D(N167), .CLK(clk), .RST(1'b0), .Q(
        round_reg[155]) );
  DFF \round_reg_reg[156]  ( .D(N168), .CLK(clk), .RST(1'b0), .Q(
        round_reg[156]) );
  DFF \round_reg_reg[157]  ( .D(N169), .CLK(clk), .RST(1'b0), .Q(
        round_reg[157]) );
  DFF \round_reg_reg[158]  ( .D(N170), .CLK(clk), .RST(1'b0), .Q(
        round_reg[158]) );
  DFF \round_reg_reg[159]  ( .D(N171), .CLK(clk), .RST(1'b0), .Q(
        round_reg[159]) );
  DFF \round_reg_reg[160]  ( .D(N172), .CLK(clk), .RST(1'b0), .Q(
        round_reg[160]) );
  DFF \round_reg_reg[161]  ( .D(N173), .CLK(clk), .RST(1'b0), .Q(
        round_reg[161]) );
  DFF \round_reg_reg[162]  ( .D(N174), .CLK(clk), .RST(1'b0), .Q(
        round_reg[162]) );
  DFF \round_reg_reg[163]  ( .D(N175), .CLK(clk), .RST(1'b0), .Q(
        round_reg[163]) );
  DFF \round_reg_reg[164]  ( .D(N176), .CLK(clk), .RST(1'b0), .Q(
        round_reg[164]) );
  DFF \round_reg_reg[165]  ( .D(N177), .CLK(clk), .RST(1'b0), .Q(
        round_reg[165]) );
  DFF \round_reg_reg[166]  ( .D(N178), .CLK(clk), .RST(1'b0), .Q(
        round_reg[166]) );
  DFF \round_reg_reg[167]  ( .D(N179), .CLK(clk), .RST(1'b0), .Q(
        round_reg[167]) );
  DFF \round_reg_reg[168]  ( .D(N180), .CLK(clk), .RST(1'b0), .Q(
        round_reg[168]) );
  DFF \round_reg_reg[169]  ( .D(N181), .CLK(clk), .RST(1'b0), .Q(
        round_reg[169]) );
  DFF \round_reg_reg[170]  ( .D(N182), .CLK(clk), .RST(1'b0), .Q(
        round_reg[170]) );
  DFF \round_reg_reg[171]  ( .D(N183), .CLK(clk), .RST(1'b0), .Q(
        round_reg[171]) );
  DFF \round_reg_reg[172]  ( .D(N184), .CLK(clk), .RST(1'b0), .Q(
        round_reg[172]) );
  DFF \round_reg_reg[173]  ( .D(N185), .CLK(clk), .RST(1'b0), .Q(
        round_reg[173]) );
  DFF \round_reg_reg[174]  ( .D(N186), .CLK(clk), .RST(1'b0), .Q(
        round_reg[174]) );
  DFF \round_reg_reg[175]  ( .D(N187), .CLK(clk), .RST(1'b0), .Q(
        round_reg[175]) );
  DFF \round_reg_reg[176]  ( .D(N188), .CLK(clk), .RST(1'b0), .Q(
        round_reg[176]) );
  DFF \round_reg_reg[177]  ( .D(N189), .CLK(clk), .RST(1'b0), .Q(
        round_reg[177]) );
  DFF \round_reg_reg[178]  ( .D(N190), .CLK(clk), .RST(1'b0), .Q(
        round_reg[178]) );
  DFF \round_reg_reg[179]  ( .D(N191), .CLK(clk), .RST(1'b0), .Q(
        round_reg[179]) );
  DFF \round_reg_reg[180]  ( .D(N192), .CLK(clk), .RST(1'b0), .Q(
        round_reg[180]) );
  DFF \round_reg_reg[181]  ( .D(N193), .CLK(clk), .RST(1'b0), .Q(
        round_reg[181]) );
  DFF \round_reg_reg[182]  ( .D(N194), .CLK(clk), .RST(1'b0), .Q(
        round_reg[182]) );
  DFF \round_reg_reg[183]  ( .D(N195), .CLK(clk), .RST(1'b0), .Q(
        round_reg[183]) );
  DFF \round_reg_reg[184]  ( .D(N196), .CLK(clk), .RST(1'b0), .Q(
        round_reg[184]) );
  DFF \round_reg_reg[185]  ( .D(N197), .CLK(clk), .RST(1'b0), .Q(
        round_reg[185]) );
  DFF \round_reg_reg[186]  ( .D(N198), .CLK(clk), .RST(1'b0), .Q(
        round_reg[186]) );
  DFF \round_reg_reg[187]  ( .D(N199), .CLK(clk), .RST(1'b0), .Q(
        round_reg[187]) );
  DFF \round_reg_reg[188]  ( .D(N200), .CLK(clk), .RST(1'b0), .Q(
        round_reg[188]) );
  DFF \round_reg_reg[189]  ( .D(N201), .CLK(clk), .RST(1'b0), .Q(
        round_reg[189]) );
  DFF \round_reg_reg[190]  ( .D(N202), .CLK(clk), .RST(1'b0), .Q(
        round_reg[190]) );
  DFF \round_reg_reg[191]  ( .D(N203), .CLK(clk), .RST(1'b0), .Q(
        round_reg[191]) );
  DFF \round_reg_reg[192]  ( .D(N204), .CLK(clk), .RST(1'b0), .Q(
        round_reg[192]) );
  DFF \round_reg_reg[193]  ( .D(N205), .CLK(clk), .RST(1'b0), .Q(
        round_reg[193]) );
  DFF \round_reg_reg[194]  ( .D(N206), .CLK(clk), .RST(1'b0), .Q(
        round_reg[194]) );
  DFF \round_reg_reg[195]  ( .D(N207), .CLK(clk), .RST(1'b0), .Q(
        round_reg[195]) );
  DFF \round_reg_reg[196]  ( .D(N208), .CLK(clk), .RST(1'b0), .Q(
        round_reg[196]) );
  DFF \round_reg_reg[197]  ( .D(N209), .CLK(clk), .RST(1'b0), .Q(
        round_reg[197]) );
  DFF \round_reg_reg[198]  ( .D(N210), .CLK(clk), .RST(1'b0), .Q(
        round_reg[198]) );
  DFF \round_reg_reg[199]  ( .D(N211), .CLK(clk), .RST(1'b0), .Q(
        round_reg[199]) );
  DFF \round_reg_reg[200]  ( .D(N212), .CLK(clk), .RST(1'b0), .Q(
        round_reg[200]) );
  DFF \round_reg_reg[201]  ( .D(N213), .CLK(clk), .RST(1'b0), .Q(
        round_reg[201]) );
  DFF \round_reg_reg[202]  ( .D(N214), .CLK(clk), .RST(1'b0), .Q(
        round_reg[202]) );
  DFF \round_reg_reg[203]  ( .D(N215), .CLK(clk), .RST(1'b0), .Q(
        round_reg[203]) );
  DFF \round_reg_reg[204]  ( .D(N216), .CLK(clk), .RST(1'b0), .Q(
        round_reg[204]) );
  DFF \round_reg_reg[205]  ( .D(N217), .CLK(clk), .RST(1'b0), .Q(
        round_reg[205]) );
  DFF \round_reg_reg[206]  ( .D(N218), .CLK(clk), .RST(1'b0), .Q(
        round_reg[206]) );
  DFF \round_reg_reg[207]  ( .D(N219), .CLK(clk), .RST(1'b0), .Q(
        round_reg[207]) );
  DFF \round_reg_reg[208]  ( .D(N220), .CLK(clk), .RST(1'b0), .Q(
        round_reg[208]) );
  DFF \round_reg_reg[209]  ( .D(N221), .CLK(clk), .RST(1'b0), .Q(
        round_reg[209]) );
  DFF \round_reg_reg[210]  ( .D(N222), .CLK(clk), .RST(1'b0), .Q(
        round_reg[210]) );
  DFF \round_reg_reg[211]  ( .D(N223), .CLK(clk), .RST(1'b0), .Q(
        round_reg[211]) );
  DFF \round_reg_reg[212]  ( .D(N224), .CLK(clk), .RST(1'b0), .Q(
        round_reg[212]) );
  DFF \round_reg_reg[213]  ( .D(N225), .CLK(clk), .RST(1'b0), .Q(
        round_reg[213]) );
  DFF \round_reg_reg[214]  ( .D(N226), .CLK(clk), .RST(1'b0), .Q(
        round_reg[214]) );
  DFF \round_reg_reg[215]  ( .D(N227), .CLK(clk), .RST(1'b0), .Q(
        round_reg[215]) );
  DFF \round_reg_reg[216]  ( .D(N228), .CLK(clk), .RST(1'b0), .Q(
        round_reg[216]) );
  DFF \round_reg_reg[217]  ( .D(N229), .CLK(clk), .RST(1'b0), .Q(
        round_reg[217]) );
  DFF \round_reg_reg[218]  ( .D(N230), .CLK(clk), .RST(1'b0), .Q(
        round_reg[218]) );
  DFF \round_reg_reg[219]  ( .D(N231), .CLK(clk), .RST(1'b0), .Q(
        round_reg[219]) );
  DFF \round_reg_reg[220]  ( .D(N232), .CLK(clk), .RST(1'b0), .Q(
        round_reg[220]) );
  DFF \round_reg_reg[221]  ( .D(N233), .CLK(clk), .RST(1'b0), .Q(
        round_reg[221]) );
  DFF \round_reg_reg[222]  ( .D(N234), .CLK(clk), .RST(1'b0), .Q(
        round_reg[222]) );
  DFF \round_reg_reg[223]  ( .D(N235), .CLK(clk), .RST(1'b0), .Q(
        round_reg[223]) );
  DFF \round_reg_reg[224]  ( .D(N236), .CLK(clk), .RST(1'b0), .Q(
        round_reg[224]) );
  DFF \round_reg_reg[225]  ( .D(N237), .CLK(clk), .RST(1'b0), .Q(
        round_reg[225]) );
  DFF \round_reg_reg[226]  ( .D(N238), .CLK(clk), .RST(1'b0), .Q(
        round_reg[226]) );
  DFF \round_reg_reg[227]  ( .D(N239), .CLK(clk), .RST(1'b0), .Q(
        round_reg[227]) );
  DFF \round_reg_reg[228]  ( .D(N240), .CLK(clk), .RST(1'b0), .Q(
        round_reg[228]) );
  DFF \round_reg_reg[229]  ( .D(N241), .CLK(clk), .RST(1'b0), .Q(
        round_reg[229]) );
  DFF \round_reg_reg[230]  ( .D(N242), .CLK(clk), .RST(1'b0), .Q(
        round_reg[230]) );
  DFF \round_reg_reg[231]  ( .D(N243), .CLK(clk), .RST(1'b0), .Q(
        round_reg[231]) );
  DFF \round_reg_reg[232]  ( .D(N244), .CLK(clk), .RST(1'b0), .Q(
        round_reg[232]) );
  DFF \round_reg_reg[233]  ( .D(N245), .CLK(clk), .RST(1'b0), .Q(
        round_reg[233]) );
  DFF \round_reg_reg[234]  ( .D(N246), .CLK(clk), .RST(1'b0), .Q(
        round_reg[234]) );
  DFF \round_reg_reg[235]  ( .D(N247), .CLK(clk), .RST(1'b0), .Q(
        round_reg[235]) );
  DFF \round_reg_reg[236]  ( .D(N248), .CLK(clk), .RST(1'b0), .Q(
        round_reg[236]) );
  DFF \round_reg_reg[237]  ( .D(N249), .CLK(clk), .RST(1'b0), .Q(
        round_reg[237]) );
  DFF \round_reg_reg[238]  ( .D(N250), .CLK(clk), .RST(1'b0), .Q(
        round_reg[238]) );
  DFF \round_reg_reg[239]  ( .D(N251), .CLK(clk), .RST(1'b0), .Q(
        round_reg[239]) );
  DFF \round_reg_reg[240]  ( .D(N252), .CLK(clk), .RST(1'b0), .Q(
        round_reg[240]) );
  DFF \round_reg_reg[241]  ( .D(N253), .CLK(clk), .RST(1'b0), .Q(
        round_reg[241]) );
  DFF \round_reg_reg[242]  ( .D(N254), .CLK(clk), .RST(1'b0), .Q(
        round_reg[242]) );
  DFF \round_reg_reg[243]  ( .D(N255), .CLK(clk), .RST(1'b0), .Q(
        round_reg[243]) );
  DFF \round_reg_reg[244]  ( .D(N256), .CLK(clk), .RST(1'b0), .Q(
        round_reg[244]) );
  DFF \round_reg_reg[245]  ( .D(N257), .CLK(clk), .RST(1'b0), .Q(
        round_reg[245]) );
  DFF \round_reg_reg[246]  ( .D(N258), .CLK(clk), .RST(1'b0), .Q(
        round_reg[246]) );
  DFF \round_reg_reg[247]  ( .D(N259), .CLK(clk), .RST(1'b0), .Q(
        round_reg[247]) );
  DFF \round_reg_reg[248]  ( .D(N260), .CLK(clk), .RST(1'b0), .Q(
        round_reg[248]) );
  DFF \round_reg_reg[249]  ( .D(N261), .CLK(clk), .RST(1'b0), .Q(
        round_reg[249]) );
  DFF \round_reg_reg[250]  ( .D(N262), .CLK(clk), .RST(1'b0), .Q(
        round_reg[250]) );
  DFF \round_reg_reg[251]  ( .D(N263), .CLK(clk), .RST(1'b0), .Q(
        round_reg[251]) );
  DFF \round_reg_reg[252]  ( .D(N264), .CLK(clk), .RST(1'b0), .Q(
        round_reg[252]) );
  DFF \round_reg_reg[253]  ( .D(N265), .CLK(clk), .RST(1'b0), .Q(
        round_reg[253]) );
  DFF \round_reg_reg[254]  ( .D(N266), .CLK(clk), .RST(1'b0), .Q(
        round_reg[254]) );
  DFF \round_reg_reg[255]  ( .D(N267), .CLK(clk), .RST(1'b0), .Q(
        round_reg[255]) );
  DFF \round_reg_reg[256]  ( .D(N268), .CLK(clk), .RST(1'b0), .Q(
        round_reg[256]) );
  DFF \round_reg_reg[257]  ( .D(N269), .CLK(clk), .RST(1'b0), .Q(
        round_reg[257]) );
  DFF \round_reg_reg[258]  ( .D(N270), .CLK(clk), .RST(1'b0), .Q(
        round_reg[258]) );
  DFF \round_reg_reg[259]  ( .D(N271), .CLK(clk), .RST(1'b0), .Q(
        round_reg[259]) );
  DFF \round_reg_reg[260]  ( .D(N272), .CLK(clk), .RST(1'b0), .Q(
        round_reg[260]) );
  DFF \round_reg_reg[261]  ( .D(N273), .CLK(clk), .RST(1'b0), .Q(
        round_reg[261]) );
  DFF \round_reg_reg[262]  ( .D(N274), .CLK(clk), .RST(1'b0), .Q(
        round_reg[262]) );
  DFF \round_reg_reg[263]  ( .D(N275), .CLK(clk), .RST(1'b0), .Q(
        round_reg[263]) );
  DFF \round_reg_reg[264]  ( .D(N276), .CLK(clk), .RST(1'b0), .Q(
        round_reg[264]) );
  DFF \round_reg_reg[265]  ( .D(N277), .CLK(clk), .RST(1'b0), .Q(
        round_reg[265]) );
  DFF \round_reg_reg[266]  ( .D(N278), .CLK(clk), .RST(1'b0), .Q(
        round_reg[266]) );
  DFF \round_reg_reg[267]  ( .D(N279), .CLK(clk), .RST(1'b0), .Q(
        round_reg[267]) );
  DFF \round_reg_reg[268]  ( .D(N280), .CLK(clk), .RST(1'b0), .Q(
        round_reg[268]) );
  DFF \round_reg_reg[269]  ( .D(N281), .CLK(clk), .RST(1'b0), .Q(
        round_reg[269]) );
  DFF \round_reg_reg[270]  ( .D(N282), .CLK(clk), .RST(1'b0), .Q(
        round_reg[270]) );
  DFF \round_reg_reg[271]  ( .D(N283), .CLK(clk), .RST(1'b0), .Q(
        round_reg[271]) );
  DFF \round_reg_reg[272]  ( .D(N284), .CLK(clk), .RST(1'b0), .Q(
        round_reg[272]) );
  DFF \round_reg_reg[273]  ( .D(N285), .CLK(clk), .RST(1'b0), .Q(
        round_reg[273]) );
  DFF \round_reg_reg[274]  ( .D(N286), .CLK(clk), .RST(1'b0), .Q(
        round_reg[274]) );
  DFF \round_reg_reg[275]  ( .D(N287), .CLK(clk), .RST(1'b0), .Q(
        round_reg[275]) );
  DFF \round_reg_reg[276]  ( .D(N288), .CLK(clk), .RST(1'b0), .Q(
        round_reg[276]) );
  DFF \round_reg_reg[277]  ( .D(N289), .CLK(clk), .RST(1'b0), .Q(
        round_reg[277]) );
  DFF \round_reg_reg[278]  ( .D(N290), .CLK(clk), .RST(1'b0), .Q(
        round_reg[278]) );
  DFF \round_reg_reg[279]  ( .D(N291), .CLK(clk), .RST(1'b0), .Q(
        round_reg[279]) );
  DFF \round_reg_reg[280]  ( .D(N292), .CLK(clk), .RST(1'b0), .Q(
        round_reg[280]) );
  DFF \round_reg_reg[281]  ( .D(N293), .CLK(clk), .RST(1'b0), .Q(
        round_reg[281]) );
  DFF \round_reg_reg[282]  ( .D(N294), .CLK(clk), .RST(1'b0), .Q(
        round_reg[282]) );
  DFF \round_reg_reg[283]  ( .D(N295), .CLK(clk), .RST(1'b0), .Q(
        round_reg[283]) );
  DFF \round_reg_reg[284]  ( .D(N296), .CLK(clk), .RST(1'b0), .Q(
        round_reg[284]) );
  DFF \round_reg_reg[285]  ( .D(N297), .CLK(clk), .RST(1'b0), .Q(
        round_reg[285]) );
  DFF \round_reg_reg[286]  ( .D(N298), .CLK(clk), .RST(1'b0), .Q(
        round_reg[286]) );
  DFF \round_reg_reg[287]  ( .D(N299), .CLK(clk), .RST(1'b0), .Q(
        round_reg[287]) );
  DFF \round_reg_reg[288]  ( .D(N300), .CLK(clk), .RST(1'b0), .Q(
        round_reg[288]) );
  DFF \round_reg_reg[289]  ( .D(N301), .CLK(clk), .RST(1'b0), .Q(
        round_reg[289]) );
  DFF \round_reg_reg[290]  ( .D(N302), .CLK(clk), .RST(1'b0), .Q(
        round_reg[290]) );
  DFF \round_reg_reg[291]  ( .D(N303), .CLK(clk), .RST(1'b0), .Q(
        round_reg[291]) );
  DFF \round_reg_reg[292]  ( .D(N304), .CLK(clk), .RST(1'b0), .Q(
        round_reg[292]) );
  DFF \round_reg_reg[293]  ( .D(N305), .CLK(clk), .RST(1'b0), .Q(
        round_reg[293]) );
  DFF \round_reg_reg[294]  ( .D(N306), .CLK(clk), .RST(1'b0), .Q(
        round_reg[294]) );
  DFF \round_reg_reg[295]  ( .D(N307), .CLK(clk), .RST(1'b0), .Q(
        round_reg[295]) );
  DFF \round_reg_reg[296]  ( .D(N308), .CLK(clk), .RST(1'b0), .Q(
        round_reg[296]) );
  DFF \round_reg_reg[297]  ( .D(N309), .CLK(clk), .RST(1'b0), .Q(
        round_reg[297]) );
  DFF \round_reg_reg[298]  ( .D(N310), .CLK(clk), .RST(1'b0), .Q(
        round_reg[298]) );
  DFF \round_reg_reg[299]  ( .D(N311), .CLK(clk), .RST(1'b0), .Q(
        round_reg[299]) );
  DFF \round_reg_reg[300]  ( .D(N312), .CLK(clk), .RST(1'b0), .Q(
        round_reg[300]) );
  DFF \round_reg_reg[301]  ( .D(N313), .CLK(clk), .RST(1'b0), .Q(
        round_reg[301]) );
  DFF \round_reg_reg[302]  ( .D(N314), .CLK(clk), .RST(1'b0), .Q(
        round_reg[302]) );
  DFF \round_reg_reg[303]  ( .D(N315), .CLK(clk), .RST(1'b0), .Q(
        round_reg[303]) );
  DFF \round_reg_reg[304]  ( .D(N316), .CLK(clk), .RST(1'b0), .Q(
        round_reg[304]) );
  DFF \round_reg_reg[305]  ( .D(N317), .CLK(clk), .RST(1'b0), .Q(
        round_reg[305]) );
  DFF \round_reg_reg[306]  ( .D(N318), .CLK(clk), .RST(1'b0), .Q(
        round_reg[306]) );
  DFF \round_reg_reg[307]  ( .D(N319), .CLK(clk), .RST(1'b0), .Q(
        round_reg[307]) );
  DFF \round_reg_reg[308]  ( .D(N320), .CLK(clk), .RST(1'b0), .Q(
        round_reg[308]) );
  DFF \round_reg_reg[309]  ( .D(N321), .CLK(clk), .RST(1'b0), .Q(
        round_reg[309]) );
  DFF \round_reg_reg[310]  ( .D(N322), .CLK(clk), .RST(1'b0), .Q(
        round_reg[310]) );
  DFF \round_reg_reg[311]  ( .D(N323), .CLK(clk), .RST(1'b0), .Q(
        round_reg[311]) );
  DFF \round_reg_reg[312]  ( .D(N324), .CLK(clk), .RST(1'b0), .Q(
        round_reg[312]) );
  DFF \round_reg_reg[313]  ( .D(N325), .CLK(clk), .RST(1'b0), .Q(
        round_reg[313]) );
  DFF \round_reg_reg[314]  ( .D(N326), .CLK(clk), .RST(1'b0), .Q(
        round_reg[314]) );
  DFF \round_reg_reg[315]  ( .D(N327), .CLK(clk), .RST(1'b0), .Q(
        round_reg[315]) );
  DFF \round_reg_reg[316]  ( .D(N328), .CLK(clk), .RST(1'b0), .Q(
        round_reg[316]) );
  DFF \round_reg_reg[317]  ( .D(N329), .CLK(clk), .RST(1'b0), .Q(
        round_reg[317]) );
  DFF \round_reg_reg[318]  ( .D(N330), .CLK(clk), .RST(1'b0), .Q(
        round_reg[318]) );
  DFF \round_reg_reg[319]  ( .D(N331), .CLK(clk), .RST(1'b0), .Q(
        round_reg[319]) );
  DFF \round_reg_reg[320]  ( .D(N332), .CLK(clk), .RST(1'b0), .Q(
        round_reg[320]) );
  DFF \round_reg_reg[321]  ( .D(N333), .CLK(clk), .RST(1'b0), .Q(
        round_reg[321]) );
  DFF \round_reg_reg[322]  ( .D(N334), .CLK(clk), .RST(1'b0), .Q(
        round_reg[322]) );
  DFF \round_reg_reg[323]  ( .D(N335), .CLK(clk), .RST(1'b0), .Q(
        round_reg[323]) );
  DFF \round_reg_reg[324]  ( .D(N336), .CLK(clk), .RST(1'b0), .Q(
        round_reg[324]) );
  DFF \round_reg_reg[325]  ( .D(N337), .CLK(clk), .RST(1'b0), .Q(
        round_reg[325]) );
  DFF \round_reg_reg[326]  ( .D(N338), .CLK(clk), .RST(1'b0), .Q(
        round_reg[326]) );
  DFF \round_reg_reg[327]  ( .D(N339), .CLK(clk), .RST(1'b0), .Q(
        round_reg[327]) );
  DFF \round_reg_reg[328]  ( .D(N340), .CLK(clk), .RST(1'b0), .Q(
        round_reg[328]) );
  DFF \round_reg_reg[329]  ( .D(N341), .CLK(clk), .RST(1'b0), .Q(
        round_reg[329]) );
  DFF \round_reg_reg[330]  ( .D(N342), .CLK(clk), .RST(1'b0), .Q(
        round_reg[330]) );
  DFF \round_reg_reg[331]  ( .D(N343), .CLK(clk), .RST(1'b0), .Q(
        round_reg[331]) );
  DFF \round_reg_reg[332]  ( .D(N344), .CLK(clk), .RST(1'b0), .Q(
        round_reg[332]) );
  DFF \round_reg_reg[333]  ( .D(N345), .CLK(clk), .RST(1'b0), .Q(
        round_reg[333]) );
  DFF \round_reg_reg[334]  ( .D(N346), .CLK(clk), .RST(1'b0), .Q(
        round_reg[334]) );
  DFF \round_reg_reg[335]  ( .D(N347), .CLK(clk), .RST(1'b0), .Q(
        round_reg[335]) );
  DFF \round_reg_reg[336]  ( .D(N348), .CLK(clk), .RST(1'b0), .Q(
        round_reg[336]) );
  DFF \round_reg_reg[337]  ( .D(N349), .CLK(clk), .RST(1'b0), .Q(
        round_reg[337]) );
  DFF \round_reg_reg[338]  ( .D(N350), .CLK(clk), .RST(1'b0), .Q(
        round_reg[338]) );
  DFF \round_reg_reg[339]  ( .D(N351), .CLK(clk), .RST(1'b0), .Q(
        round_reg[339]) );
  DFF \round_reg_reg[340]  ( .D(N352), .CLK(clk), .RST(1'b0), .Q(
        round_reg[340]) );
  DFF \round_reg_reg[341]  ( .D(N353), .CLK(clk), .RST(1'b0), .Q(
        round_reg[341]) );
  DFF \round_reg_reg[342]  ( .D(N354), .CLK(clk), .RST(1'b0), .Q(
        round_reg[342]) );
  DFF \round_reg_reg[343]  ( .D(N355), .CLK(clk), .RST(1'b0), .Q(
        round_reg[343]) );
  DFF \round_reg_reg[344]  ( .D(N356), .CLK(clk), .RST(1'b0), .Q(
        round_reg[344]) );
  DFF \round_reg_reg[345]  ( .D(N357), .CLK(clk), .RST(1'b0), .Q(
        round_reg[345]) );
  DFF \round_reg_reg[346]  ( .D(N358), .CLK(clk), .RST(1'b0), .Q(
        round_reg[346]) );
  DFF \round_reg_reg[347]  ( .D(N359), .CLK(clk), .RST(1'b0), .Q(
        round_reg[347]) );
  DFF \round_reg_reg[348]  ( .D(N360), .CLK(clk), .RST(1'b0), .Q(
        round_reg[348]) );
  DFF \round_reg_reg[349]  ( .D(N361), .CLK(clk), .RST(1'b0), .Q(
        round_reg[349]) );
  DFF \round_reg_reg[350]  ( .D(N362), .CLK(clk), .RST(1'b0), .Q(
        round_reg[350]) );
  DFF \round_reg_reg[351]  ( .D(N363), .CLK(clk), .RST(1'b0), .Q(
        round_reg[351]) );
  DFF \round_reg_reg[352]  ( .D(N364), .CLK(clk), .RST(1'b0), .Q(
        round_reg[352]) );
  DFF \round_reg_reg[353]  ( .D(N365), .CLK(clk), .RST(1'b0), .Q(
        round_reg[353]) );
  DFF \round_reg_reg[354]  ( .D(N366), .CLK(clk), .RST(1'b0), .Q(
        round_reg[354]) );
  DFF \round_reg_reg[355]  ( .D(N367), .CLK(clk), .RST(1'b0), .Q(
        round_reg[355]) );
  DFF \round_reg_reg[356]  ( .D(N368), .CLK(clk), .RST(1'b0), .Q(
        round_reg[356]) );
  DFF \round_reg_reg[357]  ( .D(N369), .CLK(clk), .RST(1'b0), .Q(
        round_reg[357]) );
  DFF \round_reg_reg[358]  ( .D(N370), .CLK(clk), .RST(1'b0), .Q(
        round_reg[358]) );
  DFF \round_reg_reg[359]  ( .D(N371), .CLK(clk), .RST(1'b0), .Q(
        round_reg[359]) );
  DFF \round_reg_reg[360]  ( .D(N372), .CLK(clk), .RST(1'b0), .Q(
        round_reg[360]) );
  DFF \round_reg_reg[361]  ( .D(N373), .CLK(clk), .RST(1'b0), .Q(
        round_reg[361]) );
  DFF \round_reg_reg[362]  ( .D(N374), .CLK(clk), .RST(1'b0), .Q(
        round_reg[362]) );
  DFF \round_reg_reg[363]  ( .D(N375), .CLK(clk), .RST(1'b0), .Q(
        round_reg[363]) );
  DFF \round_reg_reg[364]  ( .D(N376), .CLK(clk), .RST(1'b0), .Q(
        round_reg[364]) );
  DFF \round_reg_reg[365]  ( .D(N377), .CLK(clk), .RST(1'b0), .Q(
        round_reg[365]) );
  DFF \round_reg_reg[366]  ( .D(N378), .CLK(clk), .RST(1'b0), .Q(
        round_reg[366]) );
  DFF \round_reg_reg[367]  ( .D(N379), .CLK(clk), .RST(1'b0), .Q(
        round_reg[367]) );
  DFF \round_reg_reg[368]  ( .D(N380), .CLK(clk), .RST(1'b0), .Q(
        round_reg[368]) );
  DFF \round_reg_reg[369]  ( .D(N381), .CLK(clk), .RST(1'b0), .Q(
        round_reg[369]) );
  DFF \round_reg_reg[370]  ( .D(N382), .CLK(clk), .RST(1'b0), .Q(
        round_reg[370]) );
  DFF \round_reg_reg[371]  ( .D(N383), .CLK(clk), .RST(1'b0), .Q(
        round_reg[371]) );
  DFF \round_reg_reg[372]  ( .D(N384), .CLK(clk), .RST(1'b0), .Q(
        round_reg[372]) );
  DFF \round_reg_reg[373]  ( .D(N385), .CLK(clk), .RST(1'b0), .Q(
        round_reg[373]) );
  DFF \round_reg_reg[374]  ( .D(N386), .CLK(clk), .RST(1'b0), .Q(
        round_reg[374]) );
  DFF \round_reg_reg[375]  ( .D(N387), .CLK(clk), .RST(1'b0), .Q(
        round_reg[375]) );
  DFF \round_reg_reg[376]  ( .D(N388), .CLK(clk), .RST(1'b0), .Q(
        round_reg[376]) );
  DFF \round_reg_reg[377]  ( .D(N389), .CLK(clk), .RST(1'b0), .Q(
        round_reg[377]) );
  DFF \round_reg_reg[378]  ( .D(N390), .CLK(clk), .RST(1'b0), .Q(
        round_reg[378]) );
  DFF \round_reg_reg[379]  ( .D(N391), .CLK(clk), .RST(1'b0), .Q(
        round_reg[379]) );
  DFF \round_reg_reg[380]  ( .D(N392), .CLK(clk), .RST(1'b0), .Q(
        round_reg[380]) );
  DFF \round_reg_reg[381]  ( .D(N393), .CLK(clk), .RST(1'b0), .Q(
        round_reg[381]) );
  DFF \round_reg_reg[382]  ( .D(N394), .CLK(clk), .RST(1'b0), .Q(
        round_reg[382]) );
  DFF \round_reg_reg[383]  ( .D(N395), .CLK(clk), .RST(1'b0), .Q(
        round_reg[383]) );
  DFF \round_reg_reg[384]  ( .D(N396), .CLK(clk), .RST(1'b0), .Q(
        round_reg[384]) );
  DFF \round_reg_reg[385]  ( .D(N397), .CLK(clk), .RST(1'b0), .Q(
        round_reg[385]) );
  DFF \round_reg_reg[386]  ( .D(N398), .CLK(clk), .RST(1'b0), .Q(
        round_reg[386]) );
  DFF \round_reg_reg[387]  ( .D(N399), .CLK(clk), .RST(1'b0), .Q(
        round_reg[387]) );
  DFF \round_reg_reg[388]  ( .D(N400), .CLK(clk), .RST(1'b0), .Q(
        round_reg[388]) );
  DFF \round_reg_reg[389]  ( .D(N401), .CLK(clk), .RST(1'b0), .Q(
        round_reg[389]) );
  DFF \round_reg_reg[390]  ( .D(N402), .CLK(clk), .RST(1'b0), .Q(
        round_reg[390]) );
  DFF \round_reg_reg[391]  ( .D(N403), .CLK(clk), .RST(1'b0), .Q(
        round_reg[391]) );
  DFF \round_reg_reg[392]  ( .D(N404), .CLK(clk), .RST(1'b0), .Q(
        round_reg[392]) );
  DFF \round_reg_reg[393]  ( .D(N405), .CLK(clk), .RST(1'b0), .Q(
        round_reg[393]) );
  DFF \round_reg_reg[394]  ( .D(N406), .CLK(clk), .RST(1'b0), .Q(
        round_reg[394]) );
  DFF \round_reg_reg[395]  ( .D(N407), .CLK(clk), .RST(1'b0), .Q(
        round_reg[395]) );
  DFF \round_reg_reg[396]  ( .D(N408), .CLK(clk), .RST(1'b0), .Q(
        round_reg[396]) );
  DFF \round_reg_reg[397]  ( .D(N409), .CLK(clk), .RST(1'b0), .Q(
        round_reg[397]) );
  DFF \round_reg_reg[398]  ( .D(N410), .CLK(clk), .RST(1'b0), .Q(
        round_reg[398]) );
  DFF \round_reg_reg[399]  ( .D(N411), .CLK(clk), .RST(1'b0), .Q(
        round_reg[399]) );
  DFF \round_reg_reg[400]  ( .D(N412), .CLK(clk), .RST(1'b0), .Q(
        round_reg[400]) );
  DFF \round_reg_reg[401]  ( .D(N413), .CLK(clk), .RST(1'b0), .Q(
        round_reg[401]) );
  DFF \round_reg_reg[402]  ( .D(N414), .CLK(clk), .RST(1'b0), .Q(
        round_reg[402]) );
  DFF \round_reg_reg[403]  ( .D(N415), .CLK(clk), .RST(1'b0), .Q(
        round_reg[403]) );
  DFF \round_reg_reg[404]  ( .D(N416), .CLK(clk), .RST(1'b0), .Q(
        round_reg[404]) );
  DFF \round_reg_reg[405]  ( .D(N417), .CLK(clk), .RST(1'b0), .Q(
        round_reg[405]) );
  DFF \round_reg_reg[406]  ( .D(N418), .CLK(clk), .RST(1'b0), .Q(
        round_reg[406]) );
  DFF \round_reg_reg[407]  ( .D(N419), .CLK(clk), .RST(1'b0), .Q(
        round_reg[407]) );
  DFF \round_reg_reg[408]  ( .D(N420), .CLK(clk), .RST(1'b0), .Q(
        round_reg[408]) );
  DFF \round_reg_reg[409]  ( .D(N421), .CLK(clk), .RST(1'b0), .Q(
        round_reg[409]) );
  DFF \round_reg_reg[410]  ( .D(N422), .CLK(clk), .RST(1'b0), .Q(
        round_reg[410]) );
  DFF \round_reg_reg[411]  ( .D(N423), .CLK(clk), .RST(1'b0), .Q(
        round_reg[411]) );
  DFF \round_reg_reg[412]  ( .D(N424), .CLK(clk), .RST(1'b0), .Q(
        round_reg[412]) );
  DFF \round_reg_reg[413]  ( .D(N425), .CLK(clk), .RST(1'b0), .Q(
        round_reg[413]) );
  DFF \round_reg_reg[414]  ( .D(N426), .CLK(clk), .RST(1'b0), .Q(
        round_reg[414]) );
  DFF \round_reg_reg[415]  ( .D(N427), .CLK(clk), .RST(1'b0), .Q(
        round_reg[415]) );
  DFF \round_reg_reg[416]  ( .D(N428), .CLK(clk), .RST(1'b0), .Q(
        round_reg[416]) );
  DFF \round_reg_reg[417]  ( .D(N429), .CLK(clk), .RST(1'b0), .Q(
        round_reg[417]) );
  DFF \round_reg_reg[418]  ( .D(N430), .CLK(clk), .RST(1'b0), .Q(
        round_reg[418]) );
  DFF \round_reg_reg[419]  ( .D(N431), .CLK(clk), .RST(1'b0), .Q(
        round_reg[419]) );
  DFF \round_reg_reg[420]  ( .D(N432), .CLK(clk), .RST(1'b0), .Q(
        round_reg[420]) );
  DFF \round_reg_reg[421]  ( .D(N433), .CLK(clk), .RST(1'b0), .Q(
        round_reg[421]) );
  DFF \round_reg_reg[422]  ( .D(N434), .CLK(clk), .RST(1'b0), .Q(
        round_reg[422]) );
  DFF \round_reg_reg[423]  ( .D(N435), .CLK(clk), .RST(1'b0), .Q(
        round_reg[423]) );
  DFF \round_reg_reg[424]  ( .D(N436), .CLK(clk), .RST(1'b0), .Q(
        round_reg[424]) );
  DFF \round_reg_reg[425]  ( .D(N437), .CLK(clk), .RST(1'b0), .Q(
        round_reg[425]) );
  DFF \round_reg_reg[426]  ( .D(N438), .CLK(clk), .RST(1'b0), .Q(
        round_reg[426]) );
  DFF \round_reg_reg[427]  ( .D(N439), .CLK(clk), .RST(1'b0), .Q(
        round_reg[427]) );
  DFF \round_reg_reg[428]  ( .D(N440), .CLK(clk), .RST(1'b0), .Q(
        round_reg[428]) );
  DFF \round_reg_reg[429]  ( .D(N441), .CLK(clk), .RST(1'b0), .Q(
        round_reg[429]) );
  DFF \round_reg_reg[430]  ( .D(N442), .CLK(clk), .RST(1'b0), .Q(
        round_reg[430]) );
  DFF \round_reg_reg[431]  ( .D(N443), .CLK(clk), .RST(1'b0), .Q(
        round_reg[431]) );
  DFF \round_reg_reg[432]  ( .D(N444), .CLK(clk), .RST(1'b0), .Q(
        round_reg[432]) );
  DFF \round_reg_reg[433]  ( .D(N445), .CLK(clk), .RST(1'b0), .Q(
        round_reg[433]) );
  DFF \round_reg_reg[434]  ( .D(N446), .CLK(clk), .RST(1'b0), .Q(
        round_reg[434]) );
  DFF \round_reg_reg[435]  ( .D(N447), .CLK(clk), .RST(1'b0), .Q(
        round_reg[435]) );
  DFF \round_reg_reg[436]  ( .D(N448), .CLK(clk), .RST(1'b0), .Q(
        round_reg[436]) );
  DFF \round_reg_reg[437]  ( .D(N449), .CLK(clk), .RST(1'b0), .Q(
        round_reg[437]) );
  DFF \round_reg_reg[438]  ( .D(N450), .CLK(clk), .RST(1'b0), .Q(
        round_reg[438]) );
  DFF \round_reg_reg[439]  ( .D(N451), .CLK(clk), .RST(1'b0), .Q(
        round_reg[439]) );
  DFF \round_reg_reg[440]  ( .D(N452), .CLK(clk), .RST(1'b0), .Q(
        round_reg[440]) );
  DFF \round_reg_reg[441]  ( .D(N453), .CLK(clk), .RST(1'b0), .Q(
        round_reg[441]) );
  DFF \round_reg_reg[442]  ( .D(N454), .CLK(clk), .RST(1'b0), .Q(
        round_reg[442]) );
  DFF \round_reg_reg[443]  ( .D(N455), .CLK(clk), .RST(1'b0), .Q(
        round_reg[443]) );
  DFF \round_reg_reg[444]  ( .D(N456), .CLK(clk), .RST(1'b0), .Q(
        round_reg[444]) );
  DFF \round_reg_reg[445]  ( .D(N457), .CLK(clk), .RST(1'b0), .Q(
        round_reg[445]) );
  DFF \round_reg_reg[446]  ( .D(N458), .CLK(clk), .RST(1'b0), .Q(
        round_reg[446]) );
  DFF \round_reg_reg[447]  ( .D(N459), .CLK(clk), .RST(1'b0), .Q(
        round_reg[447]) );
  DFF \round_reg_reg[448]  ( .D(N460), .CLK(clk), .RST(1'b0), .Q(
        round_reg[448]) );
  DFF \round_reg_reg[449]  ( .D(N461), .CLK(clk), .RST(1'b0), .Q(
        round_reg[449]) );
  DFF \round_reg_reg[450]  ( .D(N462), .CLK(clk), .RST(1'b0), .Q(
        round_reg[450]) );
  DFF \round_reg_reg[451]  ( .D(N463), .CLK(clk), .RST(1'b0), .Q(
        round_reg[451]) );
  DFF \round_reg_reg[452]  ( .D(N464), .CLK(clk), .RST(1'b0), .Q(
        round_reg[452]) );
  DFF \round_reg_reg[453]  ( .D(N465), .CLK(clk), .RST(1'b0), .Q(
        round_reg[453]) );
  DFF \round_reg_reg[454]  ( .D(N466), .CLK(clk), .RST(1'b0), .Q(
        round_reg[454]) );
  DFF \round_reg_reg[455]  ( .D(N467), .CLK(clk), .RST(1'b0), .Q(
        round_reg[455]) );
  DFF \round_reg_reg[456]  ( .D(N468), .CLK(clk), .RST(1'b0), .Q(
        round_reg[456]) );
  DFF \round_reg_reg[457]  ( .D(N469), .CLK(clk), .RST(1'b0), .Q(
        round_reg[457]) );
  DFF \round_reg_reg[458]  ( .D(N470), .CLK(clk), .RST(1'b0), .Q(
        round_reg[458]) );
  DFF \round_reg_reg[459]  ( .D(N471), .CLK(clk), .RST(1'b0), .Q(
        round_reg[459]) );
  DFF \round_reg_reg[460]  ( .D(N472), .CLK(clk), .RST(1'b0), .Q(
        round_reg[460]) );
  DFF \round_reg_reg[461]  ( .D(N473), .CLK(clk), .RST(1'b0), .Q(
        round_reg[461]) );
  DFF \round_reg_reg[462]  ( .D(N474), .CLK(clk), .RST(1'b0), .Q(
        round_reg[462]) );
  DFF \round_reg_reg[463]  ( .D(N475), .CLK(clk), .RST(1'b0), .Q(
        round_reg[463]) );
  DFF \round_reg_reg[464]  ( .D(N476), .CLK(clk), .RST(1'b0), .Q(
        round_reg[464]) );
  DFF \round_reg_reg[465]  ( .D(N477), .CLK(clk), .RST(1'b0), .Q(
        round_reg[465]) );
  DFF \round_reg_reg[466]  ( .D(N478), .CLK(clk), .RST(1'b0), .Q(
        round_reg[466]) );
  DFF \round_reg_reg[467]  ( .D(N479), .CLK(clk), .RST(1'b0), .Q(
        round_reg[467]) );
  DFF \round_reg_reg[468]  ( .D(N480), .CLK(clk), .RST(1'b0), .Q(
        round_reg[468]) );
  DFF \round_reg_reg[469]  ( .D(N481), .CLK(clk), .RST(1'b0), .Q(
        round_reg[469]) );
  DFF \round_reg_reg[470]  ( .D(N482), .CLK(clk), .RST(1'b0), .Q(
        round_reg[470]) );
  DFF \round_reg_reg[471]  ( .D(N483), .CLK(clk), .RST(1'b0), .Q(
        round_reg[471]) );
  DFF \round_reg_reg[472]  ( .D(N484), .CLK(clk), .RST(1'b0), .Q(
        round_reg[472]) );
  DFF \round_reg_reg[473]  ( .D(N485), .CLK(clk), .RST(1'b0), .Q(
        round_reg[473]) );
  DFF \round_reg_reg[474]  ( .D(N486), .CLK(clk), .RST(1'b0), .Q(
        round_reg[474]) );
  DFF \round_reg_reg[475]  ( .D(N487), .CLK(clk), .RST(1'b0), .Q(
        round_reg[475]) );
  DFF \round_reg_reg[476]  ( .D(N488), .CLK(clk), .RST(1'b0), .Q(
        round_reg[476]) );
  DFF \round_reg_reg[477]  ( .D(N489), .CLK(clk), .RST(1'b0), .Q(
        round_reg[477]) );
  DFF \round_reg_reg[478]  ( .D(N490), .CLK(clk), .RST(1'b0), .Q(
        round_reg[478]) );
  DFF \round_reg_reg[479]  ( .D(N491), .CLK(clk), .RST(1'b0), .Q(
        round_reg[479]) );
  DFF \round_reg_reg[480]  ( .D(N492), .CLK(clk), .RST(1'b0), .Q(
        round_reg[480]) );
  DFF \round_reg_reg[481]  ( .D(N493), .CLK(clk), .RST(1'b0), .Q(
        round_reg[481]) );
  DFF \round_reg_reg[482]  ( .D(N494), .CLK(clk), .RST(1'b0), .Q(
        round_reg[482]) );
  DFF \round_reg_reg[483]  ( .D(N495), .CLK(clk), .RST(1'b0), .Q(
        round_reg[483]) );
  DFF \round_reg_reg[484]  ( .D(N496), .CLK(clk), .RST(1'b0), .Q(
        round_reg[484]) );
  DFF \round_reg_reg[485]  ( .D(N497), .CLK(clk), .RST(1'b0), .Q(
        round_reg[485]) );
  DFF \round_reg_reg[486]  ( .D(N498), .CLK(clk), .RST(1'b0), .Q(
        round_reg[486]) );
  DFF \round_reg_reg[487]  ( .D(N499), .CLK(clk), .RST(1'b0), .Q(
        round_reg[487]) );
  DFF \round_reg_reg[488]  ( .D(N500), .CLK(clk), .RST(1'b0), .Q(
        round_reg[488]) );
  DFF \round_reg_reg[489]  ( .D(N501), .CLK(clk), .RST(1'b0), .Q(
        round_reg[489]) );
  DFF \round_reg_reg[490]  ( .D(N502), .CLK(clk), .RST(1'b0), .Q(
        round_reg[490]) );
  DFF \round_reg_reg[491]  ( .D(N503), .CLK(clk), .RST(1'b0), .Q(
        round_reg[491]) );
  DFF \round_reg_reg[492]  ( .D(N504), .CLK(clk), .RST(1'b0), .Q(
        round_reg[492]) );
  DFF \round_reg_reg[493]  ( .D(N505), .CLK(clk), .RST(1'b0), .Q(
        round_reg[493]) );
  DFF \round_reg_reg[494]  ( .D(N506), .CLK(clk), .RST(1'b0), .Q(
        round_reg[494]) );
  DFF \round_reg_reg[495]  ( .D(N507), .CLK(clk), .RST(1'b0), .Q(
        round_reg[495]) );
  DFF \round_reg_reg[496]  ( .D(N508), .CLK(clk), .RST(1'b0), .Q(
        round_reg[496]) );
  DFF \round_reg_reg[497]  ( .D(N509), .CLK(clk), .RST(1'b0), .Q(
        round_reg[497]) );
  DFF \round_reg_reg[498]  ( .D(N510), .CLK(clk), .RST(1'b0), .Q(
        round_reg[498]) );
  DFF \round_reg_reg[499]  ( .D(N511), .CLK(clk), .RST(1'b0), .Q(
        round_reg[499]) );
  DFF \round_reg_reg[500]  ( .D(N512), .CLK(clk), .RST(1'b0), .Q(
        round_reg[500]) );
  DFF \round_reg_reg[501]  ( .D(N513), .CLK(clk), .RST(1'b0), .Q(
        round_reg[501]) );
  DFF \round_reg_reg[502]  ( .D(N514), .CLK(clk), .RST(1'b0), .Q(
        round_reg[502]) );
  DFF \round_reg_reg[503]  ( .D(N515), .CLK(clk), .RST(1'b0), .Q(
        round_reg[503]) );
  DFF \round_reg_reg[504]  ( .D(N516), .CLK(clk), .RST(1'b0), .Q(
        round_reg[504]) );
  DFF \round_reg_reg[505]  ( .D(N517), .CLK(clk), .RST(1'b0), .Q(
        round_reg[505]) );
  DFF \round_reg_reg[506]  ( .D(N518), .CLK(clk), .RST(1'b0), .Q(
        round_reg[506]) );
  DFF \round_reg_reg[507]  ( .D(N519), .CLK(clk), .RST(1'b0), .Q(
        round_reg[507]) );
  DFF \round_reg_reg[508]  ( .D(N520), .CLK(clk), .RST(1'b0), .Q(
        round_reg[508]) );
  DFF \round_reg_reg[509]  ( .D(N521), .CLK(clk), .RST(1'b0), .Q(
        round_reg[509]) );
  DFF \round_reg_reg[510]  ( .D(N522), .CLK(clk), .RST(1'b0), .Q(
        round_reg[510]) );
  DFF \round_reg_reg[511]  ( .D(N523), .CLK(clk), .RST(1'b0), .Q(
        round_reg[511]) );
  DFF \round_reg_reg[512]  ( .D(N524), .CLK(clk), .RST(1'b0), .Q(
        round_reg[512]) );
  DFF \round_reg_reg[513]  ( .D(N525), .CLK(clk), .RST(1'b0), .Q(
        round_reg[513]) );
  DFF \round_reg_reg[514]  ( .D(N526), .CLK(clk), .RST(1'b0), .Q(
        round_reg[514]) );
  DFF \round_reg_reg[515]  ( .D(N527), .CLK(clk), .RST(1'b0), .Q(
        round_reg[515]) );
  DFF \round_reg_reg[516]  ( .D(N528), .CLK(clk), .RST(1'b0), .Q(
        round_reg[516]) );
  DFF \round_reg_reg[517]  ( .D(N529), .CLK(clk), .RST(1'b0), .Q(
        round_reg[517]) );
  DFF \round_reg_reg[518]  ( .D(N530), .CLK(clk), .RST(1'b0), .Q(
        round_reg[518]) );
  DFF \round_reg_reg[519]  ( .D(N531), .CLK(clk), .RST(1'b0), .Q(
        round_reg[519]) );
  DFF \round_reg_reg[520]  ( .D(N532), .CLK(clk), .RST(1'b0), .Q(
        round_reg[520]) );
  DFF \round_reg_reg[521]  ( .D(N533), .CLK(clk), .RST(1'b0), .Q(
        round_reg[521]) );
  DFF \round_reg_reg[522]  ( .D(N534), .CLK(clk), .RST(1'b0), .Q(
        round_reg[522]) );
  DFF \round_reg_reg[523]  ( .D(N535), .CLK(clk), .RST(1'b0), .Q(
        round_reg[523]) );
  DFF \round_reg_reg[524]  ( .D(N536), .CLK(clk), .RST(1'b0), .Q(
        round_reg[524]) );
  DFF \round_reg_reg[525]  ( .D(N537), .CLK(clk), .RST(1'b0), .Q(
        round_reg[525]) );
  DFF \round_reg_reg[526]  ( .D(N538), .CLK(clk), .RST(1'b0), .Q(
        round_reg[526]) );
  DFF \round_reg_reg[527]  ( .D(N539), .CLK(clk), .RST(1'b0), .Q(
        round_reg[527]) );
  DFF \round_reg_reg[528]  ( .D(N540), .CLK(clk), .RST(1'b0), .Q(
        round_reg[528]) );
  DFF \round_reg_reg[529]  ( .D(N541), .CLK(clk), .RST(1'b0), .Q(
        round_reg[529]) );
  DFF \round_reg_reg[530]  ( .D(N542), .CLK(clk), .RST(1'b0), .Q(
        round_reg[530]) );
  DFF \round_reg_reg[531]  ( .D(N543), .CLK(clk), .RST(1'b0), .Q(
        round_reg[531]) );
  DFF \round_reg_reg[532]  ( .D(N544), .CLK(clk), .RST(1'b0), .Q(
        round_reg[532]) );
  DFF \round_reg_reg[533]  ( .D(N545), .CLK(clk), .RST(1'b0), .Q(
        round_reg[533]) );
  DFF \round_reg_reg[534]  ( .D(N546), .CLK(clk), .RST(1'b0), .Q(
        round_reg[534]) );
  DFF \round_reg_reg[535]  ( .D(N547), .CLK(clk), .RST(1'b0), .Q(
        round_reg[535]) );
  DFF \round_reg_reg[536]  ( .D(N548), .CLK(clk), .RST(1'b0), .Q(
        round_reg[536]) );
  DFF \round_reg_reg[537]  ( .D(N549), .CLK(clk), .RST(1'b0), .Q(
        round_reg[537]) );
  DFF \round_reg_reg[538]  ( .D(N550), .CLK(clk), .RST(1'b0), .Q(
        round_reg[538]) );
  DFF \round_reg_reg[539]  ( .D(N551), .CLK(clk), .RST(1'b0), .Q(
        round_reg[539]) );
  DFF \round_reg_reg[540]  ( .D(N552), .CLK(clk), .RST(1'b0), .Q(
        round_reg[540]) );
  DFF \round_reg_reg[541]  ( .D(N553), .CLK(clk), .RST(1'b0), .Q(
        round_reg[541]) );
  DFF \round_reg_reg[542]  ( .D(N554), .CLK(clk), .RST(1'b0), .Q(
        round_reg[542]) );
  DFF \round_reg_reg[543]  ( .D(N555), .CLK(clk), .RST(1'b0), .Q(
        round_reg[543]) );
  DFF \round_reg_reg[544]  ( .D(N556), .CLK(clk), .RST(1'b0), .Q(
        round_reg[544]) );
  DFF \round_reg_reg[545]  ( .D(N557), .CLK(clk), .RST(1'b0), .Q(
        round_reg[545]) );
  DFF \round_reg_reg[546]  ( .D(N558), .CLK(clk), .RST(1'b0), .Q(
        round_reg[546]) );
  DFF \round_reg_reg[547]  ( .D(N559), .CLK(clk), .RST(1'b0), .Q(
        round_reg[547]) );
  DFF \round_reg_reg[548]  ( .D(N560), .CLK(clk), .RST(1'b0), .Q(
        round_reg[548]) );
  DFF \round_reg_reg[549]  ( .D(N561), .CLK(clk), .RST(1'b0), .Q(
        round_reg[549]) );
  DFF \round_reg_reg[550]  ( .D(N562), .CLK(clk), .RST(1'b0), .Q(
        round_reg[550]) );
  DFF \round_reg_reg[551]  ( .D(N563), .CLK(clk), .RST(1'b0), .Q(
        round_reg[551]) );
  DFF \round_reg_reg[552]  ( .D(N564), .CLK(clk), .RST(1'b0), .Q(
        round_reg[552]) );
  DFF \round_reg_reg[553]  ( .D(N565), .CLK(clk), .RST(1'b0), .Q(
        round_reg[553]) );
  DFF \round_reg_reg[554]  ( .D(N566), .CLK(clk), .RST(1'b0), .Q(
        round_reg[554]) );
  DFF \round_reg_reg[555]  ( .D(N567), .CLK(clk), .RST(1'b0), .Q(
        round_reg[555]) );
  DFF \round_reg_reg[556]  ( .D(N568), .CLK(clk), .RST(1'b0), .Q(
        round_reg[556]) );
  DFF \round_reg_reg[557]  ( .D(N569), .CLK(clk), .RST(1'b0), .Q(
        round_reg[557]) );
  DFF \round_reg_reg[558]  ( .D(N570), .CLK(clk), .RST(1'b0), .Q(
        round_reg[558]) );
  DFF \round_reg_reg[559]  ( .D(N571), .CLK(clk), .RST(1'b0), .Q(
        round_reg[559]) );
  DFF \round_reg_reg[560]  ( .D(N572), .CLK(clk), .RST(1'b0), .Q(
        round_reg[560]) );
  DFF \round_reg_reg[561]  ( .D(N573), .CLK(clk), .RST(1'b0), .Q(
        round_reg[561]) );
  DFF \round_reg_reg[562]  ( .D(N574), .CLK(clk), .RST(1'b0), .Q(
        round_reg[562]) );
  DFF \round_reg_reg[563]  ( .D(N575), .CLK(clk), .RST(1'b0), .Q(
        round_reg[563]) );
  DFF \round_reg_reg[564]  ( .D(N576), .CLK(clk), .RST(1'b0), .Q(
        round_reg[564]) );
  DFF \round_reg_reg[565]  ( .D(N577), .CLK(clk), .RST(1'b0), .Q(
        round_reg[565]) );
  DFF \round_reg_reg[566]  ( .D(N578), .CLK(clk), .RST(1'b0), .Q(
        round_reg[566]) );
  DFF \round_reg_reg[567]  ( .D(N579), .CLK(clk), .RST(1'b0), .Q(
        round_reg[567]) );
  DFF \round_reg_reg[568]  ( .D(N580), .CLK(clk), .RST(1'b0), .Q(
        round_reg[568]) );
  DFF \round_reg_reg[569]  ( .D(N581), .CLK(clk), .RST(1'b0), .Q(
        round_reg[569]) );
  DFF \round_reg_reg[570]  ( .D(N582), .CLK(clk), .RST(1'b0), .Q(
        round_reg[570]) );
  DFF \round_reg_reg[571]  ( .D(N583), .CLK(clk), .RST(1'b0), .Q(
        round_reg[571]) );
  DFF \round_reg_reg[572]  ( .D(N584), .CLK(clk), .RST(1'b0), .Q(
        round_reg[572]) );
  DFF \round_reg_reg[573]  ( .D(N585), .CLK(clk), .RST(1'b0), .Q(
        round_reg[573]) );
  DFF \round_reg_reg[574]  ( .D(N586), .CLK(clk), .RST(1'b0), .Q(
        round_reg[574]) );
  DFF \round_reg_reg[575]  ( .D(N587), .CLK(clk), .RST(1'b0), .Q(
        round_reg[575]) );
  DFF \round_reg_reg[576]  ( .D(N588), .CLK(clk), .RST(1'b0), .Q(
        round_reg[576]) );
  DFF \round_reg_reg[577]  ( .D(N589), .CLK(clk), .RST(1'b0), .Q(
        round_reg[577]) );
  DFF \round_reg_reg[578]  ( .D(N590), .CLK(clk), .RST(1'b0), .Q(
        round_reg[578]) );
  DFF \round_reg_reg[579]  ( .D(N591), .CLK(clk), .RST(1'b0), .Q(
        round_reg[579]) );
  DFF \round_reg_reg[580]  ( .D(N592), .CLK(clk), .RST(1'b0), .Q(
        round_reg[580]) );
  DFF \round_reg_reg[581]  ( .D(N593), .CLK(clk), .RST(1'b0), .Q(
        round_reg[581]) );
  DFF \round_reg_reg[582]  ( .D(N594), .CLK(clk), .RST(1'b0), .Q(
        round_reg[582]) );
  DFF \round_reg_reg[583]  ( .D(N595), .CLK(clk), .RST(1'b0), .Q(
        round_reg[583]) );
  DFF \round_reg_reg[584]  ( .D(N596), .CLK(clk), .RST(1'b0), .Q(
        round_reg[584]) );
  DFF \round_reg_reg[585]  ( .D(N597), .CLK(clk), .RST(1'b0), .Q(
        round_reg[585]) );
  DFF \round_reg_reg[586]  ( .D(N598), .CLK(clk), .RST(1'b0), .Q(
        round_reg[586]) );
  DFF \round_reg_reg[587]  ( .D(N599), .CLK(clk), .RST(1'b0), .Q(
        round_reg[587]) );
  DFF \round_reg_reg[588]  ( .D(N600), .CLK(clk), .RST(1'b0), .Q(
        round_reg[588]) );
  DFF \round_reg_reg[589]  ( .D(N601), .CLK(clk), .RST(1'b0), .Q(
        round_reg[589]) );
  DFF \round_reg_reg[590]  ( .D(N602), .CLK(clk), .RST(1'b0), .Q(
        round_reg[590]) );
  DFF \round_reg_reg[591]  ( .D(N603), .CLK(clk), .RST(1'b0), .Q(
        round_reg[591]) );
  DFF \round_reg_reg[592]  ( .D(N604), .CLK(clk), .RST(1'b0), .Q(
        round_reg[592]) );
  DFF \round_reg_reg[593]  ( .D(N605), .CLK(clk), .RST(1'b0), .Q(
        round_reg[593]) );
  DFF \round_reg_reg[594]  ( .D(N606), .CLK(clk), .RST(1'b0), .Q(
        round_reg[594]) );
  DFF \round_reg_reg[595]  ( .D(N607), .CLK(clk), .RST(1'b0), .Q(
        round_reg[595]) );
  DFF \round_reg_reg[596]  ( .D(N608), .CLK(clk), .RST(1'b0), .Q(
        round_reg[596]) );
  DFF \round_reg_reg[597]  ( .D(N609), .CLK(clk), .RST(1'b0), .Q(
        round_reg[597]) );
  DFF \round_reg_reg[598]  ( .D(N610), .CLK(clk), .RST(1'b0), .Q(
        round_reg[598]) );
  DFF \round_reg_reg[599]  ( .D(N611), .CLK(clk), .RST(1'b0), .Q(
        round_reg[599]) );
  DFF \round_reg_reg[600]  ( .D(N612), .CLK(clk), .RST(1'b0), .Q(
        round_reg[600]) );
  DFF \round_reg_reg[601]  ( .D(N613), .CLK(clk), .RST(1'b0), .Q(
        round_reg[601]) );
  DFF \round_reg_reg[602]  ( .D(N614), .CLK(clk), .RST(1'b0), .Q(
        round_reg[602]) );
  DFF \round_reg_reg[603]  ( .D(N615), .CLK(clk), .RST(1'b0), .Q(
        round_reg[603]) );
  DFF \round_reg_reg[604]  ( .D(N616), .CLK(clk), .RST(1'b0), .Q(
        round_reg[604]) );
  DFF \round_reg_reg[605]  ( .D(N617), .CLK(clk), .RST(1'b0), .Q(
        round_reg[605]) );
  DFF \round_reg_reg[606]  ( .D(N618), .CLK(clk), .RST(1'b0), .Q(
        round_reg[606]) );
  DFF \round_reg_reg[607]  ( .D(N619), .CLK(clk), .RST(1'b0), .Q(
        round_reg[607]) );
  DFF \round_reg_reg[608]  ( .D(N620), .CLK(clk), .RST(1'b0), .Q(
        round_reg[608]) );
  DFF \round_reg_reg[609]  ( .D(N621), .CLK(clk), .RST(1'b0), .Q(
        round_reg[609]) );
  DFF \round_reg_reg[610]  ( .D(N622), .CLK(clk), .RST(1'b0), .Q(
        round_reg[610]) );
  DFF \round_reg_reg[611]  ( .D(N623), .CLK(clk), .RST(1'b0), .Q(
        round_reg[611]) );
  DFF \round_reg_reg[612]  ( .D(N624), .CLK(clk), .RST(1'b0), .Q(
        round_reg[612]) );
  DFF \round_reg_reg[613]  ( .D(N625), .CLK(clk), .RST(1'b0), .Q(
        round_reg[613]) );
  DFF \round_reg_reg[614]  ( .D(N626), .CLK(clk), .RST(1'b0), .Q(
        round_reg[614]) );
  DFF \round_reg_reg[615]  ( .D(N627), .CLK(clk), .RST(1'b0), .Q(
        round_reg[615]) );
  DFF \round_reg_reg[616]  ( .D(N628), .CLK(clk), .RST(1'b0), .Q(
        round_reg[616]) );
  DFF \round_reg_reg[617]  ( .D(N629), .CLK(clk), .RST(1'b0), .Q(
        round_reg[617]) );
  DFF \round_reg_reg[618]  ( .D(N630), .CLK(clk), .RST(1'b0), .Q(
        round_reg[618]) );
  DFF \round_reg_reg[619]  ( .D(N631), .CLK(clk), .RST(1'b0), .Q(
        round_reg[619]) );
  DFF \round_reg_reg[620]  ( .D(N632), .CLK(clk), .RST(1'b0), .Q(
        round_reg[620]) );
  DFF \round_reg_reg[621]  ( .D(N633), .CLK(clk), .RST(1'b0), .Q(
        round_reg[621]) );
  DFF \round_reg_reg[622]  ( .D(N634), .CLK(clk), .RST(1'b0), .Q(
        round_reg[622]) );
  DFF \round_reg_reg[623]  ( .D(N635), .CLK(clk), .RST(1'b0), .Q(
        round_reg[623]) );
  DFF \round_reg_reg[624]  ( .D(N636), .CLK(clk), .RST(1'b0), .Q(
        round_reg[624]) );
  DFF \round_reg_reg[625]  ( .D(N637), .CLK(clk), .RST(1'b0), .Q(
        round_reg[625]) );
  DFF \round_reg_reg[626]  ( .D(N638), .CLK(clk), .RST(1'b0), .Q(
        round_reg[626]) );
  DFF \round_reg_reg[627]  ( .D(N639), .CLK(clk), .RST(1'b0), .Q(
        round_reg[627]) );
  DFF \round_reg_reg[628]  ( .D(N640), .CLK(clk), .RST(1'b0), .Q(
        round_reg[628]) );
  DFF \round_reg_reg[629]  ( .D(N641), .CLK(clk), .RST(1'b0), .Q(
        round_reg[629]) );
  DFF \round_reg_reg[630]  ( .D(N642), .CLK(clk), .RST(1'b0), .Q(
        round_reg[630]) );
  DFF \round_reg_reg[631]  ( .D(N643), .CLK(clk), .RST(1'b0), .Q(
        round_reg[631]) );
  DFF \round_reg_reg[632]  ( .D(N644), .CLK(clk), .RST(1'b0), .Q(
        round_reg[632]) );
  DFF \round_reg_reg[633]  ( .D(N645), .CLK(clk), .RST(1'b0), .Q(
        round_reg[633]) );
  DFF \round_reg_reg[634]  ( .D(N646), .CLK(clk), .RST(1'b0), .Q(
        round_reg[634]) );
  DFF \round_reg_reg[635]  ( .D(N647), .CLK(clk), .RST(1'b0), .Q(
        round_reg[635]) );
  DFF \round_reg_reg[636]  ( .D(N648), .CLK(clk), .RST(1'b0), .Q(
        round_reg[636]) );
  DFF \round_reg_reg[637]  ( .D(N649), .CLK(clk), .RST(1'b0), .Q(
        round_reg[637]) );
  DFF \round_reg_reg[638]  ( .D(N650), .CLK(clk), .RST(1'b0), .Q(
        round_reg[638]) );
  DFF \round_reg_reg[639]  ( .D(N651), .CLK(clk), .RST(1'b0), .Q(
        round_reg[639]) );
  DFF \round_reg_reg[640]  ( .D(N652), .CLK(clk), .RST(1'b0), .Q(
        round_reg[640]) );
  DFF \round_reg_reg[641]  ( .D(N653), .CLK(clk), .RST(1'b0), .Q(
        round_reg[641]) );
  DFF \round_reg_reg[642]  ( .D(N654), .CLK(clk), .RST(1'b0), .Q(
        round_reg[642]) );
  DFF \round_reg_reg[643]  ( .D(N655), .CLK(clk), .RST(1'b0), .Q(
        round_reg[643]) );
  DFF \round_reg_reg[644]  ( .D(N656), .CLK(clk), .RST(1'b0), .Q(
        round_reg[644]) );
  DFF \round_reg_reg[645]  ( .D(N657), .CLK(clk), .RST(1'b0), .Q(
        round_reg[645]) );
  DFF \round_reg_reg[646]  ( .D(N658), .CLK(clk), .RST(1'b0), .Q(
        round_reg[646]) );
  DFF \round_reg_reg[647]  ( .D(N659), .CLK(clk), .RST(1'b0), .Q(
        round_reg[647]) );
  DFF \round_reg_reg[648]  ( .D(N660), .CLK(clk), .RST(1'b0), .Q(
        round_reg[648]) );
  DFF \round_reg_reg[649]  ( .D(N661), .CLK(clk), .RST(1'b0), .Q(
        round_reg[649]) );
  DFF \round_reg_reg[650]  ( .D(N662), .CLK(clk), .RST(1'b0), .Q(
        round_reg[650]) );
  DFF \round_reg_reg[651]  ( .D(N663), .CLK(clk), .RST(1'b0), .Q(
        round_reg[651]) );
  DFF \round_reg_reg[652]  ( .D(N664), .CLK(clk), .RST(1'b0), .Q(
        round_reg[652]) );
  DFF \round_reg_reg[653]  ( .D(N665), .CLK(clk), .RST(1'b0), .Q(
        round_reg[653]) );
  DFF \round_reg_reg[654]  ( .D(N666), .CLK(clk), .RST(1'b0), .Q(
        round_reg[654]) );
  DFF \round_reg_reg[655]  ( .D(N667), .CLK(clk), .RST(1'b0), .Q(
        round_reg[655]) );
  DFF \round_reg_reg[656]  ( .D(N668), .CLK(clk), .RST(1'b0), .Q(
        round_reg[656]) );
  DFF \round_reg_reg[657]  ( .D(N669), .CLK(clk), .RST(1'b0), .Q(
        round_reg[657]) );
  DFF \round_reg_reg[658]  ( .D(N670), .CLK(clk), .RST(1'b0), .Q(
        round_reg[658]) );
  DFF \round_reg_reg[659]  ( .D(N671), .CLK(clk), .RST(1'b0), .Q(
        round_reg[659]) );
  DFF \round_reg_reg[660]  ( .D(N672), .CLK(clk), .RST(1'b0), .Q(
        round_reg[660]) );
  DFF \round_reg_reg[661]  ( .D(N673), .CLK(clk), .RST(1'b0), .Q(
        round_reg[661]) );
  DFF \round_reg_reg[662]  ( .D(N674), .CLK(clk), .RST(1'b0), .Q(
        round_reg[662]) );
  DFF \round_reg_reg[663]  ( .D(N675), .CLK(clk), .RST(1'b0), .Q(
        round_reg[663]) );
  DFF \round_reg_reg[664]  ( .D(N676), .CLK(clk), .RST(1'b0), .Q(
        round_reg[664]) );
  DFF \round_reg_reg[665]  ( .D(N677), .CLK(clk), .RST(1'b0), .Q(
        round_reg[665]) );
  DFF \round_reg_reg[666]  ( .D(N678), .CLK(clk), .RST(1'b0), .Q(
        round_reg[666]) );
  DFF \round_reg_reg[667]  ( .D(N679), .CLK(clk), .RST(1'b0), .Q(
        round_reg[667]) );
  DFF \round_reg_reg[668]  ( .D(N680), .CLK(clk), .RST(1'b0), .Q(
        round_reg[668]) );
  DFF \round_reg_reg[669]  ( .D(N681), .CLK(clk), .RST(1'b0), .Q(
        round_reg[669]) );
  DFF \round_reg_reg[670]  ( .D(N682), .CLK(clk), .RST(1'b0), .Q(
        round_reg[670]) );
  DFF \round_reg_reg[671]  ( .D(N683), .CLK(clk), .RST(1'b0), .Q(
        round_reg[671]) );
  DFF \round_reg_reg[672]  ( .D(N684), .CLK(clk), .RST(1'b0), .Q(
        round_reg[672]) );
  DFF \round_reg_reg[673]  ( .D(N685), .CLK(clk), .RST(1'b0), .Q(
        round_reg[673]) );
  DFF \round_reg_reg[674]  ( .D(N686), .CLK(clk), .RST(1'b0), .Q(
        round_reg[674]) );
  DFF \round_reg_reg[675]  ( .D(N687), .CLK(clk), .RST(1'b0), .Q(
        round_reg[675]) );
  DFF \round_reg_reg[676]  ( .D(N688), .CLK(clk), .RST(1'b0), .Q(
        round_reg[676]) );
  DFF \round_reg_reg[677]  ( .D(N689), .CLK(clk), .RST(1'b0), .Q(
        round_reg[677]) );
  DFF \round_reg_reg[678]  ( .D(N690), .CLK(clk), .RST(1'b0), .Q(
        round_reg[678]) );
  DFF \round_reg_reg[679]  ( .D(N691), .CLK(clk), .RST(1'b0), .Q(
        round_reg[679]) );
  DFF \round_reg_reg[680]  ( .D(N692), .CLK(clk), .RST(1'b0), .Q(
        round_reg[680]) );
  DFF \round_reg_reg[681]  ( .D(N693), .CLK(clk), .RST(1'b0), .Q(
        round_reg[681]) );
  DFF \round_reg_reg[682]  ( .D(N694), .CLK(clk), .RST(1'b0), .Q(
        round_reg[682]) );
  DFF \round_reg_reg[683]  ( .D(N695), .CLK(clk), .RST(1'b0), .Q(
        round_reg[683]) );
  DFF \round_reg_reg[684]  ( .D(N696), .CLK(clk), .RST(1'b0), .Q(
        round_reg[684]) );
  DFF \round_reg_reg[685]  ( .D(N697), .CLK(clk), .RST(1'b0), .Q(
        round_reg[685]) );
  DFF \round_reg_reg[686]  ( .D(N698), .CLK(clk), .RST(1'b0), .Q(
        round_reg[686]) );
  DFF \round_reg_reg[687]  ( .D(N699), .CLK(clk), .RST(1'b0), .Q(
        round_reg[687]) );
  DFF \round_reg_reg[688]  ( .D(N700), .CLK(clk), .RST(1'b0), .Q(
        round_reg[688]) );
  DFF \round_reg_reg[689]  ( .D(N701), .CLK(clk), .RST(1'b0), .Q(
        round_reg[689]) );
  DFF \round_reg_reg[690]  ( .D(N702), .CLK(clk), .RST(1'b0), .Q(
        round_reg[690]) );
  DFF \round_reg_reg[691]  ( .D(N703), .CLK(clk), .RST(1'b0), .Q(
        round_reg[691]) );
  DFF \round_reg_reg[692]  ( .D(N704), .CLK(clk), .RST(1'b0), .Q(
        round_reg[692]) );
  DFF \round_reg_reg[693]  ( .D(N705), .CLK(clk), .RST(1'b0), .Q(
        round_reg[693]) );
  DFF \round_reg_reg[694]  ( .D(N706), .CLK(clk), .RST(1'b0), .Q(
        round_reg[694]) );
  DFF \round_reg_reg[695]  ( .D(N707), .CLK(clk), .RST(1'b0), .Q(
        round_reg[695]) );
  DFF \round_reg_reg[696]  ( .D(N708), .CLK(clk), .RST(1'b0), .Q(
        round_reg[696]) );
  DFF \round_reg_reg[697]  ( .D(N709), .CLK(clk), .RST(1'b0), .Q(
        round_reg[697]) );
  DFF \round_reg_reg[698]  ( .D(N710), .CLK(clk), .RST(1'b0), .Q(
        round_reg[698]) );
  DFF \round_reg_reg[699]  ( .D(N711), .CLK(clk), .RST(1'b0), .Q(
        round_reg[699]) );
  DFF \round_reg_reg[700]  ( .D(N712), .CLK(clk), .RST(1'b0), .Q(
        round_reg[700]) );
  DFF \round_reg_reg[701]  ( .D(N713), .CLK(clk), .RST(1'b0), .Q(
        round_reg[701]) );
  DFF \round_reg_reg[702]  ( .D(N714), .CLK(clk), .RST(1'b0), .Q(
        round_reg[702]) );
  DFF \round_reg_reg[703]  ( .D(N715), .CLK(clk), .RST(1'b0), .Q(
        round_reg[703]) );
  DFF \round_reg_reg[704]  ( .D(N716), .CLK(clk), .RST(1'b0), .Q(
        round_reg[704]) );
  DFF \round_reg_reg[705]  ( .D(N717), .CLK(clk), .RST(1'b0), .Q(
        round_reg[705]) );
  DFF \round_reg_reg[706]  ( .D(N718), .CLK(clk), .RST(1'b0), .Q(
        round_reg[706]) );
  DFF \round_reg_reg[707]  ( .D(N719), .CLK(clk), .RST(1'b0), .Q(
        round_reg[707]) );
  DFF \round_reg_reg[708]  ( .D(N720), .CLK(clk), .RST(1'b0), .Q(
        round_reg[708]) );
  DFF \round_reg_reg[709]  ( .D(N721), .CLK(clk), .RST(1'b0), .Q(
        round_reg[709]) );
  DFF \round_reg_reg[710]  ( .D(N722), .CLK(clk), .RST(1'b0), .Q(
        round_reg[710]) );
  DFF \round_reg_reg[711]  ( .D(N723), .CLK(clk), .RST(1'b0), .Q(
        round_reg[711]) );
  DFF \round_reg_reg[712]  ( .D(N724), .CLK(clk), .RST(1'b0), .Q(
        round_reg[712]) );
  DFF \round_reg_reg[713]  ( .D(N725), .CLK(clk), .RST(1'b0), .Q(
        round_reg[713]) );
  DFF \round_reg_reg[714]  ( .D(N726), .CLK(clk), .RST(1'b0), .Q(
        round_reg[714]) );
  DFF \round_reg_reg[715]  ( .D(N727), .CLK(clk), .RST(1'b0), .Q(
        round_reg[715]) );
  DFF \round_reg_reg[716]  ( .D(N728), .CLK(clk), .RST(1'b0), .Q(
        round_reg[716]) );
  DFF \round_reg_reg[717]  ( .D(N729), .CLK(clk), .RST(1'b0), .Q(
        round_reg[717]) );
  DFF \round_reg_reg[718]  ( .D(N730), .CLK(clk), .RST(1'b0), .Q(
        round_reg[718]) );
  DFF \round_reg_reg[719]  ( .D(N731), .CLK(clk), .RST(1'b0), .Q(
        round_reg[719]) );
  DFF \round_reg_reg[720]  ( .D(N732), .CLK(clk), .RST(1'b0), .Q(
        round_reg[720]) );
  DFF \round_reg_reg[721]  ( .D(N733), .CLK(clk), .RST(1'b0), .Q(
        round_reg[721]) );
  DFF \round_reg_reg[722]  ( .D(N734), .CLK(clk), .RST(1'b0), .Q(
        round_reg[722]) );
  DFF \round_reg_reg[723]  ( .D(N735), .CLK(clk), .RST(1'b0), .Q(
        round_reg[723]) );
  DFF \round_reg_reg[724]  ( .D(N736), .CLK(clk), .RST(1'b0), .Q(
        round_reg[724]) );
  DFF \round_reg_reg[725]  ( .D(N737), .CLK(clk), .RST(1'b0), .Q(
        round_reg[725]) );
  DFF \round_reg_reg[726]  ( .D(N738), .CLK(clk), .RST(1'b0), .Q(
        round_reg[726]) );
  DFF \round_reg_reg[727]  ( .D(N739), .CLK(clk), .RST(1'b0), .Q(
        round_reg[727]) );
  DFF \round_reg_reg[728]  ( .D(N740), .CLK(clk), .RST(1'b0), .Q(
        round_reg[728]) );
  DFF \round_reg_reg[729]  ( .D(N741), .CLK(clk), .RST(1'b0), .Q(
        round_reg[729]) );
  DFF \round_reg_reg[730]  ( .D(N742), .CLK(clk), .RST(1'b0), .Q(
        round_reg[730]) );
  DFF \round_reg_reg[731]  ( .D(N743), .CLK(clk), .RST(1'b0), .Q(
        round_reg[731]) );
  DFF \round_reg_reg[732]  ( .D(N744), .CLK(clk), .RST(1'b0), .Q(
        round_reg[732]) );
  DFF \round_reg_reg[733]  ( .D(N745), .CLK(clk), .RST(1'b0), .Q(
        round_reg[733]) );
  DFF \round_reg_reg[734]  ( .D(N746), .CLK(clk), .RST(1'b0), .Q(
        round_reg[734]) );
  DFF \round_reg_reg[735]  ( .D(N747), .CLK(clk), .RST(1'b0), .Q(
        round_reg[735]) );
  DFF \round_reg_reg[736]  ( .D(N748), .CLK(clk), .RST(1'b0), .Q(
        round_reg[736]) );
  DFF \round_reg_reg[737]  ( .D(N749), .CLK(clk), .RST(1'b0), .Q(
        round_reg[737]) );
  DFF \round_reg_reg[738]  ( .D(N750), .CLK(clk), .RST(1'b0), .Q(
        round_reg[738]) );
  DFF \round_reg_reg[739]  ( .D(N751), .CLK(clk), .RST(1'b0), .Q(
        round_reg[739]) );
  DFF \round_reg_reg[740]  ( .D(N752), .CLK(clk), .RST(1'b0), .Q(
        round_reg[740]) );
  DFF \round_reg_reg[741]  ( .D(N753), .CLK(clk), .RST(1'b0), .Q(
        round_reg[741]) );
  DFF \round_reg_reg[742]  ( .D(N754), .CLK(clk), .RST(1'b0), .Q(
        round_reg[742]) );
  DFF \round_reg_reg[743]  ( .D(N755), .CLK(clk), .RST(1'b0), .Q(
        round_reg[743]) );
  DFF \round_reg_reg[744]  ( .D(N756), .CLK(clk), .RST(1'b0), .Q(
        round_reg[744]) );
  DFF \round_reg_reg[745]  ( .D(N757), .CLK(clk), .RST(1'b0), .Q(
        round_reg[745]) );
  DFF \round_reg_reg[746]  ( .D(N758), .CLK(clk), .RST(1'b0), .Q(
        round_reg[746]) );
  DFF \round_reg_reg[747]  ( .D(N759), .CLK(clk), .RST(1'b0), .Q(
        round_reg[747]) );
  DFF \round_reg_reg[748]  ( .D(N760), .CLK(clk), .RST(1'b0), .Q(
        round_reg[748]) );
  DFF \round_reg_reg[749]  ( .D(N761), .CLK(clk), .RST(1'b0), .Q(
        round_reg[749]) );
  DFF \round_reg_reg[750]  ( .D(N762), .CLK(clk), .RST(1'b0), .Q(
        round_reg[750]) );
  DFF \round_reg_reg[751]  ( .D(N763), .CLK(clk), .RST(1'b0), .Q(
        round_reg[751]) );
  DFF \round_reg_reg[752]  ( .D(N764), .CLK(clk), .RST(1'b0), .Q(
        round_reg[752]) );
  DFF \round_reg_reg[753]  ( .D(N765), .CLK(clk), .RST(1'b0), .Q(
        round_reg[753]) );
  DFF \round_reg_reg[754]  ( .D(N766), .CLK(clk), .RST(1'b0), .Q(
        round_reg[754]) );
  DFF \round_reg_reg[755]  ( .D(N767), .CLK(clk), .RST(1'b0), .Q(
        round_reg[755]) );
  DFF \round_reg_reg[756]  ( .D(N768), .CLK(clk), .RST(1'b0), .Q(
        round_reg[756]) );
  DFF \round_reg_reg[757]  ( .D(N769), .CLK(clk), .RST(1'b0), .Q(
        round_reg[757]) );
  DFF \round_reg_reg[758]  ( .D(N770), .CLK(clk), .RST(1'b0), .Q(
        round_reg[758]) );
  DFF \round_reg_reg[759]  ( .D(N771), .CLK(clk), .RST(1'b0), .Q(
        round_reg[759]) );
  DFF \round_reg_reg[760]  ( .D(N772), .CLK(clk), .RST(1'b0), .Q(
        round_reg[760]) );
  DFF \round_reg_reg[761]  ( .D(N773), .CLK(clk), .RST(1'b0), .Q(
        round_reg[761]) );
  DFF \round_reg_reg[762]  ( .D(N774), .CLK(clk), .RST(1'b0), .Q(
        round_reg[762]) );
  DFF \round_reg_reg[763]  ( .D(N775), .CLK(clk), .RST(1'b0), .Q(
        round_reg[763]) );
  DFF \round_reg_reg[764]  ( .D(N776), .CLK(clk), .RST(1'b0), .Q(
        round_reg[764]) );
  DFF \round_reg_reg[765]  ( .D(N777), .CLK(clk), .RST(1'b0), .Q(
        round_reg[765]) );
  DFF \round_reg_reg[766]  ( .D(N778), .CLK(clk), .RST(1'b0), .Q(
        round_reg[766]) );
  DFF \round_reg_reg[767]  ( .D(N779), .CLK(clk), .RST(1'b0), .Q(
        round_reg[767]) );
  DFF \round_reg_reg[768]  ( .D(N780), .CLK(clk), .RST(1'b0), .Q(
        round_reg[768]) );
  DFF \round_reg_reg[769]  ( .D(N781), .CLK(clk), .RST(1'b0), .Q(
        round_reg[769]) );
  DFF \round_reg_reg[770]  ( .D(N782), .CLK(clk), .RST(1'b0), .Q(
        round_reg[770]) );
  DFF \round_reg_reg[771]  ( .D(N783), .CLK(clk), .RST(1'b0), .Q(
        round_reg[771]) );
  DFF \round_reg_reg[772]  ( .D(N784), .CLK(clk), .RST(1'b0), .Q(
        round_reg[772]) );
  DFF \round_reg_reg[773]  ( .D(N785), .CLK(clk), .RST(1'b0), .Q(
        round_reg[773]) );
  DFF \round_reg_reg[774]  ( .D(N786), .CLK(clk), .RST(1'b0), .Q(
        round_reg[774]) );
  DFF \round_reg_reg[775]  ( .D(N787), .CLK(clk), .RST(1'b0), .Q(
        round_reg[775]) );
  DFF \round_reg_reg[776]  ( .D(N788), .CLK(clk), .RST(1'b0), .Q(
        round_reg[776]) );
  DFF \round_reg_reg[777]  ( .D(N789), .CLK(clk), .RST(1'b0), .Q(
        round_reg[777]) );
  DFF \round_reg_reg[778]  ( .D(N790), .CLK(clk), .RST(1'b0), .Q(
        round_reg[778]) );
  DFF \round_reg_reg[779]  ( .D(N791), .CLK(clk), .RST(1'b0), .Q(
        round_reg[779]) );
  DFF \round_reg_reg[780]  ( .D(N792), .CLK(clk), .RST(1'b0), .Q(
        round_reg[780]) );
  DFF \round_reg_reg[781]  ( .D(N793), .CLK(clk), .RST(1'b0), .Q(
        round_reg[781]) );
  DFF \round_reg_reg[782]  ( .D(N794), .CLK(clk), .RST(1'b0), .Q(
        round_reg[782]) );
  DFF \round_reg_reg[783]  ( .D(N795), .CLK(clk), .RST(1'b0), .Q(
        round_reg[783]) );
  DFF \round_reg_reg[784]  ( .D(N796), .CLK(clk), .RST(1'b0), .Q(
        round_reg[784]) );
  DFF \round_reg_reg[785]  ( .D(N797), .CLK(clk), .RST(1'b0), .Q(
        round_reg[785]) );
  DFF \round_reg_reg[786]  ( .D(N798), .CLK(clk), .RST(1'b0), .Q(
        round_reg[786]) );
  DFF \round_reg_reg[787]  ( .D(N799), .CLK(clk), .RST(1'b0), .Q(
        round_reg[787]) );
  DFF \round_reg_reg[788]  ( .D(N800), .CLK(clk), .RST(1'b0), .Q(
        round_reg[788]) );
  DFF \round_reg_reg[789]  ( .D(N801), .CLK(clk), .RST(1'b0), .Q(
        round_reg[789]) );
  DFF \round_reg_reg[790]  ( .D(N802), .CLK(clk), .RST(1'b0), .Q(
        round_reg[790]) );
  DFF \round_reg_reg[791]  ( .D(N803), .CLK(clk), .RST(1'b0), .Q(
        round_reg[791]) );
  DFF \round_reg_reg[792]  ( .D(N804), .CLK(clk), .RST(1'b0), .Q(
        round_reg[792]) );
  DFF \round_reg_reg[793]  ( .D(N805), .CLK(clk), .RST(1'b0), .Q(
        round_reg[793]) );
  DFF \round_reg_reg[794]  ( .D(N806), .CLK(clk), .RST(1'b0), .Q(
        round_reg[794]) );
  DFF \round_reg_reg[795]  ( .D(N807), .CLK(clk), .RST(1'b0), .Q(
        round_reg[795]) );
  DFF \round_reg_reg[796]  ( .D(N808), .CLK(clk), .RST(1'b0), .Q(
        round_reg[796]) );
  DFF \round_reg_reg[797]  ( .D(N809), .CLK(clk), .RST(1'b0), .Q(
        round_reg[797]) );
  DFF \round_reg_reg[798]  ( .D(N810), .CLK(clk), .RST(1'b0), .Q(
        round_reg[798]) );
  DFF \round_reg_reg[799]  ( .D(N811), .CLK(clk), .RST(1'b0), .Q(
        round_reg[799]) );
  DFF \round_reg_reg[800]  ( .D(N812), .CLK(clk), .RST(1'b0), .Q(
        round_reg[800]) );
  DFF \round_reg_reg[801]  ( .D(N813), .CLK(clk), .RST(1'b0), .Q(
        round_reg[801]) );
  DFF \round_reg_reg[802]  ( .D(N814), .CLK(clk), .RST(1'b0), .Q(
        round_reg[802]) );
  DFF \round_reg_reg[803]  ( .D(N815), .CLK(clk), .RST(1'b0), .Q(
        round_reg[803]) );
  DFF \round_reg_reg[804]  ( .D(N816), .CLK(clk), .RST(1'b0), .Q(
        round_reg[804]) );
  DFF \round_reg_reg[805]  ( .D(N817), .CLK(clk), .RST(1'b0), .Q(
        round_reg[805]) );
  DFF \round_reg_reg[806]  ( .D(N818), .CLK(clk), .RST(1'b0), .Q(
        round_reg[806]) );
  DFF \round_reg_reg[807]  ( .D(N819), .CLK(clk), .RST(1'b0), .Q(
        round_reg[807]) );
  DFF \round_reg_reg[808]  ( .D(N820), .CLK(clk), .RST(1'b0), .Q(
        round_reg[808]) );
  DFF \round_reg_reg[809]  ( .D(N821), .CLK(clk), .RST(1'b0), .Q(
        round_reg[809]) );
  DFF \round_reg_reg[810]  ( .D(N822), .CLK(clk), .RST(1'b0), .Q(
        round_reg[810]) );
  DFF \round_reg_reg[811]  ( .D(N823), .CLK(clk), .RST(1'b0), .Q(
        round_reg[811]) );
  DFF \round_reg_reg[812]  ( .D(N824), .CLK(clk), .RST(1'b0), .Q(
        round_reg[812]) );
  DFF \round_reg_reg[813]  ( .D(N825), .CLK(clk), .RST(1'b0), .Q(
        round_reg[813]) );
  DFF \round_reg_reg[814]  ( .D(N826), .CLK(clk), .RST(1'b0), .Q(
        round_reg[814]) );
  DFF \round_reg_reg[815]  ( .D(N827), .CLK(clk), .RST(1'b0), .Q(
        round_reg[815]) );
  DFF \round_reg_reg[816]  ( .D(N828), .CLK(clk), .RST(1'b0), .Q(
        round_reg[816]) );
  DFF \round_reg_reg[817]  ( .D(N829), .CLK(clk), .RST(1'b0), .Q(
        round_reg[817]) );
  DFF \round_reg_reg[818]  ( .D(N830), .CLK(clk), .RST(1'b0), .Q(
        round_reg[818]) );
  DFF \round_reg_reg[819]  ( .D(N831), .CLK(clk), .RST(1'b0), .Q(
        round_reg[819]) );
  DFF \round_reg_reg[820]  ( .D(N832), .CLK(clk), .RST(1'b0), .Q(
        round_reg[820]) );
  DFF \round_reg_reg[821]  ( .D(N833), .CLK(clk), .RST(1'b0), .Q(
        round_reg[821]) );
  DFF \round_reg_reg[822]  ( .D(N834), .CLK(clk), .RST(1'b0), .Q(
        round_reg[822]) );
  DFF \round_reg_reg[823]  ( .D(N835), .CLK(clk), .RST(1'b0), .Q(
        round_reg[823]) );
  DFF \round_reg_reg[824]  ( .D(N836), .CLK(clk), .RST(1'b0), .Q(
        round_reg[824]) );
  DFF \round_reg_reg[825]  ( .D(N837), .CLK(clk), .RST(1'b0), .Q(
        round_reg[825]) );
  DFF \round_reg_reg[826]  ( .D(N838), .CLK(clk), .RST(1'b0), .Q(
        round_reg[826]) );
  DFF \round_reg_reg[827]  ( .D(N839), .CLK(clk), .RST(1'b0), .Q(
        round_reg[827]) );
  DFF \round_reg_reg[828]  ( .D(N840), .CLK(clk), .RST(1'b0), .Q(
        round_reg[828]) );
  DFF \round_reg_reg[829]  ( .D(N841), .CLK(clk), .RST(1'b0), .Q(
        round_reg[829]) );
  DFF \round_reg_reg[830]  ( .D(N842), .CLK(clk), .RST(1'b0), .Q(
        round_reg[830]) );
  DFF \round_reg_reg[831]  ( .D(N843), .CLK(clk), .RST(1'b0), .Q(
        round_reg[831]) );
  DFF \round_reg_reg[832]  ( .D(N844), .CLK(clk), .RST(1'b0), .Q(
        round_reg[832]) );
  DFF \round_reg_reg[833]  ( .D(N845), .CLK(clk), .RST(1'b0), .Q(
        round_reg[833]) );
  DFF \round_reg_reg[834]  ( .D(N846), .CLK(clk), .RST(1'b0), .Q(
        round_reg[834]) );
  DFF \round_reg_reg[835]  ( .D(N847), .CLK(clk), .RST(1'b0), .Q(
        round_reg[835]) );
  DFF \round_reg_reg[836]  ( .D(N848), .CLK(clk), .RST(1'b0), .Q(
        round_reg[836]) );
  DFF \round_reg_reg[837]  ( .D(N849), .CLK(clk), .RST(1'b0), .Q(
        round_reg[837]) );
  DFF \round_reg_reg[838]  ( .D(N850), .CLK(clk), .RST(1'b0), .Q(
        round_reg[838]) );
  DFF \round_reg_reg[839]  ( .D(N851), .CLK(clk), .RST(1'b0), .Q(
        round_reg[839]) );
  DFF \round_reg_reg[840]  ( .D(N852), .CLK(clk), .RST(1'b0), .Q(
        round_reg[840]) );
  DFF \round_reg_reg[841]  ( .D(N853), .CLK(clk), .RST(1'b0), .Q(
        round_reg[841]) );
  DFF \round_reg_reg[842]  ( .D(N854), .CLK(clk), .RST(1'b0), .Q(
        round_reg[842]) );
  DFF \round_reg_reg[843]  ( .D(N855), .CLK(clk), .RST(1'b0), .Q(
        round_reg[843]) );
  DFF \round_reg_reg[844]  ( .D(N856), .CLK(clk), .RST(1'b0), .Q(
        round_reg[844]) );
  DFF \round_reg_reg[845]  ( .D(N857), .CLK(clk), .RST(1'b0), .Q(
        round_reg[845]) );
  DFF \round_reg_reg[846]  ( .D(N858), .CLK(clk), .RST(1'b0), .Q(
        round_reg[846]) );
  DFF \round_reg_reg[847]  ( .D(N859), .CLK(clk), .RST(1'b0), .Q(
        round_reg[847]) );
  DFF \round_reg_reg[848]  ( .D(N860), .CLK(clk), .RST(1'b0), .Q(
        round_reg[848]) );
  DFF \round_reg_reg[849]  ( .D(N861), .CLK(clk), .RST(1'b0), .Q(
        round_reg[849]) );
  DFF \round_reg_reg[850]  ( .D(N862), .CLK(clk), .RST(1'b0), .Q(
        round_reg[850]) );
  DFF \round_reg_reg[851]  ( .D(N863), .CLK(clk), .RST(1'b0), .Q(
        round_reg[851]) );
  DFF \round_reg_reg[852]  ( .D(N864), .CLK(clk), .RST(1'b0), .Q(
        round_reg[852]) );
  DFF \round_reg_reg[853]  ( .D(N865), .CLK(clk), .RST(1'b0), .Q(
        round_reg[853]) );
  DFF \round_reg_reg[854]  ( .D(N866), .CLK(clk), .RST(1'b0), .Q(
        round_reg[854]) );
  DFF \round_reg_reg[855]  ( .D(N867), .CLK(clk), .RST(1'b0), .Q(
        round_reg[855]) );
  DFF \round_reg_reg[856]  ( .D(N868), .CLK(clk), .RST(1'b0), .Q(
        round_reg[856]) );
  DFF \round_reg_reg[857]  ( .D(N869), .CLK(clk), .RST(1'b0), .Q(
        round_reg[857]) );
  DFF \round_reg_reg[858]  ( .D(N870), .CLK(clk), .RST(1'b0), .Q(
        round_reg[858]) );
  DFF \round_reg_reg[859]  ( .D(N871), .CLK(clk), .RST(1'b0), .Q(
        round_reg[859]) );
  DFF \round_reg_reg[860]  ( .D(N872), .CLK(clk), .RST(1'b0), .Q(
        round_reg[860]) );
  DFF \round_reg_reg[861]  ( .D(N873), .CLK(clk), .RST(1'b0), .Q(
        round_reg[861]) );
  DFF \round_reg_reg[862]  ( .D(N874), .CLK(clk), .RST(1'b0), .Q(
        round_reg[862]) );
  DFF \round_reg_reg[863]  ( .D(N875), .CLK(clk), .RST(1'b0), .Q(
        round_reg[863]) );
  DFF \round_reg_reg[864]  ( .D(N876), .CLK(clk), .RST(1'b0), .Q(
        round_reg[864]) );
  DFF \round_reg_reg[865]  ( .D(N877), .CLK(clk), .RST(1'b0), .Q(
        round_reg[865]) );
  DFF \round_reg_reg[866]  ( .D(N878), .CLK(clk), .RST(1'b0), .Q(
        round_reg[866]) );
  DFF \round_reg_reg[867]  ( .D(N879), .CLK(clk), .RST(1'b0), .Q(
        round_reg[867]) );
  DFF \round_reg_reg[868]  ( .D(N880), .CLK(clk), .RST(1'b0), .Q(
        round_reg[868]) );
  DFF \round_reg_reg[869]  ( .D(N881), .CLK(clk), .RST(1'b0), .Q(
        round_reg[869]) );
  DFF \round_reg_reg[870]  ( .D(N882), .CLK(clk), .RST(1'b0), .Q(
        round_reg[870]) );
  DFF \round_reg_reg[871]  ( .D(N883), .CLK(clk), .RST(1'b0), .Q(
        round_reg[871]) );
  DFF \round_reg_reg[872]  ( .D(N884), .CLK(clk), .RST(1'b0), .Q(
        round_reg[872]) );
  DFF \round_reg_reg[873]  ( .D(N885), .CLK(clk), .RST(1'b0), .Q(
        round_reg[873]) );
  DFF \round_reg_reg[874]  ( .D(N886), .CLK(clk), .RST(1'b0), .Q(
        round_reg[874]) );
  DFF \round_reg_reg[875]  ( .D(N887), .CLK(clk), .RST(1'b0), .Q(
        round_reg[875]) );
  DFF \round_reg_reg[876]  ( .D(N888), .CLK(clk), .RST(1'b0), .Q(
        round_reg[876]) );
  DFF \round_reg_reg[877]  ( .D(N889), .CLK(clk), .RST(1'b0), .Q(
        round_reg[877]) );
  DFF \round_reg_reg[878]  ( .D(N890), .CLK(clk), .RST(1'b0), .Q(
        round_reg[878]) );
  DFF \round_reg_reg[879]  ( .D(N891), .CLK(clk), .RST(1'b0), .Q(
        round_reg[879]) );
  DFF \round_reg_reg[880]  ( .D(N892), .CLK(clk), .RST(1'b0), .Q(
        round_reg[880]) );
  DFF \round_reg_reg[881]  ( .D(N893), .CLK(clk), .RST(1'b0), .Q(
        round_reg[881]) );
  DFF \round_reg_reg[882]  ( .D(N894), .CLK(clk), .RST(1'b0), .Q(
        round_reg[882]) );
  DFF \round_reg_reg[883]  ( .D(N895), .CLK(clk), .RST(1'b0), .Q(
        round_reg[883]) );
  DFF \round_reg_reg[884]  ( .D(N896), .CLK(clk), .RST(1'b0), .Q(
        round_reg[884]) );
  DFF \round_reg_reg[885]  ( .D(N897), .CLK(clk), .RST(1'b0), .Q(
        round_reg[885]) );
  DFF \round_reg_reg[886]  ( .D(N898), .CLK(clk), .RST(1'b0), .Q(
        round_reg[886]) );
  DFF \round_reg_reg[887]  ( .D(N899), .CLK(clk), .RST(1'b0), .Q(
        round_reg[887]) );
  DFF \round_reg_reg[888]  ( .D(N900), .CLK(clk), .RST(1'b0), .Q(
        round_reg[888]) );
  DFF \round_reg_reg[889]  ( .D(N901), .CLK(clk), .RST(1'b0), .Q(
        round_reg[889]) );
  DFF \round_reg_reg[890]  ( .D(N902), .CLK(clk), .RST(1'b0), .Q(
        round_reg[890]) );
  DFF \round_reg_reg[891]  ( .D(N903), .CLK(clk), .RST(1'b0), .Q(
        round_reg[891]) );
  DFF \round_reg_reg[892]  ( .D(N904), .CLK(clk), .RST(1'b0), .Q(
        round_reg[892]) );
  DFF \round_reg_reg[893]  ( .D(N905), .CLK(clk), .RST(1'b0), .Q(
        round_reg[893]) );
  DFF \round_reg_reg[894]  ( .D(N906), .CLK(clk), .RST(1'b0), .Q(
        round_reg[894]) );
  DFF \round_reg_reg[895]  ( .D(N907), .CLK(clk), .RST(1'b0), .Q(
        round_reg[895]) );
  DFF \round_reg_reg[896]  ( .D(N908), .CLK(clk), .RST(1'b0), .Q(
        round_reg[896]) );
  DFF \round_reg_reg[897]  ( .D(N909), .CLK(clk), .RST(1'b0), .Q(
        round_reg[897]) );
  DFF \round_reg_reg[898]  ( .D(N910), .CLK(clk), .RST(1'b0), .Q(
        round_reg[898]) );
  DFF \round_reg_reg[899]  ( .D(N911), .CLK(clk), .RST(1'b0), .Q(
        round_reg[899]) );
  DFF \round_reg_reg[900]  ( .D(N912), .CLK(clk), .RST(1'b0), .Q(
        round_reg[900]) );
  DFF \round_reg_reg[901]  ( .D(N913), .CLK(clk), .RST(1'b0), .Q(
        round_reg[901]) );
  DFF \round_reg_reg[902]  ( .D(N914), .CLK(clk), .RST(1'b0), .Q(
        round_reg[902]) );
  DFF \round_reg_reg[903]  ( .D(N915), .CLK(clk), .RST(1'b0), .Q(
        round_reg[903]) );
  DFF \round_reg_reg[904]  ( .D(N916), .CLK(clk), .RST(1'b0), .Q(
        round_reg[904]) );
  DFF \round_reg_reg[905]  ( .D(N917), .CLK(clk), .RST(1'b0), .Q(
        round_reg[905]) );
  DFF \round_reg_reg[906]  ( .D(N918), .CLK(clk), .RST(1'b0), .Q(
        round_reg[906]) );
  DFF \round_reg_reg[907]  ( .D(N919), .CLK(clk), .RST(1'b0), .Q(
        round_reg[907]) );
  DFF \round_reg_reg[908]  ( .D(N920), .CLK(clk), .RST(1'b0), .Q(
        round_reg[908]) );
  DFF \round_reg_reg[909]  ( .D(N921), .CLK(clk), .RST(1'b0), .Q(
        round_reg[909]) );
  DFF \round_reg_reg[910]  ( .D(N922), .CLK(clk), .RST(1'b0), .Q(
        round_reg[910]) );
  DFF \round_reg_reg[911]  ( .D(N923), .CLK(clk), .RST(1'b0), .Q(
        round_reg[911]) );
  DFF \round_reg_reg[912]  ( .D(N924), .CLK(clk), .RST(1'b0), .Q(
        round_reg[912]) );
  DFF \round_reg_reg[913]  ( .D(N925), .CLK(clk), .RST(1'b0), .Q(
        round_reg[913]) );
  DFF \round_reg_reg[914]  ( .D(N926), .CLK(clk), .RST(1'b0), .Q(
        round_reg[914]) );
  DFF \round_reg_reg[915]  ( .D(N927), .CLK(clk), .RST(1'b0), .Q(
        round_reg[915]) );
  DFF \round_reg_reg[916]  ( .D(N928), .CLK(clk), .RST(1'b0), .Q(
        round_reg[916]) );
  DFF \round_reg_reg[917]  ( .D(N929), .CLK(clk), .RST(1'b0), .Q(
        round_reg[917]) );
  DFF \round_reg_reg[918]  ( .D(N930), .CLK(clk), .RST(1'b0), .Q(
        round_reg[918]) );
  DFF \round_reg_reg[919]  ( .D(N931), .CLK(clk), .RST(1'b0), .Q(
        round_reg[919]) );
  DFF \round_reg_reg[920]  ( .D(N932), .CLK(clk), .RST(1'b0), .Q(
        round_reg[920]) );
  DFF \round_reg_reg[921]  ( .D(N933), .CLK(clk), .RST(1'b0), .Q(
        round_reg[921]) );
  DFF \round_reg_reg[922]  ( .D(N934), .CLK(clk), .RST(1'b0), .Q(
        round_reg[922]) );
  DFF \round_reg_reg[923]  ( .D(N935), .CLK(clk), .RST(1'b0), .Q(
        round_reg[923]) );
  DFF \round_reg_reg[924]  ( .D(N936), .CLK(clk), .RST(1'b0), .Q(
        round_reg[924]) );
  DFF \round_reg_reg[925]  ( .D(N937), .CLK(clk), .RST(1'b0), .Q(
        round_reg[925]) );
  DFF \round_reg_reg[926]  ( .D(N938), .CLK(clk), .RST(1'b0), .Q(
        round_reg[926]) );
  DFF \round_reg_reg[927]  ( .D(N939), .CLK(clk), .RST(1'b0), .Q(
        round_reg[927]) );
  DFF \round_reg_reg[928]  ( .D(N940), .CLK(clk), .RST(1'b0), .Q(
        round_reg[928]) );
  DFF \round_reg_reg[929]  ( .D(N941), .CLK(clk), .RST(1'b0), .Q(
        round_reg[929]) );
  DFF \round_reg_reg[930]  ( .D(N942), .CLK(clk), .RST(1'b0), .Q(
        round_reg[930]) );
  DFF \round_reg_reg[931]  ( .D(N943), .CLK(clk), .RST(1'b0), .Q(
        round_reg[931]) );
  DFF \round_reg_reg[932]  ( .D(N944), .CLK(clk), .RST(1'b0), .Q(
        round_reg[932]) );
  DFF \round_reg_reg[933]  ( .D(N945), .CLK(clk), .RST(1'b0), .Q(
        round_reg[933]) );
  DFF \round_reg_reg[934]  ( .D(N946), .CLK(clk), .RST(1'b0), .Q(
        round_reg[934]) );
  DFF \round_reg_reg[935]  ( .D(N947), .CLK(clk), .RST(1'b0), .Q(
        round_reg[935]) );
  DFF \round_reg_reg[936]  ( .D(N948), .CLK(clk), .RST(1'b0), .Q(
        round_reg[936]) );
  DFF \round_reg_reg[937]  ( .D(N949), .CLK(clk), .RST(1'b0), .Q(
        round_reg[937]) );
  DFF \round_reg_reg[938]  ( .D(N950), .CLK(clk), .RST(1'b0), .Q(
        round_reg[938]) );
  DFF \round_reg_reg[939]  ( .D(N951), .CLK(clk), .RST(1'b0), .Q(
        round_reg[939]) );
  DFF \round_reg_reg[940]  ( .D(N952), .CLK(clk), .RST(1'b0), .Q(
        round_reg[940]) );
  DFF \round_reg_reg[941]  ( .D(N953), .CLK(clk), .RST(1'b0), .Q(
        round_reg[941]) );
  DFF \round_reg_reg[942]  ( .D(N954), .CLK(clk), .RST(1'b0), .Q(
        round_reg[942]) );
  DFF \round_reg_reg[943]  ( .D(N955), .CLK(clk), .RST(1'b0), .Q(
        round_reg[943]) );
  DFF \round_reg_reg[944]  ( .D(N956), .CLK(clk), .RST(1'b0), .Q(
        round_reg[944]) );
  DFF \round_reg_reg[945]  ( .D(N957), .CLK(clk), .RST(1'b0), .Q(
        round_reg[945]) );
  DFF \round_reg_reg[946]  ( .D(N958), .CLK(clk), .RST(1'b0), .Q(
        round_reg[946]) );
  DFF \round_reg_reg[947]  ( .D(N959), .CLK(clk), .RST(1'b0), .Q(
        round_reg[947]) );
  DFF \round_reg_reg[948]  ( .D(N960), .CLK(clk), .RST(1'b0), .Q(
        round_reg[948]) );
  DFF \round_reg_reg[949]  ( .D(N961), .CLK(clk), .RST(1'b0), .Q(
        round_reg[949]) );
  DFF \round_reg_reg[950]  ( .D(N962), .CLK(clk), .RST(1'b0), .Q(
        round_reg[950]) );
  DFF \round_reg_reg[951]  ( .D(N963), .CLK(clk), .RST(1'b0), .Q(
        round_reg[951]) );
  DFF \round_reg_reg[952]  ( .D(N964), .CLK(clk), .RST(1'b0), .Q(
        round_reg[952]) );
  DFF \round_reg_reg[953]  ( .D(N965), .CLK(clk), .RST(1'b0), .Q(
        round_reg[953]) );
  DFF \round_reg_reg[954]  ( .D(N966), .CLK(clk), .RST(1'b0), .Q(
        round_reg[954]) );
  DFF \round_reg_reg[955]  ( .D(N967), .CLK(clk), .RST(1'b0), .Q(
        round_reg[955]) );
  DFF \round_reg_reg[956]  ( .D(N968), .CLK(clk), .RST(1'b0), .Q(
        round_reg[956]) );
  DFF \round_reg_reg[957]  ( .D(N969), .CLK(clk), .RST(1'b0), .Q(
        round_reg[957]) );
  DFF \round_reg_reg[958]  ( .D(N970), .CLK(clk), .RST(1'b0), .Q(
        round_reg[958]) );
  DFF \round_reg_reg[959]  ( .D(N971), .CLK(clk), .RST(1'b0), .Q(
        round_reg[959]) );
  DFF \round_reg_reg[960]  ( .D(N972), .CLK(clk), .RST(1'b0), .Q(
        round_reg[960]) );
  DFF \round_reg_reg[961]  ( .D(N973), .CLK(clk), .RST(1'b0), .Q(
        round_reg[961]) );
  DFF \round_reg_reg[962]  ( .D(N974), .CLK(clk), .RST(1'b0), .Q(
        round_reg[962]) );
  DFF \round_reg_reg[963]  ( .D(N975), .CLK(clk), .RST(1'b0), .Q(
        round_reg[963]) );
  DFF \round_reg_reg[964]  ( .D(N976), .CLK(clk), .RST(1'b0), .Q(
        round_reg[964]) );
  DFF \round_reg_reg[965]  ( .D(N977), .CLK(clk), .RST(1'b0), .Q(
        round_reg[965]) );
  DFF \round_reg_reg[966]  ( .D(N978), .CLK(clk), .RST(1'b0), .Q(
        round_reg[966]) );
  DFF \round_reg_reg[967]  ( .D(N979), .CLK(clk), .RST(1'b0), .Q(
        round_reg[967]) );
  DFF \round_reg_reg[968]  ( .D(N980), .CLK(clk), .RST(1'b0), .Q(
        round_reg[968]) );
  DFF \round_reg_reg[969]  ( .D(N981), .CLK(clk), .RST(1'b0), .Q(
        round_reg[969]) );
  DFF \round_reg_reg[970]  ( .D(N982), .CLK(clk), .RST(1'b0), .Q(
        round_reg[970]) );
  DFF \round_reg_reg[971]  ( .D(N983), .CLK(clk), .RST(1'b0), .Q(
        round_reg[971]) );
  DFF \round_reg_reg[972]  ( .D(N984), .CLK(clk), .RST(1'b0), .Q(
        round_reg[972]) );
  DFF \round_reg_reg[973]  ( .D(N985), .CLK(clk), .RST(1'b0), .Q(
        round_reg[973]) );
  DFF \round_reg_reg[974]  ( .D(N986), .CLK(clk), .RST(1'b0), .Q(
        round_reg[974]) );
  DFF \round_reg_reg[975]  ( .D(N987), .CLK(clk), .RST(1'b0), .Q(
        round_reg[975]) );
  DFF \round_reg_reg[976]  ( .D(N988), .CLK(clk), .RST(1'b0), .Q(
        round_reg[976]) );
  DFF \round_reg_reg[977]  ( .D(N989), .CLK(clk), .RST(1'b0), .Q(
        round_reg[977]) );
  DFF \round_reg_reg[978]  ( .D(N990), .CLK(clk), .RST(1'b0), .Q(
        round_reg[978]) );
  DFF \round_reg_reg[979]  ( .D(N991), .CLK(clk), .RST(1'b0), .Q(
        round_reg[979]) );
  DFF \round_reg_reg[980]  ( .D(N992), .CLK(clk), .RST(1'b0), .Q(
        round_reg[980]) );
  DFF \round_reg_reg[981]  ( .D(N993), .CLK(clk), .RST(1'b0), .Q(
        round_reg[981]) );
  DFF \round_reg_reg[982]  ( .D(N994), .CLK(clk), .RST(1'b0), .Q(
        round_reg[982]) );
  DFF \round_reg_reg[983]  ( .D(N995), .CLK(clk), .RST(1'b0), .Q(
        round_reg[983]) );
  DFF \round_reg_reg[984]  ( .D(N996), .CLK(clk), .RST(1'b0), .Q(
        round_reg[984]) );
  DFF \round_reg_reg[985]  ( .D(N997), .CLK(clk), .RST(1'b0), .Q(
        round_reg[985]) );
  DFF \round_reg_reg[986]  ( .D(N998), .CLK(clk), .RST(1'b0), .Q(
        round_reg[986]) );
  DFF \round_reg_reg[987]  ( .D(N999), .CLK(clk), .RST(1'b0), .Q(
        round_reg[987]) );
  DFF \round_reg_reg[988]  ( .D(N1000), .CLK(clk), .RST(1'b0), .Q(
        round_reg[988]) );
  DFF \round_reg_reg[989]  ( .D(N1001), .CLK(clk), .RST(1'b0), .Q(
        round_reg[989]) );
  DFF \round_reg_reg[990]  ( .D(N1002), .CLK(clk), .RST(1'b0), .Q(
        round_reg[990]) );
  DFF \round_reg_reg[991]  ( .D(N1003), .CLK(clk), .RST(1'b0), .Q(
        round_reg[991]) );
  DFF \round_reg_reg[992]  ( .D(N1004), .CLK(clk), .RST(1'b0), .Q(
        round_reg[992]) );
  DFF \round_reg_reg[993]  ( .D(N1005), .CLK(clk), .RST(1'b0), .Q(
        round_reg[993]) );
  DFF \round_reg_reg[994]  ( .D(N1006), .CLK(clk), .RST(1'b0), .Q(
        round_reg[994]) );
  DFF \round_reg_reg[995]  ( .D(N1007), .CLK(clk), .RST(1'b0), .Q(
        round_reg[995]) );
  DFF \round_reg_reg[996]  ( .D(N1008), .CLK(clk), .RST(1'b0), .Q(
        round_reg[996]) );
  DFF \round_reg_reg[997]  ( .D(N1009), .CLK(clk), .RST(1'b0), .Q(
        round_reg[997]) );
  DFF \round_reg_reg[998]  ( .D(N1010), .CLK(clk), .RST(1'b0), .Q(
        round_reg[998]) );
  DFF \round_reg_reg[999]  ( .D(N1011), .CLK(clk), .RST(1'b0), .Q(
        round_reg[999]) );
  DFF \round_reg_reg[1000]  ( .D(N1012), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1000]) );
  DFF \round_reg_reg[1001]  ( .D(N1013), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1001]) );
  DFF \round_reg_reg[1002]  ( .D(N1014), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1002]) );
  DFF \round_reg_reg[1003]  ( .D(N1015), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1003]) );
  DFF \round_reg_reg[1004]  ( .D(N1016), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1004]) );
  DFF \round_reg_reg[1005]  ( .D(N1017), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1005]) );
  DFF \round_reg_reg[1006]  ( .D(N1018), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1006]) );
  DFF \round_reg_reg[1007]  ( .D(N1019), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1007]) );
  DFF \round_reg_reg[1008]  ( .D(N1020), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1008]) );
  DFF \round_reg_reg[1009]  ( .D(N1021), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1009]) );
  DFF \round_reg_reg[1010]  ( .D(N1022), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1010]) );
  DFF \round_reg_reg[1011]  ( .D(N1023), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1011]) );
  DFF \round_reg_reg[1012]  ( .D(N1024), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1012]) );
  DFF \round_reg_reg[1013]  ( .D(N1025), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1013]) );
  DFF \round_reg_reg[1014]  ( .D(N1026), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1014]) );
  DFF \round_reg_reg[1015]  ( .D(N1027), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1015]) );
  DFF \round_reg_reg[1016]  ( .D(N1028), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1016]) );
  DFF \round_reg_reg[1017]  ( .D(N1029), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1017]) );
  DFF \round_reg_reg[1018]  ( .D(N1030), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1018]) );
  DFF \round_reg_reg[1019]  ( .D(N1031), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1019]) );
  DFF \round_reg_reg[1020]  ( .D(N1032), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1020]) );
  DFF \round_reg_reg[1021]  ( .D(N1033), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1021]) );
  DFF \round_reg_reg[1022]  ( .D(N1034), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1022]) );
  DFF \round_reg_reg[1023]  ( .D(N1035), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1023]) );
  DFF \round_reg_reg[1024]  ( .D(N1036), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1024]) );
  DFF \round_reg_reg[1025]  ( .D(N1037), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1025]) );
  DFF \round_reg_reg[1026]  ( .D(N1038), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1026]) );
  DFF \round_reg_reg[1027]  ( .D(N1039), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1027]) );
  DFF \round_reg_reg[1028]  ( .D(N1040), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1028]) );
  DFF \round_reg_reg[1029]  ( .D(N1041), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1029]) );
  DFF \round_reg_reg[1030]  ( .D(N1042), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1030]) );
  DFF \round_reg_reg[1031]  ( .D(N1043), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1031]) );
  DFF \round_reg_reg[1032]  ( .D(N1044), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1032]) );
  DFF \round_reg_reg[1033]  ( .D(N1045), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1033]) );
  DFF \round_reg_reg[1034]  ( .D(N1046), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1034]) );
  DFF \round_reg_reg[1035]  ( .D(N1047), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1035]) );
  DFF \round_reg_reg[1036]  ( .D(N1048), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1036]) );
  DFF \round_reg_reg[1037]  ( .D(N1049), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1037]) );
  DFF \round_reg_reg[1038]  ( .D(N1050), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1038]) );
  DFF \round_reg_reg[1039]  ( .D(N1051), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1039]) );
  DFF \round_reg_reg[1040]  ( .D(N1052), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1040]) );
  DFF \round_reg_reg[1041]  ( .D(N1053), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1041]) );
  DFF \round_reg_reg[1042]  ( .D(N1054), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1042]) );
  DFF \round_reg_reg[1043]  ( .D(N1055), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1043]) );
  DFF \round_reg_reg[1044]  ( .D(N1056), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1044]) );
  DFF \round_reg_reg[1045]  ( .D(N1057), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1045]) );
  DFF \round_reg_reg[1046]  ( .D(N1058), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1046]) );
  DFF \round_reg_reg[1047]  ( .D(N1059), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1047]) );
  DFF \round_reg_reg[1048]  ( .D(N1060), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1048]) );
  DFF \round_reg_reg[1049]  ( .D(N1061), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1049]) );
  DFF \round_reg_reg[1050]  ( .D(N1062), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1050]) );
  DFF \round_reg_reg[1051]  ( .D(N1063), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1051]) );
  DFF \round_reg_reg[1052]  ( .D(N1064), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1052]) );
  DFF \round_reg_reg[1053]  ( .D(N1065), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1053]) );
  DFF \round_reg_reg[1054]  ( .D(N1066), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1054]) );
  DFF \round_reg_reg[1055]  ( .D(N1067), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1055]) );
  DFF \round_reg_reg[1056]  ( .D(N1068), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1056]) );
  DFF \round_reg_reg[1057]  ( .D(N1069), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1057]) );
  DFF \round_reg_reg[1058]  ( .D(N1070), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1058]) );
  DFF \round_reg_reg[1059]  ( .D(N1071), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1059]) );
  DFF \round_reg_reg[1060]  ( .D(N1072), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1060]) );
  DFF \round_reg_reg[1061]  ( .D(N1073), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1061]) );
  DFF \round_reg_reg[1062]  ( .D(N1074), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1062]) );
  DFF \round_reg_reg[1063]  ( .D(N1075), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1063]) );
  DFF \round_reg_reg[1064]  ( .D(N1076), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1064]) );
  DFF \round_reg_reg[1065]  ( .D(N1077), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1065]) );
  DFF \round_reg_reg[1066]  ( .D(N1078), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1066]) );
  DFF \round_reg_reg[1067]  ( .D(N1079), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1067]) );
  DFF \round_reg_reg[1068]  ( .D(N1080), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1068]) );
  DFF \round_reg_reg[1069]  ( .D(N1081), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1069]) );
  DFF \round_reg_reg[1070]  ( .D(N1082), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1070]) );
  DFF \round_reg_reg[1071]  ( .D(N1083), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1071]) );
  DFF \round_reg_reg[1072]  ( .D(N1084), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1072]) );
  DFF \round_reg_reg[1073]  ( .D(N1085), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1073]) );
  DFF \round_reg_reg[1074]  ( .D(N1086), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1074]) );
  DFF \round_reg_reg[1075]  ( .D(N1087), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1075]) );
  DFF \round_reg_reg[1076]  ( .D(N1088), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1076]) );
  DFF \round_reg_reg[1077]  ( .D(N1089), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1077]) );
  DFF \round_reg_reg[1078]  ( .D(N1090), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1078]) );
  DFF \round_reg_reg[1079]  ( .D(N1091), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1079]) );
  DFF \round_reg_reg[1080]  ( .D(N1092), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1080]) );
  DFF \round_reg_reg[1081]  ( .D(N1093), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1081]) );
  DFF \round_reg_reg[1082]  ( .D(N1094), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1082]) );
  DFF \round_reg_reg[1083]  ( .D(N1095), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1083]) );
  DFF \round_reg_reg[1084]  ( .D(N1096), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1084]) );
  DFF \round_reg_reg[1085]  ( .D(N1097), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1085]) );
  DFF \round_reg_reg[1086]  ( .D(N1098), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1086]) );
  DFF \round_reg_reg[1087]  ( .D(N1099), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1087]) );
  DFF \round_reg_reg[1088]  ( .D(N1100), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1088]) );
  DFF \round_reg_reg[1089]  ( .D(N1101), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1089]) );
  DFF \round_reg_reg[1090]  ( .D(N1102), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1090]) );
  DFF \round_reg_reg[1091]  ( .D(N1103), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1091]) );
  DFF \round_reg_reg[1092]  ( .D(N1104), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1092]) );
  DFF \round_reg_reg[1093]  ( .D(N1105), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1093]) );
  DFF \round_reg_reg[1094]  ( .D(N1106), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1094]) );
  DFF \round_reg_reg[1095]  ( .D(N1107), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1095]) );
  DFF \round_reg_reg[1096]  ( .D(N1108), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1096]) );
  DFF \round_reg_reg[1097]  ( .D(N1109), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1097]) );
  DFF \round_reg_reg[1098]  ( .D(N1110), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1098]) );
  DFF \round_reg_reg[1099]  ( .D(N1111), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1099]) );
  DFF \round_reg_reg[1100]  ( .D(N1112), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1100]) );
  DFF \round_reg_reg[1101]  ( .D(N1113), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1101]) );
  DFF \round_reg_reg[1102]  ( .D(N1114), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1102]) );
  DFF \round_reg_reg[1103]  ( .D(N1115), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1103]) );
  DFF \round_reg_reg[1104]  ( .D(N1116), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1104]) );
  DFF \round_reg_reg[1105]  ( .D(N1117), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1105]) );
  DFF \round_reg_reg[1106]  ( .D(N1118), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1106]) );
  DFF \round_reg_reg[1107]  ( .D(N1119), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1107]) );
  DFF \round_reg_reg[1108]  ( .D(N1120), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1108]) );
  DFF \round_reg_reg[1109]  ( .D(N1121), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1109]) );
  DFF \round_reg_reg[1110]  ( .D(N1122), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1110]) );
  DFF \round_reg_reg[1111]  ( .D(N1123), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1111]) );
  DFF \round_reg_reg[1112]  ( .D(N1124), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1112]) );
  DFF \round_reg_reg[1113]  ( .D(N1125), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1113]) );
  DFF \round_reg_reg[1114]  ( .D(N1126), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1114]) );
  DFF \round_reg_reg[1115]  ( .D(N1127), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1115]) );
  DFF \round_reg_reg[1116]  ( .D(N1128), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1116]) );
  DFF \round_reg_reg[1117]  ( .D(N1129), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1117]) );
  DFF \round_reg_reg[1118]  ( .D(N1130), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1118]) );
  DFF \round_reg_reg[1119]  ( .D(N1131), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1119]) );
  DFF \round_reg_reg[1120]  ( .D(N1132), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1120]) );
  DFF \round_reg_reg[1121]  ( .D(N1133), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1121]) );
  DFF \round_reg_reg[1122]  ( .D(N1134), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1122]) );
  DFF \round_reg_reg[1123]  ( .D(N1135), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1123]) );
  DFF \round_reg_reg[1124]  ( .D(N1136), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1124]) );
  DFF \round_reg_reg[1125]  ( .D(N1137), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1125]) );
  DFF \round_reg_reg[1126]  ( .D(N1138), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1126]) );
  DFF \round_reg_reg[1127]  ( .D(N1139), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1127]) );
  DFF \round_reg_reg[1128]  ( .D(N1140), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1128]) );
  DFF \round_reg_reg[1129]  ( .D(N1141), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1129]) );
  DFF \round_reg_reg[1130]  ( .D(N1142), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1130]) );
  DFF \round_reg_reg[1131]  ( .D(N1143), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1131]) );
  DFF \round_reg_reg[1132]  ( .D(N1144), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1132]) );
  DFF \round_reg_reg[1133]  ( .D(N1145), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1133]) );
  DFF \round_reg_reg[1134]  ( .D(N1146), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1134]) );
  DFF \round_reg_reg[1135]  ( .D(N1147), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1135]) );
  DFF \round_reg_reg[1136]  ( .D(N1148), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1136]) );
  DFF \round_reg_reg[1137]  ( .D(N1149), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1137]) );
  DFF \round_reg_reg[1138]  ( .D(N1150), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1138]) );
  DFF \round_reg_reg[1139]  ( .D(N1151), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1139]) );
  DFF \round_reg_reg[1140]  ( .D(N1152), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1140]) );
  DFF \round_reg_reg[1141]  ( .D(N1153), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1141]) );
  DFF \round_reg_reg[1142]  ( .D(N1154), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1142]) );
  DFF \round_reg_reg[1143]  ( .D(N1155), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1143]) );
  DFF \round_reg_reg[1144]  ( .D(N1156), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1144]) );
  DFF \round_reg_reg[1145]  ( .D(N1157), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1145]) );
  DFF \round_reg_reg[1146]  ( .D(N1158), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1146]) );
  DFF \round_reg_reg[1147]  ( .D(N1159), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1147]) );
  DFF \round_reg_reg[1148]  ( .D(N1160), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1148]) );
  DFF \round_reg_reg[1149]  ( .D(N1161), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1149]) );
  DFF \round_reg_reg[1150]  ( .D(N1162), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1150]) );
  DFF \round_reg_reg[1151]  ( .D(N1163), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1151]) );
  DFF \round_reg_reg[1152]  ( .D(N1164), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1152]) );
  DFF \round_reg_reg[1153]  ( .D(N1165), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1153]) );
  DFF \round_reg_reg[1154]  ( .D(N1166), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1154]) );
  DFF \round_reg_reg[1155]  ( .D(N1167), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1155]) );
  DFF \round_reg_reg[1156]  ( .D(N1168), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1156]) );
  DFF \round_reg_reg[1157]  ( .D(N1169), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1157]) );
  DFF \round_reg_reg[1158]  ( .D(N1170), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1158]) );
  DFF \round_reg_reg[1159]  ( .D(N1171), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1159]) );
  DFF \round_reg_reg[1160]  ( .D(N1172), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1160]) );
  DFF \round_reg_reg[1161]  ( .D(N1173), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1161]) );
  DFF \round_reg_reg[1162]  ( .D(N1174), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1162]) );
  DFF \round_reg_reg[1163]  ( .D(N1175), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1163]) );
  DFF \round_reg_reg[1164]  ( .D(N1176), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1164]) );
  DFF \round_reg_reg[1165]  ( .D(N1177), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1165]) );
  DFF \round_reg_reg[1166]  ( .D(N1178), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1166]) );
  DFF \round_reg_reg[1167]  ( .D(N1179), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1167]) );
  DFF \round_reg_reg[1168]  ( .D(N1180), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1168]) );
  DFF \round_reg_reg[1169]  ( .D(N1181), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1169]) );
  DFF \round_reg_reg[1170]  ( .D(N1182), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1170]) );
  DFF \round_reg_reg[1171]  ( .D(N1183), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1171]) );
  DFF \round_reg_reg[1172]  ( .D(N1184), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1172]) );
  DFF \round_reg_reg[1173]  ( .D(N1185), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1173]) );
  DFF \round_reg_reg[1174]  ( .D(N1186), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1174]) );
  DFF \round_reg_reg[1175]  ( .D(N1187), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1175]) );
  DFF \round_reg_reg[1176]  ( .D(N1188), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1176]) );
  DFF \round_reg_reg[1177]  ( .D(N1189), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1177]) );
  DFF \round_reg_reg[1178]  ( .D(N1190), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1178]) );
  DFF \round_reg_reg[1179]  ( .D(N1191), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1179]) );
  DFF \round_reg_reg[1180]  ( .D(N1192), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1180]) );
  DFF \round_reg_reg[1181]  ( .D(N1193), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1181]) );
  DFF \round_reg_reg[1182]  ( .D(N1194), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1182]) );
  DFF \round_reg_reg[1183]  ( .D(N1195), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1183]) );
  DFF \round_reg_reg[1184]  ( .D(N1196), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1184]) );
  DFF \round_reg_reg[1185]  ( .D(N1197), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1185]) );
  DFF \round_reg_reg[1186]  ( .D(N1198), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1186]) );
  DFF \round_reg_reg[1187]  ( .D(N1199), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1187]) );
  DFF \round_reg_reg[1188]  ( .D(N1200), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1188]) );
  DFF \round_reg_reg[1189]  ( .D(N1201), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1189]) );
  DFF \round_reg_reg[1190]  ( .D(N1202), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1190]) );
  DFF \round_reg_reg[1191]  ( .D(N1203), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1191]) );
  DFF \round_reg_reg[1192]  ( .D(N1204), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1192]) );
  DFF \round_reg_reg[1193]  ( .D(N1205), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1193]) );
  DFF \round_reg_reg[1194]  ( .D(N1206), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1194]) );
  DFF \round_reg_reg[1195]  ( .D(N1207), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1195]) );
  DFF \round_reg_reg[1196]  ( .D(N1208), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1196]) );
  DFF \round_reg_reg[1197]  ( .D(N1209), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1197]) );
  DFF \round_reg_reg[1198]  ( .D(N1210), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1198]) );
  DFF \round_reg_reg[1199]  ( .D(N1211), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1199]) );
  DFF \round_reg_reg[1200]  ( .D(N1212), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1200]) );
  DFF \round_reg_reg[1201]  ( .D(N1213), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1201]) );
  DFF \round_reg_reg[1202]  ( .D(N1214), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1202]) );
  DFF \round_reg_reg[1203]  ( .D(N1215), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1203]) );
  DFF \round_reg_reg[1204]  ( .D(N1216), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1204]) );
  DFF \round_reg_reg[1205]  ( .D(N1217), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1205]) );
  DFF \round_reg_reg[1206]  ( .D(N1218), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1206]) );
  DFF \round_reg_reg[1207]  ( .D(N1219), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1207]) );
  DFF \round_reg_reg[1208]  ( .D(N1220), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1208]) );
  DFF \round_reg_reg[1209]  ( .D(N1221), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1209]) );
  DFF \round_reg_reg[1210]  ( .D(N1222), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1210]) );
  DFF \round_reg_reg[1211]  ( .D(N1223), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1211]) );
  DFF \round_reg_reg[1212]  ( .D(N1224), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1212]) );
  DFF \round_reg_reg[1213]  ( .D(N1225), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1213]) );
  DFF \round_reg_reg[1214]  ( .D(N1226), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1214]) );
  DFF \round_reg_reg[1215]  ( .D(N1227), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1215]) );
  DFF \round_reg_reg[1216]  ( .D(N1228), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1216]) );
  DFF \round_reg_reg[1217]  ( .D(N1229), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1217]) );
  DFF \round_reg_reg[1218]  ( .D(N1230), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1218]) );
  DFF \round_reg_reg[1219]  ( .D(N1231), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1219]) );
  DFF \round_reg_reg[1220]  ( .D(N1232), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1220]) );
  DFF \round_reg_reg[1221]  ( .D(N1233), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1221]) );
  DFF \round_reg_reg[1222]  ( .D(N1234), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1222]) );
  DFF \round_reg_reg[1223]  ( .D(N1235), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1223]) );
  DFF \round_reg_reg[1224]  ( .D(N1236), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1224]) );
  DFF \round_reg_reg[1225]  ( .D(N1237), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1225]) );
  DFF \round_reg_reg[1226]  ( .D(N1238), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1226]) );
  DFF \round_reg_reg[1227]  ( .D(N1239), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1227]) );
  DFF \round_reg_reg[1228]  ( .D(N1240), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1228]) );
  DFF \round_reg_reg[1229]  ( .D(N1241), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1229]) );
  DFF \round_reg_reg[1230]  ( .D(N1242), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1230]) );
  DFF \round_reg_reg[1231]  ( .D(N1243), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1231]) );
  DFF \round_reg_reg[1232]  ( .D(N1244), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1232]) );
  DFF \round_reg_reg[1233]  ( .D(N1245), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1233]) );
  DFF \round_reg_reg[1234]  ( .D(N1246), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1234]) );
  DFF \round_reg_reg[1235]  ( .D(N1247), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1235]) );
  DFF \round_reg_reg[1236]  ( .D(N1248), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1236]) );
  DFF \round_reg_reg[1237]  ( .D(N1249), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1237]) );
  DFF \round_reg_reg[1238]  ( .D(N1250), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1238]) );
  DFF \round_reg_reg[1239]  ( .D(N1251), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1239]) );
  DFF \round_reg_reg[1240]  ( .D(N1252), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1240]) );
  DFF \round_reg_reg[1241]  ( .D(N1253), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1241]) );
  DFF \round_reg_reg[1242]  ( .D(N1254), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1242]) );
  DFF \round_reg_reg[1243]  ( .D(N1255), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1243]) );
  DFF \round_reg_reg[1244]  ( .D(N1256), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1244]) );
  DFF \round_reg_reg[1245]  ( .D(N1257), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1245]) );
  DFF \round_reg_reg[1246]  ( .D(N1258), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1246]) );
  DFF \round_reg_reg[1247]  ( .D(N1259), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1247]) );
  DFF \round_reg_reg[1248]  ( .D(N1260), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1248]) );
  DFF \round_reg_reg[1249]  ( .D(N1261), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1249]) );
  DFF \round_reg_reg[1250]  ( .D(N1262), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1250]) );
  DFF \round_reg_reg[1251]  ( .D(N1263), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1251]) );
  DFF \round_reg_reg[1252]  ( .D(N1264), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1252]) );
  DFF \round_reg_reg[1253]  ( .D(N1265), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1253]) );
  DFF \round_reg_reg[1254]  ( .D(N1266), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1254]) );
  DFF \round_reg_reg[1255]  ( .D(N1267), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1255]) );
  DFF \round_reg_reg[1256]  ( .D(N1268), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1256]) );
  DFF \round_reg_reg[1257]  ( .D(N1269), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1257]) );
  DFF \round_reg_reg[1258]  ( .D(N1270), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1258]) );
  DFF \round_reg_reg[1259]  ( .D(N1271), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1259]) );
  DFF \round_reg_reg[1260]  ( .D(N1272), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1260]) );
  DFF \round_reg_reg[1261]  ( .D(N1273), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1261]) );
  DFF \round_reg_reg[1262]  ( .D(N1274), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1262]) );
  DFF \round_reg_reg[1263]  ( .D(N1275), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1263]) );
  DFF \round_reg_reg[1264]  ( .D(N1276), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1264]) );
  DFF \round_reg_reg[1265]  ( .D(N1277), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1265]) );
  DFF \round_reg_reg[1266]  ( .D(N1278), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1266]) );
  DFF \round_reg_reg[1267]  ( .D(N1279), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1267]) );
  DFF \round_reg_reg[1268]  ( .D(N1280), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1268]) );
  DFF \round_reg_reg[1269]  ( .D(N1281), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1269]) );
  DFF \round_reg_reg[1270]  ( .D(N1282), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1270]) );
  DFF \round_reg_reg[1271]  ( .D(N1283), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1271]) );
  DFF \round_reg_reg[1272]  ( .D(N1284), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1272]) );
  DFF \round_reg_reg[1273]  ( .D(N1285), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1273]) );
  DFF \round_reg_reg[1274]  ( .D(N1286), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1274]) );
  DFF \round_reg_reg[1275]  ( .D(N1287), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1275]) );
  DFF \round_reg_reg[1276]  ( .D(N1288), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1276]) );
  DFF \round_reg_reg[1277]  ( .D(N1289), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1277]) );
  DFF \round_reg_reg[1278]  ( .D(N1290), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1278]) );
  DFF \round_reg_reg[1279]  ( .D(N1291), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1279]) );
  DFF \round_reg_reg[1280]  ( .D(N1292), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1280]) );
  DFF \round_reg_reg[1281]  ( .D(N1293), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1281]) );
  DFF \round_reg_reg[1282]  ( .D(N1294), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1282]) );
  DFF \round_reg_reg[1283]  ( .D(N1295), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1283]) );
  DFF \round_reg_reg[1284]  ( .D(N1296), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1284]) );
  DFF \round_reg_reg[1285]  ( .D(N1297), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1285]) );
  DFF \round_reg_reg[1286]  ( .D(N1298), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1286]) );
  DFF \round_reg_reg[1287]  ( .D(N1299), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1287]) );
  DFF \round_reg_reg[1288]  ( .D(N1300), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1288]) );
  DFF \round_reg_reg[1289]  ( .D(N1301), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1289]) );
  DFF \round_reg_reg[1290]  ( .D(N1302), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1290]) );
  DFF \round_reg_reg[1291]  ( .D(N1303), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1291]) );
  DFF \round_reg_reg[1292]  ( .D(N1304), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1292]) );
  DFF \round_reg_reg[1293]  ( .D(N1305), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1293]) );
  DFF \round_reg_reg[1294]  ( .D(N1306), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1294]) );
  DFF \round_reg_reg[1295]  ( .D(N1307), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1295]) );
  DFF \round_reg_reg[1296]  ( .D(N1308), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1296]) );
  DFF \round_reg_reg[1297]  ( .D(N1309), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1297]) );
  DFF \round_reg_reg[1298]  ( .D(N1310), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1298]) );
  DFF \round_reg_reg[1299]  ( .D(N1311), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1299]) );
  DFF \round_reg_reg[1300]  ( .D(N1312), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1300]) );
  DFF \round_reg_reg[1301]  ( .D(N1313), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1301]) );
  DFF \round_reg_reg[1302]  ( .D(N1314), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1302]) );
  DFF \round_reg_reg[1303]  ( .D(N1315), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1303]) );
  DFF \round_reg_reg[1304]  ( .D(N1316), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1304]) );
  DFF \round_reg_reg[1305]  ( .D(N1317), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1305]) );
  DFF \round_reg_reg[1306]  ( .D(N1318), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1306]) );
  DFF \round_reg_reg[1307]  ( .D(N1319), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1307]) );
  DFF \round_reg_reg[1308]  ( .D(N1320), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1308]) );
  DFF \round_reg_reg[1309]  ( .D(N1321), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1309]) );
  DFF \round_reg_reg[1310]  ( .D(N1322), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1310]) );
  DFF \round_reg_reg[1311]  ( .D(N1323), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1311]) );
  DFF \round_reg_reg[1312]  ( .D(N1324), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1312]) );
  DFF \round_reg_reg[1313]  ( .D(N1325), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1313]) );
  DFF \round_reg_reg[1314]  ( .D(N1326), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1314]) );
  DFF \round_reg_reg[1315]  ( .D(N1327), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1315]) );
  DFF \round_reg_reg[1316]  ( .D(N1328), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1316]) );
  DFF \round_reg_reg[1317]  ( .D(N1329), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1317]) );
  DFF \round_reg_reg[1318]  ( .D(N1330), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1318]) );
  DFF \round_reg_reg[1319]  ( .D(N1331), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1319]) );
  DFF \round_reg_reg[1320]  ( .D(N1332), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1320]) );
  DFF \round_reg_reg[1321]  ( .D(N1333), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1321]) );
  DFF \round_reg_reg[1322]  ( .D(N1334), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1322]) );
  DFF \round_reg_reg[1323]  ( .D(N1335), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1323]) );
  DFF \round_reg_reg[1324]  ( .D(N1336), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1324]) );
  DFF \round_reg_reg[1325]  ( .D(N1337), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1325]) );
  DFF \round_reg_reg[1326]  ( .D(N1338), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1326]) );
  DFF \round_reg_reg[1327]  ( .D(N1339), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1327]) );
  DFF \round_reg_reg[1328]  ( .D(N1340), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1328]) );
  DFF \round_reg_reg[1329]  ( .D(N1341), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1329]) );
  DFF \round_reg_reg[1330]  ( .D(N1342), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1330]) );
  DFF \round_reg_reg[1331]  ( .D(N1343), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1331]) );
  DFF \round_reg_reg[1332]  ( .D(N1344), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1332]) );
  DFF \round_reg_reg[1333]  ( .D(N1345), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1333]) );
  DFF \round_reg_reg[1334]  ( .D(N1346), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1334]) );
  DFF \round_reg_reg[1335]  ( .D(N1347), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1335]) );
  DFF \round_reg_reg[1336]  ( .D(N1348), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1336]) );
  DFF \round_reg_reg[1337]  ( .D(N1349), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1337]) );
  DFF \round_reg_reg[1338]  ( .D(N1350), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1338]) );
  DFF \round_reg_reg[1339]  ( .D(N1351), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1339]) );
  DFF \round_reg_reg[1340]  ( .D(N1352), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1340]) );
  DFF \round_reg_reg[1341]  ( .D(N1353), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1341]) );
  DFF \round_reg_reg[1342]  ( .D(N1354), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1342]) );
  DFF \round_reg_reg[1343]  ( .D(N1355), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1343]) );
  DFF \round_reg_reg[1344]  ( .D(N1356), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1344]) );
  DFF \round_reg_reg[1345]  ( .D(N1357), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1345]) );
  DFF \round_reg_reg[1346]  ( .D(N1358), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1346]) );
  DFF \round_reg_reg[1347]  ( .D(N1359), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1347]) );
  DFF \round_reg_reg[1348]  ( .D(N1360), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1348]) );
  DFF \round_reg_reg[1349]  ( .D(N1361), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1349]) );
  DFF \round_reg_reg[1350]  ( .D(N1362), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1350]) );
  DFF \round_reg_reg[1351]  ( .D(N1363), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1351]) );
  DFF \round_reg_reg[1352]  ( .D(N1364), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1352]) );
  DFF \round_reg_reg[1353]  ( .D(N1365), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1353]) );
  DFF \round_reg_reg[1354]  ( .D(N1366), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1354]) );
  DFF \round_reg_reg[1355]  ( .D(N1367), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1355]) );
  DFF \round_reg_reg[1356]  ( .D(N1368), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1356]) );
  DFF \round_reg_reg[1357]  ( .D(N1369), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1357]) );
  DFF \round_reg_reg[1358]  ( .D(N1370), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1358]) );
  DFF \round_reg_reg[1359]  ( .D(N1371), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1359]) );
  DFF \round_reg_reg[1360]  ( .D(N1372), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1360]) );
  DFF \round_reg_reg[1361]  ( .D(N1373), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1361]) );
  DFF \round_reg_reg[1362]  ( .D(N1374), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1362]) );
  DFF \round_reg_reg[1363]  ( .D(N1375), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1363]) );
  DFF \round_reg_reg[1364]  ( .D(N1376), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1364]) );
  DFF \round_reg_reg[1365]  ( .D(N1377), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1365]) );
  DFF \round_reg_reg[1366]  ( .D(N1378), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1366]) );
  DFF \round_reg_reg[1367]  ( .D(N1379), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1367]) );
  DFF \round_reg_reg[1368]  ( .D(N1380), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1368]) );
  DFF \round_reg_reg[1369]  ( .D(N1381), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1369]) );
  DFF \round_reg_reg[1370]  ( .D(N1382), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1370]) );
  DFF \round_reg_reg[1371]  ( .D(N1383), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1371]) );
  DFF \round_reg_reg[1372]  ( .D(N1384), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1372]) );
  DFF \round_reg_reg[1373]  ( .D(N1385), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1373]) );
  DFF \round_reg_reg[1374]  ( .D(N1386), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1374]) );
  DFF \round_reg_reg[1375]  ( .D(N1387), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1375]) );
  DFF \round_reg_reg[1376]  ( .D(N1388), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1376]) );
  DFF \round_reg_reg[1377]  ( .D(N1389), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1377]) );
  DFF \round_reg_reg[1378]  ( .D(N1390), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1378]) );
  DFF \round_reg_reg[1379]  ( .D(N1391), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1379]) );
  DFF \round_reg_reg[1380]  ( .D(N1392), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1380]) );
  DFF \round_reg_reg[1381]  ( .D(N1393), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1381]) );
  DFF \round_reg_reg[1382]  ( .D(N1394), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1382]) );
  DFF \round_reg_reg[1383]  ( .D(N1395), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1383]) );
  DFF \round_reg_reg[1384]  ( .D(N1396), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1384]) );
  DFF \round_reg_reg[1385]  ( .D(N1397), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1385]) );
  DFF \round_reg_reg[1386]  ( .D(N1398), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1386]) );
  DFF \round_reg_reg[1387]  ( .D(N1399), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1387]) );
  DFF \round_reg_reg[1388]  ( .D(N1400), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1388]) );
  DFF \round_reg_reg[1389]  ( .D(N1401), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1389]) );
  DFF \round_reg_reg[1390]  ( .D(N1402), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1390]) );
  DFF \round_reg_reg[1391]  ( .D(N1403), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1391]) );
  DFF \round_reg_reg[1392]  ( .D(N1404), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1392]) );
  DFF \round_reg_reg[1393]  ( .D(N1405), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1393]) );
  DFF \round_reg_reg[1394]  ( .D(N1406), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1394]) );
  DFF \round_reg_reg[1395]  ( .D(N1407), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1395]) );
  DFF \round_reg_reg[1396]  ( .D(N1408), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1396]) );
  DFF \round_reg_reg[1397]  ( .D(N1409), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1397]) );
  DFF \round_reg_reg[1398]  ( .D(N1410), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1398]) );
  DFF \round_reg_reg[1399]  ( .D(N1411), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1399]) );
  DFF \round_reg_reg[1400]  ( .D(N1412), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1400]) );
  DFF \round_reg_reg[1401]  ( .D(N1413), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1401]) );
  DFF \round_reg_reg[1402]  ( .D(N1414), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1402]) );
  DFF \round_reg_reg[1403]  ( .D(N1415), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1403]) );
  DFF \round_reg_reg[1404]  ( .D(N1416), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1404]) );
  DFF \round_reg_reg[1405]  ( .D(N1417), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1405]) );
  DFF \round_reg_reg[1406]  ( .D(N1418), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1406]) );
  DFF \round_reg_reg[1407]  ( .D(N1419), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1407]) );
  DFF \round_reg_reg[1408]  ( .D(N1420), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1408]) );
  DFF \round_reg_reg[1409]  ( .D(N1421), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1409]) );
  DFF \round_reg_reg[1410]  ( .D(N1422), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1410]) );
  DFF \round_reg_reg[1411]  ( .D(N1423), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1411]) );
  DFF \round_reg_reg[1412]  ( .D(N1424), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1412]) );
  DFF \round_reg_reg[1413]  ( .D(N1425), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1413]) );
  DFF \round_reg_reg[1414]  ( .D(N1426), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1414]) );
  DFF \round_reg_reg[1415]  ( .D(N1427), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1415]) );
  DFF \round_reg_reg[1416]  ( .D(N1428), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1416]) );
  DFF \round_reg_reg[1417]  ( .D(N1429), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1417]) );
  DFF \round_reg_reg[1418]  ( .D(N1430), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1418]) );
  DFF \round_reg_reg[1419]  ( .D(N1431), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1419]) );
  DFF \round_reg_reg[1420]  ( .D(N1432), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1420]) );
  DFF \round_reg_reg[1421]  ( .D(N1433), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1421]) );
  DFF \round_reg_reg[1422]  ( .D(N1434), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1422]) );
  DFF \round_reg_reg[1423]  ( .D(N1435), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1423]) );
  DFF \round_reg_reg[1424]  ( .D(N1436), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1424]) );
  DFF \round_reg_reg[1425]  ( .D(N1437), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1425]) );
  DFF \round_reg_reg[1426]  ( .D(N1438), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1426]) );
  DFF \round_reg_reg[1427]  ( .D(N1439), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1427]) );
  DFF \round_reg_reg[1428]  ( .D(N1440), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1428]) );
  DFF \round_reg_reg[1429]  ( .D(N1441), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1429]) );
  DFF \round_reg_reg[1430]  ( .D(N1442), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1430]) );
  DFF \round_reg_reg[1431]  ( .D(N1443), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1431]) );
  DFF \round_reg_reg[1432]  ( .D(N1444), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1432]) );
  DFF \round_reg_reg[1433]  ( .D(N1445), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1433]) );
  DFF \round_reg_reg[1434]  ( .D(N1446), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1434]) );
  DFF \round_reg_reg[1435]  ( .D(N1447), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1435]) );
  DFF \round_reg_reg[1436]  ( .D(N1448), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1436]) );
  DFF \round_reg_reg[1437]  ( .D(N1449), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1437]) );
  DFF \round_reg_reg[1438]  ( .D(N1450), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1438]) );
  DFF \round_reg_reg[1439]  ( .D(N1451), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1439]) );
  DFF \round_reg_reg[1440]  ( .D(N1452), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1440]) );
  DFF \round_reg_reg[1441]  ( .D(N1453), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1441]) );
  DFF \round_reg_reg[1442]  ( .D(N1454), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1442]) );
  DFF \round_reg_reg[1443]  ( .D(N1455), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1443]) );
  DFF \round_reg_reg[1444]  ( .D(N1456), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1444]) );
  DFF \round_reg_reg[1445]  ( .D(N1457), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1445]) );
  DFF \round_reg_reg[1446]  ( .D(N1458), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1446]) );
  DFF \round_reg_reg[1447]  ( .D(N1459), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1447]) );
  DFF \round_reg_reg[1448]  ( .D(N1460), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1448]) );
  DFF \round_reg_reg[1449]  ( .D(N1461), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1449]) );
  DFF \round_reg_reg[1450]  ( .D(N1462), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1450]) );
  DFF \round_reg_reg[1451]  ( .D(N1463), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1451]) );
  DFF \round_reg_reg[1452]  ( .D(N1464), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1452]) );
  DFF \round_reg_reg[1453]  ( .D(N1465), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1453]) );
  DFF \round_reg_reg[1454]  ( .D(N1466), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1454]) );
  DFF \round_reg_reg[1455]  ( .D(N1467), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1455]) );
  DFF \round_reg_reg[1456]  ( .D(N1468), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1456]) );
  DFF \round_reg_reg[1457]  ( .D(N1469), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1457]) );
  DFF \round_reg_reg[1458]  ( .D(N1470), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1458]) );
  DFF \round_reg_reg[1459]  ( .D(N1471), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1459]) );
  DFF \round_reg_reg[1460]  ( .D(N1472), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1460]) );
  DFF \round_reg_reg[1461]  ( .D(N1473), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1461]) );
  DFF \round_reg_reg[1462]  ( .D(N1474), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1462]) );
  DFF \round_reg_reg[1463]  ( .D(N1475), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1463]) );
  DFF \round_reg_reg[1464]  ( .D(N1476), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1464]) );
  DFF \round_reg_reg[1465]  ( .D(N1477), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1465]) );
  DFF \round_reg_reg[1466]  ( .D(N1478), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1466]) );
  DFF \round_reg_reg[1467]  ( .D(N1479), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1467]) );
  DFF \round_reg_reg[1468]  ( .D(N1480), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1468]) );
  DFF \round_reg_reg[1469]  ( .D(N1481), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1469]) );
  DFF \round_reg_reg[1470]  ( .D(N1482), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1470]) );
  DFF \round_reg_reg[1471]  ( .D(N1483), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1471]) );
  DFF \round_reg_reg[1472]  ( .D(N1484), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1472]) );
  DFF \round_reg_reg[1473]  ( .D(N1485), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1473]) );
  DFF \round_reg_reg[1474]  ( .D(N1486), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1474]) );
  DFF \round_reg_reg[1475]  ( .D(N1487), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1475]) );
  DFF \round_reg_reg[1476]  ( .D(N1488), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1476]) );
  DFF \round_reg_reg[1477]  ( .D(N1489), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1477]) );
  DFF \round_reg_reg[1478]  ( .D(N1490), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1478]) );
  DFF \round_reg_reg[1479]  ( .D(N1491), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1479]) );
  DFF \round_reg_reg[1480]  ( .D(N1492), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1480]) );
  DFF \round_reg_reg[1481]  ( .D(N1493), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1481]) );
  DFF \round_reg_reg[1482]  ( .D(N1494), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1482]) );
  DFF \round_reg_reg[1483]  ( .D(N1495), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1483]) );
  DFF \round_reg_reg[1484]  ( .D(N1496), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1484]) );
  DFF \round_reg_reg[1485]  ( .D(N1497), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1485]) );
  DFF \round_reg_reg[1486]  ( .D(N1498), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1486]) );
  DFF \round_reg_reg[1487]  ( .D(N1499), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1487]) );
  DFF \round_reg_reg[1488]  ( .D(N1500), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1488]) );
  DFF \round_reg_reg[1489]  ( .D(N1501), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1489]) );
  DFF \round_reg_reg[1490]  ( .D(N1502), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1490]) );
  DFF \round_reg_reg[1491]  ( .D(N1503), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1491]) );
  DFF \round_reg_reg[1492]  ( .D(N1504), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1492]) );
  DFF \round_reg_reg[1493]  ( .D(N1505), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1493]) );
  DFF \round_reg_reg[1494]  ( .D(N1506), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1494]) );
  DFF \round_reg_reg[1495]  ( .D(N1507), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1495]) );
  DFF \round_reg_reg[1496]  ( .D(N1508), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1496]) );
  DFF \round_reg_reg[1497]  ( .D(N1509), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1497]) );
  DFF \round_reg_reg[1498]  ( .D(N1510), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1498]) );
  DFF \round_reg_reg[1499]  ( .D(N1511), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1499]) );
  DFF \round_reg_reg[1500]  ( .D(N1512), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1500]) );
  DFF \round_reg_reg[1501]  ( .D(N1513), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1501]) );
  DFF \round_reg_reg[1502]  ( .D(N1514), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1502]) );
  DFF \round_reg_reg[1503]  ( .D(N1515), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1503]) );
  DFF \round_reg_reg[1504]  ( .D(N1516), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1504]) );
  DFF \round_reg_reg[1505]  ( .D(N1517), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1505]) );
  DFF \round_reg_reg[1506]  ( .D(N1518), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1506]) );
  DFF \round_reg_reg[1507]  ( .D(N1519), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1507]) );
  DFF \round_reg_reg[1508]  ( .D(N1520), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1508]) );
  DFF \round_reg_reg[1509]  ( .D(N1521), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1509]) );
  DFF \round_reg_reg[1510]  ( .D(N1522), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1510]) );
  DFF \round_reg_reg[1511]  ( .D(N1523), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1511]) );
  DFF \round_reg_reg[1512]  ( .D(N1524), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1512]) );
  DFF \round_reg_reg[1513]  ( .D(N1525), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1513]) );
  DFF \round_reg_reg[1514]  ( .D(N1526), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1514]) );
  DFF \round_reg_reg[1515]  ( .D(N1527), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1515]) );
  DFF \round_reg_reg[1516]  ( .D(N1528), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1516]) );
  DFF \round_reg_reg[1517]  ( .D(N1529), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1517]) );
  DFF \round_reg_reg[1518]  ( .D(N1530), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1518]) );
  DFF \round_reg_reg[1519]  ( .D(N1531), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1519]) );
  DFF \round_reg_reg[1520]  ( .D(N1532), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1520]) );
  DFF \round_reg_reg[1521]  ( .D(N1533), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1521]) );
  DFF \round_reg_reg[1522]  ( .D(N1534), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1522]) );
  DFF \round_reg_reg[1523]  ( .D(N1535), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1523]) );
  DFF \round_reg_reg[1524]  ( .D(N1536), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1524]) );
  DFF \round_reg_reg[1525]  ( .D(N1537), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1525]) );
  DFF \round_reg_reg[1526]  ( .D(N1538), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1526]) );
  DFF \round_reg_reg[1527]  ( .D(N1539), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1527]) );
  DFF \round_reg_reg[1528]  ( .D(N1540), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1528]) );
  DFF \round_reg_reg[1529]  ( .D(N1541), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1529]) );
  DFF \round_reg_reg[1530]  ( .D(N1542), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1530]) );
  DFF \round_reg_reg[1531]  ( .D(N1543), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1531]) );
  DFF \round_reg_reg[1532]  ( .D(N1544), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1532]) );
  DFF \round_reg_reg[1533]  ( .D(N1545), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1533]) );
  DFF \round_reg_reg[1534]  ( .D(N1546), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1534]) );
  DFF \round_reg_reg[1535]  ( .D(N1547), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1535]) );
  DFF \round_reg_reg[1536]  ( .D(N1548), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1536]) );
  DFF \round_reg_reg[1537]  ( .D(N1549), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1537]) );
  DFF \round_reg_reg[1538]  ( .D(N1550), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1538]) );
  DFF \round_reg_reg[1539]  ( .D(N1551), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1539]) );
  DFF \round_reg_reg[1540]  ( .D(N1552), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1540]) );
  DFF \round_reg_reg[1541]  ( .D(N1553), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1541]) );
  DFF \round_reg_reg[1542]  ( .D(N1554), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1542]) );
  DFF \round_reg_reg[1543]  ( .D(N1555), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1543]) );
  DFF \round_reg_reg[1544]  ( .D(N1556), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1544]) );
  DFF \round_reg_reg[1545]  ( .D(N1557), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1545]) );
  DFF \round_reg_reg[1546]  ( .D(N1558), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1546]) );
  DFF \round_reg_reg[1547]  ( .D(N1559), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1547]) );
  DFF \round_reg_reg[1548]  ( .D(N1560), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1548]) );
  DFF \round_reg_reg[1549]  ( .D(N1561), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1549]) );
  DFF \round_reg_reg[1550]  ( .D(N1562), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1550]) );
  DFF \round_reg_reg[1551]  ( .D(N1563), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1551]) );
  DFF \round_reg_reg[1552]  ( .D(N1564), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1552]) );
  DFF \round_reg_reg[1553]  ( .D(N1565), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1553]) );
  DFF \round_reg_reg[1554]  ( .D(N1566), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1554]) );
  DFF \round_reg_reg[1555]  ( .D(N1567), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1555]) );
  DFF \round_reg_reg[1556]  ( .D(N1568), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1556]) );
  DFF \round_reg_reg[1557]  ( .D(N1569), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1557]) );
  DFF \round_reg_reg[1558]  ( .D(N1570), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1558]) );
  DFF \round_reg_reg[1559]  ( .D(N1571), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1559]) );
  DFF \round_reg_reg[1560]  ( .D(N1572), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1560]) );
  DFF \round_reg_reg[1561]  ( .D(N1573), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1561]) );
  DFF \round_reg_reg[1562]  ( .D(N1574), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1562]) );
  DFF \round_reg_reg[1563]  ( .D(N1575), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1563]) );
  DFF \round_reg_reg[1564]  ( .D(N1576), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1564]) );
  DFF \round_reg_reg[1565]  ( .D(N1577), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1565]) );
  DFF \round_reg_reg[1566]  ( .D(N1578), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1566]) );
  DFF \round_reg_reg[1567]  ( .D(N1579), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1567]) );
  DFF \round_reg_reg[1568]  ( .D(N1580), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1568]) );
  DFF \round_reg_reg[1569]  ( .D(N1581), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1569]) );
  DFF \round_reg_reg[1570]  ( .D(N1582), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1570]) );
  DFF \round_reg_reg[1571]  ( .D(N1583), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1571]) );
  DFF \round_reg_reg[1572]  ( .D(N1584), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1572]) );
  DFF \round_reg_reg[1573]  ( .D(N1585), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1573]) );
  DFF \round_reg_reg[1574]  ( .D(N1586), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1574]) );
  DFF \round_reg_reg[1575]  ( .D(N1587), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1575]) );
  DFF \round_reg_reg[1576]  ( .D(N1588), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1576]) );
  DFF \round_reg_reg[1577]  ( .D(N1589), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1577]) );
  DFF \round_reg_reg[1578]  ( .D(N1590), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1578]) );
  DFF \round_reg_reg[1579]  ( .D(N1591), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1579]) );
  DFF \round_reg_reg[1580]  ( .D(N1592), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1580]) );
  DFF \round_reg_reg[1581]  ( .D(N1593), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1581]) );
  DFF \round_reg_reg[1582]  ( .D(N1594), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1582]) );
  DFF \round_reg_reg[1583]  ( .D(N1595), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1583]) );
  DFF \round_reg_reg[1584]  ( .D(N1596), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1584]) );
  DFF \round_reg_reg[1585]  ( .D(N1597), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1585]) );
  DFF \round_reg_reg[1586]  ( .D(N1598), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1586]) );
  DFF \round_reg_reg[1587]  ( .D(N1599), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1587]) );
  DFF \round_reg_reg[1588]  ( .D(N1600), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1588]) );
  DFF \round_reg_reg[1589]  ( .D(N1601), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1589]) );
  DFF \round_reg_reg[1590]  ( .D(N1602), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1590]) );
  DFF \round_reg_reg[1591]  ( .D(N1603), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1591]) );
  DFF \round_reg_reg[1592]  ( .D(N1604), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1592]) );
  DFF \round_reg_reg[1593]  ( .D(N1605), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1593]) );
  DFF \round_reg_reg[1594]  ( .D(N1606), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1594]) );
  DFF \round_reg_reg[1595]  ( .D(N1607), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1595]) );
  DFF \round_reg_reg[1596]  ( .D(N1608), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1596]) );
  DFF \round_reg_reg[1597]  ( .D(N1609), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1597]) );
  DFF \round_reg_reg[1598]  ( .D(N1610), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1598]) );
  DFF \round_reg_reg[1599]  ( .D(N1611), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1599]) );
  IV U5993 ( .A(rst), .Z(n2763) );
  ANDN U5995 ( .B(rc_i[3]), .A(rst), .Z(N10) );
  ANDN U5996 ( .B(out[88]), .A(rst), .Z(N100) );
  ANDN U5997 ( .B(out[988]), .A(rst), .Z(N1000) );
  ANDN U5998 ( .B(out[989]), .A(rst), .Z(N1001) );
  ANDN U5999 ( .B(out[990]), .A(rst), .Z(N1002) );
  ANDN U6000 ( .B(out[991]), .A(rst), .Z(N1003) );
  ANDN U6001 ( .B(out[992]), .A(rst), .Z(N1004) );
  ANDN U6002 ( .B(out[993]), .A(rst), .Z(N1005) );
  ANDN U6003 ( .B(out[994]), .A(rst), .Z(N1006) );
  ANDN U6004 ( .B(out[995]), .A(rst), .Z(N1007) );
  ANDN U6005 ( .B(out[996]), .A(rst), .Z(N1008) );
  ANDN U6006 ( .B(out[997]), .A(rst), .Z(N1009) );
  ANDN U6007 ( .B(out[89]), .A(rst), .Z(N101) );
  ANDN U6008 ( .B(out[998]), .A(rst), .Z(N1010) );
  ANDN U6009 ( .B(out[999]), .A(rst), .Z(N1011) );
  ANDN U6010 ( .B(out[1000]), .A(rst), .Z(N1012) );
  ANDN U6011 ( .B(out[1001]), .A(rst), .Z(N1013) );
  ANDN U6012 ( .B(out[1002]), .A(rst), .Z(N1014) );
  ANDN U6013 ( .B(out[1003]), .A(rst), .Z(N1015) );
  ANDN U6014 ( .B(out[1004]), .A(rst), .Z(N1016) );
  ANDN U6015 ( .B(out[1005]), .A(rst), .Z(N1017) );
  ANDN U6016 ( .B(out[1006]), .A(rst), .Z(N1018) );
  ANDN U6017 ( .B(out[1007]), .A(rst), .Z(N1019) );
  ANDN U6018 ( .B(out[90]), .A(rst), .Z(N102) );
  ANDN U6019 ( .B(out[1008]), .A(rst), .Z(N1020) );
  ANDN U6020 ( .B(out[1009]), .A(rst), .Z(N1021) );
  ANDN U6021 ( .B(out[1010]), .A(rst), .Z(N1022) );
  ANDN U6022 ( .B(out[1011]), .A(rst), .Z(N1023) );
  ANDN U6023 ( .B(out[1012]), .A(rst), .Z(N1024) );
  ANDN U6024 ( .B(out[1013]), .A(rst), .Z(N1025) );
  ANDN U6025 ( .B(out[1014]), .A(rst), .Z(N1026) );
  ANDN U6026 ( .B(out[1015]), .A(rst), .Z(N1027) );
  ANDN U6027 ( .B(out[1016]), .A(rst), .Z(N1028) );
  ANDN U6028 ( .B(out[1017]), .A(rst), .Z(N1029) );
  ANDN U6029 ( .B(out[91]), .A(rst), .Z(N103) );
  ANDN U6030 ( .B(out[1018]), .A(rst), .Z(N1030) );
  ANDN U6031 ( .B(out[1019]), .A(rst), .Z(N1031) );
  ANDN U6032 ( .B(out[1020]), .A(rst), .Z(N1032) );
  ANDN U6033 ( .B(out[1021]), .A(rst), .Z(N1033) );
  ANDN U6034 ( .B(out[1022]), .A(rst), .Z(N1034) );
  ANDN U6035 ( .B(out[1023]), .A(rst), .Z(N1035) );
  ANDN U6036 ( .B(out[1024]), .A(rst), .Z(N1036) );
  ANDN U6037 ( .B(out[1025]), .A(rst), .Z(N1037) );
  ANDN U6038 ( .B(out[1026]), .A(rst), .Z(N1038) );
  ANDN U6039 ( .B(out[1027]), .A(rst), .Z(N1039) );
  ANDN U6040 ( .B(out[92]), .A(rst), .Z(N104) );
  ANDN U6041 ( .B(out[1028]), .A(rst), .Z(N1040) );
  ANDN U6042 ( .B(out[1029]), .A(rst), .Z(N1041) );
  ANDN U6043 ( .B(out[1030]), .A(rst), .Z(N1042) );
  ANDN U6044 ( .B(out[1031]), .A(rst), .Z(N1043) );
  ANDN U6045 ( .B(out[1032]), .A(rst), .Z(N1044) );
  ANDN U6046 ( .B(out[1033]), .A(rst), .Z(N1045) );
  ANDN U6047 ( .B(out[1034]), .A(rst), .Z(N1046) );
  ANDN U6048 ( .B(out[1035]), .A(rst), .Z(N1047) );
  ANDN U6049 ( .B(out[1036]), .A(rst), .Z(N1048) );
  ANDN U6050 ( .B(out[1037]), .A(rst), .Z(N1049) );
  ANDN U6051 ( .B(out[93]), .A(rst), .Z(N105) );
  ANDN U6052 ( .B(out[1038]), .A(rst), .Z(N1050) );
  ANDN U6053 ( .B(out[1039]), .A(rst), .Z(N1051) );
  ANDN U6054 ( .B(out[1040]), .A(rst), .Z(N1052) );
  ANDN U6055 ( .B(out[1041]), .A(rst), .Z(N1053) );
  ANDN U6056 ( .B(out[1042]), .A(rst), .Z(N1054) );
  ANDN U6057 ( .B(out[1043]), .A(rst), .Z(N1055) );
  ANDN U6058 ( .B(out[1044]), .A(rst), .Z(N1056) );
  ANDN U6059 ( .B(out[1045]), .A(rst), .Z(N1057) );
  ANDN U6060 ( .B(out[1046]), .A(rst), .Z(N1058) );
  ANDN U6061 ( .B(out[1047]), .A(rst), .Z(N1059) );
  ANDN U6062 ( .B(out[94]), .A(rst), .Z(N106) );
  ANDN U6063 ( .B(out[1048]), .A(rst), .Z(N1060) );
  ANDN U6064 ( .B(out[1049]), .A(rst), .Z(N1061) );
  ANDN U6065 ( .B(out[1050]), .A(rst), .Z(N1062) );
  ANDN U6066 ( .B(out[1051]), .A(rst), .Z(N1063) );
  ANDN U6067 ( .B(out[1052]), .A(rst), .Z(N1064) );
  ANDN U6068 ( .B(out[1053]), .A(rst), .Z(N1065) );
  ANDN U6069 ( .B(out[1054]), .A(rst), .Z(N1066) );
  ANDN U6070 ( .B(out[1055]), .A(rst), .Z(N1067) );
  ANDN U6071 ( .B(out[1056]), .A(rst), .Z(N1068) );
  ANDN U6072 ( .B(out[1057]), .A(rst), .Z(N1069) );
  ANDN U6073 ( .B(out[95]), .A(rst), .Z(N107) );
  ANDN U6074 ( .B(out[1058]), .A(rst), .Z(N1070) );
  ANDN U6075 ( .B(out[1059]), .A(rst), .Z(N1071) );
  ANDN U6076 ( .B(out[1060]), .A(rst), .Z(N1072) );
  ANDN U6077 ( .B(out[1061]), .A(rst), .Z(N1073) );
  ANDN U6078 ( .B(out[1062]), .A(rst), .Z(N1074) );
  ANDN U6079 ( .B(out[1063]), .A(rst), .Z(N1075) );
  ANDN U6080 ( .B(out[1064]), .A(rst), .Z(N1076) );
  ANDN U6081 ( .B(out[1065]), .A(rst), .Z(N1077) );
  ANDN U6082 ( .B(out[1066]), .A(rst), .Z(N1078) );
  ANDN U6083 ( .B(out[1067]), .A(rst), .Z(N1079) );
  ANDN U6084 ( .B(out[96]), .A(rst), .Z(N108) );
  ANDN U6085 ( .B(out[1068]), .A(rst), .Z(N1080) );
  ANDN U6086 ( .B(out[1069]), .A(rst), .Z(N1081) );
  ANDN U6087 ( .B(out[1070]), .A(rst), .Z(N1082) );
  ANDN U6088 ( .B(out[1071]), .A(rst), .Z(N1083) );
  ANDN U6089 ( .B(out[1072]), .A(rst), .Z(N1084) );
  ANDN U6090 ( .B(out[1073]), .A(rst), .Z(N1085) );
  ANDN U6091 ( .B(out[1074]), .A(rst), .Z(N1086) );
  ANDN U6092 ( .B(out[1075]), .A(rst), .Z(N1087) );
  ANDN U6093 ( .B(out[1076]), .A(rst), .Z(N1088) );
  ANDN U6094 ( .B(out[1077]), .A(rst), .Z(N1089) );
  ANDN U6095 ( .B(out[97]), .A(rst), .Z(N109) );
  ANDN U6096 ( .B(out[1078]), .A(rst), .Z(N1090) );
  ANDN U6097 ( .B(out[1079]), .A(rst), .Z(N1091) );
  ANDN U6098 ( .B(out[1080]), .A(rst), .Z(N1092) );
  ANDN U6099 ( .B(out[1081]), .A(rst), .Z(N1093) );
  ANDN U6100 ( .B(out[1082]), .A(rst), .Z(N1094) );
  ANDN U6101 ( .B(out[1083]), .A(rst), .Z(N1095) );
  ANDN U6102 ( .B(out[1084]), .A(rst), .Z(N1096) );
  ANDN U6103 ( .B(out[1085]), .A(rst), .Z(N1097) );
  ANDN U6104 ( .B(out[1086]), .A(rst), .Z(N1098) );
  ANDN U6105 ( .B(out[1087]), .A(rst), .Z(N1099) );
  ANDN U6106 ( .B(rc_i[4]), .A(rst), .Z(N11) );
  ANDN U6107 ( .B(out[98]), .A(rst), .Z(N110) );
  ANDN U6108 ( .B(out[1088]), .A(rst), .Z(N1100) );
  ANDN U6109 ( .B(out[1089]), .A(rst), .Z(N1101) );
  ANDN U6110 ( .B(out[1090]), .A(rst), .Z(N1102) );
  ANDN U6111 ( .B(out[1091]), .A(rst), .Z(N1103) );
  ANDN U6112 ( .B(out[1092]), .A(rst), .Z(N1104) );
  ANDN U6113 ( .B(out[1093]), .A(rst), .Z(N1105) );
  ANDN U6114 ( .B(out[1094]), .A(rst), .Z(N1106) );
  ANDN U6115 ( .B(out[1095]), .A(rst), .Z(N1107) );
  ANDN U6116 ( .B(out[1096]), .A(rst), .Z(N1108) );
  ANDN U6117 ( .B(out[1097]), .A(rst), .Z(N1109) );
  ANDN U6118 ( .B(out[99]), .A(rst), .Z(N111) );
  ANDN U6119 ( .B(out[1098]), .A(rst), .Z(N1110) );
  ANDN U6120 ( .B(out[1099]), .A(rst), .Z(N1111) );
  ANDN U6121 ( .B(out[1100]), .A(rst), .Z(N1112) );
  ANDN U6122 ( .B(out[1101]), .A(rst), .Z(N1113) );
  ANDN U6123 ( .B(out[1102]), .A(rst), .Z(N1114) );
  ANDN U6124 ( .B(out[1103]), .A(rst), .Z(N1115) );
  ANDN U6125 ( .B(out[1104]), .A(rst), .Z(N1116) );
  ANDN U6126 ( .B(out[1105]), .A(rst), .Z(N1117) );
  ANDN U6127 ( .B(out[1106]), .A(rst), .Z(N1118) );
  ANDN U6128 ( .B(out[1107]), .A(rst), .Z(N1119) );
  ANDN U6129 ( .B(out[100]), .A(rst), .Z(N112) );
  ANDN U6130 ( .B(out[1108]), .A(rst), .Z(N1120) );
  ANDN U6131 ( .B(out[1109]), .A(rst), .Z(N1121) );
  ANDN U6132 ( .B(out[1110]), .A(rst), .Z(N1122) );
  ANDN U6133 ( .B(out[1111]), .A(rst), .Z(N1123) );
  ANDN U6134 ( .B(out[1112]), .A(rst), .Z(N1124) );
  ANDN U6135 ( .B(out[1113]), .A(rst), .Z(N1125) );
  ANDN U6136 ( .B(out[1114]), .A(rst), .Z(N1126) );
  ANDN U6137 ( .B(out[1115]), .A(rst), .Z(N1127) );
  ANDN U6138 ( .B(out[1116]), .A(rst), .Z(N1128) );
  ANDN U6139 ( .B(out[1117]), .A(rst), .Z(N1129) );
  ANDN U6140 ( .B(out[101]), .A(rst), .Z(N113) );
  ANDN U6141 ( .B(out[1118]), .A(rst), .Z(N1130) );
  ANDN U6142 ( .B(out[1119]), .A(rst), .Z(N1131) );
  ANDN U6143 ( .B(out[1120]), .A(rst), .Z(N1132) );
  ANDN U6144 ( .B(out[1121]), .A(rst), .Z(N1133) );
  ANDN U6145 ( .B(out[1122]), .A(rst), .Z(N1134) );
  ANDN U6146 ( .B(out[1123]), .A(rst), .Z(N1135) );
  ANDN U6147 ( .B(out[1124]), .A(rst), .Z(N1136) );
  ANDN U6148 ( .B(out[1125]), .A(rst), .Z(N1137) );
  ANDN U6149 ( .B(out[1126]), .A(rst), .Z(N1138) );
  ANDN U6150 ( .B(out[1127]), .A(rst), .Z(N1139) );
  ANDN U6151 ( .B(out[102]), .A(rst), .Z(N114) );
  ANDN U6152 ( .B(out[1128]), .A(rst), .Z(N1140) );
  ANDN U6153 ( .B(out[1129]), .A(rst), .Z(N1141) );
  ANDN U6154 ( .B(out[1130]), .A(rst), .Z(N1142) );
  ANDN U6155 ( .B(out[1131]), .A(rst), .Z(N1143) );
  ANDN U6156 ( .B(out[1132]), .A(rst), .Z(N1144) );
  ANDN U6157 ( .B(out[1133]), .A(rst), .Z(N1145) );
  ANDN U6158 ( .B(out[1134]), .A(rst), .Z(N1146) );
  ANDN U6159 ( .B(out[1135]), .A(rst), .Z(N1147) );
  ANDN U6160 ( .B(out[1136]), .A(rst), .Z(N1148) );
  ANDN U6161 ( .B(out[1137]), .A(rst), .Z(N1149) );
  ANDN U6162 ( .B(out[103]), .A(rst), .Z(N115) );
  ANDN U6163 ( .B(out[1138]), .A(rst), .Z(N1150) );
  ANDN U6164 ( .B(out[1139]), .A(rst), .Z(N1151) );
  ANDN U6165 ( .B(out[1140]), .A(rst), .Z(N1152) );
  ANDN U6166 ( .B(out[1141]), .A(rst), .Z(N1153) );
  ANDN U6167 ( .B(out[1142]), .A(rst), .Z(N1154) );
  ANDN U6168 ( .B(out[1143]), .A(rst), .Z(N1155) );
  ANDN U6169 ( .B(out[1144]), .A(rst), .Z(N1156) );
  ANDN U6170 ( .B(out[1145]), .A(rst), .Z(N1157) );
  ANDN U6171 ( .B(out[1146]), .A(rst), .Z(N1158) );
  ANDN U6172 ( .B(out[1147]), .A(rst), .Z(N1159) );
  ANDN U6173 ( .B(out[104]), .A(rst), .Z(N116) );
  ANDN U6174 ( .B(out[1148]), .A(rst), .Z(N1160) );
  ANDN U6175 ( .B(out[1149]), .A(rst), .Z(N1161) );
  ANDN U6176 ( .B(out[1150]), .A(rst), .Z(N1162) );
  ANDN U6177 ( .B(out[1151]), .A(rst), .Z(N1163) );
  ANDN U6178 ( .B(out[1152]), .A(rst), .Z(N1164) );
  ANDN U6179 ( .B(out[1153]), .A(rst), .Z(N1165) );
  ANDN U6180 ( .B(out[1154]), .A(rst), .Z(N1166) );
  ANDN U6181 ( .B(out[1155]), .A(rst), .Z(N1167) );
  ANDN U6182 ( .B(out[1156]), .A(rst), .Z(N1168) );
  ANDN U6183 ( .B(out[1157]), .A(rst), .Z(N1169) );
  ANDN U6184 ( .B(out[105]), .A(rst), .Z(N117) );
  ANDN U6185 ( .B(out[1158]), .A(rst), .Z(N1170) );
  ANDN U6186 ( .B(out[1159]), .A(rst), .Z(N1171) );
  ANDN U6187 ( .B(out[1160]), .A(rst), .Z(N1172) );
  ANDN U6188 ( .B(out[1161]), .A(rst), .Z(N1173) );
  ANDN U6189 ( .B(out[1162]), .A(rst), .Z(N1174) );
  ANDN U6190 ( .B(out[1163]), .A(rst), .Z(N1175) );
  ANDN U6191 ( .B(out[1164]), .A(rst), .Z(N1176) );
  ANDN U6192 ( .B(out[1165]), .A(rst), .Z(N1177) );
  ANDN U6193 ( .B(out[1166]), .A(rst), .Z(N1178) );
  ANDN U6194 ( .B(out[1167]), .A(rst), .Z(N1179) );
  ANDN U6195 ( .B(out[106]), .A(rst), .Z(N118) );
  ANDN U6196 ( .B(out[1168]), .A(rst), .Z(N1180) );
  ANDN U6197 ( .B(out[1169]), .A(rst), .Z(N1181) );
  ANDN U6198 ( .B(out[1170]), .A(rst), .Z(N1182) );
  ANDN U6199 ( .B(out[1171]), .A(rst), .Z(N1183) );
  ANDN U6200 ( .B(out[1172]), .A(rst), .Z(N1184) );
  ANDN U6201 ( .B(out[1173]), .A(rst), .Z(N1185) );
  ANDN U6202 ( .B(out[1174]), .A(rst), .Z(N1186) );
  ANDN U6203 ( .B(out[1175]), .A(rst), .Z(N1187) );
  ANDN U6204 ( .B(out[1176]), .A(rst), .Z(N1188) );
  ANDN U6205 ( .B(out[1177]), .A(rst), .Z(N1189) );
  ANDN U6206 ( .B(out[107]), .A(rst), .Z(N119) );
  ANDN U6207 ( .B(out[1178]), .A(rst), .Z(N1190) );
  ANDN U6208 ( .B(out[1179]), .A(rst), .Z(N1191) );
  ANDN U6209 ( .B(out[1180]), .A(rst), .Z(N1192) );
  ANDN U6210 ( .B(out[1181]), .A(rst), .Z(N1193) );
  ANDN U6211 ( .B(out[1182]), .A(rst), .Z(N1194) );
  ANDN U6212 ( .B(out[1183]), .A(rst), .Z(N1195) );
  ANDN U6213 ( .B(out[1184]), .A(rst), .Z(N1196) );
  ANDN U6214 ( .B(out[1185]), .A(rst), .Z(N1197) );
  ANDN U6215 ( .B(out[1186]), .A(rst), .Z(N1198) );
  ANDN U6216 ( .B(out[1187]), .A(rst), .Z(N1199) );
  ANDN U6217 ( .B(out[0]), .A(rst), .Z(N12) );
  ANDN U6218 ( .B(out[108]), .A(rst), .Z(N120) );
  ANDN U6219 ( .B(out[1188]), .A(rst), .Z(N1200) );
  ANDN U6220 ( .B(out[1189]), .A(rst), .Z(N1201) );
  ANDN U6221 ( .B(out[1190]), .A(rst), .Z(N1202) );
  ANDN U6222 ( .B(out[1191]), .A(rst), .Z(N1203) );
  ANDN U6223 ( .B(out[1192]), .A(rst), .Z(N1204) );
  ANDN U6224 ( .B(out[1193]), .A(rst), .Z(N1205) );
  ANDN U6225 ( .B(out[1194]), .A(rst), .Z(N1206) );
  ANDN U6226 ( .B(out[1195]), .A(rst), .Z(N1207) );
  ANDN U6227 ( .B(out[1196]), .A(rst), .Z(N1208) );
  ANDN U6228 ( .B(out[1197]), .A(rst), .Z(N1209) );
  ANDN U6229 ( .B(out[109]), .A(rst), .Z(N121) );
  ANDN U6230 ( .B(out[1198]), .A(rst), .Z(N1210) );
  ANDN U6231 ( .B(out[1199]), .A(rst), .Z(N1211) );
  ANDN U6232 ( .B(out[1200]), .A(rst), .Z(N1212) );
  ANDN U6233 ( .B(out[1201]), .A(rst), .Z(N1213) );
  ANDN U6234 ( .B(out[1202]), .A(rst), .Z(N1214) );
  ANDN U6235 ( .B(out[1203]), .A(rst), .Z(N1215) );
  ANDN U6236 ( .B(out[1204]), .A(rst), .Z(N1216) );
  ANDN U6237 ( .B(out[1205]), .A(rst), .Z(N1217) );
  ANDN U6238 ( .B(out[1206]), .A(rst), .Z(N1218) );
  ANDN U6239 ( .B(out[1207]), .A(rst), .Z(N1219) );
  ANDN U6240 ( .B(out[110]), .A(rst), .Z(N122) );
  ANDN U6241 ( .B(out[1208]), .A(rst), .Z(N1220) );
  ANDN U6242 ( .B(out[1209]), .A(rst), .Z(N1221) );
  ANDN U6243 ( .B(out[1210]), .A(rst), .Z(N1222) );
  ANDN U6244 ( .B(out[1211]), .A(rst), .Z(N1223) );
  ANDN U6245 ( .B(out[1212]), .A(rst), .Z(N1224) );
  ANDN U6246 ( .B(out[1213]), .A(rst), .Z(N1225) );
  ANDN U6247 ( .B(out[1214]), .A(rst), .Z(N1226) );
  ANDN U6248 ( .B(out[1215]), .A(rst), .Z(N1227) );
  ANDN U6249 ( .B(out[1216]), .A(rst), .Z(N1228) );
  ANDN U6250 ( .B(out[1217]), .A(rst), .Z(N1229) );
  ANDN U6251 ( .B(out[111]), .A(rst), .Z(N123) );
  ANDN U6252 ( .B(out[1218]), .A(rst), .Z(N1230) );
  ANDN U6253 ( .B(out[1219]), .A(rst), .Z(N1231) );
  ANDN U6254 ( .B(out[1220]), .A(rst), .Z(N1232) );
  ANDN U6255 ( .B(out[1221]), .A(rst), .Z(N1233) );
  ANDN U6256 ( .B(out[1222]), .A(rst), .Z(N1234) );
  ANDN U6257 ( .B(out[1223]), .A(rst), .Z(N1235) );
  ANDN U6258 ( .B(out[1224]), .A(rst), .Z(N1236) );
  ANDN U6259 ( .B(out[1225]), .A(rst), .Z(N1237) );
  ANDN U6260 ( .B(out[1226]), .A(rst), .Z(N1238) );
  ANDN U6261 ( .B(out[1227]), .A(rst), .Z(N1239) );
  ANDN U6262 ( .B(out[112]), .A(rst), .Z(N124) );
  ANDN U6263 ( .B(out[1228]), .A(rst), .Z(N1240) );
  ANDN U6264 ( .B(out[1229]), .A(rst), .Z(N1241) );
  ANDN U6265 ( .B(out[1230]), .A(rst), .Z(N1242) );
  ANDN U6266 ( .B(out[1231]), .A(rst), .Z(N1243) );
  ANDN U6267 ( .B(out[1232]), .A(rst), .Z(N1244) );
  ANDN U6268 ( .B(out[1233]), .A(rst), .Z(N1245) );
  ANDN U6269 ( .B(out[1234]), .A(rst), .Z(N1246) );
  ANDN U6270 ( .B(out[1235]), .A(rst), .Z(N1247) );
  ANDN U6271 ( .B(out[1236]), .A(rst), .Z(N1248) );
  ANDN U6272 ( .B(out[1237]), .A(rst), .Z(N1249) );
  ANDN U6273 ( .B(out[113]), .A(rst), .Z(N125) );
  ANDN U6274 ( .B(out[1238]), .A(rst), .Z(N1250) );
  ANDN U6275 ( .B(out[1239]), .A(rst), .Z(N1251) );
  ANDN U6276 ( .B(out[1240]), .A(rst), .Z(N1252) );
  ANDN U6277 ( .B(out[1241]), .A(rst), .Z(N1253) );
  ANDN U6278 ( .B(out[1242]), .A(rst), .Z(N1254) );
  ANDN U6279 ( .B(out[1243]), .A(rst), .Z(N1255) );
  ANDN U6280 ( .B(out[1244]), .A(rst), .Z(N1256) );
  ANDN U6281 ( .B(out[1245]), .A(rst), .Z(N1257) );
  ANDN U6282 ( .B(out[1246]), .A(rst), .Z(N1258) );
  ANDN U6283 ( .B(out[1247]), .A(rst), .Z(N1259) );
  ANDN U6284 ( .B(out[114]), .A(rst), .Z(N126) );
  ANDN U6285 ( .B(out[1248]), .A(rst), .Z(N1260) );
  ANDN U6286 ( .B(out[1249]), .A(rst), .Z(N1261) );
  ANDN U6287 ( .B(out[1250]), .A(rst), .Z(N1262) );
  ANDN U6288 ( .B(out[1251]), .A(rst), .Z(N1263) );
  ANDN U6289 ( .B(out[1252]), .A(rst), .Z(N1264) );
  ANDN U6290 ( .B(out[1253]), .A(rst), .Z(N1265) );
  ANDN U6291 ( .B(out[1254]), .A(rst), .Z(N1266) );
  ANDN U6292 ( .B(out[1255]), .A(rst), .Z(N1267) );
  ANDN U6293 ( .B(out[1256]), .A(rst), .Z(N1268) );
  ANDN U6294 ( .B(out[1257]), .A(rst), .Z(N1269) );
  ANDN U6295 ( .B(out[115]), .A(rst), .Z(N127) );
  ANDN U6296 ( .B(out[1258]), .A(rst), .Z(N1270) );
  ANDN U6297 ( .B(out[1259]), .A(rst), .Z(N1271) );
  ANDN U6298 ( .B(out[1260]), .A(rst), .Z(N1272) );
  ANDN U6299 ( .B(out[1261]), .A(rst), .Z(N1273) );
  ANDN U6300 ( .B(out[1262]), .A(rst), .Z(N1274) );
  ANDN U6301 ( .B(out[1263]), .A(rst), .Z(N1275) );
  ANDN U6302 ( .B(out[1264]), .A(rst), .Z(N1276) );
  ANDN U6303 ( .B(out[1265]), .A(rst), .Z(N1277) );
  ANDN U6304 ( .B(out[1266]), .A(rst), .Z(N1278) );
  ANDN U6305 ( .B(out[1267]), .A(rst), .Z(N1279) );
  ANDN U6306 ( .B(out[116]), .A(rst), .Z(N128) );
  ANDN U6307 ( .B(out[1268]), .A(rst), .Z(N1280) );
  ANDN U6308 ( .B(out[1269]), .A(rst), .Z(N1281) );
  ANDN U6309 ( .B(out[1270]), .A(rst), .Z(N1282) );
  ANDN U6310 ( .B(out[1271]), .A(rst), .Z(N1283) );
  ANDN U6311 ( .B(out[1272]), .A(rst), .Z(N1284) );
  ANDN U6312 ( .B(out[1273]), .A(rst), .Z(N1285) );
  ANDN U6313 ( .B(out[1274]), .A(rst), .Z(N1286) );
  ANDN U6314 ( .B(out[1275]), .A(rst), .Z(N1287) );
  ANDN U6315 ( .B(out[1276]), .A(rst), .Z(N1288) );
  ANDN U6316 ( .B(out[1277]), .A(rst), .Z(N1289) );
  ANDN U6317 ( .B(out[117]), .A(rst), .Z(N129) );
  ANDN U6318 ( .B(out[1278]), .A(rst), .Z(N1290) );
  ANDN U6319 ( .B(out[1279]), .A(rst), .Z(N1291) );
  ANDN U6320 ( .B(out[1280]), .A(rst), .Z(N1292) );
  ANDN U6321 ( .B(out[1281]), .A(rst), .Z(N1293) );
  ANDN U6322 ( .B(out[1282]), .A(rst), .Z(N1294) );
  ANDN U6323 ( .B(out[1283]), .A(rst), .Z(N1295) );
  ANDN U6324 ( .B(out[1284]), .A(rst), .Z(N1296) );
  ANDN U6325 ( .B(out[1285]), .A(rst), .Z(N1297) );
  ANDN U6326 ( .B(out[1286]), .A(rst), .Z(N1298) );
  ANDN U6327 ( .B(out[1287]), .A(rst), .Z(N1299) );
  ANDN U6328 ( .B(out[1]), .A(rst), .Z(N13) );
  ANDN U6329 ( .B(out[118]), .A(rst), .Z(N130) );
  ANDN U6330 ( .B(out[1288]), .A(rst), .Z(N1300) );
  ANDN U6331 ( .B(out[1289]), .A(rst), .Z(N1301) );
  ANDN U6332 ( .B(out[1290]), .A(rst), .Z(N1302) );
  ANDN U6333 ( .B(out[1291]), .A(rst), .Z(N1303) );
  ANDN U6334 ( .B(out[1292]), .A(rst), .Z(N1304) );
  ANDN U6335 ( .B(out[1293]), .A(rst), .Z(N1305) );
  ANDN U6336 ( .B(out[1294]), .A(rst), .Z(N1306) );
  ANDN U6337 ( .B(out[1295]), .A(rst), .Z(N1307) );
  ANDN U6338 ( .B(out[1296]), .A(rst), .Z(N1308) );
  ANDN U6339 ( .B(out[1297]), .A(rst), .Z(N1309) );
  ANDN U6340 ( .B(out[119]), .A(rst), .Z(N131) );
  ANDN U6341 ( .B(out[1298]), .A(rst), .Z(N1310) );
  ANDN U6342 ( .B(out[1299]), .A(rst), .Z(N1311) );
  ANDN U6343 ( .B(out[1300]), .A(rst), .Z(N1312) );
  ANDN U6344 ( .B(out[1301]), .A(rst), .Z(N1313) );
  ANDN U6345 ( .B(out[1302]), .A(rst), .Z(N1314) );
  ANDN U6346 ( .B(out[1303]), .A(rst), .Z(N1315) );
  ANDN U6347 ( .B(out[1304]), .A(rst), .Z(N1316) );
  ANDN U6348 ( .B(out[1305]), .A(rst), .Z(N1317) );
  ANDN U6349 ( .B(out[1306]), .A(rst), .Z(N1318) );
  ANDN U6350 ( .B(out[1307]), .A(rst), .Z(N1319) );
  ANDN U6351 ( .B(out[120]), .A(rst), .Z(N132) );
  ANDN U6352 ( .B(out[1308]), .A(rst), .Z(N1320) );
  ANDN U6353 ( .B(out[1309]), .A(rst), .Z(N1321) );
  ANDN U6354 ( .B(out[1310]), .A(rst), .Z(N1322) );
  ANDN U6355 ( .B(out[1311]), .A(rst), .Z(N1323) );
  ANDN U6356 ( .B(out[1312]), .A(rst), .Z(N1324) );
  ANDN U6357 ( .B(out[1313]), .A(rst), .Z(N1325) );
  ANDN U6358 ( .B(out[1314]), .A(rst), .Z(N1326) );
  ANDN U6359 ( .B(out[1315]), .A(rst), .Z(N1327) );
  ANDN U6360 ( .B(out[1316]), .A(rst), .Z(N1328) );
  ANDN U6361 ( .B(out[1317]), .A(rst), .Z(N1329) );
  ANDN U6362 ( .B(out[121]), .A(rst), .Z(N133) );
  ANDN U6363 ( .B(out[1318]), .A(rst), .Z(N1330) );
  ANDN U6364 ( .B(out[1319]), .A(rst), .Z(N1331) );
  ANDN U6365 ( .B(out[1320]), .A(rst), .Z(N1332) );
  ANDN U6366 ( .B(out[1321]), .A(rst), .Z(N1333) );
  ANDN U6367 ( .B(out[1322]), .A(rst), .Z(N1334) );
  ANDN U6368 ( .B(out[1323]), .A(rst), .Z(N1335) );
  ANDN U6369 ( .B(out[1324]), .A(rst), .Z(N1336) );
  ANDN U6370 ( .B(out[1325]), .A(rst), .Z(N1337) );
  ANDN U6371 ( .B(out[1326]), .A(rst), .Z(N1338) );
  ANDN U6372 ( .B(out[1327]), .A(rst), .Z(N1339) );
  ANDN U6373 ( .B(out[122]), .A(rst), .Z(N134) );
  ANDN U6374 ( .B(out[1328]), .A(rst), .Z(N1340) );
  ANDN U6375 ( .B(out[1329]), .A(rst), .Z(N1341) );
  ANDN U6376 ( .B(out[1330]), .A(rst), .Z(N1342) );
  ANDN U6377 ( .B(out[1331]), .A(rst), .Z(N1343) );
  ANDN U6378 ( .B(out[1332]), .A(rst), .Z(N1344) );
  ANDN U6379 ( .B(out[1333]), .A(rst), .Z(N1345) );
  ANDN U6380 ( .B(out[1334]), .A(rst), .Z(N1346) );
  ANDN U6381 ( .B(out[1335]), .A(rst), .Z(N1347) );
  ANDN U6382 ( .B(out[1336]), .A(rst), .Z(N1348) );
  ANDN U6383 ( .B(out[1337]), .A(rst), .Z(N1349) );
  ANDN U6384 ( .B(out[123]), .A(rst), .Z(N135) );
  ANDN U6385 ( .B(out[1338]), .A(rst), .Z(N1350) );
  ANDN U6386 ( .B(out[1339]), .A(rst), .Z(N1351) );
  ANDN U6387 ( .B(out[1340]), .A(rst), .Z(N1352) );
  ANDN U6388 ( .B(out[1341]), .A(rst), .Z(N1353) );
  ANDN U6389 ( .B(out[1342]), .A(rst), .Z(N1354) );
  ANDN U6390 ( .B(out[1343]), .A(rst), .Z(N1355) );
  ANDN U6391 ( .B(out[1344]), .A(rst), .Z(N1356) );
  ANDN U6392 ( .B(out[1345]), .A(rst), .Z(N1357) );
  ANDN U6393 ( .B(out[1346]), .A(rst), .Z(N1358) );
  ANDN U6394 ( .B(out[1347]), .A(rst), .Z(N1359) );
  ANDN U6395 ( .B(out[124]), .A(rst), .Z(N136) );
  ANDN U6396 ( .B(out[1348]), .A(rst), .Z(N1360) );
  ANDN U6397 ( .B(out[1349]), .A(rst), .Z(N1361) );
  ANDN U6398 ( .B(out[1350]), .A(rst), .Z(N1362) );
  ANDN U6399 ( .B(out[1351]), .A(rst), .Z(N1363) );
  ANDN U6400 ( .B(out[1352]), .A(rst), .Z(N1364) );
  ANDN U6401 ( .B(out[1353]), .A(rst), .Z(N1365) );
  ANDN U6402 ( .B(out[1354]), .A(rst), .Z(N1366) );
  ANDN U6403 ( .B(out[1355]), .A(rst), .Z(N1367) );
  ANDN U6404 ( .B(out[1356]), .A(rst), .Z(N1368) );
  ANDN U6405 ( .B(out[1357]), .A(rst), .Z(N1369) );
  ANDN U6406 ( .B(out[125]), .A(rst), .Z(N137) );
  ANDN U6407 ( .B(out[1358]), .A(rst), .Z(N1370) );
  ANDN U6408 ( .B(out[1359]), .A(rst), .Z(N1371) );
  ANDN U6409 ( .B(out[1360]), .A(rst), .Z(N1372) );
  ANDN U6410 ( .B(out[1361]), .A(rst), .Z(N1373) );
  ANDN U6411 ( .B(out[1362]), .A(rst), .Z(N1374) );
  ANDN U6412 ( .B(out[1363]), .A(rst), .Z(N1375) );
  ANDN U6413 ( .B(out[1364]), .A(rst), .Z(N1376) );
  ANDN U6414 ( .B(out[1365]), .A(rst), .Z(N1377) );
  ANDN U6415 ( .B(out[1366]), .A(rst), .Z(N1378) );
  ANDN U6416 ( .B(out[1367]), .A(rst), .Z(N1379) );
  ANDN U6417 ( .B(out[126]), .A(rst), .Z(N138) );
  ANDN U6418 ( .B(out[1368]), .A(rst), .Z(N1380) );
  ANDN U6419 ( .B(out[1369]), .A(rst), .Z(N1381) );
  ANDN U6420 ( .B(out[1370]), .A(rst), .Z(N1382) );
  ANDN U6421 ( .B(out[1371]), .A(rst), .Z(N1383) );
  ANDN U6422 ( .B(out[1372]), .A(rst), .Z(N1384) );
  ANDN U6423 ( .B(out[1373]), .A(rst), .Z(N1385) );
  ANDN U6424 ( .B(out[1374]), .A(rst), .Z(N1386) );
  ANDN U6425 ( .B(out[1375]), .A(rst), .Z(N1387) );
  ANDN U6426 ( .B(out[1376]), .A(rst), .Z(N1388) );
  ANDN U6427 ( .B(out[1377]), .A(rst), .Z(N1389) );
  ANDN U6428 ( .B(out[127]), .A(rst), .Z(N139) );
  ANDN U6429 ( .B(out[1378]), .A(rst), .Z(N1390) );
  ANDN U6430 ( .B(out[1379]), .A(rst), .Z(N1391) );
  ANDN U6431 ( .B(out[1380]), .A(rst), .Z(N1392) );
  ANDN U6432 ( .B(out[1381]), .A(rst), .Z(N1393) );
  ANDN U6433 ( .B(out[1382]), .A(rst), .Z(N1394) );
  ANDN U6434 ( .B(out[1383]), .A(rst), .Z(N1395) );
  ANDN U6435 ( .B(out[1384]), .A(rst), .Z(N1396) );
  ANDN U6436 ( .B(out[1385]), .A(rst), .Z(N1397) );
  ANDN U6437 ( .B(out[1386]), .A(rst), .Z(N1398) );
  ANDN U6438 ( .B(out[1387]), .A(rst), .Z(N1399) );
  ANDN U6439 ( .B(out[2]), .A(rst), .Z(N14) );
  ANDN U6440 ( .B(out[128]), .A(rst), .Z(N140) );
  ANDN U6441 ( .B(out[1388]), .A(rst), .Z(N1400) );
  ANDN U6442 ( .B(out[1389]), .A(rst), .Z(N1401) );
  ANDN U6443 ( .B(out[1390]), .A(rst), .Z(N1402) );
  ANDN U6444 ( .B(out[1391]), .A(rst), .Z(N1403) );
  ANDN U6445 ( .B(out[1392]), .A(rst), .Z(N1404) );
  ANDN U6446 ( .B(out[1393]), .A(rst), .Z(N1405) );
  ANDN U6447 ( .B(out[1394]), .A(rst), .Z(N1406) );
  ANDN U6448 ( .B(out[1395]), .A(rst), .Z(N1407) );
  ANDN U6449 ( .B(out[1396]), .A(rst), .Z(N1408) );
  ANDN U6450 ( .B(out[1397]), .A(rst), .Z(N1409) );
  ANDN U6451 ( .B(out[129]), .A(rst), .Z(N141) );
  ANDN U6452 ( .B(out[1398]), .A(rst), .Z(N1410) );
  ANDN U6453 ( .B(out[1399]), .A(rst), .Z(N1411) );
  ANDN U6454 ( .B(out[1400]), .A(rst), .Z(N1412) );
  ANDN U6455 ( .B(out[1401]), .A(rst), .Z(N1413) );
  ANDN U6456 ( .B(out[1402]), .A(rst), .Z(N1414) );
  ANDN U6457 ( .B(out[1403]), .A(rst), .Z(N1415) );
  ANDN U6458 ( .B(out[1404]), .A(rst), .Z(N1416) );
  ANDN U6459 ( .B(out[1405]), .A(rst), .Z(N1417) );
  ANDN U6460 ( .B(out[1406]), .A(rst), .Z(N1418) );
  ANDN U6461 ( .B(out[1407]), .A(rst), .Z(N1419) );
  ANDN U6462 ( .B(out[130]), .A(rst), .Z(N142) );
  ANDN U6463 ( .B(out[1408]), .A(rst), .Z(N1420) );
  ANDN U6464 ( .B(out[1409]), .A(rst), .Z(N1421) );
  ANDN U6465 ( .B(out[1410]), .A(rst), .Z(N1422) );
  ANDN U6466 ( .B(out[1411]), .A(rst), .Z(N1423) );
  ANDN U6467 ( .B(out[1412]), .A(rst), .Z(N1424) );
  ANDN U6468 ( .B(out[1413]), .A(rst), .Z(N1425) );
  ANDN U6469 ( .B(out[1414]), .A(rst), .Z(N1426) );
  ANDN U6470 ( .B(out[1415]), .A(rst), .Z(N1427) );
  ANDN U6471 ( .B(out[1416]), .A(rst), .Z(N1428) );
  ANDN U6472 ( .B(out[1417]), .A(rst), .Z(N1429) );
  ANDN U6473 ( .B(out[131]), .A(rst), .Z(N143) );
  ANDN U6474 ( .B(out[1418]), .A(rst), .Z(N1430) );
  ANDN U6475 ( .B(out[1419]), .A(rst), .Z(N1431) );
  ANDN U6476 ( .B(out[1420]), .A(rst), .Z(N1432) );
  ANDN U6477 ( .B(out[1421]), .A(rst), .Z(N1433) );
  ANDN U6478 ( .B(out[1422]), .A(rst), .Z(N1434) );
  ANDN U6479 ( .B(out[1423]), .A(rst), .Z(N1435) );
  ANDN U6480 ( .B(out[1424]), .A(rst), .Z(N1436) );
  ANDN U6481 ( .B(out[1425]), .A(rst), .Z(N1437) );
  ANDN U6482 ( .B(out[1426]), .A(rst), .Z(N1438) );
  ANDN U6483 ( .B(out[1427]), .A(rst), .Z(N1439) );
  ANDN U6484 ( .B(out[132]), .A(rst), .Z(N144) );
  ANDN U6485 ( .B(out[1428]), .A(rst), .Z(N1440) );
  ANDN U6486 ( .B(out[1429]), .A(rst), .Z(N1441) );
  ANDN U6487 ( .B(out[1430]), .A(rst), .Z(N1442) );
  ANDN U6488 ( .B(out[1431]), .A(rst), .Z(N1443) );
  ANDN U6489 ( .B(out[1432]), .A(rst), .Z(N1444) );
  ANDN U6490 ( .B(out[1433]), .A(rst), .Z(N1445) );
  ANDN U6491 ( .B(out[1434]), .A(rst), .Z(N1446) );
  ANDN U6492 ( .B(out[1435]), .A(rst), .Z(N1447) );
  ANDN U6493 ( .B(out[1436]), .A(rst), .Z(N1448) );
  ANDN U6494 ( .B(out[1437]), .A(rst), .Z(N1449) );
  ANDN U6495 ( .B(out[133]), .A(rst), .Z(N145) );
  ANDN U6496 ( .B(out[1438]), .A(rst), .Z(N1450) );
  ANDN U6497 ( .B(out[1439]), .A(rst), .Z(N1451) );
  ANDN U6498 ( .B(out[1440]), .A(rst), .Z(N1452) );
  ANDN U6499 ( .B(out[1441]), .A(rst), .Z(N1453) );
  ANDN U6500 ( .B(out[1442]), .A(rst), .Z(N1454) );
  ANDN U6501 ( .B(out[1443]), .A(rst), .Z(N1455) );
  ANDN U6502 ( .B(out[1444]), .A(rst), .Z(N1456) );
  ANDN U6503 ( .B(out[1445]), .A(rst), .Z(N1457) );
  ANDN U6504 ( .B(out[1446]), .A(rst), .Z(N1458) );
  ANDN U6505 ( .B(out[1447]), .A(rst), .Z(N1459) );
  ANDN U6506 ( .B(out[134]), .A(rst), .Z(N146) );
  ANDN U6507 ( .B(out[1448]), .A(rst), .Z(N1460) );
  ANDN U6508 ( .B(out[1449]), .A(rst), .Z(N1461) );
  ANDN U6509 ( .B(out[1450]), .A(rst), .Z(N1462) );
  ANDN U6510 ( .B(out[1451]), .A(rst), .Z(N1463) );
  ANDN U6511 ( .B(out[1452]), .A(rst), .Z(N1464) );
  ANDN U6512 ( .B(out[1453]), .A(rst), .Z(N1465) );
  ANDN U6513 ( .B(out[1454]), .A(rst), .Z(N1466) );
  ANDN U6514 ( .B(out[1455]), .A(rst), .Z(N1467) );
  ANDN U6515 ( .B(out[1456]), .A(rst), .Z(N1468) );
  ANDN U6516 ( .B(out[1457]), .A(rst), .Z(N1469) );
  ANDN U6517 ( .B(out[135]), .A(rst), .Z(N147) );
  ANDN U6518 ( .B(out[1458]), .A(rst), .Z(N1470) );
  ANDN U6519 ( .B(out[1459]), .A(rst), .Z(N1471) );
  ANDN U6520 ( .B(out[1460]), .A(rst), .Z(N1472) );
  ANDN U6521 ( .B(out[1461]), .A(rst), .Z(N1473) );
  ANDN U6522 ( .B(out[1462]), .A(rst), .Z(N1474) );
  ANDN U6523 ( .B(out[1463]), .A(rst), .Z(N1475) );
  ANDN U6524 ( .B(out[1464]), .A(rst), .Z(N1476) );
  ANDN U6525 ( .B(out[1465]), .A(rst), .Z(N1477) );
  ANDN U6526 ( .B(out[1466]), .A(rst), .Z(N1478) );
  ANDN U6527 ( .B(out[1467]), .A(rst), .Z(N1479) );
  ANDN U6528 ( .B(out[136]), .A(rst), .Z(N148) );
  ANDN U6529 ( .B(out[1468]), .A(rst), .Z(N1480) );
  ANDN U6530 ( .B(out[1469]), .A(rst), .Z(N1481) );
  ANDN U6531 ( .B(out[1470]), .A(rst), .Z(N1482) );
  ANDN U6532 ( .B(out[1471]), .A(rst), .Z(N1483) );
  ANDN U6533 ( .B(out[1472]), .A(rst), .Z(N1484) );
  ANDN U6534 ( .B(out[1473]), .A(rst), .Z(N1485) );
  ANDN U6535 ( .B(out[1474]), .A(rst), .Z(N1486) );
  ANDN U6536 ( .B(out[1475]), .A(rst), .Z(N1487) );
  ANDN U6537 ( .B(out[1476]), .A(rst), .Z(N1488) );
  ANDN U6538 ( .B(out[1477]), .A(rst), .Z(N1489) );
  ANDN U6539 ( .B(out[137]), .A(rst), .Z(N149) );
  ANDN U6540 ( .B(out[1478]), .A(rst), .Z(N1490) );
  ANDN U6541 ( .B(out[1479]), .A(rst), .Z(N1491) );
  ANDN U6542 ( .B(out[1480]), .A(rst), .Z(N1492) );
  ANDN U6543 ( .B(out[1481]), .A(rst), .Z(N1493) );
  ANDN U6544 ( .B(out[1482]), .A(rst), .Z(N1494) );
  ANDN U6545 ( .B(out[1483]), .A(rst), .Z(N1495) );
  ANDN U6546 ( .B(out[1484]), .A(rst), .Z(N1496) );
  ANDN U6547 ( .B(out[1485]), .A(rst), .Z(N1497) );
  ANDN U6548 ( .B(out[1486]), .A(rst), .Z(N1498) );
  ANDN U6549 ( .B(out[1487]), .A(rst), .Z(N1499) );
  ANDN U6550 ( .B(out[3]), .A(rst), .Z(N15) );
  ANDN U6551 ( .B(out[138]), .A(rst), .Z(N150) );
  ANDN U6552 ( .B(out[1488]), .A(rst), .Z(N1500) );
  ANDN U6553 ( .B(out[1489]), .A(rst), .Z(N1501) );
  ANDN U6554 ( .B(out[1490]), .A(rst), .Z(N1502) );
  ANDN U6555 ( .B(out[1491]), .A(rst), .Z(N1503) );
  ANDN U6556 ( .B(out[1492]), .A(rst), .Z(N1504) );
  ANDN U6557 ( .B(out[1493]), .A(rst), .Z(N1505) );
  ANDN U6558 ( .B(out[1494]), .A(rst), .Z(N1506) );
  ANDN U6559 ( .B(out[1495]), .A(rst), .Z(N1507) );
  ANDN U6560 ( .B(out[1496]), .A(rst), .Z(N1508) );
  ANDN U6561 ( .B(out[1497]), .A(rst), .Z(N1509) );
  ANDN U6562 ( .B(out[139]), .A(rst), .Z(N151) );
  ANDN U6563 ( .B(out[1498]), .A(rst), .Z(N1510) );
  ANDN U6564 ( .B(out[1499]), .A(rst), .Z(N1511) );
  ANDN U6565 ( .B(out[1500]), .A(rst), .Z(N1512) );
  ANDN U6566 ( .B(out[1501]), .A(rst), .Z(N1513) );
  ANDN U6567 ( .B(out[1502]), .A(rst), .Z(N1514) );
  ANDN U6568 ( .B(out[1503]), .A(rst), .Z(N1515) );
  ANDN U6569 ( .B(out[1504]), .A(rst), .Z(N1516) );
  ANDN U6570 ( .B(out[1505]), .A(rst), .Z(N1517) );
  ANDN U6571 ( .B(out[1506]), .A(rst), .Z(N1518) );
  ANDN U6572 ( .B(out[1507]), .A(rst), .Z(N1519) );
  ANDN U6573 ( .B(out[140]), .A(rst), .Z(N152) );
  ANDN U6574 ( .B(out[1508]), .A(rst), .Z(N1520) );
  ANDN U6575 ( .B(out[1509]), .A(rst), .Z(N1521) );
  ANDN U6576 ( .B(out[1510]), .A(rst), .Z(N1522) );
  ANDN U6577 ( .B(out[1511]), .A(rst), .Z(N1523) );
  ANDN U6578 ( .B(out[1512]), .A(rst), .Z(N1524) );
  ANDN U6579 ( .B(out[1513]), .A(rst), .Z(N1525) );
  ANDN U6580 ( .B(out[1514]), .A(rst), .Z(N1526) );
  ANDN U6581 ( .B(out[1515]), .A(rst), .Z(N1527) );
  ANDN U6582 ( .B(out[1516]), .A(rst), .Z(N1528) );
  ANDN U6583 ( .B(out[1517]), .A(rst), .Z(N1529) );
  ANDN U6584 ( .B(out[141]), .A(rst), .Z(N153) );
  ANDN U6585 ( .B(out[1518]), .A(rst), .Z(N1530) );
  ANDN U6586 ( .B(out[1519]), .A(rst), .Z(N1531) );
  ANDN U6587 ( .B(out[1520]), .A(rst), .Z(N1532) );
  ANDN U6588 ( .B(out[1521]), .A(rst), .Z(N1533) );
  ANDN U6589 ( .B(out[1522]), .A(rst), .Z(N1534) );
  ANDN U6590 ( .B(out[1523]), .A(rst), .Z(N1535) );
  ANDN U6591 ( .B(out[1524]), .A(rst), .Z(N1536) );
  ANDN U6592 ( .B(out[1525]), .A(rst), .Z(N1537) );
  ANDN U6593 ( .B(out[1526]), .A(rst), .Z(N1538) );
  ANDN U6594 ( .B(out[1527]), .A(rst), .Z(N1539) );
  ANDN U6595 ( .B(out[142]), .A(rst), .Z(N154) );
  ANDN U6596 ( .B(out[1528]), .A(rst), .Z(N1540) );
  ANDN U6597 ( .B(out[1529]), .A(rst), .Z(N1541) );
  ANDN U6598 ( .B(out[1530]), .A(rst), .Z(N1542) );
  ANDN U6599 ( .B(out[1531]), .A(rst), .Z(N1543) );
  ANDN U6600 ( .B(out[1532]), .A(rst), .Z(N1544) );
  ANDN U6601 ( .B(out[1533]), .A(rst), .Z(N1545) );
  ANDN U6602 ( .B(out[1534]), .A(rst), .Z(N1546) );
  ANDN U6603 ( .B(out[1535]), .A(rst), .Z(N1547) );
  ANDN U6604 ( .B(out[1536]), .A(rst), .Z(N1548) );
  ANDN U6605 ( .B(out[1537]), .A(rst), .Z(N1549) );
  ANDN U6606 ( .B(out[143]), .A(rst), .Z(N155) );
  ANDN U6607 ( .B(out[1538]), .A(rst), .Z(N1550) );
  ANDN U6608 ( .B(out[1539]), .A(rst), .Z(N1551) );
  ANDN U6609 ( .B(out[1540]), .A(rst), .Z(N1552) );
  ANDN U6610 ( .B(out[1541]), .A(rst), .Z(N1553) );
  ANDN U6611 ( .B(out[1542]), .A(rst), .Z(N1554) );
  ANDN U6612 ( .B(out[1543]), .A(rst), .Z(N1555) );
  ANDN U6613 ( .B(out[1544]), .A(rst), .Z(N1556) );
  ANDN U6614 ( .B(out[1545]), .A(rst), .Z(N1557) );
  ANDN U6615 ( .B(out[1546]), .A(rst), .Z(N1558) );
  ANDN U6616 ( .B(out[1547]), .A(rst), .Z(N1559) );
  ANDN U6617 ( .B(out[144]), .A(rst), .Z(N156) );
  ANDN U6618 ( .B(out[1548]), .A(rst), .Z(N1560) );
  ANDN U6619 ( .B(out[1549]), .A(rst), .Z(N1561) );
  ANDN U6620 ( .B(out[1550]), .A(rst), .Z(N1562) );
  ANDN U6621 ( .B(out[1551]), .A(rst), .Z(N1563) );
  ANDN U6622 ( .B(out[1552]), .A(rst), .Z(N1564) );
  ANDN U6623 ( .B(out[1553]), .A(rst), .Z(N1565) );
  ANDN U6624 ( .B(out[1554]), .A(rst), .Z(N1566) );
  ANDN U6625 ( .B(out[1555]), .A(rst), .Z(N1567) );
  ANDN U6626 ( .B(out[1556]), .A(rst), .Z(N1568) );
  ANDN U6627 ( .B(out[1557]), .A(rst), .Z(N1569) );
  ANDN U6628 ( .B(out[145]), .A(rst), .Z(N157) );
  ANDN U6629 ( .B(out[1558]), .A(rst), .Z(N1570) );
  ANDN U6630 ( .B(out[1559]), .A(rst), .Z(N1571) );
  ANDN U6631 ( .B(out[1560]), .A(rst), .Z(N1572) );
  ANDN U6632 ( .B(out[1561]), .A(rst), .Z(N1573) );
  ANDN U6633 ( .B(out[1562]), .A(rst), .Z(N1574) );
  ANDN U6634 ( .B(out[1563]), .A(rst), .Z(N1575) );
  ANDN U6635 ( .B(out[1564]), .A(rst), .Z(N1576) );
  ANDN U6636 ( .B(out[1565]), .A(rst), .Z(N1577) );
  ANDN U6637 ( .B(out[1566]), .A(rst), .Z(N1578) );
  ANDN U6638 ( .B(out[1567]), .A(rst), .Z(N1579) );
  ANDN U6639 ( .B(out[146]), .A(rst), .Z(N158) );
  ANDN U6640 ( .B(out[1568]), .A(rst), .Z(N1580) );
  ANDN U6641 ( .B(out[1569]), .A(rst), .Z(N1581) );
  ANDN U6642 ( .B(out[1570]), .A(rst), .Z(N1582) );
  ANDN U6643 ( .B(out[1571]), .A(rst), .Z(N1583) );
  ANDN U6644 ( .B(out[1572]), .A(rst), .Z(N1584) );
  ANDN U6645 ( .B(out[1573]), .A(rst), .Z(N1585) );
  ANDN U6646 ( .B(out[1574]), .A(rst), .Z(N1586) );
  ANDN U6647 ( .B(out[1575]), .A(rst), .Z(N1587) );
  ANDN U6648 ( .B(out[1576]), .A(rst), .Z(N1588) );
  ANDN U6649 ( .B(out[1577]), .A(rst), .Z(N1589) );
  ANDN U6650 ( .B(out[147]), .A(rst), .Z(N159) );
  ANDN U6651 ( .B(out[1578]), .A(rst), .Z(N1590) );
  ANDN U6652 ( .B(out[1579]), .A(rst), .Z(N1591) );
  ANDN U6653 ( .B(out[1580]), .A(rst), .Z(N1592) );
  ANDN U6654 ( .B(out[1581]), .A(rst), .Z(N1593) );
  ANDN U6655 ( .B(out[1582]), .A(rst), .Z(N1594) );
  ANDN U6656 ( .B(out[1583]), .A(rst), .Z(N1595) );
  ANDN U6657 ( .B(out[1584]), .A(rst), .Z(N1596) );
  ANDN U6658 ( .B(out[1585]), .A(rst), .Z(N1597) );
  ANDN U6659 ( .B(out[1586]), .A(rst), .Z(N1598) );
  ANDN U6660 ( .B(out[1587]), .A(rst), .Z(N1599) );
  ANDN U6661 ( .B(out[4]), .A(rst), .Z(N16) );
  ANDN U6662 ( .B(out[148]), .A(rst), .Z(N160) );
  ANDN U6663 ( .B(out[1588]), .A(rst), .Z(N1600) );
  ANDN U6664 ( .B(out[1589]), .A(rst), .Z(N1601) );
  ANDN U6665 ( .B(out[1590]), .A(rst), .Z(N1602) );
  ANDN U6666 ( .B(out[1591]), .A(rst), .Z(N1603) );
  ANDN U6667 ( .B(out[1592]), .A(rst), .Z(N1604) );
  ANDN U6668 ( .B(out[1593]), .A(rst), .Z(N1605) );
  ANDN U6669 ( .B(out[1594]), .A(rst), .Z(N1606) );
  ANDN U6670 ( .B(out[1595]), .A(rst), .Z(N1607) );
  ANDN U6671 ( .B(out[1596]), .A(rst), .Z(N1608) );
  ANDN U6672 ( .B(out[1597]), .A(rst), .Z(N1609) );
  ANDN U6673 ( .B(out[149]), .A(rst), .Z(N161) );
  ANDN U6674 ( .B(out[1598]), .A(rst), .Z(N1610) );
  ANDN U6675 ( .B(out[1599]), .A(rst), .Z(N1611) );
  ANDN U6676 ( .B(out[150]), .A(rst), .Z(N162) );
  ANDN U6677 ( .B(out[151]), .A(rst), .Z(N163) );
  ANDN U6678 ( .B(out[152]), .A(rst), .Z(N164) );
  ANDN U6679 ( .B(out[153]), .A(rst), .Z(N165) );
  ANDN U6680 ( .B(out[154]), .A(rst), .Z(N166) );
  ANDN U6681 ( .B(out[155]), .A(rst), .Z(N167) );
  ANDN U6682 ( .B(out[156]), .A(rst), .Z(N168) );
  ANDN U6683 ( .B(out[157]), .A(rst), .Z(N169) );
  ANDN U6684 ( .B(out[5]), .A(rst), .Z(N17) );
  ANDN U6685 ( .B(out[158]), .A(rst), .Z(N170) );
  ANDN U6686 ( .B(out[159]), .A(rst), .Z(N171) );
  ANDN U6687 ( .B(out[160]), .A(rst), .Z(N172) );
  ANDN U6688 ( .B(out[161]), .A(rst), .Z(N173) );
  ANDN U6689 ( .B(out[162]), .A(rst), .Z(N174) );
  ANDN U6690 ( .B(out[163]), .A(rst), .Z(N175) );
  ANDN U6691 ( .B(out[164]), .A(rst), .Z(N176) );
  ANDN U6692 ( .B(out[165]), .A(rst), .Z(N177) );
  ANDN U6693 ( .B(out[166]), .A(rst), .Z(N178) );
  ANDN U6694 ( .B(out[167]), .A(rst), .Z(N179) );
  ANDN U6695 ( .B(out[6]), .A(rst), .Z(N18) );
  ANDN U6696 ( .B(out[168]), .A(rst), .Z(N180) );
  ANDN U6697 ( .B(out[169]), .A(rst), .Z(N181) );
  ANDN U6698 ( .B(out[170]), .A(rst), .Z(N182) );
  ANDN U6699 ( .B(out[171]), .A(rst), .Z(N183) );
  ANDN U6700 ( .B(out[172]), .A(rst), .Z(N184) );
  ANDN U6701 ( .B(out[173]), .A(rst), .Z(N185) );
  ANDN U6702 ( .B(out[174]), .A(rst), .Z(N186) );
  ANDN U6703 ( .B(out[175]), .A(rst), .Z(N187) );
  ANDN U6704 ( .B(out[176]), .A(rst), .Z(N188) );
  ANDN U6705 ( .B(out[177]), .A(rst), .Z(N189) );
  ANDN U6706 ( .B(out[7]), .A(rst), .Z(N19) );
  ANDN U6707 ( .B(out[178]), .A(rst), .Z(N190) );
  ANDN U6708 ( .B(out[179]), .A(rst), .Z(N191) );
  ANDN U6709 ( .B(out[180]), .A(rst), .Z(N192) );
  ANDN U6710 ( .B(out[181]), .A(rst), .Z(N193) );
  ANDN U6711 ( .B(out[182]), .A(rst), .Z(N194) );
  ANDN U6712 ( .B(out[183]), .A(rst), .Z(N195) );
  ANDN U6713 ( .B(out[184]), .A(rst), .Z(N196) );
  ANDN U6714 ( .B(out[185]), .A(rst), .Z(N197) );
  ANDN U6715 ( .B(out[186]), .A(rst), .Z(N198) );
  ANDN U6716 ( .B(out[187]), .A(rst), .Z(N199) );
  ANDN U6717 ( .B(out[8]), .A(rst), .Z(N20) );
  ANDN U6718 ( .B(out[188]), .A(rst), .Z(N200) );
  ANDN U6719 ( .B(out[189]), .A(rst), .Z(N201) );
  ANDN U6720 ( .B(out[190]), .A(rst), .Z(N202) );
  ANDN U6721 ( .B(out[191]), .A(rst), .Z(N203) );
  ANDN U6722 ( .B(out[192]), .A(rst), .Z(N204) );
  ANDN U6723 ( .B(out[193]), .A(rst), .Z(N205) );
  ANDN U6724 ( .B(out[194]), .A(rst), .Z(N206) );
  ANDN U6725 ( .B(out[195]), .A(rst), .Z(N207) );
  ANDN U6726 ( .B(out[196]), .A(rst), .Z(N208) );
  ANDN U6727 ( .B(out[197]), .A(rst), .Z(N209) );
  ANDN U6728 ( .B(out[9]), .A(rst), .Z(N21) );
  ANDN U6729 ( .B(out[198]), .A(rst), .Z(N210) );
  ANDN U6730 ( .B(out[199]), .A(rst), .Z(N211) );
  ANDN U6731 ( .B(out[200]), .A(rst), .Z(N212) );
  ANDN U6732 ( .B(out[201]), .A(rst), .Z(N213) );
  ANDN U6733 ( .B(out[202]), .A(rst), .Z(N214) );
  ANDN U6734 ( .B(out[203]), .A(rst), .Z(N215) );
  ANDN U6735 ( .B(out[204]), .A(rst), .Z(N216) );
  ANDN U6736 ( .B(out[205]), .A(rst), .Z(N217) );
  ANDN U6737 ( .B(out[206]), .A(rst), .Z(N218) );
  ANDN U6738 ( .B(out[207]), .A(rst), .Z(N219) );
  ANDN U6739 ( .B(out[10]), .A(rst), .Z(N22) );
  ANDN U6740 ( .B(out[208]), .A(rst), .Z(N220) );
  ANDN U6741 ( .B(out[209]), .A(rst), .Z(N221) );
  ANDN U6742 ( .B(out[210]), .A(rst), .Z(N222) );
  ANDN U6743 ( .B(out[211]), .A(rst), .Z(N223) );
  ANDN U6744 ( .B(out[212]), .A(rst), .Z(N224) );
  ANDN U6745 ( .B(out[213]), .A(rst), .Z(N225) );
  ANDN U6746 ( .B(out[214]), .A(rst), .Z(N226) );
  ANDN U6747 ( .B(out[215]), .A(rst), .Z(N227) );
  ANDN U6748 ( .B(out[216]), .A(rst), .Z(N228) );
  ANDN U6749 ( .B(out[217]), .A(rst), .Z(N229) );
  ANDN U6750 ( .B(out[11]), .A(rst), .Z(N23) );
  ANDN U6751 ( .B(out[218]), .A(rst), .Z(N230) );
  ANDN U6752 ( .B(out[219]), .A(rst), .Z(N231) );
  ANDN U6753 ( .B(out[220]), .A(rst), .Z(N232) );
  ANDN U6754 ( .B(out[221]), .A(rst), .Z(N233) );
  ANDN U6755 ( .B(out[222]), .A(rst), .Z(N234) );
  ANDN U6756 ( .B(out[223]), .A(rst), .Z(N235) );
  ANDN U6757 ( .B(out[224]), .A(rst), .Z(N236) );
  ANDN U6758 ( .B(out[225]), .A(rst), .Z(N237) );
  ANDN U6759 ( .B(out[226]), .A(rst), .Z(N238) );
  ANDN U6760 ( .B(out[227]), .A(rst), .Z(N239) );
  ANDN U6761 ( .B(out[12]), .A(rst), .Z(N24) );
  ANDN U6762 ( .B(out[228]), .A(rst), .Z(N240) );
  ANDN U6763 ( .B(out[229]), .A(rst), .Z(N241) );
  ANDN U6764 ( .B(out[230]), .A(rst), .Z(N242) );
  ANDN U6765 ( .B(out[231]), .A(rst), .Z(N243) );
  ANDN U6766 ( .B(out[232]), .A(rst), .Z(N244) );
  ANDN U6767 ( .B(out[233]), .A(rst), .Z(N245) );
  ANDN U6768 ( .B(out[234]), .A(rst), .Z(N246) );
  ANDN U6769 ( .B(out[235]), .A(rst), .Z(N247) );
  ANDN U6770 ( .B(out[236]), .A(rst), .Z(N248) );
  ANDN U6771 ( .B(out[237]), .A(rst), .Z(N249) );
  ANDN U6772 ( .B(out[13]), .A(rst), .Z(N25) );
  ANDN U6773 ( .B(out[238]), .A(rst), .Z(N250) );
  ANDN U6774 ( .B(out[239]), .A(rst), .Z(N251) );
  ANDN U6775 ( .B(out[240]), .A(rst), .Z(N252) );
  ANDN U6776 ( .B(out[241]), .A(rst), .Z(N253) );
  ANDN U6777 ( .B(out[242]), .A(rst), .Z(N254) );
  ANDN U6778 ( .B(out[243]), .A(rst), .Z(N255) );
  ANDN U6779 ( .B(out[244]), .A(rst), .Z(N256) );
  ANDN U6780 ( .B(out[245]), .A(rst), .Z(N257) );
  ANDN U6781 ( .B(out[246]), .A(rst), .Z(N258) );
  ANDN U6782 ( .B(out[247]), .A(rst), .Z(N259) );
  ANDN U6783 ( .B(out[14]), .A(rst), .Z(N26) );
  ANDN U6784 ( .B(out[248]), .A(rst), .Z(N260) );
  ANDN U6785 ( .B(out[249]), .A(rst), .Z(N261) );
  ANDN U6786 ( .B(out[250]), .A(rst), .Z(N262) );
  ANDN U6787 ( .B(out[251]), .A(rst), .Z(N263) );
  ANDN U6788 ( .B(out[252]), .A(rst), .Z(N264) );
  ANDN U6789 ( .B(out[253]), .A(rst), .Z(N265) );
  ANDN U6790 ( .B(out[254]), .A(rst), .Z(N266) );
  ANDN U6791 ( .B(out[255]), .A(rst), .Z(N267) );
  ANDN U6792 ( .B(out[256]), .A(rst), .Z(N268) );
  ANDN U6793 ( .B(out[257]), .A(rst), .Z(N269) );
  ANDN U6794 ( .B(out[15]), .A(rst), .Z(N27) );
  ANDN U6795 ( .B(out[258]), .A(rst), .Z(N270) );
  ANDN U6796 ( .B(out[259]), .A(rst), .Z(N271) );
  ANDN U6797 ( .B(out[260]), .A(rst), .Z(N272) );
  ANDN U6798 ( .B(out[261]), .A(rst), .Z(N273) );
  ANDN U6799 ( .B(out[262]), .A(rst), .Z(N274) );
  ANDN U6800 ( .B(out[263]), .A(rst), .Z(N275) );
  ANDN U6801 ( .B(out[264]), .A(rst), .Z(N276) );
  ANDN U6802 ( .B(out[265]), .A(rst), .Z(N277) );
  ANDN U6803 ( .B(out[266]), .A(rst), .Z(N278) );
  ANDN U6804 ( .B(out[267]), .A(rst), .Z(N279) );
  ANDN U6805 ( .B(out[16]), .A(rst), .Z(N28) );
  ANDN U6806 ( .B(out[268]), .A(rst), .Z(N280) );
  ANDN U6807 ( .B(out[269]), .A(rst), .Z(N281) );
  ANDN U6808 ( .B(out[270]), .A(rst), .Z(N282) );
  ANDN U6809 ( .B(out[271]), .A(rst), .Z(N283) );
  ANDN U6810 ( .B(out[272]), .A(rst), .Z(N284) );
  ANDN U6811 ( .B(out[273]), .A(rst), .Z(N285) );
  ANDN U6812 ( .B(out[274]), .A(rst), .Z(N286) );
  ANDN U6813 ( .B(out[275]), .A(rst), .Z(N287) );
  ANDN U6814 ( .B(out[276]), .A(rst), .Z(N288) );
  ANDN U6815 ( .B(out[277]), .A(rst), .Z(N289) );
  ANDN U6816 ( .B(out[17]), .A(rst), .Z(N29) );
  ANDN U6817 ( .B(out[278]), .A(rst), .Z(N290) );
  ANDN U6818 ( .B(out[279]), .A(rst), .Z(N291) );
  ANDN U6819 ( .B(out[280]), .A(rst), .Z(N292) );
  ANDN U6820 ( .B(out[281]), .A(rst), .Z(N293) );
  ANDN U6821 ( .B(out[282]), .A(rst), .Z(N294) );
  ANDN U6822 ( .B(out[283]), .A(rst), .Z(N295) );
  ANDN U6823 ( .B(out[284]), .A(rst), .Z(N296) );
  ANDN U6824 ( .B(out[285]), .A(rst), .Z(N297) );
  ANDN U6825 ( .B(out[286]), .A(rst), .Z(N298) );
  ANDN U6826 ( .B(out[287]), .A(rst), .Z(N299) );
  ANDN U6827 ( .B(out[18]), .A(rst), .Z(N30) );
  ANDN U6828 ( .B(out[288]), .A(rst), .Z(N300) );
  ANDN U6829 ( .B(out[289]), .A(rst), .Z(N301) );
  ANDN U6830 ( .B(out[290]), .A(rst), .Z(N302) );
  ANDN U6831 ( .B(out[291]), .A(rst), .Z(N303) );
  ANDN U6832 ( .B(out[292]), .A(rst), .Z(N304) );
  ANDN U6833 ( .B(out[293]), .A(rst), .Z(N305) );
  ANDN U6834 ( .B(out[294]), .A(rst), .Z(N306) );
  ANDN U6835 ( .B(out[295]), .A(rst), .Z(N307) );
  ANDN U6836 ( .B(out[296]), .A(rst), .Z(N308) );
  ANDN U6837 ( .B(out[297]), .A(rst), .Z(N309) );
  ANDN U6838 ( .B(out[19]), .A(rst), .Z(N31) );
  ANDN U6839 ( .B(out[298]), .A(rst), .Z(N310) );
  ANDN U6840 ( .B(out[299]), .A(rst), .Z(N311) );
  ANDN U6841 ( .B(out[300]), .A(rst), .Z(N312) );
  ANDN U6842 ( .B(out[301]), .A(rst), .Z(N313) );
  ANDN U6843 ( .B(out[302]), .A(rst), .Z(N314) );
  ANDN U6844 ( .B(out[303]), .A(rst), .Z(N315) );
  ANDN U6845 ( .B(out[304]), .A(rst), .Z(N316) );
  ANDN U6846 ( .B(out[305]), .A(rst), .Z(N317) );
  ANDN U6847 ( .B(out[306]), .A(rst), .Z(N318) );
  ANDN U6848 ( .B(out[307]), .A(rst), .Z(N319) );
  ANDN U6849 ( .B(out[20]), .A(rst), .Z(N32) );
  ANDN U6850 ( .B(out[308]), .A(rst), .Z(N320) );
  ANDN U6851 ( .B(out[309]), .A(rst), .Z(N321) );
  ANDN U6852 ( .B(out[310]), .A(rst), .Z(N322) );
  ANDN U6853 ( .B(out[311]), .A(rst), .Z(N323) );
  ANDN U6854 ( .B(out[312]), .A(rst), .Z(N324) );
  ANDN U6855 ( .B(out[313]), .A(rst), .Z(N325) );
  ANDN U6856 ( .B(out[314]), .A(rst), .Z(N326) );
  ANDN U6857 ( .B(out[315]), .A(rst), .Z(N327) );
  ANDN U6858 ( .B(out[316]), .A(rst), .Z(N328) );
  ANDN U6859 ( .B(out[317]), .A(rst), .Z(N329) );
  ANDN U6860 ( .B(out[21]), .A(rst), .Z(N33) );
  ANDN U6861 ( .B(out[318]), .A(rst), .Z(N330) );
  ANDN U6862 ( .B(out[319]), .A(rst), .Z(N331) );
  ANDN U6863 ( .B(out[320]), .A(rst), .Z(N332) );
  ANDN U6864 ( .B(out[321]), .A(rst), .Z(N333) );
  ANDN U6865 ( .B(out[322]), .A(rst), .Z(N334) );
  ANDN U6866 ( .B(out[323]), .A(rst), .Z(N335) );
  ANDN U6867 ( .B(out[324]), .A(rst), .Z(N336) );
  ANDN U6868 ( .B(out[325]), .A(rst), .Z(N337) );
  ANDN U6869 ( .B(out[326]), .A(rst), .Z(N338) );
  ANDN U6870 ( .B(out[327]), .A(rst), .Z(N339) );
  ANDN U6871 ( .B(out[22]), .A(rst), .Z(N34) );
  ANDN U6872 ( .B(out[328]), .A(rst), .Z(N340) );
  ANDN U6873 ( .B(out[329]), .A(rst), .Z(N341) );
  ANDN U6874 ( .B(out[330]), .A(rst), .Z(N342) );
  ANDN U6875 ( .B(out[331]), .A(rst), .Z(N343) );
  ANDN U6876 ( .B(out[332]), .A(rst), .Z(N344) );
  ANDN U6877 ( .B(out[333]), .A(rst), .Z(N345) );
  ANDN U6878 ( .B(out[334]), .A(rst), .Z(N346) );
  ANDN U6879 ( .B(out[335]), .A(rst), .Z(N347) );
  ANDN U6880 ( .B(out[336]), .A(rst), .Z(N348) );
  ANDN U6881 ( .B(out[337]), .A(rst), .Z(N349) );
  ANDN U6882 ( .B(out[23]), .A(rst), .Z(N35) );
  ANDN U6883 ( .B(out[338]), .A(rst), .Z(N350) );
  ANDN U6884 ( .B(out[339]), .A(rst), .Z(N351) );
  ANDN U6885 ( .B(out[340]), .A(rst), .Z(N352) );
  ANDN U6886 ( .B(out[341]), .A(rst), .Z(N353) );
  ANDN U6887 ( .B(out[342]), .A(rst), .Z(N354) );
  ANDN U6888 ( .B(out[343]), .A(rst), .Z(N355) );
  ANDN U6889 ( .B(out[344]), .A(rst), .Z(N356) );
  ANDN U6890 ( .B(out[345]), .A(rst), .Z(N357) );
  ANDN U6891 ( .B(out[346]), .A(rst), .Z(N358) );
  ANDN U6892 ( .B(out[347]), .A(rst), .Z(N359) );
  ANDN U6893 ( .B(out[24]), .A(rst), .Z(N36) );
  ANDN U6894 ( .B(out[348]), .A(rst), .Z(N360) );
  ANDN U6895 ( .B(out[349]), .A(rst), .Z(N361) );
  ANDN U6896 ( .B(out[350]), .A(rst), .Z(N362) );
  ANDN U6897 ( .B(out[351]), .A(rst), .Z(N363) );
  ANDN U6898 ( .B(out[352]), .A(rst), .Z(N364) );
  ANDN U6899 ( .B(out[353]), .A(rst), .Z(N365) );
  ANDN U6900 ( .B(out[354]), .A(rst), .Z(N366) );
  ANDN U6901 ( .B(out[355]), .A(rst), .Z(N367) );
  ANDN U6902 ( .B(out[356]), .A(rst), .Z(N368) );
  ANDN U6903 ( .B(out[357]), .A(rst), .Z(N369) );
  ANDN U6904 ( .B(out[25]), .A(rst), .Z(N37) );
  ANDN U6905 ( .B(out[358]), .A(rst), .Z(N370) );
  ANDN U6906 ( .B(out[359]), .A(rst), .Z(N371) );
  ANDN U6907 ( .B(out[360]), .A(rst), .Z(N372) );
  ANDN U6908 ( .B(out[361]), .A(rst), .Z(N373) );
  ANDN U6909 ( .B(out[362]), .A(rst), .Z(N374) );
  ANDN U6910 ( .B(out[363]), .A(rst), .Z(N375) );
  ANDN U6911 ( .B(out[364]), .A(rst), .Z(N376) );
  ANDN U6912 ( .B(out[365]), .A(rst), .Z(N377) );
  ANDN U6913 ( .B(out[366]), .A(rst), .Z(N378) );
  ANDN U6914 ( .B(out[367]), .A(rst), .Z(N379) );
  ANDN U6915 ( .B(out[26]), .A(rst), .Z(N38) );
  ANDN U6916 ( .B(out[368]), .A(rst), .Z(N380) );
  ANDN U6917 ( .B(out[369]), .A(rst), .Z(N381) );
  ANDN U6918 ( .B(out[370]), .A(rst), .Z(N382) );
  ANDN U6919 ( .B(out[371]), .A(rst), .Z(N383) );
  ANDN U6920 ( .B(out[372]), .A(rst), .Z(N384) );
  ANDN U6921 ( .B(out[373]), .A(rst), .Z(N385) );
  ANDN U6922 ( .B(out[374]), .A(rst), .Z(N386) );
  ANDN U6923 ( .B(out[375]), .A(rst), .Z(N387) );
  ANDN U6924 ( .B(out[376]), .A(rst), .Z(N388) );
  ANDN U6925 ( .B(out[377]), .A(rst), .Z(N389) );
  ANDN U6926 ( .B(out[27]), .A(rst), .Z(N39) );
  ANDN U6927 ( .B(out[378]), .A(rst), .Z(N390) );
  ANDN U6928 ( .B(out[379]), .A(rst), .Z(N391) );
  ANDN U6929 ( .B(out[380]), .A(rst), .Z(N392) );
  ANDN U6930 ( .B(out[381]), .A(rst), .Z(N393) );
  ANDN U6931 ( .B(out[382]), .A(rst), .Z(N394) );
  ANDN U6932 ( .B(out[383]), .A(rst), .Z(N395) );
  ANDN U6933 ( .B(out[384]), .A(rst), .Z(N396) );
  ANDN U6934 ( .B(out[385]), .A(rst), .Z(N397) );
  ANDN U6935 ( .B(out[386]), .A(rst), .Z(N398) );
  ANDN U6936 ( .B(out[387]), .A(rst), .Z(N399) );
  ANDN U6937 ( .B(out[28]), .A(rst), .Z(N40) );
  ANDN U6938 ( .B(out[388]), .A(rst), .Z(N400) );
  ANDN U6939 ( .B(out[389]), .A(rst), .Z(N401) );
  ANDN U6940 ( .B(out[390]), .A(rst), .Z(N402) );
  ANDN U6941 ( .B(out[391]), .A(rst), .Z(N403) );
  ANDN U6942 ( .B(out[392]), .A(rst), .Z(N404) );
  ANDN U6943 ( .B(out[393]), .A(rst), .Z(N405) );
  ANDN U6944 ( .B(out[394]), .A(rst), .Z(N406) );
  ANDN U6945 ( .B(out[395]), .A(rst), .Z(N407) );
  ANDN U6946 ( .B(out[396]), .A(rst), .Z(N408) );
  ANDN U6947 ( .B(out[397]), .A(rst), .Z(N409) );
  ANDN U6948 ( .B(out[29]), .A(rst), .Z(N41) );
  ANDN U6949 ( .B(out[398]), .A(rst), .Z(N410) );
  ANDN U6950 ( .B(out[399]), .A(rst), .Z(N411) );
  ANDN U6951 ( .B(out[400]), .A(rst), .Z(N412) );
  ANDN U6952 ( .B(out[401]), .A(rst), .Z(N413) );
  ANDN U6953 ( .B(out[402]), .A(rst), .Z(N414) );
  ANDN U6954 ( .B(out[403]), .A(rst), .Z(N415) );
  ANDN U6955 ( .B(out[404]), .A(rst), .Z(N416) );
  ANDN U6956 ( .B(out[405]), .A(rst), .Z(N417) );
  ANDN U6957 ( .B(out[406]), .A(rst), .Z(N418) );
  ANDN U6958 ( .B(out[407]), .A(rst), .Z(N419) );
  ANDN U6959 ( .B(out[30]), .A(rst), .Z(N42) );
  ANDN U6960 ( .B(out[408]), .A(rst), .Z(N420) );
  ANDN U6961 ( .B(out[409]), .A(rst), .Z(N421) );
  ANDN U6962 ( .B(out[410]), .A(rst), .Z(N422) );
  ANDN U6963 ( .B(out[411]), .A(rst), .Z(N423) );
  ANDN U6964 ( .B(out[412]), .A(rst), .Z(N424) );
  ANDN U6965 ( .B(out[413]), .A(rst), .Z(N425) );
  ANDN U6966 ( .B(out[414]), .A(rst), .Z(N426) );
  ANDN U6967 ( .B(out[415]), .A(rst), .Z(N427) );
  ANDN U6968 ( .B(out[416]), .A(rst), .Z(N428) );
  ANDN U6969 ( .B(out[417]), .A(rst), .Z(N429) );
  ANDN U6970 ( .B(out[31]), .A(rst), .Z(N43) );
  ANDN U6971 ( .B(out[418]), .A(rst), .Z(N430) );
  ANDN U6972 ( .B(out[419]), .A(rst), .Z(N431) );
  ANDN U6973 ( .B(out[420]), .A(rst), .Z(N432) );
  ANDN U6974 ( .B(out[421]), .A(rst), .Z(N433) );
  ANDN U6975 ( .B(out[422]), .A(rst), .Z(N434) );
  ANDN U6976 ( .B(out[423]), .A(rst), .Z(N435) );
  ANDN U6977 ( .B(out[424]), .A(rst), .Z(N436) );
  ANDN U6978 ( .B(out[425]), .A(rst), .Z(N437) );
  ANDN U6979 ( .B(out[426]), .A(rst), .Z(N438) );
  ANDN U6980 ( .B(out[427]), .A(rst), .Z(N439) );
  ANDN U6981 ( .B(out[32]), .A(rst), .Z(N44) );
  ANDN U6982 ( .B(out[428]), .A(rst), .Z(N440) );
  ANDN U6983 ( .B(out[429]), .A(rst), .Z(N441) );
  ANDN U6984 ( .B(out[430]), .A(rst), .Z(N442) );
  ANDN U6985 ( .B(out[431]), .A(rst), .Z(N443) );
  ANDN U6986 ( .B(out[432]), .A(rst), .Z(N444) );
  ANDN U6987 ( .B(out[433]), .A(rst), .Z(N445) );
  ANDN U6988 ( .B(out[434]), .A(rst), .Z(N446) );
  ANDN U6989 ( .B(out[435]), .A(rst), .Z(N447) );
  ANDN U6990 ( .B(out[436]), .A(rst), .Z(N448) );
  ANDN U6991 ( .B(out[437]), .A(rst), .Z(N449) );
  ANDN U6992 ( .B(out[33]), .A(rst), .Z(N45) );
  ANDN U6993 ( .B(out[438]), .A(rst), .Z(N450) );
  ANDN U6994 ( .B(out[439]), .A(rst), .Z(N451) );
  ANDN U6995 ( .B(out[440]), .A(rst), .Z(N452) );
  ANDN U6996 ( .B(out[441]), .A(rst), .Z(N453) );
  ANDN U6997 ( .B(out[442]), .A(rst), .Z(N454) );
  ANDN U6998 ( .B(out[443]), .A(rst), .Z(N455) );
  ANDN U6999 ( .B(out[444]), .A(rst), .Z(N456) );
  ANDN U7000 ( .B(out[445]), .A(rst), .Z(N457) );
  ANDN U7001 ( .B(out[446]), .A(rst), .Z(N458) );
  ANDN U7002 ( .B(out[447]), .A(rst), .Z(N459) );
  ANDN U7003 ( .B(out[34]), .A(rst), .Z(N46) );
  ANDN U7004 ( .B(out[448]), .A(rst), .Z(N460) );
  ANDN U7005 ( .B(out[449]), .A(rst), .Z(N461) );
  ANDN U7006 ( .B(out[450]), .A(rst), .Z(N462) );
  ANDN U7007 ( .B(out[451]), .A(rst), .Z(N463) );
  ANDN U7008 ( .B(out[452]), .A(rst), .Z(N464) );
  ANDN U7009 ( .B(out[453]), .A(rst), .Z(N465) );
  ANDN U7010 ( .B(out[454]), .A(rst), .Z(N466) );
  ANDN U7011 ( .B(out[455]), .A(rst), .Z(N467) );
  ANDN U7012 ( .B(out[456]), .A(rst), .Z(N468) );
  ANDN U7013 ( .B(out[457]), .A(rst), .Z(N469) );
  ANDN U7014 ( .B(out[35]), .A(rst), .Z(N47) );
  ANDN U7015 ( .B(out[458]), .A(rst), .Z(N470) );
  ANDN U7016 ( .B(out[459]), .A(rst), .Z(N471) );
  ANDN U7017 ( .B(out[460]), .A(rst), .Z(N472) );
  ANDN U7018 ( .B(out[461]), .A(rst), .Z(N473) );
  ANDN U7019 ( .B(out[462]), .A(rst), .Z(N474) );
  ANDN U7020 ( .B(out[463]), .A(rst), .Z(N475) );
  ANDN U7021 ( .B(out[464]), .A(rst), .Z(N476) );
  ANDN U7022 ( .B(out[465]), .A(rst), .Z(N477) );
  ANDN U7023 ( .B(out[466]), .A(rst), .Z(N478) );
  ANDN U7024 ( .B(out[467]), .A(rst), .Z(N479) );
  ANDN U7025 ( .B(out[36]), .A(rst), .Z(N48) );
  ANDN U7026 ( .B(out[468]), .A(rst), .Z(N480) );
  ANDN U7027 ( .B(out[469]), .A(rst), .Z(N481) );
  ANDN U7028 ( .B(out[470]), .A(rst), .Z(N482) );
  ANDN U7029 ( .B(out[471]), .A(rst), .Z(N483) );
  ANDN U7030 ( .B(out[472]), .A(rst), .Z(N484) );
  ANDN U7031 ( .B(out[473]), .A(rst), .Z(N485) );
  ANDN U7032 ( .B(out[474]), .A(rst), .Z(N486) );
  ANDN U7033 ( .B(out[475]), .A(rst), .Z(N487) );
  ANDN U7034 ( .B(out[476]), .A(rst), .Z(N488) );
  ANDN U7035 ( .B(out[477]), .A(rst), .Z(N489) );
  ANDN U7036 ( .B(out[37]), .A(rst), .Z(N49) );
  ANDN U7037 ( .B(out[478]), .A(rst), .Z(N490) );
  ANDN U7038 ( .B(out[479]), .A(rst), .Z(N491) );
  ANDN U7039 ( .B(out[480]), .A(rst), .Z(N492) );
  ANDN U7040 ( .B(out[481]), .A(rst), .Z(N493) );
  ANDN U7041 ( .B(out[482]), .A(rst), .Z(N494) );
  ANDN U7042 ( .B(out[483]), .A(rst), .Z(N495) );
  ANDN U7043 ( .B(out[484]), .A(rst), .Z(N496) );
  ANDN U7044 ( .B(out[485]), .A(rst), .Z(N497) );
  ANDN U7045 ( .B(out[486]), .A(rst), .Z(N498) );
  ANDN U7046 ( .B(out[487]), .A(rst), .Z(N499) );
  ANDN U7047 ( .B(out[38]), .A(rst), .Z(N50) );
  ANDN U7048 ( .B(out[488]), .A(rst), .Z(N500) );
  ANDN U7049 ( .B(out[489]), .A(rst), .Z(N501) );
  ANDN U7050 ( .B(out[490]), .A(rst), .Z(N502) );
  ANDN U7051 ( .B(out[491]), .A(rst), .Z(N503) );
  ANDN U7052 ( .B(out[492]), .A(rst), .Z(N504) );
  ANDN U7053 ( .B(out[493]), .A(rst), .Z(N505) );
  ANDN U7054 ( .B(out[494]), .A(rst), .Z(N506) );
  ANDN U7055 ( .B(out[495]), .A(rst), .Z(N507) );
  ANDN U7056 ( .B(out[496]), .A(rst), .Z(N508) );
  ANDN U7057 ( .B(out[497]), .A(rst), .Z(N509) );
  ANDN U7058 ( .B(out[39]), .A(rst), .Z(N51) );
  ANDN U7059 ( .B(out[498]), .A(rst), .Z(N510) );
  ANDN U7060 ( .B(out[499]), .A(rst), .Z(N511) );
  ANDN U7061 ( .B(out[500]), .A(rst), .Z(N512) );
  ANDN U7062 ( .B(out[501]), .A(rst), .Z(N513) );
  ANDN U7063 ( .B(out[502]), .A(rst), .Z(N514) );
  ANDN U7064 ( .B(out[503]), .A(rst), .Z(N515) );
  ANDN U7065 ( .B(out[504]), .A(rst), .Z(N516) );
  ANDN U7066 ( .B(out[505]), .A(rst), .Z(N517) );
  ANDN U7067 ( .B(out[506]), .A(rst), .Z(N518) );
  ANDN U7068 ( .B(out[507]), .A(rst), .Z(N519) );
  ANDN U7069 ( .B(out[40]), .A(rst), .Z(N52) );
  ANDN U7070 ( .B(out[508]), .A(rst), .Z(N520) );
  ANDN U7071 ( .B(out[509]), .A(rst), .Z(N521) );
  ANDN U7072 ( .B(out[510]), .A(rst), .Z(N522) );
  ANDN U7073 ( .B(out[511]), .A(rst), .Z(N523) );
  ANDN U7074 ( .B(out[512]), .A(rst), .Z(N524) );
  ANDN U7075 ( .B(out[513]), .A(rst), .Z(N525) );
  ANDN U7076 ( .B(out[514]), .A(rst), .Z(N526) );
  ANDN U7077 ( .B(out[515]), .A(rst), .Z(N527) );
  ANDN U7078 ( .B(out[516]), .A(rst), .Z(N528) );
  ANDN U7079 ( .B(out[517]), .A(rst), .Z(N529) );
  ANDN U7080 ( .B(out[41]), .A(rst), .Z(N53) );
  ANDN U7081 ( .B(out[518]), .A(rst), .Z(N530) );
  ANDN U7082 ( .B(out[519]), .A(rst), .Z(N531) );
  ANDN U7083 ( .B(out[520]), .A(rst), .Z(N532) );
  ANDN U7084 ( .B(out[521]), .A(rst), .Z(N533) );
  ANDN U7085 ( .B(out[522]), .A(rst), .Z(N534) );
  ANDN U7086 ( .B(out[523]), .A(rst), .Z(N535) );
  ANDN U7087 ( .B(out[524]), .A(rst), .Z(N536) );
  ANDN U7088 ( .B(out[525]), .A(rst), .Z(N537) );
  ANDN U7089 ( .B(out[526]), .A(rst), .Z(N538) );
  ANDN U7090 ( .B(out[527]), .A(rst), .Z(N539) );
  ANDN U7091 ( .B(out[42]), .A(rst), .Z(N54) );
  ANDN U7092 ( .B(out[528]), .A(rst), .Z(N540) );
  ANDN U7093 ( .B(out[529]), .A(rst), .Z(N541) );
  ANDN U7094 ( .B(out[530]), .A(rst), .Z(N542) );
  ANDN U7095 ( .B(out[531]), .A(rst), .Z(N543) );
  ANDN U7096 ( .B(out[532]), .A(rst), .Z(N544) );
  ANDN U7097 ( .B(out[533]), .A(rst), .Z(N545) );
  ANDN U7098 ( .B(out[534]), .A(rst), .Z(N546) );
  ANDN U7099 ( .B(out[535]), .A(rst), .Z(N547) );
  ANDN U7100 ( .B(out[536]), .A(rst), .Z(N548) );
  ANDN U7101 ( .B(out[537]), .A(rst), .Z(N549) );
  ANDN U7102 ( .B(out[43]), .A(rst), .Z(N55) );
  ANDN U7103 ( .B(out[538]), .A(rst), .Z(N550) );
  ANDN U7104 ( .B(out[539]), .A(rst), .Z(N551) );
  ANDN U7105 ( .B(out[540]), .A(rst), .Z(N552) );
  ANDN U7106 ( .B(out[541]), .A(rst), .Z(N553) );
  ANDN U7107 ( .B(out[542]), .A(rst), .Z(N554) );
  ANDN U7108 ( .B(out[543]), .A(rst), .Z(N555) );
  ANDN U7109 ( .B(out[544]), .A(rst), .Z(N556) );
  ANDN U7110 ( .B(out[545]), .A(rst), .Z(N557) );
  ANDN U7111 ( .B(out[546]), .A(rst), .Z(N558) );
  ANDN U7112 ( .B(out[547]), .A(rst), .Z(N559) );
  ANDN U7113 ( .B(out[44]), .A(rst), .Z(N56) );
  ANDN U7114 ( .B(out[548]), .A(rst), .Z(N560) );
  ANDN U7115 ( .B(out[549]), .A(rst), .Z(N561) );
  ANDN U7116 ( .B(out[550]), .A(rst), .Z(N562) );
  ANDN U7117 ( .B(out[551]), .A(rst), .Z(N563) );
  ANDN U7118 ( .B(out[552]), .A(rst), .Z(N564) );
  ANDN U7119 ( .B(out[553]), .A(rst), .Z(N565) );
  ANDN U7120 ( .B(out[554]), .A(rst), .Z(N566) );
  ANDN U7121 ( .B(out[555]), .A(rst), .Z(N567) );
  ANDN U7122 ( .B(out[556]), .A(rst), .Z(N568) );
  ANDN U7123 ( .B(out[557]), .A(rst), .Z(N569) );
  ANDN U7124 ( .B(out[45]), .A(rst), .Z(N57) );
  ANDN U7125 ( .B(out[558]), .A(rst), .Z(N570) );
  ANDN U7126 ( .B(out[559]), .A(rst), .Z(N571) );
  ANDN U7127 ( .B(out[560]), .A(rst), .Z(N572) );
  ANDN U7128 ( .B(out[561]), .A(rst), .Z(N573) );
  ANDN U7129 ( .B(out[562]), .A(rst), .Z(N574) );
  ANDN U7130 ( .B(out[563]), .A(rst), .Z(N575) );
  ANDN U7131 ( .B(out[564]), .A(rst), .Z(N576) );
  ANDN U7132 ( .B(out[565]), .A(rst), .Z(N577) );
  ANDN U7133 ( .B(out[566]), .A(rst), .Z(N578) );
  ANDN U7134 ( .B(out[567]), .A(rst), .Z(N579) );
  ANDN U7135 ( .B(out[46]), .A(rst), .Z(N58) );
  ANDN U7136 ( .B(out[568]), .A(rst), .Z(N580) );
  ANDN U7137 ( .B(out[569]), .A(rst), .Z(N581) );
  ANDN U7138 ( .B(out[570]), .A(rst), .Z(N582) );
  ANDN U7139 ( .B(out[571]), .A(rst), .Z(N583) );
  ANDN U7140 ( .B(out[572]), .A(rst), .Z(N584) );
  ANDN U7141 ( .B(out[573]), .A(rst), .Z(N585) );
  ANDN U7142 ( .B(out[574]), .A(rst), .Z(N586) );
  ANDN U7143 ( .B(out[575]), .A(rst), .Z(N587) );
  ANDN U7144 ( .B(out[576]), .A(rst), .Z(N588) );
  ANDN U7145 ( .B(out[577]), .A(rst), .Z(N589) );
  ANDN U7146 ( .B(out[47]), .A(rst), .Z(N59) );
  ANDN U7147 ( .B(out[578]), .A(rst), .Z(N590) );
  ANDN U7148 ( .B(out[579]), .A(rst), .Z(N591) );
  ANDN U7149 ( .B(out[580]), .A(rst), .Z(N592) );
  ANDN U7150 ( .B(out[581]), .A(rst), .Z(N593) );
  ANDN U7151 ( .B(out[582]), .A(rst), .Z(N594) );
  ANDN U7152 ( .B(out[583]), .A(rst), .Z(N595) );
  ANDN U7153 ( .B(out[584]), .A(rst), .Z(N596) );
  ANDN U7154 ( .B(out[585]), .A(rst), .Z(N597) );
  ANDN U7155 ( .B(out[586]), .A(rst), .Z(N598) );
  ANDN U7156 ( .B(out[587]), .A(rst), .Z(N599) );
  NOR U7157 ( .A(rst), .B(init), .Z(N6) );
  ANDN U7158 ( .B(out[48]), .A(rst), .Z(N60) );
  ANDN U7159 ( .B(out[588]), .A(rst), .Z(N600) );
  ANDN U7160 ( .B(out[589]), .A(rst), .Z(N601) );
  ANDN U7161 ( .B(out[590]), .A(rst), .Z(N602) );
  ANDN U7162 ( .B(out[591]), .A(rst), .Z(N603) );
  ANDN U7163 ( .B(out[592]), .A(rst), .Z(N604) );
  ANDN U7164 ( .B(out[593]), .A(rst), .Z(N605) );
  ANDN U7165 ( .B(out[594]), .A(rst), .Z(N606) );
  ANDN U7166 ( .B(out[595]), .A(rst), .Z(N607) );
  ANDN U7167 ( .B(out[596]), .A(rst), .Z(N608) );
  ANDN U7168 ( .B(out[597]), .A(rst), .Z(N609) );
  ANDN U7169 ( .B(out[49]), .A(rst), .Z(N61) );
  ANDN U7170 ( .B(out[598]), .A(rst), .Z(N610) );
  ANDN U7171 ( .B(out[599]), .A(rst), .Z(N611) );
  ANDN U7172 ( .B(out[600]), .A(rst), .Z(N612) );
  ANDN U7173 ( .B(out[601]), .A(rst), .Z(N613) );
  ANDN U7174 ( .B(out[602]), .A(rst), .Z(N614) );
  ANDN U7175 ( .B(out[603]), .A(rst), .Z(N615) );
  ANDN U7176 ( .B(out[604]), .A(rst), .Z(N616) );
  ANDN U7177 ( .B(out[605]), .A(rst), .Z(N617) );
  ANDN U7178 ( .B(out[606]), .A(rst), .Z(N618) );
  ANDN U7179 ( .B(out[607]), .A(rst), .Z(N619) );
  ANDN U7180 ( .B(out[50]), .A(rst), .Z(N62) );
  ANDN U7181 ( .B(out[608]), .A(rst), .Z(N620) );
  ANDN U7182 ( .B(out[609]), .A(rst), .Z(N621) );
  ANDN U7183 ( .B(out[610]), .A(rst), .Z(N622) );
  ANDN U7184 ( .B(out[611]), .A(rst), .Z(N623) );
  ANDN U7185 ( .B(out[612]), .A(rst), .Z(N624) );
  ANDN U7186 ( .B(out[613]), .A(rst), .Z(N625) );
  ANDN U7187 ( .B(out[614]), .A(rst), .Z(N626) );
  ANDN U7188 ( .B(out[615]), .A(rst), .Z(N627) );
  ANDN U7189 ( .B(out[616]), .A(rst), .Z(N628) );
  ANDN U7190 ( .B(out[617]), .A(rst), .Z(N629) );
  ANDN U7191 ( .B(out[51]), .A(rst), .Z(N63) );
  ANDN U7192 ( .B(out[618]), .A(rst), .Z(N630) );
  ANDN U7193 ( .B(out[619]), .A(rst), .Z(N631) );
  ANDN U7194 ( .B(out[620]), .A(rst), .Z(N632) );
  ANDN U7195 ( .B(out[621]), .A(rst), .Z(N633) );
  ANDN U7196 ( .B(out[622]), .A(rst), .Z(N634) );
  ANDN U7197 ( .B(out[623]), .A(rst), .Z(N635) );
  ANDN U7198 ( .B(out[624]), .A(rst), .Z(N636) );
  ANDN U7199 ( .B(out[625]), .A(rst), .Z(N637) );
  ANDN U7200 ( .B(out[626]), .A(rst), .Z(N638) );
  ANDN U7201 ( .B(out[627]), .A(rst), .Z(N639) );
  ANDN U7202 ( .B(out[52]), .A(rst), .Z(N64) );
  ANDN U7203 ( .B(out[628]), .A(rst), .Z(N640) );
  ANDN U7204 ( .B(out[629]), .A(rst), .Z(N641) );
  ANDN U7205 ( .B(out[630]), .A(rst), .Z(N642) );
  ANDN U7206 ( .B(out[631]), .A(rst), .Z(N643) );
  ANDN U7207 ( .B(out[632]), .A(rst), .Z(N644) );
  ANDN U7208 ( .B(out[633]), .A(rst), .Z(N645) );
  ANDN U7209 ( .B(out[634]), .A(rst), .Z(N646) );
  ANDN U7210 ( .B(out[635]), .A(rst), .Z(N647) );
  ANDN U7211 ( .B(out[636]), .A(rst), .Z(N648) );
  ANDN U7212 ( .B(out[637]), .A(rst), .Z(N649) );
  ANDN U7213 ( .B(out[53]), .A(rst), .Z(N65) );
  ANDN U7214 ( .B(out[638]), .A(rst), .Z(N650) );
  ANDN U7215 ( .B(out[639]), .A(rst), .Z(N651) );
  ANDN U7216 ( .B(out[640]), .A(rst), .Z(N652) );
  ANDN U7217 ( .B(out[641]), .A(rst), .Z(N653) );
  ANDN U7218 ( .B(out[642]), .A(rst), .Z(N654) );
  ANDN U7219 ( .B(out[643]), .A(rst), .Z(N655) );
  ANDN U7220 ( .B(out[644]), .A(rst), .Z(N656) );
  ANDN U7221 ( .B(out[645]), .A(rst), .Z(N657) );
  ANDN U7222 ( .B(out[646]), .A(rst), .Z(N658) );
  ANDN U7223 ( .B(out[647]), .A(rst), .Z(N659) );
  ANDN U7224 ( .B(out[54]), .A(rst), .Z(N66) );
  ANDN U7225 ( .B(out[648]), .A(rst), .Z(N660) );
  ANDN U7226 ( .B(out[649]), .A(rst), .Z(N661) );
  ANDN U7227 ( .B(out[650]), .A(rst), .Z(N662) );
  ANDN U7228 ( .B(out[651]), .A(rst), .Z(N663) );
  ANDN U7229 ( .B(out[652]), .A(rst), .Z(N664) );
  ANDN U7230 ( .B(out[653]), .A(rst), .Z(N665) );
  ANDN U7231 ( .B(out[654]), .A(rst), .Z(N666) );
  ANDN U7232 ( .B(out[655]), .A(rst), .Z(N667) );
  ANDN U7233 ( .B(out[656]), .A(rst), .Z(N668) );
  ANDN U7234 ( .B(out[657]), .A(rst), .Z(N669) );
  ANDN U7235 ( .B(out[55]), .A(rst), .Z(N67) );
  ANDN U7236 ( .B(out[658]), .A(rst), .Z(N670) );
  ANDN U7237 ( .B(out[659]), .A(rst), .Z(N671) );
  ANDN U7238 ( .B(out[660]), .A(rst), .Z(N672) );
  ANDN U7239 ( .B(out[661]), .A(rst), .Z(N673) );
  ANDN U7240 ( .B(out[662]), .A(rst), .Z(N674) );
  ANDN U7241 ( .B(out[663]), .A(rst), .Z(N675) );
  ANDN U7242 ( .B(out[664]), .A(rst), .Z(N676) );
  ANDN U7243 ( .B(out[665]), .A(rst), .Z(N677) );
  ANDN U7244 ( .B(out[666]), .A(rst), .Z(N678) );
  ANDN U7245 ( .B(out[667]), .A(rst), .Z(N679) );
  ANDN U7246 ( .B(out[56]), .A(rst), .Z(N68) );
  ANDN U7247 ( .B(out[668]), .A(rst), .Z(N680) );
  ANDN U7248 ( .B(out[669]), .A(rst), .Z(N681) );
  ANDN U7249 ( .B(out[670]), .A(rst), .Z(N682) );
  ANDN U7250 ( .B(out[671]), .A(rst), .Z(N683) );
  ANDN U7251 ( .B(out[672]), .A(rst), .Z(N684) );
  ANDN U7252 ( .B(out[673]), .A(rst), .Z(N685) );
  ANDN U7253 ( .B(out[674]), .A(rst), .Z(N686) );
  ANDN U7254 ( .B(out[675]), .A(rst), .Z(N687) );
  ANDN U7255 ( .B(out[676]), .A(rst), .Z(N688) );
  ANDN U7256 ( .B(out[677]), .A(rst), .Z(N689) );
  ANDN U7257 ( .B(out[57]), .A(rst), .Z(N69) );
  ANDN U7258 ( .B(out[678]), .A(rst), .Z(N690) );
  ANDN U7259 ( .B(out[679]), .A(rst), .Z(N691) );
  ANDN U7260 ( .B(out[680]), .A(rst), .Z(N692) );
  ANDN U7261 ( .B(out[681]), .A(rst), .Z(N693) );
  ANDN U7262 ( .B(out[682]), .A(rst), .Z(N694) );
  ANDN U7263 ( .B(out[683]), .A(rst), .Z(N695) );
  ANDN U7264 ( .B(out[684]), .A(rst), .Z(N696) );
  ANDN U7265 ( .B(out[685]), .A(rst), .Z(N697) );
  ANDN U7266 ( .B(out[686]), .A(rst), .Z(N698) );
  ANDN U7267 ( .B(out[687]), .A(rst), .Z(N699) );
  ANDN U7268 ( .B(rc_i[0]), .A(rst), .Z(N7) );
  ANDN U7269 ( .B(out[58]), .A(rst), .Z(N70) );
  ANDN U7270 ( .B(out[688]), .A(rst), .Z(N700) );
  ANDN U7271 ( .B(out[689]), .A(rst), .Z(N701) );
  ANDN U7272 ( .B(out[690]), .A(rst), .Z(N702) );
  ANDN U7273 ( .B(out[691]), .A(rst), .Z(N703) );
  ANDN U7274 ( .B(out[692]), .A(rst), .Z(N704) );
  ANDN U7275 ( .B(out[693]), .A(rst), .Z(N705) );
  ANDN U7276 ( .B(out[694]), .A(rst), .Z(N706) );
  ANDN U7277 ( .B(out[695]), .A(rst), .Z(N707) );
  ANDN U7278 ( .B(out[696]), .A(rst), .Z(N708) );
  ANDN U7279 ( .B(out[697]), .A(rst), .Z(N709) );
  ANDN U7280 ( .B(out[59]), .A(rst), .Z(N71) );
  ANDN U7281 ( .B(out[698]), .A(rst), .Z(N710) );
  ANDN U7282 ( .B(out[699]), .A(rst), .Z(N711) );
  ANDN U7283 ( .B(out[700]), .A(rst), .Z(N712) );
  ANDN U7284 ( .B(out[701]), .A(rst), .Z(N713) );
  ANDN U7285 ( .B(out[702]), .A(rst), .Z(N714) );
  ANDN U7286 ( .B(out[703]), .A(rst), .Z(N715) );
  ANDN U7287 ( .B(out[704]), .A(rst), .Z(N716) );
  ANDN U7288 ( .B(out[705]), .A(rst), .Z(N717) );
  ANDN U7289 ( .B(out[706]), .A(rst), .Z(N718) );
  ANDN U7290 ( .B(out[707]), .A(rst), .Z(N719) );
  ANDN U7291 ( .B(out[60]), .A(rst), .Z(N72) );
  ANDN U7292 ( .B(out[708]), .A(rst), .Z(N720) );
  ANDN U7293 ( .B(out[709]), .A(rst), .Z(N721) );
  ANDN U7294 ( .B(out[710]), .A(rst), .Z(N722) );
  ANDN U7295 ( .B(out[711]), .A(rst), .Z(N723) );
  ANDN U7296 ( .B(out[712]), .A(rst), .Z(N724) );
  ANDN U7297 ( .B(out[713]), .A(rst), .Z(N725) );
  ANDN U7298 ( .B(out[714]), .A(rst), .Z(N726) );
  ANDN U7299 ( .B(out[715]), .A(rst), .Z(N727) );
  ANDN U7300 ( .B(out[716]), .A(rst), .Z(N728) );
  ANDN U7301 ( .B(out[717]), .A(rst), .Z(N729) );
  ANDN U7302 ( .B(out[61]), .A(rst), .Z(N73) );
  ANDN U7303 ( .B(out[718]), .A(rst), .Z(N730) );
  ANDN U7304 ( .B(out[719]), .A(rst), .Z(N731) );
  ANDN U7305 ( .B(out[720]), .A(rst), .Z(N732) );
  ANDN U7306 ( .B(out[721]), .A(rst), .Z(N733) );
  ANDN U7307 ( .B(out[722]), .A(rst), .Z(N734) );
  ANDN U7308 ( .B(out[723]), .A(rst), .Z(N735) );
  ANDN U7309 ( .B(out[724]), .A(rst), .Z(N736) );
  ANDN U7310 ( .B(out[725]), .A(rst), .Z(N737) );
  ANDN U7311 ( .B(out[726]), .A(rst), .Z(N738) );
  ANDN U7312 ( .B(out[727]), .A(rst), .Z(N739) );
  ANDN U7313 ( .B(out[62]), .A(rst), .Z(N74) );
  ANDN U7314 ( .B(out[728]), .A(rst), .Z(N740) );
  ANDN U7315 ( .B(out[729]), .A(rst), .Z(N741) );
  ANDN U7316 ( .B(out[730]), .A(rst), .Z(N742) );
  ANDN U7317 ( .B(out[731]), .A(rst), .Z(N743) );
  ANDN U7318 ( .B(out[732]), .A(rst), .Z(N744) );
  ANDN U7319 ( .B(out[733]), .A(rst), .Z(N745) );
  ANDN U7320 ( .B(out[734]), .A(rst), .Z(N746) );
  ANDN U7321 ( .B(out[735]), .A(rst), .Z(N747) );
  ANDN U7322 ( .B(out[736]), .A(rst), .Z(N748) );
  ANDN U7323 ( .B(out[737]), .A(rst), .Z(N749) );
  ANDN U7324 ( .B(out[63]), .A(rst), .Z(N75) );
  ANDN U7325 ( .B(out[738]), .A(rst), .Z(N750) );
  ANDN U7326 ( .B(out[739]), .A(rst), .Z(N751) );
  ANDN U7327 ( .B(out[740]), .A(rst), .Z(N752) );
  ANDN U7328 ( .B(out[741]), .A(rst), .Z(N753) );
  ANDN U7329 ( .B(out[742]), .A(rst), .Z(N754) );
  ANDN U7330 ( .B(out[743]), .A(rst), .Z(N755) );
  ANDN U7331 ( .B(out[744]), .A(rst), .Z(N756) );
  ANDN U7332 ( .B(out[745]), .A(rst), .Z(N757) );
  ANDN U7333 ( .B(out[746]), .A(rst), .Z(N758) );
  ANDN U7334 ( .B(out[747]), .A(rst), .Z(N759) );
  ANDN U7335 ( .B(out[64]), .A(rst), .Z(N76) );
  ANDN U7336 ( .B(out[748]), .A(rst), .Z(N760) );
  ANDN U7337 ( .B(out[749]), .A(rst), .Z(N761) );
  ANDN U7338 ( .B(out[750]), .A(rst), .Z(N762) );
  ANDN U7339 ( .B(out[751]), .A(rst), .Z(N763) );
  ANDN U7340 ( .B(out[752]), .A(rst), .Z(N764) );
  ANDN U7341 ( .B(out[753]), .A(rst), .Z(N765) );
  ANDN U7342 ( .B(out[754]), .A(rst), .Z(N766) );
  ANDN U7343 ( .B(out[755]), .A(rst), .Z(N767) );
  ANDN U7344 ( .B(out[756]), .A(rst), .Z(N768) );
  ANDN U7345 ( .B(out[757]), .A(rst), .Z(N769) );
  ANDN U7346 ( .B(out[65]), .A(rst), .Z(N77) );
  ANDN U7347 ( .B(out[758]), .A(rst), .Z(N770) );
  ANDN U7348 ( .B(out[759]), .A(rst), .Z(N771) );
  ANDN U7349 ( .B(out[760]), .A(rst), .Z(N772) );
  ANDN U7350 ( .B(out[761]), .A(rst), .Z(N773) );
  ANDN U7351 ( .B(out[762]), .A(rst), .Z(N774) );
  ANDN U7352 ( .B(out[763]), .A(rst), .Z(N775) );
  ANDN U7353 ( .B(out[764]), .A(rst), .Z(N776) );
  ANDN U7354 ( .B(out[765]), .A(rst), .Z(N777) );
  ANDN U7355 ( .B(out[766]), .A(rst), .Z(N778) );
  ANDN U7356 ( .B(out[767]), .A(rst), .Z(N779) );
  ANDN U7357 ( .B(out[66]), .A(rst), .Z(N78) );
  ANDN U7358 ( .B(out[768]), .A(rst), .Z(N780) );
  ANDN U7359 ( .B(out[769]), .A(rst), .Z(N781) );
  ANDN U7360 ( .B(out[770]), .A(rst), .Z(N782) );
  ANDN U7361 ( .B(out[771]), .A(rst), .Z(N783) );
  ANDN U7362 ( .B(out[772]), .A(rst), .Z(N784) );
  ANDN U7363 ( .B(out[773]), .A(rst), .Z(N785) );
  ANDN U7364 ( .B(out[774]), .A(rst), .Z(N786) );
  ANDN U7365 ( .B(out[775]), .A(rst), .Z(N787) );
  ANDN U7366 ( .B(out[776]), .A(rst), .Z(N788) );
  ANDN U7367 ( .B(out[777]), .A(rst), .Z(N789) );
  ANDN U7368 ( .B(out[67]), .A(rst), .Z(N79) );
  ANDN U7369 ( .B(out[778]), .A(rst), .Z(N790) );
  ANDN U7370 ( .B(out[779]), .A(rst), .Z(N791) );
  ANDN U7371 ( .B(out[780]), .A(rst), .Z(N792) );
  ANDN U7372 ( .B(out[781]), .A(rst), .Z(N793) );
  ANDN U7373 ( .B(out[782]), .A(rst), .Z(N794) );
  ANDN U7374 ( .B(out[783]), .A(rst), .Z(N795) );
  ANDN U7375 ( .B(out[784]), .A(rst), .Z(N796) );
  ANDN U7376 ( .B(out[785]), .A(rst), .Z(N797) );
  ANDN U7377 ( .B(out[786]), .A(rst), .Z(N798) );
  ANDN U7378 ( .B(out[787]), .A(rst), .Z(N799) );
  ANDN U7379 ( .B(rc_i[1]), .A(rst), .Z(N8) );
  ANDN U7380 ( .B(out[68]), .A(rst), .Z(N80) );
  ANDN U7381 ( .B(out[788]), .A(rst), .Z(N800) );
  ANDN U7382 ( .B(out[789]), .A(rst), .Z(N801) );
  ANDN U7383 ( .B(out[790]), .A(rst), .Z(N802) );
  ANDN U7384 ( .B(out[791]), .A(rst), .Z(N803) );
  ANDN U7385 ( .B(out[792]), .A(rst), .Z(N804) );
  ANDN U7386 ( .B(out[793]), .A(rst), .Z(N805) );
  ANDN U7387 ( .B(out[794]), .A(rst), .Z(N806) );
  ANDN U7388 ( .B(out[795]), .A(rst), .Z(N807) );
  ANDN U7389 ( .B(out[796]), .A(rst), .Z(N808) );
  ANDN U7390 ( .B(out[797]), .A(rst), .Z(N809) );
  ANDN U7391 ( .B(out[69]), .A(rst), .Z(N81) );
  ANDN U7392 ( .B(out[798]), .A(rst), .Z(N810) );
  ANDN U7393 ( .B(out[799]), .A(rst), .Z(N811) );
  ANDN U7394 ( .B(out[800]), .A(rst), .Z(N812) );
  ANDN U7395 ( .B(out[801]), .A(rst), .Z(N813) );
  ANDN U7396 ( .B(out[802]), .A(rst), .Z(N814) );
  ANDN U7397 ( .B(out[803]), .A(rst), .Z(N815) );
  ANDN U7398 ( .B(out[804]), .A(rst), .Z(N816) );
  ANDN U7399 ( .B(out[805]), .A(rst), .Z(N817) );
  ANDN U7400 ( .B(out[806]), .A(rst), .Z(N818) );
  ANDN U7401 ( .B(out[807]), .A(rst), .Z(N819) );
  ANDN U7402 ( .B(out[70]), .A(rst), .Z(N82) );
  ANDN U7403 ( .B(out[808]), .A(rst), .Z(N820) );
  ANDN U7404 ( .B(out[809]), .A(rst), .Z(N821) );
  ANDN U7405 ( .B(out[810]), .A(rst), .Z(N822) );
  ANDN U7406 ( .B(out[811]), .A(rst), .Z(N823) );
  ANDN U7407 ( .B(out[812]), .A(rst), .Z(N824) );
  ANDN U7408 ( .B(out[813]), .A(rst), .Z(N825) );
  ANDN U7409 ( .B(out[814]), .A(rst), .Z(N826) );
  ANDN U7410 ( .B(out[815]), .A(rst), .Z(N827) );
  ANDN U7411 ( .B(out[816]), .A(rst), .Z(N828) );
  ANDN U7412 ( .B(out[817]), .A(rst), .Z(N829) );
  ANDN U7413 ( .B(out[71]), .A(rst), .Z(N83) );
  ANDN U7414 ( .B(out[818]), .A(rst), .Z(N830) );
  ANDN U7415 ( .B(out[819]), .A(rst), .Z(N831) );
  ANDN U7416 ( .B(out[820]), .A(rst), .Z(N832) );
  ANDN U7417 ( .B(out[821]), .A(rst), .Z(N833) );
  ANDN U7418 ( .B(out[822]), .A(rst), .Z(N834) );
  ANDN U7419 ( .B(out[823]), .A(rst), .Z(N835) );
  ANDN U7420 ( .B(out[824]), .A(rst), .Z(N836) );
  ANDN U7421 ( .B(out[825]), .A(rst), .Z(N837) );
  ANDN U7422 ( .B(out[826]), .A(rst), .Z(N838) );
  ANDN U7423 ( .B(out[827]), .A(rst), .Z(N839) );
  ANDN U7424 ( .B(out[72]), .A(rst), .Z(N84) );
  ANDN U7425 ( .B(out[828]), .A(rst), .Z(N840) );
  ANDN U7426 ( .B(out[829]), .A(rst), .Z(N841) );
  ANDN U7427 ( .B(out[830]), .A(rst), .Z(N842) );
  ANDN U7428 ( .B(out[831]), .A(rst), .Z(N843) );
  ANDN U7429 ( .B(out[832]), .A(rst), .Z(N844) );
  ANDN U7430 ( .B(out[833]), .A(rst), .Z(N845) );
  ANDN U7431 ( .B(out[834]), .A(rst), .Z(N846) );
  ANDN U7432 ( .B(out[835]), .A(rst), .Z(N847) );
  ANDN U7433 ( .B(out[836]), .A(rst), .Z(N848) );
  ANDN U7434 ( .B(out[837]), .A(rst), .Z(N849) );
  ANDN U7435 ( .B(out[73]), .A(rst), .Z(N85) );
  ANDN U7436 ( .B(out[838]), .A(rst), .Z(N850) );
  ANDN U7437 ( .B(out[839]), .A(rst), .Z(N851) );
  ANDN U7438 ( .B(out[840]), .A(rst), .Z(N852) );
  ANDN U7439 ( .B(out[841]), .A(rst), .Z(N853) );
  ANDN U7440 ( .B(out[842]), .A(rst), .Z(N854) );
  ANDN U7441 ( .B(out[843]), .A(rst), .Z(N855) );
  ANDN U7442 ( .B(out[844]), .A(rst), .Z(N856) );
  ANDN U7443 ( .B(out[845]), .A(rst), .Z(N857) );
  ANDN U7444 ( .B(out[846]), .A(rst), .Z(N858) );
  ANDN U7445 ( .B(out[847]), .A(rst), .Z(N859) );
  ANDN U7446 ( .B(out[74]), .A(rst), .Z(N86) );
  ANDN U7447 ( .B(out[848]), .A(rst), .Z(N860) );
  ANDN U7448 ( .B(out[849]), .A(rst), .Z(N861) );
  ANDN U7449 ( .B(out[850]), .A(rst), .Z(N862) );
  ANDN U7450 ( .B(out[851]), .A(rst), .Z(N863) );
  ANDN U7451 ( .B(out[852]), .A(rst), .Z(N864) );
  ANDN U7452 ( .B(out[853]), .A(rst), .Z(N865) );
  ANDN U7453 ( .B(out[854]), .A(rst), .Z(N866) );
  ANDN U7454 ( .B(out[855]), .A(rst), .Z(N867) );
  ANDN U7455 ( .B(out[856]), .A(rst), .Z(N868) );
  ANDN U7456 ( .B(out[857]), .A(rst), .Z(N869) );
  ANDN U7457 ( .B(out[75]), .A(rst), .Z(N87) );
  ANDN U7458 ( .B(out[858]), .A(rst), .Z(N870) );
  ANDN U7459 ( .B(out[859]), .A(rst), .Z(N871) );
  ANDN U7460 ( .B(out[860]), .A(rst), .Z(N872) );
  ANDN U7461 ( .B(out[861]), .A(rst), .Z(N873) );
  ANDN U7462 ( .B(out[862]), .A(rst), .Z(N874) );
  ANDN U7463 ( .B(out[863]), .A(rst), .Z(N875) );
  ANDN U7464 ( .B(out[864]), .A(rst), .Z(N876) );
  ANDN U7465 ( .B(out[865]), .A(rst), .Z(N877) );
  ANDN U7466 ( .B(out[866]), .A(rst), .Z(N878) );
  ANDN U7467 ( .B(out[867]), .A(rst), .Z(N879) );
  ANDN U7468 ( .B(out[76]), .A(rst), .Z(N88) );
  ANDN U7469 ( .B(out[868]), .A(rst), .Z(N880) );
  ANDN U7470 ( .B(out[869]), .A(rst), .Z(N881) );
  ANDN U7471 ( .B(out[870]), .A(rst), .Z(N882) );
  ANDN U7472 ( .B(out[871]), .A(rst), .Z(N883) );
  ANDN U7473 ( .B(out[872]), .A(rst), .Z(N884) );
  ANDN U7474 ( .B(out[873]), .A(rst), .Z(N885) );
  ANDN U7475 ( .B(out[874]), .A(rst), .Z(N886) );
  ANDN U7476 ( .B(out[875]), .A(rst), .Z(N887) );
  ANDN U7477 ( .B(out[876]), .A(rst), .Z(N888) );
  ANDN U7478 ( .B(out[877]), .A(rst), .Z(N889) );
  ANDN U7479 ( .B(out[77]), .A(rst), .Z(N89) );
  ANDN U7480 ( .B(out[878]), .A(rst), .Z(N890) );
  ANDN U7481 ( .B(out[879]), .A(rst), .Z(N891) );
  ANDN U7482 ( .B(out[880]), .A(rst), .Z(N892) );
  ANDN U7483 ( .B(out[881]), .A(rst), .Z(N893) );
  ANDN U7484 ( .B(out[882]), .A(rst), .Z(N894) );
  ANDN U7485 ( .B(out[883]), .A(rst), .Z(N895) );
  ANDN U7486 ( .B(out[884]), .A(rst), .Z(N896) );
  ANDN U7487 ( .B(out[885]), .A(rst), .Z(N897) );
  ANDN U7488 ( .B(out[886]), .A(rst), .Z(N898) );
  ANDN U7489 ( .B(out[887]), .A(rst), .Z(N899) );
  ANDN U7490 ( .B(rc_i[2]), .A(rst), .Z(N9) );
  ANDN U7491 ( .B(out[78]), .A(rst), .Z(N90) );
  ANDN U7492 ( .B(out[888]), .A(rst), .Z(N900) );
  ANDN U7493 ( .B(out[889]), .A(rst), .Z(N901) );
  ANDN U7494 ( .B(out[890]), .A(rst), .Z(N902) );
  ANDN U7495 ( .B(out[891]), .A(rst), .Z(N903) );
  ANDN U7496 ( .B(out[892]), .A(rst), .Z(N904) );
  ANDN U7497 ( .B(out[893]), .A(rst), .Z(N905) );
  ANDN U7498 ( .B(out[894]), .A(rst), .Z(N906) );
  ANDN U7499 ( .B(out[895]), .A(rst), .Z(N907) );
  ANDN U7500 ( .B(out[896]), .A(rst), .Z(N908) );
  ANDN U7501 ( .B(out[897]), .A(rst), .Z(N909) );
  ANDN U7502 ( .B(out[79]), .A(rst), .Z(N91) );
  ANDN U7503 ( .B(out[898]), .A(rst), .Z(N910) );
  ANDN U7504 ( .B(out[899]), .A(rst), .Z(N911) );
  ANDN U7505 ( .B(out[900]), .A(rst), .Z(N912) );
  ANDN U7506 ( .B(out[901]), .A(rst), .Z(N913) );
  ANDN U7507 ( .B(out[902]), .A(rst), .Z(N914) );
  ANDN U7508 ( .B(out[903]), .A(rst), .Z(N915) );
  ANDN U7509 ( .B(out[904]), .A(rst), .Z(N916) );
  ANDN U7510 ( .B(out[905]), .A(rst), .Z(N917) );
  ANDN U7511 ( .B(out[906]), .A(rst), .Z(N918) );
  ANDN U7512 ( .B(out[907]), .A(rst), .Z(N919) );
  ANDN U7513 ( .B(out[80]), .A(rst), .Z(N92) );
  ANDN U7514 ( .B(out[908]), .A(rst), .Z(N920) );
  ANDN U7515 ( .B(out[909]), .A(rst), .Z(N921) );
  ANDN U7516 ( .B(out[910]), .A(rst), .Z(N922) );
  ANDN U7517 ( .B(out[911]), .A(rst), .Z(N923) );
  ANDN U7518 ( .B(out[912]), .A(rst), .Z(N924) );
  ANDN U7519 ( .B(out[913]), .A(rst), .Z(N925) );
  ANDN U7520 ( .B(out[914]), .A(rst), .Z(N926) );
  ANDN U7521 ( .B(out[915]), .A(rst), .Z(N927) );
  ANDN U7522 ( .B(out[916]), .A(rst), .Z(N928) );
  ANDN U7523 ( .B(out[917]), .A(rst), .Z(N929) );
  ANDN U7524 ( .B(out[81]), .A(rst), .Z(N93) );
  ANDN U7525 ( .B(out[918]), .A(rst), .Z(N930) );
  ANDN U7526 ( .B(out[919]), .A(rst), .Z(N931) );
  ANDN U7527 ( .B(out[920]), .A(rst), .Z(N932) );
  ANDN U7528 ( .B(out[921]), .A(rst), .Z(N933) );
  ANDN U7529 ( .B(out[922]), .A(rst), .Z(N934) );
  ANDN U7530 ( .B(out[923]), .A(rst), .Z(N935) );
  ANDN U7531 ( .B(out[924]), .A(rst), .Z(N936) );
  ANDN U7532 ( .B(out[925]), .A(rst), .Z(N937) );
  ANDN U7533 ( .B(out[926]), .A(rst), .Z(N938) );
  ANDN U7534 ( .B(out[927]), .A(rst), .Z(N939) );
  ANDN U7535 ( .B(out[82]), .A(rst), .Z(N94) );
  ANDN U7536 ( .B(out[928]), .A(rst), .Z(N940) );
  ANDN U7537 ( .B(out[929]), .A(rst), .Z(N941) );
  ANDN U7538 ( .B(out[930]), .A(rst), .Z(N942) );
  ANDN U7539 ( .B(out[931]), .A(rst), .Z(N943) );
  ANDN U7540 ( .B(out[932]), .A(rst), .Z(N944) );
  ANDN U7541 ( .B(out[933]), .A(rst), .Z(N945) );
  ANDN U7542 ( .B(out[934]), .A(rst), .Z(N946) );
  ANDN U7543 ( .B(out[935]), .A(rst), .Z(N947) );
  ANDN U7544 ( .B(out[936]), .A(rst), .Z(N948) );
  ANDN U7545 ( .B(out[937]), .A(rst), .Z(N949) );
  ANDN U7546 ( .B(out[83]), .A(rst), .Z(N95) );
  ANDN U7547 ( .B(out[938]), .A(rst), .Z(N950) );
  ANDN U7548 ( .B(out[939]), .A(rst), .Z(N951) );
  ANDN U7549 ( .B(out[940]), .A(rst), .Z(N952) );
  ANDN U7550 ( .B(out[941]), .A(rst), .Z(N953) );
  ANDN U7551 ( .B(out[942]), .A(rst), .Z(N954) );
  ANDN U7552 ( .B(out[943]), .A(rst), .Z(N955) );
  ANDN U7553 ( .B(out[944]), .A(rst), .Z(N956) );
  ANDN U7554 ( .B(out[945]), .A(rst), .Z(N957) );
  ANDN U7555 ( .B(out[946]), .A(rst), .Z(N958) );
  ANDN U7556 ( .B(out[947]), .A(rst), .Z(N959) );
  ANDN U7557 ( .B(out[84]), .A(rst), .Z(N96) );
  ANDN U7558 ( .B(out[948]), .A(rst), .Z(N960) );
  ANDN U7559 ( .B(out[949]), .A(rst), .Z(N961) );
  ANDN U7560 ( .B(out[950]), .A(rst), .Z(N962) );
  ANDN U7561 ( .B(out[951]), .A(rst), .Z(N963) );
  ANDN U7562 ( .B(out[952]), .A(rst), .Z(N964) );
  ANDN U7563 ( .B(out[953]), .A(rst), .Z(N965) );
  ANDN U7564 ( .B(out[954]), .A(rst), .Z(N966) );
  ANDN U7565 ( .B(out[955]), .A(rst), .Z(N967) );
  ANDN U7566 ( .B(out[956]), .A(rst), .Z(N968) );
  ANDN U7567 ( .B(out[957]), .A(rst), .Z(N969) );
  ANDN U7568 ( .B(out[85]), .A(rst), .Z(N97) );
  ANDN U7569 ( .B(out[958]), .A(rst), .Z(N970) );
  ANDN U7570 ( .B(out[959]), .A(rst), .Z(N971) );
  ANDN U7571 ( .B(out[960]), .A(rst), .Z(N972) );
  ANDN U7572 ( .B(out[961]), .A(rst), .Z(N973) );
  ANDN U7573 ( .B(out[962]), .A(rst), .Z(N974) );
  ANDN U7574 ( .B(out[963]), .A(rst), .Z(N975) );
  ANDN U7575 ( .B(out[964]), .A(rst), .Z(N976) );
  ANDN U7576 ( .B(out[965]), .A(rst), .Z(N977) );
  ANDN U7577 ( .B(out[966]), .A(rst), .Z(N978) );
  ANDN U7578 ( .B(out[967]), .A(rst), .Z(N979) );
  ANDN U7579 ( .B(out[86]), .A(rst), .Z(N98) );
  ANDN U7580 ( .B(out[968]), .A(rst), .Z(N980) );
  ANDN U7581 ( .B(out[969]), .A(rst), .Z(N981) );
  ANDN U7582 ( .B(out[970]), .A(rst), .Z(N982) );
  ANDN U7583 ( .B(out[971]), .A(rst), .Z(N983) );
  ANDN U7584 ( .B(out[972]), .A(rst), .Z(N984) );
  ANDN U7585 ( .B(out[973]), .A(rst), .Z(N985) );
  ANDN U7586 ( .B(out[974]), .A(rst), .Z(N986) );
  ANDN U7587 ( .B(out[975]), .A(rst), .Z(N987) );
  ANDN U7588 ( .B(out[976]), .A(rst), .Z(N988) );
  ANDN U7589 ( .B(out[977]), .A(rst), .Z(N989) );
  ANDN U7590 ( .B(out[87]), .A(rst), .Z(N99) );
  ANDN U7591 ( .B(out[978]), .A(rst), .Z(N990) );
  ANDN U7592 ( .B(out[979]), .A(rst), .Z(N991) );
  ANDN U7593 ( .B(out[980]), .A(rst), .Z(N992) );
  ANDN U7594 ( .B(out[981]), .A(rst), .Z(N993) );
  ANDN U7595 ( .B(out[982]), .A(rst), .Z(N994) );
  ANDN U7596 ( .B(out[983]), .A(rst), .Z(N995) );
  ANDN U7597 ( .B(out[984]), .A(rst), .Z(N996) );
  ANDN U7598 ( .B(out[985]), .A(rst), .Z(N997) );
  ANDN U7599 ( .B(out[986]), .A(rst), .Z(N998) );
  ANDN U7600 ( .B(out[987]), .A(rst), .Z(N999) );
  OR U7601 ( .A(rc_i[1]), .B(rc_i[3]), .Z(\RCONST[3].rconst_/N10 ) );
  OR U7602 ( .A(rc_i[0]), .B(\RCONST[3].rconst_/N10 ), .Z(
        \RCONST[2].rconst_/N62 ) );
  OR U7603 ( .A(rc_i[5]), .B(\RCONST[2].rconst_/N62 ), .Z(\rc[3][15] ) );
  OR U7604 ( .A(rc_i[3]), .B(rc_i[2]), .Z(\RCONST[1].rconst_/N26 ) );
  OR U7605 ( .A(rc_i[4]), .B(\RCONST[1].rconst_/N26 ), .Z(\rc[3][1] ) );
  OR U7606 ( .A(rc_i[2]), .B(\RCONST[3].rconst_/N10 ), .Z(
        \RCONST[0].rconst_/N25 ) );
  OR U7607 ( .A(rc_i[4]), .B(\RCONST[0].rconst_/N25 ), .Z(
        \RCONST[0].rconst_/N17 ) );
  NOR U7608 ( .A(rc_i[5]), .B(rc_i[2]), .Z(n2764) );
  NANDN U7609 ( .A(rc_i[1]), .B(n2764), .Z(\RCONST[2].rconst_/N57 ) );
  NANDN U7610 ( .A(\RCONST[3].rconst_/N10 ), .B(n2764), .Z(\rc[2][0] ) );
  OR U7611 ( .A(rc_i[5]), .B(rc_i[4]), .Z(\RCONST[0].rconst_/N67 ) );
  OR U7612 ( .A(rc_i[5]), .B(rc_i[3]), .Z(\RCONST[0].rconst_/N56 ) );
  OR U7613 ( .A(rc_i[4]), .B(\RCONST[0].rconst_/N56 ), .Z(
        \RCONST[1].rconst_/N68 ) );
  OR U7614 ( .A(\RCONST[3].rconst_/N10 ), .B(\RCONST[0].rconst_/N67 ), .Z(
        \RCONST[0].rconst_/N48 ) );
  OR U7615 ( .A(rc_i[0]), .B(rc_i[3]), .Z(\RCONST[1].rconst_/N15 ) );
  OR U7616 ( .A(rc_i[5]), .B(rc_i[0]), .Z(\RCONST[1].rconst_/N49 ) );
  OR U7617 ( .A(rc_i[0]), .B(rc_i[4]), .Z(\RCONST[2].rconst_/N18 ) );
  OR U7618 ( .A(\RCONST[2].rconst_/N18 ), .B(\RCONST[1].rconst_/N26 ), .Z(
        \RCONST[2].rconst_/N28 ) );
  OR U7619 ( .A(\RCONST[0].rconst_/N25 ), .B(\RCONST[2].rconst_/N18 ), .Z(
        \RCONST[2].rconst_/N47 ) );
  NANDN U7620 ( .A(\RCONST[2].rconst_/N18 ), .B(n2764), .Z(\rc[3][31] ) );
  OR U7621 ( .A(\RCONST[1].rconst_/N49 ), .B(\rc[3][1] ), .Z(\rc[1][7] ) );
  OR U7622 ( .A(rc_i[4]), .B(\RCONST[2].rconst_/N57 ), .Z(\rc[3][3] ) );
  OR U7623 ( .A(\RCONST[2].rconst_/N62 ), .B(\RCONST[0].rconst_/N67 ), .Z(
        \rc[3][63] ) );
  NAND U7624 ( .A(init), .B(round_reg[0]), .Z(n2766) );
  NANDN U7625 ( .A(init), .B(in[0]), .Z(n2765) );
  NAND U7626 ( .A(n2766), .B(n2765), .Z(\round_in[0][0] ) );
  AND U7627 ( .A(round_reg[1000]), .B(init), .Z(\round_in[0][1000] ) );
  AND U7628 ( .A(round_reg[1001]), .B(init), .Z(\round_in[0][1001] ) );
  AND U7629 ( .A(round_reg[1002]), .B(init), .Z(\round_in[0][1002] ) );
  AND U7630 ( .A(round_reg[1003]), .B(init), .Z(\round_in[0][1003] ) );
  AND U7631 ( .A(round_reg[1004]), .B(init), .Z(\round_in[0][1004] ) );
  AND U7632 ( .A(round_reg[1005]), .B(init), .Z(\round_in[0][1005] ) );
  AND U7633 ( .A(round_reg[1006]), .B(init), .Z(\round_in[0][1006] ) );
  AND U7634 ( .A(round_reg[1007]), .B(init), .Z(\round_in[0][1007] ) );
  AND U7635 ( .A(round_reg[1008]), .B(init), .Z(\round_in[0][1008] ) );
  AND U7636 ( .A(round_reg[1009]), .B(init), .Z(\round_in[0][1009] ) );
  NAND U7637 ( .A(init), .B(round_reg[100]), .Z(n2768) );
  NANDN U7638 ( .A(init), .B(in[100]), .Z(n2767) );
  NAND U7639 ( .A(n2768), .B(n2767), .Z(\round_in[0][100] ) );
  AND U7640 ( .A(round_reg[1010]), .B(init), .Z(\round_in[0][1010] ) );
  AND U7641 ( .A(round_reg[1011]), .B(init), .Z(\round_in[0][1011] ) );
  AND U7642 ( .A(round_reg[1012]), .B(init), .Z(\round_in[0][1012] ) );
  AND U7643 ( .A(round_reg[1013]), .B(init), .Z(\round_in[0][1013] ) );
  AND U7644 ( .A(round_reg[1014]), .B(init), .Z(\round_in[0][1014] ) );
  AND U7645 ( .A(round_reg[1015]), .B(init), .Z(\round_in[0][1015] ) );
  AND U7646 ( .A(round_reg[1016]), .B(init), .Z(\round_in[0][1016] ) );
  AND U7647 ( .A(round_reg[1017]), .B(init), .Z(\round_in[0][1017] ) );
  AND U7648 ( .A(round_reg[1018]), .B(init), .Z(\round_in[0][1018] ) );
  AND U7649 ( .A(round_reg[1019]), .B(init), .Z(\round_in[0][1019] ) );
  NAND U7650 ( .A(init), .B(round_reg[101]), .Z(n2770) );
  NANDN U7651 ( .A(init), .B(in[101]), .Z(n2769) );
  NAND U7652 ( .A(n2770), .B(n2769), .Z(\round_in[0][101] ) );
  AND U7653 ( .A(round_reg[1020]), .B(init), .Z(\round_in[0][1020] ) );
  AND U7654 ( .A(round_reg[1021]), .B(init), .Z(\round_in[0][1021] ) );
  AND U7655 ( .A(round_reg[1022]), .B(init), .Z(\round_in[0][1022] ) );
  AND U7656 ( .A(round_reg[1023]), .B(init), .Z(\round_in[0][1023] ) );
  AND U7657 ( .A(round_reg[1024]), .B(init), .Z(\round_in[0][1024] ) );
  AND U7658 ( .A(round_reg[1025]), .B(init), .Z(\round_in[0][1025] ) );
  AND U7659 ( .A(round_reg[1026]), .B(init), .Z(\round_in[0][1026] ) );
  AND U7660 ( .A(round_reg[1027]), .B(init), .Z(\round_in[0][1027] ) );
  AND U7661 ( .A(round_reg[1028]), .B(init), .Z(\round_in[0][1028] ) );
  AND U7662 ( .A(round_reg[1029]), .B(init), .Z(\round_in[0][1029] ) );
  NAND U7663 ( .A(init), .B(round_reg[102]), .Z(n2772) );
  NANDN U7664 ( .A(init), .B(in[102]), .Z(n2771) );
  NAND U7665 ( .A(n2772), .B(n2771), .Z(\round_in[0][102] ) );
  AND U7666 ( .A(round_reg[1030]), .B(init), .Z(\round_in[0][1030] ) );
  AND U7667 ( .A(round_reg[1031]), .B(init), .Z(\round_in[0][1031] ) );
  AND U7668 ( .A(round_reg[1032]), .B(init), .Z(\round_in[0][1032] ) );
  AND U7669 ( .A(round_reg[1033]), .B(init), .Z(\round_in[0][1033] ) );
  AND U7670 ( .A(round_reg[1034]), .B(init), .Z(\round_in[0][1034] ) );
  AND U7671 ( .A(round_reg[1035]), .B(init), .Z(\round_in[0][1035] ) );
  AND U7672 ( .A(round_reg[1036]), .B(init), .Z(\round_in[0][1036] ) );
  AND U7673 ( .A(round_reg[1037]), .B(init), .Z(\round_in[0][1037] ) );
  AND U7674 ( .A(round_reg[1038]), .B(init), .Z(\round_in[0][1038] ) );
  AND U7675 ( .A(round_reg[1039]), .B(init), .Z(\round_in[0][1039] ) );
  NAND U7676 ( .A(init), .B(round_reg[103]), .Z(n2774) );
  NANDN U7677 ( .A(init), .B(in[103]), .Z(n2773) );
  NAND U7678 ( .A(n2774), .B(n2773), .Z(\round_in[0][103] ) );
  AND U7679 ( .A(round_reg[1040]), .B(init), .Z(\round_in[0][1040] ) );
  AND U7680 ( .A(round_reg[1041]), .B(init), .Z(\round_in[0][1041] ) );
  AND U7681 ( .A(round_reg[1042]), .B(init), .Z(\round_in[0][1042] ) );
  AND U7682 ( .A(round_reg[1043]), .B(init), .Z(\round_in[0][1043] ) );
  AND U7683 ( .A(round_reg[1044]), .B(init), .Z(\round_in[0][1044] ) );
  AND U7684 ( .A(round_reg[1045]), .B(init), .Z(\round_in[0][1045] ) );
  AND U7685 ( .A(round_reg[1046]), .B(init), .Z(\round_in[0][1046] ) );
  AND U7686 ( .A(round_reg[1047]), .B(init), .Z(\round_in[0][1047] ) );
  AND U7687 ( .A(round_reg[1048]), .B(init), .Z(\round_in[0][1048] ) );
  AND U7688 ( .A(round_reg[1049]), .B(init), .Z(\round_in[0][1049] ) );
  NAND U7689 ( .A(init), .B(round_reg[104]), .Z(n2776) );
  NANDN U7690 ( .A(init), .B(in[104]), .Z(n2775) );
  NAND U7691 ( .A(n2776), .B(n2775), .Z(\round_in[0][104] ) );
  AND U7692 ( .A(round_reg[1050]), .B(init), .Z(\round_in[0][1050] ) );
  AND U7693 ( .A(round_reg[1051]), .B(init), .Z(\round_in[0][1051] ) );
  AND U7694 ( .A(round_reg[1052]), .B(init), .Z(\round_in[0][1052] ) );
  AND U7695 ( .A(round_reg[1053]), .B(init), .Z(\round_in[0][1053] ) );
  AND U7696 ( .A(round_reg[1054]), .B(init), .Z(\round_in[0][1054] ) );
  AND U7697 ( .A(round_reg[1055]), .B(init), .Z(\round_in[0][1055] ) );
  AND U7698 ( .A(round_reg[1056]), .B(init), .Z(\round_in[0][1056] ) );
  AND U7699 ( .A(round_reg[1057]), .B(init), .Z(\round_in[0][1057] ) );
  AND U7700 ( .A(round_reg[1058]), .B(init), .Z(\round_in[0][1058] ) );
  AND U7701 ( .A(round_reg[1059]), .B(init), .Z(\round_in[0][1059] ) );
  NAND U7702 ( .A(init), .B(round_reg[105]), .Z(n2778) );
  NANDN U7703 ( .A(init), .B(in[105]), .Z(n2777) );
  NAND U7704 ( .A(n2778), .B(n2777), .Z(\round_in[0][105] ) );
  AND U7705 ( .A(round_reg[1060]), .B(init), .Z(\round_in[0][1060] ) );
  AND U7706 ( .A(round_reg[1061]), .B(init), .Z(\round_in[0][1061] ) );
  AND U7707 ( .A(round_reg[1062]), .B(init), .Z(\round_in[0][1062] ) );
  AND U7708 ( .A(round_reg[1063]), .B(init), .Z(\round_in[0][1063] ) );
  AND U7709 ( .A(round_reg[1064]), .B(init), .Z(\round_in[0][1064] ) );
  AND U7710 ( .A(round_reg[1065]), .B(init), .Z(\round_in[0][1065] ) );
  AND U7711 ( .A(round_reg[1066]), .B(init), .Z(\round_in[0][1066] ) );
  AND U7712 ( .A(round_reg[1067]), .B(init), .Z(\round_in[0][1067] ) );
  AND U7713 ( .A(round_reg[1068]), .B(init), .Z(\round_in[0][1068] ) );
  AND U7714 ( .A(round_reg[1069]), .B(init), .Z(\round_in[0][1069] ) );
  NAND U7715 ( .A(init), .B(round_reg[106]), .Z(n2780) );
  NANDN U7716 ( .A(init), .B(in[106]), .Z(n2779) );
  NAND U7717 ( .A(n2780), .B(n2779), .Z(\round_in[0][106] ) );
  AND U7718 ( .A(round_reg[1070]), .B(init), .Z(\round_in[0][1070] ) );
  AND U7719 ( .A(round_reg[1071]), .B(init), .Z(\round_in[0][1071] ) );
  AND U7720 ( .A(round_reg[1072]), .B(init), .Z(\round_in[0][1072] ) );
  AND U7721 ( .A(round_reg[1073]), .B(init), .Z(\round_in[0][1073] ) );
  AND U7722 ( .A(round_reg[1074]), .B(init), .Z(\round_in[0][1074] ) );
  AND U7723 ( .A(round_reg[1075]), .B(init), .Z(\round_in[0][1075] ) );
  AND U7724 ( .A(round_reg[1076]), .B(init), .Z(\round_in[0][1076] ) );
  AND U7725 ( .A(round_reg[1077]), .B(init), .Z(\round_in[0][1077] ) );
  AND U7726 ( .A(round_reg[1078]), .B(init), .Z(\round_in[0][1078] ) );
  AND U7727 ( .A(round_reg[1079]), .B(init), .Z(\round_in[0][1079] ) );
  NAND U7728 ( .A(init), .B(round_reg[107]), .Z(n2782) );
  NANDN U7729 ( .A(init), .B(in[107]), .Z(n2781) );
  NAND U7730 ( .A(n2782), .B(n2781), .Z(\round_in[0][107] ) );
  AND U7731 ( .A(round_reg[1080]), .B(init), .Z(\round_in[0][1080] ) );
  AND U7732 ( .A(round_reg[1081]), .B(init), .Z(\round_in[0][1081] ) );
  AND U7733 ( .A(round_reg[1082]), .B(init), .Z(\round_in[0][1082] ) );
  AND U7734 ( .A(round_reg[1083]), .B(init), .Z(\round_in[0][1083] ) );
  AND U7735 ( .A(round_reg[1084]), .B(init), .Z(\round_in[0][1084] ) );
  AND U7736 ( .A(round_reg[1085]), .B(init), .Z(\round_in[0][1085] ) );
  AND U7737 ( .A(round_reg[1086]), .B(init), .Z(\round_in[0][1086] ) );
  AND U7738 ( .A(round_reg[1087]), .B(init), .Z(\round_in[0][1087] ) );
  AND U7739 ( .A(round_reg[1088]), .B(init), .Z(\round_in[0][1088] ) );
  AND U7740 ( .A(round_reg[1089]), .B(init), .Z(\round_in[0][1089] ) );
  NAND U7741 ( .A(init), .B(round_reg[108]), .Z(n2784) );
  NANDN U7742 ( .A(init), .B(in[108]), .Z(n2783) );
  NAND U7743 ( .A(n2784), .B(n2783), .Z(\round_in[0][108] ) );
  AND U7744 ( .A(round_reg[1090]), .B(init), .Z(\round_in[0][1090] ) );
  AND U7745 ( .A(round_reg[1091]), .B(init), .Z(\round_in[0][1091] ) );
  AND U7746 ( .A(round_reg[1092]), .B(init), .Z(\round_in[0][1092] ) );
  AND U7747 ( .A(round_reg[1093]), .B(init), .Z(\round_in[0][1093] ) );
  AND U7748 ( .A(round_reg[1094]), .B(init), .Z(\round_in[0][1094] ) );
  AND U7749 ( .A(round_reg[1095]), .B(init), .Z(\round_in[0][1095] ) );
  AND U7750 ( .A(round_reg[1096]), .B(init), .Z(\round_in[0][1096] ) );
  AND U7751 ( .A(round_reg[1097]), .B(init), .Z(\round_in[0][1097] ) );
  AND U7752 ( .A(round_reg[1098]), .B(init), .Z(\round_in[0][1098] ) );
  AND U7753 ( .A(round_reg[1099]), .B(init), .Z(\round_in[0][1099] ) );
  NAND U7754 ( .A(init), .B(round_reg[109]), .Z(n2786) );
  NANDN U7755 ( .A(init), .B(in[109]), .Z(n2785) );
  NAND U7756 ( .A(n2786), .B(n2785), .Z(\round_in[0][109] ) );
  NAND U7757 ( .A(init), .B(round_reg[10]), .Z(n2788) );
  NANDN U7758 ( .A(init), .B(in[10]), .Z(n2787) );
  NAND U7759 ( .A(n2788), .B(n2787), .Z(\round_in[0][10] ) );
  AND U7760 ( .A(round_reg[1100]), .B(init), .Z(\round_in[0][1100] ) );
  AND U7761 ( .A(round_reg[1101]), .B(init), .Z(\round_in[0][1101] ) );
  AND U7762 ( .A(round_reg[1102]), .B(init), .Z(\round_in[0][1102] ) );
  AND U7763 ( .A(round_reg[1103]), .B(init), .Z(\round_in[0][1103] ) );
  AND U7764 ( .A(round_reg[1104]), .B(init), .Z(\round_in[0][1104] ) );
  AND U7765 ( .A(round_reg[1105]), .B(init), .Z(\round_in[0][1105] ) );
  AND U7766 ( .A(round_reg[1106]), .B(init), .Z(\round_in[0][1106] ) );
  AND U7767 ( .A(round_reg[1107]), .B(init), .Z(\round_in[0][1107] ) );
  AND U7768 ( .A(round_reg[1108]), .B(init), .Z(\round_in[0][1108] ) );
  AND U7769 ( .A(round_reg[1109]), .B(init), .Z(\round_in[0][1109] ) );
  NAND U7770 ( .A(init), .B(round_reg[110]), .Z(n2790) );
  NANDN U7771 ( .A(init), .B(in[110]), .Z(n2789) );
  NAND U7772 ( .A(n2790), .B(n2789), .Z(\round_in[0][110] ) );
  AND U7773 ( .A(round_reg[1110]), .B(init), .Z(\round_in[0][1110] ) );
  AND U7774 ( .A(round_reg[1111]), .B(init), .Z(\round_in[0][1111] ) );
  AND U7775 ( .A(round_reg[1112]), .B(init), .Z(\round_in[0][1112] ) );
  AND U7776 ( .A(round_reg[1113]), .B(init), .Z(\round_in[0][1113] ) );
  AND U7777 ( .A(round_reg[1114]), .B(init), .Z(\round_in[0][1114] ) );
  AND U7778 ( .A(round_reg[1115]), .B(init), .Z(\round_in[0][1115] ) );
  AND U7779 ( .A(round_reg[1116]), .B(init), .Z(\round_in[0][1116] ) );
  AND U7780 ( .A(round_reg[1117]), .B(init), .Z(\round_in[0][1117] ) );
  AND U7781 ( .A(round_reg[1118]), .B(init), .Z(\round_in[0][1118] ) );
  AND U7782 ( .A(round_reg[1119]), .B(init), .Z(\round_in[0][1119] ) );
  NAND U7783 ( .A(init), .B(round_reg[111]), .Z(n2792) );
  NANDN U7784 ( .A(init), .B(in[111]), .Z(n2791) );
  NAND U7785 ( .A(n2792), .B(n2791), .Z(\round_in[0][111] ) );
  AND U7786 ( .A(round_reg[1120]), .B(init), .Z(\round_in[0][1120] ) );
  AND U7787 ( .A(round_reg[1121]), .B(init), .Z(\round_in[0][1121] ) );
  AND U7788 ( .A(round_reg[1122]), .B(init), .Z(\round_in[0][1122] ) );
  AND U7789 ( .A(round_reg[1123]), .B(init), .Z(\round_in[0][1123] ) );
  AND U7790 ( .A(round_reg[1124]), .B(init), .Z(\round_in[0][1124] ) );
  AND U7791 ( .A(round_reg[1125]), .B(init), .Z(\round_in[0][1125] ) );
  AND U7792 ( .A(round_reg[1126]), .B(init), .Z(\round_in[0][1126] ) );
  AND U7793 ( .A(round_reg[1127]), .B(init), .Z(\round_in[0][1127] ) );
  AND U7794 ( .A(round_reg[1128]), .B(init), .Z(\round_in[0][1128] ) );
  AND U7795 ( .A(round_reg[1129]), .B(init), .Z(\round_in[0][1129] ) );
  NAND U7796 ( .A(init), .B(round_reg[112]), .Z(n2794) );
  NANDN U7797 ( .A(init), .B(in[112]), .Z(n2793) );
  NAND U7798 ( .A(n2794), .B(n2793), .Z(\round_in[0][112] ) );
  AND U7799 ( .A(round_reg[1130]), .B(init), .Z(\round_in[0][1130] ) );
  AND U7800 ( .A(round_reg[1131]), .B(init), .Z(\round_in[0][1131] ) );
  AND U7801 ( .A(round_reg[1132]), .B(init), .Z(\round_in[0][1132] ) );
  AND U7802 ( .A(round_reg[1133]), .B(init), .Z(\round_in[0][1133] ) );
  AND U7803 ( .A(round_reg[1134]), .B(init), .Z(\round_in[0][1134] ) );
  AND U7804 ( .A(round_reg[1135]), .B(init), .Z(\round_in[0][1135] ) );
  AND U7805 ( .A(round_reg[1136]), .B(init), .Z(\round_in[0][1136] ) );
  AND U7806 ( .A(round_reg[1137]), .B(init), .Z(\round_in[0][1137] ) );
  AND U7807 ( .A(round_reg[1138]), .B(init), .Z(\round_in[0][1138] ) );
  AND U7808 ( .A(round_reg[1139]), .B(init), .Z(\round_in[0][1139] ) );
  NAND U7809 ( .A(init), .B(round_reg[113]), .Z(n2796) );
  NANDN U7810 ( .A(init), .B(in[113]), .Z(n2795) );
  NAND U7811 ( .A(n2796), .B(n2795), .Z(\round_in[0][113] ) );
  AND U7812 ( .A(round_reg[1140]), .B(init), .Z(\round_in[0][1140] ) );
  AND U7813 ( .A(round_reg[1141]), .B(init), .Z(\round_in[0][1141] ) );
  AND U7814 ( .A(round_reg[1142]), .B(init), .Z(\round_in[0][1142] ) );
  AND U7815 ( .A(round_reg[1143]), .B(init), .Z(\round_in[0][1143] ) );
  AND U7816 ( .A(round_reg[1144]), .B(init), .Z(\round_in[0][1144] ) );
  AND U7817 ( .A(round_reg[1145]), .B(init), .Z(\round_in[0][1145] ) );
  AND U7818 ( .A(round_reg[1146]), .B(init), .Z(\round_in[0][1146] ) );
  AND U7819 ( .A(round_reg[1147]), .B(init), .Z(\round_in[0][1147] ) );
  AND U7820 ( .A(round_reg[1148]), .B(init), .Z(\round_in[0][1148] ) );
  AND U7821 ( .A(round_reg[1149]), .B(init), .Z(\round_in[0][1149] ) );
  NAND U7822 ( .A(init), .B(round_reg[114]), .Z(n2798) );
  NANDN U7823 ( .A(init), .B(in[114]), .Z(n2797) );
  NAND U7824 ( .A(n2798), .B(n2797), .Z(\round_in[0][114] ) );
  AND U7825 ( .A(round_reg[1150]), .B(init), .Z(\round_in[0][1150] ) );
  AND U7826 ( .A(round_reg[1151]), .B(init), .Z(\round_in[0][1151] ) );
  AND U7827 ( .A(round_reg[1152]), .B(init), .Z(\round_in[0][1152] ) );
  AND U7828 ( .A(round_reg[1153]), .B(init), .Z(\round_in[0][1153] ) );
  AND U7829 ( .A(round_reg[1154]), .B(init), .Z(\round_in[0][1154] ) );
  AND U7830 ( .A(round_reg[1155]), .B(init), .Z(\round_in[0][1155] ) );
  AND U7831 ( .A(round_reg[1156]), .B(init), .Z(\round_in[0][1156] ) );
  AND U7832 ( .A(round_reg[1157]), .B(init), .Z(\round_in[0][1157] ) );
  AND U7833 ( .A(round_reg[1158]), .B(init), .Z(\round_in[0][1158] ) );
  AND U7834 ( .A(round_reg[1159]), .B(init), .Z(\round_in[0][1159] ) );
  NAND U7835 ( .A(init), .B(round_reg[115]), .Z(n2800) );
  NANDN U7836 ( .A(init), .B(in[115]), .Z(n2799) );
  NAND U7837 ( .A(n2800), .B(n2799), .Z(\round_in[0][115] ) );
  AND U7838 ( .A(round_reg[1160]), .B(init), .Z(\round_in[0][1160] ) );
  AND U7839 ( .A(round_reg[1161]), .B(init), .Z(\round_in[0][1161] ) );
  AND U7840 ( .A(round_reg[1162]), .B(init), .Z(\round_in[0][1162] ) );
  AND U7841 ( .A(round_reg[1163]), .B(init), .Z(\round_in[0][1163] ) );
  AND U7842 ( .A(round_reg[1164]), .B(init), .Z(\round_in[0][1164] ) );
  AND U7843 ( .A(round_reg[1165]), .B(init), .Z(\round_in[0][1165] ) );
  AND U7844 ( .A(round_reg[1166]), .B(init), .Z(\round_in[0][1166] ) );
  AND U7845 ( .A(round_reg[1167]), .B(init), .Z(\round_in[0][1167] ) );
  AND U7846 ( .A(round_reg[1168]), .B(init), .Z(\round_in[0][1168] ) );
  AND U7847 ( .A(round_reg[1169]), .B(init), .Z(\round_in[0][1169] ) );
  NAND U7848 ( .A(init), .B(round_reg[116]), .Z(n2802) );
  NANDN U7849 ( .A(init), .B(in[116]), .Z(n2801) );
  NAND U7850 ( .A(n2802), .B(n2801), .Z(\round_in[0][116] ) );
  AND U7851 ( .A(round_reg[1170]), .B(init), .Z(\round_in[0][1170] ) );
  AND U7852 ( .A(round_reg[1171]), .B(init), .Z(\round_in[0][1171] ) );
  AND U7853 ( .A(round_reg[1172]), .B(init), .Z(\round_in[0][1172] ) );
  AND U7854 ( .A(round_reg[1173]), .B(init), .Z(\round_in[0][1173] ) );
  AND U7855 ( .A(round_reg[1174]), .B(init), .Z(\round_in[0][1174] ) );
  AND U7856 ( .A(round_reg[1175]), .B(init), .Z(\round_in[0][1175] ) );
  AND U7857 ( .A(round_reg[1176]), .B(init), .Z(\round_in[0][1176] ) );
  AND U7858 ( .A(round_reg[1177]), .B(init), .Z(\round_in[0][1177] ) );
  AND U7859 ( .A(round_reg[1178]), .B(init), .Z(\round_in[0][1178] ) );
  AND U7860 ( .A(round_reg[1179]), .B(init), .Z(\round_in[0][1179] ) );
  NAND U7861 ( .A(init), .B(round_reg[117]), .Z(n2804) );
  NANDN U7862 ( .A(init), .B(in[117]), .Z(n2803) );
  NAND U7863 ( .A(n2804), .B(n2803), .Z(\round_in[0][117] ) );
  AND U7864 ( .A(round_reg[1180]), .B(init), .Z(\round_in[0][1180] ) );
  AND U7865 ( .A(round_reg[1181]), .B(init), .Z(\round_in[0][1181] ) );
  AND U7866 ( .A(round_reg[1182]), .B(init), .Z(\round_in[0][1182] ) );
  AND U7867 ( .A(round_reg[1183]), .B(init), .Z(\round_in[0][1183] ) );
  AND U7868 ( .A(round_reg[1184]), .B(init), .Z(\round_in[0][1184] ) );
  AND U7869 ( .A(round_reg[1185]), .B(init), .Z(\round_in[0][1185] ) );
  AND U7870 ( .A(round_reg[1186]), .B(init), .Z(\round_in[0][1186] ) );
  AND U7871 ( .A(round_reg[1187]), .B(init), .Z(\round_in[0][1187] ) );
  AND U7872 ( .A(round_reg[1188]), .B(init), .Z(\round_in[0][1188] ) );
  AND U7873 ( .A(round_reg[1189]), .B(init), .Z(\round_in[0][1189] ) );
  NAND U7874 ( .A(init), .B(round_reg[118]), .Z(n2806) );
  NANDN U7875 ( .A(init), .B(in[118]), .Z(n2805) );
  NAND U7876 ( .A(n2806), .B(n2805), .Z(\round_in[0][118] ) );
  AND U7877 ( .A(round_reg[1190]), .B(init), .Z(\round_in[0][1190] ) );
  AND U7878 ( .A(round_reg[1191]), .B(init), .Z(\round_in[0][1191] ) );
  AND U7879 ( .A(round_reg[1192]), .B(init), .Z(\round_in[0][1192] ) );
  AND U7880 ( .A(round_reg[1193]), .B(init), .Z(\round_in[0][1193] ) );
  AND U7881 ( .A(round_reg[1194]), .B(init), .Z(\round_in[0][1194] ) );
  AND U7882 ( .A(round_reg[1195]), .B(init), .Z(\round_in[0][1195] ) );
  AND U7883 ( .A(round_reg[1196]), .B(init), .Z(\round_in[0][1196] ) );
  AND U7884 ( .A(round_reg[1197]), .B(init), .Z(\round_in[0][1197] ) );
  AND U7885 ( .A(round_reg[1198]), .B(init), .Z(\round_in[0][1198] ) );
  AND U7886 ( .A(round_reg[1199]), .B(init), .Z(\round_in[0][1199] ) );
  NAND U7887 ( .A(init), .B(round_reg[119]), .Z(n2808) );
  NANDN U7888 ( .A(init), .B(in[119]), .Z(n2807) );
  NAND U7889 ( .A(n2808), .B(n2807), .Z(\round_in[0][119] ) );
  NAND U7890 ( .A(init), .B(round_reg[11]), .Z(n2810) );
  NANDN U7891 ( .A(init), .B(in[11]), .Z(n2809) );
  NAND U7892 ( .A(n2810), .B(n2809), .Z(\round_in[0][11] ) );
  AND U7893 ( .A(round_reg[1200]), .B(init), .Z(\round_in[0][1200] ) );
  AND U7894 ( .A(round_reg[1201]), .B(init), .Z(\round_in[0][1201] ) );
  AND U7895 ( .A(round_reg[1202]), .B(init), .Z(\round_in[0][1202] ) );
  AND U7896 ( .A(round_reg[1203]), .B(init), .Z(\round_in[0][1203] ) );
  AND U7897 ( .A(round_reg[1204]), .B(init), .Z(\round_in[0][1204] ) );
  AND U7898 ( .A(round_reg[1205]), .B(init), .Z(\round_in[0][1205] ) );
  AND U7899 ( .A(round_reg[1206]), .B(init), .Z(\round_in[0][1206] ) );
  AND U7900 ( .A(round_reg[1207]), .B(init), .Z(\round_in[0][1207] ) );
  AND U7901 ( .A(round_reg[1208]), .B(init), .Z(\round_in[0][1208] ) );
  AND U7902 ( .A(round_reg[1209]), .B(init), .Z(\round_in[0][1209] ) );
  NAND U7903 ( .A(init), .B(round_reg[120]), .Z(n2812) );
  NANDN U7904 ( .A(init), .B(in[120]), .Z(n2811) );
  NAND U7905 ( .A(n2812), .B(n2811), .Z(\round_in[0][120] ) );
  AND U7906 ( .A(round_reg[1210]), .B(init), .Z(\round_in[0][1210] ) );
  AND U7907 ( .A(round_reg[1211]), .B(init), .Z(\round_in[0][1211] ) );
  AND U7908 ( .A(round_reg[1212]), .B(init), .Z(\round_in[0][1212] ) );
  AND U7909 ( .A(round_reg[1213]), .B(init), .Z(\round_in[0][1213] ) );
  AND U7910 ( .A(round_reg[1214]), .B(init), .Z(\round_in[0][1214] ) );
  AND U7911 ( .A(round_reg[1215]), .B(init), .Z(\round_in[0][1215] ) );
  AND U7912 ( .A(round_reg[1216]), .B(init), .Z(\round_in[0][1216] ) );
  AND U7913 ( .A(round_reg[1217]), .B(init), .Z(\round_in[0][1217] ) );
  AND U7914 ( .A(round_reg[1218]), .B(init), .Z(\round_in[0][1218] ) );
  AND U7915 ( .A(round_reg[1219]), .B(init), .Z(\round_in[0][1219] ) );
  NAND U7916 ( .A(init), .B(round_reg[121]), .Z(n2814) );
  NANDN U7917 ( .A(init), .B(in[121]), .Z(n2813) );
  NAND U7918 ( .A(n2814), .B(n2813), .Z(\round_in[0][121] ) );
  AND U7919 ( .A(round_reg[1220]), .B(init), .Z(\round_in[0][1220] ) );
  AND U7920 ( .A(round_reg[1221]), .B(init), .Z(\round_in[0][1221] ) );
  AND U7921 ( .A(round_reg[1222]), .B(init), .Z(\round_in[0][1222] ) );
  AND U7922 ( .A(round_reg[1223]), .B(init), .Z(\round_in[0][1223] ) );
  AND U7923 ( .A(round_reg[1224]), .B(init), .Z(\round_in[0][1224] ) );
  AND U7924 ( .A(round_reg[1225]), .B(init), .Z(\round_in[0][1225] ) );
  AND U7925 ( .A(round_reg[1226]), .B(init), .Z(\round_in[0][1226] ) );
  AND U7926 ( .A(round_reg[1227]), .B(init), .Z(\round_in[0][1227] ) );
  AND U7927 ( .A(round_reg[1228]), .B(init), .Z(\round_in[0][1228] ) );
  AND U7928 ( .A(round_reg[1229]), .B(init), .Z(\round_in[0][1229] ) );
  NAND U7929 ( .A(init), .B(round_reg[122]), .Z(n2816) );
  NANDN U7930 ( .A(init), .B(in[122]), .Z(n2815) );
  NAND U7931 ( .A(n2816), .B(n2815), .Z(\round_in[0][122] ) );
  AND U7932 ( .A(round_reg[1230]), .B(init), .Z(\round_in[0][1230] ) );
  AND U7933 ( .A(round_reg[1231]), .B(init), .Z(\round_in[0][1231] ) );
  AND U7934 ( .A(round_reg[1232]), .B(init), .Z(\round_in[0][1232] ) );
  AND U7935 ( .A(round_reg[1233]), .B(init), .Z(\round_in[0][1233] ) );
  AND U7936 ( .A(round_reg[1234]), .B(init), .Z(\round_in[0][1234] ) );
  AND U7937 ( .A(round_reg[1235]), .B(init), .Z(\round_in[0][1235] ) );
  AND U7938 ( .A(round_reg[1236]), .B(init), .Z(\round_in[0][1236] ) );
  AND U7939 ( .A(round_reg[1237]), .B(init), .Z(\round_in[0][1237] ) );
  AND U7940 ( .A(round_reg[1238]), .B(init), .Z(\round_in[0][1238] ) );
  AND U7941 ( .A(round_reg[1239]), .B(init), .Z(\round_in[0][1239] ) );
  NAND U7942 ( .A(init), .B(round_reg[123]), .Z(n2818) );
  NANDN U7943 ( .A(init), .B(in[123]), .Z(n2817) );
  NAND U7944 ( .A(n2818), .B(n2817), .Z(\round_in[0][123] ) );
  AND U7945 ( .A(round_reg[1240]), .B(init), .Z(\round_in[0][1240] ) );
  AND U7946 ( .A(round_reg[1241]), .B(init), .Z(\round_in[0][1241] ) );
  AND U7947 ( .A(round_reg[1242]), .B(init), .Z(\round_in[0][1242] ) );
  AND U7948 ( .A(round_reg[1243]), .B(init), .Z(\round_in[0][1243] ) );
  AND U7949 ( .A(round_reg[1244]), .B(init), .Z(\round_in[0][1244] ) );
  AND U7950 ( .A(round_reg[1245]), .B(init), .Z(\round_in[0][1245] ) );
  AND U7951 ( .A(round_reg[1246]), .B(init), .Z(\round_in[0][1246] ) );
  AND U7952 ( .A(round_reg[1247]), .B(init), .Z(\round_in[0][1247] ) );
  AND U7953 ( .A(round_reg[1248]), .B(init), .Z(\round_in[0][1248] ) );
  AND U7954 ( .A(round_reg[1249]), .B(init), .Z(\round_in[0][1249] ) );
  NAND U7955 ( .A(init), .B(round_reg[124]), .Z(n2820) );
  NANDN U7956 ( .A(init), .B(in[124]), .Z(n2819) );
  NAND U7957 ( .A(n2820), .B(n2819), .Z(\round_in[0][124] ) );
  AND U7958 ( .A(round_reg[1250]), .B(init), .Z(\round_in[0][1250] ) );
  AND U7959 ( .A(round_reg[1251]), .B(init), .Z(\round_in[0][1251] ) );
  AND U7960 ( .A(round_reg[1252]), .B(init), .Z(\round_in[0][1252] ) );
  AND U7961 ( .A(round_reg[1253]), .B(init), .Z(\round_in[0][1253] ) );
  AND U7962 ( .A(round_reg[1254]), .B(init), .Z(\round_in[0][1254] ) );
  AND U7963 ( .A(round_reg[1255]), .B(init), .Z(\round_in[0][1255] ) );
  AND U7964 ( .A(round_reg[1256]), .B(init), .Z(\round_in[0][1256] ) );
  AND U7965 ( .A(round_reg[1257]), .B(init), .Z(\round_in[0][1257] ) );
  AND U7966 ( .A(round_reg[1258]), .B(init), .Z(\round_in[0][1258] ) );
  AND U7967 ( .A(round_reg[1259]), .B(init), .Z(\round_in[0][1259] ) );
  NAND U7968 ( .A(init), .B(round_reg[125]), .Z(n2822) );
  NANDN U7969 ( .A(init), .B(in[125]), .Z(n2821) );
  NAND U7970 ( .A(n2822), .B(n2821), .Z(\round_in[0][125] ) );
  AND U7971 ( .A(round_reg[1260]), .B(init), .Z(\round_in[0][1260] ) );
  AND U7972 ( .A(round_reg[1261]), .B(init), .Z(\round_in[0][1261] ) );
  AND U7973 ( .A(round_reg[1262]), .B(init), .Z(\round_in[0][1262] ) );
  AND U7974 ( .A(round_reg[1263]), .B(init), .Z(\round_in[0][1263] ) );
  AND U7975 ( .A(round_reg[1264]), .B(init), .Z(\round_in[0][1264] ) );
  AND U7976 ( .A(round_reg[1265]), .B(init), .Z(\round_in[0][1265] ) );
  AND U7977 ( .A(round_reg[1266]), .B(init), .Z(\round_in[0][1266] ) );
  AND U7978 ( .A(round_reg[1267]), .B(init), .Z(\round_in[0][1267] ) );
  AND U7979 ( .A(round_reg[1268]), .B(init), .Z(\round_in[0][1268] ) );
  AND U7980 ( .A(round_reg[1269]), .B(init), .Z(\round_in[0][1269] ) );
  NAND U7981 ( .A(init), .B(round_reg[126]), .Z(n2824) );
  NANDN U7982 ( .A(init), .B(in[126]), .Z(n2823) );
  NAND U7983 ( .A(n2824), .B(n2823), .Z(\round_in[0][126] ) );
  AND U7984 ( .A(round_reg[1270]), .B(init), .Z(\round_in[0][1270] ) );
  AND U7985 ( .A(round_reg[1271]), .B(init), .Z(\round_in[0][1271] ) );
  AND U7986 ( .A(round_reg[1272]), .B(init), .Z(\round_in[0][1272] ) );
  AND U7987 ( .A(round_reg[1273]), .B(init), .Z(\round_in[0][1273] ) );
  AND U7988 ( .A(round_reg[1274]), .B(init), .Z(\round_in[0][1274] ) );
  AND U7989 ( .A(round_reg[1275]), .B(init), .Z(\round_in[0][1275] ) );
  AND U7990 ( .A(round_reg[1276]), .B(init), .Z(\round_in[0][1276] ) );
  AND U7991 ( .A(round_reg[1277]), .B(init), .Z(\round_in[0][1277] ) );
  AND U7992 ( .A(round_reg[1278]), .B(init), .Z(\round_in[0][1278] ) );
  AND U7993 ( .A(round_reg[1279]), .B(init), .Z(\round_in[0][1279] ) );
  NAND U7994 ( .A(init), .B(round_reg[127]), .Z(n2826) );
  NANDN U7995 ( .A(init), .B(in[127]), .Z(n2825) );
  NAND U7996 ( .A(n2826), .B(n2825), .Z(\round_in[0][127] ) );
  AND U7997 ( .A(round_reg[1280]), .B(init), .Z(\round_in[0][1280] ) );
  AND U7998 ( .A(round_reg[1281]), .B(init), .Z(\round_in[0][1281] ) );
  AND U7999 ( .A(round_reg[1282]), .B(init), .Z(\round_in[0][1282] ) );
  AND U8000 ( .A(round_reg[1283]), .B(init), .Z(\round_in[0][1283] ) );
  AND U8001 ( .A(round_reg[1284]), .B(init), .Z(\round_in[0][1284] ) );
  AND U8002 ( .A(round_reg[1285]), .B(init), .Z(\round_in[0][1285] ) );
  AND U8003 ( .A(round_reg[1286]), .B(init), .Z(\round_in[0][1286] ) );
  AND U8004 ( .A(round_reg[1287]), .B(init), .Z(\round_in[0][1287] ) );
  AND U8005 ( .A(round_reg[1288]), .B(init), .Z(\round_in[0][1288] ) );
  AND U8006 ( .A(round_reg[1289]), .B(init), .Z(\round_in[0][1289] ) );
  NAND U8007 ( .A(init), .B(round_reg[128]), .Z(n2828) );
  NANDN U8008 ( .A(init), .B(in[128]), .Z(n2827) );
  NAND U8009 ( .A(n2828), .B(n2827), .Z(\round_in[0][128] ) );
  AND U8010 ( .A(round_reg[1290]), .B(init), .Z(\round_in[0][1290] ) );
  AND U8011 ( .A(round_reg[1291]), .B(init), .Z(\round_in[0][1291] ) );
  AND U8012 ( .A(round_reg[1292]), .B(init), .Z(\round_in[0][1292] ) );
  AND U8013 ( .A(round_reg[1293]), .B(init), .Z(\round_in[0][1293] ) );
  AND U8014 ( .A(round_reg[1294]), .B(init), .Z(\round_in[0][1294] ) );
  AND U8015 ( .A(round_reg[1295]), .B(init), .Z(\round_in[0][1295] ) );
  AND U8016 ( .A(round_reg[1296]), .B(init), .Z(\round_in[0][1296] ) );
  AND U8017 ( .A(round_reg[1297]), .B(init), .Z(\round_in[0][1297] ) );
  AND U8018 ( .A(round_reg[1298]), .B(init), .Z(\round_in[0][1298] ) );
  AND U8019 ( .A(round_reg[1299]), .B(init), .Z(\round_in[0][1299] ) );
  NAND U8020 ( .A(init), .B(round_reg[129]), .Z(n2830) );
  NANDN U8021 ( .A(init), .B(in[129]), .Z(n2829) );
  NAND U8022 ( .A(n2830), .B(n2829), .Z(\round_in[0][129] ) );
  NAND U8023 ( .A(init), .B(round_reg[12]), .Z(n2832) );
  NANDN U8024 ( .A(init), .B(in[12]), .Z(n2831) );
  NAND U8025 ( .A(n2832), .B(n2831), .Z(\round_in[0][12] ) );
  AND U8026 ( .A(round_reg[1300]), .B(init), .Z(\round_in[0][1300] ) );
  AND U8027 ( .A(round_reg[1301]), .B(init), .Z(\round_in[0][1301] ) );
  AND U8028 ( .A(round_reg[1302]), .B(init), .Z(\round_in[0][1302] ) );
  AND U8029 ( .A(round_reg[1303]), .B(init), .Z(\round_in[0][1303] ) );
  AND U8030 ( .A(round_reg[1304]), .B(init), .Z(\round_in[0][1304] ) );
  AND U8031 ( .A(round_reg[1305]), .B(init), .Z(\round_in[0][1305] ) );
  AND U8032 ( .A(round_reg[1306]), .B(init), .Z(\round_in[0][1306] ) );
  AND U8033 ( .A(round_reg[1307]), .B(init), .Z(\round_in[0][1307] ) );
  AND U8034 ( .A(round_reg[1308]), .B(init), .Z(\round_in[0][1308] ) );
  AND U8035 ( .A(round_reg[1309]), .B(init), .Z(\round_in[0][1309] ) );
  NAND U8036 ( .A(init), .B(round_reg[130]), .Z(n2834) );
  NANDN U8037 ( .A(init), .B(in[130]), .Z(n2833) );
  NAND U8038 ( .A(n2834), .B(n2833), .Z(\round_in[0][130] ) );
  AND U8039 ( .A(round_reg[1310]), .B(init), .Z(\round_in[0][1310] ) );
  AND U8040 ( .A(round_reg[1311]), .B(init), .Z(\round_in[0][1311] ) );
  AND U8041 ( .A(round_reg[1312]), .B(init), .Z(\round_in[0][1312] ) );
  AND U8042 ( .A(round_reg[1313]), .B(init), .Z(\round_in[0][1313] ) );
  AND U8043 ( .A(round_reg[1314]), .B(init), .Z(\round_in[0][1314] ) );
  AND U8044 ( .A(round_reg[1315]), .B(init), .Z(\round_in[0][1315] ) );
  AND U8045 ( .A(round_reg[1316]), .B(init), .Z(\round_in[0][1316] ) );
  AND U8046 ( .A(round_reg[1317]), .B(init), .Z(\round_in[0][1317] ) );
  AND U8047 ( .A(round_reg[1318]), .B(init), .Z(\round_in[0][1318] ) );
  AND U8048 ( .A(round_reg[1319]), .B(init), .Z(\round_in[0][1319] ) );
  NAND U8049 ( .A(init), .B(round_reg[131]), .Z(n2836) );
  NANDN U8050 ( .A(init), .B(in[131]), .Z(n2835) );
  NAND U8051 ( .A(n2836), .B(n2835), .Z(\round_in[0][131] ) );
  AND U8052 ( .A(round_reg[1320]), .B(init), .Z(\round_in[0][1320] ) );
  AND U8053 ( .A(round_reg[1321]), .B(init), .Z(\round_in[0][1321] ) );
  AND U8054 ( .A(round_reg[1322]), .B(init), .Z(\round_in[0][1322] ) );
  AND U8055 ( .A(round_reg[1323]), .B(init), .Z(\round_in[0][1323] ) );
  AND U8056 ( .A(round_reg[1324]), .B(init), .Z(\round_in[0][1324] ) );
  AND U8057 ( .A(round_reg[1325]), .B(init), .Z(\round_in[0][1325] ) );
  AND U8058 ( .A(round_reg[1326]), .B(init), .Z(\round_in[0][1326] ) );
  AND U8059 ( .A(round_reg[1327]), .B(init), .Z(\round_in[0][1327] ) );
  AND U8060 ( .A(round_reg[1328]), .B(init), .Z(\round_in[0][1328] ) );
  AND U8061 ( .A(round_reg[1329]), .B(init), .Z(\round_in[0][1329] ) );
  NAND U8062 ( .A(init), .B(round_reg[132]), .Z(n2838) );
  NANDN U8063 ( .A(init), .B(in[132]), .Z(n2837) );
  NAND U8064 ( .A(n2838), .B(n2837), .Z(\round_in[0][132] ) );
  AND U8065 ( .A(round_reg[1330]), .B(init), .Z(\round_in[0][1330] ) );
  AND U8066 ( .A(round_reg[1331]), .B(init), .Z(\round_in[0][1331] ) );
  AND U8067 ( .A(round_reg[1332]), .B(init), .Z(\round_in[0][1332] ) );
  AND U8068 ( .A(round_reg[1333]), .B(init), .Z(\round_in[0][1333] ) );
  AND U8069 ( .A(round_reg[1334]), .B(init), .Z(\round_in[0][1334] ) );
  AND U8070 ( .A(round_reg[1335]), .B(init), .Z(\round_in[0][1335] ) );
  AND U8071 ( .A(round_reg[1336]), .B(init), .Z(\round_in[0][1336] ) );
  AND U8072 ( .A(round_reg[1337]), .B(init), .Z(\round_in[0][1337] ) );
  AND U8073 ( .A(round_reg[1338]), .B(init), .Z(\round_in[0][1338] ) );
  AND U8074 ( .A(round_reg[1339]), .B(init), .Z(\round_in[0][1339] ) );
  NAND U8075 ( .A(init), .B(round_reg[133]), .Z(n2840) );
  NANDN U8076 ( .A(init), .B(in[133]), .Z(n2839) );
  NAND U8077 ( .A(n2840), .B(n2839), .Z(\round_in[0][133] ) );
  AND U8078 ( .A(round_reg[1340]), .B(init), .Z(\round_in[0][1340] ) );
  AND U8079 ( .A(round_reg[1341]), .B(init), .Z(\round_in[0][1341] ) );
  AND U8080 ( .A(round_reg[1342]), .B(init), .Z(\round_in[0][1342] ) );
  AND U8081 ( .A(round_reg[1343]), .B(init), .Z(\round_in[0][1343] ) );
  AND U8082 ( .A(round_reg[1344]), .B(init), .Z(\round_in[0][1344] ) );
  AND U8083 ( .A(round_reg[1345]), .B(init), .Z(\round_in[0][1345] ) );
  AND U8084 ( .A(round_reg[1346]), .B(init), .Z(\round_in[0][1346] ) );
  AND U8085 ( .A(round_reg[1347]), .B(init), .Z(\round_in[0][1347] ) );
  AND U8086 ( .A(round_reg[1348]), .B(init), .Z(\round_in[0][1348] ) );
  AND U8087 ( .A(round_reg[1349]), .B(init), .Z(\round_in[0][1349] ) );
  NAND U8088 ( .A(init), .B(round_reg[134]), .Z(n2842) );
  NANDN U8089 ( .A(init), .B(in[134]), .Z(n2841) );
  NAND U8090 ( .A(n2842), .B(n2841), .Z(\round_in[0][134] ) );
  AND U8091 ( .A(round_reg[1350]), .B(init), .Z(\round_in[0][1350] ) );
  AND U8092 ( .A(round_reg[1351]), .B(init), .Z(\round_in[0][1351] ) );
  AND U8093 ( .A(round_reg[1352]), .B(init), .Z(\round_in[0][1352] ) );
  AND U8094 ( .A(round_reg[1353]), .B(init), .Z(\round_in[0][1353] ) );
  AND U8095 ( .A(round_reg[1354]), .B(init), .Z(\round_in[0][1354] ) );
  AND U8096 ( .A(round_reg[1355]), .B(init), .Z(\round_in[0][1355] ) );
  AND U8097 ( .A(round_reg[1356]), .B(init), .Z(\round_in[0][1356] ) );
  AND U8098 ( .A(round_reg[1357]), .B(init), .Z(\round_in[0][1357] ) );
  AND U8099 ( .A(round_reg[1358]), .B(init), .Z(\round_in[0][1358] ) );
  AND U8100 ( .A(round_reg[1359]), .B(init), .Z(\round_in[0][1359] ) );
  NAND U8101 ( .A(init), .B(round_reg[135]), .Z(n2844) );
  NANDN U8102 ( .A(init), .B(in[135]), .Z(n2843) );
  NAND U8103 ( .A(n2844), .B(n2843), .Z(\round_in[0][135] ) );
  AND U8104 ( .A(round_reg[1360]), .B(init), .Z(\round_in[0][1360] ) );
  AND U8105 ( .A(round_reg[1361]), .B(init), .Z(\round_in[0][1361] ) );
  AND U8106 ( .A(round_reg[1362]), .B(init), .Z(\round_in[0][1362] ) );
  AND U8107 ( .A(round_reg[1363]), .B(init), .Z(\round_in[0][1363] ) );
  AND U8108 ( .A(round_reg[1364]), .B(init), .Z(\round_in[0][1364] ) );
  AND U8109 ( .A(round_reg[1365]), .B(init), .Z(\round_in[0][1365] ) );
  AND U8110 ( .A(round_reg[1366]), .B(init), .Z(\round_in[0][1366] ) );
  AND U8111 ( .A(round_reg[1367]), .B(init), .Z(\round_in[0][1367] ) );
  AND U8112 ( .A(round_reg[1368]), .B(init), .Z(\round_in[0][1368] ) );
  AND U8113 ( .A(round_reg[1369]), .B(init), .Z(\round_in[0][1369] ) );
  NAND U8114 ( .A(init), .B(round_reg[136]), .Z(n2846) );
  NANDN U8115 ( .A(init), .B(in[136]), .Z(n2845) );
  NAND U8116 ( .A(n2846), .B(n2845), .Z(\round_in[0][136] ) );
  AND U8117 ( .A(round_reg[1370]), .B(init), .Z(\round_in[0][1370] ) );
  AND U8118 ( .A(round_reg[1371]), .B(init), .Z(\round_in[0][1371] ) );
  AND U8119 ( .A(round_reg[1372]), .B(init), .Z(\round_in[0][1372] ) );
  AND U8120 ( .A(round_reg[1373]), .B(init), .Z(\round_in[0][1373] ) );
  AND U8121 ( .A(round_reg[1374]), .B(init), .Z(\round_in[0][1374] ) );
  AND U8122 ( .A(round_reg[1375]), .B(init), .Z(\round_in[0][1375] ) );
  AND U8123 ( .A(round_reg[1376]), .B(init), .Z(\round_in[0][1376] ) );
  AND U8124 ( .A(round_reg[1377]), .B(init), .Z(\round_in[0][1377] ) );
  AND U8125 ( .A(round_reg[1378]), .B(init), .Z(\round_in[0][1378] ) );
  AND U8126 ( .A(round_reg[1379]), .B(init), .Z(\round_in[0][1379] ) );
  NAND U8127 ( .A(init), .B(round_reg[137]), .Z(n2848) );
  NANDN U8128 ( .A(init), .B(in[137]), .Z(n2847) );
  NAND U8129 ( .A(n2848), .B(n2847), .Z(\round_in[0][137] ) );
  AND U8130 ( .A(round_reg[1380]), .B(init), .Z(\round_in[0][1380] ) );
  AND U8131 ( .A(round_reg[1381]), .B(init), .Z(\round_in[0][1381] ) );
  AND U8132 ( .A(round_reg[1382]), .B(init), .Z(\round_in[0][1382] ) );
  AND U8133 ( .A(round_reg[1383]), .B(init), .Z(\round_in[0][1383] ) );
  AND U8134 ( .A(round_reg[1384]), .B(init), .Z(\round_in[0][1384] ) );
  AND U8135 ( .A(round_reg[1385]), .B(init), .Z(\round_in[0][1385] ) );
  AND U8136 ( .A(round_reg[1386]), .B(init), .Z(\round_in[0][1386] ) );
  AND U8137 ( .A(round_reg[1387]), .B(init), .Z(\round_in[0][1387] ) );
  AND U8138 ( .A(round_reg[1388]), .B(init), .Z(\round_in[0][1388] ) );
  AND U8139 ( .A(round_reg[1389]), .B(init), .Z(\round_in[0][1389] ) );
  NAND U8140 ( .A(init), .B(round_reg[138]), .Z(n2850) );
  NANDN U8141 ( .A(init), .B(in[138]), .Z(n2849) );
  NAND U8142 ( .A(n2850), .B(n2849), .Z(\round_in[0][138] ) );
  AND U8143 ( .A(round_reg[1390]), .B(init), .Z(\round_in[0][1390] ) );
  AND U8144 ( .A(round_reg[1391]), .B(init), .Z(\round_in[0][1391] ) );
  AND U8145 ( .A(round_reg[1392]), .B(init), .Z(\round_in[0][1392] ) );
  AND U8146 ( .A(round_reg[1393]), .B(init), .Z(\round_in[0][1393] ) );
  AND U8147 ( .A(round_reg[1394]), .B(init), .Z(\round_in[0][1394] ) );
  AND U8148 ( .A(round_reg[1395]), .B(init), .Z(\round_in[0][1395] ) );
  AND U8149 ( .A(round_reg[1396]), .B(init), .Z(\round_in[0][1396] ) );
  AND U8150 ( .A(round_reg[1397]), .B(init), .Z(\round_in[0][1397] ) );
  AND U8151 ( .A(round_reg[1398]), .B(init), .Z(\round_in[0][1398] ) );
  AND U8152 ( .A(round_reg[1399]), .B(init), .Z(\round_in[0][1399] ) );
  NAND U8153 ( .A(init), .B(round_reg[139]), .Z(n2852) );
  NANDN U8154 ( .A(init), .B(in[139]), .Z(n2851) );
  NAND U8155 ( .A(n2852), .B(n2851), .Z(\round_in[0][139] ) );
  NAND U8156 ( .A(init), .B(round_reg[13]), .Z(n2854) );
  NANDN U8157 ( .A(init), .B(in[13]), .Z(n2853) );
  NAND U8158 ( .A(n2854), .B(n2853), .Z(\round_in[0][13] ) );
  AND U8159 ( .A(round_reg[1400]), .B(init), .Z(\round_in[0][1400] ) );
  AND U8160 ( .A(round_reg[1401]), .B(init), .Z(\round_in[0][1401] ) );
  AND U8161 ( .A(round_reg[1402]), .B(init), .Z(\round_in[0][1402] ) );
  AND U8162 ( .A(round_reg[1403]), .B(init), .Z(\round_in[0][1403] ) );
  AND U8163 ( .A(round_reg[1404]), .B(init), .Z(\round_in[0][1404] ) );
  AND U8164 ( .A(round_reg[1405]), .B(init), .Z(\round_in[0][1405] ) );
  AND U8165 ( .A(round_reg[1406]), .B(init), .Z(\round_in[0][1406] ) );
  AND U8166 ( .A(round_reg[1407]), .B(init), .Z(\round_in[0][1407] ) );
  AND U8167 ( .A(round_reg[1408]), .B(init), .Z(\round_in[0][1408] ) );
  AND U8168 ( .A(round_reg[1409]), .B(init), .Z(\round_in[0][1409] ) );
  NAND U8169 ( .A(init), .B(round_reg[140]), .Z(n2856) );
  NANDN U8170 ( .A(init), .B(in[140]), .Z(n2855) );
  NAND U8171 ( .A(n2856), .B(n2855), .Z(\round_in[0][140] ) );
  AND U8172 ( .A(round_reg[1410]), .B(init), .Z(\round_in[0][1410] ) );
  AND U8173 ( .A(round_reg[1411]), .B(init), .Z(\round_in[0][1411] ) );
  AND U8174 ( .A(round_reg[1412]), .B(init), .Z(\round_in[0][1412] ) );
  AND U8175 ( .A(round_reg[1413]), .B(init), .Z(\round_in[0][1413] ) );
  AND U8176 ( .A(round_reg[1414]), .B(init), .Z(\round_in[0][1414] ) );
  AND U8177 ( .A(round_reg[1415]), .B(init), .Z(\round_in[0][1415] ) );
  AND U8178 ( .A(round_reg[1416]), .B(init), .Z(\round_in[0][1416] ) );
  AND U8179 ( .A(round_reg[1417]), .B(init), .Z(\round_in[0][1417] ) );
  AND U8180 ( .A(round_reg[1418]), .B(init), .Z(\round_in[0][1418] ) );
  AND U8181 ( .A(round_reg[1419]), .B(init), .Z(\round_in[0][1419] ) );
  NAND U8182 ( .A(init), .B(round_reg[141]), .Z(n2858) );
  NANDN U8183 ( .A(init), .B(in[141]), .Z(n2857) );
  NAND U8184 ( .A(n2858), .B(n2857), .Z(\round_in[0][141] ) );
  AND U8185 ( .A(round_reg[1420]), .B(init), .Z(\round_in[0][1420] ) );
  AND U8186 ( .A(round_reg[1421]), .B(init), .Z(\round_in[0][1421] ) );
  AND U8187 ( .A(round_reg[1422]), .B(init), .Z(\round_in[0][1422] ) );
  AND U8188 ( .A(round_reg[1423]), .B(init), .Z(\round_in[0][1423] ) );
  AND U8189 ( .A(round_reg[1424]), .B(init), .Z(\round_in[0][1424] ) );
  AND U8190 ( .A(round_reg[1425]), .B(init), .Z(\round_in[0][1425] ) );
  AND U8191 ( .A(round_reg[1426]), .B(init), .Z(\round_in[0][1426] ) );
  AND U8192 ( .A(round_reg[1427]), .B(init), .Z(\round_in[0][1427] ) );
  AND U8193 ( .A(round_reg[1428]), .B(init), .Z(\round_in[0][1428] ) );
  AND U8194 ( .A(round_reg[1429]), .B(init), .Z(\round_in[0][1429] ) );
  NAND U8195 ( .A(init), .B(round_reg[142]), .Z(n2860) );
  NANDN U8196 ( .A(init), .B(in[142]), .Z(n2859) );
  NAND U8197 ( .A(n2860), .B(n2859), .Z(\round_in[0][142] ) );
  AND U8198 ( .A(round_reg[1430]), .B(init), .Z(\round_in[0][1430] ) );
  AND U8199 ( .A(round_reg[1431]), .B(init), .Z(\round_in[0][1431] ) );
  AND U8200 ( .A(round_reg[1432]), .B(init), .Z(\round_in[0][1432] ) );
  AND U8201 ( .A(round_reg[1433]), .B(init), .Z(\round_in[0][1433] ) );
  AND U8202 ( .A(round_reg[1434]), .B(init), .Z(\round_in[0][1434] ) );
  AND U8203 ( .A(round_reg[1435]), .B(init), .Z(\round_in[0][1435] ) );
  AND U8204 ( .A(round_reg[1436]), .B(init), .Z(\round_in[0][1436] ) );
  AND U8205 ( .A(round_reg[1437]), .B(init), .Z(\round_in[0][1437] ) );
  AND U8206 ( .A(round_reg[1438]), .B(init), .Z(\round_in[0][1438] ) );
  AND U8207 ( .A(round_reg[1439]), .B(init), .Z(\round_in[0][1439] ) );
  NAND U8208 ( .A(init), .B(round_reg[143]), .Z(n2862) );
  NANDN U8209 ( .A(init), .B(in[143]), .Z(n2861) );
  NAND U8210 ( .A(n2862), .B(n2861), .Z(\round_in[0][143] ) );
  AND U8211 ( .A(round_reg[1440]), .B(init), .Z(\round_in[0][1440] ) );
  AND U8212 ( .A(round_reg[1441]), .B(init), .Z(\round_in[0][1441] ) );
  AND U8213 ( .A(round_reg[1442]), .B(init), .Z(\round_in[0][1442] ) );
  AND U8214 ( .A(round_reg[1443]), .B(init), .Z(\round_in[0][1443] ) );
  AND U8215 ( .A(round_reg[1444]), .B(init), .Z(\round_in[0][1444] ) );
  AND U8216 ( .A(round_reg[1445]), .B(init), .Z(\round_in[0][1445] ) );
  AND U8217 ( .A(round_reg[1446]), .B(init), .Z(\round_in[0][1446] ) );
  AND U8218 ( .A(round_reg[1447]), .B(init), .Z(\round_in[0][1447] ) );
  AND U8219 ( .A(round_reg[1448]), .B(init), .Z(\round_in[0][1448] ) );
  AND U8220 ( .A(round_reg[1449]), .B(init), .Z(\round_in[0][1449] ) );
  NAND U8221 ( .A(init), .B(round_reg[144]), .Z(n2864) );
  NANDN U8222 ( .A(init), .B(in[144]), .Z(n2863) );
  NAND U8223 ( .A(n2864), .B(n2863), .Z(\round_in[0][144] ) );
  AND U8224 ( .A(round_reg[1450]), .B(init), .Z(\round_in[0][1450] ) );
  AND U8225 ( .A(round_reg[1451]), .B(init), .Z(\round_in[0][1451] ) );
  AND U8226 ( .A(round_reg[1452]), .B(init), .Z(\round_in[0][1452] ) );
  AND U8227 ( .A(round_reg[1453]), .B(init), .Z(\round_in[0][1453] ) );
  AND U8228 ( .A(round_reg[1454]), .B(init), .Z(\round_in[0][1454] ) );
  AND U8229 ( .A(round_reg[1455]), .B(init), .Z(\round_in[0][1455] ) );
  AND U8230 ( .A(round_reg[1456]), .B(init), .Z(\round_in[0][1456] ) );
  AND U8231 ( .A(round_reg[1457]), .B(init), .Z(\round_in[0][1457] ) );
  AND U8232 ( .A(round_reg[1458]), .B(init), .Z(\round_in[0][1458] ) );
  AND U8233 ( .A(round_reg[1459]), .B(init), .Z(\round_in[0][1459] ) );
  NAND U8234 ( .A(init), .B(round_reg[145]), .Z(n2866) );
  NANDN U8235 ( .A(init), .B(in[145]), .Z(n2865) );
  NAND U8236 ( .A(n2866), .B(n2865), .Z(\round_in[0][145] ) );
  AND U8237 ( .A(round_reg[1460]), .B(init), .Z(\round_in[0][1460] ) );
  AND U8238 ( .A(round_reg[1461]), .B(init), .Z(\round_in[0][1461] ) );
  AND U8239 ( .A(round_reg[1462]), .B(init), .Z(\round_in[0][1462] ) );
  AND U8240 ( .A(round_reg[1463]), .B(init), .Z(\round_in[0][1463] ) );
  AND U8241 ( .A(round_reg[1464]), .B(init), .Z(\round_in[0][1464] ) );
  AND U8242 ( .A(round_reg[1465]), .B(init), .Z(\round_in[0][1465] ) );
  AND U8243 ( .A(round_reg[1466]), .B(init), .Z(\round_in[0][1466] ) );
  AND U8244 ( .A(round_reg[1467]), .B(init), .Z(\round_in[0][1467] ) );
  AND U8245 ( .A(round_reg[1468]), .B(init), .Z(\round_in[0][1468] ) );
  AND U8246 ( .A(round_reg[1469]), .B(init), .Z(\round_in[0][1469] ) );
  NAND U8247 ( .A(init), .B(round_reg[146]), .Z(n2868) );
  NANDN U8248 ( .A(init), .B(in[146]), .Z(n2867) );
  NAND U8249 ( .A(n2868), .B(n2867), .Z(\round_in[0][146] ) );
  AND U8250 ( .A(round_reg[1470]), .B(init), .Z(\round_in[0][1470] ) );
  AND U8251 ( .A(round_reg[1471]), .B(init), .Z(\round_in[0][1471] ) );
  AND U8252 ( .A(round_reg[1472]), .B(init), .Z(\round_in[0][1472] ) );
  AND U8253 ( .A(round_reg[1473]), .B(init), .Z(\round_in[0][1473] ) );
  AND U8254 ( .A(round_reg[1474]), .B(init), .Z(\round_in[0][1474] ) );
  AND U8255 ( .A(round_reg[1475]), .B(init), .Z(\round_in[0][1475] ) );
  AND U8256 ( .A(round_reg[1476]), .B(init), .Z(\round_in[0][1476] ) );
  AND U8257 ( .A(round_reg[1477]), .B(init), .Z(\round_in[0][1477] ) );
  AND U8258 ( .A(round_reg[1478]), .B(init), .Z(\round_in[0][1478] ) );
  AND U8259 ( .A(round_reg[1479]), .B(init), .Z(\round_in[0][1479] ) );
  NAND U8260 ( .A(init), .B(round_reg[147]), .Z(n2870) );
  NANDN U8261 ( .A(init), .B(in[147]), .Z(n2869) );
  NAND U8262 ( .A(n2870), .B(n2869), .Z(\round_in[0][147] ) );
  AND U8263 ( .A(round_reg[1480]), .B(init), .Z(\round_in[0][1480] ) );
  AND U8264 ( .A(round_reg[1481]), .B(init), .Z(\round_in[0][1481] ) );
  AND U8265 ( .A(round_reg[1482]), .B(init), .Z(\round_in[0][1482] ) );
  AND U8266 ( .A(round_reg[1483]), .B(init), .Z(\round_in[0][1483] ) );
  AND U8267 ( .A(round_reg[1484]), .B(init), .Z(\round_in[0][1484] ) );
  AND U8268 ( .A(round_reg[1485]), .B(init), .Z(\round_in[0][1485] ) );
  AND U8269 ( .A(round_reg[1486]), .B(init), .Z(\round_in[0][1486] ) );
  AND U8270 ( .A(round_reg[1487]), .B(init), .Z(\round_in[0][1487] ) );
  AND U8271 ( .A(round_reg[1488]), .B(init), .Z(\round_in[0][1488] ) );
  AND U8272 ( .A(round_reg[1489]), .B(init), .Z(\round_in[0][1489] ) );
  NAND U8273 ( .A(init), .B(round_reg[148]), .Z(n2872) );
  NANDN U8274 ( .A(init), .B(in[148]), .Z(n2871) );
  NAND U8275 ( .A(n2872), .B(n2871), .Z(\round_in[0][148] ) );
  AND U8276 ( .A(round_reg[1490]), .B(init), .Z(\round_in[0][1490] ) );
  AND U8277 ( .A(round_reg[1491]), .B(init), .Z(\round_in[0][1491] ) );
  AND U8278 ( .A(round_reg[1492]), .B(init), .Z(\round_in[0][1492] ) );
  AND U8279 ( .A(round_reg[1493]), .B(init), .Z(\round_in[0][1493] ) );
  AND U8280 ( .A(round_reg[1494]), .B(init), .Z(\round_in[0][1494] ) );
  AND U8281 ( .A(round_reg[1495]), .B(init), .Z(\round_in[0][1495] ) );
  AND U8282 ( .A(round_reg[1496]), .B(init), .Z(\round_in[0][1496] ) );
  AND U8283 ( .A(round_reg[1497]), .B(init), .Z(\round_in[0][1497] ) );
  AND U8284 ( .A(round_reg[1498]), .B(init), .Z(\round_in[0][1498] ) );
  AND U8285 ( .A(round_reg[1499]), .B(init), .Z(\round_in[0][1499] ) );
  NAND U8286 ( .A(init), .B(round_reg[149]), .Z(n2874) );
  NANDN U8287 ( .A(init), .B(in[149]), .Z(n2873) );
  NAND U8288 ( .A(n2874), .B(n2873), .Z(\round_in[0][149] ) );
  NAND U8289 ( .A(init), .B(round_reg[14]), .Z(n2876) );
  NANDN U8290 ( .A(init), .B(in[14]), .Z(n2875) );
  NAND U8291 ( .A(n2876), .B(n2875), .Z(\round_in[0][14] ) );
  AND U8292 ( .A(round_reg[1500]), .B(init), .Z(\round_in[0][1500] ) );
  AND U8293 ( .A(round_reg[1501]), .B(init), .Z(\round_in[0][1501] ) );
  AND U8294 ( .A(round_reg[1502]), .B(init), .Z(\round_in[0][1502] ) );
  AND U8295 ( .A(round_reg[1503]), .B(init), .Z(\round_in[0][1503] ) );
  AND U8296 ( .A(round_reg[1504]), .B(init), .Z(\round_in[0][1504] ) );
  AND U8297 ( .A(round_reg[1505]), .B(init), .Z(\round_in[0][1505] ) );
  AND U8298 ( .A(round_reg[1506]), .B(init), .Z(\round_in[0][1506] ) );
  AND U8299 ( .A(round_reg[1507]), .B(init), .Z(\round_in[0][1507] ) );
  AND U8300 ( .A(round_reg[1508]), .B(init), .Z(\round_in[0][1508] ) );
  AND U8301 ( .A(round_reg[1509]), .B(init), .Z(\round_in[0][1509] ) );
  NAND U8302 ( .A(init), .B(round_reg[150]), .Z(n2878) );
  NANDN U8303 ( .A(init), .B(in[150]), .Z(n2877) );
  NAND U8304 ( .A(n2878), .B(n2877), .Z(\round_in[0][150] ) );
  AND U8305 ( .A(round_reg[1510]), .B(init), .Z(\round_in[0][1510] ) );
  AND U8306 ( .A(round_reg[1511]), .B(init), .Z(\round_in[0][1511] ) );
  AND U8307 ( .A(round_reg[1512]), .B(init), .Z(\round_in[0][1512] ) );
  AND U8308 ( .A(round_reg[1513]), .B(init), .Z(\round_in[0][1513] ) );
  AND U8309 ( .A(round_reg[1514]), .B(init), .Z(\round_in[0][1514] ) );
  AND U8310 ( .A(round_reg[1515]), .B(init), .Z(\round_in[0][1515] ) );
  AND U8311 ( .A(round_reg[1516]), .B(init), .Z(\round_in[0][1516] ) );
  AND U8312 ( .A(round_reg[1517]), .B(init), .Z(\round_in[0][1517] ) );
  AND U8313 ( .A(round_reg[1518]), .B(init), .Z(\round_in[0][1518] ) );
  AND U8314 ( .A(round_reg[1519]), .B(init), .Z(\round_in[0][1519] ) );
  NAND U8315 ( .A(init), .B(round_reg[151]), .Z(n2880) );
  NANDN U8316 ( .A(init), .B(in[151]), .Z(n2879) );
  NAND U8317 ( .A(n2880), .B(n2879), .Z(\round_in[0][151] ) );
  AND U8318 ( .A(round_reg[1520]), .B(init), .Z(\round_in[0][1520] ) );
  AND U8319 ( .A(round_reg[1521]), .B(init), .Z(\round_in[0][1521] ) );
  AND U8320 ( .A(round_reg[1522]), .B(init), .Z(\round_in[0][1522] ) );
  AND U8321 ( .A(round_reg[1523]), .B(init), .Z(\round_in[0][1523] ) );
  AND U8322 ( .A(round_reg[1524]), .B(init), .Z(\round_in[0][1524] ) );
  AND U8323 ( .A(round_reg[1525]), .B(init), .Z(\round_in[0][1525] ) );
  AND U8324 ( .A(round_reg[1526]), .B(init), .Z(\round_in[0][1526] ) );
  AND U8325 ( .A(round_reg[1527]), .B(init), .Z(\round_in[0][1527] ) );
  AND U8326 ( .A(round_reg[1528]), .B(init), .Z(\round_in[0][1528] ) );
  AND U8327 ( .A(round_reg[1529]), .B(init), .Z(\round_in[0][1529] ) );
  NAND U8328 ( .A(init), .B(round_reg[152]), .Z(n2882) );
  NANDN U8329 ( .A(init), .B(in[152]), .Z(n2881) );
  NAND U8330 ( .A(n2882), .B(n2881), .Z(\round_in[0][152] ) );
  AND U8331 ( .A(round_reg[1530]), .B(init), .Z(\round_in[0][1530] ) );
  AND U8332 ( .A(round_reg[1531]), .B(init), .Z(\round_in[0][1531] ) );
  AND U8333 ( .A(round_reg[1532]), .B(init), .Z(\round_in[0][1532] ) );
  AND U8334 ( .A(round_reg[1533]), .B(init), .Z(\round_in[0][1533] ) );
  AND U8335 ( .A(round_reg[1534]), .B(init), .Z(\round_in[0][1534] ) );
  AND U8336 ( .A(round_reg[1535]), .B(init), .Z(\round_in[0][1535] ) );
  AND U8337 ( .A(round_reg[1536]), .B(init), .Z(\round_in[0][1536] ) );
  AND U8338 ( .A(round_reg[1537]), .B(init), .Z(\round_in[0][1537] ) );
  AND U8339 ( .A(round_reg[1538]), .B(init), .Z(\round_in[0][1538] ) );
  AND U8340 ( .A(round_reg[1539]), .B(init), .Z(\round_in[0][1539] ) );
  NAND U8341 ( .A(init), .B(round_reg[153]), .Z(n2884) );
  NANDN U8342 ( .A(init), .B(in[153]), .Z(n2883) );
  NAND U8343 ( .A(n2884), .B(n2883), .Z(\round_in[0][153] ) );
  AND U8344 ( .A(round_reg[1540]), .B(init), .Z(\round_in[0][1540] ) );
  AND U8345 ( .A(round_reg[1541]), .B(init), .Z(\round_in[0][1541] ) );
  AND U8346 ( .A(round_reg[1542]), .B(init), .Z(\round_in[0][1542] ) );
  AND U8347 ( .A(round_reg[1543]), .B(init), .Z(\round_in[0][1543] ) );
  AND U8348 ( .A(round_reg[1544]), .B(init), .Z(\round_in[0][1544] ) );
  AND U8349 ( .A(round_reg[1545]), .B(init), .Z(\round_in[0][1545] ) );
  AND U8350 ( .A(round_reg[1546]), .B(init), .Z(\round_in[0][1546] ) );
  AND U8351 ( .A(round_reg[1547]), .B(init), .Z(\round_in[0][1547] ) );
  AND U8352 ( .A(round_reg[1548]), .B(init), .Z(\round_in[0][1548] ) );
  AND U8353 ( .A(round_reg[1549]), .B(init), .Z(\round_in[0][1549] ) );
  NAND U8354 ( .A(init), .B(round_reg[154]), .Z(n2886) );
  NANDN U8355 ( .A(init), .B(in[154]), .Z(n2885) );
  NAND U8356 ( .A(n2886), .B(n2885), .Z(\round_in[0][154] ) );
  AND U8357 ( .A(round_reg[1550]), .B(init), .Z(\round_in[0][1550] ) );
  AND U8358 ( .A(round_reg[1551]), .B(init), .Z(\round_in[0][1551] ) );
  AND U8359 ( .A(round_reg[1552]), .B(init), .Z(\round_in[0][1552] ) );
  AND U8360 ( .A(round_reg[1553]), .B(init), .Z(\round_in[0][1553] ) );
  AND U8361 ( .A(round_reg[1554]), .B(init), .Z(\round_in[0][1554] ) );
  AND U8362 ( .A(round_reg[1555]), .B(init), .Z(\round_in[0][1555] ) );
  AND U8363 ( .A(round_reg[1556]), .B(init), .Z(\round_in[0][1556] ) );
  AND U8364 ( .A(round_reg[1557]), .B(init), .Z(\round_in[0][1557] ) );
  AND U8365 ( .A(round_reg[1558]), .B(init), .Z(\round_in[0][1558] ) );
  AND U8366 ( .A(round_reg[1559]), .B(init), .Z(\round_in[0][1559] ) );
  NAND U8367 ( .A(init), .B(round_reg[155]), .Z(n2888) );
  NANDN U8368 ( .A(init), .B(in[155]), .Z(n2887) );
  NAND U8369 ( .A(n2888), .B(n2887), .Z(\round_in[0][155] ) );
  AND U8370 ( .A(round_reg[1560]), .B(init), .Z(\round_in[0][1560] ) );
  AND U8371 ( .A(round_reg[1561]), .B(init), .Z(\round_in[0][1561] ) );
  AND U8372 ( .A(round_reg[1562]), .B(init), .Z(\round_in[0][1562] ) );
  AND U8373 ( .A(round_reg[1563]), .B(init), .Z(\round_in[0][1563] ) );
  AND U8374 ( .A(round_reg[1564]), .B(init), .Z(\round_in[0][1564] ) );
  AND U8375 ( .A(round_reg[1565]), .B(init), .Z(\round_in[0][1565] ) );
  AND U8376 ( .A(round_reg[1566]), .B(init), .Z(\round_in[0][1566] ) );
  AND U8377 ( .A(round_reg[1567]), .B(init), .Z(\round_in[0][1567] ) );
  AND U8378 ( .A(round_reg[1568]), .B(init), .Z(\round_in[0][1568] ) );
  AND U8379 ( .A(round_reg[1569]), .B(init), .Z(\round_in[0][1569] ) );
  NAND U8380 ( .A(init), .B(round_reg[156]), .Z(n2890) );
  NANDN U8381 ( .A(init), .B(in[156]), .Z(n2889) );
  NAND U8382 ( .A(n2890), .B(n2889), .Z(\round_in[0][156] ) );
  AND U8383 ( .A(round_reg[1570]), .B(init), .Z(\round_in[0][1570] ) );
  AND U8384 ( .A(round_reg[1571]), .B(init), .Z(\round_in[0][1571] ) );
  AND U8385 ( .A(round_reg[1572]), .B(init), .Z(\round_in[0][1572] ) );
  AND U8386 ( .A(round_reg[1573]), .B(init), .Z(\round_in[0][1573] ) );
  AND U8387 ( .A(round_reg[1574]), .B(init), .Z(\round_in[0][1574] ) );
  AND U8388 ( .A(round_reg[1575]), .B(init), .Z(\round_in[0][1575] ) );
  AND U8389 ( .A(round_reg[1576]), .B(init), .Z(\round_in[0][1576] ) );
  AND U8390 ( .A(round_reg[1577]), .B(init), .Z(\round_in[0][1577] ) );
  AND U8391 ( .A(round_reg[1578]), .B(init), .Z(\round_in[0][1578] ) );
  AND U8392 ( .A(round_reg[1579]), .B(init), .Z(\round_in[0][1579] ) );
  NAND U8393 ( .A(init), .B(round_reg[157]), .Z(n2892) );
  NANDN U8394 ( .A(init), .B(in[157]), .Z(n2891) );
  NAND U8395 ( .A(n2892), .B(n2891), .Z(\round_in[0][157] ) );
  AND U8396 ( .A(round_reg[1580]), .B(init), .Z(\round_in[0][1580] ) );
  AND U8397 ( .A(round_reg[1581]), .B(init), .Z(\round_in[0][1581] ) );
  AND U8398 ( .A(round_reg[1582]), .B(init), .Z(\round_in[0][1582] ) );
  AND U8399 ( .A(round_reg[1583]), .B(init), .Z(\round_in[0][1583] ) );
  AND U8400 ( .A(round_reg[1584]), .B(init), .Z(\round_in[0][1584] ) );
  AND U8401 ( .A(round_reg[1585]), .B(init), .Z(\round_in[0][1585] ) );
  AND U8402 ( .A(round_reg[1586]), .B(init), .Z(\round_in[0][1586] ) );
  AND U8403 ( .A(round_reg[1587]), .B(init), .Z(\round_in[0][1587] ) );
  AND U8404 ( .A(round_reg[1588]), .B(init), .Z(\round_in[0][1588] ) );
  AND U8405 ( .A(round_reg[1589]), .B(init), .Z(\round_in[0][1589] ) );
  NAND U8406 ( .A(init), .B(round_reg[158]), .Z(n2894) );
  NANDN U8407 ( .A(init), .B(in[158]), .Z(n2893) );
  NAND U8408 ( .A(n2894), .B(n2893), .Z(\round_in[0][158] ) );
  AND U8409 ( .A(round_reg[1590]), .B(init), .Z(\round_in[0][1590] ) );
  AND U8410 ( .A(round_reg[1591]), .B(init), .Z(\round_in[0][1591] ) );
  AND U8411 ( .A(round_reg[1592]), .B(init), .Z(\round_in[0][1592] ) );
  AND U8412 ( .A(round_reg[1593]), .B(init), .Z(\round_in[0][1593] ) );
  AND U8413 ( .A(round_reg[1594]), .B(init), .Z(\round_in[0][1594] ) );
  AND U8414 ( .A(round_reg[1595]), .B(init), .Z(\round_in[0][1595] ) );
  AND U8415 ( .A(round_reg[1596]), .B(init), .Z(\round_in[0][1596] ) );
  AND U8416 ( .A(round_reg[1597]), .B(init), .Z(\round_in[0][1597] ) );
  AND U8417 ( .A(round_reg[1598]), .B(init), .Z(\round_in[0][1598] ) );
  AND U8418 ( .A(round_reg[1599]), .B(init), .Z(\round_in[0][1599] ) );
  NAND U8419 ( .A(init), .B(round_reg[159]), .Z(n2896) );
  NANDN U8420 ( .A(init), .B(in[159]), .Z(n2895) );
  NAND U8421 ( .A(n2896), .B(n2895), .Z(\round_in[0][159] ) );
  NAND U8422 ( .A(init), .B(round_reg[15]), .Z(n2898) );
  NANDN U8423 ( .A(init), .B(in[15]), .Z(n2897) );
  NAND U8424 ( .A(n2898), .B(n2897), .Z(\round_in[0][15] ) );
  NAND U8425 ( .A(init), .B(round_reg[160]), .Z(n2900) );
  NANDN U8426 ( .A(init), .B(in[160]), .Z(n2899) );
  NAND U8427 ( .A(n2900), .B(n2899), .Z(\round_in[0][160] ) );
  NAND U8428 ( .A(init), .B(round_reg[161]), .Z(n2902) );
  NANDN U8429 ( .A(init), .B(in[161]), .Z(n2901) );
  NAND U8430 ( .A(n2902), .B(n2901), .Z(\round_in[0][161] ) );
  NAND U8431 ( .A(init), .B(round_reg[162]), .Z(n2904) );
  NANDN U8432 ( .A(init), .B(in[162]), .Z(n2903) );
  NAND U8433 ( .A(n2904), .B(n2903), .Z(\round_in[0][162] ) );
  NAND U8434 ( .A(init), .B(round_reg[163]), .Z(n2906) );
  NANDN U8435 ( .A(init), .B(in[163]), .Z(n2905) );
  NAND U8436 ( .A(n2906), .B(n2905), .Z(\round_in[0][163] ) );
  NAND U8437 ( .A(init), .B(round_reg[164]), .Z(n2908) );
  NANDN U8438 ( .A(init), .B(in[164]), .Z(n2907) );
  NAND U8439 ( .A(n2908), .B(n2907), .Z(\round_in[0][164] ) );
  NAND U8440 ( .A(init), .B(round_reg[165]), .Z(n2910) );
  NANDN U8441 ( .A(init), .B(in[165]), .Z(n2909) );
  NAND U8442 ( .A(n2910), .B(n2909), .Z(\round_in[0][165] ) );
  NAND U8443 ( .A(init), .B(round_reg[166]), .Z(n2912) );
  NANDN U8444 ( .A(init), .B(in[166]), .Z(n2911) );
  NAND U8445 ( .A(n2912), .B(n2911), .Z(\round_in[0][166] ) );
  NAND U8446 ( .A(init), .B(round_reg[167]), .Z(n2914) );
  NANDN U8447 ( .A(init), .B(in[167]), .Z(n2913) );
  NAND U8448 ( .A(n2914), .B(n2913), .Z(\round_in[0][167] ) );
  NAND U8449 ( .A(init), .B(round_reg[168]), .Z(n2916) );
  NANDN U8450 ( .A(init), .B(in[168]), .Z(n2915) );
  NAND U8451 ( .A(n2916), .B(n2915), .Z(\round_in[0][168] ) );
  NAND U8452 ( .A(init), .B(round_reg[169]), .Z(n2918) );
  NANDN U8453 ( .A(init), .B(in[169]), .Z(n2917) );
  NAND U8454 ( .A(n2918), .B(n2917), .Z(\round_in[0][169] ) );
  NAND U8455 ( .A(init), .B(round_reg[16]), .Z(n2920) );
  NANDN U8456 ( .A(init), .B(in[16]), .Z(n2919) );
  NAND U8457 ( .A(n2920), .B(n2919), .Z(\round_in[0][16] ) );
  NAND U8458 ( .A(init), .B(round_reg[170]), .Z(n2922) );
  NANDN U8459 ( .A(init), .B(in[170]), .Z(n2921) );
  NAND U8460 ( .A(n2922), .B(n2921), .Z(\round_in[0][170] ) );
  NAND U8461 ( .A(init), .B(round_reg[171]), .Z(n2924) );
  NANDN U8462 ( .A(init), .B(in[171]), .Z(n2923) );
  NAND U8463 ( .A(n2924), .B(n2923), .Z(\round_in[0][171] ) );
  NAND U8464 ( .A(init), .B(round_reg[172]), .Z(n2926) );
  NANDN U8465 ( .A(init), .B(in[172]), .Z(n2925) );
  NAND U8466 ( .A(n2926), .B(n2925), .Z(\round_in[0][172] ) );
  NAND U8467 ( .A(init), .B(round_reg[173]), .Z(n2928) );
  NANDN U8468 ( .A(init), .B(in[173]), .Z(n2927) );
  NAND U8469 ( .A(n2928), .B(n2927), .Z(\round_in[0][173] ) );
  NAND U8470 ( .A(init), .B(round_reg[174]), .Z(n2930) );
  NANDN U8471 ( .A(init), .B(in[174]), .Z(n2929) );
  NAND U8472 ( .A(n2930), .B(n2929), .Z(\round_in[0][174] ) );
  NAND U8473 ( .A(init), .B(round_reg[175]), .Z(n2932) );
  NANDN U8474 ( .A(init), .B(in[175]), .Z(n2931) );
  NAND U8475 ( .A(n2932), .B(n2931), .Z(\round_in[0][175] ) );
  NAND U8476 ( .A(init), .B(round_reg[176]), .Z(n2934) );
  NANDN U8477 ( .A(init), .B(in[176]), .Z(n2933) );
  NAND U8478 ( .A(n2934), .B(n2933), .Z(\round_in[0][176] ) );
  NAND U8479 ( .A(init), .B(round_reg[177]), .Z(n2936) );
  NANDN U8480 ( .A(init), .B(in[177]), .Z(n2935) );
  NAND U8481 ( .A(n2936), .B(n2935), .Z(\round_in[0][177] ) );
  NAND U8482 ( .A(init), .B(round_reg[178]), .Z(n2938) );
  NANDN U8483 ( .A(init), .B(in[178]), .Z(n2937) );
  NAND U8484 ( .A(n2938), .B(n2937), .Z(\round_in[0][178] ) );
  NAND U8485 ( .A(init), .B(round_reg[179]), .Z(n2940) );
  NANDN U8486 ( .A(init), .B(in[179]), .Z(n2939) );
  NAND U8487 ( .A(n2940), .B(n2939), .Z(\round_in[0][179] ) );
  NAND U8488 ( .A(init), .B(round_reg[17]), .Z(n2942) );
  NANDN U8489 ( .A(init), .B(in[17]), .Z(n2941) );
  NAND U8490 ( .A(n2942), .B(n2941), .Z(\round_in[0][17] ) );
  NAND U8491 ( .A(init), .B(round_reg[180]), .Z(n2944) );
  NANDN U8492 ( .A(init), .B(in[180]), .Z(n2943) );
  NAND U8493 ( .A(n2944), .B(n2943), .Z(\round_in[0][180] ) );
  NAND U8494 ( .A(init), .B(round_reg[181]), .Z(n2946) );
  NANDN U8495 ( .A(init), .B(in[181]), .Z(n2945) );
  NAND U8496 ( .A(n2946), .B(n2945), .Z(\round_in[0][181] ) );
  NAND U8497 ( .A(init), .B(round_reg[182]), .Z(n2948) );
  NANDN U8498 ( .A(init), .B(in[182]), .Z(n2947) );
  NAND U8499 ( .A(n2948), .B(n2947), .Z(\round_in[0][182] ) );
  NAND U8500 ( .A(init), .B(round_reg[183]), .Z(n2950) );
  NANDN U8501 ( .A(init), .B(in[183]), .Z(n2949) );
  NAND U8502 ( .A(n2950), .B(n2949), .Z(\round_in[0][183] ) );
  NAND U8503 ( .A(init), .B(round_reg[184]), .Z(n2952) );
  NANDN U8504 ( .A(init), .B(in[184]), .Z(n2951) );
  NAND U8505 ( .A(n2952), .B(n2951), .Z(\round_in[0][184] ) );
  NAND U8506 ( .A(init), .B(round_reg[185]), .Z(n2954) );
  NANDN U8507 ( .A(init), .B(in[185]), .Z(n2953) );
  NAND U8508 ( .A(n2954), .B(n2953), .Z(\round_in[0][185] ) );
  NAND U8509 ( .A(init), .B(round_reg[186]), .Z(n2956) );
  NANDN U8510 ( .A(init), .B(in[186]), .Z(n2955) );
  NAND U8511 ( .A(n2956), .B(n2955), .Z(\round_in[0][186] ) );
  NAND U8512 ( .A(init), .B(round_reg[187]), .Z(n2958) );
  NANDN U8513 ( .A(init), .B(in[187]), .Z(n2957) );
  NAND U8514 ( .A(n2958), .B(n2957), .Z(\round_in[0][187] ) );
  NAND U8515 ( .A(init), .B(round_reg[188]), .Z(n2960) );
  NANDN U8516 ( .A(init), .B(in[188]), .Z(n2959) );
  NAND U8517 ( .A(n2960), .B(n2959), .Z(\round_in[0][188] ) );
  NAND U8518 ( .A(init), .B(round_reg[189]), .Z(n2962) );
  NANDN U8519 ( .A(init), .B(in[189]), .Z(n2961) );
  NAND U8520 ( .A(n2962), .B(n2961), .Z(\round_in[0][189] ) );
  NAND U8521 ( .A(init), .B(round_reg[18]), .Z(n2964) );
  NANDN U8522 ( .A(init), .B(in[18]), .Z(n2963) );
  NAND U8523 ( .A(n2964), .B(n2963), .Z(\round_in[0][18] ) );
  NAND U8524 ( .A(init), .B(round_reg[190]), .Z(n2966) );
  NANDN U8525 ( .A(init), .B(in[190]), .Z(n2965) );
  NAND U8526 ( .A(n2966), .B(n2965), .Z(\round_in[0][190] ) );
  NAND U8527 ( .A(init), .B(round_reg[191]), .Z(n2968) );
  NANDN U8528 ( .A(init), .B(in[191]), .Z(n2967) );
  NAND U8529 ( .A(n2968), .B(n2967), .Z(\round_in[0][191] ) );
  NAND U8530 ( .A(init), .B(round_reg[192]), .Z(n2970) );
  NANDN U8531 ( .A(init), .B(in[192]), .Z(n2969) );
  NAND U8532 ( .A(n2970), .B(n2969), .Z(\round_in[0][192] ) );
  NAND U8533 ( .A(init), .B(round_reg[193]), .Z(n2972) );
  NANDN U8534 ( .A(init), .B(in[193]), .Z(n2971) );
  NAND U8535 ( .A(n2972), .B(n2971), .Z(\round_in[0][193] ) );
  NAND U8536 ( .A(init), .B(round_reg[194]), .Z(n2974) );
  NANDN U8537 ( .A(init), .B(in[194]), .Z(n2973) );
  NAND U8538 ( .A(n2974), .B(n2973), .Z(\round_in[0][194] ) );
  NAND U8539 ( .A(init), .B(round_reg[195]), .Z(n2976) );
  NANDN U8540 ( .A(init), .B(in[195]), .Z(n2975) );
  NAND U8541 ( .A(n2976), .B(n2975), .Z(\round_in[0][195] ) );
  NAND U8542 ( .A(init), .B(round_reg[196]), .Z(n2978) );
  NANDN U8543 ( .A(init), .B(in[196]), .Z(n2977) );
  NAND U8544 ( .A(n2978), .B(n2977), .Z(\round_in[0][196] ) );
  NAND U8545 ( .A(init), .B(round_reg[197]), .Z(n2980) );
  NANDN U8546 ( .A(init), .B(in[197]), .Z(n2979) );
  NAND U8547 ( .A(n2980), .B(n2979), .Z(\round_in[0][197] ) );
  NAND U8548 ( .A(init), .B(round_reg[198]), .Z(n2982) );
  NANDN U8549 ( .A(init), .B(in[198]), .Z(n2981) );
  NAND U8550 ( .A(n2982), .B(n2981), .Z(\round_in[0][198] ) );
  NAND U8551 ( .A(init), .B(round_reg[199]), .Z(n2984) );
  NANDN U8552 ( .A(init), .B(in[199]), .Z(n2983) );
  NAND U8553 ( .A(n2984), .B(n2983), .Z(\round_in[0][199] ) );
  NAND U8554 ( .A(init), .B(round_reg[19]), .Z(n2986) );
  NANDN U8555 ( .A(init), .B(in[19]), .Z(n2985) );
  NAND U8556 ( .A(n2986), .B(n2985), .Z(\round_in[0][19] ) );
  NAND U8557 ( .A(init), .B(round_reg[1]), .Z(n2988) );
  NANDN U8558 ( .A(init), .B(in[1]), .Z(n2987) );
  NAND U8559 ( .A(n2988), .B(n2987), .Z(\round_in[0][1] ) );
  NAND U8560 ( .A(init), .B(round_reg[200]), .Z(n2990) );
  NANDN U8561 ( .A(init), .B(in[200]), .Z(n2989) );
  NAND U8562 ( .A(n2990), .B(n2989), .Z(\round_in[0][200] ) );
  NAND U8563 ( .A(init), .B(round_reg[201]), .Z(n2992) );
  NANDN U8564 ( .A(init), .B(in[201]), .Z(n2991) );
  NAND U8565 ( .A(n2992), .B(n2991), .Z(\round_in[0][201] ) );
  NAND U8566 ( .A(init), .B(round_reg[202]), .Z(n2994) );
  NANDN U8567 ( .A(init), .B(in[202]), .Z(n2993) );
  NAND U8568 ( .A(n2994), .B(n2993), .Z(\round_in[0][202] ) );
  NAND U8569 ( .A(init), .B(round_reg[203]), .Z(n2996) );
  NANDN U8570 ( .A(init), .B(in[203]), .Z(n2995) );
  NAND U8571 ( .A(n2996), .B(n2995), .Z(\round_in[0][203] ) );
  NAND U8572 ( .A(init), .B(round_reg[204]), .Z(n2998) );
  NANDN U8573 ( .A(init), .B(in[204]), .Z(n2997) );
  NAND U8574 ( .A(n2998), .B(n2997), .Z(\round_in[0][204] ) );
  NAND U8575 ( .A(init), .B(round_reg[205]), .Z(n3000) );
  NANDN U8576 ( .A(init), .B(in[205]), .Z(n2999) );
  NAND U8577 ( .A(n3000), .B(n2999), .Z(\round_in[0][205] ) );
  NAND U8578 ( .A(init), .B(round_reg[206]), .Z(n3002) );
  NANDN U8579 ( .A(init), .B(in[206]), .Z(n3001) );
  NAND U8580 ( .A(n3002), .B(n3001), .Z(\round_in[0][206] ) );
  NAND U8581 ( .A(init), .B(round_reg[207]), .Z(n3004) );
  NANDN U8582 ( .A(init), .B(in[207]), .Z(n3003) );
  NAND U8583 ( .A(n3004), .B(n3003), .Z(\round_in[0][207] ) );
  NAND U8584 ( .A(init), .B(round_reg[208]), .Z(n3006) );
  NANDN U8585 ( .A(init), .B(in[208]), .Z(n3005) );
  NAND U8586 ( .A(n3006), .B(n3005), .Z(\round_in[0][208] ) );
  NAND U8587 ( .A(init), .B(round_reg[209]), .Z(n3008) );
  NANDN U8588 ( .A(init), .B(in[209]), .Z(n3007) );
  NAND U8589 ( .A(n3008), .B(n3007), .Z(\round_in[0][209] ) );
  NAND U8590 ( .A(init), .B(round_reg[20]), .Z(n3010) );
  NANDN U8591 ( .A(init), .B(in[20]), .Z(n3009) );
  NAND U8592 ( .A(n3010), .B(n3009), .Z(\round_in[0][20] ) );
  NAND U8593 ( .A(init), .B(round_reg[210]), .Z(n3012) );
  NANDN U8594 ( .A(init), .B(in[210]), .Z(n3011) );
  NAND U8595 ( .A(n3012), .B(n3011), .Z(\round_in[0][210] ) );
  NAND U8596 ( .A(init), .B(round_reg[211]), .Z(n3014) );
  NANDN U8597 ( .A(init), .B(in[211]), .Z(n3013) );
  NAND U8598 ( .A(n3014), .B(n3013), .Z(\round_in[0][211] ) );
  NAND U8599 ( .A(init), .B(round_reg[212]), .Z(n3016) );
  NANDN U8600 ( .A(init), .B(in[212]), .Z(n3015) );
  NAND U8601 ( .A(n3016), .B(n3015), .Z(\round_in[0][212] ) );
  NAND U8602 ( .A(init), .B(round_reg[213]), .Z(n3018) );
  NANDN U8603 ( .A(init), .B(in[213]), .Z(n3017) );
  NAND U8604 ( .A(n3018), .B(n3017), .Z(\round_in[0][213] ) );
  NAND U8605 ( .A(init), .B(round_reg[214]), .Z(n3020) );
  NANDN U8606 ( .A(init), .B(in[214]), .Z(n3019) );
  NAND U8607 ( .A(n3020), .B(n3019), .Z(\round_in[0][214] ) );
  NAND U8608 ( .A(init), .B(round_reg[215]), .Z(n3022) );
  NANDN U8609 ( .A(init), .B(in[215]), .Z(n3021) );
  NAND U8610 ( .A(n3022), .B(n3021), .Z(\round_in[0][215] ) );
  NAND U8611 ( .A(init), .B(round_reg[216]), .Z(n3024) );
  NANDN U8612 ( .A(init), .B(in[216]), .Z(n3023) );
  NAND U8613 ( .A(n3024), .B(n3023), .Z(\round_in[0][216] ) );
  NAND U8614 ( .A(init), .B(round_reg[217]), .Z(n3026) );
  NANDN U8615 ( .A(init), .B(in[217]), .Z(n3025) );
  NAND U8616 ( .A(n3026), .B(n3025), .Z(\round_in[0][217] ) );
  NAND U8617 ( .A(init), .B(round_reg[218]), .Z(n3028) );
  NANDN U8618 ( .A(init), .B(in[218]), .Z(n3027) );
  NAND U8619 ( .A(n3028), .B(n3027), .Z(\round_in[0][218] ) );
  NAND U8620 ( .A(init), .B(round_reg[219]), .Z(n3030) );
  NANDN U8621 ( .A(init), .B(in[219]), .Z(n3029) );
  NAND U8622 ( .A(n3030), .B(n3029), .Z(\round_in[0][219] ) );
  NAND U8623 ( .A(init), .B(round_reg[21]), .Z(n3032) );
  NANDN U8624 ( .A(init), .B(in[21]), .Z(n3031) );
  NAND U8625 ( .A(n3032), .B(n3031), .Z(\round_in[0][21] ) );
  NAND U8626 ( .A(init), .B(round_reg[220]), .Z(n3034) );
  NANDN U8627 ( .A(init), .B(in[220]), .Z(n3033) );
  NAND U8628 ( .A(n3034), .B(n3033), .Z(\round_in[0][220] ) );
  NAND U8629 ( .A(init), .B(round_reg[221]), .Z(n3036) );
  NANDN U8630 ( .A(init), .B(in[221]), .Z(n3035) );
  NAND U8631 ( .A(n3036), .B(n3035), .Z(\round_in[0][221] ) );
  NAND U8632 ( .A(init), .B(round_reg[222]), .Z(n3038) );
  NANDN U8633 ( .A(init), .B(in[222]), .Z(n3037) );
  NAND U8634 ( .A(n3038), .B(n3037), .Z(\round_in[0][222] ) );
  NAND U8635 ( .A(init), .B(round_reg[223]), .Z(n3040) );
  NANDN U8636 ( .A(init), .B(in[223]), .Z(n3039) );
  NAND U8637 ( .A(n3040), .B(n3039), .Z(\round_in[0][223] ) );
  NAND U8638 ( .A(init), .B(round_reg[224]), .Z(n3042) );
  NANDN U8639 ( .A(init), .B(in[224]), .Z(n3041) );
  NAND U8640 ( .A(n3042), .B(n3041), .Z(\round_in[0][224] ) );
  NAND U8641 ( .A(init), .B(round_reg[225]), .Z(n3044) );
  NANDN U8642 ( .A(init), .B(in[225]), .Z(n3043) );
  NAND U8643 ( .A(n3044), .B(n3043), .Z(\round_in[0][225] ) );
  NAND U8644 ( .A(init), .B(round_reg[226]), .Z(n3046) );
  NANDN U8645 ( .A(init), .B(in[226]), .Z(n3045) );
  NAND U8646 ( .A(n3046), .B(n3045), .Z(\round_in[0][226] ) );
  NAND U8647 ( .A(init), .B(round_reg[227]), .Z(n3048) );
  NANDN U8648 ( .A(init), .B(in[227]), .Z(n3047) );
  NAND U8649 ( .A(n3048), .B(n3047), .Z(\round_in[0][227] ) );
  NAND U8650 ( .A(init), .B(round_reg[228]), .Z(n3050) );
  NANDN U8651 ( .A(init), .B(in[228]), .Z(n3049) );
  NAND U8652 ( .A(n3050), .B(n3049), .Z(\round_in[0][228] ) );
  NAND U8653 ( .A(init), .B(round_reg[229]), .Z(n3052) );
  NANDN U8654 ( .A(init), .B(in[229]), .Z(n3051) );
  NAND U8655 ( .A(n3052), .B(n3051), .Z(\round_in[0][229] ) );
  NAND U8656 ( .A(init), .B(round_reg[22]), .Z(n3054) );
  NANDN U8657 ( .A(init), .B(in[22]), .Z(n3053) );
  NAND U8658 ( .A(n3054), .B(n3053), .Z(\round_in[0][22] ) );
  NAND U8659 ( .A(init), .B(round_reg[230]), .Z(n3056) );
  NANDN U8660 ( .A(init), .B(in[230]), .Z(n3055) );
  NAND U8661 ( .A(n3056), .B(n3055), .Z(\round_in[0][230] ) );
  NAND U8662 ( .A(init), .B(round_reg[231]), .Z(n3058) );
  NANDN U8663 ( .A(init), .B(in[231]), .Z(n3057) );
  NAND U8664 ( .A(n3058), .B(n3057), .Z(\round_in[0][231] ) );
  NAND U8665 ( .A(init), .B(round_reg[232]), .Z(n3060) );
  NANDN U8666 ( .A(init), .B(in[232]), .Z(n3059) );
  NAND U8667 ( .A(n3060), .B(n3059), .Z(\round_in[0][232] ) );
  NAND U8668 ( .A(init), .B(round_reg[233]), .Z(n3062) );
  NANDN U8669 ( .A(init), .B(in[233]), .Z(n3061) );
  NAND U8670 ( .A(n3062), .B(n3061), .Z(\round_in[0][233] ) );
  NAND U8671 ( .A(init), .B(round_reg[234]), .Z(n3064) );
  NANDN U8672 ( .A(init), .B(in[234]), .Z(n3063) );
  NAND U8673 ( .A(n3064), .B(n3063), .Z(\round_in[0][234] ) );
  NAND U8674 ( .A(init), .B(round_reg[235]), .Z(n3066) );
  NANDN U8675 ( .A(init), .B(in[235]), .Z(n3065) );
  NAND U8676 ( .A(n3066), .B(n3065), .Z(\round_in[0][235] ) );
  NAND U8677 ( .A(init), .B(round_reg[236]), .Z(n3068) );
  NANDN U8678 ( .A(init), .B(in[236]), .Z(n3067) );
  NAND U8679 ( .A(n3068), .B(n3067), .Z(\round_in[0][236] ) );
  NAND U8680 ( .A(init), .B(round_reg[237]), .Z(n3070) );
  NANDN U8681 ( .A(init), .B(in[237]), .Z(n3069) );
  NAND U8682 ( .A(n3070), .B(n3069), .Z(\round_in[0][237] ) );
  NAND U8683 ( .A(init), .B(round_reg[238]), .Z(n3072) );
  NANDN U8684 ( .A(init), .B(in[238]), .Z(n3071) );
  NAND U8685 ( .A(n3072), .B(n3071), .Z(\round_in[0][238] ) );
  NAND U8686 ( .A(init), .B(round_reg[239]), .Z(n3074) );
  NANDN U8687 ( .A(init), .B(in[239]), .Z(n3073) );
  NAND U8688 ( .A(n3074), .B(n3073), .Z(\round_in[0][239] ) );
  NAND U8689 ( .A(init), .B(round_reg[23]), .Z(n3076) );
  NANDN U8690 ( .A(init), .B(in[23]), .Z(n3075) );
  NAND U8691 ( .A(n3076), .B(n3075), .Z(\round_in[0][23] ) );
  NAND U8692 ( .A(init), .B(round_reg[240]), .Z(n3078) );
  NANDN U8693 ( .A(init), .B(in[240]), .Z(n3077) );
  NAND U8694 ( .A(n3078), .B(n3077), .Z(\round_in[0][240] ) );
  NAND U8695 ( .A(init), .B(round_reg[241]), .Z(n3080) );
  NANDN U8696 ( .A(init), .B(in[241]), .Z(n3079) );
  NAND U8697 ( .A(n3080), .B(n3079), .Z(\round_in[0][241] ) );
  NAND U8698 ( .A(init), .B(round_reg[242]), .Z(n3082) );
  NANDN U8699 ( .A(init), .B(in[242]), .Z(n3081) );
  NAND U8700 ( .A(n3082), .B(n3081), .Z(\round_in[0][242] ) );
  NAND U8701 ( .A(init), .B(round_reg[243]), .Z(n3084) );
  NANDN U8702 ( .A(init), .B(in[243]), .Z(n3083) );
  NAND U8703 ( .A(n3084), .B(n3083), .Z(\round_in[0][243] ) );
  NAND U8704 ( .A(init), .B(round_reg[244]), .Z(n3086) );
  NANDN U8705 ( .A(init), .B(in[244]), .Z(n3085) );
  NAND U8706 ( .A(n3086), .B(n3085), .Z(\round_in[0][244] ) );
  NAND U8707 ( .A(init), .B(round_reg[245]), .Z(n3088) );
  NANDN U8708 ( .A(init), .B(in[245]), .Z(n3087) );
  NAND U8709 ( .A(n3088), .B(n3087), .Z(\round_in[0][245] ) );
  NAND U8710 ( .A(init), .B(round_reg[246]), .Z(n3090) );
  NANDN U8711 ( .A(init), .B(in[246]), .Z(n3089) );
  NAND U8712 ( .A(n3090), .B(n3089), .Z(\round_in[0][246] ) );
  NAND U8713 ( .A(init), .B(round_reg[247]), .Z(n3092) );
  NANDN U8714 ( .A(init), .B(in[247]), .Z(n3091) );
  NAND U8715 ( .A(n3092), .B(n3091), .Z(\round_in[0][247] ) );
  NAND U8716 ( .A(init), .B(round_reg[248]), .Z(n3094) );
  NANDN U8717 ( .A(init), .B(in[248]), .Z(n3093) );
  NAND U8718 ( .A(n3094), .B(n3093), .Z(\round_in[0][248] ) );
  NAND U8719 ( .A(init), .B(round_reg[249]), .Z(n3096) );
  NANDN U8720 ( .A(init), .B(in[249]), .Z(n3095) );
  NAND U8721 ( .A(n3096), .B(n3095), .Z(\round_in[0][249] ) );
  NAND U8722 ( .A(init), .B(round_reg[24]), .Z(n3098) );
  NANDN U8723 ( .A(init), .B(in[24]), .Z(n3097) );
  NAND U8724 ( .A(n3098), .B(n3097), .Z(\round_in[0][24] ) );
  NAND U8725 ( .A(init), .B(round_reg[250]), .Z(n3100) );
  NANDN U8726 ( .A(init), .B(in[250]), .Z(n3099) );
  NAND U8727 ( .A(n3100), .B(n3099), .Z(\round_in[0][250] ) );
  NAND U8728 ( .A(init), .B(round_reg[251]), .Z(n3102) );
  NANDN U8729 ( .A(init), .B(in[251]), .Z(n3101) );
  NAND U8730 ( .A(n3102), .B(n3101), .Z(\round_in[0][251] ) );
  NAND U8731 ( .A(init), .B(round_reg[252]), .Z(n3104) );
  NANDN U8732 ( .A(init), .B(in[252]), .Z(n3103) );
  NAND U8733 ( .A(n3104), .B(n3103), .Z(\round_in[0][252] ) );
  NAND U8734 ( .A(init), .B(round_reg[253]), .Z(n3106) );
  NANDN U8735 ( .A(init), .B(in[253]), .Z(n3105) );
  NAND U8736 ( .A(n3106), .B(n3105), .Z(\round_in[0][253] ) );
  NAND U8737 ( .A(init), .B(round_reg[254]), .Z(n3108) );
  NANDN U8738 ( .A(init), .B(in[254]), .Z(n3107) );
  NAND U8739 ( .A(n3108), .B(n3107), .Z(\round_in[0][254] ) );
  NAND U8740 ( .A(init), .B(round_reg[255]), .Z(n3110) );
  NANDN U8741 ( .A(init), .B(in[255]), .Z(n3109) );
  NAND U8742 ( .A(n3110), .B(n3109), .Z(\round_in[0][255] ) );
  NAND U8743 ( .A(init), .B(round_reg[256]), .Z(n3112) );
  NANDN U8744 ( .A(init), .B(in[256]), .Z(n3111) );
  NAND U8745 ( .A(n3112), .B(n3111), .Z(\round_in[0][256] ) );
  NAND U8746 ( .A(init), .B(round_reg[257]), .Z(n3114) );
  NANDN U8747 ( .A(init), .B(in[257]), .Z(n3113) );
  NAND U8748 ( .A(n3114), .B(n3113), .Z(\round_in[0][257] ) );
  NAND U8749 ( .A(init), .B(round_reg[258]), .Z(n3116) );
  NANDN U8750 ( .A(init), .B(in[258]), .Z(n3115) );
  NAND U8751 ( .A(n3116), .B(n3115), .Z(\round_in[0][258] ) );
  NAND U8752 ( .A(init), .B(round_reg[259]), .Z(n3118) );
  NANDN U8753 ( .A(init), .B(in[259]), .Z(n3117) );
  NAND U8754 ( .A(n3118), .B(n3117), .Z(\round_in[0][259] ) );
  NAND U8755 ( .A(init), .B(round_reg[25]), .Z(n3120) );
  NANDN U8756 ( .A(init), .B(in[25]), .Z(n3119) );
  NAND U8757 ( .A(n3120), .B(n3119), .Z(\round_in[0][25] ) );
  NAND U8758 ( .A(init), .B(round_reg[260]), .Z(n3122) );
  NANDN U8759 ( .A(init), .B(in[260]), .Z(n3121) );
  NAND U8760 ( .A(n3122), .B(n3121), .Z(\round_in[0][260] ) );
  NAND U8761 ( .A(init), .B(round_reg[261]), .Z(n3124) );
  NANDN U8762 ( .A(init), .B(in[261]), .Z(n3123) );
  NAND U8763 ( .A(n3124), .B(n3123), .Z(\round_in[0][261] ) );
  NAND U8764 ( .A(init), .B(round_reg[262]), .Z(n3126) );
  NANDN U8765 ( .A(init), .B(in[262]), .Z(n3125) );
  NAND U8766 ( .A(n3126), .B(n3125), .Z(\round_in[0][262] ) );
  NAND U8767 ( .A(init), .B(round_reg[263]), .Z(n3128) );
  NANDN U8768 ( .A(init), .B(in[263]), .Z(n3127) );
  NAND U8769 ( .A(n3128), .B(n3127), .Z(\round_in[0][263] ) );
  NAND U8770 ( .A(init), .B(round_reg[264]), .Z(n3130) );
  NANDN U8771 ( .A(init), .B(in[264]), .Z(n3129) );
  NAND U8772 ( .A(n3130), .B(n3129), .Z(\round_in[0][264] ) );
  NAND U8773 ( .A(init), .B(round_reg[265]), .Z(n3132) );
  NANDN U8774 ( .A(init), .B(in[265]), .Z(n3131) );
  NAND U8775 ( .A(n3132), .B(n3131), .Z(\round_in[0][265] ) );
  NAND U8776 ( .A(init), .B(round_reg[266]), .Z(n3134) );
  NANDN U8777 ( .A(init), .B(in[266]), .Z(n3133) );
  NAND U8778 ( .A(n3134), .B(n3133), .Z(\round_in[0][266] ) );
  NAND U8779 ( .A(init), .B(round_reg[267]), .Z(n3136) );
  NANDN U8780 ( .A(init), .B(in[267]), .Z(n3135) );
  NAND U8781 ( .A(n3136), .B(n3135), .Z(\round_in[0][267] ) );
  NAND U8782 ( .A(init), .B(round_reg[268]), .Z(n3138) );
  NANDN U8783 ( .A(init), .B(in[268]), .Z(n3137) );
  NAND U8784 ( .A(n3138), .B(n3137), .Z(\round_in[0][268] ) );
  NAND U8785 ( .A(init), .B(round_reg[269]), .Z(n3140) );
  NANDN U8786 ( .A(init), .B(in[269]), .Z(n3139) );
  NAND U8787 ( .A(n3140), .B(n3139), .Z(\round_in[0][269] ) );
  NAND U8788 ( .A(init), .B(round_reg[26]), .Z(n3142) );
  NANDN U8789 ( .A(init), .B(in[26]), .Z(n3141) );
  NAND U8790 ( .A(n3142), .B(n3141), .Z(\round_in[0][26] ) );
  NAND U8791 ( .A(init), .B(round_reg[270]), .Z(n3144) );
  NANDN U8792 ( .A(init), .B(in[270]), .Z(n3143) );
  NAND U8793 ( .A(n3144), .B(n3143), .Z(\round_in[0][270] ) );
  NAND U8794 ( .A(init), .B(round_reg[271]), .Z(n3146) );
  NANDN U8795 ( .A(init), .B(in[271]), .Z(n3145) );
  NAND U8796 ( .A(n3146), .B(n3145), .Z(\round_in[0][271] ) );
  NAND U8797 ( .A(init), .B(round_reg[272]), .Z(n3148) );
  NANDN U8798 ( .A(init), .B(in[272]), .Z(n3147) );
  NAND U8799 ( .A(n3148), .B(n3147), .Z(\round_in[0][272] ) );
  NAND U8800 ( .A(init), .B(round_reg[273]), .Z(n3150) );
  NANDN U8801 ( .A(init), .B(in[273]), .Z(n3149) );
  NAND U8802 ( .A(n3150), .B(n3149), .Z(\round_in[0][273] ) );
  NAND U8803 ( .A(init), .B(round_reg[274]), .Z(n3152) );
  NANDN U8804 ( .A(init), .B(in[274]), .Z(n3151) );
  NAND U8805 ( .A(n3152), .B(n3151), .Z(\round_in[0][274] ) );
  NAND U8806 ( .A(init), .B(round_reg[275]), .Z(n3154) );
  NANDN U8807 ( .A(init), .B(in[275]), .Z(n3153) );
  NAND U8808 ( .A(n3154), .B(n3153), .Z(\round_in[0][275] ) );
  NAND U8809 ( .A(init), .B(round_reg[276]), .Z(n3156) );
  NANDN U8810 ( .A(init), .B(in[276]), .Z(n3155) );
  NAND U8811 ( .A(n3156), .B(n3155), .Z(\round_in[0][276] ) );
  NAND U8812 ( .A(init), .B(round_reg[277]), .Z(n3158) );
  NANDN U8813 ( .A(init), .B(in[277]), .Z(n3157) );
  NAND U8814 ( .A(n3158), .B(n3157), .Z(\round_in[0][277] ) );
  NAND U8815 ( .A(init), .B(round_reg[278]), .Z(n3160) );
  NANDN U8816 ( .A(init), .B(in[278]), .Z(n3159) );
  NAND U8817 ( .A(n3160), .B(n3159), .Z(\round_in[0][278] ) );
  NAND U8818 ( .A(init), .B(round_reg[279]), .Z(n3162) );
  NANDN U8819 ( .A(init), .B(in[279]), .Z(n3161) );
  NAND U8820 ( .A(n3162), .B(n3161), .Z(\round_in[0][279] ) );
  NAND U8821 ( .A(init), .B(round_reg[27]), .Z(n3164) );
  NANDN U8822 ( .A(init), .B(in[27]), .Z(n3163) );
  NAND U8823 ( .A(n3164), .B(n3163), .Z(\round_in[0][27] ) );
  NAND U8824 ( .A(init), .B(round_reg[280]), .Z(n3166) );
  NANDN U8825 ( .A(init), .B(in[280]), .Z(n3165) );
  NAND U8826 ( .A(n3166), .B(n3165), .Z(\round_in[0][280] ) );
  NAND U8827 ( .A(init), .B(round_reg[281]), .Z(n3168) );
  NANDN U8828 ( .A(init), .B(in[281]), .Z(n3167) );
  NAND U8829 ( .A(n3168), .B(n3167), .Z(\round_in[0][281] ) );
  NAND U8830 ( .A(init), .B(round_reg[282]), .Z(n3170) );
  NANDN U8831 ( .A(init), .B(in[282]), .Z(n3169) );
  NAND U8832 ( .A(n3170), .B(n3169), .Z(\round_in[0][282] ) );
  NAND U8833 ( .A(init), .B(round_reg[283]), .Z(n3172) );
  NANDN U8834 ( .A(init), .B(in[283]), .Z(n3171) );
  NAND U8835 ( .A(n3172), .B(n3171), .Z(\round_in[0][283] ) );
  NAND U8836 ( .A(init), .B(round_reg[284]), .Z(n3174) );
  NANDN U8837 ( .A(init), .B(in[284]), .Z(n3173) );
  NAND U8838 ( .A(n3174), .B(n3173), .Z(\round_in[0][284] ) );
  NAND U8839 ( .A(init), .B(round_reg[285]), .Z(n3176) );
  NANDN U8840 ( .A(init), .B(in[285]), .Z(n3175) );
  NAND U8841 ( .A(n3176), .B(n3175), .Z(\round_in[0][285] ) );
  NAND U8842 ( .A(init), .B(round_reg[286]), .Z(n3178) );
  NANDN U8843 ( .A(init), .B(in[286]), .Z(n3177) );
  NAND U8844 ( .A(n3178), .B(n3177), .Z(\round_in[0][286] ) );
  NAND U8845 ( .A(init), .B(round_reg[287]), .Z(n3180) );
  NANDN U8846 ( .A(init), .B(in[287]), .Z(n3179) );
  NAND U8847 ( .A(n3180), .B(n3179), .Z(\round_in[0][287] ) );
  NAND U8848 ( .A(init), .B(round_reg[288]), .Z(n3182) );
  NANDN U8849 ( .A(init), .B(in[288]), .Z(n3181) );
  NAND U8850 ( .A(n3182), .B(n3181), .Z(\round_in[0][288] ) );
  NAND U8851 ( .A(init), .B(round_reg[289]), .Z(n3184) );
  NANDN U8852 ( .A(init), .B(in[289]), .Z(n3183) );
  NAND U8853 ( .A(n3184), .B(n3183), .Z(\round_in[0][289] ) );
  NAND U8854 ( .A(init), .B(round_reg[28]), .Z(n3186) );
  NANDN U8855 ( .A(init), .B(in[28]), .Z(n3185) );
  NAND U8856 ( .A(n3186), .B(n3185), .Z(\round_in[0][28] ) );
  NAND U8857 ( .A(init), .B(round_reg[290]), .Z(n3188) );
  NANDN U8858 ( .A(init), .B(in[290]), .Z(n3187) );
  NAND U8859 ( .A(n3188), .B(n3187), .Z(\round_in[0][290] ) );
  NAND U8860 ( .A(init), .B(round_reg[291]), .Z(n3190) );
  NANDN U8861 ( .A(init), .B(in[291]), .Z(n3189) );
  NAND U8862 ( .A(n3190), .B(n3189), .Z(\round_in[0][291] ) );
  NAND U8863 ( .A(init), .B(round_reg[292]), .Z(n3192) );
  NANDN U8864 ( .A(init), .B(in[292]), .Z(n3191) );
  NAND U8865 ( .A(n3192), .B(n3191), .Z(\round_in[0][292] ) );
  NAND U8866 ( .A(init), .B(round_reg[293]), .Z(n3194) );
  NANDN U8867 ( .A(init), .B(in[293]), .Z(n3193) );
  NAND U8868 ( .A(n3194), .B(n3193), .Z(\round_in[0][293] ) );
  NAND U8869 ( .A(init), .B(round_reg[294]), .Z(n3196) );
  NANDN U8870 ( .A(init), .B(in[294]), .Z(n3195) );
  NAND U8871 ( .A(n3196), .B(n3195), .Z(\round_in[0][294] ) );
  NAND U8872 ( .A(init), .B(round_reg[295]), .Z(n3198) );
  NANDN U8873 ( .A(init), .B(in[295]), .Z(n3197) );
  NAND U8874 ( .A(n3198), .B(n3197), .Z(\round_in[0][295] ) );
  NAND U8875 ( .A(init), .B(round_reg[296]), .Z(n3200) );
  NANDN U8876 ( .A(init), .B(in[296]), .Z(n3199) );
  NAND U8877 ( .A(n3200), .B(n3199), .Z(\round_in[0][296] ) );
  NAND U8878 ( .A(init), .B(round_reg[297]), .Z(n3202) );
  NANDN U8879 ( .A(init), .B(in[297]), .Z(n3201) );
  NAND U8880 ( .A(n3202), .B(n3201), .Z(\round_in[0][297] ) );
  NAND U8881 ( .A(init), .B(round_reg[298]), .Z(n3204) );
  NANDN U8882 ( .A(init), .B(in[298]), .Z(n3203) );
  NAND U8883 ( .A(n3204), .B(n3203), .Z(\round_in[0][298] ) );
  NAND U8884 ( .A(init), .B(round_reg[299]), .Z(n3206) );
  NANDN U8885 ( .A(init), .B(in[299]), .Z(n3205) );
  NAND U8886 ( .A(n3206), .B(n3205), .Z(\round_in[0][299] ) );
  NAND U8887 ( .A(init), .B(round_reg[29]), .Z(n3208) );
  NANDN U8888 ( .A(init), .B(in[29]), .Z(n3207) );
  NAND U8889 ( .A(n3208), .B(n3207), .Z(\round_in[0][29] ) );
  NAND U8890 ( .A(init), .B(round_reg[2]), .Z(n3210) );
  NANDN U8891 ( .A(init), .B(in[2]), .Z(n3209) );
  NAND U8892 ( .A(n3210), .B(n3209), .Z(\round_in[0][2] ) );
  NAND U8893 ( .A(init), .B(round_reg[300]), .Z(n3212) );
  NANDN U8894 ( .A(init), .B(in[300]), .Z(n3211) );
  NAND U8895 ( .A(n3212), .B(n3211), .Z(\round_in[0][300] ) );
  NAND U8896 ( .A(init), .B(round_reg[301]), .Z(n3214) );
  NANDN U8897 ( .A(init), .B(in[301]), .Z(n3213) );
  NAND U8898 ( .A(n3214), .B(n3213), .Z(\round_in[0][301] ) );
  NAND U8899 ( .A(init), .B(round_reg[302]), .Z(n3216) );
  NANDN U8900 ( .A(init), .B(in[302]), .Z(n3215) );
  NAND U8901 ( .A(n3216), .B(n3215), .Z(\round_in[0][302] ) );
  NAND U8902 ( .A(init), .B(round_reg[303]), .Z(n3218) );
  NANDN U8903 ( .A(init), .B(in[303]), .Z(n3217) );
  NAND U8904 ( .A(n3218), .B(n3217), .Z(\round_in[0][303] ) );
  NAND U8905 ( .A(init), .B(round_reg[304]), .Z(n3220) );
  NANDN U8906 ( .A(init), .B(in[304]), .Z(n3219) );
  NAND U8907 ( .A(n3220), .B(n3219), .Z(\round_in[0][304] ) );
  NAND U8908 ( .A(init), .B(round_reg[305]), .Z(n3222) );
  NANDN U8909 ( .A(init), .B(in[305]), .Z(n3221) );
  NAND U8910 ( .A(n3222), .B(n3221), .Z(\round_in[0][305] ) );
  NAND U8911 ( .A(init), .B(round_reg[306]), .Z(n3224) );
  NANDN U8912 ( .A(init), .B(in[306]), .Z(n3223) );
  NAND U8913 ( .A(n3224), .B(n3223), .Z(\round_in[0][306] ) );
  NAND U8914 ( .A(init), .B(round_reg[307]), .Z(n3226) );
  NANDN U8915 ( .A(init), .B(in[307]), .Z(n3225) );
  NAND U8916 ( .A(n3226), .B(n3225), .Z(\round_in[0][307] ) );
  NAND U8917 ( .A(init), .B(round_reg[308]), .Z(n3228) );
  NANDN U8918 ( .A(init), .B(in[308]), .Z(n3227) );
  NAND U8919 ( .A(n3228), .B(n3227), .Z(\round_in[0][308] ) );
  NAND U8920 ( .A(init), .B(round_reg[309]), .Z(n3230) );
  NANDN U8921 ( .A(init), .B(in[309]), .Z(n3229) );
  NAND U8922 ( .A(n3230), .B(n3229), .Z(\round_in[0][309] ) );
  NAND U8923 ( .A(init), .B(round_reg[30]), .Z(n3232) );
  NANDN U8924 ( .A(init), .B(in[30]), .Z(n3231) );
  NAND U8925 ( .A(n3232), .B(n3231), .Z(\round_in[0][30] ) );
  NAND U8926 ( .A(init), .B(round_reg[310]), .Z(n3234) );
  NANDN U8927 ( .A(init), .B(in[310]), .Z(n3233) );
  NAND U8928 ( .A(n3234), .B(n3233), .Z(\round_in[0][310] ) );
  NAND U8929 ( .A(init), .B(round_reg[311]), .Z(n3236) );
  NANDN U8930 ( .A(init), .B(in[311]), .Z(n3235) );
  NAND U8931 ( .A(n3236), .B(n3235), .Z(\round_in[0][311] ) );
  NAND U8932 ( .A(init), .B(round_reg[312]), .Z(n3238) );
  NANDN U8933 ( .A(init), .B(in[312]), .Z(n3237) );
  NAND U8934 ( .A(n3238), .B(n3237), .Z(\round_in[0][312] ) );
  NAND U8935 ( .A(init), .B(round_reg[313]), .Z(n3240) );
  NANDN U8936 ( .A(init), .B(in[313]), .Z(n3239) );
  NAND U8937 ( .A(n3240), .B(n3239), .Z(\round_in[0][313] ) );
  NAND U8938 ( .A(init), .B(round_reg[314]), .Z(n3242) );
  NANDN U8939 ( .A(init), .B(in[314]), .Z(n3241) );
  NAND U8940 ( .A(n3242), .B(n3241), .Z(\round_in[0][314] ) );
  NAND U8941 ( .A(init), .B(round_reg[315]), .Z(n3244) );
  NANDN U8942 ( .A(init), .B(in[315]), .Z(n3243) );
  NAND U8943 ( .A(n3244), .B(n3243), .Z(\round_in[0][315] ) );
  NAND U8944 ( .A(init), .B(round_reg[316]), .Z(n3246) );
  NANDN U8945 ( .A(init), .B(in[316]), .Z(n3245) );
  NAND U8946 ( .A(n3246), .B(n3245), .Z(\round_in[0][316] ) );
  NAND U8947 ( .A(init), .B(round_reg[317]), .Z(n3248) );
  NANDN U8948 ( .A(init), .B(in[317]), .Z(n3247) );
  NAND U8949 ( .A(n3248), .B(n3247), .Z(\round_in[0][317] ) );
  NAND U8950 ( .A(init), .B(round_reg[318]), .Z(n3250) );
  NANDN U8951 ( .A(init), .B(in[318]), .Z(n3249) );
  NAND U8952 ( .A(n3250), .B(n3249), .Z(\round_in[0][318] ) );
  NAND U8953 ( .A(init), .B(round_reg[319]), .Z(n3252) );
  NANDN U8954 ( .A(init), .B(in[319]), .Z(n3251) );
  NAND U8955 ( .A(n3252), .B(n3251), .Z(\round_in[0][319] ) );
  NAND U8956 ( .A(init), .B(round_reg[31]), .Z(n3254) );
  NANDN U8957 ( .A(init), .B(in[31]), .Z(n3253) );
  NAND U8958 ( .A(n3254), .B(n3253), .Z(\round_in[0][31] ) );
  NAND U8959 ( .A(init), .B(round_reg[320]), .Z(n3256) );
  NANDN U8960 ( .A(init), .B(in[320]), .Z(n3255) );
  NAND U8961 ( .A(n3256), .B(n3255), .Z(\round_in[0][320] ) );
  NAND U8962 ( .A(init), .B(round_reg[321]), .Z(n3258) );
  NANDN U8963 ( .A(init), .B(in[321]), .Z(n3257) );
  NAND U8964 ( .A(n3258), .B(n3257), .Z(\round_in[0][321] ) );
  NAND U8965 ( .A(init), .B(round_reg[322]), .Z(n3260) );
  NANDN U8966 ( .A(init), .B(in[322]), .Z(n3259) );
  NAND U8967 ( .A(n3260), .B(n3259), .Z(\round_in[0][322] ) );
  NAND U8968 ( .A(init), .B(round_reg[323]), .Z(n3262) );
  NANDN U8969 ( .A(init), .B(in[323]), .Z(n3261) );
  NAND U8970 ( .A(n3262), .B(n3261), .Z(\round_in[0][323] ) );
  NAND U8971 ( .A(init), .B(round_reg[324]), .Z(n3264) );
  NANDN U8972 ( .A(init), .B(in[324]), .Z(n3263) );
  NAND U8973 ( .A(n3264), .B(n3263), .Z(\round_in[0][324] ) );
  NAND U8974 ( .A(init), .B(round_reg[325]), .Z(n3266) );
  NANDN U8975 ( .A(init), .B(in[325]), .Z(n3265) );
  NAND U8976 ( .A(n3266), .B(n3265), .Z(\round_in[0][325] ) );
  NAND U8977 ( .A(init), .B(round_reg[326]), .Z(n3268) );
  NANDN U8978 ( .A(init), .B(in[326]), .Z(n3267) );
  NAND U8979 ( .A(n3268), .B(n3267), .Z(\round_in[0][326] ) );
  NAND U8980 ( .A(init), .B(round_reg[327]), .Z(n3270) );
  NANDN U8981 ( .A(init), .B(in[327]), .Z(n3269) );
  NAND U8982 ( .A(n3270), .B(n3269), .Z(\round_in[0][327] ) );
  NAND U8983 ( .A(init), .B(round_reg[328]), .Z(n3272) );
  NANDN U8984 ( .A(init), .B(in[328]), .Z(n3271) );
  NAND U8985 ( .A(n3272), .B(n3271), .Z(\round_in[0][328] ) );
  NAND U8986 ( .A(init), .B(round_reg[329]), .Z(n3274) );
  NANDN U8987 ( .A(init), .B(in[329]), .Z(n3273) );
  NAND U8988 ( .A(n3274), .B(n3273), .Z(\round_in[0][329] ) );
  NAND U8989 ( .A(init), .B(round_reg[32]), .Z(n3276) );
  NANDN U8990 ( .A(init), .B(in[32]), .Z(n3275) );
  NAND U8991 ( .A(n3276), .B(n3275), .Z(\round_in[0][32] ) );
  NAND U8992 ( .A(init), .B(round_reg[330]), .Z(n3278) );
  NANDN U8993 ( .A(init), .B(in[330]), .Z(n3277) );
  NAND U8994 ( .A(n3278), .B(n3277), .Z(\round_in[0][330] ) );
  NAND U8995 ( .A(init), .B(round_reg[331]), .Z(n3280) );
  NANDN U8996 ( .A(init), .B(in[331]), .Z(n3279) );
  NAND U8997 ( .A(n3280), .B(n3279), .Z(\round_in[0][331] ) );
  NAND U8998 ( .A(init), .B(round_reg[332]), .Z(n3282) );
  NANDN U8999 ( .A(init), .B(in[332]), .Z(n3281) );
  NAND U9000 ( .A(n3282), .B(n3281), .Z(\round_in[0][332] ) );
  NAND U9001 ( .A(init), .B(round_reg[333]), .Z(n3284) );
  NANDN U9002 ( .A(init), .B(in[333]), .Z(n3283) );
  NAND U9003 ( .A(n3284), .B(n3283), .Z(\round_in[0][333] ) );
  NAND U9004 ( .A(init), .B(round_reg[334]), .Z(n3286) );
  NANDN U9005 ( .A(init), .B(in[334]), .Z(n3285) );
  NAND U9006 ( .A(n3286), .B(n3285), .Z(\round_in[0][334] ) );
  NAND U9007 ( .A(init), .B(round_reg[335]), .Z(n3288) );
  NANDN U9008 ( .A(init), .B(in[335]), .Z(n3287) );
  NAND U9009 ( .A(n3288), .B(n3287), .Z(\round_in[0][335] ) );
  NAND U9010 ( .A(init), .B(round_reg[336]), .Z(n3290) );
  NANDN U9011 ( .A(init), .B(in[336]), .Z(n3289) );
  NAND U9012 ( .A(n3290), .B(n3289), .Z(\round_in[0][336] ) );
  NAND U9013 ( .A(init), .B(round_reg[337]), .Z(n3292) );
  NANDN U9014 ( .A(init), .B(in[337]), .Z(n3291) );
  NAND U9015 ( .A(n3292), .B(n3291), .Z(\round_in[0][337] ) );
  NAND U9016 ( .A(init), .B(round_reg[338]), .Z(n3294) );
  NANDN U9017 ( .A(init), .B(in[338]), .Z(n3293) );
  NAND U9018 ( .A(n3294), .B(n3293), .Z(\round_in[0][338] ) );
  NAND U9019 ( .A(init), .B(round_reg[339]), .Z(n3296) );
  NANDN U9020 ( .A(init), .B(in[339]), .Z(n3295) );
  NAND U9021 ( .A(n3296), .B(n3295), .Z(\round_in[0][339] ) );
  NAND U9022 ( .A(init), .B(round_reg[33]), .Z(n3298) );
  NANDN U9023 ( .A(init), .B(in[33]), .Z(n3297) );
  NAND U9024 ( .A(n3298), .B(n3297), .Z(\round_in[0][33] ) );
  NAND U9025 ( .A(init), .B(round_reg[340]), .Z(n3300) );
  NANDN U9026 ( .A(init), .B(in[340]), .Z(n3299) );
  NAND U9027 ( .A(n3300), .B(n3299), .Z(\round_in[0][340] ) );
  NAND U9028 ( .A(init), .B(round_reg[341]), .Z(n3302) );
  NANDN U9029 ( .A(init), .B(in[341]), .Z(n3301) );
  NAND U9030 ( .A(n3302), .B(n3301), .Z(\round_in[0][341] ) );
  NAND U9031 ( .A(init), .B(round_reg[342]), .Z(n3304) );
  NANDN U9032 ( .A(init), .B(in[342]), .Z(n3303) );
  NAND U9033 ( .A(n3304), .B(n3303), .Z(\round_in[0][342] ) );
  NAND U9034 ( .A(init), .B(round_reg[343]), .Z(n3306) );
  NANDN U9035 ( .A(init), .B(in[343]), .Z(n3305) );
  NAND U9036 ( .A(n3306), .B(n3305), .Z(\round_in[0][343] ) );
  NAND U9037 ( .A(init), .B(round_reg[344]), .Z(n3308) );
  NANDN U9038 ( .A(init), .B(in[344]), .Z(n3307) );
  NAND U9039 ( .A(n3308), .B(n3307), .Z(\round_in[0][344] ) );
  NAND U9040 ( .A(init), .B(round_reg[345]), .Z(n3310) );
  NANDN U9041 ( .A(init), .B(in[345]), .Z(n3309) );
  NAND U9042 ( .A(n3310), .B(n3309), .Z(\round_in[0][345] ) );
  NAND U9043 ( .A(init), .B(round_reg[346]), .Z(n3312) );
  NANDN U9044 ( .A(init), .B(in[346]), .Z(n3311) );
  NAND U9045 ( .A(n3312), .B(n3311), .Z(\round_in[0][346] ) );
  NAND U9046 ( .A(init), .B(round_reg[347]), .Z(n3314) );
  NANDN U9047 ( .A(init), .B(in[347]), .Z(n3313) );
  NAND U9048 ( .A(n3314), .B(n3313), .Z(\round_in[0][347] ) );
  NAND U9049 ( .A(init), .B(round_reg[348]), .Z(n3316) );
  NANDN U9050 ( .A(init), .B(in[348]), .Z(n3315) );
  NAND U9051 ( .A(n3316), .B(n3315), .Z(\round_in[0][348] ) );
  NAND U9052 ( .A(init), .B(round_reg[349]), .Z(n3318) );
  NANDN U9053 ( .A(init), .B(in[349]), .Z(n3317) );
  NAND U9054 ( .A(n3318), .B(n3317), .Z(\round_in[0][349] ) );
  NAND U9055 ( .A(init), .B(round_reg[34]), .Z(n3320) );
  NANDN U9056 ( .A(init), .B(in[34]), .Z(n3319) );
  NAND U9057 ( .A(n3320), .B(n3319), .Z(\round_in[0][34] ) );
  NAND U9058 ( .A(init), .B(round_reg[350]), .Z(n3322) );
  NANDN U9059 ( .A(init), .B(in[350]), .Z(n3321) );
  NAND U9060 ( .A(n3322), .B(n3321), .Z(\round_in[0][350] ) );
  NAND U9061 ( .A(init), .B(round_reg[351]), .Z(n3324) );
  NANDN U9062 ( .A(init), .B(in[351]), .Z(n3323) );
  NAND U9063 ( .A(n3324), .B(n3323), .Z(\round_in[0][351] ) );
  NAND U9064 ( .A(init), .B(round_reg[352]), .Z(n3326) );
  NANDN U9065 ( .A(init), .B(in[352]), .Z(n3325) );
  NAND U9066 ( .A(n3326), .B(n3325), .Z(\round_in[0][352] ) );
  NAND U9067 ( .A(init), .B(round_reg[353]), .Z(n3328) );
  NANDN U9068 ( .A(init), .B(in[353]), .Z(n3327) );
  NAND U9069 ( .A(n3328), .B(n3327), .Z(\round_in[0][353] ) );
  NAND U9070 ( .A(init), .B(round_reg[354]), .Z(n3330) );
  NANDN U9071 ( .A(init), .B(in[354]), .Z(n3329) );
  NAND U9072 ( .A(n3330), .B(n3329), .Z(\round_in[0][354] ) );
  NAND U9073 ( .A(init), .B(round_reg[355]), .Z(n3332) );
  NANDN U9074 ( .A(init), .B(in[355]), .Z(n3331) );
  NAND U9075 ( .A(n3332), .B(n3331), .Z(\round_in[0][355] ) );
  NAND U9076 ( .A(init), .B(round_reg[356]), .Z(n3334) );
  NANDN U9077 ( .A(init), .B(in[356]), .Z(n3333) );
  NAND U9078 ( .A(n3334), .B(n3333), .Z(\round_in[0][356] ) );
  NAND U9079 ( .A(init), .B(round_reg[357]), .Z(n3336) );
  NANDN U9080 ( .A(init), .B(in[357]), .Z(n3335) );
  NAND U9081 ( .A(n3336), .B(n3335), .Z(\round_in[0][357] ) );
  NAND U9082 ( .A(init), .B(round_reg[358]), .Z(n3338) );
  NANDN U9083 ( .A(init), .B(in[358]), .Z(n3337) );
  NAND U9084 ( .A(n3338), .B(n3337), .Z(\round_in[0][358] ) );
  NAND U9085 ( .A(init), .B(round_reg[359]), .Z(n3340) );
  NANDN U9086 ( .A(init), .B(in[359]), .Z(n3339) );
  NAND U9087 ( .A(n3340), .B(n3339), .Z(\round_in[0][359] ) );
  NAND U9088 ( .A(init), .B(round_reg[35]), .Z(n3342) );
  NANDN U9089 ( .A(init), .B(in[35]), .Z(n3341) );
  NAND U9090 ( .A(n3342), .B(n3341), .Z(\round_in[0][35] ) );
  NAND U9091 ( .A(init), .B(round_reg[360]), .Z(n3344) );
  NANDN U9092 ( .A(init), .B(in[360]), .Z(n3343) );
  NAND U9093 ( .A(n3344), .B(n3343), .Z(\round_in[0][360] ) );
  NAND U9094 ( .A(init), .B(round_reg[361]), .Z(n3346) );
  NANDN U9095 ( .A(init), .B(in[361]), .Z(n3345) );
  NAND U9096 ( .A(n3346), .B(n3345), .Z(\round_in[0][361] ) );
  NAND U9097 ( .A(init), .B(round_reg[362]), .Z(n3348) );
  NANDN U9098 ( .A(init), .B(in[362]), .Z(n3347) );
  NAND U9099 ( .A(n3348), .B(n3347), .Z(\round_in[0][362] ) );
  NAND U9100 ( .A(init), .B(round_reg[363]), .Z(n3350) );
  NANDN U9101 ( .A(init), .B(in[363]), .Z(n3349) );
  NAND U9102 ( .A(n3350), .B(n3349), .Z(\round_in[0][363] ) );
  NAND U9103 ( .A(init), .B(round_reg[364]), .Z(n3352) );
  NANDN U9104 ( .A(init), .B(in[364]), .Z(n3351) );
  NAND U9105 ( .A(n3352), .B(n3351), .Z(\round_in[0][364] ) );
  NAND U9106 ( .A(init), .B(round_reg[365]), .Z(n3354) );
  NANDN U9107 ( .A(init), .B(in[365]), .Z(n3353) );
  NAND U9108 ( .A(n3354), .B(n3353), .Z(\round_in[0][365] ) );
  NAND U9109 ( .A(init), .B(round_reg[366]), .Z(n3356) );
  NANDN U9110 ( .A(init), .B(in[366]), .Z(n3355) );
  NAND U9111 ( .A(n3356), .B(n3355), .Z(\round_in[0][366] ) );
  NAND U9112 ( .A(init), .B(round_reg[367]), .Z(n3358) );
  NANDN U9113 ( .A(init), .B(in[367]), .Z(n3357) );
  NAND U9114 ( .A(n3358), .B(n3357), .Z(\round_in[0][367] ) );
  NAND U9115 ( .A(init), .B(round_reg[368]), .Z(n3360) );
  NANDN U9116 ( .A(init), .B(in[368]), .Z(n3359) );
  NAND U9117 ( .A(n3360), .B(n3359), .Z(\round_in[0][368] ) );
  NAND U9118 ( .A(init), .B(round_reg[369]), .Z(n3362) );
  NANDN U9119 ( .A(init), .B(in[369]), .Z(n3361) );
  NAND U9120 ( .A(n3362), .B(n3361), .Z(\round_in[0][369] ) );
  NAND U9121 ( .A(init), .B(round_reg[36]), .Z(n3364) );
  NANDN U9122 ( .A(init), .B(in[36]), .Z(n3363) );
  NAND U9123 ( .A(n3364), .B(n3363), .Z(\round_in[0][36] ) );
  NAND U9124 ( .A(init), .B(round_reg[370]), .Z(n3366) );
  NANDN U9125 ( .A(init), .B(in[370]), .Z(n3365) );
  NAND U9126 ( .A(n3366), .B(n3365), .Z(\round_in[0][370] ) );
  NAND U9127 ( .A(init), .B(round_reg[371]), .Z(n3368) );
  NANDN U9128 ( .A(init), .B(in[371]), .Z(n3367) );
  NAND U9129 ( .A(n3368), .B(n3367), .Z(\round_in[0][371] ) );
  NAND U9130 ( .A(init), .B(round_reg[372]), .Z(n3370) );
  NANDN U9131 ( .A(init), .B(in[372]), .Z(n3369) );
  NAND U9132 ( .A(n3370), .B(n3369), .Z(\round_in[0][372] ) );
  NAND U9133 ( .A(init), .B(round_reg[373]), .Z(n3372) );
  NANDN U9134 ( .A(init), .B(in[373]), .Z(n3371) );
  NAND U9135 ( .A(n3372), .B(n3371), .Z(\round_in[0][373] ) );
  NAND U9136 ( .A(init), .B(round_reg[374]), .Z(n3374) );
  NANDN U9137 ( .A(init), .B(in[374]), .Z(n3373) );
  NAND U9138 ( .A(n3374), .B(n3373), .Z(\round_in[0][374] ) );
  NAND U9139 ( .A(init), .B(round_reg[375]), .Z(n3376) );
  NANDN U9140 ( .A(init), .B(in[375]), .Z(n3375) );
  NAND U9141 ( .A(n3376), .B(n3375), .Z(\round_in[0][375] ) );
  NAND U9142 ( .A(init), .B(round_reg[376]), .Z(n3378) );
  NANDN U9143 ( .A(init), .B(in[376]), .Z(n3377) );
  NAND U9144 ( .A(n3378), .B(n3377), .Z(\round_in[0][376] ) );
  NAND U9145 ( .A(init), .B(round_reg[377]), .Z(n3380) );
  NANDN U9146 ( .A(init), .B(in[377]), .Z(n3379) );
  NAND U9147 ( .A(n3380), .B(n3379), .Z(\round_in[0][377] ) );
  NAND U9148 ( .A(init), .B(round_reg[378]), .Z(n3382) );
  NANDN U9149 ( .A(init), .B(in[378]), .Z(n3381) );
  NAND U9150 ( .A(n3382), .B(n3381), .Z(\round_in[0][378] ) );
  NAND U9151 ( .A(init), .B(round_reg[379]), .Z(n3384) );
  NANDN U9152 ( .A(init), .B(in[379]), .Z(n3383) );
  NAND U9153 ( .A(n3384), .B(n3383), .Z(\round_in[0][379] ) );
  NAND U9154 ( .A(init), .B(round_reg[37]), .Z(n3386) );
  NANDN U9155 ( .A(init), .B(in[37]), .Z(n3385) );
  NAND U9156 ( .A(n3386), .B(n3385), .Z(\round_in[0][37] ) );
  NAND U9157 ( .A(init), .B(round_reg[380]), .Z(n3388) );
  NANDN U9158 ( .A(init), .B(in[380]), .Z(n3387) );
  NAND U9159 ( .A(n3388), .B(n3387), .Z(\round_in[0][380] ) );
  NAND U9160 ( .A(init), .B(round_reg[381]), .Z(n3390) );
  NANDN U9161 ( .A(init), .B(in[381]), .Z(n3389) );
  NAND U9162 ( .A(n3390), .B(n3389), .Z(\round_in[0][381] ) );
  NAND U9163 ( .A(init), .B(round_reg[382]), .Z(n3392) );
  NANDN U9164 ( .A(init), .B(in[382]), .Z(n3391) );
  NAND U9165 ( .A(n3392), .B(n3391), .Z(\round_in[0][382] ) );
  NAND U9166 ( .A(init), .B(round_reg[383]), .Z(n3394) );
  NANDN U9167 ( .A(init), .B(in[383]), .Z(n3393) );
  NAND U9168 ( .A(n3394), .B(n3393), .Z(\round_in[0][383] ) );
  NAND U9169 ( .A(init), .B(round_reg[384]), .Z(n3396) );
  NANDN U9170 ( .A(init), .B(in[384]), .Z(n3395) );
  NAND U9171 ( .A(n3396), .B(n3395), .Z(\round_in[0][384] ) );
  NAND U9172 ( .A(init), .B(round_reg[385]), .Z(n3398) );
  NANDN U9173 ( .A(init), .B(in[385]), .Z(n3397) );
  NAND U9174 ( .A(n3398), .B(n3397), .Z(\round_in[0][385] ) );
  NAND U9175 ( .A(init), .B(round_reg[386]), .Z(n3400) );
  NANDN U9176 ( .A(init), .B(in[386]), .Z(n3399) );
  NAND U9177 ( .A(n3400), .B(n3399), .Z(\round_in[0][386] ) );
  NAND U9178 ( .A(init), .B(round_reg[387]), .Z(n3402) );
  NANDN U9179 ( .A(init), .B(in[387]), .Z(n3401) );
  NAND U9180 ( .A(n3402), .B(n3401), .Z(\round_in[0][387] ) );
  NAND U9181 ( .A(init), .B(round_reg[388]), .Z(n3404) );
  NANDN U9182 ( .A(init), .B(in[388]), .Z(n3403) );
  NAND U9183 ( .A(n3404), .B(n3403), .Z(\round_in[0][388] ) );
  NAND U9184 ( .A(init), .B(round_reg[389]), .Z(n3406) );
  NANDN U9185 ( .A(init), .B(in[389]), .Z(n3405) );
  NAND U9186 ( .A(n3406), .B(n3405), .Z(\round_in[0][389] ) );
  NAND U9187 ( .A(init), .B(round_reg[38]), .Z(n3408) );
  NANDN U9188 ( .A(init), .B(in[38]), .Z(n3407) );
  NAND U9189 ( .A(n3408), .B(n3407), .Z(\round_in[0][38] ) );
  NAND U9190 ( .A(init), .B(round_reg[390]), .Z(n3410) );
  NANDN U9191 ( .A(init), .B(in[390]), .Z(n3409) );
  NAND U9192 ( .A(n3410), .B(n3409), .Z(\round_in[0][390] ) );
  NAND U9193 ( .A(init), .B(round_reg[391]), .Z(n3412) );
  NANDN U9194 ( .A(init), .B(in[391]), .Z(n3411) );
  NAND U9195 ( .A(n3412), .B(n3411), .Z(\round_in[0][391] ) );
  NAND U9196 ( .A(init), .B(round_reg[392]), .Z(n3414) );
  NANDN U9197 ( .A(init), .B(in[392]), .Z(n3413) );
  NAND U9198 ( .A(n3414), .B(n3413), .Z(\round_in[0][392] ) );
  NAND U9199 ( .A(init), .B(round_reg[393]), .Z(n3416) );
  NANDN U9200 ( .A(init), .B(in[393]), .Z(n3415) );
  NAND U9201 ( .A(n3416), .B(n3415), .Z(\round_in[0][393] ) );
  NAND U9202 ( .A(init), .B(round_reg[394]), .Z(n3418) );
  NANDN U9203 ( .A(init), .B(in[394]), .Z(n3417) );
  NAND U9204 ( .A(n3418), .B(n3417), .Z(\round_in[0][394] ) );
  NAND U9205 ( .A(init), .B(round_reg[395]), .Z(n3420) );
  NANDN U9206 ( .A(init), .B(in[395]), .Z(n3419) );
  NAND U9207 ( .A(n3420), .B(n3419), .Z(\round_in[0][395] ) );
  NAND U9208 ( .A(init), .B(round_reg[396]), .Z(n3422) );
  NANDN U9209 ( .A(init), .B(in[396]), .Z(n3421) );
  NAND U9210 ( .A(n3422), .B(n3421), .Z(\round_in[0][396] ) );
  NAND U9211 ( .A(init), .B(round_reg[397]), .Z(n3424) );
  NANDN U9212 ( .A(init), .B(in[397]), .Z(n3423) );
  NAND U9213 ( .A(n3424), .B(n3423), .Z(\round_in[0][397] ) );
  NAND U9214 ( .A(init), .B(round_reg[398]), .Z(n3426) );
  NANDN U9215 ( .A(init), .B(in[398]), .Z(n3425) );
  NAND U9216 ( .A(n3426), .B(n3425), .Z(\round_in[0][398] ) );
  NAND U9217 ( .A(init), .B(round_reg[399]), .Z(n3428) );
  NANDN U9218 ( .A(init), .B(in[399]), .Z(n3427) );
  NAND U9219 ( .A(n3428), .B(n3427), .Z(\round_in[0][399] ) );
  NAND U9220 ( .A(init), .B(round_reg[39]), .Z(n3430) );
  NANDN U9221 ( .A(init), .B(in[39]), .Z(n3429) );
  NAND U9222 ( .A(n3430), .B(n3429), .Z(\round_in[0][39] ) );
  NAND U9223 ( .A(init), .B(round_reg[3]), .Z(n3432) );
  NANDN U9224 ( .A(init), .B(in[3]), .Z(n3431) );
  NAND U9225 ( .A(n3432), .B(n3431), .Z(\round_in[0][3] ) );
  NAND U9226 ( .A(init), .B(round_reg[400]), .Z(n3434) );
  NANDN U9227 ( .A(init), .B(in[400]), .Z(n3433) );
  NAND U9228 ( .A(n3434), .B(n3433), .Z(\round_in[0][400] ) );
  NAND U9229 ( .A(init), .B(round_reg[401]), .Z(n3436) );
  NANDN U9230 ( .A(init), .B(in[401]), .Z(n3435) );
  NAND U9231 ( .A(n3436), .B(n3435), .Z(\round_in[0][401] ) );
  NAND U9232 ( .A(init), .B(round_reg[402]), .Z(n3438) );
  NANDN U9233 ( .A(init), .B(in[402]), .Z(n3437) );
  NAND U9234 ( .A(n3438), .B(n3437), .Z(\round_in[0][402] ) );
  NAND U9235 ( .A(init), .B(round_reg[403]), .Z(n3440) );
  NANDN U9236 ( .A(init), .B(in[403]), .Z(n3439) );
  NAND U9237 ( .A(n3440), .B(n3439), .Z(\round_in[0][403] ) );
  NAND U9238 ( .A(init), .B(round_reg[404]), .Z(n3442) );
  NANDN U9239 ( .A(init), .B(in[404]), .Z(n3441) );
  NAND U9240 ( .A(n3442), .B(n3441), .Z(\round_in[0][404] ) );
  NAND U9241 ( .A(init), .B(round_reg[405]), .Z(n3444) );
  NANDN U9242 ( .A(init), .B(in[405]), .Z(n3443) );
  NAND U9243 ( .A(n3444), .B(n3443), .Z(\round_in[0][405] ) );
  NAND U9244 ( .A(init), .B(round_reg[406]), .Z(n3446) );
  NANDN U9245 ( .A(init), .B(in[406]), .Z(n3445) );
  NAND U9246 ( .A(n3446), .B(n3445), .Z(\round_in[0][406] ) );
  NAND U9247 ( .A(init), .B(round_reg[407]), .Z(n3448) );
  NANDN U9248 ( .A(init), .B(in[407]), .Z(n3447) );
  NAND U9249 ( .A(n3448), .B(n3447), .Z(\round_in[0][407] ) );
  NAND U9250 ( .A(init), .B(round_reg[408]), .Z(n3450) );
  NANDN U9251 ( .A(init), .B(in[408]), .Z(n3449) );
  NAND U9252 ( .A(n3450), .B(n3449), .Z(\round_in[0][408] ) );
  NAND U9253 ( .A(init), .B(round_reg[409]), .Z(n3452) );
  NANDN U9254 ( .A(init), .B(in[409]), .Z(n3451) );
  NAND U9255 ( .A(n3452), .B(n3451), .Z(\round_in[0][409] ) );
  NAND U9256 ( .A(init), .B(round_reg[40]), .Z(n3454) );
  NANDN U9257 ( .A(init), .B(in[40]), .Z(n3453) );
  NAND U9258 ( .A(n3454), .B(n3453), .Z(\round_in[0][40] ) );
  NAND U9259 ( .A(init), .B(round_reg[410]), .Z(n3456) );
  NANDN U9260 ( .A(init), .B(in[410]), .Z(n3455) );
  NAND U9261 ( .A(n3456), .B(n3455), .Z(\round_in[0][410] ) );
  NAND U9262 ( .A(init), .B(round_reg[411]), .Z(n3458) );
  NANDN U9263 ( .A(init), .B(in[411]), .Z(n3457) );
  NAND U9264 ( .A(n3458), .B(n3457), .Z(\round_in[0][411] ) );
  NAND U9265 ( .A(init), .B(round_reg[412]), .Z(n3460) );
  NANDN U9266 ( .A(init), .B(in[412]), .Z(n3459) );
  NAND U9267 ( .A(n3460), .B(n3459), .Z(\round_in[0][412] ) );
  NAND U9268 ( .A(init), .B(round_reg[413]), .Z(n3462) );
  NANDN U9269 ( .A(init), .B(in[413]), .Z(n3461) );
  NAND U9270 ( .A(n3462), .B(n3461), .Z(\round_in[0][413] ) );
  NAND U9271 ( .A(init), .B(round_reg[414]), .Z(n3464) );
  NANDN U9272 ( .A(init), .B(in[414]), .Z(n3463) );
  NAND U9273 ( .A(n3464), .B(n3463), .Z(\round_in[0][414] ) );
  NAND U9274 ( .A(init), .B(round_reg[415]), .Z(n3466) );
  NANDN U9275 ( .A(init), .B(in[415]), .Z(n3465) );
  NAND U9276 ( .A(n3466), .B(n3465), .Z(\round_in[0][415] ) );
  NAND U9277 ( .A(init), .B(round_reg[416]), .Z(n3468) );
  NANDN U9278 ( .A(init), .B(in[416]), .Z(n3467) );
  NAND U9279 ( .A(n3468), .B(n3467), .Z(\round_in[0][416] ) );
  NAND U9280 ( .A(init), .B(round_reg[417]), .Z(n3470) );
  NANDN U9281 ( .A(init), .B(in[417]), .Z(n3469) );
  NAND U9282 ( .A(n3470), .B(n3469), .Z(\round_in[0][417] ) );
  NAND U9283 ( .A(init), .B(round_reg[418]), .Z(n3472) );
  NANDN U9284 ( .A(init), .B(in[418]), .Z(n3471) );
  NAND U9285 ( .A(n3472), .B(n3471), .Z(\round_in[0][418] ) );
  NAND U9286 ( .A(init), .B(round_reg[419]), .Z(n3474) );
  NANDN U9287 ( .A(init), .B(in[419]), .Z(n3473) );
  NAND U9288 ( .A(n3474), .B(n3473), .Z(\round_in[0][419] ) );
  NAND U9289 ( .A(init), .B(round_reg[41]), .Z(n3476) );
  NANDN U9290 ( .A(init), .B(in[41]), .Z(n3475) );
  NAND U9291 ( .A(n3476), .B(n3475), .Z(\round_in[0][41] ) );
  NAND U9292 ( .A(init), .B(round_reg[420]), .Z(n3478) );
  NANDN U9293 ( .A(init), .B(in[420]), .Z(n3477) );
  NAND U9294 ( .A(n3478), .B(n3477), .Z(\round_in[0][420] ) );
  NAND U9295 ( .A(init), .B(round_reg[421]), .Z(n3480) );
  NANDN U9296 ( .A(init), .B(in[421]), .Z(n3479) );
  NAND U9297 ( .A(n3480), .B(n3479), .Z(\round_in[0][421] ) );
  NAND U9298 ( .A(init), .B(round_reg[422]), .Z(n3482) );
  NANDN U9299 ( .A(init), .B(in[422]), .Z(n3481) );
  NAND U9300 ( .A(n3482), .B(n3481), .Z(\round_in[0][422] ) );
  NAND U9301 ( .A(init), .B(round_reg[423]), .Z(n3484) );
  NANDN U9302 ( .A(init), .B(in[423]), .Z(n3483) );
  NAND U9303 ( .A(n3484), .B(n3483), .Z(\round_in[0][423] ) );
  NAND U9304 ( .A(init), .B(round_reg[424]), .Z(n3486) );
  NANDN U9305 ( .A(init), .B(in[424]), .Z(n3485) );
  NAND U9306 ( .A(n3486), .B(n3485), .Z(\round_in[0][424] ) );
  NAND U9307 ( .A(init), .B(round_reg[425]), .Z(n3488) );
  NANDN U9308 ( .A(init), .B(in[425]), .Z(n3487) );
  NAND U9309 ( .A(n3488), .B(n3487), .Z(\round_in[0][425] ) );
  NAND U9310 ( .A(init), .B(round_reg[426]), .Z(n3490) );
  NANDN U9311 ( .A(init), .B(in[426]), .Z(n3489) );
  NAND U9312 ( .A(n3490), .B(n3489), .Z(\round_in[0][426] ) );
  NAND U9313 ( .A(init), .B(round_reg[427]), .Z(n3492) );
  NANDN U9314 ( .A(init), .B(in[427]), .Z(n3491) );
  NAND U9315 ( .A(n3492), .B(n3491), .Z(\round_in[0][427] ) );
  NAND U9316 ( .A(init), .B(round_reg[428]), .Z(n3494) );
  NANDN U9317 ( .A(init), .B(in[428]), .Z(n3493) );
  NAND U9318 ( .A(n3494), .B(n3493), .Z(\round_in[0][428] ) );
  NAND U9319 ( .A(init), .B(round_reg[429]), .Z(n3496) );
  NANDN U9320 ( .A(init), .B(in[429]), .Z(n3495) );
  NAND U9321 ( .A(n3496), .B(n3495), .Z(\round_in[0][429] ) );
  NAND U9322 ( .A(init), .B(round_reg[42]), .Z(n3498) );
  NANDN U9323 ( .A(init), .B(in[42]), .Z(n3497) );
  NAND U9324 ( .A(n3498), .B(n3497), .Z(\round_in[0][42] ) );
  NAND U9325 ( .A(init), .B(round_reg[430]), .Z(n3500) );
  NANDN U9326 ( .A(init), .B(in[430]), .Z(n3499) );
  NAND U9327 ( .A(n3500), .B(n3499), .Z(\round_in[0][430] ) );
  NAND U9328 ( .A(init), .B(round_reg[431]), .Z(n3502) );
  NANDN U9329 ( .A(init), .B(in[431]), .Z(n3501) );
  NAND U9330 ( .A(n3502), .B(n3501), .Z(\round_in[0][431] ) );
  NAND U9331 ( .A(init), .B(round_reg[432]), .Z(n3504) );
  NANDN U9332 ( .A(init), .B(in[432]), .Z(n3503) );
  NAND U9333 ( .A(n3504), .B(n3503), .Z(\round_in[0][432] ) );
  NAND U9334 ( .A(init), .B(round_reg[433]), .Z(n3506) );
  NANDN U9335 ( .A(init), .B(in[433]), .Z(n3505) );
  NAND U9336 ( .A(n3506), .B(n3505), .Z(\round_in[0][433] ) );
  NAND U9337 ( .A(init), .B(round_reg[434]), .Z(n3508) );
  NANDN U9338 ( .A(init), .B(in[434]), .Z(n3507) );
  NAND U9339 ( .A(n3508), .B(n3507), .Z(\round_in[0][434] ) );
  NAND U9340 ( .A(init), .B(round_reg[435]), .Z(n3510) );
  NANDN U9341 ( .A(init), .B(in[435]), .Z(n3509) );
  NAND U9342 ( .A(n3510), .B(n3509), .Z(\round_in[0][435] ) );
  NAND U9343 ( .A(init), .B(round_reg[436]), .Z(n3512) );
  NANDN U9344 ( .A(init), .B(in[436]), .Z(n3511) );
  NAND U9345 ( .A(n3512), .B(n3511), .Z(\round_in[0][436] ) );
  NAND U9346 ( .A(init), .B(round_reg[437]), .Z(n3514) );
  NANDN U9347 ( .A(init), .B(in[437]), .Z(n3513) );
  NAND U9348 ( .A(n3514), .B(n3513), .Z(\round_in[0][437] ) );
  NAND U9349 ( .A(init), .B(round_reg[438]), .Z(n3516) );
  NANDN U9350 ( .A(init), .B(in[438]), .Z(n3515) );
  NAND U9351 ( .A(n3516), .B(n3515), .Z(\round_in[0][438] ) );
  NAND U9352 ( .A(init), .B(round_reg[439]), .Z(n3518) );
  NANDN U9353 ( .A(init), .B(in[439]), .Z(n3517) );
  NAND U9354 ( .A(n3518), .B(n3517), .Z(\round_in[0][439] ) );
  NAND U9355 ( .A(init), .B(round_reg[43]), .Z(n3520) );
  NANDN U9356 ( .A(init), .B(in[43]), .Z(n3519) );
  NAND U9357 ( .A(n3520), .B(n3519), .Z(\round_in[0][43] ) );
  NAND U9358 ( .A(init), .B(round_reg[440]), .Z(n3522) );
  NANDN U9359 ( .A(init), .B(in[440]), .Z(n3521) );
  NAND U9360 ( .A(n3522), .B(n3521), .Z(\round_in[0][440] ) );
  NAND U9361 ( .A(init), .B(round_reg[441]), .Z(n3524) );
  NANDN U9362 ( .A(init), .B(in[441]), .Z(n3523) );
  NAND U9363 ( .A(n3524), .B(n3523), .Z(\round_in[0][441] ) );
  NAND U9364 ( .A(init), .B(round_reg[442]), .Z(n3526) );
  NANDN U9365 ( .A(init), .B(in[442]), .Z(n3525) );
  NAND U9366 ( .A(n3526), .B(n3525), .Z(\round_in[0][442] ) );
  NAND U9367 ( .A(init), .B(round_reg[443]), .Z(n3528) );
  NANDN U9368 ( .A(init), .B(in[443]), .Z(n3527) );
  NAND U9369 ( .A(n3528), .B(n3527), .Z(\round_in[0][443] ) );
  NAND U9370 ( .A(init), .B(round_reg[444]), .Z(n3530) );
  NANDN U9371 ( .A(init), .B(in[444]), .Z(n3529) );
  NAND U9372 ( .A(n3530), .B(n3529), .Z(\round_in[0][444] ) );
  NAND U9373 ( .A(init), .B(round_reg[445]), .Z(n3532) );
  NANDN U9374 ( .A(init), .B(in[445]), .Z(n3531) );
  NAND U9375 ( .A(n3532), .B(n3531), .Z(\round_in[0][445] ) );
  NAND U9376 ( .A(init), .B(round_reg[446]), .Z(n3534) );
  NANDN U9377 ( .A(init), .B(in[446]), .Z(n3533) );
  NAND U9378 ( .A(n3534), .B(n3533), .Z(\round_in[0][446] ) );
  NAND U9379 ( .A(init), .B(round_reg[447]), .Z(n3536) );
  NANDN U9380 ( .A(init), .B(in[447]), .Z(n3535) );
  NAND U9381 ( .A(n3536), .B(n3535), .Z(\round_in[0][447] ) );
  NAND U9382 ( .A(init), .B(round_reg[448]), .Z(n3538) );
  NANDN U9383 ( .A(init), .B(in[448]), .Z(n3537) );
  NAND U9384 ( .A(n3538), .B(n3537), .Z(\round_in[0][448] ) );
  NAND U9385 ( .A(init), .B(round_reg[449]), .Z(n3540) );
  NANDN U9386 ( .A(init), .B(in[449]), .Z(n3539) );
  NAND U9387 ( .A(n3540), .B(n3539), .Z(\round_in[0][449] ) );
  NAND U9388 ( .A(init), .B(round_reg[44]), .Z(n3542) );
  NANDN U9389 ( .A(init), .B(in[44]), .Z(n3541) );
  NAND U9390 ( .A(n3542), .B(n3541), .Z(\round_in[0][44] ) );
  NAND U9391 ( .A(init), .B(round_reg[450]), .Z(n3544) );
  NANDN U9392 ( .A(init), .B(in[450]), .Z(n3543) );
  NAND U9393 ( .A(n3544), .B(n3543), .Z(\round_in[0][450] ) );
  NAND U9394 ( .A(init), .B(round_reg[451]), .Z(n3546) );
  NANDN U9395 ( .A(init), .B(in[451]), .Z(n3545) );
  NAND U9396 ( .A(n3546), .B(n3545), .Z(\round_in[0][451] ) );
  NAND U9397 ( .A(init), .B(round_reg[452]), .Z(n3548) );
  NANDN U9398 ( .A(init), .B(in[452]), .Z(n3547) );
  NAND U9399 ( .A(n3548), .B(n3547), .Z(\round_in[0][452] ) );
  NAND U9400 ( .A(init), .B(round_reg[453]), .Z(n3550) );
  NANDN U9401 ( .A(init), .B(in[453]), .Z(n3549) );
  NAND U9402 ( .A(n3550), .B(n3549), .Z(\round_in[0][453] ) );
  NAND U9403 ( .A(init), .B(round_reg[454]), .Z(n3552) );
  NANDN U9404 ( .A(init), .B(in[454]), .Z(n3551) );
  NAND U9405 ( .A(n3552), .B(n3551), .Z(\round_in[0][454] ) );
  NAND U9406 ( .A(init), .B(round_reg[455]), .Z(n3554) );
  NANDN U9407 ( .A(init), .B(in[455]), .Z(n3553) );
  NAND U9408 ( .A(n3554), .B(n3553), .Z(\round_in[0][455] ) );
  NAND U9409 ( .A(init), .B(round_reg[456]), .Z(n3556) );
  NANDN U9410 ( .A(init), .B(in[456]), .Z(n3555) );
  NAND U9411 ( .A(n3556), .B(n3555), .Z(\round_in[0][456] ) );
  NAND U9412 ( .A(init), .B(round_reg[457]), .Z(n3558) );
  NANDN U9413 ( .A(init), .B(in[457]), .Z(n3557) );
  NAND U9414 ( .A(n3558), .B(n3557), .Z(\round_in[0][457] ) );
  NAND U9415 ( .A(init), .B(round_reg[458]), .Z(n3560) );
  NANDN U9416 ( .A(init), .B(in[458]), .Z(n3559) );
  NAND U9417 ( .A(n3560), .B(n3559), .Z(\round_in[0][458] ) );
  NAND U9418 ( .A(init), .B(round_reg[459]), .Z(n3562) );
  NANDN U9419 ( .A(init), .B(in[459]), .Z(n3561) );
  NAND U9420 ( .A(n3562), .B(n3561), .Z(\round_in[0][459] ) );
  NAND U9421 ( .A(init), .B(round_reg[45]), .Z(n3564) );
  NANDN U9422 ( .A(init), .B(in[45]), .Z(n3563) );
  NAND U9423 ( .A(n3564), .B(n3563), .Z(\round_in[0][45] ) );
  NAND U9424 ( .A(init), .B(round_reg[460]), .Z(n3566) );
  NANDN U9425 ( .A(init), .B(in[460]), .Z(n3565) );
  NAND U9426 ( .A(n3566), .B(n3565), .Z(\round_in[0][460] ) );
  NAND U9427 ( .A(init), .B(round_reg[461]), .Z(n3568) );
  NANDN U9428 ( .A(init), .B(in[461]), .Z(n3567) );
  NAND U9429 ( .A(n3568), .B(n3567), .Z(\round_in[0][461] ) );
  NAND U9430 ( .A(init), .B(round_reg[462]), .Z(n3570) );
  NANDN U9431 ( .A(init), .B(in[462]), .Z(n3569) );
  NAND U9432 ( .A(n3570), .B(n3569), .Z(\round_in[0][462] ) );
  NAND U9433 ( .A(init), .B(round_reg[463]), .Z(n3572) );
  NANDN U9434 ( .A(init), .B(in[463]), .Z(n3571) );
  NAND U9435 ( .A(n3572), .B(n3571), .Z(\round_in[0][463] ) );
  NAND U9436 ( .A(init), .B(round_reg[464]), .Z(n3574) );
  NANDN U9437 ( .A(init), .B(in[464]), .Z(n3573) );
  NAND U9438 ( .A(n3574), .B(n3573), .Z(\round_in[0][464] ) );
  NAND U9439 ( .A(init), .B(round_reg[465]), .Z(n3576) );
  NANDN U9440 ( .A(init), .B(in[465]), .Z(n3575) );
  NAND U9441 ( .A(n3576), .B(n3575), .Z(\round_in[0][465] ) );
  NAND U9442 ( .A(init), .B(round_reg[466]), .Z(n3578) );
  NANDN U9443 ( .A(init), .B(in[466]), .Z(n3577) );
  NAND U9444 ( .A(n3578), .B(n3577), .Z(\round_in[0][466] ) );
  NAND U9445 ( .A(init), .B(round_reg[467]), .Z(n3580) );
  NANDN U9446 ( .A(init), .B(in[467]), .Z(n3579) );
  NAND U9447 ( .A(n3580), .B(n3579), .Z(\round_in[0][467] ) );
  NAND U9448 ( .A(init), .B(round_reg[468]), .Z(n3582) );
  NANDN U9449 ( .A(init), .B(in[468]), .Z(n3581) );
  NAND U9450 ( .A(n3582), .B(n3581), .Z(\round_in[0][468] ) );
  NAND U9451 ( .A(init), .B(round_reg[469]), .Z(n3584) );
  NANDN U9452 ( .A(init), .B(in[469]), .Z(n3583) );
  NAND U9453 ( .A(n3584), .B(n3583), .Z(\round_in[0][469] ) );
  NAND U9454 ( .A(init), .B(round_reg[46]), .Z(n3586) );
  NANDN U9455 ( .A(init), .B(in[46]), .Z(n3585) );
  NAND U9456 ( .A(n3586), .B(n3585), .Z(\round_in[0][46] ) );
  NAND U9457 ( .A(init), .B(round_reg[470]), .Z(n3588) );
  NANDN U9458 ( .A(init), .B(in[470]), .Z(n3587) );
  NAND U9459 ( .A(n3588), .B(n3587), .Z(\round_in[0][470] ) );
  NAND U9460 ( .A(init), .B(round_reg[471]), .Z(n3590) );
  NANDN U9461 ( .A(init), .B(in[471]), .Z(n3589) );
  NAND U9462 ( .A(n3590), .B(n3589), .Z(\round_in[0][471] ) );
  NAND U9463 ( .A(init), .B(round_reg[472]), .Z(n3592) );
  NANDN U9464 ( .A(init), .B(in[472]), .Z(n3591) );
  NAND U9465 ( .A(n3592), .B(n3591), .Z(\round_in[0][472] ) );
  NAND U9466 ( .A(init), .B(round_reg[473]), .Z(n3594) );
  NANDN U9467 ( .A(init), .B(in[473]), .Z(n3593) );
  NAND U9468 ( .A(n3594), .B(n3593), .Z(\round_in[0][473] ) );
  NAND U9469 ( .A(init), .B(round_reg[474]), .Z(n3596) );
  NANDN U9470 ( .A(init), .B(in[474]), .Z(n3595) );
  NAND U9471 ( .A(n3596), .B(n3595), .Z(\round_in[0][474] ) );
  NAND U9472 ( .A(init), .B(round_reg[475]), .Z(n3598) );
  NANDN U9473 ( .A(init), .B(in[475]), .Z(n3597) );
  NAND U9474 ( .A(n3598), .B(n3597), .Z(\round_in[0][475] ) );
  NAND U9475 ( .A(init), .B(round_reg[476]), .Z(n3600) );
  NANDN U9476 ( .A(init), .B(in[476]), .Z(n3599) );
  NAND U9477 ( .A(n3600), .B(n3599), .Z(\round_in[0][476] ) );
  NAND U9478 ( .A(init), .B(round_reg[477]), .Z(n3602) );
  NANDN U9479 ( .A(init), .B(in[477]), .Z(n3601) );
  NAND U9480 ( .A(n3602), .B(n3601), .Z(\round_in[0][477] ) );
  NAND U9481 ( .A(init), .B(round_reg[478]), .Z(n3604) );
  NANDN U9482 ( .A(init), .B(in[478]), .Z(n3603) );
  NAND U9483 ( .A(n3604), .B(n3603), .Z(\round_in[0][478] ) );
  NAND U9484 ( .A(init), .B(round_reg[479]), .Z(n3606) );
  NANDN U9485 ( .A(init), .B(in[479]), .Z(n3605) );
  NAND U9486 ( .A(n3606), .B(n3605), .Z(\round_in[0][479] ) );
  NAND U9487 ( .A(init), .B(round_reg[47]), .Z(n3608) );
  NANDN U9488 ( .A(init), .B(in[47]), .Z(n3607) );
  NAND U9489 ( .A(n3608), .B(n3607), .Z(\round_in[0][47] ) );
  NAND U9490 ( .A(init), .B(round_reg[480]), .Z(n3610) );
  NANDN U9491 ( .A(init), .B(in[480]), .Z(n3609) );
  NAND U9492 ( .A(n3610), .B(n3609), .Z(\round_in[0][480] ) );
  NAND U9493 ( .A(init), .B(round_reg[481]), .Z(n3612) );
  NANDN U9494 ( .A(init), .B(in[481]), .Z(n3611) );
  NAND U9495 ( .A(n3612), .B(n3611), .Z(\round_in[0][481] ) );
  NAND U9496 ( .A(init), .B(round_reg[482]), .Z(n3614) );
  NANDN U9497 ( .A(init), .B(in[482]), .Z(n3613) );
  NAND U9498 ( .A(n3614), .B(n3613), .Z(\round_in[0][482] ) );
  NAND U9499 ( .A(init), .B(round_reg[483]), .Z(n3616) );
  NANDN U9500 ( .A(init), .B(in[483]), .Z(n3615) );
  NAND U9501 ( .A(n3616), .B(n3615), .Z(\round_in[0][483] ) );
  NAND U9502 ( .A(init), .B(round_reg[484]), .Z(n3618) );
  NANDN U9503 ( .A(init), .B(in[484]), .Z(n3617) );
  NAND U9504 ( .A(n3618), .B(n3617), .Z(\round_in[0][484] ) );
  NAND U9505 ( .A(init), .B(round_reg[485]), .Z(n3620) );
  NANDN U9506 ( .A(init), .B(in[485]), .Z(n3619) );
  NAND U9507 ( .A(n3620), .B(n3619), .Z(\round_in[0][485] ) );
  NAND U9508 ( .A(init), .B(round_reg[486]), .Z(n3622) );
  NANDN U9509 ( .A(init), .B(in[486]), .Z(n3621) );
  NAND U9510 ( .A(n3622), .B(n3621), .Z(\round_in[0][486] ) );
  NAND U9511 ( .A(init), .B(round_reg[487]), .Z(n3624) );
  NANDN U9512 ( .A(init), .B(in[487]), .Z(n3623) );
  NAND U9513 ( .A(n3624), .B(n3623), .Z(\round_in[0][487] ) );
  NAND U9514 ( .A(init), .B(round_reg[488]), .Z(n3626) );
  NANDN U9515 ( .A(init), .B(in[488]), .Z(n3625) );
  NAND U9516 ( .A(n3626), .B(n3625), .Z(\round_in[0][488] ) );
  NAND U9517 ( .A(init), .B(round_reg[489]), .Z(n3628) );
  NANDN U9518 ( .A(init), .B(in[489]), .Z(n3627) );
  NAND U9519 ( .A(n3628), .B(n3627), .Z(\round_in[0][489] ) );
  NAND U9520 ( .A(init), .B(round_reg[48]), .Z(n3630) );
  NANDN U9521 ( .A(init), .B(in[48]), .Z(n3629) );
  NAND U9522 ( .A(n3630), .B(n3629), .Z(\round_in[0][48] ) );
  NAND U9523 ( .A(init), .B(round_reg[490]), .Z(n3632) );
  NANDN U9524 ( .A(init), .B(in[490]), .Z(n3631) );
  NAND U9525 ( .A(n3632), .B(n3631), .Z(\round_in[0][490] ) );
  NAND U9526 ( .A(init), .B(round_reg[491]), .Z(n3634) );
  NANDN U9527 ( .A(init), .B(in[491]), .Z(n3633) );
  NAND U9528 ( .A(n3634), .B(n3633), .Z(\round_in[0][491] ) );
  NAND U9529 ( .A(init), .B(round_reg[492]), .Z(n3636) );
  NANDN U9530 ( .A(init), .B(in[492]), .Z(n3635) );
  NAND U9531 ( .A(n3636), .B(n3635), .Z(\round_in[0][492] ) );
  NAND U9532 ( .A(init), .B(round_reg[493]), .Z(n3638) );
  NANDN U9533 ( .A(init), .B(in[493]), .Z(n3637) );
  NAND U9534 ( .A(n3638), .B(n3637), .Z(\round_in[0][493] ) );
  NAND U9535 ( .A(init), .B(round_reg[494]), .Z(n3640) );
  NANDN U9536 ( .A(init), .B(in[494]), .Z(n3639) );
  NAND U9537 ( .A(n3640), .B(n3639), .Z(\round_in[0][494] ) );
  NAND U9538 ( .A(init), .B(round_reg[495]), .Z(n3642) );
  NANDN U9539 ( .A(init), .B(in[495]), .Z(n3641) );
  NAND U9540 ( .A(n3642), .B(n3641), .Z(\round_in[0][495] ) );
  NAND U9541 ( .A(init), .B(round_reg[496]), .Z(n3644) );
  NANDN U9542 ( .A(init), .B(in[496]), .Z(n3643) );
  NAND U9543 ( .A(n3644), .B(n3643), .Z(\round_in[0][496] ) );
  NAND U9544 ( .A(init), .B(round_reg[497]), .Z(n3646) );
  NANDN U9545 ( .A(init), .B(in[497]), .Z(n3645) );
  NAND U9546 ( .A(n3646), .B(n3645), .Z(\round_in[0][497] ) );
  NAND U9547 ( .A(init), .B(round_reg[498]), .Z(n3648) );
  NANDN U9548 ( .A(init), .B(in[498]), .Z(n3647) );
  NAND U9549 ( .A(n3648), .B(n3647), .Z(\round_in[0][498] ) );
  NAND U9550 ( .A(init), .B(round_reg[499]), .Z(n3650) );
  NANDN U9551 ( .A(init), .B(in[499]), .Z(n3649) );
  NAND U9552 ( .A(n3650), .B(n3649), .Z(\round_in[0][499] ) );
  NAND U9553 ( .A(init), .B(round_reg[49]), .Z(n3652) );
  NANDN U9554 ( .A(init), .B(in[49]), .Z(n3651) );
  NAND U9555 ( .A(n3652), .B(n3651), .Z(\round_in[0][49] ) );
  NAND U9556 ( .A(init), .B(round_reg[4]), .Z(n3654) );
  NANDN U9557 ( .A(init), .B(in[4]), .Z(n3653) );
  NAND U9558 ( .A(n3654), .B(n3653), .Z(\round_in[0][4] ) );
  NAND U9559 ( .A(init), .B(round_reg[500]), .Z(n3656) );
  NANDN U9560 ( .A(init), .B(in[500]), .Z(n3655) );
  NAND U9561 ( .A(n3656), .B(n3655), .Z(\round_in[0][500] ) );
  NAND U9562 ( .A(init), .B(round_reg[501]), .Z(n3658) );
  NANDN U9563 ( .A(init), .B(in[501]), .Z(n3657) );
  NAND U9564 ( .A(n3658), .B(n3657), .Z(\round_in[0][501] ) );
  NAND U9565 ( .A(init), .B(round_reg[502]), .Z(n3660) );
  NANDN U9566 ( .A(init), .B(in[502]), .Z(n3659) );
  NAND U9567 ( .A(n3660), .B(n3659), .Z(\round_in[0][502] ) );
  NAND U9568 ( .A(init), .B(round_reg[503]), .Z(n3662) );
  NANDN U9569 ( .A(init), .B(in[503]), .Z(n3661) );
  NAND U9570 ( .A(n3662), .B(n3661), .Z(\round_in[0][503] ) );
  NAND U9571 ( .A(init), .B(round_reg[504]), .Z(n3664) );
  NANDN U9572 ( .A(init), .B(in[504]), .Z(n3663) );
  NAND U9573 ( .A(n3664), .B(n3663), .Z(\round_in[0][504] ) );
  NAND U9574 ( .A(init), .B(round_reg[505]), .Z(n3666) );
  NANDN U9575 ( .A(init), .B(in[505]), .Z(n3665) );
  NAND U9576 ( .A(n3666), .B(n3665), .Z(\round_in[0][505] ) );
  NAND U9577 ( .A(init), .B(round_reg[506]), .Z(n3668) );
  NANDN U9578 ( .A(init), .B(in[506]), .Z(n3667) );
  NAND U9579 ( .A(n3668), .B(n3667), .Z(\round_in[0][506] ) );
  NAND U9580 ( .A(init), .B(round_reg[507]), .Z(n3670) );
  NANDN U9581 ( .A(init), .B(in[507]), .Z(n3669) );
  NAND U9582 ( .A(n3670), .B(n3669), .Z(\round_in[0][507] ) );
  NAND U9583 ( .A(init), .B(round_reg[508]), .Z(n3672) );
  NANDN U9584 ( .A(init), .B(in[508]), .Z(n3671) );
  NAND U9585 ( .A(n3672), .B(n3671), .Z(\round_in[0][508] ) );
  NAND U9586 ( .A(init), .B(round_reg[509]), .Z(n3674) );
  NANDN U9587 ( .A(init), .B(in[509]), .Z(n3673) );
  NAND U9588 ( .A(n3674), .B(n3673), .Z(\round_in[0][509] ) );
  NAND U9589 ( .A(init), .B(round_reg[50]), .Z(n3676) );
  NANDN U9590 ( .A(init), .B(in[50]), .Z(n3675) );
  NAND U9591 ( .A(n3676), .B(n3675), .Z(\round_in[0][50] ) );
  NAND U9592 ( .A(init), .B(round_reg[510]), .Z(n3678) );
  NANDN U9593 ( .A(init), .B(in[510]), .Z(n3677) );
  NAND U9594 ( .A(n3678), .B(n3677), .Z(\round_in[0][510] ) );
  NAND U9595 ( .A(init), .B(round_reg[511]), .Z(n3680) );
  NANDN U9596 ( .A(init), .B(in[511]), .Z(n3679) );
  NAND U9597 ( .A(n3680), .B(n3679), .Z(\round_in[0][511] ) );
  NAND U9598 ( .A(init), .B(round_reg[512]), .Z(n3682) );
  NANDN U9599 ( .A(init), .B(in[512]), .Z(n3681) );
  NAND U9600 ( .A(n3682), .B(n3681), .Z(\round_in[0][512] ) );
  NAND U9601 ( .A(init), .B(round_reg[513]), .Z(n3684) );
  NANDN U9602 ( .A(init), .B(in[513]), .Z(n3683) );
  NAND U9603 ( .A(n3684), .B(n3683), .Z(\round_in[0][513] ) );
  NAND U9604 ( .A(init), .B(round_reg[514]), .Z(n3686) );
  NANDN U9605 ( .A(init), .B(in[514]), .Z(n3685) );
  NAND U9606 ( .A(n3686), .B(n3685), .Z(\round_in[0][514] ) );
  NAND U9607 ( .A(init), .B(round_reg[515]), .Z(n3688) );
  NANDN U9608 ( .A(init), .B(in[515]), .Z(n3687) );
  NAND U9609 ( .A(n3688), .B(n3687), .Z(\round_in[0][515] ) );
  NAND U9610 ( .A(init), .B(round_reg[516]), .Z(n3690) );
  NANDN U9611 ( .A(init), .B(in[516]), .Z(n3689) );
  NAND U9612 ( .A(n3690), .B(n3689), .Z(\round_in[0][516] ) );
  NAND U9613 ( .A(init), .B(round_reg[517]), .Z(n3692) );
  NANDN U9614 ( .A(init), .B(in[517]), .Z(n3691) );
  NAND U9615 ( .A(n3692), .B(n3691), .Z(\round_in[0][517] ) );
  NAND U9616 ( .A(init), .B(round_reg[518]), .Z(n3694) );
  NANDN U9617 ( .A(init), .B(in[518]), .Z(n3693) );
  NAND U9618 ( .A(n3694), .B(n3693), .Z(\round_in[0][518] ) );
  NAND U9619 ( .A(init), .B(round_reg[519]), .Z(n3696) );
  NANDN U9620 ( .A(init), .B(in[519]), .Z(n3695) );
  NAND U9621 ( .A(n3696), .B(n3695), .Z(\round_in[0][519] ) );
  NAND U9622 ( .A(init), .B(round_reg[51]), .Z(n3698) );
  NANDN U9623 ( .A(init), .B(in[51]), .Z(n3697) );
  NAND U9624 ( .A(n3698), .B(n3697), .Z(\round_in[0][51] ) );
  NAND U9625 ( .A(init), .B(round_reg[520]), .Z(n3700) );
  NANDN U9626 ( .A(init), .B(in[520]), .Z(n3699) );
  NAND U9627 ( .A(n3700), .B(n3699), .Z(\round_in[0][520] ) );
  NAND U9628 ( .A(init), .B(round_reg[521]), .Z(n3702) );
  NANDN U9629 ( .A(init), .B(in[521]), .Z(n3701) );
  NAND U9630 ( .A(n3702), .B(n3701), .Z(\round_in[0][521] ) );
  NAND U9631 ( .A(init), .B(round_reg[522]), .Z(n3704) );
  NANDN U9632 ( .A(init), .B(in[522]), .Z(n3703) );
  NAND U9633 ( .A(n3704), .B(n3703), .Z(\round_in[0][522] ) );
  NAND U9634 ( .A(init), .B(round_reg[523]), .Z(n3706) );
  NANDN U9635 ( .A(init), .B(in[523]), .Z(n3705) );
  NAND U9636 ( .A(n3706), .B(n3705), .Z(\round_in[0][523] ) );
  NAND U9637 ( .A(init), .B(round_reg[524]), .Z(n3708) );
  NANDN U9638 ( .A(init), .B(in[524]), .Z(n3707) );
  NAND U9639 ( .A(n3708), .B(n3707), .Z(\round_in[0][524] ) );
  NAND U9640 ( .A(init), .B(round_reg[525]), .Z(n3710) );
  NANDN U9641 ( .A(init), .B(in[525]), .Z(n3709) );
  NAND U9642 ( .A(n3710), .B(n3709), .Z(\round_in[0][525] ) );
  NAND U9643 ( .A(init), .B(round_reg[526]), .Z(n3712) );
  NANDN U9644 ( .A(init), .B(in[526]), .Z(n3711) );
  NAND U9645 ( .A(n3712), .B(n3711), .Z(\round_in[0][526] ) );
  NAND U9646 ( .A(init), .B(round_reg[527]), .Z(n3714) );
  NANDN U9647 ( .A(init), .B(in[527]), .Z(n3713) );
  NAND U9648 ( .A(n3714), .B(n3713), .Z(\round_in[0][527] ) );
  NAND U9649 ( .A(init), .B(round_reg[528]), .Z(n3716) );
  NANDN U9650 ( .A(init), .B(in[528]), .Z(n3715) );
  NAND U9651 ( .A(n3716), .B(n3715), .Z(\round_in[0][528] ) );
  NAND U9652 ( .A(init), .B(round_reg[529]), .Z(n3718) );
  NANDN U9653 ( .A(init), .B(in[529]), .Z(n3717) );
  NAND U9654 ( .A(n3718), .B(n3717), .Z(\round_in[0][529] ) );
  NAND U9655 ( .A(init), .B(round_reg[52]), .Z(n3720) );
  NANDN U9656 ( .A(init), .B(in[52]), .Z(n3719) );
  NAND U9657 ( .A(n3720), .B(n3719), .Z(\round_in[0][52] ) );
  NAND U9658 ( .A(init), .B(round_reg[530]), .Z(n3722) );
  NANDN U9659 ( .A(init), .B(in[530]), .Z(n3721) );
  NAND U9660 ( .A(n3722), .B(n3721), .Z(\round_in[0][530] ) );
  NAND U9661 ( .A(init), .B(round_reg[531]), .Z(n3724) );
  NANDN U9662 ( .A(init), .B(in[531]), .Z(n3723) );
  NAND U9663 ( .A(n3724), .B(n3723), .Z(\round_in[0][531] ) );
  NAND U9664 ( .A(init), .B(round_reg[532]), .Z(n3726) );
  NANDN U9665 ( .A(init), .B(in[532]), .Z(n3725) );
  NAND U9666 ( .A(n3726), .B(n3725), .Z(\round_in[0][532] ) );
  NAND U9667 ( .A(init), .B(round_reg[533]), .Z(n3728) );
  NANDN U9668 ( .A(init), .B(in[533]), .Z(n3727) );
  NAND U9669 ( .A(n3728), .B(n3727), .Z(\round_in[0][533] ) );
  NAND U9670 ( .A(init), .B(round_reg[534]), .Z(n3730) );
  NANDN U9671 ( .A(init), .B(in[534]), .Z(n3729) );
  NAND U9672 ( .A(n3730), .B(n3729), .Z(\round_in[0][534] ) );
  NAND U9673 ( .A(init), .B(round_reg[535]), .Z(n3732) );
  NANDN U9674 ( .A(init), .B(in[535]), .Z(n3731) );
  NAND U9675 ( .A(n3732), .B(n3731), .Z(\round_in[0][535] ) );
  NAND U9676 ( .A(init), .B(round_reg[536]), .Z(n3734) );
  NANDN U9677 ( .A(init), .B(in[536]), .Z(n3733) );
  NAND U9678 ( .A(n3734), .B(n3733), .Z(\round_in[0][536] ) );
  NAND U9679 ( .A(init), .B(round_reg[537]), .Z(n3736) );
  NANDN U9680 ( .A(init), .B(in[537]), .Z(n3735) );
  NAND U9681 ( .A(n3736), .B(n3735), .Z(\round_in[0][537] ) );
  NAND U9682 ( .A(init), .B(round_reg[538]), .Z(n3738) );
  NANDN U9683 ( .A(init), .B(in[538]), .Z(n3737) );
  NAND U9684 ( .A(n3738), .B(n3737), .Z(\round_in[0][538] ) );
  NAND U9685 ( .A(init), .B(round_reg[539]), .Z(n3740) );
  NANDN U9686 ( .A(init), .B(in[539]), .Z(n3739) );
  NAND U9687 ( .A(n3740), .B(n3739), .Z(\round_in[0][539] ) );
  NAND U9688 ( .A(init), .B(round_reg[53]), .Z(n3742) );
  NANDN U9689 ( .A(init), .B(in[53]), .Z(n3741) );
  NAND U9690 ( .A(n3742), .B(n3741), .Z(\round_in[0][53] ) );
  NAND U9691 ( .A(init), .B(round_reg[540]), .Z(n3744) );
  NANDN U9692 ( .A(init), .B(in[540]), .Z(n3743) );
  NAND U9693 ( .A(n3744), .B(n3743), .Z(\round_in[0][540] ) );
  NAND U9694 ( .A(init), .B(round_reg[541]), .Z(n3746) );
  NANDN U9695 ( .A(init), .B(in[541]), .Z(n3745) );
  NAND U9696 ( .A(n3746), .B(n3745), .Z(\round_in[0][541] ) );
  NAND U9697 ( .A(init), .B(round_reg[542]), .Z(n3748) );
  NANDN U9698 ( .A(init), .B(in[542]), .Z(n3747) );
  NAND U9699 ( .A(n3748), .B(n3747), .Z(\round_in[0][542] ) );
  NAND U9700 ( .A(init), .B(round_reg[543]), .Z(n3750) );
  NANDN U9701 ( .A(init), .B(in[543]), .Z(n3749) );
  NAND U9702 ( .A(n3750), .B(n3749), .Z(\round_in[0][543] ) );
  NAND U9703 ( .A(init), .B(round_reg[544]), .Z(n3752) );
  NANDN U9704 ( .A(init), .B(in[544]), .Z(n3751) );
  NAND U9705 ( .A(n3752), .B(n3751), .Z(\round_in[0][544] ) );
  NAND U9706 ( .A(init), .B(round_reg[545]), .Z(n3754) );
  NANDN U9707 ( .A(init), .B(in[545]), .Z(n3753) );
  NAND U9708 ( .A(n3754), .B(n3753), .Z(\round_in[0][545] ) );
  NAND U9709 ( .A(init), .B(round_reg[546]), .Z(n3756) );
  NANDN U9710 ( .A(init), .B(in[546]), .Z(n3755) );
  NAND U9711 ( .A(n3756), .B(n3755), .Z(\round_in[0][546] ) );
  NAND U9712 ( .A(init), .B(round_reg[547]), .Z(n3758) );
  NANDN U9713 ( .A(init), .B(in[547]), .Z(n3757) );
  NAND U9714 ( .A(n3758), .B(n3757), .Z(\round_in[0][547] ) );
  NAND U9715 ( .A(init), .B(round_reg[548]), .Z(n3760) );
  NANDN U9716 ( .A(init), .B(in[548]), .Z(n3759) );
  NAND U9717 ( .A(n3760), .B(n3759), .Z(\round_in[0][548] ) );
  NAND U9718 ( .A(init), .B(round_reg[549]), .Z(n3762) );
  NANDN U9719 ( .A(init), .B(in[549]), .Z(n3761) );
  NAND U9720 ( .A(n3762), .B(n3761), .Z(\round_in[0][549] ) );
  NAND U9721 ( .A(init), .B(round_reg[54]), .Z(n3764) );
  NANDN U9722 ( .A(init), .B(in[54]), .Z(n3763) );
  NAND U9723 ( .A(n3764), .B(n3763), .Z(\round_in[0][54] ) );
  NAND U9724 ( .A(init), .B(round_reg[550]), .Z(n3766) );
  NANDN U9725 ( .A(init), .B(in[550]), .Z(n3765) );
  NAND U9726 ( .A(n3766), .B(n3765), .Z(\round_in[0][550] ) );
  NAND U9727 ( .A(init), .B(round_reg[551]), .Z(n3768) );
  NANDN U9728 ( .A(init), .B(in[551]), .Z(n3767) );
  NAND U9729 ( .A(n3768), .B(n3767), .Z(\round_in[0][551] ) );
  NAND U9730 ( .A(init), .B(round_reg[552]), .Z(n3770) );
  NANDN U9731 ( .A(init), .B(in[552]), .Z(n3769) );
  NAND U9732 ( .A(n3770), .B(n3769), .Z(\round_in[0][552] ) );
  NAND U9733 ( .A(init), .B(round_reg[553]), .Z(n3772) );
  NANDN U9734 ( .A(init), .B(in[553]), .Z(n3771) );
  NAND U9735 ( .A(n3772), .B(n3771), .Z(\round_in[0][553] ) );
  NAND U9736 ( .A(init), .B(round_reg[554]), .Z(n3774) );
  NANDN U9737 ( .A(init), .B(in[554]), .Z(n3773) );
  NAND U9738 ( .A(n3774), .B(n3773), .Z(\round_in[0][554] ) );
  NAND U9739 ( .A(init), .B(round_reg[555]), .Z(n3776) );
  NANDN U9740 ( .A(init), .B(in[555]), .Z(n3775) );
  NAND U9741 ( .A(n3776), .B(n3775), .Z(\round_in[0][555] ) );
  NAND U9742 ( .A(init), .B(round_reg[556]), .Z(n3778) );
  NANDN U9743 ( .A(init), .B(in[556]), .Z(n3777) );
  NAND U9744 ( .A(n3778), .B(n3777), .Z(\round_in[0][556] ) );
  NAND U9745 ( .A(init), .B(round_reg[557]), .Z(n3780) );
  NANDN U9746 ( .A(init), .B(in[557]), .Z(n3779) );
  NAND U9747 ( .A(n3780), .B(n3779), .Z(\round_in[0][557] ) );
  NAND U9748 ( .A(init), .B(round_reg[558]), .Z(n3782) );
  NANDN U9749 ( .A(init), .B(in[558]), .Z(n3781) );
  NAND U9750 ( .A(n3782), .B(n3781), .Z(\round_in[0][558] ) );
  NAND U9751 ( .A(init), .B(round_reg[559]), .Z(n3784) );
  NANDN U9752 ( .A(init), .B(in[559]), .Z(n3783) );
  NAND U9753 ( .A(n3784), .B(n3783), .Z(\round_in[0][559] ) );
  NAND U9754 ( .A(init), .B(round_reg[55]), .Z(n3786) );
  NANDN U9755 ( .A(init), .B(in[55]), .Z(n3785) );
  NAND U9756 ( .A(n3786), .B(n3785), .Z(\round_in[0][55] ) );
  NAND U9757 ( .A(init), .B(round_reg[560]), .Z(n3788) );
  NANDN U9758 ( .A(init), .B(in[560]), .Z(n3787) );
  NAND U9759 ( .A(n3788), .B(n3787), .Z(\round_in[0][560] ) );
  NAND U9760 ( .A(init), .B(round_reg[561]), .Z(n3790) );
  NANDN U9761 ( .A(init), .B(in[561]), .Z(n3789) );
  NAND U9762 ( .A(n3790), .B(n3789), .Z(\round_in[0][561] ) );
  NAND U9763 ( .A(init), .B(round_reg[562]), .Z(n3792) );
  NANDN U9764 ( .A(init), .B(in[562]), .Z(n3791) );
  NAND U9765 ( .A(n3792), .B(n3791), .Z(\round_in[0][562] ) );
  NAND U9766 ( .A(init), .B(round_reg[563]), .Z(n3794) );
  NANDN U9767 ( .A(init), .B(in[563]), .Z(n3793) );
  NAND U9768 ( .A(n3794), .B(n3793), .Z(\round_in[0][563] ) );
  NAND U9769 ( .A(init), .B(round_reg[564]), .Z(n3796) );
  NANDN U9770 ( .A(init), .B(in[564]), .Z(n3795) );
  NAND U9771 ( .A(n3796), .B(n3795), .Z(\round_in[0][564] ) );
  NAND U9772 ( .A(init), .B(round_reg[565]), .Z(n3798) );
  NANDN U9773 ( .A(init), .B(in[565]), .Z(n3797) );
  NAND U9774 ( .A(n3798), .B(n3797), .Z(\round_in[0][565] ) );
  NAND U9775 ( .A(init), .B(round_reg[566]), .Z(n3800) );
  NANDN U9776 ( .A(init), .B(in[566]), .Z(n3799) );
  NAND U9777 ( .A(n3800), .B(n3799), .Z(\round_in[0][566] ) );
  NAND U9778 ( .A(init), .B(round_reg[567]), .Z(n3802) );
  NANDN U9779 ( .A(init), .B(in[567]), .Z(n3801) );
  NAND U9780 ( .A(n3802), .B(n3801), .Z(\round_in[0][567] ) );
  NAND U9781 ( .A(init), .B(round_reg[568]), .Z(n3804) );
  NANDN U9782 ( .A(init), .B(in[568]), .Z(n3803) );
  NAND U9783 ( .A(n3804), .B(n3803), .Z(\round_in[0][568] ) );
  NAND U9784 ( .A(init), .B(round_reg[569]), .Z(n3806) );
  NANDN U9785 ( .A(init), .B(in[569]), .Z(n3805) );
  NAND U9786 ( .A(n3806), .B(n3805), .Z(\round_in[0][569] ) );
  NAND U9787 ( .A(init), .B(round_reg[56]), .Z(n3808) );
  NANDN U9788 ( .A(init), .B(in[56]), .Z(n3807) );
  NAND U9789 ( .A(n3808), .B(n3807), .Z(\round_in[0][56] ) );
  NAND U9790 ( .A(init), .B(round_reg[570]), .Z(n3810) );
  NANDN U9791 ( .A(init), .B(in[570]), .Z(n3809) );
  NAND U9792 ( .A(n3810), .B(n3809), .Z(\round_in[0][570] ) );
  NAND U9793 ( .A(init), .B(round_reg[571]), .Z(n3812) );
  NANDN U9794 ( .A(init), .B(in[571]), .Z(n3811) );
  NAND U9795 ( .A(n3812), .B(n3811), .Z(\round_in[0][571] ) );
  NAND U9796 ( .A(init), .B(round_reg[572]), .Z(n3814) );
  NANDN U9797 ( .A(init), .B(in[572]), .Z(n3813) );
  NAND U9798 ( .A(n3814), .B(n3813), .Z(\round_in[0][572] ) );
  NAND U9799 ( .A(init), .B(round_reg[573]), .Z(n3816) );
  NANDN U9800 ( .A(init), .B(in[573]), .Z(n3815) );
  NAND U9801 ( .A(n3816), .B(n3815), .Z(\round_in[0][573] ) );
  NAND U9802 ( .A(init), .B(round_reg[574]), .Z(n3818) );
  NANDN U9803 ( .A(init), .B(in[574]), .Z(n3817) );
  NAND U9804 ( .A(n3818), .B(n3817), .Z(\round_in[0][574] ) );
  NAND U9805 ( .A(init), .B(round_reg[575]), .Z(n3820) );
  NANDN U9806 ( .A(init), .B(in[575]), .Z(n3819) );
  NAND U9807 ( .A(n3820), .B(n3819), .Z(\round_in[0][575] ) );
  AND U9808 ( .A(round_reg[576]), .B(init), .Z(\round_in[0][576] ) );
  AND U9809 ( .A(round_reg[577]), .B(init), .Z(\round_in[0][577] ) );
  AND U9810 ( .A(round_reg[578]), .B(init), .Z(\round_in[0][578] ) );
  AND U9811 ( .A(round_reg[579]), .B(init), .Z(\round_in[0][579] ) );
  NAND U9812 ( .A(init), .B(round_reg[57]), .Z(n3822) );
  NANDN U9813 ( .A(init), .B(in[57]), .Z(n3821) );
  NAND U9814 ( .A(n3822), .B(n3821), .Z(\round_in[0][57] ) );
  AND U9815 ( .A(round_reg[580]), .B(init), .Z(\round_in[0][580] ) );
  AND U9816 ( .A(round_reg[581]), .B(init), .Z(\round_in[0][581] ) );
  AND U9817 ( .A(round_reg[582]), .B(init), .Z(\round_in[0][582] ) );
  AND U9818 ( .A(round_reg[583]), .B(init), .Z(\round_in[0][583] ) );
  AND U9819 ( .A(round_reg[584]), .B(init), .Z(\round_in[0][584] ) );
  AND U9820 ( .A(round_reg[585]), .B(init), .Z(\round_in[0][585] ) );
  AND U9821 ( .A(round_reg[586]), .B(init), .Z(\round_in[0][586] ) );
  AND U9822 ( .A(round_reg[587]), .B(init), .Z(\round_in[0][587] ) );
  AND U9823 ( .A(round_reg[588]), .B(init), .Z(\round_in[0][588] ) );
  AND U9824 ( .A(round_reg[589]), .B(init), .Z(\round_in[0][589] ) );
  NAND U9825 ( .A(init), .B(round_reg[58]), .Z(n3824) );
  NANDN U9826 ( .A(init), .B(in[58]), .Z(n3823) );
  NAND U9827 ( .A(n3824), .B(n3823), .Z(\round_in[0][58] ) );
  AND U9828 ( .A(round_reg[590]), .B(init), .Z(\round_in[0][590] ) );
  AND U9829 ( .A(round_reg[591]), .B(init), .Z(\round_in[0][591] ) );
  AND U9830 ( .A(round_reg[592]), .B(init), .Z(\round_in[0][592] ) );
  AND U9831 ( .A(round_reg[593]), .B(init), .Z(\round_in[0][593] ) );
  AND U9832 ( .A(round_reg[594]), .B(init), .Z(\round_in[0][594] ) );
  AND U9833 ( .A(round_reg[595]), .B(init), .Z(\round_in[0][595] ) );
  AND U9834 ( .A(round_reg[596]), .B(init), .Z(\round_in[0][596] ) );
  AND U9835 ( .A(round_reg[597]), .B(init), .Z(\round_in[0][597] ) );
  AND U9836 ( .A(round_reg[598]), .B(init), .Z(\round_in[0][598] ) );
  AND U9837 ( .A(round_reg[599]), .B(init), .Z(\round_in[0][599] ) );
  NAND U9838 ( .A(init), .B(round_reg[59]), .Z(n3826) );
  NANDN U9839 ( .A(init), .B(in[59]), .Z(n3825) );
  NAND U9840 ( .A(n3826), .B(n3825), .Z(\round_in[0][59] ) );
  NAND U9841 ( .A(init), .B(round_reg[5]), .Z(n3828) );
  NANDN U9842 ( .A(init), .B(in[5]), .Z(n3827) );
  NAND U9843 ( .A(n3828), .B(n3827), .Z(\round_in[0][5] ) );
  AND U9844 ( .A(round_reg[600]), .B(init), .Z(\round_in[0][600] ) );
  AND U9845 ( .A(round_reg[601]), .B(init), .Z(\round_in[0][601] ) );
  AND U9846 ( .A(round_reg[602]), .B(init), .Z(\round_in[0][602] ) );
  AND U9847 ( .A(round_reg[603]), .B(init), .Z(\round_in[0][603] ) );
  AND U9848 ( .A(round_reg[604]), .B(init), .Z(\round_in[0][604] ) );
  AND U9849 ( .A(round_reg[605]), .B(init), .Z(\round_in[0][605] ) );
  AND U9850 ( .A(round_reg[606]), .B(init), .Z(\round_in[0][606] ) );
  AND U9851 ( .A(round_reg[607]), .B(init), .Z(\round_in[0][607] ) );
  AND U9852 ( .A(round_reg[608]), .B(init), .Z(\round_in[0][608] ) );
  AND U9853 ( .A(round_reg[609]), .B(init), .Z(\round_in[0][609] ) );
  NAND U9854 ( .A(init), .B(round_reg[60]), .Z(n3830) );
  NANDN U9855 ( .A(init), .B(in[60]), .Z(n3829) );
  NAND U9856 ( .A(n3830), .B(n3829), .Z(\round_in[0][60] ) );
  AND U9857 ( .A(round_reg[610]), .B(init), .Z(\round_in[0][610] ) );
  AND U9858 ( .A(round_reg[611]), .B(init), .Z(\round_in[0][611] ) );
  AND U9859 ( .A(round_reg[612]), .B(init), .Z(\round_in[0][612] ) );
  AND U9860 ( .A(round_reg[613]), .B(init), .Z(\round_in[0][613] ) );
  AND U9861 ( .A(round_reg[614]), .B(init), .Z(\round_in[0][614] ) );
  AND U9862 ( .A(round_reg[615]), .B(init), .Z(\round_in[0][615] ) );
  AND U9863 ( .A(round_reg[616]), .B(init), .Z(\round_in[0][616] ) );
  AND U9864 ( .A(round_reg[617]), .B(init), .Z(\round_in[0][617] ) );
  AND U9865 ( .A(round_reg[618]), .B(init), .Z(\round_in[0][618] ) );
  AND U9866 ( .A(round_reg[619]), .B(init), .Z(\round_in[0][619] ) );
  NAND U9867 ( .A(init), .B(round_reg[61]), .Z(n3832) );
  NANDN U9868 ( .A(init), .B(in[61]), .Z(n3831) );
  NAND U9869 ( .A(n3832), .B(n3831), .Z(\round_in[0][61] ) );
  AND U9870 ( .A(round_reg[620]), .B(init), .Z(\round_in[0][620] ) );
  AND U9871 ( .A(round_reg[621]), .B(init), .Z(\round_in[0][621] ) );
  AND U9872 ( .A(round_reg[622]), .B(init), .Z(\round_in[0][622] ) );
  AND U9873 ( .A(round_reg[623]), .B(init), .Z(\round_in[0][623] ) );
  AND U9874 ( .A(round_reg[624]), .B(init), .Z(\round_in[0][624] ) );
  AND U9875 ( .A(round_reg[625]), .B(init), .Z(\round_in[0][625] ) );
  AND U9876 ( .A(round_reg[626]), .B(init), .Z(\round_in[0][626] ) );
  AND U9877 ( .A(round_reg[627]), .B(init), .Z(\round_in[0][627] ) );
  AND U9878 ( .A(round_reg[628]), .B(init), .Z(\round_in[0][628] ) );
  AND U9879 ( .A(round_reg[629]), .B(init), .Z(\round_in[0][629] ) );
  NAND U9880 ( .A(init), .B(round_reg[62]), .Z(n3834) );
  NANDN U9881 ( .A(init), .B(in[62]), .Z(n3833) );
  NAND U9882 ( .A(n3834), .B(n3833), .Z(\round_in[0][62] ) );
  AND U9883 ( .A(round_reg[630]), .B(init), .Z(\round_in[0][630] ) );
  AND U9884 ( .A(round_reg[631]), .B(init), .Z(\round_in[0][631] ) );
  AND U9885 ( .A(round_reg[632]), .B(init), .Z(\round_in[0][632] ) );
  AND U9886 ( .A(round_reg[633]), .B(init), .Z(\round_in[0][633] ) );
  AND U9887 ( .A(round_reg[634]), .B(init), .Z(\round_in[0][634] ) );
  AND U9888 ( .A(round_reg[635]), .B(init), .Z(\round_in[0][635] ) );
  AND U9889 ( .A(round_reg[636]), .B(init), .Z(\round_in[0][636] ) );
  AND U9890 ( .A(round_reg[637]), .B(init), .Z(\round_in[0][637] ) );
  AND U9891 ( .A(round_reg[638]), .B(init), .Z(\round_in[0][638] ) );
  AND U9892 ( .A(round_reg[639]), .B(init), .Z(\round_in[0][639] ) );
  NAND U9893 ( .A(init), .B(round_reg[63]), .Z(n3836) );
  NANDN U9894 ( .A(init), .B(in[63]), .Z(n3835) );
  NAND U9895 ( .A(n3836), .B(n3835), .Z(\round_in[0][63] ) );
  AND U9896 ( .A(round_reg[640]), .B(init), .Z(\round_in[0][640] ) );
  AND U9897 ( .A(round_reg[641]), .B(init), .Z(\round_in[0][641] ) );
  AND U9898 ( .A(round_reg[642]), .B(init), .Z(\round_in[0][642] ) );
  AND U9899 ( .A(round_reg[643]), .B(init), .Z(\round_in[0][643] ) );
  AND U9900 ( .A(round_reg[644]), .B(init), .Z(\round_in[0][644] ) );
  AND U9901 ( .A(round_reg[645]), .B(init), .Z(\round_in[0][645] ) );
  AND U9902 ( .A(round_reg[646]), .B(init), .Z(\round_in[0][646] ) );
  AND U9903 ( .A(round_reg[647]), .B(init), .Z(\round_in[0][647] ) );
  AND U9904 ( .A(round_reg[648]), .B(init), .Z(\round_in[0][648] ) );
  AND U9905 ( .A(round_reg[649]), .B(init), .Z(\round_in[0][649] ) );
  NAND U9906 ( .A(init), .B(round_reg[64]), .Z(n3838) );
  NANDN U9907 ( .A(init), .B(in[64]), .Z(n3837) );
  NAND U9908 ( .A(n3838), .B(n3837), .Z(\round_in[0][64] ) );
  AND U9909 ( .A(round_reg[650]), .B(init), .Z(\round_in[0][650] ) );
  AND U9910 ( .A(round_reg[651]), .B(init), .Z(\round_in[0][651] ) );
  AND U9911 ( .A(round_reg[652]), .B(init), .Z(\round_in[0][652] ) );
  AND U9912 ( .A(round_reg[653]), .B(init), .Z(\round_in[0][653] ) );
  AND U9913 ( .A(round_reg[654]), .B(init), .Z(\round_in[0][654] ) );
  AND U9914 ( .A(round_reg[655]), .B(init), .Z(\round_in[0][655] ) );
  AND U9915 ( .A(round_reg[656]), .B(init), .Z(\round_in[0][656] ) );
  AND U9916 ( .A(round_reg[657]), .B(init), .Z(\round_in[0][657] ) );
  AND U9917 ( .A(round_reg[658]), .B(init), .Z(\round_in[0][658] ) );
  AND U9918 ( .A(round_reg[659]), .B(init), .Z(\round_in[0][659] ) );
  NAND U9919 ( .A(init), .B(round_reg[65]), .Z(n3840) );
  NANDN U9920 ( .A(init), .B(in[65]), .Z(n3839) );
  NAND U9921 ( .A(n3840), .B(n3839), .Z(\round_in[0][65] ) );
  AND U9922 ( .A(round_reg[660]), .B(init), .Z(\round_in[0][660] ) );
  AND U9923 ( .A(round_reg[661]), .B(init), .Z(\round_in[0][661] ) );
  AND U9924 ( .A(round_reg[662]), .B(init), .Z(\round_in[0][662] ) );
  AND U9925 ( .A(round_reg[663]), .B(init), .Z(\round_in[0][663] ) );
  AND U9926 ( .A(round_reg[664]), .B(init), .Z(\round_in[0][664] ) );
  AND U9927 ( .A(round_reg[665]), .B(init), .Z(\round_in[0][665] ) );
  AND U9928 ( .A(round_reg[666]), .B(init), .Z(\round_in[0][666] ) );
  AND U9929 ( .A(round_reg[667]), .B(init), .Z(\round_in[0][667] ) );
  AND U9930 ( .A(round_reg[668]), .B(init), .Z(\round_in[0][668] ) );
  AND U9931 ( .A(round_reg[669]), .B(init), .Z(\round_in[0][669] ) );
  NAND U9932 ( .A(init), .B(round_reg[66]), .Z(n3842) );
  NANDN U9933 ( .A(init), .B(in[66]), .Z(n3841) );
  NAND U9934 ( .A(n3842), .B(n3841), .Z(\round_in[0][66] ) );
  AND U9935 ( .A(round_reg[670]), .B(init), .Z(\round_in[0][670] ) );
  AND U9936 ( .A(round_reg[671]), .B(init), .Z(\round_in[0][671] ) );
  AND U9937 ( .A(round_reg[672]), .B(init), .Z(\round_in[0][672] ) );
  AND U9938 ( .A(round_reg[673]), .B(init), .Z(\round_in[0][673] ) );
  AND U9939 ( .A(round_reg[674]), .B(init), .Z(\round_in[0][674] ) );
  AND U9940 ( .A(round_reg[675]), .B(init), .Z(\round_in[0][675] ) );
  AND U9941 ( .A(round_reg[676]), .B(init), .Z(\round_in[0][676] ) );
  AND U9942 ( .A(round_reg[677]), .B(init), .Z(\round_in[0][677] ) );
  AND U9943 ( .A(round_reg[678]), .B(init), .Z(\round_in[0][678] ) );
  AND U9944 ( .A(round_reg[679]), .B(init), .Z(\round_in[0][679] ) );
  NAND U9945 ( .A(init), .B(round_reg[67]), .Z(n3844) );
  NANDN U9946 ( .A(init), .B(in[67]), .Z(n3843) );
  NAND U9947 ( .A(n3844), .B(n3843), .Z(\round_in[0][67] ) );
  AND U9948 ( .A(round_reg[680]), .B(init), .Z(\round_in[0][680] ) );
  AND U9949 ( .A(round_reg[681]), .B(init), .Z(\round_in[0][681] ) );
  AND U9950 ( .A(round_reg[682]), .B(init), .Z(\round_in[0][682] ) );
  AND U9951 ( .A(round_reg[683]), .B(init), .Z(\round_in[0][683] ) );
  AND U9952 ( .A(round_reg[684]), .B(init), .Z(\round_in[0][684] ) );
  AND U9953 ( .A(round_reg[685]), .B(init), .Z(\round_in[0][685] ) );
  AND U9954 ( .A(round_reg[686]), .B(init), .Z(\round_in[0][686] ) );
  AND U9955 ( .A(round_reg[687]), .B(init), .Z(\round_in[0][687] ) );
  AND U9956 ( .A(round_reg[688]), .B(init), .Z(\round_in[0][688] ) );
  AND U9957 ( .A(round_reg[689]), .B(init), .Z(\round_in[0][689] ) );
  NAND U9958 ( .A(init), .B(round_reg[68]), .Z(n3846) );
  NANDN U9959 ( .A(init), .B(in[68]), .Z(n3845) );
  NAND U9960 ( .A(n3846), .B(n3845), .Z(\round_in[0][68] ) );
  AND U9961 ( .A(round_reg[690]), .B(init), .Z(\round_in[0][690] ) );
  AND U9962 ( .A(round_reg[691]), .B(init), .Z(\round_in[0][691] ) );
  AND U9963 ( .A(round_reg[692]), .B(init), .Z(\round_in[0][692] ) );
  AND U9964 ( .A(round_reg[693]), .B(init), .Z(\round_in[0][693] ) );
  AND U9965 ( .A(round_reg[694]), .B(init), .Z(\round_in[0][694] ) );
  AND U9966 ( .A(round_reg[695]), .B(init), .Z(\round_in[0][695] ) );
  AND U9967 ( .A(round_reg[696]), .B(init), .Z(\round_in[0][696] ) );
  AND U9968 ( .A(round_reg[697]), .B(init), .Z(\round_in[0][697] ) );
  AND U9969 ( .A(round_reg[698]), .B(init), .Z(\round_in[0][698] ) );
  AND U9970 ( .A(round_reg[699]), .B(init), .Z(\round_in[0][699] ) );
  NAND U9971 ( .A(init), .B(round_reg[69]), .Z(n3848) );
  NANDN U9972 ( .A(init), .B(in[69]), .Z(n3847) );
  NAND U9973 ( .A(n3848), .B(n3847), .Z(\round_in[0][69] ) );
  NAND U9974 ( .A(init), .B(round_reg[6]), .Z(n3850) );
  NANDN U9975 ( .A(init), .B(in[6]), .Z(n3849) );
  NAND U9976 ( .A(n3850), .B(n3849), .Z(\round_in[0][6] ) );
  AND U9977 ( .A(round_reg[700]), .B(init), .Z(\round_in[0][700] ) );
  AND U9978 ( .A(round_reg[701]), .B(init), .Z(\round_in[0][701] ) );
  AND U9979 ( .A(round_reg[702]), .B(init), .Z(\round_in[0][702] ) );
  AND U9980 ( .A(round_reg[703]), .B(init), .Z(\round_in[0][703] ) );
  AND U9981 ( .A(round_reg[704]), .B(init), .Z(\round_in[0][704] ) );
  AND U9982 ( .A(round_reg[705]), .B(init), .Z(\round_in[0][705] ) );
  AND U9983 ( .A(round_reg[706]), .B(init), .Z(\round_in[0][706] ) );
  AND U9984 ( .A(round_reg[707]), .B(init), .Z(\round_in[0][707] ) );
  AND U9985 ( .A(round_reg[708]), .B(init), .Z(\round_in[0][708] ) );
  AND U9986 ( .A(round_reg[709]), .B(init), .Z(\round_in[0][709] ) );
  NAND U9987 ( .A(init), .B(round_reg[70]), .Z(n3852) );
  NANDN U9988 ( .A(init), .B(in[70]), .Z(n3851) );
  NAND U9989 ( .A(n3852), .B(n3851), .Z(\round_in[0][70] ) );
  AND U9990 ( .A(round_reg[710]), .B(init), .Z(\round_in[0][710] ) );
  AND U9991 ( .A(round_reg[711]), .B(init), .Z(\round_in[0][711] ) );
  AND U9992 ( .A(round_reg[712]), .B(init), .Z(\round_in[0][712] ) );
  AND U9993 ( .A(round_reg[713]), .B(init), .Z(\round_in[0][713] ) );
  AND U9994 ( .A(round_reg[714]), .B(init), .Z(\round_in[0][714] ) );
  AND U9995 ( .A(round_reg[715]), .B(init), .Z(\round_in[0][715] ) );
  AND U9996 ( .A(round_reg[716]), .B(init), .Z(\round_in[0][716] ) );
  AND U9997 ( .A(round_reg[717]), .B(init), .Z(\round_in[0][717] ) );
  AND U9998 ( .A(round_reg[718]), .B(init), .Z(\round_in[0][718] ) );
  AND U9999 ( .A(round_reg[719]), .B(init), .Z(\round_in[0][719] ) );
  NAND U10000 ( .A(init), .B(round_reg[71]), .Z(n3854) );
  NANDN U10001 ( .A(init), .B(in[71]), .Z(n3853) );
  NAND U10002 ( .A(n3854), .B(n3853), .Z(\round_in[0][71] ) );
  AND U10003 ( .A(round_reg[720]), .B(init), .Z(\round_in[0][720] ) );
  AND U10004 ( .A(round_reg[721]), .B(init), .Z(\round_in[0][721] ) );
  AND U10005 ( .A(round_reg[722]), .B(init), .Z(\round_in[0][722] ) );
  AND U10006 ( .A(round_reg[723]), .B(init), .Z(\round_in[0][723] ) );
  AND U10007 ( .A(round_reg[724]), .B(init), .Z(\round_in[0][724] ) );
  AND U10008 ( .A(round_reg[725]), .B(init), .Z(\round_in[0][725] ) );
  AND U10009 ( .A(round_reg[726]), .B(init), .Z(\round_in[0][726] ) );
  AND U10010 ( .A(round_reg[727]), .B(init), .Z(\round_in[0][727] ) );
  AND U10011 ( .A(round_reg[728]), .B(init), .Z(\round_in[0][728] ) );
  AND U10012 ( .A(round_reg[729]), .B(init), .Z(\round_in[0][729] ) );
  NAND U10013 ( .A(init), .B(round_reg[72]), .Z(n3856) );
  NANDN U10014 ( .A(init), .B(in[72]), .Z(n3855) );
  NAND U10015 ( .A(n3856), .B(n3855), .Z(\round_in[0][72] ) );
  AND U10016 ( .A(round_reg[730]), .B(init), .Z(\round_in[0][730] ) );
  AND U10017 ( .A(round_reg[731]), .B(init), .Z(\round_in[0][731] ) );
  AND U10018 ( .A(round_reg[732]), .B(init), .Z(\round_in[0][732] ) );
  AND U10019 ( .A(round_reg[733]), .B(init), .Z(\round_in[0][733] ) );
  AND U10020 ( .A(round_reg[734]), .B(init), .Z(\round_in[0][734] ) );
  AND U10021 ( .A(round_reg[735]), .B(init), .Z(\round_in[0][735] ) );
  AND U10022 ( .A(round_reg[736]), .B(init), .Z(\round_in[0][736] ) );
  AND U10023 ( .A(round_reg[737]), .B(init), .Z(\round_in[0][737] ) );
  AND U10024 ( .A(round_reg[738]), .B(init), .Z(\round_in[0][738] ) );
  AND U10025 ( .A(round_reg[739]), .B(init), .Z(\round_in[0][739] ) );
  NAND U10026 ( .A(init), .B(round_reg[73]), .Z(n3858) );
  NANDN U10027 ( .A(init), .B(in[73]), .Z(n3857) );
  NAND U10028 ( .A(n3858), .B(n3857), .Z(\round_in[0][73] ) );
  AND U10029 ( .A(round_reg[740]), .B(init), .Z(\round_in[0][740] ) );
  AND U10030 ( .A(round_reg[741]), .B(init), .Z(\round_in[0][741] ) );
  AND U10031 ( .A(round_reg[742]), .B(init), .Z(\round_in[0][742] ) );
  AND U10032 ( .A(round_reg[743]), .B(init), .Z(\round_in[0][743] ) );
  AND U10033 ( .A(round_reg[744]), .B(init), .Z(\round_in[0][744] ) );
  AND U10034 ( .A(round_reg[745]), .B(init), .Z(\round_in[0][745] ) );
  AND U10035 ( .A(round_reg[746]), .B(init), .Z(\round_in[0][746] ) );
  AND U10036 ( .A(round_reg[747]), .B(init), .Z(\round_in[0][747] ) );
  AND U10037 ( .A(round_reg[748]), .B(init), .Z(\round_in[0][748] ) );
  AND U10038 ( .A(round_reg[749]), .B(init), .Z(\round_in[0][749] ) );
  NAND U10039 ( .A(init), .B(round_reg[74]), .Z(n3860) );
  NANDN U10040 ( .A(init), .B(in[74]), .Z(n3859) );
  NAND U10041 ( .A(n3860), .B(n3859), .Z(\round_in[0][74] ) );
  AND U10042 ( .A(round_reg[750]), .B(init), .Z(\round_in[0][750] ) );
  AND U10043 ( .A(round_reg[751]), .B(init), .Z(\round_in[0][751] ) );
  AND U10044 ( .A(round_reg[752]), .B(init), .Z(\round_in[0][752] ) );
  AND U10045 ( .A(round_reg[753]), .B(init), .Z(\round_in[0][753] ) );
  AND U10046 ( .A(round_reg[754]), .B(init), .Z(\round_in[0][754] ) );
  AND U10047 ( .A(round_reg[755]), .B(init), .Z(\round_in[0][755] ) );
  AND U10048 ( .A(round_reg[756]), .B(init), .Z(\round_in[0][756] ) );
  AND U10049 ( .A(round_reg[757]), .B(init), .Z(\round_in[0][757] ) );
  AND U10050 ( .A(round_reg[758]), .B(init), .Z(\round_in[0][758] ) );
  AND U10051 ( .A(round_reg[759]), .B(init), .Z(\round_in[0][759] ) );
  NAND U10052 ( .A(init), .B(round_reg[75]), .Z(n3862) );
  NANDN U10053 ( .A(init), .B(in[75]), .Z(n3861) );
  NAND U10054 ( .A(n3862), .B(n3861), .Z(\round_in[0][75] ) );
  AND U10055 ( .A(round_reg[760]), .B(init), .Z(\round_in[0][760] ) );
  AND U10056 ( .A(round_reg[761]), .B(init), .Z(\round_in[0][761] ) );
  AND U10057 ( .A(round_reg[762]), .B(init), .Z(\round_in[0][762] ) );
  AND U10058 ( .A(round_reg[763]), .B(init), .Z(\round_in[0][763] ) );
  AND U10059 ( .A(round_reg[764]), .B(init), .Z(\round_in[0][764] ) );
  AND U10060 ( .A(round_reg[765]), .B(init), .Z(\round_in[0][765] ) );
  AND U10061 ( .A(round_reg[766]), .B(init), .Z(\round_in[0][766] ) );
  AND U10062 ( .A(round_reg[767]), .B(init), .Z(\round_in[0][767] ) );
  AND U10063 ( .A(round_reg[768]), .B(init), .Z(\round_in[0][768] ) );
  AND U10064 ( .A(round_reg[769]), .B(init), .Z(\round_in[0][769] ) );
  NAND U10065 ( .A(init), .B(round_reg[76]), .Z(n3864) );
  NANDN U10066 ( .A(init), .B(in[76]), .Z(n3863) );
  NAND U10067 ( .A(n3864), .B(n3863), .Z(\round_in[0][76] ) );
  AND U10068 ( .A(round_reg[770]), .B(init), .Z(\round_in[0][770] ) );
  AND U10069 ( .A(round_reg[771]), .B(init), .Z(\round_in[0][771] ) );
  AND U10070 ( .A(round_reg[772]), .B(init), .Z(\round_in[0][772] ) );
  AND U10071 ( .A(round_reg[773]), .B(init), .Z(\round_in[0][773] ) );
  AND U10072 ( .A(round_reg[774]), .B(init), .Z(\round_in[0][774] ) );
  AND U10073 ( .A(round_reg[775]), .B(init), .Z(\round_in[0][775] ) );
  AND U10074 ( .A(round_reg[776]), .B(init), .Z(\round_in[0][776] ) );
  AND U10075 ( .A(round_reg[777]), .B(init), .Z(\round_in[0][777] ) );
  AND U10076 ( .A(round_reg[778]), .B(init), .Z(\round_in[0][778] ) );
  AND U10077 ( .A(round_reg[779]), .B(init), .Z(\round_in[0][779] ) );
  NAND U10078 ( .A(init), .B(round_reg[77]), .Z(n3866) );
  NANDN U10079 ( .A(init), .B(in[77]), .Z(n3865) );
  NAND U10080 ( .A(n3866), .B(n3865), .Z(\round_in[0][77] ) );
  AND U10081 ( .A(round_reg[780]), .B(init), .Z(\round_in[0][780] ) );
  AND U10082 ( .A(round_reg[781]), .B(init), .Z(\round_in[0][781] ) );
  AND U10083 ( .A(round_reg[782]), .B(init), .Z(\round_in[0][782] ) );
  AND U10084 ( .A(round_reg[783]), .B(init), .Z(\round_in[0][783] ) );
  AND U10085 ( .A(round_reg[784]), .B(init), .Z(\round_in[0][784] ) );
  AND U10086 ( .A(round_reg[785]), .B(init), .Z(\round_in[0][785] ) );
  AND U10087 ( .A(round_reg[786]), .B(init), .Z(\round_in[0][786] ) );
  AND U10088 ( .A(round_reg[787]), .B(init), .Z(\round_in[0][787] ) );
  AND U10089 ( .A(round_reg[788]), .B(init), .Z(\round_in[0][788] ) );
  AND U10090 ( .A(round_reg[789]), .B(init), .Z(\round_in[0][789] ) );
  NAND U10091 ( .A(init), .B(round_reg[78]), .Z(n3868) );
  NANDN U10092 ( .A(init), .B(in[78]), .Z(n3867) );
  NAND U10093 ( .A(n3868), .B(n3867), .Z(\round_in[0][78] ) );
  AND U10094 ( .A(round_reg[790]), .B(init), .Z(\round_in[0][790] ) );
  AND U10095 ( .A(round_reg[791]), .B(init), .Z(\round_in[0][791] ) );
  AND U10096 ( .A(round_reg[792]), .B(init), .Z(\round_in[0][792] ) );
  AND U10097 ( .A(round_reg[793]), .B(init), .Z(\round_in[0][793] ) );
  AND U10098 ( .A(round_reg[794]), .B(init), .Z(\round_in[0][794] ) );
  AND U10099 ( .A(round_reg[795]), .B(init), .Z(\round_in[0][795] ) );
  AND U10100 ( .A(round_reg[796]), .B(init), .Z(\round_in[0][796] ) );
  AND U10101 ( .A(round_reg[797]), .B(init), .Z(\round_in[0][797] ) );
  AND U10102 ( .A(round_reg[798]), .B(init), .Z(\round_in[0][798] ) );
  AND U10103 ( .A(round_reg[799]), .B(init), .Z(\round_in[0][799] ) );
  NAND U10104 ( .A(init), .B(round_reg[79]), .Z(n3870) );
  NANDN U10105 ( .A(init), .B(in[79]), .Z(n3869) );
  NAND U10106 ( .A(n3870), .B(n3869), .Z(\round_in[0][79] ) );
  NAND U10107 ( .A(init), .B(round_reg[7]), .Z(n3872) );
  NANDN U10108 ( .A(init), .B(in[7]), .Z(n3871) );
  NAND U10109 ( .A(n3872), .B(n3871), .Z(\round_in[0][7] ) );
  AND U10110 ( .A(round_reg[800]), .B(init), .Z(\round_in[0][800] ) );
  AND U10111 ( .A(round_reg[801]), .B(init), .Z(\round_in[0][801] ) );
  AND U10112 ( .A(round_reg[802]), .B(init), .Z(\round_in[0][802] ) );
  AND U10113 ( .A(round_reg[803]), .B(init), .Z(\round_in[0][803] ) );
  AND U10114 ( .A(round_reg[804]), .B(init), .Z(\round_in[0][804] ) );
  AND U10115 ( .A(round_reg[805]), .B(init), .Z(\round_in[0][805] ) );
  AND U10116 ( .A(round_reg[806]), .B(init), .Z(\round_in[0][806] ) );
  AND U10117 ( .A(round_reg[807]), .B(init), .Z(\round_in[0][807] ) );
  AND U10118 ( .A(round_reg[808]), .B(init), .Z(\round_in[0][808] ) );
  AND U10119 ( .A(round_reg[809]), .B(init), .Z(\round_in[0][809] ) );
  NAND U10120 ( .A(init), .B(round_reg[80]), .Z(n3874) );
  NANDN U10121 ( .A(init), .B(in[80]), .Z(n3873) );
  NAND U10122 ( .A(n3874), .B(n3873), .Z(\round_in[0][80] ) );
  AND U10123 ( .A(round_reg[810]), .B(init), .Z(\round_in[0][810] ) );
  AND U10124 ( .A(round_reg[811]), .B(init), .Z(\round_in[0][811] ) );
  AND U10125 ( .A(round_reg[812]), .B(init), .Z(\round_in[0][812] ) );
  AND U10126 ( .A(round_reg[813]), .B(init), .Z(\round_in[0][813] ) );
  AND U10127 ( .A(round_reg[814]), .B(init), .Z(\round_in[0][814] ) );
  AND U10128 ( .A(round_reg[815]), .B(init), .Z(\round_in[0][815] ) );
  AND U10129 ( .A(round_reg[816]), .B(init), .Z(\round_in[0][816] ) );
  AND U10130 ( .A(round_reg[817]), .B(init), .Z(\round_in[0][817] ) );
  AND U10131 ( .A(round_reg[818]), .B(init), .Z(\round_in[0][818] ) );
  AND U10132 ( .A(round_reg[819]), .B(init), .Z(\round_in[0][819] ) );
  NAND U10133 ( .A(init), .B(round_reg[81]), .Z(n3876) );
  NANDN U10134 ( .A(init), .B(in[81]), .Z(n3875) );
  NAND U10135 ( .A(n3876), .B(n3875), .Z(\round_in[0][81] ) );
  AND U10136 ( .A(round_reg[820]), .B(init), .Z(\round_in[0][820] ) );
  AND U10137 ( .A(round_reg[821]), .B(init), .Z(\round_in[0][821] ) );
  AND U10138 ( .A(round_reg[822]), .B(init), .Z(\round_in[0][822] ) );
  AND U10139 ( .A(round_reg[823]), .B(init), .Z(\round_in[0][823] ) );
  AND U10140 ( .A(round_reg[824]), .B(init), .Z(\round_in[0][824] ) );
  AND U10141 ( .A(round_reg[825]), .B(init), .Z(\round_in[0][825] ) );
  AND U10142 ( .A(round_reg[826]), .B(init), .Z(\round_in[0][826] ) );
  AND U10143 ( .A(round_reg[827]), .B(init), .Z(\round_in[0][827] ) );
  AND U10144 ( .A(round_reg[828]), .B(init), .Z(\round_in[0][828] ) );
  AND U10145 ( .A(round_reg[829]), .B(init), .Z(\round_in[0][829] ) );
  NAND U10146 ( .A(init), .B(round_reg[82]), .Z(n3878) );
  NANDN U10147 ( .A(init), .B(in[82]), .Z(n3877) );
  NAND U10148 ( .A(n3878), .B(n3877), .Z(\round_in[0][82] ) );
  AND U10149 ( .A(round_reg[830]), .B(init), .Z(\round_in[0][830] ) );
  AND U10150 ( .A(round_reg[831]), .B(init), .Z(\round_in[0][831] ) );
  AND U10151 ( .A(round_reg[832]), .B(init), .Z(\round_in[0][832] ) );
  AND U10152 ( .A(round_reg[833]), .B(init), .Z(\round_in[0][833] ) );
  AND U10153 ( .A(round_reg[834]), .B(init), .Z(\round_in[0][834] ) );
  AND U10154 ( .A(round_reg[835]), .B(init), .Z(\round_in[0][835] ) );
  AND U10155 ( .A(round_reg[836]), .B(init), .Z(\round_in[0][836] ) );
  AND U10156 ( .A(round_reg[837]), .B(init), .Z(\round_in[0][837] ) );
  AND U10157 ( .A(round_reg[838]), .B(init), .Z(\round_in[0][838] ) );
  AND U10158 ( .A(round_reg[839]), .B(init), .Z(\round_in[0][839] ) );
  NAND U10159 ( .A(init), .B(round_reg[83]), .Z(n3880) );
  NANDN U10160 ( .A(init), .B(in[83]), .Z(n3879) );
  NAND U10161 ( .A(n3880), .B(n3879), .Z(\round_in[0][83] ) );
  AND U10162 ( .A(round_reg[840]), .B(init), .Z(\round_in[0][840] ) );
  AND U10163 ( .A(round_reg[841]), .B(init), .Z(\round_in[0][841] ) );
  AND U10164 ( .A(round_reg[842]), .B(init), .Z(\round_in[0][842] ) );
  AND U10165 ( .A(round_reg[843]), .B(init), .Z(\round_in[0][843] ) );
  AND U10166 ( .A(round_reg[844]), .B(init), .Z(\round_in[0][844] ) );
  AND U10167 ( .A(round_reg[845]), .B(init), .Z(\round_in[0][845] ) );
  AND U10168 ( .A(round_reg[846]), .B(init), .Z(\round_in[0][846] ) );
  AND U10169 ( .A(round_reg[847]), .B(init), .Z(\round_in[0][847] ) );
  AND U10170 ( .A(round_reg[848]), .B(init), .Z(\round_in[0][848] ) );
  AND U10171 ( .A(round_reg[849]), .B(init), .Z(\round_in[0][849] ) );
  NAND U10172 ( .A(init), .B(round_reg[84]), .Z(n3882) );
  NANDN U10173 ( .A(init), .B(in[84]), .Z(n3881) );
  NAND U10174 ( .A(n3882), .B(n3881), .Z(\round_in[0][84] ) );
  AND U10175 ( .A(round_reg[850]), .B(init), .Z(\round_in[0][850] ) );
  AND U10176 ( .A(round_reg[851]), .B(init), .Z(\round_in[0][851] ) );
  AND U10177 ( .A(round_reg[852]), .B(init), .Z(\round_in[0][852] ) );
  AND U10178 ( .A(round_reg[853]), .B(init), .Z(\round_in[0][853] ) );
  AND U10179 ( .A(round_reg[854]), .B(init), .Z(\round_in[0][854] ) );
  AND U10180 ( .A(round_reg[855]), .B(init), .Z(\round_in[0][855] ) );
  AND U10181 ( .A(round_reg[856]), .B(init), .Z(\round_in[0][856] ) );
  AND U10182 ( .A(round_reg[857]), .B(init), .Z(\round_in[0][857] ) );
  AND U10183 ( .A(round_reg[858]), .B(init), .Z(\round_in[0][858] ) );
  AND U10184 ( .A(round_reg[859]), .B(init), .Z(\round_in[0][859] ) );
  NAND U10185 ( .A(init), .B(round_reg[85]), .Z(n3884) );
  NANDN U10186 ( .A(init), .B(in[85]), .Z(n3883) );
  NAND U10187 ( .A(n3884), .B(n3883), .Z(\round_in[0][85] ) );
  AND U10188 ( .A(round_reg[860]), .B(init), .Z(\round_in[0][860] ) );
  AND U10189 ( .A(round_reg[861]), .B(init), .Z(\round_in[0][861] ) );
  AND U10190 ( .A(round_reg[862]), .B(init), .Z(\round_in[0][862] ) );
  AND U10191 ( .A(round_reg[863]), .B(init), .Z(\round_in[0][863] ) );
  AND U10192 ( .A(round_reg[864]), .B(init), .Z(\round_in[0][864] ) );
  AND U10193 ( .A(round_reg[865]), .B(init), .Z(\round_in[0][865] ) );
  AND U10194 ( .A(round_reg[866]), .B(init), .Z(\round_in[0][866] ) );
  AND U10195 ( .A(round_reg[867]), .B(init), .Z(\round_in[0][867] ) );
  AND U10196 ( .A(round_reg[868]), .B(init), .Z(\round_in[0][868] ) );
  AND U10197 ( .A(round_reg[869]), .B(init), .Z(\round_in[0][869] ) );
  NAND U10198 ( .A(init), .B(round_reg[86]), .Z(n3886) );
  NANDN U10199 ( .A(init), .B(in[86]), .Z(n3885) );
  NAND U10200 ( .A(n3886), .B(n3885), .Z(\round_in[0][86] ) );
  AND U10201 ( .A(round_reg[870]), .B(init), .Z(\round_in[0][870] ) );
  AND U10202 ( .A(round_reg[871]), .B(init), .Z(\round_in[0][871] ) );
  AND U10203 ( .A(round_reg[872]), .B(init), .Z(\round_in[0][872] ) );
  AND U10204 ( .A(round_reg[873]), .B(init), .Z(\round_in[0][873] ) );
  AND U10205 ( .A(round_reg[874]), .B(init), .Z(\round_in[0][874] ) );
  AND U10206 ( .A(round_reg[875]), .B(init), .Z(\round_in[0][875] ) );
  AND U10207 ( .A(round_reg[876]), .B(init), .Z(\round_in[0][876] ) );
  AND U10208 ( .A(round_reg[877]), .B(init), .Z(\round_in[0][877] ) );
  AND U10209 ( .A(round_reg[878]), .B(init), .Z(\round_in[0][878] ) );
  AND U10210 ( .A(round_reg[879]), .B(init), .Z(\round_in[0][879] ) );
  NAND U10211 ( .A(init), .B(round_reg[87]), .Z(n3888) );
  NANDN U10212 ( .A(init), .B(in[87]), .Z(n3887) );
  NAND U10213 ( .A(n3888), .B(n3887), .Z(\round_in[0][87] ) );
  AND U10214 ( .A(round_reg[880]), .B(init), .Z(\round_in[0][880] ) );
  AND U10215 ( .A(round_reg[881]), .B(init), .Z(\round_in[0][881] ) );
  AND U10216 ( .A(round_reg[882]), .B(init), .Z(\round_in[0][882] ) );
  AND U10217 ( .A(round_reg[883]), .B(init), .Z(\round_in[0][883] ) );
  AND U10218 ( .A(round_reg[884]), .B(init), .Z(\round_in[0][884] ) );
  AND U10219 ( .A(round_reg[885]), .B(init), .Z(\round_in[0][885] ) );
  AND U10220 ( .A(round_reg[886]), .B(init), .Z(\round_in[0][886] ) );
  AND U10221 ( .A(round_reg[887]), .B(init), .Z(\round_in[0][887] ) );
  AND U10222 ( .A(round_reg[888]), .B(init), .Z(\round_in[0][888] ) );
  AND U10223 ( .A(round_reg[889]), .B(init), .Z(\round_in[0][889] ) );
  NAND U10224 ( .A(init), .B(round_reg[88]), .Z(n3890) );
  NANDN U10225 ( .A(init), .B(in[88]), .Z(n3889) );
  NAND U10226 ( .A(n3890), .B(n3889), .Z(\round_in[0][88] ) );
  AND U10227 ( .A(round_reg[890]), .B(init), .Z(\round_in[0][890] ) );
  AND U10228 ( .A(round_reg[891]), .B(init), .Z(\round_in[0][891] ) );
  AND U10229 ( .A(round_reg[892]), .B(init), .Z(\round_in[0][892] ) );
  AND U10230 ( .A(round_reg[893]), .B(init), .Z(\round_in[0][893] ) );
  AND U10231 ( .A(round_reg[894]), .B(init), .Z(\round_in[0][894] ) );
  AND U10232 ( .A(round_reg[895]), .B(init), .Z(\round_in[0][895] ) );
  AND U10233 ( .A(round_reg[896]), .B(init), .Z(\round_in[0][896] ) );
  AND U10234 ( .A(round_reg[897]), .B(init), .Z(\round_in[0][897] ) );
  AND U10235 ( .A(round_reg[898]), .B(init), .Z(\round_in[0][898] ) );
  AND U10236 ( .A(round_reg[899]), .B(init), .Z(\round_in[0][899] ) );
  NAND U10237 ( .A(init), .B(round_reg[89]), .Z(n3892) );
  NANDN U10238 ( .A(init), .B(in[89]), .Z(n3891) );
  NAND U10239 ( .A(n3892), .B(n3891), .Z(\round_in[0][89] ) );
  NAND U10240 ( .A(init), .B(round_reg[8]), .Z(n3894) );
  NANDN U10241 ( .A(init), .B(in[8]), .Z(n3893) );
  NAND U10242 ( .A(n3894), .B(n3893), .Z(\round_in[0][8] ) );
  AND U10243 ( .A(round_reg[900]), .B(init), .Z(\round_in[0][900] ) );
  AND U10244 ( .A(round_reg[901]), .B(init), .Z(\round_in[0][901] ) );
  AND U10245 ( .A(round_reg[902]), .B(init), .Z(\round_in[0][902] ) );
  AND U10246 ( .A(round_reg[903]), .B(init), .Z(\round_in[0][903] ) );
  AND U10247 ( .A(round_reg[904]), .B(init), .Z(\round_in[0][904] ) );
  AND U10248 ( .A(round_reg[905]), .B(init), .Z(\round_in[0][905] ) );
  AND U10249 ( .A(round_reg[906]), .B(init), .Z(\round_in[0][906] ) );
  AND U10250 ( .A(round_reg[907]), .B(init), .Z(\round_in[0][907] ) );
  AND U10251 ( .A(round_reg[908]), .B(init), .Z(\round_in[0][908] ) );
  AND U10252 ( .A(round_reg[909]), .B(init), .Z(\round_in[0][909] ) );
  NAND U10253 ( .A(init), .B(round_reg[90]), .Z(n3896) );
  NANDN U10254 ( .A(init), .B(in[90]), .Z(n3895) );
  NAND U10255 ( .A(n3896), .B(n3895), .Z(\round_in[0][90] ) );
  AND U10256 ( .A(round_reg[910]), .B(init), .Z(\round_in[0][910] ) );
  AND U10257 ( .A(round_reg[911]), .B(init), .Z(\round_in[0][911] ) );
  AND U10258 ( .A(round_reg[912]), .B(init), .Z(\round_in[0][912] ) );
  AND U10259 ( .A(round_reg[913]), .B(init), .Z(\round_in[0][913] ) );
  AND U10260 ( .A(round_reg[914]), .B(init), .Z(\round_in[0][914] ) );
  AND U10261 ( .A(round_reg[915]), .B(init), .Z(\round_in[0][915] ) );
  AND U10262 ( .A(round_reg[916]), .B(init), .Z(\round_in[0][916] ) );
  AND U10263 ( .A(round_reg[917]), .B(init), .Z(\round_in[0][917] ) );
  AND U10264 ( .A(round_reg[918]), .B(init), .Z(\round_in[0][918] ) );
  AND U10265 ( .A(round_reg[919]), .B(init), .Z(\round_in[0][919] ) );
  NAND U10266 ( .A(init), .B(round_reg[91]), .Z(n3898) );
  NANDN U10267 ( .A(init), .B(in[91]), .Z(n3897) );
  NAND U10268 ( .A(n3898), .B(n3897), .Z(\round_in[0][91] ) );
  AND U10269 ( .A(round_reg[920]), .B(init), .Z(\round_in[0][920] ) );
  AND U10270 ( .A(round_reg[921]), .B(init), .Z(\round_in[0][921] ) );
  AND U10271 ( .A(round_reg[922]), .B(init), .Z(\round_in[0][922] ) );
  AND U10272 ( .A(round_reg[923]), .B(init), .Z(\round_in[0][923] ) );
  AND U10273 ( .A(round_reg[924]), .B(init), .Z(\round_in[0][924] ) );
  AND U10274 ( .A(round_reg[925]), .B(init), .Z(\round_in[0][925] ) );
  AND U10275 ( .A(round_reg[926]), .B(init), .Z(\round_in[0][926] ) );
  AND U10276 ( .A(round_reg[927]), .B(init), .Z(\round_in[0][927] ) );
  AND U10277 ( .A(round_reg[928]), .B(init), .Z(\round_in[0][928] ) );
  AND U10278 ( .A(round_reg[929]), .B(init), .Z(\round_in[0][929] ) );
  NAND U10279 ( .A(init), .B(round_reg[92]), .Z(n3900) );
  NANDN U10280 ( .A(init), .B(in[92]), .Z(n3899) );
  NAND U10281 ( .A(n3900), .B(n3899), .Z(\round_in[0][92] ) );
  AND U10282 ( .A(round_reg[930]), .B(init), .Z(\round_in[0][930] ) );
  AND U10283 ( .A(round_reg[931]), .B(init), .Z(\round_in[0][931] ) );
  AND U10284 ( .A(round_reg[932]), .B(init), .Z(\round_in[0][932] ) );
  AND U10285 ( .A(round_reg[933]), .B(init), .Z(\round_in[0][933] ) );
  AND U10286 ( .A(round_reg[934]), .B(init), .Z(\round_in[0][934] ) );
  AND U10287 ( .A(round_reg[935]), .B(init), .Z(\round_in[0][935] ) );
  AND U10288 ( .A(round_reg[936]), .B(init), .Z(\round_in[0][936] ) );
  AND U10289 ( .A(round_reg[937]), .B(init), .Z(\round_in[0][937] ) );
  AND U10290 ( .A(round_reg[938]), .B(init), .Z(\round_in[0][938] ) );
  AND U10291 ( .A(round_reg[939]), .B(init), .Z(\round_in[0][939] ) );
  NAND U10292 ( .A(init), .B(round_reg[93]), .Z(n3902) );
  NANDN U10293 ( .A(init), .B(in[93]), .Z(n3901) );
  NAND U10294 ( .A(n3902), .B(n3901), .Z(\round_in[0][93] ) );
  AND U10295 ( .A(round_reg[940]), .B(init), .Z(\round_in[0][940] ) );
  AND U10296 ( .A(round_reg[941]), .B(init), .Z(\round_in[0][941] ) );
  AND U10297 ( .A(round_reg[942]), .B(init), .Z(\round_in[0][942] ) );
  AND U10298 ( .A(round_reg[943]), .B(init), .Z(\round_in[0][943] ) );
  AND U10299 ( .A(round_reg[944]), .B(init), .Z(\round_in[0][944] ) );
  AND U10300 ( .A(round_reg[945]), .B(init), .Z(\round_in[0][945] ) );
  AND U10301 ( .A(round_reg[946]), .B(init), .Z(\round_in[0][946] ) );
  AND U10302 ( .A(round_reg[947]), .B(init), .Z(\round_in[0][947] ) );
  AND U10303 ( .A(round_reg[948]), .B(init), .Z(\round_in[0][948] ) );
  AND U10304 ( .A(round_reg[949]), .B(init), .Z(\round_in[0][949] ) );
  NAND U10305 ( .A(init), .B(round_reg[94]), .Z(n3904) );
  NANDN U10306 ( .A(init), .B(in[94]), .Z(n3903) );
  NAND U10307 ( .A(n3904), .B(n3903), .Z(\round_in[0][94] ) );
  AND U10308 ( .A(round_reg[950]), .B(init), .Z(\round_in[0][950] ) );
  AND U10309 ( .A(round_reg[951]), .B(init), .Z(\round_in[0][951] ) );
  AND U10310 ( .A(round_reg[952]), .B(init), .Z(\round_in[0][952] ) );
  AND U10311 ( .A(round_reg[953]), .B(init), .Z(\round_in[0][953] ) );
  AND U10312 ( .A(round_reg[954]), .B(init), .Z(\round_in[0][954] ) );
  AND U10313 ( .A(round_reg[955]), .B(init), .Z(\round_in[0][955] ) );
  AND U10314 ( .A(round_reg[956]), .B(init), .Z(\round_in[0][956] ) );
  AND U10315 ( .A(round_reg[957]), .B(init), .Z(\round_in[0][957] ) );
  AND U10316 ( .A(round_reg[958]), .B(init), .Z(\round_in[0][958] ) );
  AND U10317 ( .A(round_reg[959]), .B(init), .Z(\round_in[0][959] ) );
  NAND U10318 ( .A(init), .B(round_reg[95]), .Z(n3906) );
  NANDN U10319 ( .A(init), .B(in[95]), .Z(n3905) );
  NAND U10320 ( .A(n3906), .B(n3905), .Z(\round_in[0][95] ) );
  AND U10321 ( .A(round_reg[960]), .B(init), .Z(\round_in[0][960] ) );
  AND U10322 ( .A(round_reg[961]), .B(init), .Z(\round_in[0][961] ) );
  AND U10323 ( .A(round_reg[962]), .B(init), .Z(\round_in[0][962] ) );
  AND U10324 ( .A(round_reg[963]), .B(init), .Z(\round_in[0][963] ) );
  AND U10325 ( .A(round_reg[964]), .B(init), .Z(\round_in[0][964] ) );
  AND U10326 ( .A(round_reg[965]), .B(init), .Z(\round_in[0][965] ) );
  AND U10327 ( .A(round_reg[966]), .B(init), .Z(\round_in[0][966] ) );
  AND U10328 ( .A(round_reg[967]), .B(init), .Z(\round_in[0][967] ) );
  AND U10329 ( .A(round_reg[968]), .B(init), .Z(\round_in[0][968] ) );
  AND U10330 ( .A(round_reg[969]), .B(init), .Z(\round_in[0][969] ) );
  NAND U10331 ( .A(init), .B(round_reg[96]), .Z(n3908) );
  NANDN U10332 ( .A(init), .B(in[96]), .Z(n3907) );
  NAND U10333 ( .A(n3908), .B(n3907), .Z(\round_in[0][96] ) );
  AND U10334 ( .A(round_reg[970]), .B(init), .Z(\round_in[0][970] ) );
  AND U10335 ( .A(round_reg[971]), .B(init), .Z(\round_in[0][971] ) );
  AND U10336 ( .A(round_reg[972]), .B(init), .Z(\round_in[0][972] ) );
  AND U10337 ( .A(round_reg[973]), .B(init), .Z(\round_in[0][973] ) );
  AND U10338 ( .A(round_reg[974]), .B(init), .Z(\round_in[0][974] ) );
  AND U10339 ( .A(round_reg[975]), .B(init), .Z(\round_in[0][975] ) );
  AND U10340 ( .A(round_reg[976]), .B(init), .Z(\round_in[0][976] ) );
  AND U10341 ( .A(round_reg[977]), .B(init), .Z(\round_in[0][977] ) );
  AND U10342 ( .A(round_reg[978]), .B(init), .Z(\round_in[0][978] ) );
  AND U10343 ( .A(round_reg[979]), .B(init), .Z(\round_in[0][979] ) );
  NAND U10344 ( .A(init), .B(round_reg[97]), .Z(n3910) );
  NANDN U10345 ( .A(init), .B(in[97]), .Z(n3909) );
  NAND U10346 ( .A(n3910), .B(n3909), .Z(\round_in[0][97] ) );
  AND U10347 ( .A(round_reg[980]), .B(init), .Z(\round_in[0][980] ) );
  AND U10348 ( .A(round_reg[981]), .B(init), .Z(\round_in[0][981] ) );
  AND U10349 ( .A(round_reg[982]), .B(init), .Z(\round_in[0][982] ) );
  AND U10350 ( .A(round_reg[983]), .B(init), .Z(\round_in[0][983] ) );
  AND U10351 ( .A(round_reg[984]), .B(init), .Z(\round_in[0][984] ) );
  AND U10352 ( .A(round_reg[985]), .B(init), .Z(\round_in[0][985] ) );
  AND U10353 ( .A(round_reg[986]), .B(init), .Z(\round_in[0][986] ) );
  AND U10354 ( .A(round_reg[987]), .B(init), .Z(\round_in[0][987] ) );
  AND U10355 ( .A(round_reg[988]), .B(init), .Z(\round_in[0][988] ) );
  AND U10356 ( .A(round_reg[989]), .B(init), .Z(\round_in[0][989] ) );
  NAND U10357 ( .A(init), .B(round_reg[98]), .Z(n3912) );
  NANDN U10358 ( .A(init), .B(in[98]), .Z(n3911) );
  NAND U10359 ( .A(n3912), .B(n3911), .Z(\round_in[0][98] ) );
  AND U10360 ( .A(round_reg[990]), .B(init), .Z(\round_in[0][990] ) );
  AND U10361 ( .A(round_reg[991]), .B(init), .Z(\round_in[0][991] ) );
  AND U10362 ( .A(round_reg[992]), .B(init), .Z(\round_in[0][992] ) );
  AND U10363 ( .A(round_reg[993]), .B(init), .Z(\round_in[0][993] ) );
  AND U10364 ( .A(round_reg[994]), .B(init), .Z(\round_in[0][994] ) );
  AND U10365 ( .A(round_reg[995]), .B(init), .Z(\round_in[0][995] ) );
  AND U10366 ( .A(round_reg[996]), .B(init), .Z(\round_in[0][996] ) );
  AND U10367 ( .A(round_reg[997]), .B(init), .Z(\round_in[0][997] ) );
  AND U10368 ( .A(round_reg[998]), .B(init), .Z(\round_in[0][998] ) );
  AND U10369 ( .A(round_reg[999]), .B(init), .Z(\round_in[0][999] ) );
  NAND U10370 ( .A(init), .B(round_reg[99]), .Z(n3914) );
  NANDN U10371 ( .A(init), .B(in[99]), .Z(n3913) );
  NAND U10372 ( .A(n3914), .B(n3913), .Z(\round_in[0][99] ) );
  NAND U10373 ( .A(init), .B(round_reg[9]), .Z(n3916) );
  NANDN U10374 ( .A(init), .B(in[9]), .Z(n3915) );
  NAND U10375 ( .A(n3916), .B(n3915), .Z(\round_in[0][9] ) );
endmodule

