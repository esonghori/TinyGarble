
module matrixMult_N_M_1_N5_M8 ( clk, rst, x, y, o );
  input [39:0] x;
  input [199:0] y;
  output [39:0] o;
  input clk, rst;
  wire   N9, N10, N11, N12, N13, N14, N15, N16, N25, N26, N27, N28, N29, N30,
         N31, N32, N41, N42, N43, N44, N45, N46, N47, N48, N57, N58, N59, N60,
         N61, N62, N63, N64, N73, N74, N75, N76, N77, N78, N79, N80, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870;

  DFF \oi_reg[0][7]  ( .D(N16), .CLK(clk), .RST(rst), .Q(o[7]) );
  DFF \oi_reg[0][6]  ( .D(N15), .CLK(clk), .RST(rst), .Q(o[6]) );
  DFF \oi_reg[0][5]  ( .D(N14), .CLK(clk), .RST(rst), .Q(o[5]) );
  DFF \oi_reg[0][4]  ( .D(N13), .CLK(clk), .RST(rst), .Q(o[4]) );
  DFF \oi_reg[0][3]  ( .D(N12), .CLK(clk), .RST(rst), .Q(o[3]) );
  DFF \oi_reg[0][2]  ( .D(N11), .CLK(clk), .RST(rst), .Q(o[2]) );
  DFF \oi_reg[0][1]  ( .D(N10), .CLK(clk), .RST(rst), .Q(o[1]) );
  DFF \oi_reg[0][0]  ( .D(N9), .CLK(clk), .RST(rst), .Q(o[0]) );
  DFF \oi_reg[1][7]  ( .D(N32), .CLK(clk), .RST(rst), .Q(o[15]) );
  DFF \oi_reg[1][6]  ( .D(N31), .CLK(clk), .RST(rst), .Q(o[14]) );
  DFF \oi_reg[1][5]  ( .D(N30), .CLK(clk), .RST(rst), .Q(o[13]) );
  DFF \oi_reg[1][4]  ( .D(N29), .CLK(clk), .RST(rst), .Q(o[12]) );
  DFF \oi_reg[1][3]  ( .D(N28), .CLK(clk), .RST(rst), .Q(o[11]) );
  DFF \oi_reg[1][2]  ( .D(N27), .CLK(clk), .RST(rst), .Q(o[10]) );
  DFF \oi_reg[1][1]  ( .D(N26), .CLK(clk), .RST(rst), .Q(o[9]) );
  DFF \oi_reg[1][0]  ( .D(N25), .CLK(clk), .RST(rst), .Q(o[8]) );
  DFF \oi_reg[2][7]  ( .D(N48), .CLK(clk), .RST(rst), .Q(o[23]) );
  DFF \oi_reg[2][6]  ( .D(N47), .CLK(clk), .RST(rst), .Q(o[22]) );
  DFF \oi_reg[2][5]  ( .D(N46), .CLK(clk), .RST(rst), .Q(o[21]) );
  DFF \oi_reg[2][4]  ( .D(N45), .CLK(clk), .RST(rst), .Q(o[20]) );
  DFF \oi_reg[2][3]  ( .D(N44), .CLK(clk), .RST(rst), .Q(o[19]) );
  DFF \oi_reg[2][2]  ( .D(N43), .CLK(clk), .RST(rst), .Q(o[18]) );
  DFF \oi_reg[2][1]  ( .D(N42), .CLK(clk), .RST(rst), .Q(o[17]) );
  DFF \oi_reg[2][0]  ( .D(N41), .CLK(clk), .RST(rst), .Q(o[16]) );
  DFF \oi_reg[3][7]  ( .D(N64), .CLK(clk), .RST(rst), .Q(o[31]) );
  DFF \oi_reg[3][6]  ( .D(N63), .CLK(clk), .RST(rst), .Q(o[30]) );
  DFF \oi_reg[3][5]  ( .D(N62), .CLK(clk), .RST(rst), .Q(o[29]) );
  DFF \oi_reg[3][4]  ( .D(N61), .CLK(clk), .RST(rst), .Q(o[28]) );
  DFF \oi_reg[3][3]  ( .D(N60), .CLK(clk), .RST(rst), .Q(o[27]) );
  DFF \oi_reg[3][2]  ( .D(N59), .CLK(clk), .RST(rst), .Q(o[26]) );
  DFF \oi_reg[3][1]  ( .D(N58), .CLK(clk), .RST(rst), .Q(o[25]) );
  DFF \oi_reg[3][0]  ( .D(N57), .CLK(clk), .RST(rst), .Q(o[24]) );
  DFF \oi_reg[4][7]  ( .D(N80), .CLK(clk), .RST(rst), .Q(o[39]) );
  DFF \oi_reg[4][6]  ( .D(N79), .CLK(clk), .RST(rst), .Q(o[38]) );
  DFF \oi_reg[4][5]  ( .D(N78), .CLK(clk), .RST(rst), .Q(o[37]) );
  DFF \oi_reg[4][4]  ( .D(N77), .CLK(clk), .RST(rst), .Q(o[36]) );
  DFF \oi_reg[4][3]  ( .D(N76), .CLK(clk), .RST(rst), .Q(o[35]) );
  DFF \oi_reg[4][2]  ( .D(N75), .CLK(clk), .RST(rst), .Q(o[34]) );
  DFF \oi_reg[4][1]  ( .D(N74), .CLK(clk), .RST(rst), .Q(o[33]) );
  DFF \oi_reg[4][0]  ( .D(N73), .CLK(clk), .RST(rst), .Q(o[32]) );
  NAND U3 ( .A(n793), .B(n794), .Z(n1) );
  XOR U4 ( .A(n793), .B(n794), .Z(n2) );
  NANDN U5 ( .A(n792), .B(n2), .Z(n3) );
  NAND U6 ( .A(n1), .B(n3), .Z(n806) );
  NAND U7 ( .A(n665), .B(n666), .Z(n4) );
  XOR U8 ( .A(n665), .B(n666), .Z(n5) );
  NANDN U9 ( .A(n664), .B(n5), .Z(n6) );
  NAND U10 ( .A(n4), .B(n6), .Z(n678) );
  NAND U11 ( .A(n537), .B(n538), .Z(n7) );
  XOR U12 ( .A(n537), .B(n538), .Z(n8) );
  NANDN U13 ( .A(n536), .B(n8), .Z(n9) );
  NAND U14 ( .A(n7), .B(n9), .Z(n550) );
  NAND U15 ( .A(n409), .B(n410), .Z(n10) );
  XOR U16 ( .A(n409), .B(n410), .Z(n11) );
  NANDN U17 ( .A(n408), .B(n11), .Z(n12) );
  NAND U18 ( .A(n10), .B(n12), .Z(n422) );
  NAND U19 ( .A(n281), .B(n282), .Z(n13) );
  XOR U20 ( .A(n281), .B(n282), .Z(n14) );
  NANDN U21 ( .A(n280), .B(n14), .Z(n15) );
  NAND U22 ( .A(n13), .B(n15), .Z(n294) );
  XOR U23 ( .A(n855), .B(n854), .Z(n16) );
  XNOR U24 ( .A(n857), .B(n16), .Z(n827) );
  XOR U25 ( .A(n727), .B(n726), .Z(n17) );
  XNOR U26 ( .A(n729), .B(n17), .Z(n699) );
  XOR U27 ( .A(n599), .B(n598), .Z(n18) );
  XNOR U28 ( .A(n601), .B(n18), .Z(n571) );
  XOR U29 ( .A(n471), .B(n470), .Z(n19) );
  XNOR U30 ( .A(n473), .B(n19), .Z(n443) );
  XOR U31 ( .A(n343), .B(n342), .Z(n20) );
  XNOR U32 ( .A(n345), .B(n20), .Z(n315) );
  NAND U33 ( .A(n790), .B(n791), .Z(n21) );
  XOR U34 ( .A(n790), .B(n791), .Z(n22) );
  NANDN U35 ( .A(n789), .B(n22), .Z(n23) );
  NAND U36 ( .A(n21), .B(n23), .Z(n805) );
  NAND U37 ( .A(n662), .B(n663), .Z(n24) );
  XOR U38 ( .A(n662), .B(n663), .Z(n25) );
  NANDN U39 ( .A(n661), .B(n25), .Z(n26) );
  NAND U40 ( .A(n24), .B(n26), .Z(n677) );
  NAND U41 ( .A(n534), .B(n535), .Z(n27) );
  XOR U42 ( .A(n534), .B(n535), .Z(n28) );
  NANDN U43 ( .A(n533), .B(n28), .Z(n29) );
  NAND U44 ( .A(n27), .B(n29), .Z(n549) );
  NAND U45 ( .A(n406), .B(n407), .Z(n30) );
  XOR U46 ( .A(n406), .B(n407), .Z(n31) );
  NANDN U47 ( .A(n405), .B(n31), .Z(n32) );
  NAND U48 ( .A(n30), .B(n32), .Z(n421) );
  NAND U49 ( .A(n278), .B(n279), .Z(n33) );
  XOR U50 ( .A(n278), .B(n279), .Z(n34) );
  NANDN U51 ( .A(n277), .B(n34), .Z(n35) );
  NAND U52 ( .A(n33), .B(n35), .Z(n293) );
  NAND U53 ( .A(n815), .B(n816), .Z(n36) );
  XOR U54 ( .A(n815), .B(n816), .Z(n37) );
  NANDN U55 ( .A(n814), .B(n37), .Z(n38) );
  NAND U56 ( .A(n36), .B(n38), .Z(n861) );
  NAND U57 ( .A(n687), .B(n688), .Z(n39) );
  XOR U58 ( .A(n687), .B(n688), .Z(n40) );
  NANDN U59 ( .A(n686), .B(n40), .Z(n41) );
  NAND U60 ( .A(n39), .B(n41), .Z(n733) );
  NAND U61 ( .A(n559), .B(n560), .Z(n42) );
  XOR U62 ( .A(n559), .B(n560), .Z(n43) );
  NANDN U63 ( .A(n558), .B(n43), .Z(n44) );
  NAND U64 ( .A(n42), .B(n44), .Z(n605) );
  NAND U65 ( .A(n431), .B(n432), .Z(n45) );
  XOR U66 ( .A(n431), .B(n432), .Z(n46) );
  NANDN U67 ( .A(n430), .B(n46), .Z(n47) );
  NAND U68 ( .A(n45), .B(n47), .Z(n477) );
  NAND U69 ( .A(n303), .B(n304), .Z(n48) );
  XOR U70 ( .A(n303), .B(n304), .Z(n49) );
  NANDN U71 ( .A(n302), .B(n49), .Z(n50) );
  NAND U72 ( .A(n48), .B(n50), .Z(n349) );
  NAND U73 ( .A(n821), .B(n819), .Z(n51) );
  XOR U74 ( .A(n821), .B(n819), .Z(n52) );
  NANDN U75 ( .A(n820), .B(n52), .Z(n53) );
  NAND U76 ( .A(n51), .B(n53), .Z(n824) );
  NAND U77 ( .A(n693), .B(n691), .Z(n54) );
  XOR U78 ( .A(n693), .B(n691), .Z(n55) );
  NANDN U79 ( .A(n692), .B(n55), .Z(n56) );
  NAND U80 ( .A(n54), .B(n56), .Z(n696) );
  NAND U81 ( .A(n565), .B(n563), .Z(n57) );
  XOR U82 ( .A(n565), .B(n563), .Z(n58) );
  NANDN U83 ( .A(n564), .B(n58), .Z(n59) );
  NAND U84 ( .A(n57), .B(n59), .Z(n568) );
  NAND U85 ( .A(n437), .B(n435), .Z(n60) );
  XOR U86 ( .A(n437), .B(n435), .Z(n61) );
  NANDN U87 ( .A(n436), .B(n61), .Z(n62) );
  NAND U88 ( .A(n60), .B(n62), .Z(n440) );
  NAND U89 ( .A(n309), .B(n307), .Z(n63) );
  XOR U90 ( .A(n309), .B(n307), .Z(n64) );
  NANDN U91 ( .A(n308), .B(n64), .Z(n65) );
  NAND U92 ( .A(n63), .B(n65), .Z(n312) );
  NAND U93 ( .A(n781), .B(n782), .Z(n66) );
  XOR U94 ( .A(n781), .B(n782), .Z(n67) );
  NANDN U95 ( .A(n780), .B(n67), .Z(n68) );
  NAND U96 ( .A(n66), .B(n68), .Z(n800) );
  NAND U97 ( .A(n812), .B(n813), .Z(n69) );
  XOR U98 ( .A(n812), .B(n813), .Z(n70) );
  NANDN U99 ( .A(n811), .B(n70), .Z(n71) );
  NAND U100 ( .A(n69), .B(n71), .Z(n862) );
  NAND U101 ( .A(n653), .B(n654), .Z(n72) );
  XOR U102 ( .A(n653), .B(n654), .Z(n73) );
  NANDN U103 ( .A(n652), .B(n73), .Z(n74) );
  NAND U104 ( .A(n72), .B(n74), .Z(n672) );
  NAND U105 ( .A(n684), .B(n685), .Z(n75) );
  XOR U106 ( .A(n684), .B(n685), .Z(n76) );
  NANDN U107 ( .A(n683), .B(n76), .Z(n77) );
  NAND U108 ( .A(n75), .B(n77), .Z(n734) );
  NAND U109 ( .A(n525), .B(n526), .Z(n78) );
  XOR U110 ( .A(n525), .B(n526), .Z(n79) );
  NANDN U111 ( .A(n524), .B(n79), .Z(n80) );
  NAND U112 ( .A(n78), .B(n80), .Z(n544) );
  NAND U113 ( .A(n556), .B(n557), .Z(n81) );
  XOR U114 ( .A(n556), .B(n557), .Z(n82) );
  NANDN U115 ( .A(n555), .B(n82), .Z(n83) );
  NAND U116 ( .A(n81), .B(n83), .Z(n606) );
  NAND U117 ( .A(n397), .B(n398), .Z(n84) );
  XOR U118 ( .A(n397), .B(n398), .Z(n85) );
  NANDN U119 ( .A(n396), .B(n85), .Z(n86) );
  NAND U120 ( .A(n84), .B(n86), .Z(n416) );
  NAND U121 ( .A(n428), .B(n429), .Z(n87) );
  XOR U122 ( .A(n428), .B(n429), .Z(n88) );
  NANDN U123 ( .A(n427), .B(n88), .Z(n89) );
  NAND U124 ( .A(n87), .B(n89), .Z(n478) );
  NAND U125 ( .A(n269), .B(n270), .Z(n90) );
  XOR U126 ( .A(n269), .B(n270), .Z(n91) );
  NANDN U127 ( .A(n268), .B(n91), .Z(n92) );
  NAND U128 ( .A(n90), .B(n92), .Z(n288) );
  NAND U129 ( .A(n300), .B(n301), .Z(n93) );
  XOR U130 ( .A(n300), .B(n301), .Z(n94) );
  NANDN U131 ( .A(n299), .B(n94), .Z(n95) );
  NAND U132 ( .A(n93), .B(n95), .Z(n350) );
  XOR U133 ( .A(n827), .B(n826), .Z(n825) );
  XOR U134 ( .A(n699), .B(n698), .Z(n697) );
  XOR U135 ( .A(n571), .B(n570), .Z(n569) );
  XOR U136 ( .A(n443), .B(n442), .Z(n441) );
  XOR U137 ( .A(n315), .B(n314), .Z(n313) );
  NAND U138 ( .A(n776), .B(n774), .Z(n96) );
  XOR U139 ( .A(n776), .B(n774), .Z(n97) );
  NANDN U140 ( .A(n775), .B(n97), .Z(n98) );
  NAND U141 ( .A(n96), .B(n98), .Z(n782) );
  NAND U142 ( .A(n648), .B(n646), .Z(n99) );
  XOR U143 ( .A(n648), .B(n646), .Z(n100) );
  NANDN U144 ( .A(n647), .B(n100), .Z(n101) );
  NAND U145 ( .A(n99), .B(n101), .Z(n654) );
  NAND U146 ( .A(n520), .B(n518), .Z(n102) );
  XOR U147 ( .A(n520), .B(n518), .Z(n103) );
  NANDN U148 ( .A(n519), .B(n103), .Z(n104) );
  NAND U149 ( .A(n102), .B(n104), .Z(n526) );
  NAND U150 ( .A(n392), .B(n390), .Z(n105) );
  XOR U151 ( .A(n392), .B(n390), .Z(n106) );
  NANDN U152 ( .A(n391), .B(n106), .Z(n107) );
  NAND U153 ( .A(n105), .B(n107), .Z(n398) );
  NAND U154 ( .A(n264), .B(n262), .Z(n108) );
  XOR U155 ( .A(n264), .B(n262), .Z(n109) );
  NANDN U156 ( .A(n263), .B(n109), .Z(n110) );
  NAND U157 ( .A(n108), .B(n110), .Z(n270) );
  XOR U158 ( .A(n868), .B(n867), .Z(n866) );
  NANDN U159 ( .A(n859), .B(n860), .Z(n864) );
  XOR U160 ( .A(n740), .B(n739), .Z(n738) );
  NANDN U161 ( .A(n731), .B(n732), .Z(n736) );
  XOR U162 ( .A(n612), .B(n611), .Z(n610) );
  NANDN U163 ( .A(n603), .B(n604), .Z(n608) );
  XOR U164 ( .A(n484), .B(n483), .Z(n482) );
  NANDN U165 ( .A(n475), .B(n476), .Z(n480) );
  XOR U166 ( .A(n356), .B(n355), .Z(n354) );
  NANDN U167 ( .A(n347), .B(n348), .Z(n352) );
  NAND U168 ( .A(n754), .B(n752), .Z(n111) );
  XOR U169 ( .A(n754), .B(n752), .Z(n112) );
  NANDN U170 ( .A(n753), .B(n112), .Z(n113) );
  NAND U171 ( .A(n111), .B(n113), .Z(n768) );
  XOR U172 ( .A(n766), .B(n764), .Z(n114) );
  NANDN U173 ( .A(n765), .B(n114), .Z(n115) );
  NAND U174 ( .A(n766), .B(n764), .Z(n116) );
  AND U175 ( .A(n115), .B(n116), .Z(n784) );
  NAND U176 ( .A(n626), .B(n624), .Z(n117) );
  XOR U177 ( .A(n626), .B(n624), .Z(n118) );
  NANDN U178 ( .A(n625), .B(n118), .Z(n119) );
  NAND U179 ( .A(n117), .B(n119), .Z(n640) );
  XOR U180 ( .A(n638), .B(n636), .Z(n120) );
  NANDN U181 ( .A(n637), .B(n120), .Z(n121) );
  NAND U182 ( .A(n638), .B(n636), .Z(n122) );
  AND U183 ( .A(n121), .B(n122), .Z(n656) );
  NAND U184 ( .A(n498), .B(n496), .Z(n123) );
  XOR U185 ( .A(n498), .B(n496), .Z(n124) );
  NANDN U186 ( .A(n497), .B(n124), .Z(n125) );
  NAND U187 ( .A(n123), .B(n125), .Z(n512) );
  XOR U188 ( .A(n510), .B(n508), .Z(n126) );
  NANDN U189 ( .A(n509), .B(n126), .Z(n127) );
  NAND U190 ( .A(n510), .B(n508), .Z(n128) );
  AND U191 ( .A(n127), .B(n128), .Z(n528) );
  NAND U192 ( .A(n370), .B(n368), .Z(n129) );
  XOR U193 ( .A(n370), .B(n368), .Z(n130) );
  NANDN U194 ( .A(n369), .B(n130), .Z(n131) );
  NAND U195 ( .A(n129), .B(n131), .Z(n384) );
  XOR U196 ( .A(n382), .B(n380), .Z(n132) );
  NANDN U197 ( .A(n381), .B(n132), .Z(n133) );
  NAND U198 ( .A(n382), .B(n380), .Z(n134) );
  AND U199 ( .A(n133), .B(n134), .Z(n400) );
  NAND U200 ( .A(n242), .B(n240), .Z(n135) );
  XOR U201 ( .A(n242), .B(n240), .Z(n136) );
  NANDN U202 ( .A(n241), .B(n136), .Z(n137) );
  NAND U203 ( .A(n135), .B(n137), .Z(n256) );
  XOR U204 ( .A(n254), .B(n252), .Z(n138) );
  NANDN U205 ( .A(n253), .B(n138), .Z(n139) );
  NAND U206 ( .A(n254), .B(n252), .Z(n140) );
  AND U207 ( .A(n139), .B(n140), .Z(n272) );
  AND U208 ( .A(n870), .B(n869), .Z(n141) );
  NAND U209 ( .A(n864), .B(n863), .Z(n142) );
  XNOR U210 ( .A(n141), .B(n142), .Z(n143) );
  NAND U211 ( .A(n855), .B(n854), .Z(n144) );
  NAND U212 ( .A(n858), .B(n144), .Z(n145) );
  XNOR U213 ( .A(n143), .B(n145), .Z(n146) );
  NAND U214 ( .A(n827), .B(n826), .Z(n147) );
  NAND U215 ( .A(n828), .B(n829), .Z(n148) );
  AND U216 ( .A(n147), .B(n148), .Z(n149) );
  AND U217 ( .A(n853), .B(n852), .Z(n150) );
  XNOR U218 ( .A(n847), .B(n846), .Z(n151) );
  XNOR U219 ( .A(n150), .B(n151), .Z(n152) );
  XNOR U220 ( .A(n149), .B(n152), .Z(n153) );
  XNOR U221 ( .A(n146), .B(n153), .Z(n154) );
  NANDN U222 ( .A(n823), .B(n824), .Z(n155) );
  XNOR U223 ( .A(n823), .B(n824), .Z(n156) );
  NAND U224 ( .A(n825), .B(n156), .Z(n157) );
  AND U225 ( .A(n155), .B(n157), .Z(n158) );
  XNOR U226 ( .A(n154), .B(n158), .Z(N80) );
  AND U227 ( .A(n742), .B(n741), .Z(n159) );
  NAND U228 ( .A(n736), .B(n735), .Z(n160) );
  XNOR U229 ( .A(n159), .B(n160), .Z(n161) );
  NAND U230 ( .A(n727), .B(n726), .Z(n162) );
  NAND U231 ( .A(n730), .B(n162), .Z(n163) );
  XNOR U232 ( .A(n161), .B(n163), .Z(n164) );
  NAND U233 ( .A(n699), .B(n698), .Z(n165) );
  NAND U234 ( .A(n700), .B(n701), .Z(n166) );
  AND U235 ( .A(n165), .B(n166), .Z(n167) );
  AND U236 ( .A(n725), .B(n724), .Z(n168) );
  XNOR U237 ( .A(n719), .B(n718), .Z(n169) );
  XNOR U238 ( .A(n168), .B(n169), .Z(n170) );
  XNOR U239 ( .A(n167), .B(n170), .Z(n171) );
  XNOR U240 ( .A(n164), .B(n171), .Z(n172) );
  NANDN U241 ( .A(n695), .B(n696), .Z(n173) );
  XNOR U242 ( .A(n695), .B(n696), .Z(n174) );
  NAND U243 ( .A(n697), .B(n174), .Z(n175) );
  AND U244 ( .A(n173), .B(n175), .Z(n176) );
  XNOR U245 ( .A(n172), .B(n176), .Z(N64) );
  AND U246 ( .A(n614), .B(n613), .Z(n177) );
  NAND U247 ( .A(n608), .B(n607), .Z(n178) );
  XNOR U248 ( .A(n177), .B(n178), .Z(n179) );
  NAND U249 ( .A(n599), .B(n598), .Z(n180) );
  NAND U250 ( .A(n602), .B(n180), .Z(n181) );
  XNOR U251 ( .A(n179), .B(n181), .Z(n182) );
  NAND U252 ( .A(n571), .B(n570), .Z(n183) );
  NAND U253 ( .A(n572), .B(n573), .Z(n184) );
  AND U254 ( .A(n183), .B(n184), .Z(n185) );
  AND U255 ( .A(n597), .B(n596), .Z(n186) );
  XNOR U256 ( .A(n591), .B(n590), .Z(n187) );
  XNOR U257 ( .A(n186), .B(n187), .Z(n188) );
  XNOR U258 ( .A(n185), .B(n188), .Z(n189) );
  XNOR U259 ( .A(n182), .B(n189), .Z(n190) );
  NANDN U260 ( .A(n567), .B(n568), .Z(n191) );
  XNOR U261 ( .A(n567), .B(n568), .Z(n192) );
  NAND U262 ( .A(n569), .B(n192), .Z(n193) );
  AND U263 ( .A(n191), .B(n193), .Z(n194) );
  XNOR U264 ( .A(n190), .B(n194), .Z(N48) );
  AND U265 ( .A(n486), .B(n485), .Z(n195) );
  NAND U266 ( .A(n480), .B(n479), .Z(n196) );
  XNOR U267 ( .A(n195), .B(n196), .Z(n197) );
  NAND U268 ( .A(n471), .B(n470), .Z(n198) );
  NAND U269 ( .A(n474), .B(n198), .Z(n199) );
  XNOR U270 ( .A(n197), .B(n199), .Z(n200) );
  NAND U271 ( .A(n443), .B(n442), .Z(n201) );
  NAND U272 ( .A(n444), .B(n445), .Z(n202) );
  AND U273 ( .A(n201), .B(n202), .Z(n203) );
  AND U274 ( .A(n469), .B(n468), .Z(n204) );
  XNOR U275 ( .A(n463), .B(n462), .Z(n205) );
  XNOR U276 ( .A(n204), .B(n205), .Z(n206) );
  XNOR U277 ( .A(n203), .B(n206), .Z(n207) );
  XNOR U278 ( .A(n200), .B(n207), .Z(n208) );
  NANDN U279 ( .A(n439), .B(n440), .Z(n209) );
  XNOR U280 ( .A(n439), .B(n440), .Z(n210) );
  NAND U281 ( .A(n441), .B(n210), .Z(n211) );
  AND U282 ( .A(n209), .B(n211), .Z(n212) );
  XNOR U283 ( .A(n208), .B(n212), .Z(N32) );
  NAND U284 ( .A(n315), .B(n314), .Z(n213) );
  NAND U285 ( .A(n316), .B(n317), .Z(n214) );
  AND U286 ( .A(n213), .B(n214), .Z(n215) );
  AND U287 ( .A(n341), .B(n340), .Z(n216) );
  XNOR U288 ( .A(n335), .B(n334), .Z(n217) );
  XNOR U289 ( .A(n216), .B(n217), .Z(n218) );
  AND U290 ( .A(n358), .B(n357), .Z(n219) );
  NAND U291 ( .A(n352), .B(n351), .Z(n220) );
  XNOR U292 ( .A(n219), .B(n220), .Z(n221) );
  NAND U293 ( .A(n343), .B(n342), .Z(n222) );
  NAND U294 ( .A(n346), .B(n222), .Z(n223) );
  XNOR U295 ( .A(n221), .B(n223), .Z(n224) );
  XNOR U296 ( .A(n215), .B(n218), .Z(n225) );
  XNOR U297 ( .A(n224), .B(n225), .Z(n226) );
  NANDN U298 ( .A(n311), .B(n312), .Z(n227) );
  XNOR U299 ( .A(n311), .B(n312), .Z(n228) );
  NAND U300 ( .A(n313), .B(n228), .Z(n229) );
  AND U301 ( .A(n227), .B(n229), .Z(n230) );
  XNOR U302 ( .A(n226), .B(n230), .Z(N16) );
  AND U303 ( .A(x[32]), .B(y[160]), .Z(n231) );
  XOR U304 ( .A(n231), .B(o[0]), .Z(N9) );
  AND U305 ( .A(x[32]), .B(y[161]), .Z(n238) );
  XOR U306 ( .A(n238), .B(o[1]), .Z(n233) );
  NAND U307 ( .A(x[33]), .B(y[160]), .Z(n232) );
  XNOR U308 ( .A(n233), .B(n232), .Z(n235) );
  NAND U309 ( .A(n231), .B(o[0]), .Z(n234) );
  XNOR U310 ( .A(n235), .B(n234), .Z(N10) );
  NANDN U311 ( .A(n233), .B(n232), .Z(n237) );
  NAND U312 ( .A(n235), .B(n234), .Z(n236) );
  AND U313 ( .A(n237), .B(n236), .Z(n244) );
  AND U314 ( .A(x[32]), .B(y[162]), .Z(n249) );
  XNOR U315 ( .A(n249), .B(o[2]), .Z(n243) );
  XNOR U316 ( .A(n244), .B(n243), .Z(n246) );
  NAND U317 ( .A(y[161]), .B(x[33]), .Z(n241) );
  AND U318 ( .A(n238), .B(o[1]), .Z(n242) );
  AND U319 ( .A(y[160]), .B(x[34]), .Z(n240) );
  XNOR U320 ( .A(n242), .B(n240), .Z(n239) );
  XNOR U321 ( .A(n241), .B(n239), .Z(n245) );
  XNOR U322 ( .A(n246), .B(n245), .Z(N11) );
  NANDN U323 ( .A(n244), .B(n243), .Z(n248) );
  NAND U324 ( .A(n246), .B(n245), .Z(n247) );
  NAND U325 ( .A(n248), .B(n247), .Z(n255) );
  XNOR U326 ( .A(n256), .B(n255), .Z(n258) );
  NAND U327 ( .A(y[160]), .B(x[35]), .Z(n263) );
  AND U328 ( .A(n249), .B(o[2]), .Z(n264) );
  AND U329 ( .A(x[32]), .B(y[163]), .Z(n262) );
  XNOR U330 ( .A(n264), .B(n262), .Z(n250) );
  XNOR U331 ( .A(n263), .B(n250), .Z(n254) );
  NAND U332 ( .A(y[161]), .B(x[34]), .Z(n265) );
  XNOR U333 ( .A(o[3]), .B(n265), .Z(n253) );
  NAND U334 ( .A(x[33]), .B(y[162]), .Z(n252) );
  XOR U335 ( .A(n253), .B(n252), .Z(n251) );
  XNOR U336 ( .A(n254), .B(n251), .Z(n257) );
  XNOR U337 ( .A(n258), .B(n257), .Z(N12) );
  NANDN U338 ( .A(n256), .B(n255), .Z(n260) );
  NAND U339 ( .A(n258), .B(n257), .Z(n259) );
  NAND U340 ( .A(n260), .B(n259), .Z(n271) );
  XNOR U341 ( .A(n272), .B(n271), .Z(n274) );
  NAND U342 ( .A(y[162]), .B(x[34]), .Z(n280) );
  NAND U343 ( .A(y[161]), .B(x[35]), .Z(n283) );
  XNOR U344 ( .A(o[4]), .B(n283), .Z(n282) );
  AND U345 ( .A(x[33]), .B(y[163]), .Z(n281) );
  XNOR U346 ( .A(n282), .B(n281), .Z(n261) );
  XNOR U347 ( .A(n280), .B(n261), .Z(n268) );
  NAND U348 ( .A(y[160]), .B(x[36]), .Z(n278) );
  ANDN U349 ( .B(o[3]), .A(n265), .Z(n277) );
  NAND U350 ( .A(x[32]), .B(y[164]), .Z(n279) );
  XOR U351 ( .A(n277), .B(n279), .Z(n266) );
  XOR U352 ( .A(n278), .B(n266), .Z(n269) );
  XNOR U353 ( .A(n270), .B(n269), .Z(n267) );
  XNOR U354 ( .A(n268), .B(n267), .Z(n273) );
  XNOR U355 ( .A(n274), .B(n273), .Z(N13) );
  NANDN U356 ( .A(n272), .B(n271), .Z(n276) );
  NAND U357 ( .A(n274), .B(n273), .Z(n275) );
  NAND U358 ( .A(n276), .B(n275), .Z(n287) );
  XNOR U359 ( .A(n288), .B(n287), .Z(n290) );
  XNOR U360 ( .A(n293), .B(n294), .Z(n296) );
  NAND U361 ( .A(y[160]), .B(x[37]), .Z(n308) );
  ANDN U362 ( .B(o[4]), .A(n283), .Z(n309) );
  AND U363 ( .A(x[32]), .B(y[165]), .Z(n307) );
  XNOR U364 ( .A(n309), .B(n307), .Z(n284) );
  XOR U365 ( .A(n308), .B(n284), .Z(n301) );
  NAND U366 ( .A(x[33]), .B(y[164]), .Z(n302) );
  NAND U367 ( .A(y[161]), .B(x[36]), .Z(n305) );
  XNOR U368 ( .A(o[5]), .B(n305), .Z(n304) );
  AND U369 ( .A(y[162]), .B(x[35]), .Z(n303) );
  XNOR U370 ( .A(n304), .B(n303), .Z(n285) );
  XOR U371 ( .A(n302), .B(n285), .Z(n300) );
  NAND U372 ( .A(x[34]), .B(y[163]), .Z(n299) );
  XOR U373 ( .A(n300), .B(n299), .Z(n286) );
  XOR U374 ( .A(n301), .B(n286), .Z(n295) );
  XOR U375 ( .A(n296), .B(n295), .Z(n289) );
  XNOR U376 ( .A(n290), .B(n289), .Z(N14) );
  NANDN U377 ( .A(n288), .B(n287), .Z(n292) );
  NAND U378 ( .A(n290), .B(n289), .Z(n291) );
  NAND U379 ( .A(n292), .B(n291), .Z(n356) );
  NANDN U380 ( .A(n294), .B(n293), .Z(n298) );
  NAND U381 ( .A(n296), .B(n295), .Z(n297) );
  NAND U382 ( .A(n298), .B(n297), .Z(n355) );
  XOR U383 ( .A(n350), .B(n349), .Z(n348) );
  NAND U384 ( .A(y[160]), .B(x[38]), .Z(n337) );
  ANDN U385 ( .B(o[5]), .A(n305), .Z(n336) );
  NAND U386 ( .A(x[32]), .B(y[166]), .Z(n339) );
  XOR U387 ( .A(n336), .B(n339), .Z(n306) );
  XNOR U388 ( .A(n337), .B(n306), .Z(n311) );
  AND U389 ( .A(x[34]), .B(y[164]), .Z(n317) );
  AND U390 ( .A(y[163]), .B(x[35]), .Z(n316) );
  XOR U391 ( .A(n317), .B(n316), .Z(n314) );
  AND U392 ( .A(y[161]), .B(x[37]), .Z(n318) );
  XOR U393 ( .A(n318), .B(o[6]), .Z(n342) );
  NAND U394 ( .A(x[33]), .B(y[165]), .Z(n345) );
  AND U395 ( .A(y[162]), .B(x[36]), .Z(n343) );
  XNOR U396 ( .A(n313), .B(n312), .Z(n310) );
  XOR U397 ( .A(n311), .B(n310), .Z(n347) );
  XNOR U398 ( .A(n348), .B(n347), .Z(n353) );
  XNOR U399 ( .A(n354), .B(n353), .Z(N15) );
  AND U400 ( .A(x[39]), .B(y[160]), .Z(n327) );
  AND U401 ( .A(n318), .B(o[6]), .Z(n325) );
  AND U402 ( .A(x[36]), .B(y[163]), .Z(n323) );
  AND U403 ( .A(y[164]), .B(x[35]), .Z(n320) );
  NAND U404 ( .A(y[165]), .B(x[34]), .Z(n319) );
  XNOR U405 ( .A(n320), .B(n319), .Z(n321) );
  XNOR U406 ( .A(o[7]), .B(n321), .Z(n322) );
  XNOR U407 ( .A(n323), .B(n322), .Z(n324) );
  XNOR U408 ( .A(n325), .B(n324), .Z(n326) );
  XNOR U409 ( .A(n327), .B(n326), .Z(n335) );
  AND U410 ( .A(x[37]), .B(y[162]), .Z(n329) );
  NAND U411 ( .A(x[38]), .B(y[161]), .Z(n328) );
  XNOR U412 ( .A(n329), .B(n328), .Z(n333) );
  AND U413 ( .A(y[166]), .B(x[33]), .Z(n331) );
  NAND U414 ( .A(y[167]), .B(x[32]), .Z(n330) );
  XNOR U415 ( .A(n331), .B(n330), .Z(n332) );
  XNOR U416 ( .A(n333), .B(n332), .Z(n334) );
  NANDN U417 ( .A(n337), .B(n336), .Z(n341) );
  ANDN U418 ( .B(n337), .A(n336), .Z(n338) );
  OR U419 ( .A(n339), .B(n338), .Z(n340) );
  NOR U420 ( .A(n343), .B(n342), .Z(n344) );
  OR U421 ( .A(n345), .B(n344), .Z(n346) );
  OR U422 ( .A(n350), .B(n349), .Z(n351) );
  NAND U423 ( .A(n354), .B(n353), .Z(n358) );
  NAND U424 ( .A(n356), .B(n355), .Z(n357) );
  AND U425 ( .A(x[32]), .B(y[168]), .Z(n359) );
  XOR U426 ( .A(n359), .B(o[8]), .Z(N25) );
  AND U427 ( .A(x[32]), .B(y[169]), .Z(n366) );
  XOR U428 ( .A(n366), .B(o[9]), .Z(n361) );
  NAND U429 ( .A(x[33]), .B(y[168]), .Z(n360) );
  XNOR U430 ( .A(n361), .B(n360), .Z(n363) );
  NAND U431 ( .A(n359), .B(o[8]), .Z(n362) );
  XNOR U432 ( .A(n363), .B(n362), .Z(N26) );
  NANDN U433 ( .A(n361), .B(n360), .Z(n365) );
  NAND U434 ( .A(n363), .B(n362), .Z(n364) );
  AND U435 ( .A(n365), .B(n364), .Z(n372) );
  AND U436 ( .A(x[32]), .B(y[170]), .Z(n377) );
  XNOR U437 ( .A(n377), .B(o[10]), .Z(n371) );
  XNOR U438 ( .A(n372), .B(n371), .Z(n374) );
  NAND U439 ( .A(x[33]), .B(y[169]), .Z(n369) );
  AND U440 ( .A(n366), .B(o[9]), .Z(n370) );
  AND U441 ( .A(x[34]), .B(y[168]), .Z(n368) );
  XNOR U442 ( .A(n370), .B(n368), .Z(n367) );
  XNOR U443 ( .A(n369), .B(n367), .Z(n373) );
  XNOR U444 ( .A(n374), .B(n373), .Z(N27) );
  NANDN U445 ( .A(n372), .B(n371), .Z(n376) );
  NAND U446 ( .A(n374), .B(n373), .Z(n375) );
  NAND U447 ( .A(n376), .B(n375), .Z(n383) );
  XNOR U448 ( .A(n384), .B(n383), .Z(n386) );
  NAND U449 ( .A(x[35]), .B(y[168]), .Z(n391) );
  AND U450 ( .A(n377), .B(o[10]), .Z(n392) );
  AND U451 ( .A(x[32]), .B(y[171]), .Z(n390) );
  XNOR U452 ( .A(n392), .B(n390), .Z(n378) );
  XNOR U453 ( .A(n391), .B(n378), .Z(n382) );
  NAND U454 ( .A(x[34]), .B(y[169]), .Z(n393) );
  XNOR U455 ( .A(o[11]), .B(n393), .Z(n381) );
  NAND U456 ( .A(x[33]), .B(y[170]), .Z(n380) );
  XOR U457 ( .A(n381), .B(n380), .Z(n379) );
  XNOR U458 ( .A(n382), .B(n379), .Z(n385) );
  XNOR U459 ( .A(n386), .B(n385), .Z(N28) );
  NANDN U460 ( .A(n384), .B(n383), .Z(n388) );
  NAND U461 ( .A(n386), .B(n385), .Z(n387) );
  NAND U462 ( .A(n388), .B(n387), .Z(n399) );
  XNOR U463 ( .A(n400), .B(n399), .Z(n402) );
  NAND U464 ( .A(x[34]), .B(y[170]), .Z(n408) );
  NAND U465 ( .A(x[35]), .B(y[169]), .Z(n411) );
  XNOR U466 ( .A(o[12]), .B(n411), .Z(n410) );
  AND U467 ( .A(x[33]), .B(y[171]), .Z(n409) );
  XNOR U468 ( .A(n410), .B(n409), .Z(n389) );
  XNOR U469 ( .A(n408), .B(n389), .Z(n396) );
  NAND U470 ( .A(x[36]), .B(y[168]), .Z(n406) );
  ANDN U471 ( .B(o[11]), .A(n393), .Z(n405) );
  NAND U472 ( .A(x[32]), .B(y[172]), .Z(n407) );
  XOR U473 ( .A(n405), .B(n407), .Z(n394) );
  XOR U474 ( .A(n406), .B(n394), .Z(n397) );
  XNOR U475 ( .A(n398), .B(n397), .Z(n395) );
  XNOR U476 ( .A(n396), .B(n395), .Z(n401) );
  XNOR U477 ( .A(n402), .B(n401), .Z(N29) );
  NANDN U478 ( .A(n400), .B(n399), .Z(n404) );
  NAND U479 ( .A(n402), .B(n401), .Z(n403) );
  NAND U480 ( .A(n404), .B(n403), .Z(n415) );
  XNOR U481 ( .A(n416), .B(n415), .Z(n418) );
  XNOR U482 ( .A(n421), .B(n422), .Z(n424) );
  NAND U483 ( .A(x[37]), .B(y[168]), .Z(n436) );
  ANDN U484 ( .B(o[12]), .A(n411), .Z(n437) );
  AND U485 ( .A(x[32]), .B(y[173]), .Z(n435) );
  XNOR U486 ( .A(n437), .B(n435), .Z(n412) );
  XOR U487 ( .A(n436), .B(n412), .Z(n429) );
  NAND U488 ( .A(x[33]), .B(y[172]), .Z(n430) );
  NAND U489 ( .A(x[36]), .B(y[169]), .Z(n433) );
  XNOR U490 ( .A(o[13]), .B(n433), .Z(n432) );
  AND U491 ( .A(x[35]), .B(y[170]), .Z(n431) );
  XNOR U492 ( .A(n432), .B(n431), .Z(n413) );
  XOR U493 ( .A(n430), .B(n413), .Z(n428) );
  NAND U494 ( .A(x[34]), .B(y[171]), .Z(n427) );
  XOR U495 ( .A(n428), .B(n427), .Z(n414) );
  XOR U496 ( .A(n429), .B(n414), .Z(n423) );
  XOR U497 ( .A(n424), .B(n423), .Z(n417) );
  XNOR U498 ( .A(n418), .B(n417), .Z(N30) );
  NANDN U499 ( .A(n416), .B(n415), .Z(n420) );
  NAND U500 ( .A(n418), .B(n417), .Z(n419) );
  NAND U501 ( .A(n420), .B(n419), .Z(n484) );
  NANDN U502 ( .A(n422), .B(n421), .Z(n426) );
  NAND U503 ( .A(n424), .B(n423), .Z(n425) );
  NAND U504 ( .A(n426), .B(n425), .Z(n483) );
  XOR U505 ( .A(n478), .B(n477), .Z(n476) );
  NAND U506 ( .A(x[38]), .B(y[168]), .Z(n465) );
  ANDN U507 ( .B(o[13]), .A(n433), .Z(n464) );
  NAND U508 ( .A(x[32]), .B(y[174]), .Z(n467) );
  XOR U509 ( .A(n464), .B(n467), .Z(n434) );
  XNOR U510 ( .A(n465), .B(n434), .Z(n439) );
  AND U511 ( .A(x[34]), .B(y[172]), .Z(n445) );
  AND U512 ( .A(x[35]), .B(y[171]), .Z(n444) );
  XOR U513 ( .A(n445), .B(n444), .Z(n442) );
  AND U514 ( .A(x[37]), .B(y[169]), .Z(n446) );
  XOR U515 ( .A(n446), .B(o[14]), .Z(n470) );
  NAND U516 ( .A(x[33]), .B(y[173]), .Z(n473) );
  AND U517 ( .A(x[36]), .B(y[170]), .Z(n471) );
  XNOR U518 ( .A(n441), .B(n440), .Z(n438) );
  XOR U519 ( .A(n439), .B(n438), .Z(n475) );
  XNOR U520 ( .A(n476), .B(n475), .Z(n481) );
  XNOR U521 ( .A(n482), .B(n481), .Z(N31) );
  AND U522 ( .A(y[175]), .B(x[32]), .Z(n455) );
  AND U523 ( .A(n446), .B(o[14]), .Z(n453) );
  AND U524 ( .A(y[171]), .B(x[36]), .Z(n451) );
  AND U525 ( .A(y[172]), .B(x[35]), .Z(n448) );
  NAND U526 ( .A(y[173]), .B(x[34]), .Z(n447) );
  XNOR U527 ( .A(n448), .B(n447), .Z(n449) );
  XNOR U528 ( .A(o[15]), .B(n449), .Z(n450) );
  XNOR U529 ( .A(n451), .B(n450), .Z(n452) );
  XNOR U530 ( .A(n453), .B(n452), .Z(n454) );
  XNOR U531 ( .A(n455), .B(n454), .Z(n463) );
  AND U532 ( .A(y[169]), .B(x[38]), .Z(n457) );
  NAND U533 ( .A(y[170]), .B(x[37]), .Z(n456) );
  XNOR U534 ( .A(n457), .B(n456), .Z(n461) );
  AND U535 ( .A(y[168]), .B(x[39]), .Z(n459) );
  NAND U536 ( .A(y[174]), .B(x[33]), .Z(n458) );
  XNOR U537 ( .A(n459), .B(n458), .Z(n460) );
  XNOR U538 ( .A(n461), .B(n460), .Z(n462) );
  NANDN U539 ( .A(n465), .B(n464), .Z(n469) );
  ANDN U540 ( .B(n465), .A(n464), .Z(n466) );
  OR U541 ( .A(n467), .B(n466), .Z(n468) );
  NOR U542 ( .A(n471), .B(n470), .Z(n472) );
  OR U543 ( .A(n473), .B(n472), .Z(n474) );
  OR U544 ( .A(n478), .B(n477), .Z(n479) );
  NAND U545 ( .A(n482), .B(n481), .Z(n486) );
  NAND U546 ( .A(n484), .B(n483), .Z(n485) );
  AND U547 ( .A(x[32]), .B(y[176]), .Z(n487) );
  XOR U548 ( .A(n487), .B(o[16]), .Z(N41) );
  AND U549 ( .A(x[32]), .B(y[177]), .Z(n494) );
  XOR U550 ( .A(n494), .B(o[17]), .Z(n489) );
  NAND U551 ( .A(x[33]), .B(y[176]), .Z(n488) );
  XNOR U552 ( .A(n489), .B(n488), .Z(n491) );
  NAND U553 ( .A(n487), .B(o[16]), .Z(n490) );
  XNOR U554 ( .A(n491), .B(n490), .Z(N42) );
  NANDN U555 ( .A(n489), .B(n488), .Z(n493) );
  NAND U556 ( .A(n491), .B(n490), .Z(n492) );
  AND U557 ( .A(n493), .B(n492), .Z(n500) );
  AND U558 ( .A(x[32]), .B(y[178]), .Z(n505) );
  XNOR U559 ( .A(n505), .B(o[18]), .Z(n499) );
  XNOR U560 ( .A(n500), .B(n499), .Z(n502) );
  NAND U561 ( .A(x[33]), .B(y[177]), .Z(n497) );
  AND U562 ( .A(n494), .B(o[17]), .Z(n498) );
  AND U563 ( .A(x[34]), .B(y[176]), .Z(n496) );
  XNOR U564 ( .A(n498), .B(n496), .Z(n495) );
  XNOR U565 ( .A(n497), .B(n495), .Z(n501) );
  XNOR U566 ( .A(n502), .B(n501), .Z(N43) );
  NANDN U567 ( .A(n500), .B(n499), .Z(n504) );
  NAND U568 ( .A(n502), .B(n501), .Z(n503) );
  NAND U569 ( .A(n504), .B(n503), .Z(n511) );
  XNOR U570 ( .A(n512), .B(n511), .Z(n514) );
  NAND U571 ( .A(x[35]), .B(y[176]), .Z(n519) );
  AND U572 ( .A(n505), .B(o[18]), .Z(n520) );
  AND U573 ( .A(x[32]), .B(y[179]), .Z(n518) );
  XNOR U574 ( .A(n520), .B(n518), .Z(n506) );
  XNOR U575 ( .A(n519), .B(n506), .Z(n510) );
  NAND U576 ( .A(x[34]), .B(y[177]), .Z(n521) );
  XNOR U577 ( .A(o[19]), .B(n521), .Z(n509) );
  NAND U578 ( .A(x[33]), .B(y[178]), .Z(n508) );
  XOR U579 ( .A(n509), .B(n508), .Z(n507) );
  XNOR U580 ( .A(n510), .B(n507), .Z(n513) );
  XNOR U581 ( .A(n514), .B(n513), .Z(N44) );
  NANDN U582 ( .A(n512), .B(n511), .Z(n516) );
  NAND U583 ( .A(n514), .B(n513), .Z(n515) );
  NAND U584 ( .A(n516), .B(n515), .Z(n527) );
  XNOR U585 ( .A(n528), .B(n527), .Z(n530) );
  NAND U586 ( .A(x[34]), .B(y[178]), .Z(n536) );
  NAND U587 ( .A(x[35]), .B(y[177]), .Z(n539) );
  XNOR U588 ( .A(o[20]), .B(n539), .Z(n538) );
  AND U589 ( .A(x[33]), .B(y[179]), .Z(n537) );
  XNOR U590 ( .A(n538), .B(n537), .Z(n517) );
  XNOR U591 ( .A(n536), .B(n517), .Z(n524) );
  NAND U592 ( .A(x[36]), .B(y[176]), .Z(n534) );
  ANDN U593 ( .B(o[19]), .A(n521), .Z(n533) );
  NAND U594 ( .A(x[32]), .B(y[180]), .Z(n535) );
  XOR U595 ( .A(n533), .B(n535), .Z(n522) );
  XOR U596 ( .A(n534), .B(n522), .Z(n525) );
  XNOR U597 ( .A(n526), .B(n525), .Z(n523) );
  XNOR U598 ( .A(n524), .B(n523), .Z(n529) );
  XNOR U599 ( .A(n530), .B(n529), .Z(N45) );
  NANDN U600 ( .A(n528), .B(n527), .Z(n532) );
  NAND U601 ( .A(n530), .B(n529), .Z(n531) );
  NAND U602 ( .A(n532), .B(n531), .Z(n543) );
  XNOR U603 ( .A(n544), .B(n543), .Z(n546) );
  XNOR U604 ( .A(n549), .B(n550), .Z(n552) );
  NAND U605 ( .A(x[37]), .B(y[176]), .Z(n564) );
  ANDN U606 ( .B(o[20]), .A(n539), .Z(n565) );
  AND U607 ( .A(x[32]), .B(y[181]), .Z(n563) );
  XNOR U608 ( .A(n565), .B(n563), .Z(n540) );
  XOR U609 ( .A(n564), .B(n540), .Z(n557) );
  NAND U610 ( .A(x[33]), .B(y[180]), .Z(n558) );
  NAND U611 ( .A(x[36]), .B(y[177]), .Z(n561) );
  XNOR U612 ( .A(o[21]), .B(n561), .Z(n560) );
  AND U613 ( .A(x[35]), .B(y[178]), .Z(n559) );
  XNOR U614 ( .A(n560), .B(n559), .Z(n541) );
  XOR U615 ( .A(n558), .B(n541), .Z(n556) );
  NAND U616 ( .A(x[34]), .B(y[179]), .Z(n555) );
  XOR U617 ( .A(n556), .B(n555), .Z(n542) );
  XOR U618 ( .A(n557), .B(n542), .Z(n551) );
  XOR U619 ( .A(n552), .B(n551), .Z(n545) );
  XNOR U620 ( .A(n546), .B(n545), .Z(N46) );
  NANDN U621 ( .A(n544), .B(n543), .Z(n548) );
  NAND U622 ( .A(n546), .B(n545), .Z(n547) );
  NAND U623 ( .A(n548), .B(n547), .Z(n612) );
  NANDN U624 ( .A(n550), .B(n549), .Z(n554) );
  NAND U625 ( .A(n552), .B(n551), .Z(n553) );
  NAND U626 ( .A(n554), .B(n553), .Z(n611) );
  XOR U627 ( .A(n606), .B(n605), .Z(n604) );
  NAND U628 ( .A(x[38]), .B(y[176]), .Z(n593) );
  ANDN U629 ( .B(o[21]), .A(n561), .Z(n592) );
  NAND U630 ( .A(x[32]), .B(y[182]), .Z(n595) );
  XOR U631 ( .A(n592), .B(n595), .Z(n562) );
  XNOR U632 ( .A(n593), .B(n562), .Z(n567) );
  AND U633 ( .A(x[34]), .B(y[180]), .Z(n573) );
  AND U634 ( .A(x[35]), .B(y[179]), .Z(n572) );
  XOR U635 ( .A(n573), .B(n572), .Z(n570) );
  AND U636 ( .A(x[37]), .B(y[177]), .Z(n574) );
  XOR U637 ( .A(n574), .B(o[22]), .Z(n598) );
  NAND U638 ( .A(x[33]), .B(y[181]), .Z(n601) );
  AND U639 ( .A(x[36]), .B(y[178]), .Z(n599) );
  XNOR U640 ( .A(n569), .B(n568), .Z(n566) );
  XOR U641 ( .A(n567), .B(n566), .Z(n603) );
  XNOR U642 ( .A(n604), .B(n603), .Z(n609) );
  XNOR U643 ( .A(n610), .B(n609), .Z(N47) );
  AND U644 ( .A(y[183]), .B(x[32]), .Z(n583) );
  AND U645 ( .A(n574), .B(o[22]), .Z(n581) );
  AND U646 ( .A(y[179]), .B(x[36]), .Z(n579) );
  AND U647 ( .A(y[180]), .B(x[35]), .Z(n576) );
  NAND U648 ( .A(y[181]), .B(x[34]), .Z(n575) );
  XNOR U649 ( .A(n576), .B(n575), .Z(n577) );
  XNOR U650 ( .A(o[23]), .B(n577), .Z(n578) );
  XNOR U651 ( .A(n579), .B(n578), .Z(n580) );
  XNOR U652 ( .A(n581), .B(n580), .Z(n582) );
  XNOR U653 ( .A(n583), .B(n582), .Z(n591) );
  AND U654 ( .A(y[177]), .B(x[38]), .Z(n585) );
  NAND U655 ( .A(y[178]), .B(x[37]), .Z(n584) );
  XNOR U656 ( .A(n585), .B(n584), .Z(n589) );
  AND U657 ( .A(y[176]), .B(x[39]), .Z(n587) );
  NAND U658 ( .A(y[182]), .B(x[33]), .Z(n586) );
  XNOR U659 ( .A(n587), .B(n586), .Z(n588) );
  XNOR U660 ( .A(n589), .B(n588), .Z(n590) );
  NANDN U661 ( .A(n593), .B(n592), .Z(n597) );
  ANDN U662 ( .B(n593), .A(n592), .Z(n594) );
  OR U663 ( .A(n595), .B(n594), .Z(n596) );
  NOR U664 ( .A(n599), .B(n598), .Z(n600) );
  OR U665 ( .A(n601), .B(n600), .Z(n602) );
  OR U666 ( .A(n606), .B(n605), .Z(n607) );
  NAND U667 ( .A(n610), .B(n609), .Z(n614) );
  NAND U668 ( .A(n612), .B(n611), .Z(n613) );
  AND U669 ( .A(x[32]), .B(y[184]), .Z(n615) );
  XOR U670 ( .A(n615), .B(o[24]), .Z(N57) );
  AND U671 ( .A(x[32]), .B(y[185]), .Z(n622) );
  XOR U672 ( .A(n622), .B(o[25]), .Z(n617) );
  NAND U673 ( .A(x[33]), .B(y[184]), .Z(n616) );
  XNOR U674 ( .A(n617), .B(n616), .Z(n619) );
  NAND U675 ( .A(n615), .B(o[24]), .Z(n618) );
  XNOR U676 ( .A(n619), .B(n618), .Z(N58) );
  NANDN U677 ( .A(n617), .B(n616), .Z(n621) );
  NAND U678 ( .A(n619), .B(n618), .Z(n620) );
  AND U679 ( .A(n621), .B(n620), .Z(n628) );
  AND U680 ( .A(x[32]), .B(y[186]), .Z(n633) );
  XNOR U681 ( .A(n633), .B(o[26]), .Z(n627) );
  XNOR U682 ( .A(n628), .B(n627), .Z(n630) );
  NAND U683 ( .A(x[33]), .B(y[185]), .Z(n625) );
  AND U684 ( .A(n622), .B(o[25]), .Z(n626) );
  AND U685 ( .A(x[34]), .B(y[184]), .Z(n624) );
  XNOR U686 ( .A(n626), .B(n624), .Z(n623) );
  XNOR U687 ( .A(n625), .B(n623), .Z(n629) );
  XNOR U688 ( .A(n630), .B(n629), .Z(N59) );
  NANDN U689 ( .A(n628), .B(n627), .Z(n632) );
  NAND U690 ( .A(n630), .B(n629), .Z(n631) );
  NAND U691 ( .A(n632), .B(n631), .Z(n639) );
  XNOR U692 ( .A(n640), .B(n639), .Z(n642) );
  NAND U693 ( .A(x[35]), .B(y[184]), .Z(n647) );
  AND U694 ( .A(n633), .B(o[26]), .Z(n648) );
  AND U695 ( .A(x[32]), .B(y[187]), .Z(n646) );
  XNOR U696 ( .A(n648), .B(n646), .Z(n634) );
  XNOR U697 ( .A(n647), .B(n634), .Z(n638) );
  NAND U698 ( .A(x[34]), .B(y[185]), .Z(n649) );
  XNOR U699 ( .A(o[27]), .B(n649), .Z(n637) );
  NAND U700 ( .A(x[33]), .B(y[186]), .Z(n636) );
  XOR U701 ( .A(n637), .B(n636), .Z(n635) );
  XNOR U702 ( .A(n638), .B(n635), .Z(n641) );
  XNOR U703 ( .A(n642), .B(n641), .Z(N60) );
  NANDN U704 ( .A(n640), .B(n639), .Z(n644) );
  NAND U705 ( .A(n642), .B(n641), .Z(n643) );
  NAND U706 ( .A(n644), .B(n643), .Z(n655) );
  XNOR U707 ( .A(n656), .B(n655), .Z(n658) );
  NAND U708 ( .A(x[34]), .B(y[186]), .Z(n664) );
  NAND U709 ( .A(x[35]), .B(y[185]), .Z(n667) );
  XNOR U710 ( .A(o[28]), .B(n667), .Z(n666) );
  AND U711 ( .A(x[33]), .B(y[187]), .Z(n665) );
  XNOR U712 ( .A(n666), .B(n665), .Z(n645) );
  XNOR U713 ( .A(n664), .B(n645), .Z(n652) );
  NAND U714 ( .A(x[36]), .B(y[184]), .Z(n662) );
  ANDN U715 ( .B(o[27]), .A(n649), .Z(n661) );
  NAND U716 ( .A(x[32]), .B(y[188]), .Z(n663) );
  XOR U717 ( .A(n661), .B(n663), .Z(n650) );
  XOR U718 ( .A(n662), .B(n650), .Z(n653) );
  XNOR U719 ( .A(n654), .B(n653), .Z(n651) );
  XNOR U720 ( .A(n652), .B(n651), .Z(n657) );
  XNOR U721 ( .A(n658), .B(n657), .Z(N61) );
  NANDN U722 ( .A(n656), .B(n655), .Z(n660) );
  NAND U723 ( .A(n658), .B(n657), .Z(n659) );
  NAND U724 ( .A(n660), .B(n659), .Z(n671) );
  XNOR U725 ( .A(n672), .B(n671), .Z(n674) );
  XNOR U726 ( .A(n677), .B(n678), .Z(n680) );
  NAND U727 ( .A(x[37]), .B(y[184]), .Z(n692) );
  ANDN U728 ( .B(o[28]), .A(n667), .Z(n693) );
  AND U729 ( .A(x[32]), .B(y[189]), .Z(n691) );
  XNOR U730 ( .A(n693), .B(n691), .Z(n668) );
  XOR U731 ( .A(n692), .B(n668), .Z(n685) );
  NAND U732 ( .A(x[33]), .B(y[188]), .Z(n686) );
  NAND U733 ( .A(x[36]), .B(y[185]), .Z(n689) );
  XNOR U734 ( .A(o[29]), .B(n689), .Z(n688) );
  AND U735 ( .A(x[35]), .B(y[186]), .Z(n687) );
  XNOR U736 ( .A(n688), .B(n687), .Z(n669) );
  XOR U737 ( .A(n686), .B(n669), .Z(n684) );
  NAND U738 ( .A(x[34]), .B(y[187]), .Z(n683) );
  XOR U739 ( .A(n684), .B(n683), .Z(n670) );
  XOR U740 ( .A(n685), .B(n670), .Z(n679) );
  XOR U741 ( .A(n680), .B(n679), .Z(n673) );
  XNOR U742 ( .A(n674), .B(n673), .Z(N62) );
  NANDN U743 ( .A(n672), .B(n671), .Z(n676) );
  NAND U744 ( .A(n674), .B(n673), .Z(n675) );
  NAND U745 ( .A(n676), .B(n675), .Z(n740) );
  NANDN U746 ( .A(n678), .B(n677), .Z(n682) );
  NAND U747 ( .A(n680), .B(n679), .Z(n681) );
  NAND U748 ( .A(n682), .B(n681), .Z(n739) );
  XOR U749 ( .A(n734), .B(n733), .Z(n732) );
  NAND U750 ( .A(x[38]), .B(y[184]), .Z(n721) );
  ANDN U751 ( .B(o[29]), .A(n689), .Z(n720) );
  NAND U752 ( .A(x[32]), .B(y[190]), .Z(n723) );
  XOR U753 ( .A(n720), .B(n723), .Z(n690) );
  XNOR U754 ( .A(n721), .B(n690), .Z(n695) );
  AND U755 ( .A(x[34]), .B(y[188]), .Z(n701) );
  AND U756 ( .A(x[35]), .B(y[187]), .Z(n700) );
  XOR U757 ( .A(n701), .B(n700), .Z(n698) );
  AND U758 ( .A(x[37]), .B(y[185]), .Z(n702) );
  XOR U759 ( .A(n702), .B(o[30]), .Z(n726) );
  NAND U760 ( .A(x[33]), .B(y[189]), .Z(n729) );
  AND U761 ( .A(x[36]), .B(y[186]), .Z(n727) );
  XNOR U762 ( .A(n697), .B(n696), .Z(n694) );
  XOR U763 ( .A(n695), .B(n694), .Z(n731) );
  XNOR U764 ( .A(n732), .B(n731), .Z(n737) );
  XNOR U765 ( .A(n738), .B(n737), .Z(N63) );
  AND U766 ( .A(y[191]), .B(x[32]), .Z(n711) );
  AND U767 ( .A(n702), .B(o[30]), .Z(n709) );
  AND U768 ( .A(y[187]), .B(x[36]), .Z(n707) );
  AND U769 ( .A(y[188]), .B(x[35]), .Z(n704) );
  NAND U770 ( .A(y[189]), .B(x[34]), .Z(n703) );
  XNOR U771 ( .A(n704), .B(n703), .Z(n705) );
  XNOR U772 ( .A(o[31]), .B(n705), .Z(n706) );
  XNOR U773 ( .A(n707), .B(n706), .Z(n708) );
  XNOR U774 ( .A(n709), .B(n708), .Z(n710) );
  XNOR U775 ( .A(n711), .B(n710), .Z(n719) );
  AND U776 ( .A(y[185]), .B(x[38]), .Z(n713) );
  NAND U777 ( .A(y[186]), .B(x[37]), .Z(n712) );
  XNOR U778 ( .A(n713), .B(n712), .Z(n717) );
  AND U779 ( .A(y[184]), .B(x[39]), .Z(n715) );
  NAND U780 ( .A(y[190]), .B(x[33]), .Z(n714) );
  XNOR U781 ( .A(n715), .B(n714), .Z(n716) );
  XNOR U782 ( .A(n717), .B(n716), .Z(n718) );
  NANDN U783 ( .A(n721), .B(n720), .Z(n725) );
  ANDN U784 ( .B(n721), .A(n720), .Z(n722) );
  OR U785 ( .A(n723), .B(n722), .Z(n724) );
  NOR U786 ( .A(n727), .B(n726), .Z(n728) );
  OR U787 ( .A(n729), .B(n728), .Z(n730) );
  OR U788 ( .A(n734), .B(n733), .Z(n735) );
  NAND U789 ( .A(n738), .B(n737), .Z(n742) );
  NAND U790 ( .A(n740), .B(n739), .Z(n741) );
  AND U791 ( .A(x[32]), .B(y[192]), .Z(n743) );
  XOR U792 ( .A(n743), .B(o[32]), .Z(N73) );
  AND U793 ( .A(x[32]), .B(y[193]), .Z(n750) );
  XOR U794 ( .A(n750), .B(o[33]), .Z(n745) );
  NAND U795 ( .A(x[33]), .B(y[192]), .Z(n744) );
  XNOR U796 ( .A(n745), .B(n744), .Z(n747) );
  NAND U797 ( .A(n743), .B(o[32]), .Z(n746) );
  XNOR U798 ( .A(n747), .B(n746), .Z(N74) );
  NANDN U799 ( .A(n745), .B(n744), .Z(n749) );
  NAND U800 ( .A(n747), .B(n746), .Z(n748) );
  AND U801 ( .A(n749), .B(n748), .Z(n756) );
  AND U802 ( .A(x[32]), .B(y[194]), .Z(n761) );
  XNOR U803 ( .A(n761), .B(o[34]), .Z(n755) );
  XNOR U804 ( .A(n756), .B(n755), .Z(n758) );
  NAND U805 ( .A(x[33]), .B(y[193]), .Z(n753) );
  AND U806 ( .A(n750), .B(o[33]), .Z(n754) );
  AND U807 ( .A(x[34]), .B(y[192]), .Z(n752) );
  XNOR U808 ( .A(n754), .B(n752), .Z(n751) );
  XNOR U809 ( .A(n753), .B(n751), .Z(n757) );
  XNOR U810 ( .A(n758), .B(n757), .Z(N75) );
  NANDN U811 ( .A(n756), .B(n755), .Z(n760) );
  NAND U812 ( .A(n758), .B(n757), .Z(n759) );
  NAND U813 ( .A(n760), .B(n759), .Z(n767) );
  XNOR U814 ( .A(n768), .B(n767), .Z(n770) );
  NAND U815 ( .A(x[35]), .B(y[192]), .Z(n775) );
  AND U816 ( .A(n761), .B(o[34]), .Z(n776) );
  AND U817 ( .A(x[32]), .B(y[195]), .Z(n774) );
  XNOR U818 ( .A(n776), .B(n774), .Z(n762) );
  XNOR U819 ( .A(n775), .B(n762), .Z(n766) );
  NAND U820 ( .A(x[34]), .B(y[193]), .Z(n777) );
  XNOR U821 ( .A(o[35]), .B(n777), .Z(n765) );
  NAND U822 ( .A(x[33]), .B(y[194]), .Z(n764) );
  XOR U823 ( .A(n765), .B(n764), .Z(n763) );
  XNOR U824 ( .A(n766), .B(n763), .Z(n769) );
  XNOR U825 ( .A(n770), .B(n769), .Z(N76) );
  NANDN U826 ( .A(n768), .B(n767), .Z(n772) );
  NAND U827 ( .A(n770), .B(n769), .Z(n771) );
  NAND U828 ( .A(n772), .B(n771), .Z(n783) );
  XNOR U829 ( .A(n784), .B(n783), .Z(n786) );
  NAND U830 ( .A(x[34]), .B(y[194]), .Z(n792) );
  NAND U831 ( .A(x[35]), .B(y[193]), .Z(n795) );
  XNOR U832 ( .A(o[36]), .B(n795), .Z(n794) );
  AND U833 ( .A(x[33]), .B(y[195]), .Z(n793) );
  XNOR U834 ( .A(n794), .B(n793), .Z(n773) );
  XNOR U835 ( .A(n792), .B(n773), .Z(n780) );
  NAND U836 ( .A(x[36]), .B(y[192]), .Z(n790) );
  ANDN U837 ( .B(o[35]), .A(n777), .Z(n789) );
  NAND U838 ( .A(x[32]), .B(y[196]), .Z(n791) );
  XOR U839 ( .A(n789), .B(n791), .Z(n778) );
  XOR U840 ( .A(n790), .B(n778), .Z(n781) );
  XNOR U841 ( .A(n782), .B(n781), .Z(n779) );
  XNOR U842 ( .A(n780), .B(n779), .Z(n785) );
  XNOR U843 ( .A(n786), .B(n785), .Z(N77) );
  NANDN U844 ( .A(n784), .B(n783), .Z(n788) );
  NAND U845 ( .A(n786), .B(n785), .Z(n787) );
  NAND U846 ( .A(n788), .B(n787), .Z(n799) );
  XNOR U847 ( .A(n800), .B(n799), .Z(n802) );
  XNOR U848 ( .A(n805), .B(n806), .Z(n808) );
  NAND U849 ( .A(x[37]), .B(y[192]), .Z(n820) );
  ANDN U850 ( .B(o[36]), .A(n795), .Z(n821) );
  AND U851 ( .A(x[32]), .B(y[197]), .Z(n819) );
  XNOR U852 ( .A(n821), .B(n819), .Z(n796) );
  XOR U853 ( .A(n820), .B(n796), .Z(n813) );
  NAND U854 ( .A(x[33]), .B(y[196]), .Z(n814) );
  NAND U855 ( .A(x[36]), .B(y[193]), .Z(n817) );
  XNOR U856 ( .A(o[37]), .B(n817), .Z(n816) );
  AND U857 ( .A(x[35]), .B(y[194]), .Z(n815) );
  XNOR U858 ( .A(n816), .B(n815), .Z(n797) );
  XOR U859 ( .A(n814), .B(n797), .Z(n812) );
  NAND U860 ( .A(x[34]), .B(y[195]), .Z(n811) );
  XOR U861 ( .A(n812), .B(n811), .Z(n798) );
  XOR U862 ( .A(n813), .B(n798), .Z(n807) );
  XOR U863 ( .A(n808), .B(n807), .Z(n801) );
  XNOR U864 ( .A(n802), .B(n801), .Z(N78) );
  NANDN U865 ( .A(n800), .B(n799), .Z(n804) );
  NAND U866 ( .A(n802), .B(n801), .Z(n803) );
  NAND U867 ( .A(n804), .B(n803), .Z(n868) );
  NANDN U868 ( .A(n806), .B(n805), .Z(n810) );
  NAND U869 ( .A(n808), .B(n807), .Z(n809) );
  NAND U870 ( .A(n810), .B(n809), .Z(n867) );
  XOR U871 ( .A(n862), .B(n861), .Z(n860) );
  NAND U872 ( .A(x[38]), .B(y[192]), .Z(n849) );
  ANDN U873 ( .B(o[37]), .A(n817), .Z(n848) );
  NAND U874 ( .A(x[32]), .B(y[198]), .Z(n851) );
  XOR U875 ( .A(n848), .B(n851), .Z(n818) );
  XNOR U876 ( .A(n849), .B(n818), .Z(n823) );
  AND U877 ( .A(x[34]), .B(y[196]), .Z(n829) );
  AND U878 ( .A(x[35]), .B(y[195]), .Z(n828) );
  XOR U879 ( .A(n829), .B(n828), .Z(n826) );
  AND U880 ( .A(x[37]), .B(y[193]), .Z(n830) );
  XOR U881 ( .A(n830), .B(o[38]), .Z(n854) );
  NAND U882 ( .A(x[33]), .B(y[197]), .Z(n857) );
  AND U883 ( .A(x[36]), .B(y[194]), .Z(n855) );
  XNOR U884 ( .A(n825), .B(n824), .Z(n822) );
  XOR U885 ( .A(n823), .B(n822), .Z(n859) );
  XNOR U886 ( .A(n860), .B(n859), .Z(n865) );
  XNOR U887 ( .A(n866), .B(n865), .Z(N79) );
  AND U888 ( .A(y[199]), .B(x[32]), .Z(n839) );
  AND U889 ( .A(n830), .B(o[38]), .Z(n837) );
  AND U890 ( .A(y[195]), .B(x[36]), .Z(n835) );
  AND U891 ( .A(y[196]), .B(x[35]), .Z(n832) );
  NAND U892 ( .A(y[197]), .B(x[34]), .Z(n831) );
  XNOR U893 ( .A(n832), .B(n831), .Z(n833) );
  XNOR U894 ( .A(o[39]), .B(n833), .Z(n834) );
  XNOR U895 ( .A(n835), .B(n834), .Z(n836) );
  XNOR U896 ( .A(n837), .B(n836), .Z(n838) );
  XNOR U897 ( .A(n839), .B(n838), .Z(n847) );
  AND U898 ( .A(y[193]), .B(x[38]), .Z(n841) );
  NAND U899 ( .A(y[194]), .B(x[37]), .Z(n840) );
  XNOR U900 ( .A(n841), .B(n840), .Z(n845) );
  AND U901 ( .A(y[192]), .B(x[39]), .Z(n843) );
  NAND U902 ( .A(y[198]), .B(x[33]), .Z(n842) );
  XNOR U903 ( .A(n843), .B(n842), .Z(n844) );
  XNOR U904 ( .A(n845), .B(n844), .Z(n846) );
  NANDN U905 ( .A(n849), .B(n848), .Z(n853) );
  ANDN U906 ( .B(n849), .A(n848), .Z(n850) );
  OR U907 ( .A(n851), .B(n850), .Z(n852) );
  NOR U908 ( .A(n855), .B(n854), .Z(n856) );
  OR U909 ( .A(n857), .B(n856), .Z(n858) );
  OR U910 ( .A(n862), .B(n861), .Z(n863) );
  NAND U911 ( .A(n866), .B(n865), .Z(n870) );
  NAND U912 ( .A(n868), .B(n867), .Z(n869) );
endmodule

